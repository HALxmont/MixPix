magic
tech sky130B
magscale 1 2
timestamp 1667844642
<< nwell >>
rect 1066 56837 68854 57403
rect 1066 55749 68854 56315
rect 1066 54661 68854 55227
rect 1066 53573 68854 54139
rect 1066 52485 68854 53051
rect 1066 51397 68854 51963
rect 1066 50309 68854 50875
rect 1066 49221 68854 49787
rect 1066 48133 68854 48699
rect 1066 47045 68854 47611
rect 1066 45957 68854 46523
rect 1066 44869 68854 45435
rect 1066 43781 68854 44347
rect 1066 42693 68854 43259
rect 1066 41605 68854 42171
rect 1066 40517 68854 41083
rect 1066 39429 68854 39995
rect 1066 38341 68854 38907
rect 1066 37253 68854 37819
rect 1066 36165 68854 36731
rect 1066 35077 68854 35643
rect 1066 33989 68854 34555
rect 1066 32901 68854 33467
rect 1066 31813 68854 32379
rect 1066 30725 68854 31291
rect 1066 29637 68854 30203
rect 1066 28549 68854 29115
rect 1066 27461 68854 28027
rect 1066 26373 68854 26939
rect 1066 25285 68854 25851
rect 1066 24197 68854 24763
rect 1066 23109 68854 23675
rect 1066 22021 68854 22587
rect 1066 20933 68854 21499
rect 1066 19845 68854 20411
rect 1066 18757 68854 19323
rect 1066 17669 68854 18235
rect 1066 16581 68854 17147
rect 1066 15493 68854 16059
rect 1066 14405 68854 14971
rect 1066 13317 68854 13883
rect 1066 12229 68854 12795
rect 1066 11141 68854 11707
rect 1066 10053 68854 10619
rect 1066 8965 68854 9531
rect 1066 7877 68854 8443
rect 1066 6789 68854 7355
rect 1066 5701 68854 6267
rect 1066 4613 68854 5179
rect 1066 3525 68854 4091
rect 1066 2437 68854 3003
<< obsli1 >>
rect 1104 2159 68816 57681
<< obsm1 >>
rect 1104 1640 68816 57712
<< metal2 >>
rect 3514 59200 3570 60000
rect 4066 59200 4122 60000
rect 4618 59200 4674 60000
rect 5170 59200 5226 60000
rect 5722 59200 5778 60000
rect 6274 59200 6330 60000
rect 6826 59200 6882 60000
rect 7378 59200 7434 60000
rect 7930 59200 7986 60000
rect 8482 59200 8538 60000
rect 9034 59200 9090 60000
rect 9586 59200 9642 60000
rect 10138 59200 10194 60000
rect 10690 59200 10746 60000
rect 11242 59200 11298 60000
rect 11794 59200 11850 60000
rect 12346 59200 12402 60000
rect 12898 59200 12954 60000
rect 13450 59200 13506 60000
rect 14002 59200 14058 60000
rect 14554 59200 14610 60000
rect 15106 59200 15162 60000
rect 15658 59200 15714 60000
rect 16210 59200 16266 60000
rect 16762 59200 16818 60000
rect 17314 59200 17370 60000
rect 17866 59200 17922 60000
rect 18418 59200 18474 60000
rect 18970 59200 19026 60000
rect 19522 59200 19578 60000
rect 20074 59200 20130 60000
rect 20626 59200 20682 60000
rect 21178 59200 21234 60000
rect 21730 59200 21786 60000
rect 22282 59200 22338 60000
rect 22834 59200 22890 60000
rect 23386 59200 23442 60000
rect 23938 59200 23994 60000
rect 24490 59200 24546 60000
rect 25042 59200 25098 60000
rect 25594 59200 25650 60000
rect 26146 59200 26202 60000
rect 26698 59200 26754 60000
rect 27250 59200 27306 60000
rect 27802 59200 27858 60000
rect 28354 59200 28410 60000
rect 28906 59200 28962 60000
rect 29458 59200 29514 60000
rect 30010 59200 30066 60000
rect 30562 59200 30618 60000
rect 31114 59200 31170 60000
rect 31666 59200 31722 60000
rect 32218 59200 32274 60000
rect 32770 59200 32826 60000
rect 33322 59200 33378 60000
rect 33874 59200 33930 60000
rect 34426 59200 34482 60000
rect 34978 59200 35034 60000
rect 35530 59200 35586 60000
rect 36082 59200 36138 60000
rect 36634 59200 36690 60000
rect 37186 59200 37242 60000
rect 37738 59200 37794 60000
rect 38290 59200 38346 60000
rect 38842 59200 38898 60000
rect 39394 59200 39450 60000
rect 39946 59200 40002 60000
rect 40498 59200 40554 60000
rect 41050 59200 41106 60000
rect 41602 59200 41658 60000
rect 42154 59200 42210 60000
rect 42706 59200 42762 60000
rect 43258 59200 43314 60000
rect 43810 59200 43866 60000
rect 44362 59200 44418 60000
rect 44914 59200 44970 60000
rect 45466 59200 45522 60000
rect 46018 59200 46074 60000
rect 46570 59200 46626 60000
rect 47122 59200 47178 60000
rect 47674 59200 47730 60000
rect 48226 59200 48282 60000
rect 48778 59200 48834 60000
rect 49330 59200 49386 60000
rect 49882 59200 49938 60000
rect 50434 59200 50490 60000
rect 50986 59200 51042 60000
rect 51538 59200 51594 60000
rect 52090 59200 52146 60000
rect 52642 59200 52698 60000
rect 53194 59200 53250 60000
rect 53746 59200 53802 60000
rect 54298 59200 54354 60000
rect 54850 59200 54906 60000
rect 55402 59200 55458 60000
rect 55954 59200 56010 60000
rect 56506 59200 56562 60000
rect 57058 59200 57114 60000
rect 57610 59200 57666 60000
rect 58162 59200 58218 60000
rect 58714 59200 58770 60000
rect 59266 59200 59322 60000
rect 59818 59200 59874 60000
rect 60370 59200 60426 60000
rect 60922 59200 60978 60000
rect 61474 59200 61530 60000
rect 62026 59200 62082 60000
rect 62578 59200 62634 60000
rect 63130 59200 63186 60000
rect 63682 59200 63738 60000
rect 64234 59200 64290 60000
rect 64786 59200 64842 60000
rect 65338 59200 65394 60000
rect 65890 59200 65946 60000
rect 66442 59200 66498 60000
rect 12346 0 12402 800
rect 12438 0 12494 800
rect 12530 0 12586 800
rect 12622 0 12678 800
rect 12714 0 12770 800
rect 12806 0 12862 800
rect 12898 0 12954 800
rect 12990 0 13046 800
rect 13082 0 13138 800
rect 13174 0 13230 800
rect 13266 0 13322 800
rect 13358 0 13414 800
rect 13450 0 13506 800
rect 13542 0 13598 800
rect 13634 0 13690 800
rect 13726 0 13782 800
rect 13818 0 13874 800
rect 13910 0 13966 800
rect 14002 0 14058 800
rect 14094 0 14150 800
rect 14186 0 14242 800
rect 14278 0 14334 800
rect 14370 0 14426 800
rect 14462 0 14518 800
rect 14554 0 14610 800
rect 14646 0 14702 800
rect 14738 0 14794 800
rect 14830 0 14886 800
rect 14922 0 14978 800
rect 15014 0 15070 800
rect 15106 0 15162 800
rect 15198 0 15254 800
rect 15290 0 15346 800
rect 15382 0 15438 800
rect 15474 0 15530 800
rect 15566 0 15622 800
rect 15658 0 15714 800
rect 15750 0 15806 800
rect 15842 0 15898 800
rect 15934 0 15990 800
rect 16026 0 16082 800
rect 16118 0 16174 800
rect 16210 0 16266 800
rect 16302 0 16358 800
rect 16394 0 16450 800
rect 16486 0 16542 800
rect 16578 0 16634 800
rect 16670 0 16726 800
rect 16762 0 16818 800
rect 16854 0 16910 800
rect 16946 0 17002 800
rect 17038 0 17094 800
rect 17130 0 17186 800
rect 17222 0 17278 800
rect 17314 0 17370 800
rect 17406 0 17462 800
rect 17498 0 17554 800
rect 17590 0 17646 800
rect 17682 0 17738 800
rect 17774 0 17830 800
rect 17866 0 17922 800
rect 17958 0 18014 800
rect 18050 0 18106 800
rect 18142 0 18198 800
rect 18234 0 18290 800
rect 18326 0 18382 800
rect 18418 0 18474 800
rect 18510 0 18566 800
rect 18602 0 18658 800
rect 18694 0 18750 800
rect 18786 0 18842 800
rect 18878 0 18934 800
rect 18970 0 19026 800
rect 19062 0 19118 800
rect 19154 0 19210 800
rect 19246 0 19302 800
rect 19338 0 19394 800
rect 19430 0 19486 800
rect 19522 0 19578 800
rect 19614 0 19670 800
rect 19706 0 19762 800
rect 19798 0 19854 800
rect 19890 0 19946 800
rect 19982 0 20038 800
rect 20074 0 20130 800
rect 20166 0 20222 800
rect 20258 0 20314 800
rect 20350 0 20406 800
rect 20442 0 20498 800
rect 20534 0 20590 800
rect 20626 0 20682 800
rect 20718 0 20774 800
rect 20810 0 20866 800
rect 20902 0 20958 800
rect 20994 0 21050 800
rect 21086 0 21142 800
rect 21178 0 21234 800
rect 21270 0 21326 800
rect 21362 0 21418 800
rect 21454 0 21510 800
rect 21546 0 21602 800
rect 21638 0 21694 800
rect 21730 0 21786 800
rect 21822 0 21878 800
rect 21914 0 21970 800
rect 22006 0 22062 800
rect 22098 0 22154 800
rect 22190 0 22246 800
rect 22282 0 22338 800
rect 22374 0 22430 800
rect 22466 0 22522 800
rect 22558 0 22614 800
rect 22650 0 22706 800
rect 22742 0 22798 800
rect 22834 0 22890 800
rect 22926 0 22982 800
rect 23018 0 23074 800
rect 23110 0 23166 800
rect 23202 0 23258 800
rect 23294 0 23350 800
rect 23386 0 23442 800
rect 23478 0 23534 800
rect 23570 0 23626 800
rect 23662 0 23718 800
rect 23754 0 23810 800
rect 23846 0 23902 800
rect 23938 0 23994 800
rect 24030 0 24086 800
rect 24122 0 24178 800
rect 24214 0 24270 800
rect 24306 0 24362 800
rect 24398 0 24454 800
rect 24490 0 24546 800
rect 24582 0 24638 800
rect 24674 0 24730 800
rect 24766 0 24822 800
rect 24858 0 24914 800
rect 24950 0 25006 800
rect 25042 0 25098 800
rect 25134 0 25190 800
rect 25226 0 25282 800
rect 25318 0 25374 800
rect 25410 0 25466 800
rect 25502 0 25558 800
rect 25594 0 25650 800
rect 25686 0 25742 800
rect 25778 0 25834 800
rect 25870 0 25926 800
rect 25962 0 26018 800
rect 26054 0 26110 800
rect 26146 0 26202 800
rect 26238 0 26294 800
rect 26330 0 26386 800
rect 26422 0 26478 800
rect 26514 0 26570 800
rect 26606 0 26662 800
rect 26698 0 26754 800
rect 26790 0 26846 800
rect 26882 0 26938 800
rect 26974 0 27030 800
rect 27066 0 27122 800
rect 27158 0 27214 800
rect 27250 0 27306 800
rect 27342 0 27398 800
rect 27434 0 27490 800
rect 27526 0 27582 800
rect 27618 0 27674 800
rect 27710 0 27766 800
rect 27802 0 27858 800
rect 27894 0 27950 800
rect 27986 0 28042 800
rect 28078 0 28134 800
rect 28170 0 28226 800
rect 28262 0 28318 800
rect 28354 0 28410 800
rect 28446 0 28502 800
rect 28538 0 28594 800
rect 28630 0 28686 800
rect 28722 0 28778 800
rect 28814 0 28870 800
rect 28906 0 28962 800
rect 28998 0 29054 800
rect 29090 0 29146 800
rect 29182 0 29238 800
rect 29274 0 29330 800
rect 29366 0 29422 800
rect 29458 0 29514 800
rect 29550 0 29606 800
rect 29642 0 29698 800
rect 29734 0 29790 800
rect 29826 0 29882 800
rect 29918 0 29974 800
rect 30010 0 30066 800
rect 30102 0 30158 800
rect 30194 0 30250 800
rect 30286 0 30342 800
rect 30378 0 30434 800
rect 30470 0 30526 800
rect 30562 0 30618 800
rect 30654 0 30710 800
rect 30746 0 30802 800
rect 30838 0 30894 800
rect 30930 0 30986 800
rect 31022 0 31078 800
rect 31114 0 31170 800
rect 31206 0 31262 800
rect 31298 0 31354 800
rect 31390 0 31446 800
rect 31482 0 31538 800
rect 31574 0 31630 800
rect 31666 0 31722 800
rect 31758 0 31814 800
rect 31850 0 31906 800
rect 31942 0 31998 800
rect 32034 0 32090 800
rect 32126 0 32182 800
rect 32218 0 32274 800
rect 32310 0 32366 800
rect 32402 0 32458 800
rect 32494 0 32550 800
rect 32586 0 32642 800
rect 32678 0 32734 800
rect 32770 0 32826 800
rect 32862 0 32918 800
rect 32954 0 33010 800
rect 33046 0 33102 800
rect 33138 0 33194 800
rect 33230 0 33286 800
rect 33322 0 33378 800
rect 33414 0 33470 800
rect 33506 0 33562 800
rect 33598 0 33654 800
rect 33690 0 33746 800
rect 33782 0 33838 800
rect 33874 0 33930 800
rect 33966 0 34022 800
rect 34058 0 34114 800
rect 34150 0 34206 800
rect 34242 0 34298 800
rect 34334 0 34390 800
rect 34426 0 34482 800
rect 34518 0 34574 800
rect 34610 0 34666 800
rect 34702 0 34758 800
rect 34794 0 34850 800
rect 34886 0 34942 800
rect 34978 0 35034 800
rect 35070 0 35126 800
rect 35162 0 35218 800
rect 35254 0 35310 800
rect 35346 0 35402 800
rect 35438 0 35494 800
rect 35530 0 35586 800
rect 35622 0 35678 800
rect 35714 0 35770 800
rect 35806 0 35862 800
rect 35898 0 35954 800
rect 35990 0 36046 800
rect 36082 0 36138 800
rect 36174 0 36230 800
rect 36266 0 36322 800
rect 36358 0 36414 800
rect 36450 0 36506 800
rect 36542 0 36598 800
rect 36634 0 36690 800
rect 36726 0 36782 800
rect 36818 0 36874 800
rect 36910 0 36966 800
rect 37002 0 37058 800
rect 37094 0 37150 800
rect 37186 0 37242 800
rect 37278 0 37334 800
rect 37370 0 37426 800
rect 37462 0 37518 800
rect 37554 0 37610 800
rect 37646 0 37702 800
rect 37738 0 37794 800
rect 37830 0 37886 800
rect 37922 0 37978 800
rect 38014 0 38070 800
rect 38106 0 38162 800
rect 38198 0 38254 800
rect 38290 0 38346 800
rect 38382 0 38438 800
rect 38474 0 38530 800
rect 38566 0 38622 800
rect 38658 0 38714 800
rect 38750 0 38806 800
rect 38842 0 38898 800
rect 38934 0 38990 800
rect 39026 0 39082 800
rect 39118 0 39174 800
rect 39210 0 39266 800
rect 39302 0 39358 800
rect 39394 0 39450 800
rect 39486 0 39542 800
rect 39578 0 39634 800
rect 39670 0 39726 800
rect 39762 0 39818 800
rect 39854 0 39910 800
rect 39946 0 40002 800
rect 40038 0 40094 800
rect 40130 0 40186 800
rect 40222 0 40278 800
rect 40314 0 40370 800
rect 40406 0 40462 800
rect 40498 0 40554 800
rect 40590 0 40646 800
rect 40682 0 40738 800
rect 40774 0 40830 800
rect 40866 0 40922 800
rect 40958 0 41014 800
rect 41050 0 41106 800
rect 41142 0 41198 800
rect 41234 0 41290 800
rect 41326 0 41382 800
rect 41418 0 41474 800
rect 41510 0 41566 800
rect 41602 0 41658 800
rect 41694 0 41750 800
rect 41786 0 41842 800
rect 41878 0 41934 800
rect 41970 0 42026 800
rect 42062 0 42118 800
rect 42154 0 42210 800
rect 42246 0 42302 800
rect 42338 0 42394 800
rect 42430 0 42486 800
rect 42522 0 42578 800
rect 42614 0 42670 800
rect 42706 0 42762 800
rect 42798 0 42854 800
rect 42890 0 42946 800
rect 42982 0 43038 800
rect 43074 0 43130 800
rect 43166 0 43222 800
rect 43258 0 43314 800
rect 43350 0 43406 800
rect 43442 0 43498 800
rect 43534 0 43590 800
rect 43626 0 43682 800
rect 43718 0 43774 800
rect 43810 0 43866 800
rect 43902 0 43958 800
rect 43994 0 44050 800
rect 44086 0 44142 800
rect 44178 0 44234 800
rect 44270 0 44326 800
rect 44362 0 44418 800
rect 44454 0 44510 800
rect 44546 0 44602 800
rect 44638 0 44694 800
rect 44730 0 44786 800
rect 44822 0 44878 800
rect 44914 0 44970 800
rect 45006 0 45062 800
rect 45098 0 45154 800
rect 45190 0 45246 800
rect 45282 0 45338 800
rect 45374 0 45430 800
rect 45466 0 45522 800
rect 45558 0 45614 800
rect 45650 0 45706 800
rect 45742 0 45798 800
rect 45834 0 45890 800
rect 45926 0 45982 800
rect 46018 0 46074 800
rect 46110 0 46166 800
rect 46202 0 46258 800
rect 46294 0 46350 800
rect 46386 0 46442 800
rect 46478 0 46534 800
rect 46570 0 46626 800
rect 46662 0 46718 800
rect 46754 0 46810 800
rect 46846 0 46902 800
rect 46938 0 46994 800
rect 47030 0 47086 800
rect 47122 0 47178 800
rect 47214 0 47270 800
rect 47306 0 47362 800
rect 47398 0 47454 800
rect 47490 0 47546 800
rect 47582 0 47638 800
rect 47674 0 47730 800
rect 47766 0 47822 800
rect 47858 0 47914 800
rect 47950 0 48006 800
rect 48042 0 48098 800
rect 48134 0 48190 800
rect 48226 0 48282 800
rect 48318 0 48374 800
rect 48410 0 48466 800
rect 48502 0 48558 800
rect 48594 0 48650 800
rect 48686 0 48742 800
rect 48778 0 48834 800
rect 48870 0 48926 800
rect 48962 0 49018 800
rect 49054 0 49110 800
rect 49146 0 49202 800
rect 49238 0 49294 800
rect 49330 0 49386 800
rect 49422 0 49478 800
rect 49514 0 49570 800
rect 49606 0 49662 800
rect 49698 0 49754 800
rect 49790 0 49846 800
rect 49882 0 49938 800
rect 49974 0 50030 800
rect 50066 0 50122 800
rect 50158 0 50214 800
rect 50250 0 50306 800
rect 50342 0 50398 800
rect 50434 0 50490 800
rect 50526 0 50582 800
rect 50618 0 50674 800
rect 50710 0 50766 800
rect 50802 0 50858 800
rect 50894 0 50950 800
rect 50986 0 51042 800
rect 51078 0 51134 800
rect 51170 0 51226 800
rect 51262 0 51318 800
rect 51354 0 51410 800
rect 51446 0 51502 800
rect 51538 0 51594 800
rect 51630 0 51686 800
rect 51722 0 51778 800
rect 51814 0 51870 800
rect 51906 0 51962 800
rect 51998 0 52054 800
rect 52090 0 52146 800
rect 52182 0 52238 800
rect 52274 0 52330 800
rect 52366 0 52422 800
rect 52458 0 52514 800
rect 52550 0 52606 800
rect 52642 0 52698 800
rect 52734 0 52790 800
rect 52826 0 52882 800
rect 52918 0 52974 800
rect 53010 0 53066 800
rect 53102 0 53158 800
rect 53194 0 53250 800
rect 53286 0 53342 800
rect 53378 0 53434 800
rect 53470 0 53526 800
rect 53562 0 53618 800
rect 53654 0 53710 800
rect 53746 0 53802 800
rect 53838 0 53894 800
rect 53930 0 53986 800
rect 54022 0 54078 800
rect 54114 0 54170 800
rect 54206 0 54262 800
rect 54298 0 54354 800
rect 54390 0 54446 800
rect 54482 0 54538 800
rect 54574 0 54630 800
rect 54666 0 54722 800
rect 54758 0 54814 800
rect 54850 0 54906 800
rect 54942 0 54998 800
rect 55034 0 55090 800
rect 55126 0 55182 800
rect 55218 0 55274 800
rect 55310 0 55366 800
rect 55402 0 55458 800
rect 55494 0 55550 800
rect 55586 0 55642 800
rect 55678 0 55734 800
rect 55770 0 55826 800
rect 55862 0 55918 800
rect 55954 0 56010 800
rect 56046 0 56102 800
rect 56138 0 56194 800
rect 56230 0 56286 800
rect 56322 0 56378 800
rect 56414 0 56470 800
rect 56506 0 56562 800
rect 56598 0 56654 800
rect 56690 0 56746 800
rect 56782 0 56838 800
rect 56874 0 56930 800
rect 56966 0 57022 800
rect 57058 0 57114 800
rect 57150 0 57206 800
rect 57242 0 57298 800
rect 57334 0 57390 800
rect 57426 0 57482 800
rect 57518 0 57574 800
rect 57610 0 57666 800
<< obsm2 >>
rect 2596 59144 3458 59242
rect 3626 59144 4010 59242
rect 4178 59144 4562 59242
rect 4730 59144 5114 59242
rect 5282 59144 5666 59242
rect 5834 59144 6218 59242
rect 6386 59144 6770 59242
rect 6938 59144 7322 59242
rect 7490 59144 7874 59242
rect 8042 59144 8426 59242
rect 8594 59144 8978 59242
rect 9146 59144 9530 59242
rect 9698 59144 10082 59242
rect 10250 59144 10634 59242
rect 10802 59144 11186 59242
rect 11354 59144 11738 59242
rect 11906 59144 12290 59242
rect 12458 59144 12842 59242
rect 13010 59144 13394 59242
rect 13562 59144 13946 59242
rect 14114 59144 14498 59242
rect 14666 59144 15050 59242
rect 15218 59144 15602 59242
rect 15770 59144 16154 59242
rect 16322 59144 16706 59242
rect 16874 59144 17258 59242
rect 17426 59144 17810 59242
rect 17978 59144 18362 59242
rect 18530 59144 18914 59242
rect 19082 59144 19466 59242
rect 19634 59144 20018 59242
rect 20186 59144 20570 59242
rect 20738 59144 21122 59242
rect 21290 59144 21674 59242
rect 21842 59144 22226 59242
rect 22394 59144 22778 59242
rect 22946 59144 23330 59242
rect 23498 59144 23882 59242
rect 24050 59144 24434 59242
rect 24602 59144 24986 59242
rect 25154 59144 25538 59242
rect 25706 59144 26090 59242
rect 26258 59144 26642 59242
rect 26810 59144 27194 59242
rect 27362 59144 27746 59242
rect 27914 59144 28298 59242
rect 28466 59144 28850 59242
rect 29018 59144 29402 59242
rect 29570 59144 29954 59242
rect 30122 59144 30506 59242
rect 30674 59144 31058 59242
rect 31226 59144 31610 59242
rect 31778 59144 32162 59242
rect 32330 59144 32714 59242
rect 32882 59144 33266 59242
rect 33434 59144 33818 59242
rect 33986 59144 34370 59242
rect 34538 59144 34922 59242
rect 35090 59144 35474 59242
rect 35642 59144 36026 59242
rect 36194 59144 36578 59242
rect 36746 59144 37130 59242
rect 37298 59144 37682 59242
rect 37850 59144 38234 59242
rect 38402 59144 38786 59242
rect 38954 59144 39338 59242
rect 39506 59144 39890 59242
rect 40058 59144 40442 59242
rect 40610 59144 40994 59242
rect 41162 59144 41546 59242
rect 41714 59144 42098 59242
rect 42266 59144 42650 59242
rect 42818 59144 43202 59242
rect 43370 59144 43754 59242
rect 43922 59144 44306 59242
rect 44474 59144 44858 59242
rect 45026 59144 45410 59242
rect 45578 59144 45962 59242
rect 46130 59144 46514 59242
rect 46682 59144 47066 59242
rect 47234 59144 47618 59242
rect 47786 59144 48170 59242
rect 48338 59144 48722 59242
rect 48890 59144 49274 59242
rect 49442 59144 49826 59242
rect 49994 59144 50378 59242
rect 50546 59144 50930 59242
rect 51098 59144 51482 59242
rect 51650 59144 52034 59242
rect 52202 59144 52586 59242
rect 52754 59144 53138 59242
rect 53306 59144 53690 59242
rect 53858 59144 54242 59242
rect 54410 59144 54794 59242
rect 54962 59144 55346 59242
rect 55514 59144 55898 59242
rect 56066 59144 56450 59242
rect 56618 59144 57002 59242
rect 57170 59144 57554 59242
rect 57722 59144 58106 59242
rect 58274 59144 58658 59242
rect 58826 59144 59210 59242
rect 59378 59144 59762 59242
rect 59930 59144 60314 59242
rect 60482 59144 60866 59242
rect 61034 59144 61418 59242
rect 61586 59144 61970 59242
rect 62138 59144 62522 59242
rect 62690 59144 63074 59242
rect 63242 59144 63626 59242
rect 63794 59144 64178 59242
rect 64346 59144 64730 59242
rect 64898 59144 65282 59242
rect 65450 59144 65834 59242
rect 66002 59144 66386 59242
rect 2596 856 66496 59144
rect 2596 734 12290 856
rect 57722 734 66496 856
<< obsm3 >>
rect 3233 2075 65966 57697
<< metal4 >>
rect 4208 2128 4528 57712
rect 19568 2128 19888 57712
rect 34928 2128 35248 57712
rect 50288 2128 50608 57712
rect 65648 2128 65968 57712
<< obsm4 >>
rect 13675 2755 13741 6085
<< labels >>
rlabel metal2 s 3514 59200 3570 60000 6 io_in[0]
port 1 nsew signal input
rlabel metal2 s 20074 59200 20130 60000 6 io_in[10]
port 2 nsew signal input
rlabel metal2 s 21730 59200 21786 60000 6 io_in[11]
port 3 nsew signal input
rlabel metal2 s 23386 59200 23442 60000 6 io_in[12]
port 4 nsew signal input
rlabel metal2 s 25042 59200 25098 60000 6 io_in[13]
port 5 nsew signal input
rlabel metal2 s 26698 59200 26754 60000 6 io_in[14]
port 6 nsew signal input
rlabel metal2 s 28354 59200 28410 60000 6 io_in[15]
port 7 nsew signal input
rlabel metal2 s 30010 59200 30066 60000 6 io_in[16]
port 8 nsew signal input
rlabel metal2 s 31666 59200 31722 60000 6 io_in[17]
port 9 nsew signal input
rlabel metal2 s 33322 59200 33378 60000 6 io_in[18]
port 10 nsew signal input
rlabel metal2 s 34978 59200 35034 60000 6 io_in[19]
port 11 nsew signal input
rlabel metal2 s 5170 59200 5226 60000 6 io_in[1]
port 12 nsew signal input
rlabel metal2 s 36634 59200 36690 60000 6 io_in[20]
port 13 nsew signal input
rlabel metal2 s 38290 59200 38346 60000 6 io_in[21]
port 14 nsew signal input
rlabel metal2 s 39946 59200 40002 60000 6 io_in[22]
port 15 nsew signal input
rlabel metal2 s 41602 59200 41658 60000 6 io_in[23]
port 16 nsew signal input
rlabel metal2 s 43258 59200 43314 60000 6 io_in[24]
port 17 nsew signal input
rlabel metal2 s 44914 59200 44970 60000 6 io_in[25]
port 18 nsew signal input
rlabel metal2 s 46570 59200 46626 60000 6 io_in[26]
port 19 nsew signal input
rlabel metal2 s 48226 59200 48282 60000 6 io_in[27]
port 20 nsew signal input
rlabel metal2 s 49882 59200 49938 60000 6 io_in[28]
port 21 nsew signal input
rlabel metal2 s 51538 59200 51594 60000 6 io_in[29]
port 22 nsew signal input
rlabel metal2 s 6826 59200 6882 60000 6 io_in[2]
port 23 nsew signal input
rlabel metal2 s 53194 59200 53250 60000 6 io_in[30]
port 24 nsew signal input
rlabel metal2 s 54850 59200 54906 60000 6 io_in[31]
port 25 nsew signal input
rlabel metal2 s 56506 59200 56562 60000 6 io_in[32]
port 26 nsew signal input
rlabel metal2 s 58162 59200 58218 60000 6 io_in[33]
port 27 nsew signal input
rlabel metal2 s 59818 59200 59874 60000 6 io_in[34]
port 28 nsew signal input
rlabel metal2 s 61474 59200 61530 60000 6 io_in[35]
port 29 nsew signal input
rlabel metal2 s 63130 59200 63186 60000 6 io_in[36]
port 30 nsew signal input
rlabel metal2 s 64786 59200 64842 60000 6 io_in[37]
port 31 nsew signal input
rlabel metal2 s 8482 59200 8538 60000 6 io_in[3]
port 32 nsew signal input
rlabel metal2 s 10138 59200 10194 60000 6 io_in[4]
port 33 nsew signal input
rlabel metal2 s 11794 59200 11850 60000 6 io_in[5]
port 34 nsew signal input
rlabel metal2 s 13450 59200 13506 60000 6 io_in[6]
port 35 nsew signal input
rlabel metal2 s 15106 59200 15162 60000 6 io_in[7]
port 36 nsew signal input
rlabel metal2 s 16762 59200 16818 60000 6 io_in[8]
port 37 nsew signal input
rlabel metal2 s 18418 59200 18474 60000 6 io_in[9]
port 38 nsew signal input
rlabel metal2 s 4066 59200 4122 60000 6 io_oeb[0]
port 39 nsew signal output
rlabel metal2 s 20626 59200 20682 60000 6 io_oeb[10]
port 40 nsew signal output
rlabel metal2 s 22282 59200 22338 60000 6 io_oeb[11]
port 41 nsew signal output
rlabel metal2 s 23938 59200 23994 60000 6 io_oeb[12]
port 42 nsew signal output
rlabel metal2 s 25594 59200 25650 60000 6 io_oeb[13]
port 43 nsew signal output
rlabel metal2 s 27250 59200 27306 60000 6 io_oeb[14]
port 44 nsew signal output
rlabel metal2 s 28906 59200 28962 60000 6 io_oeb[15]
port 45 nsew signal output
rlabel metal2 s 30562 59200 30618 60000 6 io_oeb[16]
port 46 nsew signal output
rlabel metal2 s 32218 59200 32274 60000 6 io_oeb[17]
port 47 nsew signal output
rlabel metal2 s 33874 59200 33930 60000 6 io_oeb[18]
port 48 nsew signal output
rlabel metal2 s 35530 59200 35586 60000 6 io_oeb[19]
port 49 nsew signal output
rlabel metal2 s 5722 59200 5778 60000 6 io_oeb[1]
port 50 nsew signal output
rlabel metal2 s 37186 59200 37242 60000 6 io_oeb[20]
port 51 nsew signal output
rlabel metal2 s 38842 59200 38898 60000 6 io_oeb[21]
port 52 nsew signal output
rlabel metal2 s 40498 59200 40554 60000 6 io_oeb[22]
port 53 nsew signal output
rlabel metal2 s 42154 59200 42210 60000 6 io_oeb[23]
port 54 nsew signal output
rlabel metal2 s 43810 59200 43866 60000 6 io_oeb[24]
port 55 nsew signal output
rlabel metal2 s 45466 59200 45522 60000 6 io_oeb[25]
port 56 nsew signal output
rlabel metal2 s 47122 59200 47178 60000 6 io_oeb[26]
port 57 nsew signal output
rlabel metal2 s 48778 59200 48834 60000 6 io_oeb[27]
port 58 nsew signal output
rlabel metal2 s 50434 59200 50490 60000 6 io_oeb[28]
port 59 nsew signal output
rlabel metal2 s 52090 59200 52146 60000 6 io_oeb[29]
port 60 nsew signal output
rlabel metal2 s 7378 59200 7434 60000 6 io_oeb[2]
port 61 nsew signal output
rlabel metal2 s 53746 59200 53802 60000 6 io_oeb[30]
port 62 nsew signal output
rlabel metal2 s 55402 59200 55458 60000 6 io_oeb[31]
port 63 nsew signal output
rlabel metal2 s 57058 59200 57114 60000 6 io_oeb[32]
port 64 nsew signal output
rlabel metal2 s 58714 59200 58770 60000 6 io_oeb[33]
port 65 nsew signal output
rlabel metal2 s 60370 59200 60426 60000 6 io_oeb[34]
port 66 nsew signal output
rlabel metal2 s 62026 59200 62082 60000 6 io_oeb[35]
port 67 nsew signal output
rlabel metal2 s 63682 59200 63738 60000 6 io_oeb[36]
port 68 nsew signal output
rlabel metal2 s 65338 59200 65394 60000 6 io_oeb[37]
port 69 nsew signal output
rlabel metal2 s 9034 59200 9090 60000 6 io_oeb[3]
port 70 nsew signal output
rlabel metal2 s 10690 59200 10746 60000 6 io_oeb[4]
port 71 nsew signal output
rlabel metal2 s 12346 59200 12402 60000 6 io_oeb[5]
port 72 nsew signal output
rlabel metal2 s 14002 59200 14058 60000 6 io_oeb[6]
port 73 nsew signal output
rlabel metal2 s 15658 59200 15714 60000 6 io_oeb[7]
port 74 nsew signal output
rlabel metal2 s 17314 59200 17370 60000 6 io_oeb[8]
port 75 nsew signal output
rlabel metal2 s 18970 59200 19026 60000 6 io_oeb[9]
port 76 nsew signal output
rlabel metal2 s 4618 59200 4674 60000 6 io_out[0]
port 77 nsew signal output
rlabel metal2 s 21178 59200 21234 60000 6 io_out[10]
port 78 nsew signal output
rlabel metal2 s 22834 59200 22890 60000 6 io_out[11]
port 79 nsew signal output
rlabel metal2 s 24490 59200 24546 60000 6 io_out[12]
port 80 nsew signal output
rlabel metal2 s 26146 59200 26202 60000 6 io_out[13]
port 81 nsew signal output
rlabel metal2 s 27802 59200 27858 60000 6 io_out[14]
port 82 nsew signal output
rlabel metal2 s 29458 59200 29514 60000 6 io_out[15]
port 83 nsew signal output
rlabel metal2 s 31114 59200 31170 60000 6 io_out[16]
port 84 nsew signal output
rlabel metal2 s 32770 59200 32826 60000 6 io_out[17]
port 85 nsew signal output
rlabel metal2 s 34426 59200 34482 60000 6 io_out[18]
port 86 nsew signal output
rlabel metal2 s 36082 59200 36138 60000 6 io_out[19]
port 87 nsew signal output
rlabel metal2 s 6274 59200 6330 60000 6 io_out[1]
port 88 nsew signal output
rlabel metal2 s 37738 59200 37794 60000 6 io_out[20]
port 89 nsew signal output
rlabel metal2 s 39394 59200 39450 60000 6 io_out[21]
port 90 nsew signal output
rlabel metal2 s 41050 59200 41106 60000 6 io_out[22]
port 91 nsew signal output
rlabel metal2 s 42706 59200 42762 60000 6 io_out[23]
port 92 nsew signal output
rlabel metal2 s 44362 59200 44418 60000 6 io_out[24]
port 93 nsew signal output
rlabel metal2 s 46018 59200 46074 60000 6 io_out[25]
port 94 nsew signal output
rlabel metal2 s 47674 59200 47730 60000 6 io_out[26]
port 95 nsew signal output
rlabel metal2 s 49330 59200 49386 60000 6 io_out[27]
port 96 nsew signal output
rlabel metal2 s 50986 59200 51042 60000 6 io_out[28]
port 97 nsew signal output
rlabel metal2 s 52642 59200 52698 60000 6 io_out[29]
port 98 nsew signal output
rlabel metal2 s 7930 59200 7986 60000 6 io_out[2]
port 99 nsew signal output
rlabel metal2 s 54298 59200 54354 60000 6 io_out[30]
port 100 nsew signal output
rlabel metal2 s 55954 59200 56010 60000 6 io_out[31]
port 101 nsew signal output
rlabel metal2 s 57610 59200 57666 60000 6 io_out[32]
port 102 nsew signal output
rlabel metal2 s 59266 59200 59322 60000 6 io_out[33]
port 103 nsew signal output
rlabel metal2 s 60922 59200 60978 60000 6 io_out[34]
port 104 nsew signal output
rlabel metal2 s 62578 59200 62634 60000 6 io_out[35]
port 105 nsew signal output
rlabel metal2 s 64234 59200 64290 60000 6 io_out[36]
port 106 nsew signal output
rlabel metal2 s 65890 59200 65946 60000 6 io_out[37]
port 107 nsew signal output
rlabel metal2 s 9586 59200 9642 60000 6 io_out[3]
port 108 nsew signal output
rlabel metal2 s 11242 59200 11298 60000 6 io_out[4]
port 109 nsew signal output
rlabel metal2 s 12898 59200 12954 60000 6 io_out[5]
port 110 nsew signal output
rlabel metal2 s 14554 59200 14610 60000 6 io_out[6]
port 111 nsew signal output
rlabel metal2 s 16210 59200 16266 60000 6 io_out[7]
port 112 nsew signal output
rlabel metal2 s 17866 59200 17922 60000 6 io_out[8]
port 113 nsew signal output
rlabel metal2 s 19522 59200 19578 60000 6 io_out[9]
port 114 nsew signal output
rlabel metal2 s 57426 0 57482 800 6 irq[0]
port 115 nsew signal output
rlabel metal2 s 57518 0 57574 800 6 irq[1]
port 116 nsew signal output
rlabel metal2 s 57610 0 57666 800 6 irq[2]
port 117 nsew signal output
rlabel metal2 s 22098 0 22154 800 6 la_data_in[0]
port 118 nsew signal input
rlabel metal2 s 49698 0 49754 800 6 la_data_in[100]
port 119 nsew signal input
rlabel metal2 s 49974 0 50030 800 6 la_data_in[101]
port 120 nsew signal input
rlabel metal2 s 50250 0 50306 800 6 la_data_in[102]
port 121 nsew signal input
rlabel metal2 s 50526 0 50582 800 6 la_data_in[103]
port 122 nsew signal input
rlabel metal2 s 50802 0 50858 800 6 la_data_in[104]
port 123 nsew signal input
rlabel metal2 s 51078 0 51134 800 6 la_data_in[105]
port 124 nsew signal input
rlabel metal2 s 51354 0 51410 800 6 la_data_in[106]
port 125 nsew signal input
rlabel metal2 s 51630 0 51686 800 6 la_data_in[107]
port 126 nsew signal input
rlabel metal2 s 51906 0 51962 800 6 la_data_in[108]
port 127 nsew signal input
rlabel metal2 s 52182 0 52238 800 6 la_data_in[109]
port 128 nsew signal input
rlabel metal2 s 24858 0 24914 800 6 la_data_in[10]
port 129 nsew signal input
rlabel metal2 s 52458 0 52514 800 6 la_data_in[110]
port 130 nsew signal input
rlabel metal2 s 52734 0 52790 800 6 la_data_in[111]
port 131 nsew signal input
rlabel metal2 s 53010 0 53066 800 6 la_data_in[112]
port 132 nsew signal input
rlabel metal2 s 53286 0 53342 800 6 la_data_in[113]
port 133 nsew signal input
rlabel metal2 s 53562 0 53618 800 6 la_data_in[114]
port 134 nsew signal input
rlabel metal2 s 53838 0 53894 800 6 la_data_in[115]
port 135 nsew signal input
rlabel metal2 s 54114 0 54170 800 6 la_data_in[116]
port 136 nsew signal input
rlabel metal2 s 54390 0 54446 800 6 la_data_in[117]
port 137 nsew signal input
rlabel metal2 s 54666 0 54722 800 6 la_data_in[118]
port 138 nsew signal input
rlabel metal2 s 54942 0 54998 800 6 la_data_in[119]
port 139 nsew signal input
rlabel metal2 s 25134 0 25190 800 6 la_data_in[11]
port 140 nsew signal input
rlabel metal2 s 55218 0 55274 800 6 la_data_in[120]
port 141 nsew signal input
rlabel metal2 s 55494 0 55550 800 6 la_data_in[121]
port 142 nsew signal input
rlabel metal2 s 55770 0 55826 800 6 la_data_in[122]
port 143 nsew signal input
rlabel metal2 s 56046 0 56102 800 6 la_data_in[123]
port 144 nsew signal input
rlabel metal2 s 56322 0 56378 800 6 la_data_in[124]
port 145 nsew signal input
rlabel metal2 s 56598 0 56654 800 6 la_data_in[125]
port 146 nsew signal input
rlabel metal2 s 56874 0 56930 800 6 la_data_in[126]
port 147 nsew signal input
rlabel metal2 s 57150 0 57206 800 6 la_data_in[127]
port 148 nsew signal input
rlabel metal2 s 25410 0 25466 800 6 la_data_in[12]
port 149 nsew signal input
rlabel metal2 s 25686 0 25742 800 6 la_data_in[13]
port 150 nsew signal input
rlabel metal2 s 25962 0 26018 800 6 la_data_in[14]
port 151 nsew signal input
rlabel metal2 s 26238 0 26294 800 6 la_data_in[15]
port 152 nsew signal input
rlabel metal2 s 26514 0 26570 800 6 la_data_in[16]
port 153 nsew signal input
rlabel metal2 s 26790 0 26846 800 6 la_data_in[17]
port 154 nsew signal input
rlabel metal2 s 27066 0 27122 800 6 la_data_in[18]
port 155 nsew signal input
rlabel metal2 s 27342 0 27398 800 6 la_data_in[19]
port 156 nsew signal input
rlabel metal2 s 22374 0 22430 800 6 la_data_in[1]
port 157 nsew signal input
rlabel metal2 s 27618 0 27674 800 6 la_data_in[20]
port 158 nsew signal input
rlabel metal2 s 27894 0 27950 800 6 la_data_in[21]
port 159 nsew signal input
rlabel metal2 s 28170 0 28226 800 6 la_data_in[22]
port 160 nsew signal input
rlabel metal2 s 28446 0 28502 800 6 la_data_in[23]
port 161 nsew signal input
rlabel metal2 s 28722 0 28778 800 6 la_data_in[24]
port 162 nsew signal input
rlabel metal2 s 28998 0 29054 800 6 la_data_in[25]
port 163 nsew signal input
rlabel metal2 s 29274 0 29330 800 6 la_data_in[26]
port 164 nsew signal input
rlabel metal2 s 29550 0 29606 800 6 la_data_in[27]
port 165 nsew signal input
rlabel metal2 s 29826 0 29882 800 6 la_data_in[28]
port 166 nsew signal input
rlabel metal2 s 30102 0 30158 800 6 la_data_in[29]
port 167 nsew signal input
rlabel metal2 s 22650 0 22706 800 6 la_data_in[2]
port 168 nsew signal input
rlabel metal2 s 30378 0 30434 800 6 la_data_in[30]
port 169 nsew signal input
rlabel metal2 s 30654 0 30710 800 6 la_data_in[31]
port 170 nsew signal input
rlabel metal2 s 30930 0 30986 800 6 la_data_in[32]
port 171 nsew signal input
rlabel metal2 s 31206 0 31262 800 6 la_data_in[33]
port 172 nsew signal input
rlabel metal2 s 31482 0 31538 800 6 la_data_in[34]
port 173 nsew signal input
rlabel metal2 s 31758 0 31814 800 6 la_data_in[35]
port 174 nsew signal input
rlabel metal2 s 32034 0 32090 800 6 la_data_in[36]
port 175 nsew signal input
rlabel metal2 s 32310 0 32366 800 6 la_data_in[37]
port 176 nsew signal input
rlabel metal2 s 32586 0 32642 800 6 la_data_in[38]
port 177 nsew signal input
rlabel metal2 s 32862 0 32918 800 6 la_data_in[39]
port 178 nsew signal input
rlabel metal2 s 22926 0 22982 800 6 la_data_in[3]
port 179 nsew signal input
rlabel metal2 s 33138 0 33194 800 6 la_data_in[40]
port 180 nsew signal input
rlabel metal2 s 33414 0 33470 800 6 la_data_in[41]
port 181 nsew signal input
rlabel metal2 s 33690 0 33746 800 6 la_data_in[42]
port 182 nsew signal input
rlabel metal2 s 33966 0 34022 800 6 la_data_in[43]
port 183 nsew signal input
rlabel metal2 s 34242 0 34298 800 6 la_data_in[44]
port 184 nsew signal input
rlabel metal2 s 34518 0 34574 800 6 la_data_in[45]
port 185 nsew signal input
rlabel metal2 s 34794 0 34850 800 6 la_data_in[46]
port 186 nsew signal input
rlabel metal2 s 35070 0 35126 800 6 la_data_in[47]
port 187 nsew signal input
rlabel metal2 s 35346 0 35402 800 6 la_data_in[48]
port 188 nsew signal input
rlabel metal2 s 35622 0 35678 800 6 la_data_in[49]
port 189 nsew signal input
rlabel metal2 s 23202 0 23258 800 6 la_data_in[4]
port 190 nsew signal input
rlabel metal2 s 35898 0 35954 800 6 la_data_in[50]
port 191 nsew signal input
rlabel metal2 s 36174 0 36230 800 6 la_data_in[51]
port 192 nsew signal input
rlabel metal2 s 36450 0 36506 800 6 la_data_in[52]
port 193 nsew signal input
rlabel metal2 s 36726 0 36782 800 6 la_data_in[53]
port 194 nsew signal input
rlabel metal2 s 37002 0 37058 800 6 la_data_in[54]
port 195 nsew signal input
rlabel metal2 s 37278 0 37334 800 6 la_data_in[55]
port 196 nsew signal input
rlabel metal2 s 37554 0 37610 800 6 la_data_in[56]
port 197 nsew signal input
rlabel metal2 s 37830 0 37886 800 6 la_data_in[57]
port 198 nsew signal input
rlabel metal2 s 38106 0 38162 800 6 la_data_in[58]
port 199 nsew signal input
rlabel metal2 s 38382 0 38438 800 6 la_data_in[59]
port 200 nsew signal input
rlabel metal2 s 23478 0 23534 800 6 la_data_in[5]
port 201 nsew signal input
rlabel metal2 s 38658 0 38714 800 6 la_data_in[60]
port 202 nsew signal input
rlabel metal2 s 38934 0 38990 800 6 la_data_in[61]
port 203 nsew signal input
rlabel metal2 s 39210 0 39266 800 6 la_data_in[62]
port 204 nsew signal input
rlabel metal2 s 39486 0 39542 800 6 la_data_in[63]
port 205 nsew signal input
rlabel metal2 s 39762 0 39818 800 6 la_data_in[64]
port 206 nsew signal input
rlabel metal2 s 40038 0 40094 800 6 la_data_in[65]
port 207 nsew signal input
rlabel metal2 s 40314 0 40370 800 6 la_data_in[66]
port 208 nsew signal input
rlabel metal2 s 40590 0 40646 800 6 la_data_in[67]
port 209 nsew signal input
rlabel metal2 s 40866 0 40922 800 6 la_data_in[68]
port 210 nsew signal input
rlabel metal2 s 41142 0 41198 800 6 la_data_in[69]
port 211 nsew signal input
rlabel metal2 s 23754 0 23810 800 6 la_data_in[6]
port 212 nsew signal input
rlabel metal2 s 41418 0 41474 800 6 la_data_in[70]
port 213 nsew signal input
rlabel metal2 s 41694 0 41750 800 6 la_data_in[71]
port 214 nsew signal input
rlabel metal2 s 41970 0 42026 800 6 la_data_in[72]
port 215 nsew signal input
rlabel metal2 s 42246 0 42302 800 6 la_data_in[73]
port 216 nsew signal input
rlabel metal2 s 42522 0 42578 800 6 la_data_in[74]
port 217 nsew signal input
rlabel metal2 s 42798 0 42854 800 6 la_data_in[75]
port 218 nsew signal input
rlabel metal2 s 43074 0 43130 800 6 la_data_in[76]
port 219 nsew signal input
rlabel metal2 s 43350 0 43406 800 6 la_data_in[77]
port 220 nsew signal input
rlabel metal2 s 43626 0 43682 800 6 la_data_in[78]
port 221 nsew signal input
rlabel metal2 s 43902 0 43958 800 6 la_data_in[79]
port 222 nsew signal input
rlabel metal2 s 24030 0 24086 800 6 la_data_in[7]
port 223 nsew signal input
rlabel metal2 s 44178 0 44234 800 6 la_data_in[80]
port 224 nsew signal input
rlabel metal2 s 44454 0 44510 800 6 la_data_in[81]
port 225 nsew signal input
rlabel metal2 s 44730 0 44786 800 6 la_data_in[82]
port 226 nsew signal input
rlabel metal2 s 45006 0 45062 800 6 la_data_in[83]
port 227 nsew signal input
rlabel metal2 s 45282 0 45338 800 6 la_data_in[84]
port 228 nsew signal input
rlabel metal2 s 45558 0 45614 800 6 la_data_in[85]
port 229 nsew signal input
rlabel metal2 s 45834 0 45890 800 6 la_data_in[86]
port 230 nsew signal input
rlabel metal2 s 46110 0 46166 800 6 la_data_in[87]
port 231 nsew signal input
rlabel metal2 s 46386 0 46442 800 6 la_data_in[88]
port 232 nsew signal input
rlabel metal2 s 46662 0 46718 800 6 la_data_in[89]
port 233 nsew signal input
rlabel metal2 s 24306 0 24362 800 6 la_data_in[8]
port 234 nsew signal input
rlabel metal2 s 46938 0 46994 800 6 la_data_in[90]
port 235 nsew signal input
rlabel metal2 s 47214 0 47270 800 6 la_data_in[91]
port 236 nsew signal input
rlabel metal2 s 47490 0 47546 800 6 la_data_in[92]
port 237 nsew signal input
rlabel metal2 s 47766 0 47822 800 6 la_data_in[93]
port 238 nsew signal input
rlabel metal2 s 48042 0 48098 800 6 la_data_in[94]
port 239 nsew signal input
rlabel metal2 s 48318 0 48374 800 6 la_data_in[95]
port 240 nsew signal input
rlabel metal2 s 48594 0 48650 800 6 la_data_in[96]
port 241 nsew signal input
rlabel metal2 s 48870 0 48926 800 6 la_data_in[97]
port 242 nsew signal input
rlabel metal2 s 49146 0 49202 800 6 la_data_in[98]
port 243 nsew signal input
rlabel metal2 s 49422 0 49478 800 6 la_data_in[99]
port 244 nsew signal input
rlabel metal2 s 24582 0 24638 800 6 la_data_in[9]
port 245 nsew signal input
rlabel metal2 s 22190 0 22246 800 6 la_data_out[0]
port 246 nsew signal output
rlabel metal2 s 49790 0 49846 800 6 la_data_out[100]
port 247 nsew signal output
rlabel metal2 s 50066 0 50122 800 6 la_data_out[101]
port 248 nsew signal output
rlabel metal2 s 50342 0 50398 800 6 la_data_out[102]
port 249 nsew signal output
rlabel metal2 s 50618 0 50674 800 6 la_data_out[103]
port 250 nsew signal output
rlabel metal2 s 50894 0 50950 800 6 la_data_out[104]
port 251 nsew signal output
rlabel metal2 s 51170 0 51226 800 6 la_data_out[105]
port 252 nsew signal output
rlabel metal2 s 51446 0 51502 800 6 la_data_out[106]
port 253 nsew signal output
rlabel metal2 s 51722 0 51778 800 6 la_data_out[107]
port 254 nsew signal output
rlabel metal2 s 51998 0 52054 800 6 la_data_out[108]
port 255 nsew signal output
rlabel metal2 s 52274 0 52330 800 6 la_data_out[109]
port 256 nsew signal output
rlabel metal2 s 24950 0 25006 800 6 la_data_out[10]
port 257 nsew signal output
rlabel metal2 s 52550 0 52606 800 6 la_data_out[110]
port 258 nsew signal output
rlabel metal2 s 52826 0 52882 800 6 la_data_out[111]
port 259 nsew signal output
rlabel metal2 s 53102 0 53158 800 6 la_data_out[112]
port 260 nsew signal output
rlabel metal2 s 53378 0 53434 800 6 la_data_out[113]
port 261 nsew signal output
rlabel metal2 s 53654 0 53710 800 6 la_data_out[114]
port 262 nsew signal output
rlabel metal2 s 53930 0 53986 800 6 la_data_out[115]
port 263 nsew signal output
rlabel metal2 s 54206 0 54262 800 6 la_data_out[116]
port 264 nsew signal output
rlabel metal2 s 54482 0 54538 800 6 la_data_out[117]
port 265 nsew signal output
rlabel metal2 s 54758 0 54814 800 6 la_data_out[118]
port 266 nsew signal output
rlabel metal2 s 55034 0 55090 800 6 la_data_out[119]
port 267 nsew signal output
rlabel metal2 s 25226 0 25282 800 6 la_data_out[11]
port 268 nsew signal output
rlabel metal2 s 55310 0 55366 800 6 la_data_out[120]
port 269 nsew signal output
rlabel metal2 s 55586 0 55642 800 6 la_data_out[121]
port 270 nsew signal output
rlabel metal2 s 55862 0 55918 800 6 la_data_out[122]
port 271 nsew signal output
rlabel metal2 s 56138 0 56194 800 6 la_data_out[123]
port 272 nsew signal output
rlabel metal2 s 56414 0 56470 800 6 la_data_out[124]
port 273 nsew signal output
rlabel metal2 s 56690 0 56746 800 6 la_data_out[125]
port 274 nsew signal output
rlabel metal2 s 56966 0 57022 800 6 la_data_out[126]
port 275 nsew signal output
rlabel metal2 s 57242 0 57298 800 6 la_data_out[127]
port 276 nsew signal output
rlabel metal2 s 25502 0 25558 800 6 la_data_out[12]
port 277 nsew signal output
rlabel metal2 s 25778 0 25834 800 6 la_data_out[13]
port 278 nsew signal output
rlabel metal2 s 26054 0 26110 800 6 la_data_out[14]
port 279 nsew signal output
rlabel metal2 s 26330 0 26386 800 6 la_data_out[15]
port 280 nsew signal output
rlabel metal2 s 26606 0 26662 800 6 la_data_out[16]
port 281 nsew signal output
rlabel metal2 s 26882 0 26938 800 6 la_data_out[17]
port 282 nsew signal output
rlabel metal2 s 27158 0 27214 800 6 la_data_out[18]
port 283 nsew signal output
rlabel metal2 s 27434 0 27490 800 6 la_data_out[19]
port 284 nsew signal output
rlabel metal2 s 22466 0 22522 800 6 la_data_out[1]
port 285 nsew signal output
rlabel metal2 s 27710 0 27766 800 6 la_data_out[20]
port 286 nsew signal output
rlabel metal2 s 27986 0 28042 800 6 la_data_out[21]
port 287 nsew signal output
rlabel metal2 s 28262 0 28318 800 6 la_data_out[22]
port 288 nsew signal output
rlabel metal2 s 28538 0 28594 800 6 la_data_out[23]
port 289 nsew signal output
rlabel metal2 s 28814 0 28870 800 6 la_data_out[24]
port 290 nsew signal output
rlabel metal2 s 29090 0 29146 800 6 la_data_out[25]
port 291 nsew signal output
rlabel metal2 s 29366 0 29422 800 6 la_data_out[26]
port 292 nsew signal output
rlabel metal2 s 29642 0 29698 800 6 la_data_out[27]
port 293 nsew signal output
rlabel metal2 s 29918 0 29974 800 6 la_data_out[28]
port 294 nsew signal output
rlabel metal2 s 30194 0 30250 800 6 la_data_out[29]
port 295 nsew signal output
rlabel metal2 s 22742 0 22798 800 6 la_data_out[2]
port 296 nsew signal output
rlabel metal2 s 30470 0 30526 800 6 la_data_out[30]
port 297 nsew signal output
rlabel metal2 s 30746 0 30802 800 6 la_data_out[31]
port 298 nsew signal output
rlabel metal2 s 31022 0 31078 800 6 la_data_out[32]
port 299 nsew signal output
rlabel metal2 s 31298 0 31354 800 6 la_data_out[33]
port 300 nsew signal output
rlabel metal2 s 31574 0 31630 800 6 la_data_out[34]
port 301 nsew signal output
rlabel metal2 s 31850 0 31906 800 6 la_data_out[35]
port 302 nsew signal output
rlabel metal2 s 32126 0 32182 800 6 la_data_out[36]
port 303 nsew signal output
rlabel metal2 s 32402 0 32458 800 6 la_data_out[37]
port 304 nsew signal output
rlabel metal2 s 32678 0 32734 800 6 la_data_out[38]
port 305 nsew signal output
rlabel metal2 s 32954 0 33010 800 6 la_data_out[39]
port 306 nsew signal output
rlabel metal2 s 23018 0 23074 800 6 la_data_out[3]
port 307 nsew signal output
rlabel metal2 s 33230 0 33286 800 6 la_data_out[40]
port 308 nsew signal output
rlabel metal2 s 33506 0 33562 800 6 la_data_out[41]
port 309 nsew signal output
rlabel metal2 s 33782 0 33838 800 6 la_data_out[42]
port 310 nsew signal output
rlabel metal2 s 34058 0 34114 800 6 la_data_out[43]
port 311 nsew signal output
rlabel metal2 s 34334 0 34390 800 6 la_data_out[44]
port 312 nsew signal output
rlabel metal2 s 34610 0 34666 800 6 la_data_out[45]
port 313 nsew signal output
rlabel metal2 s 34886 0 34942 800 6 la_data_out[46]
port 314 nsew signal output
rlabel metal2 s 35162 0 35218 800 6 la_data_out[47]
port 315 nsew signal output
rlabel metal2 s 35438 0 35494 800 6 la_data_out[48]
port 316 nsew signal output
rlabel metal2 s 35714 0 35770 800 6 la_data_out[49]
port 317 nsew signal output
rlabel metal2 s 23294 0 23350 800 6 la_data_out[4]
port 318 nsew signal output
rlabel metal2 s 35990 0 36046 800 6 la_data_out[50]
port 319 nsew signal output
rlabel metal2 s 36266 0 36322 800 6 la_data_out[51]
port 320 nsew signal output
rlabel metal2 s 36542 0 36598 800 6 la_data_out[52]
port 321 nsew signal output
rlabel metal2 s 36818 0 36874 800 6 la_data_out[53]
port 322 nsew signal output
rlabel metal2 s 37094 0 37150 800 6 la_data_out[54]
port 323 nsew signal output
rlabel metal2 s 37370 0 37426 800 6 la_data_out[55]
port 324 nsew signal output
rlabel metal2 s 37646 0 37702 800 6 la_data_out[56]
port 325 nsew signal output
rlabel metal2 s 37922 0 37978 800 6 la_data_out[57]
port 326 nsew signal output
rlabel metal2 s 38198 0 38254 800 6 la_data_out[58]
port 327 nsew signal output
rlabel metal2 s 38474 0 38530 800 6 la_data_out[59]
port 328 nsew signal output
rlabel metal2 s 23570 0 23626 800 6 la_data_out[5]
port 329 nsew signal output
rlabel metal2 s 38750 0 38806 800 6 la_data_out[60]
port 330 nsew signal output
rlabel metal2 s 39026 0 39082 800 6 la_data_out[61]
port 331 nsew signal output
rlabel metal2 s 39302 0 39358 800 6 la_data_out[62]
port 332 nsew signal output
rlabel metal2 s 39578 0 39634 800 6 la_data_out[63]
port 333 nsew signal output
rlabel metal2 s 39854 0 39910 800 6 la_data_out[64]
port 334 nsew signal output
rlabel metal2 s 40130 0 40186 800 6 la_data_out[65]
port 335 nsew signal output
rlabel metal2 s 40406 0 40462 800 6 la_data_out[66]
port 336 nsew signal output
rlabel metal2 s 40682 0 40738 800 6 la_data_out[67]
port 337 nsew signal output
rlabel metal2 s 40958 0 41014 800 6 la_data_out[68]
port 338 nsew signal output
rlabel metal2 s 41234 0 41290 800 6 la_data_out[69]
port 339 nsew signal output
rlabel metal2 s 23846 0 23902 800 6 la_data_out[6]
port 340 nsew signal output
rlabel metal2 s 41510 0 41566 800 6 la_data_out[70]
port 341 nsew signal output
rlabel metal2 s 41786 0 41842 800 6 la_data_out[71]
port 342 nsew signal output
rlabel metal2 s 42062 0 42118 800 6 la_data_out[72]
port 343 nsew signal output
rlabel metal2 s 42338 0 42394 800 6 la_data_out[73]
port 344 nsew signal output
rlabel metal2 s 42614 0 42670 800 6 la_data_out[74]
port 345 nsew signal output
rlabel metal2 s 42890 0 42946 800 6 la_data_out[75]
port 346 nsew signal output
rlabel metal2 s 43166 0 43222 800 6 la_data_out[76]
port 347 nsew signal output
rlabel metal2 s 43442 0 43498 800 6 la_data_out[77]
port 348 nsew signal output
rlabel metal2 s 43718 0 43774 800 6 la_data_out[78]
port 349 nsew signal output
rlabel metal2 s 43994 0 44050 800 6 la_data_out[79]
port 350 nsew signal output
rlabel metal2 s 24122 0 24178 800 6 la_data_out[7]
port 351 nsew signal output
rlabel metal2 s 44270 0 44326 800 6 la_data_out[80]
port 352 nsew signal output
rlabel metal2 s 44546 0 44602 800 6 la_data_out[81]
port 353 nsew signal output
rlabel metal2 s 44822 0 44878 800 6 la_data_out[82]
port 354 nsew signal output
rlabel metal2 s 45098 0 45154 800 6 la_data_out[83]
port 355 nsew signal output
rlabel metal2 s 45374 0 45430 800 6 la_data_out[84]
port 356 nsew signal output
rlabel metal2 s 45650 0 45706 800 6 la_data_out[85]
port 357 nsew signal output
rlabel metal2 s 45926 0 45982 800 6 la_data_out[86]
port 358 nsew signal output
rlabel metal2 s 46202 0 46258 800 6 la_data_out[87]
port 359 nsew signal output
rlabel metal2 s 46478 0 46534 800 6 la_data_out[88]
port 360 nsew signal output
rlabel metal2 s 46754 0 46810 800 6 la_data_out[89]
port 361 nsew signal output
rlabel metal2 s 24398 0 24454 800 6 la_data_out[8]
port 362 nsew signal output
rlabel metal2 s 47030 0 47086 800 6 la_data_out[90]
port 363 nsew signal output
rlabel metal2 s 47306 0 47362 800 6 la_data_out[91]
port 364 nsew signal output
rlabel metal2 s 47582 0 47638 800 6 la_data_out[92]
port 365 nsew signal output
rlabel metal2 s 47858 0 47914 800 6 la_data_out[93]
port 366 nsew signal output
rlabel metal2 s 48134 0 48190 800 6 la_data_out[94]
port 367 nsew signal output
rlabel metal2 s 48410 0 48466 800 6 la_data_out[95]
port 368 nsew signal output
rlabel metal2 s 48686 0 48742 800 6 la_data_out[96]
port 369 nsew signal output
rlabel metal2 s 48962 0 49018 800 6 la_data_out[97]
port 370 nsew signal output
rlabel metal2 s 49238 0 49294 800 6 la_data_out[98]
port 371 nsew signal output
rlabel metal2 s 49514 0 49570 800 6 la_data_out[99]
port 372 nsew signal output
rlabel metal2 s 24674 0 24730 800 6 la_data_out[9]
port 373 nsew signal output
rlabel metal2 s 22282 0 22338 800 6 la_oenb[0]
port 374 nsew signal input
rlabel metal2 s 49882 0 49938 800 6 la_oenb[100]
port 375 nsew signal input
rlabel metal2 s 50158 0 50214 800 6 la_oenb[101]
port 376 nsew signal input
rlabel metal2 s 50434 0 50490 800 6 la_oenb[102]
port 377 nsew signal input
rlabel metal2 s 50710 0 50766 800 6 la_oenb[103]
port 378 nsew signal input
rlabel metal2 s 50986 0 51042 800 6 la_oenb[104]
port 379 nsew signal input
rlabel metal2 s 51262 0 51318 800 6 la_oenb[105]
port 380 nsew signal input
rlabel metal2 s 51538 0 51594 800 6 la_oenb[106]
port 381 nsew signal input
rlabel metal2 s 51814 0 51870 800 6 la_oenb[107]
port 382 nsew signal input
rlabel metal2 s 52090 0 52146 800 6 la_oenb[108]
port 383 nsew signal input
rlabel metal2 s 52366 0 52422 800 6 la_oenb[109]
port 384 nsew signal input
rlabel metal2 s 25042 0 25098 800 6 la_oenb[10]
port 385 nsew signal input
rlabel metal2 s 52642 0 52698 800 6 la_oenb[110]
port 386 nsew signal input
rlabel metal2 s 52918 0 52974 800 6 la_oenb[111]
port 387 nsew signal input
rlabel metal2 s 53194 0 53250 800 6 la_oenb[112]
port 388 nsew signal input
rlabel metal2 s 53470 0 53526 800 6 la_oenb[113]
port 389 nsew signal input
rlabel metal2 s 53746 0 53802 800 6 la_oenb[114]
port 390 nsew signal input
rlabel metal2 s 54022 0 54078 800 6 la_oenb[115]
port 391 nsew signal input
rlabel metal2 s 54298 0 54354 800 6 la_oenb[116]
port 392 nsew signal input
rlabel metal2 s 54574 0 54630 800 6 la_oenb[117]
port 393 nsew signal input
rlabel metal2 s 54850 0 54906 800 6 la_oenb[118]
port 394 nsew signal input
rlabel metal2 s 55126 0 55182 800 6 la_oenb[119]
port 395 nsew signal input
rlabel metal2 s 25318 0 25374 800 6 la_oenb[11]
port 396 nsew signal input
rlabel metal2 s 55402 0 55458 800 6 la_oenb[120]
port 397 nsew signal input
rlabel metal2 s 55678 0 55734 800 6 la_oenb[121]
port 398 nsew signal input
rlabel metal2 s 55954 0 56010 800 6 la_oenb[122]
port 399 nsew signal input
rlabel metal2 s 56230 0 56286 800 6 la_oenb[123]
port 400 nsew signal input
rlabel metal2 s 56506 0 56562 800 6 la_oenb[124]
port 401 nsew signal input
rlabel metal2 s 56782 0 56838 800 6 la_oenb[125]
port 402 nsew signal input
rlabel metal2 s 57058 0 57114 800 6 la_oenb[126]
port 403 nsew signal input
rlabel metal2 s 57334 0 57390 800 6 la_oenb[127]
port 404 nsew signal input
rlabel metal2 s 25594 0 25650 800 6 la_oenb[12]
port 405 nsew signal input
rlabel metal2 s 25870 0 25926 800 6 la_oenb[13]
port 406 nsew signal input
rlabel metal2 s 26146 0 26202 800 6 la_oenb[14]
port 407 nsew signal input
rlabel metal2 s 26422 0 26478 800 6 la_oenb[15]
port 408 nsew signal input
rlabel metal2 s 26698 0 26754 800 6 la_oenb[16]
port 409 nsew signal input
rlabel metal2 s 26974 0 27030 800 6 la_oenb[17]
port 410 nsew signal input
rlabel metal2 s 27250 0 27306 800 6 la_oenb[18]
port 411 nsew signal input
rlabel metal2 s 27526 0 27582 800 6 la_oenb[19]
port 412 nsew signal input
rlabel metal2 s 22558 0 22614 800 6 la_oenb[1]
port 413 nsew signal input
rlabel metal2 s 27802 0 27858 800 6 la_oenb[20]
port 414 nsew signal input
rlabel metal2 s 28078 0 28134 800 6 la_oenb[21]
port 415 nsew signal input
rlabel metal2 s 28354 0 28410 800 6 la_oenb[22]
port 416 nsew signal input
rlabel metal2 s 28630 0 28686 800 6 la_oenb[23]
port 417 nsew signal input
rlabel metal2 s 28906 0 28962 800 6 la_oenb[24]
port 418 nsew signal input
rlabel metal2 s 29182 0 29238 800 6 la_oenb[25]
port 419 nsew signal input
rlabel metal2 s 29458 0 29514 800 6 la_oenb[26]
port 420 nsew signal input
rlabel metal2 s 29734 0 29790 800 6 la_oenb[27]
port 421 nsew signal input
rlabel metal2 s 30010 0 30066 800 6 la_oenb[28]
port 422 nsew signal input
rlabel metal2 s 30286 0 30342 800 6 la_oenb[29]
port 423 nsew signal input
rlabel metal2 s 22834 0 22890 800 6 la_oenb[2]
port 424 nsew signal input
rlabel metal2 s 30562 0 30618 800 6 la_oenb[30]
port 425 nsew signal input
rlabel metal2 s 30838 0 30894 800 6 la_oenb[31]
port 426 nsew signal input
rlabel metal2 s 31114 0 31170 800 6 la_oenb[32]
port 427 nsew signal input
rlabel metal2 s 31390 0 31446 800 6 la_oenb[33]
port 428 nsew signal input
rlabel metal2 s 31666 0 31722 800 6 la_oenb[34]
port 429 nsew signal input
rlabel metal2 s 31942 0 31998 800 6 la_oenb[35]
port 430 nsew signal input
rlabel metal2 s 32218 0 32274 800 6 la_oenb[36]
port 431 nsew signal input
rlabel metal2 s 32494 0 32550 800 6 la_oenb[37]
port 432 nsew signal input
rlabel metal2 s 32770 0 32826 800 6 la_oenb[38]
port 433 nsew signal input
rlabel metal2 s 33046 0 33102 800 6 la_oenb[39]
port 434 nsew signal input
rlabel metal2 s 23110 0 23166 800 6 la_oenb[3]
port 435 nsew signal input
rlabel metal2 s 33322 0 33378 800 6 la_oenb[40]
port 436 nsew signal input
rlabel metal2 s 33598 0 33654 800 6 la_oenb[41]
port 437 nsew signal input
rlabel metal2 s 33874 0 33930 800 6 la_oenb[42]
port 438 nsew signal input
rlabel metal2 s 34150 0 34206 800 6 la_oenb[43]
port 439 nsew signal input
rlabel metal2 s 34426 0 34482 800 6 la_oenb[44]
port 440 nsew signal input
rlabel metal2 s 34702 0 34758 800 6 la_oenb[45]
port 441 nsew signal input
rlabel metal2 s 34978 0 35034 800 6 la_oenb[46]
port 442 nsew signal input
rlabel metal2 s 35254 0 35310 800 6 la_oenb[47]
port 443 nsew signal input
rlabel metal2 s 35530 0 35586 800 6 la_oenb[48]
port 444 nsew signal input
rlabel metal2 s 35806 0 35862 800 6 la_oenb[49]
port 445 nsew signal input
rlabel metal2 s 23386 0 23442 800 6 la_oenb[4]
port 446 nsew signal input
rlabel metal2 s 36082 0 36138 800 6 la_oenb[50]
port 447 nsew signal input
rlabel metal2 s 36358 0 36414 800 6 la_oenb[51]
port 448 nsew signal input
rlabel metal2 s 36634 0 36690 800 6 la_oenb[52]
port 449 nsew signal input
rlabel metal2 s 36910 0 36966 800 6 la_oenb[53]
port 450 nsew signal input
rlabel metal2 s 37186 0 37242 800 6 la_oenb[54]
port 451 nsew signal input
rlabel metal2 s 37462 0 37518 800 6 la_oenb[55]
port 452 nsew signal input
rlabel metal2 s 37738 0 37794 800 6 la_oenb[56]
port 453 nsew signal input
rlabel metal2 s 38014 0 38070 800 6 la_oenb[57]
port 454 nsew signal input
rlabel metal2 s 38290 0 38346 800 6 la_oenb[58]
port 455 nsew signal input
rlabel metal2 s 38566 0 38622 800 6 la_oenb[59]
port 456 nsew signal input
rlabel metal2 s 23662 0 23718 800 6 la_oenb[5]
port 457 nsew signal input
rlabel metal2 s 38842 0 38898 800 6 la_oenb[60]
port 458 nsew signal input
rlabel metal2 s 39118 0 39174 800 6 la_oenb[61]
port 459 nsew signal input
rlabel metal2 s 39394 0 39450 800 6 la_oenb[62]
port 460 nsew signal input
rlabel metal2 s 39670 0 39726 800 6 la_oenb[63]
port 461 nsew signal input
rlabel metal2 s 39946 0 40002 800 6 la_oenb[64]
port 462 nsew signal input
rlabel metal2 s 40222 0 40278 800 6 la_oenb[65]
port 463 nsew signal input
rlabel metal2 s 40498 0 40554 800 6 la_oenb[66]
port 464 nsew signal input
rlabel metal2 s 40774 0 40830 800 6 la_oenb[67]
port 465 nsew signal input
rlabel metal2 s 41050 0 41106 800 6 la_oenb[68]
port 466 nsew signal input
rlabel metal2 s 41326 0 41382 800 6 la_oenb[69]
port 467 nsew signal input
rlabel metal2 s 23938 0 23994 800 6 la_oenb[6]
port 468 nsew signal input
rlabel metal2 s 41602 0 41658 800 6 la_oenb[70]
port 469 nsew signal input
rlabel metal2 s 41878 0 41934 800 6 la_oenb[71]
port 470 nsew signal input
rlabel metal2 s 42154 0 42210 800 6 la_oenb[72]
port 471 nsew signal input
rlabel metal2 s 42430 0 42486 800 6 la_oenb[73]
port 472 nsew signal input
rlabel metal2 s 42706 0 42762 800 6 la_oenb[74]
port 473 nsew signal input
rlabel metal2 s 42982 0 43038 800 6 la_oenb[75]
port 474 nsew signal input
rlabel metal2 s 43258 0 43314 800 6 la_oenb[76]
port 475 nsew signal input
rlabel metal2 s 43534 0 43590 800 6 la_oenb[77]
port 476 nsew signal input
rlabel metal2 s 43810 0 43866 800 6 la_oenb[78]
port 477 nsew signal input
rlabel metal2 s 44086 0 44142 800 6 la_oenb[79]
port 478 nsew signal input
rlabel metal2 s 24214 0 24270 800 6 la_oenb[7]
port 479 nsew signal input
rlabel metal2 s 44362 0 44418 800 6 la_oenb[80]
port 480 nsew signal input
rlabel metal2 s 44638 0 44694 800 6 la_oenb[81]
port 481 nsew signal input
rlabel metal2 s 44914 0 44970 800 6 la_oenb[82]
port 482 nsew signal input
rlabel metal2 s 45190 0 45246 800 6 la_oenb[83]
port 483 nsew signal input
rlabel metal2 s 45466 0 45522 800 6 la_oenb[84]
port 484 nsew signal input
rlabel metal2 s 45742 0 45798 800 6 la_oenb[85]
port 485 nsew signal input
rlabel metal2 s 46018 0 46074 800 6 la_oenb[86]
port 486 nsew signal input
rlabel metal2 s 46294 0 46350 800 6 la_oenb[87]
port 487 nsew signal input
rlabel metal2 s 46570 0 46626 800 6 la_oenb[88]
port 488 nsew signal input
rlabel metal2 s 46846 0 46902 800 6 la_oenb[89]
port 489 nsew signal input
rlabel metal2 s 24490 0 24546 800 6 la_oenb[8]
port 490 nsew signal input
rlabel metal2 s 47122 0 47178 800 6 la_oenb[90]
port 491 nsew signal input
rlabel metal2 s 47398 0 47454 800 6 la_oenb[91]
port 492 nsew signal input
rlabel metal2 s 47674 0 47730 800 6 la_oenb[92]
port 493 nsew signal input
rlabel metal2 s 47950 0 48006 800 6 la_oenb[93]
port 494 nsew signal input
rlabel metal2 s 48226 0 48282 800 6 la_oenb[94]
port 495 nsew signal input
rlabel metal2 s 48502 0 48558 800 6 la_oenb[95]
port 496 nsew signal input
rlabel metal2 s 48778 0 48834 800 6 la_oenb[96]
port 497 nsew signal input
rlabel metal2 s 49054 0 49110 800 6 la_oenb[97]
port 498 nsew signal input
rlabel metal2 s 49330 0 49386 800 6 la_oenb[98]
port 499 nsew signal input
rlabel metal2 s 49606 0 49662 800 6 la_oenb[99]
port 500 nsew signal input
rlabel metal2 s 24766 0 24822 800 6 la_oenb[9]
port 501 nsew signal input
rlabel metal2 s 66442 59200 66498 60000 6 serial_data_rlbp_out
port 502 nsew signal output
rlabel metal4 s 4208 2128 4528 57712 6 vccd1
port 503 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 57712 6 vccd1
port 503 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 57712 6 vccd1
port 503 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 57712 6 vssd1
port 504 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 57712 6 vssd1
port 504 nsew ground bidirectional
rlabel metal2 s 12346 0 12402 800 6 wb_clk_i
port 505 nsew signal input
rlabel metal2 s 12438 0 12494 800 6 wb_rst_i
port 506 nsew signal input
rlabel metal2 s 12530 0 12586 800 6 wbs_ack_o
port 507 nsew signal output
rlabel metal2 s 12898 0 12954 800 6 wbs_adr_i[0]
port 508 nsew signal input
rlabel metal2 s 16026 0 16082 800 6 wbs_adr_i[10]
port 509 nsew signal input
rlabel metal2 s 16302 0 16358 800 6 wbs_adr_i[11]
port 510 nsew signal input
rlabel metal2 s 16578 0 16634 800 6 wbs_adr_i[12]
port 511 nsew signal input
rlabel metal2 s 16854 0 16910 800 6 wbs_adr_i[13]
port 512 nsew signal input
rlabel metal2 s 17130 0 17186 800 6 wbs_adr_i[14]
port 513 nsew signal input
rlabel metal2 s 17406 0 17462 800 6 wbs_adr_i[15]
port 514 nsew signal input
rlabel metal2 s 17682 0 17738 800 6 wbs_adr_i[16]
port 515 nsew signal input
rlabel metal2 s 17958 0 18014 800 6 wbs_adr_i[17]
port 516 nsew signal input
rlabel metal2 s 18234 0 18290 800 6 wbs_adr_i[18]
port 517 nsew signal input
rlabel metal2 s 18510 0 18566 800 6 wbs_adr_i[19]
port 518 nsew signal input
rlabel metal2 s 13266 0 13322 800 6 wbs_adr_i[1]
port 519 nsew signal input
rlabel metal2 s 18786 0 18842 800 6 wbs_adr_i[20]
port 520 nsew signal input
rlabel metal2 s 19062 0 19118 800 6 wbs_adr_i[21]
port 521 nsew signal input
rlabel metal2 s 19338 0 19394 800 6 wbs_adr_i[22]
port 522 nsew signal input
rlabel metal2 s 19614 0 19670 800 6 wbs_adr_i[23]
port 523 nsew signal input
rlabel metal2 s 19890 0 19946 800 6 wbs_adr_i[24]
port 524 nsew signal input
rlabel metal2 s 20166 0 20222 800 6 wbs_adr_i[25]
port 525 nsew signal input
rlabel metal2 s 20442 0 20498 800 6 wbs_adr_i[26]
port 526 nsew signal input
rlabel metal2 s 20718 0 20774 800 6 wbs_adr_i[27]
port 527 nsew signal input
rlabel metal2 s 20994 0 21050 800 6 wbs_adr_i[28]
port 528 nsew signal input
rlabel metal2 s 21270 0 21326 800 6 wbs_adr_i[29]
port 529 nsew signal input
rlabel metal2 s 13634 0 13690 800 6 wbs_adr_i[2]
port 530 nsew signal input
rlabel metal2 s 21546 0 21602 800 6 wbs_adr_i[30]
port 531 nsew signal input
rlabel metal2 s 21822 0 21878 800 6 wbs_adr_i[31]
port 532 nsew signal input
rlabel metal2 s 14002 0 14058 800 6 wbs_adr_i[3]
port 533 nsew signal input
rlabel metal2 s 14370 0 14426 800 6 wbs_adr_i[4]
port 534 nsew signal input
rlabel metal2 s 14646 0 14702 800 6 wbs_adr_i[5]
port 535 nsew signal input
rlabel metal2 s 14922 0 14978 800 6 wbs_adr_i[6]
port 536 nsew signal input
rlabel metal2 s 15198 0 15254 800 6 wbs_adr_i[7]
port 537 nsew signal input
rlabel metal2 s 15474 0 15530 800 6 wbs_adr_i[8]
port 538 nsew signal input
rlabel metal2 s 15750 0 15806 800 6 wbs_adr_i[9]
port 539 nsew signal input
rlabel metal2 s 12622 0 12678 800 6 wbs_cyc_i
port 540 nsew signal input
rlabel metal2 s 12990 0 13046 800 6 wbs_dat_i[0]
port 541 nsew signal input
rlabel metal2 s 16118 0 16174 800 6 wbs_dat_i[10]
port 542 nsew signal input
rlabel metal2 s 16394 0 16450 800 6 wbs_dat_i[11]
port 543 nsew signal input
rlabel metal2 s 16670 0 16726 800 6 wbs_dat_i[12]
port 544 nsew signal input
rlabel metal2 s 16946 0 17002 800 6 wbs_dat_i[13]
port 545 nsew signal input
rlabel metal2 s 17222 0 17278 800 6 wbs_dat_i[14]
port 546 nsew signal input
rlabel metal2 s 17498 0 17554 800 6 wbs_dat_i[15]
port 547 nsew signal input
rlabel metal2 s 17774 0 17830 800 6 wbs_dat_i[16]
port 548 nsew signal input
rlabel metal2 s 18050 0 18106 800 6 wbs_dat_i[17]
port 549 nsew signal input
rlabel metal2 s 18326 0 18382 800 6 wbs_dat_i[18]
port 550 nsew signal input
rlabel metal2 s 18602 0 18658 800 6 wbs_dat_i[19]
port 551 nsew signal input
rlabel metal2 s 13358 0 13414 800 6 wbs_dat_i[1]
port 552 nsew signal input
rlabel metal2 s 18878 0 18934 800 6 wbs_dat_i[20]
port 553 nsew signal input
rlabel metal2 s 19154 0 19210 800 6 wbs_dat_i[21]
port 554 nsew signal input
rlabel metal2 s 19430 0 19486 800 6 wbs_dat_i[22]
port 555 nsew signal input
rlabel metal2 s 19706 0 19762 800 6 wbs_dat_i[23]
port 556 nsew signal input
rlabel metal2 s 19982 0 20038 800 6 wbs_dat_i[24]
port 557 nsew signal input
rlabel metal2 s 20258 0 20314 800 6 wbs_dat_i[25]
port 558 nsew signal input
rlabel metal2 s 20534 0 20590 800 6 wbs_dat_i[26]
port 559 nsew signal input
rlabel metal2 s 20810 0 20866 800 6 wbs_dat_i[27]
port 560 nsew signal input
rlabel metal2 s 21086 0 21142 800 6 wbs_dat_i[28]
port 561 nsew signal input
rlabel metal2 s 21362 0 21418 800 6 wbs_dat_i[29]
port 562 nsew signal input
rlabel metal2 s 13726 0 13782 800 6 wbs_dat_i[2]
port 563 nsew signal input
rlabel metal2 s 21638 0 21694 800 6 wbs_dat_i[30]
port 564 nsew signal input
rlabel metal2 s 21914 0 21970 800 6 wbs_dat_i[31]
port 565 nsew signal input
rlabel metal2 s 14094 0 14150 800 6 wbs_dat_i[3]
port 566 nsew signal input
rlabel metal2 s 14462 0 14518 800 6 wbs_dat_i[4]
port 567 nsew signal input
rlabel metal2 s 14738 0 14794 800 6 wbs_dat_i[5]
port 568 nsew signal input
rlabel metal2 s 15014 0 15070 800 6 wbs_dat_i[6]
port 569 nsew signal input
rlabel metal2 s 15290 0 15346 800 6 wbs_dat_i[7]
port 570 nsew signal input
rlabel metal2 s 15566 0 15622 800 6 wbs_dat_i[8]
port 571 nsew signal input
rlabel metal2 s 15842 0 15898 800 6 wbs_dat_i[9]
port 572 nsew signal input
rlabel metal2 s 13082 0 13138 800 6 wbs_dat_o[0]
port 573 nsew signal output
rlabel metal2 s 16210 0 16266 800 6 wbs_dat_o[10]
port 574 nsew signal output
rlabel metal2 s 16486 0 16542 800 6 wbs_dat_o[11]
port 575 nsew signal output
rlabel metal2 s 16762 0 16818 800 6 wbs_dat_o[12]
port 576 nsew signal output
rlabel metal2 s 17038 0 17094 800 6 wbs_dat_o[13]
port 577 nsew signal output
rlabel metal2 s 17314 0 17370 800 6 wbs_dat_o[14]
port 578 nsew signal output
rlabel metal2 s 17590 0 17646 800 6 wbs_dat_o[15]
port 579 nsew signal output
rlabel metal2 s 17866 0 17922 800 6 wbs_dat_o[16]
port 580 nsew signal output
rlabel metal2 s 18142 0 18198 800 6 wbs_dat_o[17]
port 581 nsew signal output
rlabel metal2 s 18418 0 18474 800 6 wbs_dat_o[18]
port 582 nsew signal output
rlabel metal2 s 18694 0 18750 800 6 wbs_dat_o[19]
port 583 nsew signal output
rlabel metal2 s 13450 0 13506 800 6 wbs_dat_o[1]
port 584 nsew signal output
rlabel metal2 s 18970 0 19026 800 6 wbs_dat_o[20]
port 585 nsew signal output
rlabel metal2 s 19246 0 19302 800 6 wbs_dat_o[21]
port 586 nsew signal output
rlabel metal2 s 19522 0 19578 800 6 wbs_dat_o[22]
port 587 nsew signal output
rlabel metal2 s 19798 0 19854 800 6 wbs_dat_o[23]
port 588 nsew signal output
rlabel metal2 s 20074 0 20130 800 6 wbs_dat_o[24]
port 589 nsew signal output
rlabel metal2 s 20350 0 20406 800 6 wbs_dat_o[25]
port 590 nsew signal output
rlabel metal2 s 20626 0 20682 800 6 wbs_dat_o[26]
port 591 nsew signal output
rlabel metal2 s 20902 0 20958 800 6 wbs_dat_o[27]
port 592 nsew signal output
rlabel metal2 s 21178 0 21234 800 6 wbs_dat_o[28]
port 593 nsew signal output
rlabel metal2 s 21454 0 21510 800 6 wbs_dat_o[29]
port 594 nsew signal output
rlabel metal2 s 13818 0 13874 800 6 wbs_dat_o[2]
port 595 nsew signal output
rlabel metal2 s 21730 0 21786 800 6 wbs_dat_o[30]
port 596 nsew signal output
rlabel metal2 s 22006 0 22062 800 6 wbs_dat_o[31]
port 597 nsew signal output
rlabel metal2 s 14186 0 14242 800 6 wbs_dat_o[3]
port 598 nsew signal output
rlabel metal2 s 14554 0 14610 800 6 wbs_dat_o[4]
port 599 nsew signal output
rlabel metal2 s 14830 0 14886 800 6 wbs_dat_o[5]
port 600 nsew signal output
rlabel metal2 s 15106 0 15162 800 6 wbs_dat_o[6]
port 601 nsew signal output
rlabel metal2 s 15382 0 15438 800 6 wbs_dat_o[7]
port 602 nsew signal output
rlabel metal2 s 15658 0 15714 800 6 wbs_dat_o[8]
port 603 nsew signal output
rlabel metal2 s 15934 0 15990 800 6 wbs_dat_o[9]
port 604 nsew signal output
rlabel metal2 s 13174 0 13230 800 6 wbs_sel_i[0]
port 605 nsew signal input
rlabel metal2 s 13542 0 13598 800 6 wbs_sel_i[1]
port 606 nsew signal input
rlabel metal2 s 13910 0 13966 800 6 wbs_sel_i[2]
port 607 nsew signal input
rlabel metal2 s 14278 0 14334 800 6 wbs_sel_i[3]
port 608 nsew signal input
rlabel metal2 s 12714 0 12770 800 6 wbs_stb_i
port 609 nsew signal input
rlabel metal2 s 12806 0 12862 800 6 wbs_we_i
port 610 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 70000 60000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 2168612
string GDS_FILE /home/mxmont/Documents/Universidad/IC-UBB/MixPix/CARAVEL_WRAPPER/MixPix/openlane/rlbp/runs/22_11_07_15_09/results/signoff/rlbp_macro.magic.gds
string GDS_START 306578
<< end >>

