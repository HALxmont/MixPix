magic
tech sky130B
magscale 1 2
timestamp 1662509196
<< viali >>
rect 4353 17153 4387 17187
rect 4997 17153 5031 17187
rect 5825 17153 5859 17187
rect 7113 17153 7147 17187
rect 7573 17153 7607 17187
rect 8401 17153 8435 17187
rect 9137 17153 9171 17187
rect 9873 17153 9907 17187
rect 10517 17153 10551 17187
rect 11897 17153 11931 17187
rect 12633 17153 12667 17187
rect 13277 17153 13311 17187
rect 14657 17153 14691 17187
rect 15485 17153 15519 17187
rect 15945 17153 15979 17187
rect 17233 17153 17267 17187
rect 18061 17153 18095 17187
rect 18705 17153 18739 17187
rect 19533 17153 19567 17187
rect 20177 17153 20211 17187
rect 21281 17153 21315 17187
rect 22293 17153 22327 17187
rect 22937 17153 22971 17187
rect 23673 17153 23707 17187
rect 25145 17153 25179 17187
rect 25605 17153 25639 17187
rect 26433 17153 26467 17187
rect 27721 17153 27755 17187
rect 28365 17153 28399 17187
rect 29009 17153 29043 17187
rect 29837 17153 29871 17187
rect 30573 17153 30607 17187
rect 31217 17153 31251 17187
rect 32137 17153 32171 17187
rect 32781 17153 32815 17187
rect 33517 17153 33551 17187
rect 34713 17153 34747 17187
rect 35357 17153 35391 17187
rect 37289 17153 37323 17187
rect 37933 17153 37967 17187
rect 38577 17153 38611 17187
rect 39865 17153 39899 17187
rect 40509 17153 40543 17187
rect 41153 17153 41187 17187
rect 42441 17153 42475 17187
rect 43729 17153 43763 17187
rect 45017 17153 45051 17187
rect 46305 17153 46339 17187
rect 47593 17153 47627 17187
rect 48237 17153 48271 17187
rect 48881 17153 48915 17187
rect 50169 17153 50203 17187
rect 50813 17153 50847 17187
rect 51457 17153 51491 17187
rect 52745 17153 52779 17187
rect 54033 17153 54067 17187
rect 55321 17153 55355 17187
rect 55965 17153 55999 17187
rect 56609 17153 56643 17187
rect 36001 17085 36035 17119
rect 45661 17085 45695 17119
rect 43085 17017 43119 17051
rect 53389 17017 53423 17051
rect 6377 16745 6411 16779
rect 11437 16745 11471 16779
rect 14197 16745 14231 16779
rect 16957 16745 16991 16779
rect 21097 16745 21131 16779
rect 24409 16745 24443 16779
rect 27077 16745 27111 16779
rect 36277 16745 36311 16779
rect 39865 16745 39899 16779
rect 43637 16745 43671 16779
rect 46397 16745 46431 16779
rect 49157 16745 49191 16779
rect 54217 16745 54251 16779
rect 17417 13889 17451 13923
rect 3341 13821 3375 13855
rect 13369 13821 13403 13855
rect 14013 13821 14047 13855
rect 11437 13277 11471 13311
rect 6745 13209 6779 13243
rect 12633 13209 12667 13243
rect 16957 13209 16991 13243
rect 2053 13141 2087 13175
rect 2697 13141 2731 13175
rect 3249 13141 3283 13175
rect 3801 13141 3835 13175
rect 5181 13141 5215 13175
rect 6009 13141 6043 13175
rect 9413 13141 9447 13175
rect 9873 13141 9907 13175
rect 10885 13141 10919 13175
rect 11897 13141 11931 13175
rect 13185 13141 13219 13175
rect 14197 13141 14231 13175
rect 15117 13141 15151 13175
rect 15669 13141 15703 13175
rect 17785 13141 17819 13175
rect 18245 13141 18279 13175
rect 22385 13141 22419 13175
rect 9505 12937 9539 12971
rect 13001 12937 13035 12971
rect 17601 12937 17635 12971
rect 13645 12869 13679 12903
rect 21925 12869 21959 12903
rect 2513 12801 2547 12835
rect 14565 12801 14599 12835
rect 15117 12801 15151 12835
rect 19349 12801 19383 12835
rect 4169 12733 4203 12767
rect 19809 12733 19843 12767
rect 21281 12733 21315 12767
rect 4629 12665 4663 12699
rect 8401 12665 8435 12699
rect 22661 12665 22695 12699
rect 1961 12597 1995 12631
rect 3065 12597 3099 12631
rect 3617 12597 3651 12631
rect 5273 12597 5307 12631
rect 5825 12597 5859 12631
rect 6469 12597 6503 12631
rect 7021 12597 7055 12631
rect 7849 12597 7883 12631
rect 8861 12597 8895 12631
rect 10425 12597 10459 12631
rect 10977 12597 11011 12631
rect 11621 12597 11655 12631
rect 12265 12597 12299 12631
rect 16129 12597 16163 12631
rect 17141 12597 17175 12631
rect 18245 12597 18279 12631
rect 18797 12597 18831 12631
rect 20729 12597 20763 12631
rect 23489 12597 23523 12631
rect 23949 12597 23983 12631
rect 6561 12393 6595 12427
rect 9229 12393 9263 12427
rect 25145 12393 25179 12427
rect 2513 12189 2547 12223
rect 5825 12189 5859 12223
rect 18061 12189 18095 12223
rect 20361 12189 20395 12223
rect 1501 12121 1535 12155
rect 4445 12121 4479 12155
rect 7757 12121 7791 12155
rect 16313 12121 16347 12155
rect 21373 12121 21407 12155
rect 23121 12121 23155 12155
rect 1961 12053 1995 12087
rect 3157 12053 3191 12087
rect 3893 12053 3927 12087
rect 5181 12053 5215 12087
rect 7205 12053 7239 12087
rect 8401 12053 8435 12087
rect 10057 12053 10091 12087
rect 10609 12053 10643 12087
rect 11253 12053 11287 12087
rect 12081 12053 12115 12087
rect 13093 12053 13127 12087
rect 14197 12053 14231 12087
rect 15025 12053 15059 12087
rect 15669 12053 15703 12087
rect 17049 12053 17083 12087
rect 18613 12053 18647 12087
rect 19257 12053 19291 12087
rect 20913 12053 20947 12087
rect 22293 12053 22327 12087
rect 23765 12053 23799 12087
rect 24409 12053 24443 12087
rect 25605 12053 25639 12087
rect 37105 12053 37139 12087
rect 2973 11849 3007 11883
rect 6929 11849 6963 11883
rect 8677 11849 8711 11883
rect 20085 11849 20119 11883
rect 23121 11849 23155 11883
rect 26249 11645 26283 11679
rect 3525 11577 3559 11611
rect 14565 11577 14599 11611
rect 18797 11577 18831 11611
rect 23673 11577 23707 11611
rect 36461 11577 36495 11611
rect 37933 11577 37967 11611
rect 1869 11509 1903 11543
rect 4077 11509 4111 11543
rect 4905 11509 4939 11543
rect 5825 11509 5859 11543
rect 7573 11509 7607 11543
rect 8125 11509 8159 11543
rect 9321 11509 9355 11543
rect 9873 11509 9907 11543
rect 10425 11509 10459 11543
rect 10977 11509 11011 11543
rect 11805 11509 11839 11543
rect 12449 11509 12483 11543
rect 12909 11509 12943 11543
rect 13645 11509 13679 11543
rect 15117 11509 15151 11543
rect 15945 11509 15979 11543
rect 16681 11509 16715 11543
rect 17233 11509 17267 11543
rect 18245 11509 18279 11543
rect 19257 11509 19291 11543
rect 20545 11509 20579 11543
rect 21281 11509 21315 11543
rect 22109 11509 22143 11543
rect 22661 11509 22695 11543
rect 24501 11509 24535 11543
rect 25053 11509 25087 11543
rect 25605 11509 25639 11543
rect 35725 11509 35759 11543
rect 37381 11509 37415 11543
rect 38393 11509 38427 11543
rect 42901 11509 42935 11543
rect 43453 11509 43487 11543
rect 25513 11305 25547 11339
rect 35725 11305 35759 11339
rect 39865 11305 39899 11339
rect 43361 11305 43395 11339
rect 2053 11237 2087 11271
rect 5917 11237 5951 11271
rect 6929 11237 6963 11271
rect 7757 11237 7791 11271
rect 9413 11237 9447 11271
rect 11069 11237 11103 11271
rect 15669 11237 15703 11271
rect 16129 11237 16163 11271
rect 20177 11237 20211 11271
rect 24869 11237 24903 11271
rect 15025 11169 15059 11203
rect 17417 11169 17451 11203
rect 21005 11169 21039 11203
rect 3157 11101 3191 11135
rect 4813 11101 4847 11135
rect 6469 11101 6503 11135
rect 7113 11101 7147 11135
rect 7941 11101 7975 11135
rect 9597 11101 9631 11135
rect 12265 11101 12299 11135
rect 12909 11101 12943 11135
rect 13369 11101 13403 11135
rect 14105 11101 14139 11135
rect 15485 11101 15519 11135
rect 16313 11101 16347 11135
rect 16773 11101 16807 11135
rect 22201 11101 22235 11135
rect 27813 11101 27847 11135
rect 4169 11033 4203 11067
rect 10057 11033 10091 11067
rect 11529 11033 11563 11067
rect 17969 11033 18003 11067
rect 18705 11033 18739 11067
rect 19349 11033 19383 11067
rect 21465 11033 21499 11067
rect 22661 11033 22695 11067
rect 25973 11033 26007 11067
rect 26617 11033 26651 11067
rect 27261 11033 27295 11067
rect 28641 11033 28675 11067
rect 29561 11033 29595 11067
rect 35173 11033 35207 11067
rect 36185 11033 36219 11067
rect 36737 11033 36771 11067
rect 37473 11033 37507 11067
rect 39129 11033 39163 11067
rect 40417 11033 40451 11067
rect 41981 11033 42015 11067
rect 42717 11033 42751 11067
rect 43913 11033 43947 11067
rect 2605 10965 2639 10999
rect 23305 10965 23339 10999
rect 23765 10965 23799 10999
rect 38117 10965 38151 10999
rect 38577 10965 38611 10999
rect 45017 10965 45051 10999
rect 1777 10761 1811 10795
rect 3985 10761 4019 10795
rect 5825 10761 5859 10795
rect 8217 10761 8251 10795
rect 25789 10761 25823 10795
rect 36553 10761 36587 10795
rect 37933 10761 37967 10795
rect 39497 10761 39531 10795
rect 41153 10761 41187 10795
rect 41797 10761 41831 10795
rect 44465 10761 44499 10795
rect 48329 10761 48363 10795
rect 48789 10761 48823 10795
rect 46949 10693 46983 10727
rect 1593 10625 1627 10659
rect 2237 10625 2271 10659
rect 3801 10625 3835 10659
rect 4721 10625 4755 10659
rect 7113 10625 7147 10659
rect 7757 10625 7791 10659
rect 8401 10625 8435 10659
rect 8953 10625 8987 10659
rect 9413 10625 9447 10659
rect 10425 10625 10459 10659
rect 10885 10625 10919 10659
rect 11805 10625 11839 10659
rect 16129 10625 16163 10659
rect 16681 10625 16715 10659
rect 17693 10625 17727 10659
rect 19901 10625 19935 10659
rect 20085 10625 20119 10659
rect 20729 10625 20763 10659
rect 22661 10625 22695 10659
rect 23489 10625 23523 10659
rect 25605 10625 25639 10659
rect 27169 10625 27203 10659
rect 29377 10625 29411 10659
rect 47593 10625 47627 10659
rect 6469 10557 6503 10591
rect 11529 10557 11563 10591
rect 17417 10557 17451 10591
rect 19717 10557 19751 10591
rect 26249 10557 26283 10591
rect 33977 10557 34011 10591
rect 38945 10557 38979 10591
rect 7573 10489 7607 10523
rect 10241 10489 10275 10523
rect 13553 10489 13587 10523
rect 15485 10489 15519 10523
rect 19257 10489 19291 10523
rect 21189 10489 21223 10523
rect 23673 10489 23707 10523
rect 30573 10489 30607 10523
rect 38393 10489 38427 10523
rect 45293 10489 45327 10523
rect 2421 10421 2455 10455
rect 3341 10421 3375 10455
rect 4905 10421 4939 10455
rect 6929 10421 6963 10455
rect 9597 10421 9631 10455
rect 12541 10421 12575 10455
rect 14197 10421 14231 10455
rect 14841 10421 14875 10455
rect 15945 10421 15979 10455
rect 16865 10421 16899 10455
rect 18429 10421 18463 10455
rect 20545 10421 20579 10455
rect 22109 10421 22143 10455
rect 22845 10421 22879 10455
rect 24593 10421 24627 10455
rect 26985 10421 27019 10455
rect 27997 10421 28031 10455
rect 28733 10421 28767 10455
rect 29561 10421 29595 10455
rect 30113 10421 30147 10455
rect 33333 10421 33367 10455
rect 34621 10421 34655 10455
rect 35541 10421 35575 10455
rect 36093 10421 36127 10455
rect 37381 10421 37415 10455
rect 40049 10421 40083 10455
rect 40601 10421 40635 10455
rect 42533 10421 42567 10455
rect 42993 10421 43027 10455
rect 44005 10421 44039 10455
rect 45845 10421 45879 10455
rect 46397 10421 46431 10455
rect 47777 10421 47811 10455
rect 10241 10217 10275 10251
rect 16681 10217 16715 10251
rect 3157 10149 3191 10183
rect 5825 10149 5859 10183
rect 17141 10149 17175 10183
rect 35265 10149 35299 10183
rect 38853 10149 38887 10183
rect 42073 10149 42107 10183
rect 3801 10081 3835 10115
rect 6285 10081 6319 10115
rect 11989 10081 12023 10115
rect 14933 10081 14967 10115
rect 20729 10081 20763 10115
rect 22569 10081 22603 10115
rect 42717 10081 42751 10115
rect 52285 10081 52319 10115
rect 1685 10013 1719 10047
rect 2329 10013 2363 10047
rect 2973 10013 3007 10047
rect 4077 10013 4111 10047
rect 5641 10013 5675 10047
rect 6561 10013 6595 10047
rect 8401 10013 8435 10047
rect 9597 10013 9631 10047
rect 10057 10013 10091 10047
rect 10701 10013 10735 10047
rect 11345 10013 11379 10047
rect 12265 10013 12299 10047
rect 14105 10013 14139 10047
rect 15209 10013 15243 10047
rect 16497 10013 16531 10047
rect 17325 10013 17359 10047
rect 18061 10013 18095 10047
rect 18521 10013 18555 10047
rect 20453 10013 20487 10047
rect 21373 10013 21407 10047
rect 22109 10013 22143 10047
rect 22845 10013 22879 10047
rect 24409 10013 24443 10047
rect 24685 10013 24719 10047
rect 26157 10013 26191 10047
rect 26433 10013 26467 10047
rect 30849 10013 30883 10047
rect 31125 10013 31159 10047
rect 33149 10013 33183 10047
rect 33425 10013 33459 10047
rect 36277 10013 36311 10047
rect 38117 10013 38151 10047
rect 38393 10013 38427 10047
rect 42257 10013 42291 10047
rect 42993 10013 43027 10047
rect 45661 10013 45695 10047
rect 46489 10013 46523 10047
rect 46765 10013 46799 10047
rect 47409 10013 47443 10047
rect 47685 10013 47719 10047
rect 48513 10013 48547 10047
rect 49249 10013 49283 10047
rect 52561 10013 52595 10047
rect 53389 10013 53423 10047
rect 28825 9945 28859 9979
rect 41061 9945 41095 9979
rect 1869 9877 1903 9911
rect 2513 9877 2547 9911
rect 4813 9877 4847 9911
rect 7297 9877 7331 9911
rect 8217 9877 8251 9911
rect 9505 9877 9539 9911
rect 10885 9877 10919 9911
rect 11529 9877 11563 9911
rect 13001 9877 13035 9911
rect 13553 9877 13587 9911
rect 14289 9877 14323 9911
rect 15945 9877 15979 9911
rect 19717 9877 19751 9911
rect 21189 9877 21223 9911
rect 21925 9877 21959 9911
rect 23581 9877 23615 9911
rect 25421 9877 25455 9911
rect 27169 9877 27203 9911
rect 27629 9877 27663 9911
rect 28365 9877 28399 9911
rect 29561 9877 29595 9911
rect 30113 9877 30147 9911
rect 32597 9877 32631 9911
rect 34161 9877 34195 9911
rect 34805 9877 34839 9911
rect 36369 9877 36403 9911
rect 37381 9877 37415 9911
rect 39865 9877 39899 9911
rect 40417 9877 40451 9911
rect 43729 9877 43763 9911
rect 44189 9877 44223 9911
rect 45017 9877 45051 9911
rect 49065 9877 49099 9911
rect 2789 9673 2823 9707
rect 4261 9673 4295 9707
rect 6377 9673 6411 9707
rect 10517 9673 10551 9707
rect 18153 9673 18187 9707
rect 19901 9673 19935 9707
rect 22385 9673 22419 9707
rect 24225 9673 24259 9707
rect 24869 9673 24903 9707
rect 26433 9673 26467 9707
rect 27997 9673 28031 9707
rect 30941 9673 30975 9707
rect 32321 9673 32355 9707
rect 33793 9673 33827 9707
rect 34253 9673 34287 9707
rect 38393 9673 38427 9707
rect 39221 9673 39255 9707
rect 43913 9673 43947 9707
rect 46489 9673 46523 9707
rect 47777 9673 47811 9707
rect 11529 9605 11563 9639
rect 13093 9605 13127 9639
rect 14933 9605 14967 9639
rect 15761 9605 15795 9639
rect 23213 9605 23247 9639
rect 23765 9605 23799 9639
rect 37749 9605 37783 9639
rect 41613 9605 41647 9639
rect 50537 9605 50571 9639
rect 53782 9605 53816 9639
rect 1777 9537 1811 9571
rect 2513 9537 2547 9571
rect 2605 9537 2639 9571
rect 3249 9537 3283 9571
rect 3525 9537 3559 9571
rect 4997 9537 5031 9571
rect 5181 9537 5215 9571
rect 5641 9537 5675 9571
rect 6561 9537 6595 9571
rect 7849 9537 7883 9571
rect 8769 9537 8803 9571
rect 9965 9537 9999 9571
rect 10701 9537 10735 9571
rect 11713 9537 11747 9571
rect 12909 9537 12943 9571
rect 14749 9537 14783 9571
rect 15577 9537 15611 9571
rect 17141 9537 17175 9571
rect 17417 9537 17451 9571
rect 19257 9537 19291 9571
rect 20637 9537 20671 9571
rect 20913 9537 20947 9571
rect 22201 9537 22235 9571
rect 23029 9537 23063 9571
rect 24409 9537 24443 9571
rect 25053 9537 25087 9571
rect 25237 9537 25271 9571
rect 26065 9537 26099 9571
rect 26249 9537 26283 9571
rect 27261 9537 27295 9571
rect 28457 9537 28491 9571
rect 28641 9537 28675 9571
rect 29285 9537 29319 9571
rect 29561 9537 29595 9571
rect 30757 9537 30791 9571
rect 32137 9537 32171 9571
rect 33057 9537 33091 9571
rect 34989 9537 35023 9571
rect 35265 9537 35299 9571
rect 36461 9537 36495 9571
rect 36737 9537 36771 9571
rect 38577 9537 38611 9571
rect 39957 9537 39991 9571
rect 40233 9537 40267 9571
rect 41429 9537 41463 9571
rect 42717 9537 42751 9571
rect 44097 9537 44131 9571
rect 44649 9537 44683 9571
rect 45661 9537 45695 9571
rect 45845 9537 45879 9571
rect 46673 9537 46707 9571
rect 47593 9537 47627 9571
rect 48329 9537 48363 9571
rect 49249 9537 49283 9571
rect 50077 9537 50111 9571
rect 51365 9537 51399 9571
rect 52009 9537 52043 9571
rect 53021 9537 53055 9571
rect 6745 9469 6779 9503
rect 8033 9469 8067 9503
rect 8493 9469 8527 9503
rect 10885 9469 10919 9503
rect 11897 9469 11931 9503
rect 12725 9469 12759 9503
rect 14565 9469 14599 9503
rect 15393 9469 15427 9503
rect 19073 9469 19107 9503
rect 22017 9469 22051 9503
rect 22845 9469 22879 9503
rect 26985 9469 27019 9503
rect 28825 9469 28859 9503
rect 32781 9469 32815 9503
rect 41245 9469 41279 9503
rect 42441 9469 42475 9503
rect 46029 9469 46063 9503
rect 48973 9469 49007 9503
rect 52745 9469 52779 9503
rect 5825 9401 5859 9435
rect 35725 9401 35759 9435
rect 44833 9401 44867 9435
rect 48513 9401 48547 9435
rect 52193 9401 52227 9435
rect 1961 9333 1995 9367
rect 4997 9333 5031 9367
rect 7665 9333 7699 9367
rect 9505 9333 9539 9367
rect 14105 9333 14139 9367
rect 19441 9333 19475 9367
rect 25237 9333 25271 9367
rect 30297 9333 30331 9367
rect 31401 9333 31435 9367
rect 37841 9333 37875 9367
rect 40693 9333 40727 9367
rect 43453 9333 43487 9367
rect 51549 9333 51583 9367
rect 2421 9129 2455 9163
rect 4169 9129 4203 9163
rect 6929 9129 6963 9163
rect 9321 9129 9355 9163
rect 12265 9129 12299 9163
rect 12909 9129 12943 9163
rect 18613 9129 18647 9163
rect 19809 9129 19843 9163
rect 20269 9129 20303 9163
rect 26341 9129 26375 9163
rect 29009 9129 29043 9163
rect 31585 9129 31619 9163
rect 32965 9129 32999 9163
rect 35265 9129 35299 9163
rect 37749 9129 37783 9163
rect 42165 9129 42199 9163
rect 42625 9129 42659 9163
rect 44465 9129 44499 9163
rect 48145 9129 48179 9163
rect 51273 9129 51307 9163
rect 1685 9061 1719 9095
rect 5641 9061 5675 9095
rect 10425 9061 10459 9095
rect 15209 9061 15243 9095
rect 15853 9061 15887 9095
rect 21833 9061 21867 9095
rect 25053 9061 25087 9095
rect 25697 9061 25731 9095
rect 33425 9061 33459 9095
rect 34713 9061 34747 9095
rect 38209 9061 38243 9095
rect 50537 9061 50571 9095
rect 3249 8993 3283 9027
rect 4629 8993 4663 9027
rect 7389 8993 7423 9027
rect 16681 8993 16715 9027
rect 20637 8993 20671 9027
rect 22293 8993 22327 9027
rect 35357 8993 35391 9027
rect 36829 8993 36863 9027
rect 39865 8993 39899 9027
rect 44097 8993 44131 9027
rect 45017 8993 45051 9027
rect 48605 8993 48639 9027
rect 52377 8993 52411 9027
rect 1593 8925 1627 8959
rect 1777 8925 1811 8959
rect 2237 8925 2271 8959
rect 2881 8925 2915 8959
rect 3065 8925 3099 8959
rect 3985 8925 4019 8959
rect 4905 8925 4939 8959
rect 6101 8925 6135 8959
rect 6745 8925 6779 8959
rect 7665 8925 7699 8959
rect 9137 8925 9171 8959
rect 9781 8925 9815 8959
rect 10609 8925 10643 8959
rect 10793 8925 10827 8959
rect 11253 8925 11287 8959
rect 11529 8925 11563 8959
rect 12725 8925 12759 8959
rect 13369 8925 13403 8959
rect 14197 8925 14231 8959
rect 14473 8925 14507 8959
rect 15669 8925 15703 8959
rect 16497 8925 16531 8959
rect 17141 8925 17175 8959
rect 17417 8925 17451 8959
rect 19625 8925 19659 8959
rect 20453 8925 20487 8959
rect 21649 8925 21683 8959
rect 22569 8925 22603 8959
rect 24869 8925 24903 8959
rect 25513 8925 25547 8959
rect 26157 8925 26191 8959
rect 27997 8925 28031 8959
rect 28181 8925 28215 8959
rect 28641 8925 28675 8959
rect 28825 8925 28859 8959
rect 30481 8925 30515 8959
rect 30757 8925 30791 8959
rect 31217 8925 31251 8959
rect 31401 8925 31435 8959
rect 32781 8925 32815 8959
rect 33609 8925 33643 8959
rect 35265 8925 35299 8959
rect 36461 8925 36495 8959
rect 36645 8925 36679 8959
rect 37381 8925 37415 8959
rect 37565 8925 37599 8959
rect 38393 8925 38427 8959
rect 38945 8925 38979 8959
rect 39129 8925 39163 8959
rect 40049 8925 40083 8959
rect 40693 8925 40727 8959
rect 41337 8925 41371 8959
rect 41981 8925 42015 8959
rect 43361 8925 43395 8959
rect 43637 8925 43671 8959
rect 44281 8925 44315 8959
rect 46397 8925 46431 8959
rect 46673 8925 46707 8959
rect 47869 8925 47903 8959
rect 47961 8925 47995 8959
rect 48881 8925 48915 8959
rect 51457 8925 51491 8959
rect 51641 8925 51675 8959
rect 52653 8925 52687 8959
rect 53481 8925 53515 8959
rect 54125 8925 54159 8959
rect 16313 8857 16347 8891
rect 26801 8857 26835 8891
rect 26985 8857 27019 8891
rect 27169 8857 27203 8891
rect 47133 8857 47167 8891
rect 50721 8857 50755 8891
rect 6285 8789 6319 8823
rect 8401 8789 8435 8823
rect 9965 8789 9999 8823
rect 13461 8789 13495 8823
rect 18153 8789 18187 8823
rect 21189 8789 21223 8823
rect 23305 8789 23339 8823
rect 23857 8789 23891 8823
rect 27997 8789 28031 8823
rect 29745 8789 29779 8823
rect 32045 8789 32079 8823
rect 34069 8789 34103 8823
rect 35633 8789 35667 8823
rect 39313 8789 39347 8823
rect 40233 8789 40267 8823
rect 40877 8789 40911 8823
rect 41521 8789 41555 8823
rect 45661 8789 45695 8823
rect 49617 8789 49651 8823
rect 53941 8789 53975 8823
rect 4721 8585 4755 8619
rect 7849 8585 7883 8619
rect 10885 8585 10919 8619
rect 12449 8585 12483 8619
rect 13369 8585 13403 8619
rect 14013 8585 14047 8619
rect 14657 8585 14691 8619
rect 18797 8585 18831 8619
rect 21097 8585 21131 8619
rect 22845 8585 22879 8619
rect 24961 8585 24995 8619
rect 27077 8585 27111 8619
rect 28549 8585 28583 8619
rect 31493 8585 31527 8619
rect 33241 8585 33275 8619
rect 34897 8585 34931 8619
rect 39037 8585 39071 8619
rect 39681 8585 39715 8619
rect 40141 8585 40175 8619
rect 43453 8585 43487 8619
rect 43913 8585 43947 8619
rect 44925 8585 44959 8619
rect 49065 8585 49099 8619
rect 51825 8585 51859 8619
rect 53113 8585 53147 8619
rect 9045 8517 9079 8551
rect 11529 8517 11563 8551
rect 48421 8517 48455 8551
rect 1593 8449 1627 8483
rect 1777 8449 1811 8483
rect 2421 8449 2455 8483
rect 3525 8449 3559 8483
rect 3709 8449 3743 8483
rect 4353 8449 4387 8483
rect 4537 8449 4571 8483
rect 5825 8449 5859 8483
rect 6653 8449 6687 8483
rect 8033 8449 8067 8483
rect 8217 8449 8251 8483
rect 9229 8449 9263 8483
rect 9321 8449 9355 8483
rect 10149 8449 10183 8483
rect 10333 8449 10367 8483
rect 10793 8449 10827 8483
rect 10977 8449 11011 8483
rect 11713 8449 11747 8483
rect 11805 8449 11839 8483
rect 12633 8449 12667 8483
rect 13829 8449 13863 8483
rect 14473 8449 14507 8483
rect 15117 8449 15151 8483
rect 15301 8449 15335 8483
rect 15945 8449 15979 8483
rect 17049 8449 17083 8483
rect 17877 8449 17911 8483
rect 18613 8449 18647 8483
rect 19441 8449 19475 8483
rect 19625 8449 19659 8483
rect 20361 8449 20395 8483
rect 22293 8449 22327 8483
rect 23029 8449 23063 8483
rect 23673 8449 23707 8483
rect 24317 8449 24351 8483
rect 24501 8449 24535 8483
rect 25697 8449 25731 8483
rect 25973 8449 26007 8483
rect 27261 8449 27295 8483
rect 27353 8449 27387 8483
rect 28365 8449 28399 8483
rect 28549 8449 28583 8483
rect 29101 8449 29135 8483
rect 30205 8449 30239 8483
rect 30849 8449 30883 8483
rect 31033 8449 31067 8483
rect 32137 8449 32171 8483
rect 33425 8449 33459 8483
rect 34253 8449 34287 8483
rect 34345 8449 34379 8483
rect 35081 8449 35115 8483
rect 35817 8449 35851 8483
rect 37841 8449 37875 8483
rect 38025 8449 38059 8483
rect 38761 8449 38795 8483
rect 38853 8449 38887 8483
rect 39497 8449 39531 8483
rect 40325 8449 40359 8483
rect 41153 8449 41187 8483
rect 42625 8449 42659 8483
rect 42809 8449 42843 8483
rect 43269 8449 43303 8483
rect 44097 8449 44131 8483
rect 44741 8449 44775 8483
rect 46213 8449 46247 8483
rect 46765 8449 46799 8483
rect 46857 8449 46891 8483
rect 49249 8449 49283 8483
rect 50077 8449 50111 8483
rect 50813 8449 50847 8483
rect 51641 8449 51675 8483
rect 52929 8449 52963 8483
rect 2605 8381 2639 8415
rect 6377 8381 6411 8415
rect 12817 8381 12851 8415
rect 15761 8381 15795 8415
rect 16129 8381 16163 8415
rect 17233 8381 17267 8415
rect 18061 8381 18095 8415
rect 20085 8381 20119 8415
rect 23213 8381 23247 8415
rect 30021 8381 30055 8415
rect 33609 8381 33643 8415
rect 35541 8381 35575 8415
rect 37289 8381 37323 8415
rect 40877 8381 40911 8415
rect 42441 8381 42475 8415
rect 45937 8381 45971 8415
rect 48237 8381 48271 8415
rect 49433 8381 49467 8415
rect 51457 8381 51491 8415
rect 52745 8381 52779 8415
rect 54677 8381 54711 8415
rect 1685 8313 1719 8347
rect 3341 8313 3375 8347
rect 10333 8313 10367 8347
rect 16865 8313 16899 8347
rect 22109 8313 22143 8347
rect 23857 8313 23891 8347
rect 24501 8313 24535 8347
rect 29561 8313 29595 8347
rect 31033 8313 31067 8347
rect 32321 8313 32355 8347
rect 38209 8313 38243 8347
rect 49893 8313 49927 8347
rect 53573 8313 53607 8347
rect 54217 8313 54251 8347
rect 2237 8245 2271 8279
rect 5641 8245 5675 8279
rect 7389 8245 7423 8279
rect 15301 8245 15335 8279
rect 17693 8245 17727 8279
rect 19257 8245 19291 8279
rect 29193 8245 29227 8279
rect 30389 8245 30423 8279
rect 34069 8245 34103 8279
rect 41889 8245 41923 8279
rect 47041 8245 47075 8279
rect 47593 8245 47627 8279
rect 50629 8245 50663 8279
rect 7757 8041 7791 8075
rect 15853 8041 15887 8075
rect 16589 8041 16623 8075
rect 18061 8041 18095 8075
rect 22753 8041 22787 8075
rect 24409 8041 24443 8075
rect 25513 8041 25547 8075
rect 26893 8041 26927 8075
rect 28457 8041 28491 8075
rect 28733 8041 28767 8075
rect 32689 8041 32723 8075
rect 35081 8041 35115 8075
rect 38393 8041 38427 8075
rect 43269 8041 43303 8075
rect 46305 8041 46339 8075
rect 46765 8041 46799 8075
rect 49617 8041 49651 8075
rect 51181 8041 51215 8075
rect 51641 8041 51675 8075
rect 4537 7973 4571 8007
rect 11437 7973 11471 8007
rect 14381 7973 14415 8007
rect 33517 7973 33551 8007
rect 40233 7973 40267 8007
rect 2881 7905 2915 7939
rect 14841 7905 14875 7939
rect 26433 7905 26467 7939
rect 34069 7905 34103 7939
rect 36369 7905 36403 7939
rect 37381 7905 37415 7939
rect 45293 7905 45327 7939
rect 48789 7905 48823 7939
rect 1869 7837 1903 7871
rect 2697 7837 2731 7871
rect 4353 7837 4387 7871
rect 4997 7837 5031 7871
rect 5641 7837 5675 7871
rect 5917 7837 5951 7871
rect 7573 7837 7607 7871
rect 8217 7837 8251 7871
rect 9229 7837 9263 7871
rect 9689 7837 9723 7871
rect 9965 7837 9999 7871
rect 12633 7837 12667 7871
rect 12909 7837 12943 7871
rect 13369 7837 13403 7871
rect 14197 7837 14231 7871
rect 15117 7837 15151 7871
rect 16773 7837 16807 7871
rect 16957 7837 16991 7871
rect 17877 7837 17911 7871
rect 18061 7837 18095 7871
rect 18521 7837 18555 7871
rect 18705 7837 18739 7871
rect 19257 7837 19291 7871
rect 20545 7837 20579 7871
rect 20821 7837 20855 7871
rect 21281 7837 21315 7871
rect 21465 7837 21499 7871
rect 22201 7837 22235 7871
rect 23673 7837 23707 7871
rect 23857 7837 23891 7871
rect 24593 7837 24627 7871
rect 24777 7837 24811 7871
rect 25881 7837 25915 7871
rect 27077 7837 27111 7871
rect 27537 7837 27571 7871
rect 27813 7837 27847 7871
rect 27905 7837 27939 7871
rect 28917 7837 28951 7871
rect 30665 7837 30699 7871
rect 31217 7837 31251 7871
rect 32045 7837 32079 7871
rect 32229 7837 32263 7871
rect 32873 7837 32907 7871
rect 33333 7837 33367 7871
rect 33517 7837 33551 7871
rect 33977 7837 34011 7871
rect 34161 7837 34195 7871
rect 34713 7837 34747 7871
rect 36645 7837 36679 7871
rect 37197 7837 37231 7871
rect 38025 7837 38059 7871
rect 38209 7837 38243 7871
rect 38853 7837 38887 7871
rect 39037 7837 39071 7871
rect 41429 7837 41463 7871
rect 41705 7837 41739 7871
rect 43085 7837 43119 7871
rect 44189 7837 44223 7871
rect 45569 7837 45603 7871
rect 46949 7837 46983 7871
rect 47777 7837 47811 7871
rect 48421 7837 48455 7871
rect 48605 7837 48639 7871
rect 49249 7837 49283 7871
rect 49433 7837 49467 7871
rect 50169 7837 50203 7871
rect 50445 7837 50479 7871
rect 53941 7837 53975 7871
rect 18613 7769 18647 7803
rect 22845 7769 22879 7803
rect 23765 7769 23799 7803
rect 25697 7769 25731 7803
rect 30021 7769 30055 7803
rect 34897 7769 34931 7803
rect 40417 7769 40451 7803
rect 42901 7769 42935 7803
rect 53389 7769 53423 7803
rect 54585 7769 54619 7803
rect 2053 7701 2087 7735
rect 2513 7701 2547 7735
rect 3893 7701 3927 7735
rect 5181 7701 5215 7735
rect 6653 7701 6687 7735
rect 8401 7701 8435 7735
rect 10701 7701 10735 7735
rect 11897 7701 11931 7735
rect 13553 7701 13587 7735
rect 19441 7701 19475 7735
rect 21649 7701 21683 7735
rect 30113 7701 30147 7735
rect 31401 7701 31435 7735
rect 31861 7701 31895 7735
rect 39221 7701 39255 7735
rect 42441 7701 42475 7735
rect 44373 7701 44407 7735
rect 47961 7701 47995 7735
rect 52193 7701 52227 7735
rect 52745 7701 52779 7735
rect 54125 7701 54159 7735
rect 55321 7701 55355 7735
rect 1777 7497 1811 7531
rect 6377 7497 6411 7531
rect 9045 7497 9079 7531
rect 10977 7497 11011 7531
rect 17693 7497 17727 7531
rect 31585 7497 31619 7531
rect 34161 7497 34195 7531
rect 46029 7497 46063 7531
rect 51365 7497 51399 7531
rect 52009 7497 52043 7531
rect 53113 7497 53147 7531
rect 11529 7429 11563 7463
rect 24409 7429 24443 7463
rect 38301 7429 38335 7463
rect 44649 7429 44683 7463
rect 1593 7361 1627 7395
rect 2421 7361 2455 7395
rect 3249 7361 3283 7395
rect 3433 7361 3467 7395
rect 4905 7361 4939 7395
rect 5641 7361 5675 7395
rect 6561 7361 6595 7395
rect 6653 7361 6687 7395
rect 7389 7361 7423 7395
rect 8309 7361 8343 7395
rect 9689 7361 9723 7395
rect 10793 7361 10827 7395
rect 11713 7361 11747 7395
rect 12449 7361 12483 7395
rect 13093 7361 13127 7395
rect 13921 7361 13955 7395
rect 14105 7361 14139 7395
rect 14197 7361 14231 7395
rect 15393 7361 15427 7395
rect 17233 7361 17267 7395
rect 17877 7361 17911 7395
rect 18337 7361 18371 7395
rect 19625 7361 19659 7395
rect 21097 7361 21131 7395
rect 21281 7361 21315 7395
rect 22109 7361 22143 7395
rect 22845 7361 22879 7395
rect 24317 7361 24351 7395
rect 24501 7361 24535 7395
rect 25697 7361 25731 7395
rect 26065 7361 26099 7395
rect 26433 7361 26467 7395
rect 29009 7361 29043 7395
rect 30205 7361 30239 7395
rect 31401 7361 31435 7395
rect 32689 7361 32723 7395
rect 33977 7361 34011 7395
rect 34621 7361 34655 7395
rect 35541 7361 35575 7395
rect 37473 7361 37507 7395
rect 37565 7361 37599 7395
rect 39221 7361 39255 7395
rect 40417 7361 40451 7395
rect 40693 7361 40727 7395
rect 42809 7361 42843 7395
rect 43545 7361 43579 7395
rect 43637 7361 43671 7395
rect 44465 7361 44499 7395
rect 45385 7361 45419 7395
rect 45569 7361 45603 7395
rect 46213 7361 46247 7395
rect 46673 7361 46707 7395
rect 48237 7361 48271 7395
rect 49341 7361 49375 7395
rect 50353 7361 50387 7395
rect 50629 7361 50663 7395
rect 52101 7361 52135 7395
rect 52929 7361 52963 7395
rect 54217 7361 54251 7395
rect 55689 7361 55723 7395
rect 56333 7361 56367 7395
rect 56517 7361 56551 7395
rect 57897 7361 57931 7395
rect 2605 7293 2639 7327
rect 5181 7293 5215 7327
rect 7573 7293 7607 7327
rect 8033 7293 8067 7327
rect 9505 7293 9539 7327
rect 9873 7293 9907 7327
rect 11897 7293 11931 7327
rect 15117 7293 15151 7327
rect 19901 7293 19935 7327
rect 22569 7293 22603 7327
rect 25053 7293 25087 7327
rect 25145 7293 25179 7327
rect 26985 7293 27019 7327
rect 27261 7293 27295 7327
rect 28641 7293 28675 7327
rect 28733 7293 28767 7327
rect 29929 7293 29963 7327
rect 32413 7293 32447 7327
rect 35265 7293 35299 7327
rect 38945 7293 38979 7327
rect 44281 7293 44315 7327
rect 45201 7293 45235 7327
rect 48053 7293 48087 7327
rect 49157 7293 49191 7327
rect 52745 7293 52779 7327
rect 53941 7293 53975 7327
rect 56425 7293 56459 7327
rect 7205 7225 7239 7259
rect 13277 7225 13311 7259
rect 38117 7225 38151 7259
rect 41429 7225 41463 7259
rect 42993 7225 43027 7259
rect 48421 7225 48455 7259
rect 2237 7157 2271 7191
rect 3065 7157 3099 7191
rect 4169 7157 4203 7191
rect 5825 7157 5859 7191
rect 12541 7157 12575 7191
rect 16129 7157 16163 7191
rect 17049 7157 17083 7191
rect 18521 7157 18555 7191
rect 19165 7157 19199 7191
rect 20913 7157 20947 7191
rect 21925 7157 21959 7191
rect 23581 7157 23615 7191
rect 33425 7157 33459 7191
rect 34713 7157 34747 7191
rect 36277 7157 36311 7191
rect 37289 7157 37323 7191
rect 39957 7157 39991 7191
rect 43821 7157 43855 7191
rect 46857 7157 46891 7191
rect 49525 7157 49559 7191
rect 54953 7157 54987 7191
rect 55873 7157 55907 7191
rect 57989 7157 58023 7191
rect 5641 6953 5675 6987
rect 6101 6953 6135 6987
rect 17969 6953 18003 6987
rect 21833 6953 21867 6987
rect 23305 6953 23339 6987
rect 29745 6953 29779 6987
rect 30573 6953 30607 6987
rect 36369 6953 36403 6987
rect 48605 6953 48639 6987
rect 51273 6953 51307 6987
rect 55873 6953 55907 6987
rect 1961 6885 1995 6919
rect 15669 6885 15703 6919
rect 23857 6885 23891 6919
rect 26985 6885 27019 6919
rect 37841 6885 37875 6919
rect 41613 6885 41647 6919
rect 56793 6885 56827 6919
rect 11069 6817 11103 6851
rect 16957 6817 16991 6851
rect 19257 6817 19291 6851
rect 22293 6817 22327 6851
rect 24409 6817 24443 6851
rect 25789 6817 25823 6851
rect 28733 6817 28767 6851
rect 31493 6817 31527 6851
rect 32045 6817 32079 6851
rect 35817 6817 35851 6851
rect 36185 6817 36219 6851
rect 39037 6817 39071 6851
rect 40233 6817 40267 6851
rect 44465 6817 44499 6851
rect 45017 6817 45051 6851
rect 52009 6817 52043 6851
rect 53849 6817 53883 6851
rect 57805 6817 57839 6851
rect 1777 6749 1811 6783
rect 2421 6749 2455 6783
rect 3249 6749 3283 6783
rect 3801 6749 3835 6783
rect 4077 6749 4111 6783
rect 5457 6749 5491 6783
rect 6285 6749 6319 6783
rect 6745 6749 6779 6783
rect 6929 6749 6963 6783
rect 7021 6749 7055 6783
rect 7113 6749 7147 6783
rect 8401 6749 8435 6783
rect 9505 6749 9539 6783
rect 10149 6749 10183 6783
rect 11345 6719 11379 6753
rect 13277 6749 13311 6783
rect 13553 6749 13587 6783
rect 14105 6749 14139 6783
rect 15025 6749 15059 6783
rect 15853 6749 15887 6783
rect 16497 6749 16531 6783
rect 17233 6749 17267 6783
rect 18705 6749 18739 6783
rect 19533 6749 19567 6783
rect 21189 6749 21223 6783
rect 21649 6749 21683 6783
rect 22569 6749 22603 6783
rect 25881 6749 25915 6783
rect 26157 6749 26191 6783
rect 29009 6749 29043 6783
rect 30021 6749 30055 6783
rect 30481 6749 30515 6783
rect 30665 6749 30699 6783
rect 31953 6749 31987 6783
rect 32413 6749 32447 6783
rect 33241 6749 33275 6783
rect 33977 6749 34011 6783
rect 36829 6749 36863 6783
rect 37105 6749 37139 6783
rect 38393 6749 38427 6783
rect 41337 6749 41371 6783
rect 42441 6749 42475 6783
rect 44189 6749 44223 6783
rect 45293 6749 45327 6783
rect 46581 6749 46615 6783
rect 46857 6749 46891 6783
rect 49341 6749 49375 6783
rect 49617 6749 49651 6783
rect 50261 6749 50295 6783
rect 50537 6749 50571 6783
rect 53573 6749 53607 6783
rect 57529 6749 57563 6783
rect 10333 6681 10367 6715
rect 24961 6681 24995 6715
rect 25145 6681 25179 6715
rect 25329 6681 25363 6715
rect 26617 6681 26651 6715
rect 26801 6681 26835 6715
rect 27537 6681 27571 6715
rect 27721 6681 27755 6715
rect 32965 6681 32999 6715
rect 35081 6681 35115 6715
rect 35265 6681 35299 6715
rect 39221 6681 39255 6715
rect 40417 6681 40451 6715
rect 41613 6681 41647 6715
rect 42625 6681 42659 6715
rect 51825 6681 51859 6715
rect 54309 6681 54343 6715
rect 55689 6681 55723 6715
rect 2605 6613 2639 6647
rect 4813 6613 4847 6647
rect 7389 6613 7423 6647
rect 8217 6613 8251 6647
rect 9321 6613 9355 6647
rect 12081 6613 12115 6647
rect 12541 6613 12575 6647
rect 14289 6613 14323 6647
rect 15209 6613 15243 6647
rect 20269 6613 20303 6647
rect 29561 6613 29595 6647
rect 33063 6613 33097 6647
rect 33149 6613 33183 6647
rect 34161 6613 34195 6647
rect 36001 6613 36035 6647
rect 38577 6613 38611 6647
rect 41429 6613 41463 6647
rect 43453 6613 43487 6647
rect 46029 6613 46063 6647
rect 47593 6613 47627 6647
rect 48053 6613 48087 6647
rect 52837 6613 52871 6647
rect 55889 6613 55923 6647
rect 56057 6613 56091 6647
rect 8309 6409 8343 6443
rect 9873 6409 9907 6443
rect 19809 6409 19843 6443
rect 23489 6409 23523 6443
rect 30757 6409 30791 6443
rect 35449 6409 35483 6443
rect 37473 6409 37507 6443
rect 40785 6409 40819 6443
rect 47685 6409 47719 6443
rect 50537 6409 50571 6443
rect 57897 6409 57931 6443
rect 15945 6341 15979 6375
rect 18581 6341 18615 6375
rect 18797 6341 18831 6375
rect 30389 6341 30423 6375
rect 30589 6341 30623 6375
rect 32137 6341 32171 6375
rect 33057 6341 33091 6375
rect 33241 6341 33275 6375
rect 33793 6341 33827 6375
rect 39773 6341 39807 6375
rect 42993 6341 43027 6375
rect 46949 6341 46983 6375
rect 2053 6273 2087 6307
rect 2513 6273 2547 6307
rect 3893 6273 3927 6307
rect 4629 6273 4663 6307
rect 4813 6273 4847 6307
rect 4908 6276 4942 6310
rect 4997 6273 5031 6307
rect 7573 6273 7607 6307
rect 9137 6273 9171 6307
rect 10321 6273 10355 6307
rect 10496 6276 10530 6310
rect 10609 6273 10643 6307
rect 10701 6273 10735 6307
rect 11529 6273 11563 6307
rect 12725 6273 12759 6307
rect 13461 6273 13495 6307
rect 13640 6273 13674 6307
rect 13737 6273 13771 6307
rect 13829 6273 13863 6307
rect 14749 6273 14783 6307
rect 14933 6273 14967 6307
rect 17417 6273 17451 6307
rect 17509 6273 17543 6307
rect 19625 6273 19659 6307
rect 20269 6273 20303 6307
rect 20545 6273 20579 6307
rect 21833 6273 21867 6307
rect 22017 6273 22051 6307
rect 22109 6273 22143 6307
rect 22201 6273 22235 6307
rect 23397 6273 23431 6307
rect 23581 6273 23615 6307
rect 24041 6273 24075 6307
rect 24225 6273 24259 6307
rect 25099 6273 25133 6307
rect 25237 6273 25271 6307
rect 25329 6273 25363 6307
rect 25513 6273 25547 6307
rect 25973 6273 26007 6307
rect 26157 6273 26191 6307
rect 27261 6273 27295 6307
rect 27905 6273 27939 6307
rect 28089 6273 28123 6307
rect 28181 6273 28215 6307
rect 28293 6273 28327 6307
rect 29285 6273 29319 6307
rect 29469 6273 29503 6307
rect 29561 6273 29595 6307
rect 29653 6273 29687 6307
rect 32229 6273 32263 6307
rect 32413 6273 32447 6307
rect 34437 6273 34471 6307
rect 34621 6273 34655 6307
rect 35265 6273 35299 6307
rect 35541 6273 35575 6307
rect 36369 6273 36403 6307
rect 37473 6273 37507 6307
rect 37565 6273 37599 6307
rect 37749 6273 37783 6307
rect 40601 6273 40635 6307
rect 41521 6273 41555 6307
rect 41705 6273 41739 6307
rect 45118 6273 45152 6307
rect 45385 6273 45419 6307
rect 46857 6273 46891 6307
rect 50077 6273 50111 6307
rect 50721 6273 50755 6307
rect 51917 6273 51951 6307
rect 53849 6273 53883 6307
rect 55413 6273 55447 6307
rect 56149 6273 56183 6307
rect 56977 6273 57011 6307
rect 58081 6273 58115 6307
rect 4169 6205 4203 6239
rect 7297 6205 7331 6239
rect 8861 6205 8895 6239
rect 17877 6205 17911 6239
rect 32505 6205 32539 6239
rect 34345 6205 34379 6239
rect 38301 6205 38335 6239
rect 40049 6205 40083 6239
rect 41797 6205 41831 6239
rect 49157 6205 49191 6239
rect 49433 6205 49467 6239
rect 52193 6205 52227 6239
rect 54125 6205 54159 6239
rect 55137 6205 55171 6239
rect 55873 6205 55907 6239
rect 2697 6137 2731 6171
rect 5273 6137 5307 6171
rect 14105 6137 14139 6171
rect 24409 6137 24443 6171
rect 26157 6137 26191 6171
rect 27445 6137 27479 6171
rect 35265 6137 35299 6171
rect 42441 6137 42475 6171
rect 44005 6137 44039 6171
rect 45845 6137 45879 6171
rect 51181 6137 51215 6171
rect 56793 6137 56827 6171
rect 1869 6069 1903 6103
rect 3157 6069 3191 6103
rect 5733 6069 5767 6103
rect 6837 6069 6871 6103
rect 10977 6069 11011 6103
rect 11713 6069 11747 6103
rect 12909 6069 12943 6103
rect 14565 6069 14599 6103
rect 16037 6069 16071 6103
rect 16773 6069 16807 6103
rect 17233 6069 17267 6103
rect 18429 6069 18463 6103
rect 18613 6069 18647 6103
rect 21281 6069 21315 6103
rect 22477 6069 22511 6103
rect 24869 6069 24903 6103
rect 28549 6069 28583 6103
rect 29929 6069 29963 6103
rect 30573 6069 30607 6103
rect 31217 6069 31251 6103
rect 32597 6069 32631 6103
rect 34805 6069 34839 6103
rect 36553 6069 36587 6103
rect 41337 6069 41371 6103
rect 49893 6069 49927 6103
rect 53113 6069 53147 6103
rect 55965 6069 55999 6103
rect 56333 6069 56367 6103
rect 1777 5865 1811 5899
rect 2421 5865 2455 5899
rect 8217 5865 8251 5899
rect 10057 5865 10091 5899
rect 17509 5865 17543 5899
rect 19625 5865 19659 5899
rect 26065 5865 26099 5899
rect 27169 5865 27203 5899
rect 29929 5865 29963 5899
rect 33149 5865 33183 5899
rect 33793 5865 33827 5899
rect 34713 5865 34747 5899
rect 35633 5865 35667 5899
rect 41324 5865 41358 5899
rect 42809 5865 42843 5899
rect 44005 5865 44039 5899
rect 51549 5865 51583 5899
rect 53573 5865 53607 5899
rect 3249 5797 3283 5831
rect 6653 5797 6687 5831
rect 31309 5797 31343 5831
rect 37841 5797 37875 5831
rect 39957 5797 39991 5831
rect 43361 5797 43395 5831
rect 46305 5797 46339 5831
rect 50261 5797 50295 5831
rect 50813 5797 50847 5831
rect 56609 5797 56643 5831
rect 14105 5729 14139 5763
rect 23121 5729 23155 5763
rect 24685 5729 24719 5763
rect 36369 5729 36403 5763
rect 41061 5729 41095 5763
rect 47869 5729 47903 5763
rect 48145 5729 48179 5763
rect 52561 5729 52595 5763
rect 57621 5729 57655 5763
rect 1593 5661 1627 5695
rect 2237 5661 2271 5695
rect 2881 5661 2915 5695
rect 3801 5661 3835 5695
rect 3980 5661 4014 5695
rect 4080 5655 4114 5689
rect 4169 5661 4203 5695
rect 5273 5661 5307 5695
rect 5540 5661 5574 5695
rect 7665 5661 7699 5695
rect 8401 5661 8435 5695
rect 9229 5661 9263 5695
rect 9873 5661 9907 5695
rect 10701 5661 10735 5695
rect 12541 5661 12575 5695
rect 13461 5661 13495 5695
rect 14361 5661 14395 5695
rect 16405 5661 16439 5695
rect 16589 5661 16623 5695
rect 16681 5661 16715 5695
rect 16819 5661 16853 5695
rect 18061 5661 18095 5695
rect 18245 5661 18279 5695
rect 18337 5661 18371 5695
rect 18429 5661 18463 5695
rect 20637 5661 20671 5695
rect 21281 5661 21315 5695
rect 22854 5661 22888 5695
rect 23857 5661 23891 5695
rect 24952 5661 24986 5695
rect 26801 5661 26835 5695
rect 28742 5661 28776 5695
rect 29009 5661 29043 5695
rect 29745 5661 29779 5695
rect 30389 5661 30423 5695
rect 32689 5661 32723 5695
rect 34897 5661 34931 5695
rect 34989 5661 35023 5695
rect 35449 5661 35483 5695
rect 36093 5661 36127 5695
rect 38577 5661 38611 5695
rect 40417 5661 40451 5695
rect 44189 5661 44223 5695
rect 45017 5661 45051 5695
rect 45661 5661 45695 5695
rect 47225 5661 47259 5695
rect 50169 5661 50203 5695
rect 52285 5661 52319 5695
rect 54125 5661 54159 5695
rect 55321 5661 55355 5695
rect 55597 5661 55631 5695
rect 57345 5661 57379 5695
rect 3065 5593 3099 5627
rect 9689 5593 9723 5627
rect 10968 5593 11002 5627
rect 13277 5593 13311 5627
rect 19257 5593 19291 5627
rect 19441 5593 19475 5627
rect 26985 5593 27019 5627
rect 29561 5593 29595 5627
rect 32422 5593 32456 5627
rect 34713 5593 34747 5627
rect 38485 5593 38519 5627
rect 4445 5525 4479 5559
rect 7481 5525 7515 5559
rect 9045 5525 9079 5559
rect 12081 5525 12115 5559
rect 12725 5525 12759 5559
rect 15485 5525 15519 5559
rect 17049 5525 17083 5559
rect 18705 5525 18739 5559
rect 21741 5525 21775 5559
rect 27629 5525 27663 5559
rect 39129 5525 39163 5559
rect 40601 5525 40635 5559
rect 45201 5525 45235 5559
rect 47317 5525 47351 5559
rect 49617 5525 49651 5559
rect 53113 5525 53147 5559
rect 54217 5525 54251 5559
rect 58081 5525 58115 5559
rect 2329 5321 2363 5355
rect 9045 5321 9079 5355
rect 16129 5321 16163 5355
rect 16681 5321 16715 5355
rect 18521 5321 18555 5355
rect 19901 5321 19935 5355
rect 24685 5321 24719 5355
rect 32505 5321 32539 5355
rect 37565 5321 37599 5355
rect 42533 5321 42567 5355
rect 46857 5321 46891 5355
rect 47593 5321 47627 5355
rect 52745 5321 52779 5355
rect 52929 5321 52963 5355
rect 54953 5321 54987 5355
rect 57897 5321 57931 5355
rect 1961 5253 1995 5287
rect 2789 5253 2823 5287
rect 3157 5253 3191 5287
rect 7910 5253 7944 5287
rect 9505 5253 9539 5287
rect 9873 5253 9907 5287
rect 15945 5253 15979 5287
rect 17794 5253 17828 5287
rect 18889 5253 18923 5287
rect 21014 5253 21048 5287
rect 33241 5253 33275 5287
rect 55321 5253 55355 5287
rect 2145 5185 2179 5219
rect 2973 5185 3007 5219
rect 3801 5185 3835 5219
rect 4445 5185 4479 5219
rect 4701 5185 4735 5219
rect 7205 5185 7239 5219
rect 7665 5185 7699 5219
rect 9689 5185 9723 5219
rect 10609 5185 10643 5219
rect 10701 5185 10735 5219
rect 10793 5185 10827 5219
rect 10989 5185 11023 5219
rect 11805 5185 11839 5219
rect 14105 5185 14139 5219
rect 14381 5185 14415 5219
rect 15761 5185 15795 5219
rect 18705 5185 18739 5219
rect 21833 5185 21867 5219
rect 23305 5185 23339 5219
rect 23561 5185 23595 5219
rect 25697 5185 25731 5219
rect 25881 5185 25915 5219
rect 25973 5185 26007 5219
rect 26985 5185 27019 5219
rect 27721 5185 27755 5219
rect 27905 5185 27939 5219
rect 27997 5185 28031 5219
rect 28457 5185 28491 5219
rect 28733 5185 28767 5219
rect 30205 5185 30239 5219
rect 30461 5185 30495 5219
rect 32321 5185 32355 5219
rect 32597 5185 32631 5219
rect 35633 5185 35667 5219
rect 37657 5185 37691 5219
rect 38761 5185 38795 5219
rect 38945 5185 38979 5219
rect 39037 5185 39071 5219
rect 39845 5185 39879 5219
rect 42625 5185 42659 5219
rect 43545 5185 43579 5219
rect 43812 5185 43846 5219
rect 45569 5185 45603 5219
rect 45753 5185 45787 5219
rect 45845 5185 45879 5219
rect 47041 5185 47075 5219
rect 49893 5185 49927 5219
rect 52101 5185 52135 5219
rect 52926 5185 52960 5219
rect 54217 5185 54251 5219
rect 54309 5185 54343 5219
rect 54861 5185 54895 5219
rect 55137 5185 55171 5219
rect 55965 5185 55999 5219
rect 56793 5185 56827 5219
rect 58081 5185 58115 5219
rect 1501 5117 1535 5151
rect 6469 5117 6503 5151
rect 11529 5117 11563 5151
rect 12817 5117 12851 5151
rect 13093 5117 13127 5151
rect 18061 5117 18095 5151
rect 21281 5117 21315 5151
rect 28549 5117 28583 5151
rect 35265 5117 35299 5151
rect 39589 5117 39623 5151
rect 49617 5117 49651 5151
rect 53389 5117 53423 5151
rect 54033 5117 54067 5151
rect 54125 5117 54159 5151
rect 56057 5117 56091 5151
rect 3985 5049 4019 5083
rect 5825 5049 5859 5083
rect 28917 5049 28951 5083
rect 33057 5049 33091 5083
rect 41429 5049 41463 5083
rect 44925 5049 44959 5083
rect 56333 5049 56367 5083
rect 7021 4981 7055 5015
rect 10333 4981 10367 5015
rect 19349 4981 19383 5015
rect 22017 4981 22051 5015
rect 22845 4981 22879 5015
rect 25513 4981 25547 5015
rect 27537 4981 27571 5015
rect 28641 4981 28675 5015
rect 29469 4981 29503 5015
rect 31585 4981 31619 5015
rect 32137 4981 32171 5015
rect 33839 4981 33873 5015
rect 36553 4981 36587 5015
rect 38577 4981 38611 5015
rect 40969 4981 41003 5015
rect 45385 4981 45419 5015
rect 48145 4981 48179 5015
rect 50353 4981 50387 5015
rect 51089 4981 51123 5015
rect 52009 4981 52043 5015
rect 53297 4981 53331 5015
rect 53849 4981 53883 5015
rect 56149 4981 56183 5015
rect 56885 4981 56919 5015
rect 4353 4777 4387 4811
rect 8217 4777 8251 4811
rect 13093 4777 13127 4811
rect 14841 4777 14875 4811
rect 23213 4777 23247 4811
rect 24593 4777 24627 4811
rect 26065 4777 26099 4811
rect 30205 4777 30239 4811
rect 30757 4777 30791 4811
rect 35265 4777 35299 4811
rect 36645 4777 36679 4811
rect 40417 4777 40451 4811
rect 43453 4777 43487 4811
rect 45201 4777 45235 4811
rect 50169 4777 50203 4811
rect 51733 4777 51767 4811
rect 53297 4777 53331 4811
rect 54769 4777 54803 4811
rect 55505 4777 55539 4811
rect 55689 4777 55723 4811
rect 6285 4709 6319 4743
rect 17877 4709 17911 4743
rect 25145 4709 25179 4743
rect 34161 4709 34195 4743
rect 38669 4709 38703 4743
rect 47317 4709 47351 4743
rect 53941 4709 53975 4743
rect 56241 4709 56275 4743
rect 1685 4641 1719 4675
rect 6837 4641 6871 4675
rect 10149 4641 10183 4675
rect 11713 4641 11747 4675
rect 14197 4641 14231 4675
rect 16773 4641 16807 4675
rect 23857 4641 23891 4675
rect 37289 4641 37323 4675
rect 40233 4641 40267 4675
rect 41797 4641 41831 4675
rect 46397 4641 46431 4675
rect 48697 4641 48731 4675
rect 57253 4641 57287 4675
rect 2513 4573 2547 4607
rect 2697 4573 2731 4607
rect 2789 4573 2823 4607
rect 2881 4573 2915 4607
rect 4261 4573 4295 4607
rect 4905 4573 4939 4607
rect 7104 4573 7138 4607
rect 9137 4573 9171 4607
rect 9781 4573 9815 4607
rect 10609 4573 10643 4607
rect 10793 4573 10827 4607
rect 10885 4573 10919 4607
rect 10977 4573 11011 4607
rect 14657 4573 14691 4607
rect 17693 4573 17727 4607
rect 18613 4573 18647 4607
rect 19533 4573 19567 4607
rect 21373 4573 21407 4607
rect 21465 4573 21499 4607
rect 21649 4573 21683 4607
rect 22569 4573 22603 4607
rect 22748 4570 22782 4604
rect 22848 4570 22882 4604
rect 22937 4573 22971 4607
rect 25329 4573 25363 4607
rect 25605 4573 25639 4607
rect 26617 4573 26651 4607
rect 28825 4573 28859 4607
rect 29561 4573 29595 4607
rect 29745 4573 29779 4607
rect 29837 4573 29871 4607
rect 29929 4573 29963 4607
rect 31217 4573 31251 4607
rect 31401 4573 31435 4607
rect 31493 4573 31527 4607
rect 31585 4573 31619 4607
rect 32781 4573 32815 4607
rect 36001 4573 36035 4607
rect 36185 4573 36219 4607
rect 36277 4573 36311 4607
rect 36369 4573 36403 4607
rect 39129 4573 39163 4607
rect 40141 4573 40175 4607
rect 41061 4573 41095 4607
rect 41337 4573 41371 4607
rect 42809 4573 42843 4607
rect 42993 4573 43027 4607
rect 43085 4573 43119 4607
rect 43177 4573 43211 4607
rect 44189 4573 44223 4607
rect 44465 4573 44499 4607
rect 45201 4573 45235 4607
rect 45293 4573 45327 4607
rect 45937 4573 45971 4607
rect 46213 4573 46247 4607
rect 48430 4573 48464 4607
rect 49157 4573 49191 4607
rect 50813 4573 50847 4607
rect 52469 4573 52503 4607
rect 52745 4573 52779 4607
rect 53481 4573 53515 4607
rect 54585 4573 54619 4607
rect 54769 4573 54803 4607
rect 56977 4573 57011 4607
rect 57713 4573 57747 4607
rect 1869 4505 1903 4539
rect 2053 4505 2087 4539
rect 3157 4505 3191 4539
rect 5172 4505 5206 4539
rect 8953 4505 8987 4539
rect 9965 4505 9999 4539
rect 11253 4505 11287 4539
rect 11958 4505 11992 4539
rect 16528 4505 16562 4539
rect 19778 4505 19812 4539
rect 24501 4505 24535 4539
rect 25513 4505 25547 4539
rect 31861 4505 31895 4539
rect 33026 4505 33060 4539
rect 37534 4505 37568 4539
rect 40417 4505 40451 4539
rect 45477 4505 45511 4539
rect 55321 4505 55355 4539
rect 9321 4437 9355 4471
rect 15393 4437 15427 4471
rect 18429 4437 18463 4471
rect 20913 4437 20947 4471
rect 21833 4437 21867 4471
rect 27905 4437 27939 4471
rect 34805 4437 34839 4471
rect 39957 4437 39991 4471
rect 40877 4437 40911 4471
rect 41245 4437 41279 4471
rect 44005 4437 44039 4471
rect 44373 4437 44407 4471
rect 45017 4437 45051 4471
rect 46029 4437 46063 4471
rect 55521 4437 55555 4471
rect 57897 4437 57931 4471
rect 7481 4233 7515 4267
rect 8033 4233 8067 4267
rect 19441 4233 19475 4267
rect 25881 4233 25915 4267
rect 28549 4233 28583 4267
rect 37289 4233 37323 4267
rect 48329 4233 48363 4267
rect 5641 4165 5675 4199
rect 10149 4165 10183 4199
rect 13737 4165 13771 4199
rect 14841 4165 14875 4199
rect 15025 4165 15059 4199
rect 18153 4165 18187 4199
rect 55873 4165 55907 4199
rect 1869 4097 1903 4131
rect 2789 4097 2823 4131
rect 2881 4100 2915 4134
rect 2973 4097 3007 4131
rect 3157 4097 3191 4131
rect 4353 4097 4387 4131
rect 5089 4097 5123 4131
rect 6745 4097 6779 4131
rect 7297 4097 7331 4131
rect 7481 4097 7515 4131
rect 9157 4097 9191 4131
rect 10379 4097 10413 4131
rect 10517 4097 10551 4131
rect 10630 4097 10664 4131
rect 10793 4097 10827 4131
rect 11796 4097 11830 4131
rect 13967 4097 14001 4131
rect 14086 4097 14120 4131
rect 14202 4097 14236 4131
rect 14381 4097 14415 4131
rect 15853 4097 15887 4131
rect 16037 4097 16071 4131
rect 16129 4097 16163 4131
rect 16937 4097 16971 4131
rect 17030 4097 17064 4131
rect 17146 4097 17180 4131
rect 17325 4097 17359 4131
rect 18797 4097 18831 4131
rect 18981 4097 19015 4131
rect 19073 4097 19107 4131
rect 19165 4097 19199 4131
rect 21025 4097 21059 4131
rect 21281 4097 21315 4131
rect 22109 4097 22143 4131
rect 22201 4097 22235 4131
rect 22293 4097 22327 4131
rect 22477 4097 22511 4131
rect 23857 4097 23891 4131
rect 24685 4097 24719 4131
rect 24869 4097 24903 4131
rect 24961 4097 24995 4131
rect 25053 4097 25087 4131
rect 25789 4097 25823 4131
rect 26065 4097 26099 4131
rect 27169 4097 27203 4131
rect 27425 4097 27459 4131
rect 29009 4097 29043 4131
rect 29193 4097 29227 4131
rect 29837 4097 29871 4131
rect 29929 4097 29963 4131
rect 30113 4097 30147 4131
rect 30297 4097 30331 4131
rect 32137 4097 32171 4131
rect 32393 4097 32427 4131
rect 34253 4097 34287 4131
rect 35265 4097 35299 4131
rect 35449 4097 35483 4131
rect 35541 4097 35575 4131
rect 35633 4097 35667 4131
rect 37565 4097 37599 4131
rect 37657 4097 37691 4131
rect 37749 4097 37783 4131
rect 37927 4097 37961 4131
rect 39037 4097 39071 4131
rect 39313 4097 39347 4131
rect 40325 4097 40359 4131
rect 40601 4097 40635 4131
rect 41061 4097 41095 4131
rect 41153 4097 41187 4131
rect 41337 4097 41371 4131
rect 42993 4097 43027 4131
rect 43177 4097 43211 4131
rect 43269 4097 43303 4131
rect 43361 4097 43395 4131
rect 44097 4097 44131 4131
rect 44281 4097 44315 4131
rect 44373 4097 44407 4131
rect 44465 4097 44499 4131
rect 49442 4097 49476 4131
rect 49709 4097 49743 4131
rect 51733 4097 51767 4131
rect 51825 4097 51859 4131
rect 52009 4097 52043 4131
rect 52193 4097 52227 4131
rect 54033 4097 54067 4131
rect 54125 4097 54159 4131
rect 54493 4097 54527 4131
rect 55137 4097 55171 4131
rect 55781 4097 55815 4131
rect 55965 4097 55999 4131
rect 57897 4097 57931 4131
rect 9413 4029 9447 4063
rect 11529 4029 11563 4063
rect 16681 4029 16715 4063
rect 18337 4029 18371 4063
rect 21833 4029 21867 4063
rect 25329 4029 25363 4063
rect 31309 4029 31343 4063
rect 31585 4029 31619 4063
rect 33977 4029 34011 4063
rect 43637 4029 43671 4063
rect 44741 4029 44775 4063
rect 45845 4029 45879 4063
rect 55321 4029 55355 4063
rect 2513 3961 2547 3995
rect 5825 3961 5859 3995
rect 12909 3961 12943 3995
rect 15669 3961 15703 3995
rect 36369 3961 36403 3995
rect 46489 3961 46523 3995
rect 50813 3961 50847 3995
rect 53389 3961 53423 3995
rect 54309 3961 54343 3995
rect 57989 3961 58023 3995
rect 2053 3893 2087 3927
rect 4169 3893 4203 3927
rect 4905 3893 4939 3927
rect 6561 3893 6595 3927
rect 19901 3893 19935 3927
rect 23305 3893 23339 3927
rect 23949 3893 23983 3927
rect 26249 3893 26283 3927
rect 33517 3893 33551 3927
rect 35909 3893 35943 3927
rect 41521 3893 41555 3927
rect 42441 3893 42475 3927
rect 45201 3893 45235 3927
rect 47593 3893 47627 3927
rect 50169 3893 50203 3927
rect 52745 3893 52779 3927
rect 54953 3893 54987 3927
rect 56517 3893 56551 3927
rect 57069 3893 57103 3927
rect 2053 3689 2087 3723
rect 2513 3689 2547 3723
rect 3893 3689 3927 3723
rect 4445 3689 4479 3723
rect 7573 3689 7607 3723
rect 13553 3689 13587 3723
rect 15393 3689 15427 3723
rect 16773 3689 16807 3723
rect 23765 3689 23799 3723
rect 26801 3689 26835 3723
rect 32689 3689 32723 3723
rect 33425 3689 33459 3723
rect 34805 3689 34839 3723
rect 40509 3689 40543 3723
rect 50813 3689 50847 3723
rect 52285 3689 52319 3723
rect 55965 3689 55999 3723
rect 57253 3689 57287 3723
rect 57805 3689 57839 3723
rect 1961 3621 1995 3655
rect 2973 3621 3007 3655
rect 6653 3621 6687 3655
rect 40049 3621 40083 3655
rect 45201 3621 45235 3655
rect 51457 3621 51491 3655
rect 1777 3553 1811 3587
rect 2605 3553 2639 3587
rect 5273 3553 5307 3587
rect 9045 3553 9079 3587
rect 10793 3553 10827 3587
rect 10977 3553 11011 3587
rect 11529 3553 11563 3587
rect 16865 3553 16899 3587
rect 25421 3553 25455 3587
rect 40417 3553 40451 3587
rect 46581 3553 46615 3587
rect 49433 3553 49467 3587
rect 53297 3553 53331 3587
rect 56609 3553 56643 3587
rect 2053 3485 2087 3519
rect 2789 3485 2823 3519
rect 4169 3485 4203 3519
rect 4261 3485 4295 3519
rect 5540 3485 5574 3519
rect 7665 3485 7699 3519
rect 7941 3485 7975 3519
rect 9321 3485 9355 3519
rect 10425 3485 10459 3519
rect 10609 3485 10643 3519
rect 13369 3485 13403 3519
rect 13553 3485 13587 3519
rect 14473 3485 14507 3519
rect 14565 3485 14599 3519
rect 14657 3485 14691 3519
rect 14841 3485 14875 3519
rect 16037 3485 16071 3519
rect 16313 3485 16347 3519
rect 16773 3485 16807 3519
rect 17049 3485 17083 3519
rect 17969 3485 18003 3519
rect 18429 3485 18463 3519
rect 19257 3485 19291 3519
rect 19533 3485 19567 3519
rect 20821 3485 20855 3519
rect 23305 3485 23339 3519
rect 24961 3485 24995 3519
rect 27445 3485 27479 3519
rect 29561 3485 29595 3519
rect 31217 3485 31251 3519
rect 33977 3485 34011 3519
rect 34713 3485 34747 3519
rect 34897 3485 34931 3519
rect 35541 3485 35575 3519
rect 37473 3485 37507 3519
rect 37933 3485 37967 3519
rect 38301 3485 38335 3519
rect 38853 3485 38887 3519
rect 40233 3485 40267 3519
rect 40969 3485 41003 3519
rect 41245 3485 41279 3519
rect 41889 3485 41923 3519
rect 42625 3485 42659 3519
rect 42809 3485 42843 3519
rect 42901 3485 42935 3519
rect 42993 3485 43027 3519
rect 43729 3485 43763 3519
rect 43913 3485 43947 3519
rect 44005 3485 44039 3519
rect 44097 3485 44131 3519
rect 47041 3485 47075 3519
rect 50169 3485 50203 3519
rect 53021 3485 53055 3519
rect 53757 3485 53791 3519
rect 54401 3485 54435 3519
rect 54585 3485 54619 3519
rect 55321 3485 55355 3519
rect 2513 3417 2547 3451
rect 3801 3417 3835 3451
rect 11796 3417 11830 3451
rect 14197 3417 14231 3451
rect 15853 3417 15887 3451
rect 25666 3417 25700 3451
rect 27997 3417 28031 3451
rect 28181 3417 28215 3451
rect 28825 3417 28859 3451
rect 29009 3417 29043 3451
rect 35808 3417 35842 3451
rect 40509 3417 40543 3451
rect 43269 3417 43303 3451
rect 46314 3417 46348 3451
rect 49166 3417 49200 3451
rect 7389 3349 7423 3383
rect 12909 3349 12943 3383
rect 16221 3349 16255 3383
rect 17233 3349 17267 3383
rect 18613 3349 18647 3383
rect 22109 3349 22143 3383
rect 23121 3349 23155 3383
rect 29791 3349 29825 3383
rect 36921 3349 36955 3383
rect 38669 3349 38703 3383
rect 41061 3349 41095 3383
rect 41429 3349 41463 3383
rect 44373 3349 44407 3383
rect 48053 3349 48087 3383
rect 1501 3145 1535 3179
rect 3065 3145 3099 3179
rect 3985 3145 4019 3179
rect 6469 3145 6503 3179
rect 7113 3145 7147 3179
rect 12449 3145 12483 3179
rect 16865 3145 16899 3179
rect 17233 3145 17267 3179
rect 22201 3145 22235 3179
rect 25237 3145 25271 3179
rect 26433 3145 26467 3179
rect 33793 3145 33827 3179
rect 36737 3145 36771 3179
rect 37289 3145 37323 3179
rect 40877 3145 40911 3179
rect 41245 3145 41279 3179
rect 52929 3145 52963 3179
rect 57897 3145 57931 3179
rect 2697 3077 2731 3111
rect 3709 3077 3743 3111
rect 4077 3077 4111 3111
rect 6929 3077 6963 3111
rect 7665 3077 7699 3111
rect 15209 3077 15243 3111
rect 15485 3077 15519 3111
rect 15945 3077 15979 3111
rect 18889 3077 18923 3111
rect 19073 3077 19107 3111
rect 19533 3077 19567 3111
rect 21281 3077 21315 3111
rect 27813 3077 27847 3111
rect 30389 3077 30423 3111
rect 31493 3077 31527 3111
rect 32505 3077 32539 3111
rect 43821 3077 43855 3111
rect 49258 3077 49292 3111
rect 2237 3009 2271 3043
rect 2881 3009 2915 3043
rect 2973 3009 3007 3043
rect 3893 3009 3927 3043
rect 4261 3009 4295 3043
rect 4905 3009 4939 3043
rect 5089 3009 5123 3043
rect 5825 3009 5859 3043
rect 7205 3009 7239 3043
rect 8769 3009 8803 3043
rect 9045 3009 9079 3043
rect 9505 3009 9539 3043
rect 11529 3009 11563 3043
rect 11805 3009 11839 3043
rect 13277 3009 13311 3043
rect 13737 3009 13771 3043
rect 14473 3009 14507 3043
rect 15393 3009 15427 3043
rect 17049 3009 17083 3043
rect 17325 3009 17359 3043
rect 18153 3009 18187 3043
rect 21833 3009 21867 3043
rect 22017 3009 22051 3043
rect 23029 3009 23063 3043
rect 23765 3009 23799 3043
rect 25513 3009 25547 3043
rect 25605 3009 25639 3043
rect 25697 3009 25731 3043
rect 25881 3009 25915 3043
rect 27721 3009 27755 3043
rect 27905 3009 27939 3043
rect 29285 3009 29319 3043
rect 30849 3009 30883 3043
rect 31033 3012 31067 3046
rect 31128 3012 31162 3046
rect 31217 3009 31251 3043
rect 34713 3009 34747 3043
rect 36001 3009 36035 3043
rect 37473 3009 37507 3043
rect 37657 3009 37691 3043
rect 37749 3009 37783 3043
rect 40141 3009 40175 3043
rect 40785 3009 40819 3043
rect 41061 3009 41095 3043
rect 41705 3009 41739 3043
rect 43177 3009 43211 3043
rect 43356 3009 43390 3043
rect 43456 3009 43490 3043
rect 43591 3009 43625 3043
rect 44281 3009 44315 3043
rect 49525 3009 49559 3043
rect 51273 3009 51307 3043
rect 52929 3009 52963 3043
rect 54125 3009 54159 3043
rect 54769 3009 54803 3043
rect 9781 2941 9815 2975
rect 11621 2941 11655 2975
rect 24777 2941 24811 2975
rect 29009 2941 29043 2975
rect 34989 2941 35023 2975
rect 47593 2941 47627 2975
rect 50629 2941 50663 2975
rect 53481 2941 53515 2975
rect 56701 2941 56735 2975
rect 2053 2873 2087 2907
rect 7665 2873 7699 2907
rect 11989 2873 12023 2907
rect 13921 2873 13955 2907
rect 14657 2873 14691 2907
rect 15945 2873 15979 2907
rect 23581 2873 23615 2907
rect 28365 2873 28399 2907
rect 38209 2873 38243 2907
rect 42441 2873 42475 2907
rect 48145 2873 48179 2907
rect 51917 2873 51951 2907
rect 55413 2873 55447 2907
rect 3249 2805 3283 2839
rect 5641 2805 5675 2839
rect 10977 2805 11011 2839
rect 11529 2805 11563 2839
rect 13093 2805 13127 2839
rect 17969 2805 18003 2839
rect 22845 2805 22879 2839
rect 26985 2805 27019 2839
rect 38853 2805 38887 2839
rect 39497 2805 39531 2839
rect 44925 2805 44959 2839
rect 45569 2805 45603 2839
rect 46213 2805 46247 2839
rect 46857 2805 46891 2839
rect 49985 2805 50019 2839
rect 56057 2805 56091 2839
rect 1869 2601 1903 2635
rect 3065 2601 3099 2635
rect 4445 2601 4479 2635
rect 6837 2601 6871 2635
rect 17877 2601 17911 2635
rect 31125 2601 31159 2635
rect 33977 2601 34011 2635
rect 35357 2601 35391 2635
rect 36737 2601 36771 2635
rect 47041 2601 47075 2635
rect 57253 2601 57287 2635
rect 6653 2533 6687 2567
rect 17049 2533 17083 2567
rect 24501 2533 24535 2567
rect 25789 2533 25823 2567
rect 29009 2533 29043 2567
rect 32137 2533 32171 2567
rect 41153 2533 41187 2567
rect 42441 2533 42475 2567
rect 46305 2533 46339 2567
rect 56609 2533 56643 2567
rect 2237 2465 2271 2499
rect 7021 2465 7055 2499
rect 9321 2465 9355 2499
rect 9413 2465 9447 2499
rect 18429 2465 18463 2499
rect 27721 2465 27755 2499
rect 30021 2465 30055 2499
rect 34713 2465 34747 2499
rect 36001 2465 36035 2499
rect 38577 2465 38611 2499
rect 39221 2465 39255 2499
rect 47593 2465 47627 2499
rect 52101 2465 52135 2499
rect 55965 2465 55999 2499
rect 2053 2397 2087 2431
rect 2697 2397 2731 2431
rect 2881 2397 2915 2431
rect 3985 2397 4019 2431
rect 5825 2397 5859 2431
rect 6837 2397 6871 2431
rect 7573 2397 7607 2431
rect 7849 2397 7883 2431
rect 9137 2397 9171 2431
rect 9229 2397 9263 2431
rect 10701 2397 10735 2431
rect 10977 2397 11011 2431
rect 11529 2397 11563 2431
rect 11805 2397 11839 2431
rect 13553 2397 13587 2431
rect 14381 2397 14415 2431
rect 15117 2397 15151 2431
rect 15853 2397 15887 2431
rect 17233 2397 17267 2431
rect 17693 2397 17727 2431
rect 18613 2397 18647 2431
rect 20269 2397 20303 2431
rect 20545 2397 20579 2431
rect 21281 2397 21315 2431
rect 21833 2397 21867 2431
rect 22017 2397 22051 2431
rect 22661 2397 22695 2431
rect 22845 2397 22879 2431
rect 22937 2397 22971 2431
rect 23765 2397 23799 2431
rect 24685 2397 24719 2431
rect 26433 2397 26467 2431
rect 26985 2397 27019 2431
rect 28365 2397 28399 2431
rect 30481 2397 30515 2431
rect 31309 2397 31343 2431
rect 31585 2397 31619 2431
rect 33241 2397 33275 2431
rect 33517 2397 33551 2431
rect 37289 2397 37323 2431
rect 37933 2397 37967 2431
rect 39865 2397 39899 2431
rect 40509 2397 40543 2431
rect 43085 2397 43119 2431
rect 43729 2397 43763 2431
rect 44373 2397 44407 2431
rect 45017 2397 45051 2431
rect 45661 2397 45695 2431
rect 48237 2397 48271 2431
rect 48881 2397 48915 2431
rect 49525 2397 49559 2431
rect 50169 2397 50203 2431
rect 50813 2397 50847 2431
rect 51457 2397 51491 2431
rect 52745 2397 52779 2431
rect 53389 2397 53423 2431
rect 54033 2397 54067 2431
rect 55321 2397 55355 2431
rect 5558 2329 5592 2363
rect 7113 2329 7147 2363
rect 8953 2329 8987 2363
rect 31493 2329 31527 2363
rect 13369 2261 13403 2295
rect 14565 2261 14599 2295
rect 15301 2261 15335 2295
rect 16037 2261 16071 2295
rect 19533 2261 19567 2295
rect 21097 2261 21131 2295
rect 22201 2261 22235 2295
rect 23581 2261 23615 2295
rect 41797 2261 41831 2295
rect 54677 2261 54711 2295
rect 57897 2261 57931 2295
<< metal1 >>
rect 1104 17434 58880 17456
rect 1104 17382 15398 17434
rect 15450 17382 15462 17434
rect 15514 17382 15526 17434
rect 15578 17382 15590 17434
rect 15642 17382 15654 17434
rect 15706 17382 29846 17434
rect 29898 17382 29910 17434
rect 29962 17382 29974 17434
rect 30026 17382 30038 17434
rect 30090 17382 30102 17434
rect 30154 17382 44294 17434
rect 44346 17382 44358 17434
rect 44410 17382 44422 17434
rect 44474 17382 44486 17434
rect 44538 17382 44550 17434
rect 44602 17382 58880 17434
rect 1104 17360 58880 17382
rect 4341 17187 4399 17193
rect 4341 17153 4353 17187
rect 4387 17184 4399 17187
rect 4430 17184 4436 17196
rect 4387 17156 4436 17184
rect 4387 17153 4399 17156
rect 4341 17147 4399 17153
rect 4430 17144 4436 17156
rect 4488 17144 4494 17196
rect 4890 17144 4896 17196
rect 4948 17184 4954 17196
rect 4985 17187 5043 17193
rect 4985 17184 4997 17187
rect 4948 17156 4997 17184
rect 4948 17144 4954 17156
rect 4985 17153 4997 17156
rect 5031 17153 5043 17187
rect 5810 17184 5816 17196
rect 5771 17156 5816 17184
rect 4985 17147 5043 17153
rect 5810 17144 5816 17156
rect 5868 17144 5874 17196
rect 7101 17187 7159 17193
rect 7101 17153 7113 17187
rect 7147 17184 7159 17187
rect 7190 17184 7196 17196
rect 7147 17156 7196 17184
rect 7147 17153 7159 17156
rect 7101 17147 7159 17153
rect 7190 17144 7196 17156
rect 7248 17144 7254 17196
rect 7561 17187 7619 17193
rect 7561 17153 7573 17187
rect 7607 17184 7619 17187
rect 7650 17184 7656 17196
rect 7607 17156 7656 17184
rect 7607 17153 7619 17156
rect 7561 17147 7619 17153
rect 7650 17144 7656 17156
rect 7708 17144 7714 17196
rect 8389 17187 8447 17193
rect 8389 17153 8401 17187
rect 8435 17184 8447 17187
rect 8570 17184 8576 17196
rect 8435 17156 8576 17184
rect 8435 17153 8447 17156
rect 8389 17147 8447 17153
rect 8570 17144 8576 17156
rect 8628 17144 8634 17196
rect 9030 17144 9036 17196
rect 9088 17184 9094 17196
rect 9125 17187 9183 17193
rect 9125 17184 9137 17187
rect 9088 17156 9137 17184
rect 9088 17144 9094 17156
rect 9125 17153 9137 17156
rect 9171 17153 9183 17187
rect 9125 17147 9183 17153
rect 9861 17187 9919 17193
rect 9861 17153 9873 17187
rect 9907 17184 9919 17187
rect 9950 17184 9956 17196
rect 9907 17156 9956 17184
rect 9907 17153 9919 17156
rect 9861 17147 9919 17153
rect 9950 17144 9956 17156
rect 10008 17144 10014 17196
rect 10410 17144 10416 17196
rect 10468 17184 10474 17196
rect 10505 17187 10563 17193
rect 10505 17184 10517 17187
rect 10468 17156 10517 17184
rect 10468 17144 10474 17156
rect 10505 17153 10517 17156
rect 10551 17153 10563 17187
rect 10505 17147 10563 17153
rect 11790 17144 11796 17196
rect 11848 17184 11854 17196
rect 11885 17187 11943 17193
rect 11885 17184 11897 17187
rect 11848 17156 11897 17184
rect 11848 17144 11854 17156
rect 11885 17153 11897 17156
rect 11931 17153 11943 17187
rect 11885 17147 11943 17153
rect 12621 17187 12679 17193
rect 12621 17153 12633 17187
rect 12667 17184 12679 17187
rect 12710 17184 12716 17196
rect 12667 17156 12716 17184
rect 12667 17153 12679 17156
rect 12621 17147 12679 17153
rect 12710 17144 12716 17156
rect 12768 17144 12774 17196
rect 13170 17144 13176 17196
rect 13228 17184 13234 17196
rect 13265 17187 13323 17193
rect 13265 17184 13277 17187
rect 13228 17156 13277 17184
rect 13228 17144 13234 17156
rect 13265 17153 13277 17156
rect 13311 17153 13323 17187
rect 13265 17147 13323 17153
rect 14550 17144 14556 17196
rect 14608 17184 14614 17196
rect 14645 17187 14703 17193
rect 14645 17184 14657 17187
rect 14608 17156 14657 17184
rect 14608 17144 14614 17156
rect 14645 17153 14657 17156
rect 14691 17153 14703 17187
rect 14645 17147 14703 17153
rect 15286 17144 15292 17196
rect 15344 17184 15350 17196
rect 15473 17187 15531 17193
rect 15473 17184 15485 17187
rect 15344 17156 15485 17184
rect 15344 17144 15350 17156
rect 15473 17153 15485 17156
rect 15519 17153 15531 17187
rect 15930 17184 15936 17196
rect 15891 17156 15936 17184
rect 15473 17147 15531 17153
rect 15930 17144 15936 17156
rect 15988 17144 15994 17196
rect 17221 17187 17279 17193
rect 17221 17153 17233 17187
rect 17267 17184 17279 17187
rect 17310 17184 17316 17196
rect 17267 17156 17316 17184
rect 17267 17153 17279 17156
rect 17221 17147 17279 17153
rect 17310 17144 17316 17156
rect 17368 17144 17374 17196
rect 18049 17187 18107 17193
rect 18049 17153 18061 17187
rect 18095 17184 18107 17187
rect 18230 17184 18236 17196
rect 18095 17156 18236 17184
rect 18095 17153 18107 17156
rect 18049 17147 18107 17153
rect 18230 17144 18236 17156
rect 18288 17144 18294 17196
rect 18690 17184 18696 17196
rect 18651 17156 18696 17184
rect 18690 17144 18696 17156
rect 18748 17144 18754 17196
rect 19521 17187 19579 17193
rect 19521 17153 19533 17187
rect 19567 17184 19579 17187
rect 19610 17184 19616 17196
rect 19567 17156 19616 17184
rect 19567 17153 19579 17156
rect 19521 17147 19579 17153
rect 19610 17144 19616 17156
rect 19668 17144 19674 17196
rect 20070 17144 20076 17196
rect 20128 17184 20134 17196
rect 20165 17187 20223 17193
rect 20165 17184 20177 17187
rect 20128 17156 20177 17184
rect 20128 17144 20134 17156
rect 20165 17153 20177 17156
rect 20211 17153 20223 17187
rect 20165 17147 20223 17153
rect 21269 17187 21327 17193
rect 21269 17153 21281 17187
rect 21315 17184 21327 17187
rect 21450 17184 21456 17196
rect 21315 17156 21456 17184
rect 21315 17153 21327 17156
rect 21269 17147 21327 17153
rect 21450 17144 21456 17156
rect 21508 17144 21514 17196
rect 22281 17187 22339 17193
rect 22281 17153 22293 17187
rect 22327 17184 22339 17187
rect 22370 17184 22376 17196
rect 22327 17156 22376 17184
rect 22327 17153 22339 17156
rect 22281 17147 22339 17153
rect 22370 17144 22376 17156
rect 22428 17144 22434 17196
rect 22830 17144 22836 17196
rect 22888 17184 22894 17196
rect 22925 17187 22983 17193
rect 22925 17184 22937 17187
rect 22888 17156 22937 17184
rect 22888 17144 22894 17156
rect 22925 17153 22937 17156
rect 22971 17153 22983 17187
rect 22925 17147 22983 17153
rect 23661 17187 23719 17193
rect 23661 17153 23673 17187
rect 23707 17184 23719 17187
rect 23750 17184 23756 17196
rect 23707 17156 23756 17184
rect 23707 17153 23719 17156
rect 23661 17147 23719 17153
rect 23750 17144 23756 17156
rect 23808 17144 23814 17196
rect 25130 17184 25136 17196
rect 25091 17156 25136 17184
rect 25130 17144 25136 17156
rect 25188 17144 25194 17196
rect 25590 17184 25596 17196
rect 25551 17156 25596 17184
rect 25590 17144 25596 17156
rect 25648 17144 25654 17196
rect 26421 17187 26479 17193
rect 26421 17153 26433 17187
rect 26467 17184 26479 17187
rect 26510 17184 26516 17196
rect 26467 17156 26516 17184
rect 26467 17153 26479 17156
rect 26421 17147 26479 17153
rect 26510 17144 26516 17156
rect 26568 17144 26574 17196
rect 27709 17187 27767 17193
rect 27709 17153 27721 17187
rect 27755 17184 27767 17187
rect 27890 17184 27896 17196
rect 27755 17156 27896 17184
rect 27755 17153 27767 17156
rect 27709 17147 27767 17153
rect 27890 17144 27896 17156
rect 27948 17144 27954 17196
rect 28350 17184 28356 17196
rect 28311 17156 28356 17184
rect 28350 17144 28356 17156
rect 28408 17144 28414 17196
rect 28997 17187 29055 17193
rect 28997 17153 29009 17187
rect 29043 17184 29055 17187
rect 29270 17184 29276 17196
rect 29043 17156 29276 17184
rect 29043 17153 29055 17156
rect 28997 17147 29055 17153
rect 29270 17144 29276 17156
rect 29328 17144 29334 17196
rect 29730 17144 29736 17196
rect 29788 17184 29794 17196
rect 29825 17187 29883 17193
rect 29825 17184 29837 17187
rect 29788 17156 29837 17184
rect 29788 17144 29794 17156
rect 29825 17153 29837 17156
rect 29871 17153 29883 17187
rect 29825 17147 29883 17153
rect 30561 17187 30619 17193
rect 30561 17153 30573 17187
rect 30607 17184 30619 17187
rect 30650 17184 30656 17196
rect 30607 17156 30656 17184
rect 30607 17153 30619 17156
rect 30561 17147 30619 17153
rect 30650 17144 30656 17156
rect 30708 17144 30714 17196
rect 31110 17144 31116 17196
rect 31168 17184 31174 17196
rect 31205 17187 31263 17193
rect 31205 17184 31217 17187
rect 31168 17156 31217 17184
rect 31168 17144 31174 17156
rect 31205 17153 31217 17156
rect 31251 17153 31263 17187
rect 31205 17147 31263 17153
rect 32030 17144 32036 17196
rect 32088 17184 32094 17196
rect 32125 17187 32183 17193
rect 32125 17184 32137 17187
rect 32088 17156 32137 17184
rect 32088 17144 32094 17156
rect 32125 17153 32137 17156
rect 32171 17153 32183 17187
rect 32125 17147 32183 17153
rect 32490 17144 32496 17196
rect 32548 17184 32554 17196
rect 32769 17187 32827 17193
rect 32769 17184 32781 17187
rect 32548 17156 32781 17184
rect 32548 17144 32554 17156
rect 32769 17153 32781 17156
rect 32815 17153 32827 17187
rect 32769 17147 32827 17153
rect 33410 17144 33416 17196
rect 33468 17184 33474 17196
rect 33505 17187 33563 17193
rect 33505 17184 33517 17187
rect 33468 17156 33517 17184
rect 33468 17144 33474 17156
rect 33505 17153 33517 17156
rect 33551 17153 33563 17187
rect 33505 17147 33563 17153
rect 33870 17144 33876 17196
rect 33928 17184 33934 17196
rect 34701 17187 34759 17193
rect 34701 17184 34713 17187
rect 33928 17156 34713 17184
rect 33928 17144 33934 17156
rect 34701 17153 34713 17156
rect 34747 17153 34759 17187
rect 34701 17147 34759 17153
rect 34790 17144 34796 17196
rect 34848 17184 34854 17196
rect 35345 17187 35403 17193
rect 35345 17184 35357 17187
rect 34848 17156 35357 17184
rect 34848 17144 34854 17156
rect 35345 17153 35357 17156
rect 35391 17153 35403 17187
rect 35345 17147 35403 17153
rect 36630 17144 36636 17196
rect 36688 17184 36694 17196
rect 37277 17187 37335 17193
rect 37277 17184 37289 17187
rect 36688 17156 37289 17184
rect 36688 17144 36694 17156
rect 37277 17153 37289 17156
rect 37323 17153 37335 17187
rect 37277 17147 37335 17153
rect 37550 17144 37556 17196
rect 37608 17184 37614 17196
rect 37921 17187 37979 17193
rect 37921 17184 37933 17187
rect 37608 17156 37933 17184
rect 37608 17144 37614 17156
rect 37921 17153 37933 17156
rect 37967 17153 37979 17187
rect 37921 17147 37979 17153
rect 38010 17144 38016 17196
rect 38068 17184 38074 17196
rect 38565 17187 38623 17193
rect 38565 17184 38577 17187
rect 38068 17156 38577 17184
rect 38068 17144 38074 17156
rect 38565 17153 38577 17156
rect 38611 17153 38623 17187
rect 38565 17147 38623 17153
rect 38930 17144 38936 17196
rect 38988 17184 38994 17196
rect 39853 17187 39911 17193
rect 39853 17184 39865 17187
rect 38988 17156 39865 17184
rect 38988 17144 38994 17156
rect 39853 17153 39865 17156
rect 39899 17153 39911 17187
rect 39853 17147 39911 17153
rect 40310 17144 40316 17196
rect 40368 17184 40374 17196
rect 40497 17187 40555 17193
rect 40497 17184 40509 17187
rect 40368 17156 40509 17184
rect 40368 17144 40374 17156
rect 40497 17153 40509 17156
rect 40543 17153 40555 17187
rect 40497 17147 40555 17153
rect 40770 17144 40776 17196
rect 40828 17184 40834 17196
rect 41141 17187 41199 17193
rect 41141 17184 41153 17187
rect 40828 17156 41153 17184
rect 40828 17144 40834 17156
rect 41141 17153 41153 17156
rect 41187 17153 41199 17187
rect 41141 17147 41199 17153
rect 41690 17144 41696 17196
rect 41748 17184 41754 17196
rect 42429 17187 42487 17193
rect 42429 17184 42441 17187
rect 41748 17156 42441 17184
rect 41748 17144 41754 17156
rect 42429 17153 42441 17156
rect 42475 17153 42487 17187
rect 42429 17147 42487 17153
rect 43070 17144 43076 17196
rect 43128 17184 43134 17196
rect 43717 17187 43775 17193
rect 43717 17184 43729 17187
rect 43128 17156 43729 17184
rect 43128 17144 43134 17156
rect 43717 17153 43729 17156
rect 43763 17153 43775 17187
rect 43717 17147 43775 17153
rect 44634 17144 44640 17196
rect 44692 17184 44698 17196
rect 45005 17187 45063 17193
rect 45005 17184 45017 17187
rect 44692 17156 45017 17184
rect 44692 17144 44698 17156
rect 45005 17153 45017 17156
rect 45051 17153 45063 17187
rect 45005 17147 45063 17153
rect 45830 17144 45836 17196
rect 45888 17184 45894 17196
rect 46293 17187 46351 17193
rect 46293 17184 46305 17187
rect 45888 17156 46305 17184
rect 45888 17144 45894 17156
rect 46293 17153 46305 17156
rect 46339 17153 46351 17187
rect 46293 17147 46351 17153
rect 47210 17144 47216 17196
rect 47268 17184 47274 17196
rect 47581 17187 47639 17193
rect 47581 17184 47593 17187
rect 47268 17156 47593 17184
rect 47268 17144 47274 17156
rect 47581 17153 47593 17156
rect 47627 17153 47639 17187
rect 47581 17147 47639 17153
rect 47670 17144 47676 17196
rect 47728 17184 47734 17196
rect 48225 17187 48283 17193
rect 48225 17184 48237 17187
rect 47728 17156 48237 17184
rect 47728 17144 47734 17156
rect 48225 17153 48237 17156
rect 48271 17153 48283 17187
rect 48225 17147 48283 17153
rect 48590 17144 48596 17196
rect 48648 17184 48654 17196
rect 48869 17187 48927 17193
rect 48869 17184 48881 17187
rect 48648 17156 48881 17184
rect 48648 17144 48654 17156
rect 48869 17153 48881 17156
rect 48915 17153 48927 17187
rect 48869 17147 48927 17153
rect 49970 17144 49976 17196
rect 50028 17184 50034 17196
rect 50157 17187 50215 17193
rect 50157 17184 50169 17187
rect 50028 17156 50169 17184
rect 50028 17144 50034 17156
rect 50157 17153 50169 17156
rect 50203 17153 50215 17187
rect 50157 17147 50215 17153
rect 50430 17144 50436 17196
rect 50488 17184 50494 17196
rect 50801 17187 50859 17193
rect 50801 17184 50813 17187
rect 50488 17156 50813 17184
rect 50488 17144 50494 17156
rect 50801 17153 50813 17156
rect 50847 17153 50859 17187
rect 50801 17147 50859 17153
rect 51350 17144 51356 17196
rect 51408 17184 51414 17196
rect 51445 17187 51503 17193
rect 51445 17184 51457 17187
rect 51408 17156 51457 17184
rect 51408 17144 51414 17156
rect 51445 17153 51457 17156
rect 51491 17153 51503 17187
rect 51445 17147 51503 17153
rect 51810 17144 51816 17196
rect 51868 17184 51874 17196
rect 52733 17187 52791 17193
rect 52733 17184 52745 17187
rect 51868 17156 52745 17184
rect 51868 17144 51874 17156
rect 52733 17153 52745 17156
rect 52779 17153 52791 17187
rect 52733 17147 52791 17153
rect 53190 17144 53196 17196
rect 53248 17184 53254 17196
rect 54021 17187 54079 17193
rect 54021 17184 54033 17187
rect 53248 17156 54033 17184
rect 53248 17144 53254 17156
rect 54021 17153 54033 17156
rect 54067 17153 54079 17187
rect 54021 17147 54079 17153
rect 54570 17144 54576 17196
rect 54628 17184 54634 17196
rect 55309 17187 55367 17193
rect 55309 17184 55321 17187
rect 54628 17156 55321 17184
rect 54628 17144 54634 17156
rect 55309 17153 55321 17156
rect 55355 17153 55367 17187
rect 55309 17147 55367 17153
rect 55490 17144 55496 17196
rect 55548 17184 55554 17196
rect 55953 17187 56011 17193
rect 55953 17184 55965 17187
rect 55548 17156 55965 17184
rect 55548 17144 55554 17156
rect 55953 17153 55965 17156
rect 55999 17153 56011 17187
rect 55953 17147 56011 17153
rect 56042 17144 56048 17196
rect 56100 17184 56106 17196
rect 56597 17187 56655 17193
rect 56597 17184 56609 17187
rect 56100 17156 56609 17184
rect 56100 17144 56106 17156
rect 56597 17153 56609 17156
rect 56643 17153 56655 17187
rect 56597 17147 56655 17153
rect 35250 17076 35256 17128
rect 35308 17116 35314 17128
rect 35989 17119 36047 17125
rect 35989 17116 36001 17119
rect 35308 17088 36001 17116
rect 35308 17076 35314 17088
rect 35989 17085 36001 17088
rect 36035 17085 36047 17119
rect 35989 17079 36047 17085
rect 44910 17076 44916 17128
rect 44968 17116 44974 17128
rect 45649 17119 45707 17125
rect 45649 17116 45661 17119
rect 44968 17088 45661 17116
rect 44968 17076 44974 17088
rect 45649 17085 45661 17088
rect 45695 17085 45707 17119
rect 45649 17079 45707 17085
rect 42150 17008 42156 17060
rect 42208 17048 42214 17060
rect 43073 17051 43131 17057
rect 43073 17048 43085 17051
rect 42208 17020 43085 17048
rect 42208 17008 42214 17020
rect 43073 17017 43085 17020
rect 43119 17017 43131 17051
rect 43073 17011 43131 17017
rect 52730 17008 52736 17060
rect 52788 17048 52794 17060
rect 53377 17051 53435 17057
rect 53377 17048 53389 17051
rect 52788 17020 53389 17048
rect 52788 17008 52794 17020
rect 53377 17017 53389 17020
rect 53423 17017 53435 17051
rect 53377 17011 53435 17017
rect 1104 16890 58880 16912
rect 1104 16838 8174 16890
rect 8226 16838 8238 16890
rect 8290 16838 8302 16890
rect 8354 16838 8366 16890
rect 8418 16838 8430 16890
rect 8482 16838 22622 16890
rect 22674 16838 22686 16890
rect 22738 16838 22750 16890
rect 22802 16838 22814 16890
rect 22866 16838 22878 16890
rect 22930 16838 37070 16890
rect 37122 16838 37134 16890
rect 37186 16838 37198 16890
rect 37250 16838 37262 16890
rect 37314 16838 37326 16890
rect 37378 16838 51518 16890
rect 51570 16838 51582 16890
rect 51634 16838 51646 16890
rect 51698 16838 51710 16890
rect 51762 16838 51774 16890
rect 51826 16838 58880 16890
rect 1104 16816 58880 16838
rect 6270 16736 6276 16788
rect 6328 16776 6334 16788
rect 6365 16779 6423 16785
rect 6365 16776 6377 16779
rect 6328 16748 6377 16776
rect 6328 16736 6334 16748
rect 6365 16745 6377 16748
rect 6411 16745 6423 16779
rect 6365 16739 6423 16745
rect 11330 16736 11336 16788
rect 11388 16776 11394 16788
rect 11425 16779 11483 16785
rect 11425 16776 11437 16779
rect 11388 16748 11437 16776
rect 11388 16736 11394 16748
rect 11425 16745 11437 16748
rect 11471 16745 11483 16779
rect 11425 16739 11483 16745
rect 14090 16736 14096 16788
rect 14148 16776 14154 16788
rect 14185 16779 14243 16785
rect 14185 16776 14197 16779
rect 14148 16748 14197 16776
rect 14148 16736 14154 16748
rect 14185 16745 14197 16748
rect 14231 16745 14243 16779
rect 14185 16739 14243 16745
rect 16850 16736 16856 16788
rect 16908 16776 16914 16788
rect 16945 16779 17003 16785
rect 16945 16776 16957 16779
rect 16908 16748 16957 16776
rect 16908 16736 16914 16748
rect 16945 16745 16957 16748
rect 16991 16745 17003 16779
rect 16945 16739 17003 16745
rect 20990 16736 20996 16788
rect 21048 16776 21054 16788
rect 21085 16779 21143 16785
rect 21085 16776 21097 16779
rect 21048 16748 21097 16776
rect 21048 16736 21054 16748
rect 21085 16745 21097 16748
rect 21131 16745 21143 16779
rect 21085 16739 21143 16745
rect 24210 16736 24216 16788
rect 24268 16776 24274 16788
rect 24397 16779 24455 16785
rect 24397 16776 24409 16779
rect 24268 16748 24409 16776
rect 24268 16736 24274 16748
rect 24397 16745 24409 16748
rect 24443 16745 24455 16779
rect 24397 16739 24455 16745
rect 26970 16736 26976 16788
rect 27028 16776 27034 16788
rect 27065 16779 27123 16785
rect 27065 16776 27077 16779
rect 27028 16748 27077 16776
rect 27028 16736 27034 16748
rect 27065 16745 27077 16748
rect 27111 16745 27123 16779
rect 27065 16739 27123 16745
rect 36170 16736 36176 16788
rect 36228 16776 36234 16788
rect 36265 16779 36323 16785
rect 36265 16776 36277 16779
rect 36228 16748 36277 16776
rect 36228 16736 36234 16748
rect 36265 16745 36277 16748
rect 36311 16745 36323 16779
rect 36265 16739 36323 16745
rect 39390 16736 39396 16788
rect 39448 16776 39454 16788
rect 39853 16779 39911 16785
rect 39853 16776 39865 16779
rect 39448 16748 39865 16776
rect 39448 16736 39454 16748
rect 39853 16745 39865 16748
rect 39899 16745 39911 16779
rect 39853 16739 39911 16745
rect 43530 16736 43536 16788
rect 43588 16776 43594 16788
rect 43625 16779 43683 16785
rect 43625 16776 43637 16779
rect 43588 16748 43637 16776
rect 43588 16736 43594 16748
rect 43625 16745 43637 16748
rect 43671 16745 43683 16779
rect 43625 16739 43683 16745
rect 46290 16736 46296 16788
rect 46348 16776 46354 16788
rect 46385 16779 46443 16785
rect 46385 16776 46397 16779
rect 46348 16748 46397 16776
rect 46348 16736 46354 16748
rect 46385 16745 46397 16748
rect 46431 16745 46443 16779
rect 46385 16739 46443 16745
rect 49050 16736 49056 16788
rect 49108 16776 49114 16788
rect 49145 16779 49203 16785
rect 49145 16776 49157 16779
rect 49108 16748 49157 16776
rect 49108 16736 49114 16748
rect 49145 16745 49157 16748
rect 49191 16745 49203 16779
rect 49145 16739 49203 16745
rect 54110 16736 54116 16788
rect 54168 16776 54174 16788
rect 54205 16779 54263 16785
rect 54205 16776 54217 16779
rect 54168 16748 54217 16776
rect 54168 16736 54174 16748
rect 54205 16745 54217 16748
rect 54251 16745 54263 16779
rect 54205 16739 54263 16745
rect 1104 16346 58880 16368
rect 1104 16294 15398 16346
rect 15450 16294 15462 16346
rect 15514 16294 15526 16346
rect 15578 16294 15590 16346
rect 15642 16294 15654 16346
rect 15706 16294 29846 16346
rect 29898 16294 29910 16346
rect 29962 16294 29974 16346
rect 30026 16294 30038 16346
rect 30090 16294 30102 16346
rect 30154 16294 44294 16346
rect 44346 16294 44358 16346
rect 44410 16294 44422 16346
rect 44474 16294 44486 16346
rect 44538 16294 44550 16346
rect 44602 16294 58880 16346
rect 1104 16272 58880 16294
rect 1104 15802 58880 15824
rect 1104 15750 8174 15802
rect 8226 15750 8238 15802
rect 8290 15750 8302 15802
rect 8354 15750 8366 15802
rect 8418 15750 8430 15802
rect 8482 15750 22622 15802
rect 22674 15750 22686 15802
rect 22738 15750 22750 15802
rect 22802 15750 22814 15802
rect 22866 15750 22878 15802
rect 22930 15750 37070 15802
rect 37122 15750 37134 15802
rect 37186 15750 37198 15802
rect 37250 15750 37262 15802
rect 37314 15750 37326 15802
rect 37378 15750 51518 15802
rect 51570 15750 51582 15802
rect 51634 15750 51646 15802
rect 51698 15750 51710 15802
rect 51762 15750 51774 15802
rect 51826 15750 58880 15802
rect 1104 15728 58880 15750
rect 1104 15258 58880 15280
rect 1104 15206 15398 15258
rect 15450 15206 15462 15258
rect 15514 15206 15526 15258
rect 15578 15206 15590 15258
rect 15642 15206 15654 15258
rect 15706 15206 29846 15258
rect 29898 15206 29910 15258
rect 29962 15206 29974 15258
rect 30026 15206 30038 15258
rect 30090 15206 30102 15258
rect 30154 15206 44294 15258
rect 44346 15206 44358 15258
rect 44410 15206 44422 15258
rect 44474 15206 44486 15258
rect 44538 15206 44550 15258
rect 44602 15206 58880 15258
rect 1104 15184 58880 15206
rect 1104 14714 58880 14736
rect 1104 14662 8174 14714
rect 8226 14662 8238 14714
rect 8290 14662 8302 14714
rect 8354 14662 8366 14714
rect 8418 14662 8430 14714
rect 8482 14662 22622 14714
rect 22674 14662 22686 14714
rect 22738 14662 22750 14714
rect 22802 14662 22814 14714
rect 22866 14662 22878 14714
rect 22930 14662 37070 14714
rect 37122 14662 37134 14714
rect 37186 14662 37198 14714
rect 37250 14662 37262 14714
rect 37314 14662 37326 14714
rect 37378 14662 51518 14714
rect 51570 14662 51582 14714
rect 51634 14662 51646 14714
rect 51698 14662 51710 14714
rect 51762 14662 51774 14714
rect 51826 14662 58880 14714
rect 1104 14640 58880 14662
rect 1104 14170 58880 14192
rect 1104 14118 15398 14170
rect 15450 14118 15462 14170
rect 15514 14118 15526 14170
rect 15578 14118 15590 14170
rect 15642 14118 15654 14170
rect 15706 14118 29846 14170
rect 29898 14118 29910 14170
rect 29962 14118 29974 14170
rect 30026 14118 30038 14170
rect 30090 14118 30102 14170
rect 30154 14118 44294 14170
rect 44346 14118 44358 14170
rect 44410 14118 44422 14170
rect 44474 14118 44486 14170
rect 44538 14118 44550 14170
rect 44602 14118 58880 14170
rect 1104 14096 58880 14118
rect 17405 13923 17463 13929
rect 17405 13889 17417 13923
rect 17451 13920 17463 13923
rect 20254 13920 20260 13932
rect 17451 13892 20260 13920
rect 17451 13889 17463 13892
rect 17405 13883 17463 13889
rect 20254 13880 20260 13892
rect 20312 13880 20318 13932
rect 3142 13812 3148 13864
rect 3200 13852 3206 13864
rect 3329 13855 3387 13861
rect 3329 13852 3341 13855
rect 3200 13824 3341 13852
rect 3200 13812 3206 13824
rect 3329 13821 3341 13824
rect 3375 13821 3387 13855
rect 13354 13852 13360 13864
rect 13315 13824 13360 13852
rect 3329 13815 3387 13821
rect 13354 13812 13360 13824
rect 13412 13812 13418 13864
rect 14001 13855 14059 13861
rect 14001 13821 14013 13855
rect 14047 13852 14059 13855
rect 25406 13852 25412 13864
rect 14047 13824 25412 13852
rect 14047 13821 14059 13824
rect 14001 13815 14059 13821
rect 25406 13812 25412 13824
rect 25464 13812 25470 13864
rect 1104 13626 58880 13648
rect 1104 13574 8174 13626
rect 8226 13574 8238 13626
rect 8290 13574 8302 13626
rect 8354 13574 8366 13626
rect 8418 13574 8430 13626
rect 8482 13574 22622 13626
rect 22674 13574 22686 13626
rect 22738 13574 22750 13626
rect 22802 13574 22814 13626
rect 22866 13574 22878 13626
rect 22930 13574 37070 13626
rect 37122 13574 37134 13626
rect 37186 13574 37198 13626
rect 37250 13574 37262 13626
rect 37314 13574 37326 13626
rect 37378 13574 51518 13626
rect 51570 13574 51582 13626
rect 51634 13574 51646 13626
rect 51698 13574 51710 13626
rect 51762 13574 51774 13626
rect 51826 13574 58880 13626
rect 1104 13552 58880 13574
rect 11422 13308 11428 13320
rect 11335 13280 11428 13308
rect 11422 13268 11428 13280
rect 11480 13308 11486 13320
rect 15194 13308 15200 13320
rect 11480 13280 15200 13308
rect 11480 13268 11486 13280
rect 15194 13268 15200 13280
rect 15252 13268 15258 13320
rect 22278 13308 22284 13320
rect 16546 13280 22284 13308
rect 5258 13200 5264 13252
rect 5316 13240 5322 13252
rect 6733 13243 6791 13249
rect 6733 13240 6745 13243
rect 5316 13212 6745 13240
rect 5316 13200 5322 13212
rect 6733 13209 6745 13212
rect 6779 13240 6791 13243
rect 9490 13240 9496 13252
rect 6779 13212 9496 13240
rect 6779 13209 6791 13212
rect 6733 13203 6791 13209
rect 9490 13200 9496 13212
rect 9548 13240 9554 13252
rect 12621 13243 12679 13249
rect 12621 13240 12633 13243
rect 9548 13212 12633 13240
rect 9548 13200 9554 13212
rect 12621 13209 12633 13212
rect 12667 13240 12679 13243
rect 12986 13240 12992 13252
rect 12667 13212 12992 13240
rect 12667 13209 12679 13212
rect 12621 13203 12679 13209
rect 12986 13200 12992 13212
rect 13044 13200 13050 13252
rect 16546 13240 16574 13280
rect 22278 13268 22284 13280
rect 22336 13268 22342 13320
rect 16942 13240 16948 13252
rect 14200 13212 16574 13240
rect 16855 13212 16948 13240
rect 14200 13184 14228 13212
rect 16942 13200 16948 13212
rect 17000 13240 17006 13252
rect 19702 13240 19708 13252
rect 17000 13212 19708 13240
rect 17000 13200 17006 13212
rect 19702 13200 19708 13212
rect 19760 13200 19766 13252
rect 1486 13132 1492 13184
rect 1544 13172 1550 13184
rect 2041 13175 2099 13181
rect 2041 13172 2053 13175
rect 1544 13144 2053 13172
rect 1544 13132 1550 13144
rect 2041 13141 2053 13144
rect 2087 13141 2099 13175
rect 2682 13172 2688 13184
rect 2643 13144 2688 13172
rect 2041 13135 2099 13141
rect 2682 13132 2688 13144
rect 2740 13132 2746 13184
rect 3234 13172 3240 13184
rect 3195 13144 3240 13172
rect 3234 13132 3240 13144
rect 3292 13132 3298 13184
rect 3786 13172 3792 13184
rect 3747 13144 3792 13172
rect 3786 13132 3792 13144
rect 3844 13132 3850 13184
rect 4982 13132 4988 13184
rect 5040 13172 5046 13184
rect 5169 13175 5227 13181
rect 5169 13172 5181 13175
rect 5040 13144 5181 13172
rect 5040 13132 5046 13144
rect 5169 13141 5181 13144
rect 5215 13141 5227 13175
rect 5169 13135 5227 13141
rect 5997 13175 6055 13181
rect 5997 13141 6009 13175
rect 6043 13172 6055 13175
rect 6270 13172 6276 13184
rect 6043 13144 6276 13172
rect 6043 13141 6055 13144
rect 5997 13135 6055 13141
rect 6270 13132 6276 13144
rect 6328 13132 6334 13184
rect 9401 13175 9459 13181
rect 9401 13141 9413 13175
rect 9447 13172 9459 13175
rect 9582 13172 9588 13184
rect 9447 13144 9588 13172
rect 9447 13141 9459 13144
rect 9401 13135 9459 13141
rect 9582 13132 9588 13144
rect 9640 13132 9646 13184
rect 9674 13132 9680 13184
rect 9732 13172 9738 13184
rect 9861 13175 9919 13181
rect 9861 13172 9873 13175
rect 9732 13144 9873 13172
rect 9732 13132 9738 13144
rect 9861 13141 9873 13144
rect 9907 13141 9919 13175
rect 9861 13135 9919 13141
rect 10873 13175 10931 13181
rect 10873 13141 10885 13175
rect 10919 13172 10931 13175
rect 11054 13172 11060 13184
rect 10919 13144 11060 13172
rect 10919 13141 10931 13144
rect 10873 13135 10931 13141
rect 11054 13132 11060 13144
rect 11112 13132 11118 13184
rect 11606 13132 11612 13184
rect 11664 13172 11670 13184
rect 11885 13175 11943 13181
rect 11885 13172 11897 13175
rect 11664 13144 11897 13172
rect 11664 13132 11670 13144
rect 11885 13141 11897 13144
rect 11931 13141 11943 13175
rect 11885 13135 11943 13141
rect 12894 13132 12900 13184
rect 12952 13172 12958 13184
rect 13173 13175 13231 13181
rect 13173 13172 13185 13175
rect 12952 13144 13185 13172
rect 12952 13132 12958 13144
rect 13173 13141 13185 13144
rect 13219 13141 13231 13175
rect 14182 13172 14188 13184
rect 14143 13144 14188 13172
rect 13173 13135 13231 13141
rect 14182 13132 14188 13144
rect 14240 13132 14246 13184
rect 15102 13172 15108 13184
rect 15063 13144 15108 13172
rect 15102 13132 15108 13144
rect 15160 13132 15166 13184
rect 15657 13175 15715 13181
rect 15657 13141 15669 13175
rect 15703 13172 15715 13175
rect 15838 13172 15844 13184
rect 15703 13144 15844 13172
rect 15703 13141 15715 13144
rect 15657 13135 15715 13141
rect 15838 13132 15844 13144
rect 15896 13132 15902 13184
rect 17770 13172 17776 13184
rect 17731 13144 17776 13172
rect 17770 13132 17776 13144
rect 17828 13132 17834 13184
rect 18046 13132 18052 13184
rect 18104 13172 18110 13184
rect 18233 13175 18291 13181
rect 18233 13172 18245 13175
rect 18104 13144 18245 13172
rect 18104 13132 18110 13144
rect 18233 13141 18245 13144
rect 18279 13141 18291 13175
rect 18233 13135 18291 13141
rect 22373 13175 22431 13181
rect 22373 13141 22385 13175
rect 22419 13172 22431 13175
rect 27798 13172 27804 13184
rect 22419 13144 27804 13172
rect 22419 13141 22431 13144
rect 22373 13135 22431 13141
rect 27798 13132 27804 13144
rect 27856 13132 27862 13184
rect 1104 13082 58880 13104
rect 1104 13030 15398 13082
rect 15450 13030 15462 13082
rect 15514 13030 15526 13082
rect 15578 13030 15590 13082
rect 15642 13030 15654 13082
rect 15706 13030 29846 13082
rect 29898 13030 29910 13082
rect 29962 13030 29974 13082
rect 30026 13030 30038 13082
rect 30090 13030 30102 13082
rect 30154 13030 44294 13082
rect 44346 13030 44358 13082
rect 44410 13030 44422 13082
rect 44474 13030 44486 13082
rect 44538 13030 44550 13082
rect 44602 13030 58880 13082
rect 1104 13008 58880 13030
rect 9490 12968 9496 12980
rect 9451 12940 9496 12968
rect 9490 12928 9496 12940
rect 9548 12928 9554 12980
rect 12986 12968 12992 12980
rect 12947 12940 12992 12968
rect 12986 12928 12992 12940
rect 13044 12928 13050 12980
rect 15102 12968 15108 12980
rect 13096 12940 15108 12968
rect 3970 12860 3976 12912
rect 4028 12900 4034 12912
rect 13096 12900 13124 12940
rect 15102 12928 15108 12940
rect 15160 12928 15166 12980
rect 15194 12928 15200 12980
rect 15252 12968 15258 12980
rect 17589 12971 17647 12977
rect 17589 12968 17601 12971
rect 15252 12940 17601 12968
rect 15252 12928 15258 12940
rect 17589 12937 17601 12940
rect 17635 12937 17647 12971
rect 17589 12931 17647 12937
rect 4028 12872 13124 12900
rect 13633 12903 13691 12909
rect 4028 12860 4034 12872
rect 13633 12869 13645 12903
rect 13679 12900 13691 12903
rect 18230 12900 18236 12912
rect 13679 12872 18236 12900
rect 13679 12869 13691 12872
rect 13633 12863 13691 12869
rect 18230 12860 18236 12872
rect 18288 12860 18294 12912
rect 21910 12900 21916 12912
rect 21823 12872 21916 12900
rect 21910 12860 21916 12872
rect 21968 12900 21974 12912
rect 25038 12900 25044 12912
rect 21968 12872 25044 12900
rect 21968 12860 21974 12872
rect 25038 12860 25044 12872
rect 25096 12860 25102 12912
rect 2501 12835 2559 12841
rect 2501 12801 2513 12835
rect 2547 12832 2559 12835
rect 5902 12832 5908 12844
rect 2547 12804 5908 12832
rect 2547 12801 2559 12804
rect 2501 12795 2559 12801
rect 5902 12792 5908 12804
rect 5960 12832 5966 12844
rect 12894 12832 12900 12844
rect 5960 12804 12900 12832
rect 5960 12792 5966 12804
rect 12894 12792 12900 12804
rect 12952 12792 12958 12844
rect 14553 12835 14611 12841
rect 14553 12801 14565 12835
rect 14599 12832 14611 12835
rect 15105 12835 15163 12841
rect 15105 12832 15117 12835
rect 14599 12804 15117 12832
rect 14599 12801 14611 12804
rect 14553 12795 14611 12801
rect 15105 12801 15117 12804
rect 15151 12832 15163 12835
rect 17218 12832 17224 12844
rect 15151 12804 17224 12832
rect 15151 12801 15163 12804
rect 15105 12795 15163 12801
rect 17218 12792 17224 12804
rect 17276 12792 17282 12844
rect 19337 12835 19395 12841
rect 19337 12801 19349 12835
rect 19383 12832 19395 12835
rect 22094 12832 22100 12844
rect 19383 12804 22100 12832
rect 19383 12801 19395 12804
rect 19337 12795 19395 12801
rect 22094 12792 22100 12804
rect 22152 12792 22158 12844
rect 4157 12767 4215 12773
rect 4157 12733 4169 12767
rect 4203 12764 4215 12767
rect 11422 12764 11428 12776
rect 4203 12736 11428 12764
rect 4203 12733 4215 12736
rect 4157 12727 4215 12733
rect 11422 12724 11428 12736
rect 11480 12724 11486 12776
rect 16942 12764 16948 12776
rect 13096 12736 16948 12764
rect 3142 12656 3148 12708
rect 3200 12696 3206 12708
rect 4617 12699 4675 12705
rect 4617 12696 4629 12699
rect 3200 12668 4629 12696
rect 3200 12656 3206 12668
rect 4617 12665 4629 12668
rect 4663 12665 4675 12699
rect 8389 12699 8447 12705
rect 8389 12696 8401 12699
rect 4617 12659 4675 12665
rect 6886 12668 8401 12696
rect 1946 12628 1952 12640
rect 1907 12600 1952 12628
rect 1946 12588 1952 12600
rect 2004 12588 2010 12640
rect 3053 12631 3111 12637
rect 3053 12597 3065 12631
rect 3099 12628 3111 12631
rect 3602 12628 3608 12640
rect 3099 12600 3608 12628
rect 3099 12597 3111 12600
rect 3053 12591 3111 12597
rect 3602 12588 3608 12600
rect 3660 12588 3666 12640
rect 5258 12628 5264 12640
rect 5219 12600 5264 12628
rect 5258 12588 5264 12600
rect 5316 12588 5322 12640
rect 5813 12631 5871 12637
rect 5813 12597 5825 12631
rect 5859 12628 5871 12631
rect 6457 12631 6515 12637
rect 6457 12628 6469 12631
rect 5859 12600 6469 12628
rect 5859 12597 5871 12600
rect 5813 12591 5871 12597
rect 6457 12597 6469 12600
rect 6503 12628 6515 12631
rect 6546 12628 6552 12640
rect 6503 12600 6552 12628
rect 6503 12597 6515 12600
rect 6457 12591 6515 12597
rect 6546 12588 6552 12600
rect 6604 12628 6610 12640
rect 6886 12628 6914 12668
rect 8389 12665 8401 12668
rect 8435 12696 8447 12699
rect 9214 12696 9220 12708
rect 8435 12668 9220 12696
rect 8435 12665 8447 12668
rect 8389 12659 8447 12665
rect 9214 12656 9220 12668
rect 9272 12696 9278 12708
rect 9272 12668 12296 12696
rect 9272 12656 9278 12668
rect 6604 12600 6914 12628
rect 6604 12588 6610 12600
rect 7006 12588 7012 12640
rect 7064 12628 7070 12640
rect 7837 12631 7895 12637
rect 7064 12600 7109 12628
rect 7064 12588 7070 12600
rect 7837 12597 7849 12631
rect 7883 12628 7895 12631
rect 7926 12628 7932 12640
rect 7883 12600 7932 12628
rect 7883 12597 7895 12600
rect 7837 12591 7895 12597
rect 7926 12588 7932 12600
rect 7984 12588 7990 12640
rect 8846 12628 8852 12640
rect 8807 12600 8852 12628
rect 8846 12588 8852 12600
rect 8904 12588 8910 12640
rect 10413 12631 10471 12637
rect 10413 12597 10425 12631
rect 10459 12628 10471 12631
rect 10962 12628 10968 12640
rect 10459 12600 10968 12628
rect 10459 12597 10471 12600
rect 10413 12591 10471 12597
rect 10962 12588 10968 12600
rect 11020 12588 11026 12640
rect 11609 12631 11667 12637
rect 11609 12597 11621 12631
rect 11655 12628 11667 12631
rect 11698 12628 11704 12640
rect 11655 12600 11704 12628
rect 11655 12597 11667 12600
rect 11609 12591 11667 12597
rect 11698 12588 11704 12600
rect 11756 12588 11762 12640
rect 12268 12637 12296 12668
rect 12253 12631 12311 12637
rect 12253 12597 12265 12631
rect 12299 12628 12311 12631
rect 13096 12628 13124 12736
rect 16942 12724 16948 12736
rect 17000 12724 17006 12776
rect 19058 12724 19064 12776
rect 19116 12764 19122 12776
rect 19797 12767 19855 12773
rect 19797 12764 19809 12767
rect 19116 12736 19809 12764
rect 19116 12724 19122 12736
rect 19797 12733 19809 12736
rect 19843 12733 19855 12767
rect 19797 12727 19855 12733
rect 21269 12767 21327 12773
rect 21269 12733 21281 12767
rect 21315 12764 21327 12767
rect 23658 12764 23664 12776
rect 21315 12736 23664 12764
rect 21315 12733 21327 12736
rect 21269 12727 21327 12733
rect 23658 12724 23664 12736
rect 23716 12724 23722 12776
rect 13170 12656 13176 12708
rect 13228 12696 13234 12708
rect 20070 12696 20076 12708
rect 13228 12668 20076 12696
rect 13228 12656 13234 12668
rect 20070 12656 20076 12668
rect 20128 12656 20134 12708
rect 22649 12699 22707 12705
rect 22649 12665 22661 12699
rect 22695 12696 22707 12699
rect 25130 12696 25136 12708
rect 22695 12668 25136 12696
rect 22695 12665 22707 12668
rect 22649 12659 22707 12665
rect 25130 12656 25136 12668
rect 25188 12656 25194 12708
rect 16114 12628 16120 12640
rect 12299 12600 13124 12628
rect 16075 12600 16120 12628
rect 12299 12597 12311 12600
rect 12253 12591 12311 12597
rect 16114 12588 16120 12600
rect 16172 12588 16178 12640
rect 17129 12631 17187 12637
rect 17129 12597 17141 12631
rect 17175 12628 17187 12631
rect 17218 12628 17224 12640
rect 17175 12600 17224 12628
rect 17175 12597 17187 12600
rect 17129 12591 17187 12597
rect 17218 12588 17224 12600
rect 17276 12588 17282 12640
rect 18230 12628 18236 12640
rect 18191 12600 18236 12628
rect 18230 12588 18236 12600
rect 18288 12588 18294 12640
rect 18785 12631 18843 12637
rect 18785 12597 18797 12631
rect 18831 12628 18843 12631
rect 19978 12628 19984 12640
rect 18831 12600 19984 12628
rect 18831 12597 18843 12600
rect 18785 12591 18843 12597
rect 19978 12588 19984 12600
rect 20036 12588 20042 12640
rect 20714 12628 20720 12640
rect 20675 12600 20720 12628
rect 20714 12588 20720 12600
rect 20772 12588 20778 12640
rect 23474 12628 23480 12640
rect 23435 12600 23480 12628
rect 23474 12588 23480 12600
rect 23532 12588 23538 12640
rect 23934 12628 23940 12640
rect 23895 12600 23940 12628
rect 23934 12588 23940 12600
rect 23992 12588 23998 12640
rect 1104 12538 58880 12560
rect 1104 12486 8174 12538
rect 8226 12486 8238 12538
rect 8290 12486 8302 12538
rect 8354 12486 8366 12538
rect 8418 12486 8430 12538
rect 8482 12486 22622 12538
rect 22674 12486 22686 12538
rect 22738 12486 22750 12538
rect 22802 12486 22814 12538
rect 22866 12486 22878 12538
rect 22930 12486 37070 12538
rect 37122 12486 37134 12538
rect 37186 12486 37198 12538
rect 37250 12486 37262 12538
rect 37314 12486 37326 12538
rect 37378 12486 51518 12538
rect 51570 12486 51582 12538
rect 51634 12486 51646 12538
rect 51698 12486 51710 12538
rect 51762 12486 51774 12538
rect 51826 12486 58880 12538
rect 1104 12464 58880 12486
rect 6546 12424 6552 12436
rect 6507 12396 6552 12424
rect 6546 12384 6552 12396
rect 6604 12384 6610 12436
rect 9214 12424 9220 12436
rect 9175 12396 9220 12424
rect 9214 12384 9220 12396
rect 9272 12384 9278 12436
rect 25130 12424 25136 12436
rect 25091 12396 25136 12424
rect 25130 12384 25136 12396
rect 25188 12384 25194 12436
rect 10962 12316 10968 12368
rect 11020 12356 11026 12368
rect 20162 12356 20168 12368
rect 11020 12328 20168 12356
rect 11020 12316 11026 12328
rect 20162 12316 20168 12328
rect 20220 12316 20226 12368
rect 1854 12180 1860 12232
rect 1912 12220 1918 12232
rect 2501 12223 2559 12229
rect 2501 12220 2513 12223
rect 1912 12192 2513 12220
rect 1912 12180 1918 12192
rect 2501 12189 2513 12192
rect 2547 12189 2559 12223
rect 3142 12220 3148 12232
rect 2501 12183 2559 12189
rect 2746 12192 3148 12220
rect 1489 12155 1547 12161
rect 1489 12121 1501 12155
rect 1535 12152 1547 12155
rect 2746 12152 2774 12192
rect 3142 12180 3148 12192
rect 3200 12220 3206 12232
rect 3326 12220 3332 12232
rect 3200 12192 3332 12220
rect 3200 12180 3206 12192
rect 3326 12180 3332 12192
rect 3384 12180 3390 12232
rect 5813 12223 5871 12229
rect 5813 12189 5825 12223
rect 5859 12220 5871 12223
rect 8570 12220 8576 12232
rect 5859 12192 8576 12220
rect 5859 12189 5871 12192
rect 5813 12183 5871 12189
rect 8570 12180 8576 12192
rect 8628 12180 8634 12232
rect 18049 12223 18107 12229
rect 18049 12189 18061 12223
rect 18095 12220 18107 12223
rect 19242 12220 19248 12232
rect 18095 12192 19248 12220
rect 18095 12189 18107 12192
rect 18049 12183 18107 12189
rect 19242 12180 19248 12192
rect 19300 12180 19306 12232
rect 20349 12223 20407 12229
rect 20349 12189 20361 12223
rect 20395 12220 20407 12223
rect 20530 12220 20536 12232
rect 20395 12192 20536 12220
rect 20395 12189 20407 12192
rect 20349 12183 20407 12189
rect 20530 12180 20536 12192
rect 20588 12180 20594 12232
rect 22462 12220 22468 12232
rect 21376 12192 22468 12220
rect 1535 12124 2774 12152
rect 4433 12155 4491 12161
rect 1535 12121 1547 12124
rect 1489 12115 1547 12121
rect 4433 12121 4445 12155
rect 4479 12152 4491 12155
rect 5902 12152 5908 12164
rect 4479 12124 5908 12152
rect 4479 12121 4491 12124
rect 4433 12115 4491 12121
rect 5902 12112 5908 12124
rect 5960 12112 5966 12164
rect 6914 12112 6920 12164
rect 6972 12152 6978 12164
rect 7745 12155 7803 12161
rect 7745 12152 7757 12155
rect 6972 12124 7757 12152
rect 6972 12112 6978 12124
rect 7745 12121 7757 12124
rect 7791 12152 7803 12155
rect 16301 12155 16359 12161
rect 7791 12124 10088 12152
rect 7791 12121 7803 12124
rect 7745 12115 7803 12121
rect 10060 12096 10088 12124
rect 16301 12121 16313 12155
rect 16347 12152 16359 12155
rect 17218 12152 17224 12164
rect 16347 12124 17224 12152
rect 16347 12121 16359 12124
rect 16301 12115 16359 12121
rect 17218 12112 17224 12124
rect 17276 12112 17282 12164
rect 20070 12112 20076 12164
rect 20128 12152 20134 12164
rect 21376 12161 21404 12192
rect 22462 12180 22468 12192
rect 22520 12180 22526 12232
rect 21361 12155 21419 12161
rect 21361 12152 21373 12155
rect 20128 12124 21373 12152
rect 20128 12112 20134 12124
rect 21361 12121 21373 12124
rect 21407 12121 21419 12155
rect 23109 12155 23167 12161
rect 23109 12152 23121 12155
rect 21361 12115 21419 12121
rect 22066 12124 23121 12152
rect 1670 12044 1676 12096
rect 1728 12084 1734 12096
rect 1949 12087 2007 12093
rect 1949 12084 1961 12087
rect 1728 12056 1961 12084
rect 1728 12044 1734 12056
rect 1949 12053 1961 12056
rect 1995 12053 2007 12087
rect 1949 12047 2007 12053
rect 2958 12044 2964 12096
rect 3016 12084 3022 12096
rect 3145 12087 3203 12093
rect 3145 12084 3157 12087
rect 3016 12056 3157 12084
rect 3016 12044 3022 12056
rect 3145 12053 3157 12056
rect 3191 12084 3203 12087
rect 3878 12084 3884 12096
rect 3191 12056 3884 12084
rect 3191 12053 3203 12056
rect 3145 12047 3203 12053
rect 3878 12044 3884 12056
rect 3936 12044 3942 12096
rect 5166 12084 5172 12096
rect 5127 12056 5172 12084
rect 5166 12044 5172 12056
rect 5224 12044 5230 12096
rect 7193 12087 7251 12093
rect 7193 12053 7205 12087
rect 7239 12084 7251 12087
rect 7834 12084 7840 12096
rect 7239 12056 7840 12084
rect 7239 12053 7251 12056
rect 7193 12047 7251 12053
rect 7834 12044 7840 12056
rect 7892 12044 7898 12096
rect 8389 12087 8447 12093
rect 8389 12053 8401 12087
rect 8435 12084 8447 12087
rect 8662 12084 8668 12096
rect 8435 12056 8668 12084
rect 8435 12053 8447 12056
rect 8389 12047 8447 12053
rect 8662 12044 8668 12056
rect 8720 12044 8726 12096
rect 10042 12084 10048 12096
rect 10003 12056 10048 12084
rect 10042 12044 10048 12056
rect 10100 12044 10106 12096
rect 10318 12044 10324 12096
rect 10376 12084 10382 12096
rect 10597 12087 10655 12093
rect 10597 12084 10609 12087
rect 10376 12056 10609 12084
rect 10376 12044 10382 12056
rect 10597 12053 10609 12056
rect 10643 12053 10655 12087
rect 10597 12047 10655 12053
rect 11146 12044 11152 12096
rect 11204 12084 11210 12096
rect 11241 12087 11299 12093
rect 11241 12084 11253 12087
rect 11204 12056 11253 12084
rect 11204 12044 11210 12056
rect 11241 12053 11253 12056
rect 11287 12053 11299 12087
rect 11241 12047 11299 12053
rect 12069 12087 12127 12093
rect 12069 12053 12081 12087
rect 12115 12084 12127 12087
rect 12434 12084 12440 12096
rect 12115 12056 12440 12084
rect 12115 12053 12127 12056
rect 12069 12047 12127 12053
rect 12434 12044 12440 12056
rect 12492 12044 12498 12096
rect 13081 12087 13139 12093
rect 13081 12053 13093 12087
rect 13127 12084 13139 12087
rect 13262 12084 13268 12096
rect 13127 12056 13268 12084
rect 13127 12053 13139 12056
rect 13081 12047 13139 12053
rect 13262 12044 13268 12056
rect 13320 12044 13326 12096
rect 14182 12084 14188 12096
rect 14143 12056 14188 12084
rect 14182 12044 14188 12056
rect 14240 12044 14246 12096
rect 14642 12044 14648 12096
rect 14700 12084 14706 12096
rect 15013 12087 15071 12093
rect 15013 12084 15025 12087
rect 14700 12056 15025 12084
rect 14700 12044 14706 12056
rect 15013 12053 15025 12056
rect 15059 12053 15071 12087
rect 15013 12047 15071 12053
rect 15657 12087 15715 12093
rect 15657 12053 15669 12087
rect 15703 12084 15715 12087
rect 16574 12084 16580 12096
rect 15703 12056 16580 12084
rect 15703 12053 15715 12056
rect 15657 12047 15715 12053
rect 16574 12044 16580 12056
rect 16632 12044 16638 12096
rect 16942 12044 16948 12096
rect 17000 12084 17006 12096
rect 17037 12087 17095 12093
rect 17037 12084 17049 12087
rect 17000 12056 17049 12084
rect 17000 12044 17006 12056
rect 17037 12053 17049 12056
rect 17083 12053 17095 12087
rect 18598 12084 18604 12096
rect 18559 12056 18604 12084
rect 17037 12047 17095 12053
rect 18598 12044 18604 12056
rect 18656 12044 18662 12096
rect 18782 12044 18788 12096
rect 18840 12084 18846 12096
rect 19245 12087 19303 12093
rect 19245 12084 19257 12087
rect 18840 12056 19257 12084
rect 18840 12044 18846 12056
rect 19245 12053 19257 12056
rect 19291 12053 19303 12087
rect 19245 12047 19303 12053
rect 19702 12044 19708 12096
rect 19760 12084 19766 12096
rect 20622 12084 20628 12096
rect 19760 12056 20628 12084
rect 19760 12044 19766 12056
rect 20622 12044 20628 12056
rect 20680 12084 20686 12096
rect 20901 12087 20959 12093
rect 20901 12084 20913 12087
rect 20680 12056 20913 12084
rect 20680 12044 20686 12056
rect 20901 12053 20913 12056
rect 20947 12084 20959 12087
rect 22066 12084 22094 12124
rect 23109 12121 23121 12124
rect 23155 12121 23167 12155
rect 23109 12115 23167 12121
rect 22278 12084 22284 12096
rect 20947 12056 22094 12084
rect 22239 12056 22284 12084
rect 20947 12053 20959 12056
rect 20901 12047 20959 12053
rect 22278 12044 22284 12056
rect 22336 12044 22342 12096
rect 23753 12087 23811 12093
rect 23753 12053 23765 12087
rect 23799 12084 23811 12087
rect 23842 12084 23848 12096
rect 23799 12056 23848 12084
rect 23799 12053 23811 12056
rect 23753 12047 23811 12053
rect 23842 12044 23848 12056
rect 23900 12044 23906 12096
rect 24026 12044 24032 12096
rect 24084 12084 24090 12096
rect 24397 12087 24455 12093
rect 24397 12084 24409 12087
rect 24084 12056 24409 12084
rect 24084 12044 24090 12056
rect 24397 12053 24409 12056
rect 24443 12053 24455 12087
rect 25590 12084 25596 12096
rect 25551 12056 25596 12084
rect 24397 12047 24455 12053
rect 25590 12044 25596 12056
rect 25648 12044 25654 12096
rect 36814 12044 36820 12096
rect 36872 12084 36878 12096
rect 37093 12087 37151 12093
rect 37093 12084 37105 12087
rect 36872 12056 37105 12084
rect 36872 12044 36878 12056
rect 37093 12053 37105 12056
rect 37139 12053 37151 12087
rect 37093 12047 37151 12053
rect 1104 11994 58880 12016
rect 1104 11942 15398 11994
rect 15450 11942 15462 11994
rect 15514 11942 15526 11994
rect 15578 11942 15590 11994
rect 15642 11942 15654 11994
rect 15706 11942 29846 11994
rect 29898 11942 29910 11994
rect 29962 11942 29974 11994
rect 30026 11942 30038 11994
rect 30090 11942 30102 11994
rect 30154 11942 44294 11994
rect 44346 11942 44358 11994
rect 44410 11942 44422 11994
rect 44474 11942 44486 11994
rect 44538 11942 44550 11994
rect 44602 11942 58880 11994
rect 1104 11920 58880 11942
rect 2958 11880 2964 11892
rect 2919 11852 2964 11880
rect 2958 11840 2964 11852
rect 3016 11840 3022 11892
rect 6914 11880 6920 11892
rect 6875 11852 6920 11880
rect 6914 11840 6920 11852
rect 6972 11840 6978 11892
rect 8570 11840 8576 11892
rect 8628 11880 8634 11892
rect 8665 11883 8723 11889
rect 8665 11880 8677 11883
rect 8628 11852 8677 11880
rect 8628 11840 8634 11852
rect 8665 11849 8677 11852
rect 8711 11849 8723 11883
rect 20070 11880 20076 11892
rect 20031 11852 20076 11880
rect 8665 11843 8723 11849
rect 20070 11840 20076 11852
rect 20128 11840 20134 11892
rect 22462 11840 22468 11892
rect 22520 11880 22526 11892
rect 23106 11880 23112 11892
rect 22520 11852 23112 11880
rect 22520 11840 22526 11852
rect 23106 11840 23112 11852
rect 23164 11840 23170 11892
rect 4246 11772 4252 11824
rect 4304 11812 4310 11824
rect 21910 11812 21916 11824
rect 4304 11784 21916 11812
rect 4304 11772 4310 11784
rect 21910 11772 21916 11784
rect 21968 11772 21974 11824
rect 11698 11704 11704 11756
rect 11756 11744 11762 11756
rect 45646 11744 45652 11756
rect 11756 11716 45652 11744
rect 11756 11704 11762 11716
rect 45646 11704 45652 11716
rect 45704 11704 45710 11756
rect 20990 11636 20996 11688
rect 21048 11676 21054 11688
rect 26237 11679 26295 11685
rect 26237 11676 26249 11679
rect 21048 11648 26249 11676
rect 21048 11636 21054 11648
rect 26237 11645 26249 11648
rect 26283 11676 26295 11679
rect 36538 11676 36544 11688
rect 26283 11648 36544 11676
rect 26283 11645 26295 11648
rect 26237 11639 26295 11645
rect 36538 11636 36544 11648
rect 36596 11636 36602 11688
rect 3418 11568 3424 11620
rect 3476 11608 3482 11620
rect 3513 11611 3571 11617
rect 3513 11608 3525 11611
rect 3476 11580 3525 11608
rect 3476 11568 3482 11580
rect 3513 11577 3525 11580
rect 3559 11608 3571 11611
rect 3602 11608 3608 11620
rect 3559 11580 3608 11608
rect 3559 11577 3571 11580
rect 3513 11571 3571 11577
rect 3602 11568 3608 11580
rect 3660 11608 3666 11620
rect 14550 11608 14556 11620
rect 3660 11580 14556 11608
rect 3660 11568 3666 11580
rect 14550 11568 14556 11580
rect 14608 11568 14614 11620
rect 16574 11568 16580 11620
rect 16632 11608 16638 11620
rect 18785 11611 18843 11617
rect 18785 11608 18797 11611
rect 16632 11580 18797 11608
rect 16632 11568 16638 11580
rect 18785 11577 18797 11580
rect 18831 11608 18843 11611
rect 23566 11608 23572 11620
rect 18831 11580 23572 11608
rect 18831 11577 18843 11580
rect 18785 11571 18843 11577
rect 23566 11568 23572 11580
rect 23624 11608 23630 11620
rect 23661 11611 23719 11617
rect 23661 11608 23673 11611
rect 23624 11580 23673 11608
rect 23624 11568 23630 11580
rect 23661 11577 23673 11580
rect 23707 11577 23719 11611
rect 23661 11571 23719 11577
rect 23750 11568 23756 11620
rect 23808 11608 23814 11620
rect 23808 11580 27384 11608
rect 23808 11568 23814 11580
rect 1578 11500 1584 11552
rect 1636 11540 1642 11552
rect 1857 11543 1915 11549
rect 1857 11540 1869 11543
rect 1636 11512 1869 11540
rect 1636 11500 1642 11512
rect 1857 11509 1869 11512
rect 1903 11509 1915 11543
rect 1857 11503 1915 11509
rect 4065 11543 4123 11549
rect 4065 11509 4077 11543
rect 4111 11540 4123 11543
rect 4338 11540 4344 11552
rect 4111 11512 4344 11540
rect 4111 11509 4123 11512
rect 4065 11503 4123 11509
rect 4338 11500 4344 11512
rect 4396 11540 4402 11552
rect 4890 11540 4896 11552
rect 4396 11512 4896 11540
rect 4396 11500 4402 11512
rect 4890 11500 4896 11512
rect 4948 11500 4954 11552
rect 5810 11540 5816 11552
rect 5771 11512 5816 11540
rect 5810 11500 5816 11512
rect 5868 11500 5874 11552
rect 7466 11500 7472 11552
rect 7524 11540 7530 11552
rect 7561 11543 7619 11549
rect 7561 11540 7573 11543
rect 7524 11512 7573 11540
rect 7524 11500 7530 11512
rect 7561 11509 7573 11512
rect 7607 11509 7619 11543
rect 7561 11503 7619 11509
rect 7650 11500 7656 11552
rect 7708 11540 7714 11552
rect 8113 11543 8171 11549
rect 8113 11540 8125 11543
rect 7708 11512 8125 11540
rect 7708 11500 7714 11512
rect 8113 11509 8125 11512
rect 8159 11509 8171 11543
rect 8113 11503 8171 11509
rect 9309 11543 9367 11549
rect 9309 11509 9321 11543
rect 9355 11540 9367 11543
rect 9674 11540 9680 11552
rect 9355 11512 9680 11540
rect 9355 11509 9367 11512
rect 9309 11503 9367 11509
rect 9674 11500 9680 11512
rect 9732 11500 9738 11552
rect 9861 11543 9919 11549
rect 9861 11509 9873 11543
rect 9907 11540 9919 11543
rect 10410 11540 10416 11552
rect 9907 11512 10416 11540
rect 9907 11509 9919 11512
rect 9861 11503 9919 11509
rect 10410 11500 10416 11512
rect 10468 11500 10474 11552
rect 10965 11543 11023 11549
rect 10965 11509 10977 11543
rect 11011 11540 11023 11543
rect 11793 11543 11851 11549
rect 11793 11540 11805 11543
rect 11011 11512 11805 11540
rect 11011 11509 11023 11512
rect 10965 11503 11023 11509
rect 11793 11509 11805 11512
rect 11839 11540 11851 11543
rect 12434 11540 12440 11552
rect 11839 11512 12440 11540
rect 11839 11509 11851 11512
rect 11793 11503 11851 11509
rect 12434 11500 12440 11512
rect 12492 11540 12498 11552
rect 12492 11512 12585 11540
rect 12492 11500 12498 11512
rect 12802 11500 12808 11552
rect 12860 11540 12866 11552
rect 12897 11543 12955 11549
rect 12897 11540 12909 11543
rect 12860 11512 12909 11540
rect 12860 11500 12866 11512
rect 12897 11509 12909 11512
rect 12943 11509 12955 11543
rect 13630 11540 13636 11552
rect 13591 11512 13636 11540
rect 12897 11503 12955 11509
rect 13630 11500 13636 11512
rect 13688 11500 13694 11552
rect 15010 11500 15016 11552
rect 15068 11540 15074 11552
rect 15105 11543 15163 11549
rect 15105 11540 15117 11543
rect 15068 11512 15117 11540
rect 15068 11500 15074 11512
rect 15105 11509 15117 11512
rect 15151 11509 15163 11543
rect 15105 11503 15163 11509
rect 15746 11500 15752 11552
rect 15804 11540 15810 11552
rect 15933 11543 15991 11549
rect 15933 11540 15945 11543
rect 15804 11512 15945 11540
rect 15804 11500 15810 11512
rect 15933 11509 15945 11512
rect 15979 11509 15991 11543
rect 15933 11503 15991 11509
rect 16298 11500 16304 11552
rect 16356 11540 16362 11552
rect 16669 11543 16727 11549
rect 16669 11540 16681 11543
rect 16356 11512 16681 11540
rect 16356 11500 16362 11512
rect 16669 11509 16681 11512
rect 16715 11509 16727 11543
rect 17218 11540 17224 11552
rect 17179 11512 17224 11540
rect 16669 11503 16727 11509
rect 17218 11500 17224 11512
rect 17276 11500 17282 11552
rect 18230 11540 18236 11552
rect 18191 11512 18236 11540
rect 18230 11500 18236 11512
rect 18288 11500 18294 11552
rect 19242 11540 19248 11552
rect 19203 11512 19248 11540
rect 19242 11500 19248 11512
rect 19300 11500 19306 11552
rect 19794 11500 19800 11552
rect 19852 11540 19858 11552
rect 20254 11540 20260 11552
rect 19852 11512 20260 11540
rect 19852 11500 19858 11512
rect 20254 11500 20260 11512
rect 20312 11540 20318 11552
rect 20533 11543 20591 11549
rect 20533 11540 20545 11543
rect 20312 11512 20545 11540
rect 20312 11500 20318 11512
rect 20533 11509 20545 11512
rect 20579 11509 20591 11543
rect 20533 11503 20591 11509
rect 21269 11543 21327 11549
rect 21269 11509 21281 11543
rect 21315 11540 21327 11543
rect 21726 11540 21732 11552
rect 21315 11512 21732 11540
rect 21315 11509 21327 11512
rect 21269 11503 21327 11509
rect 21726 11500 21732 11512
rect 21784 11500 21790 11552
rect 22094 11500 22100 11552
rect 22152 11540 22158 11552
rect 22649 11543 22707 11549
rect 22152 11512 22197 11540
rect 22152 11500 22158 11512
rect 22649 11509 22661 11543
rect 22695 11540 22707 11543
rect 23198 11540 23204 11552
rect 22695 11512 23204 11540
rect 22695 11509 22707 11512
rect 22649 11503 22707 11509
rect 23198 11500 23204 11512
rect 23256 11500 23262 11552
rect 24486 11540 24492 11552
rect 24447 11512 24492 11540
rect 24486 11500 24492 11512
rect 24544 11500 24550 11552
rect 24946 11500 24952 11552
rect 25004 11540 25010 11552
rect 25041 11543 25099 11549
rect 25041 11540 25053 11543
rect 25004 11512 25053 11540
rect 25004 11500 25010 11512
rect 25041 11509 25053 11512
rect 25087 11509 25099 11543
rect 25041 11503 25099 11509
rect 25406 11500 25412 11552
rect 25464 11540 25470 11552
rect 25593 11543 25651 11549
rect 25593 11540 25605 11543
rect 25464 11512 25605 11540
rect 25464 11500 25470 11512
rect 25593 11509 25605 11512
rect 25639 11509 25651 11543
rect 27356 11540 27384 11580
rect 27430 11568 27436 11620
rect 27488 11608 27494 11620
rect 36449 11611 36507 11617
rect 36449 11608 36461 11611
rect 27488 11580 36461 11608
rect 27488 11568 27494 11580
rect 36449 11577 36461 11580
rect 36495 11577 36507 11611
rect 36449 11571 36507 11577
rect 37921 11611 37979 11617
rect 37921 11577 37933 11611
rect 37967 11608 37979 11611
rect 41782 11608 41788 11620
rect 37967 11580 41788 11608
rect 37967 11577 37979 11580
rect 37921 11571 37979 11577
rect 41782 11568 41788 11580
rect 41840 11568 41846 11620
rect 27982 11540 27988 11552
rect 27356 11512 27988 11540
rect 25593 11503 25651 11509
rect 27982 11500 27988 11512
rect 28040 11500 28046 11552
rect 35710 11540 35716 11552
rect 35671 11512 35716 11540
rect 35710 11500 35716 11512
rect 35768 11500 35774 11552
rect 37369 11543 37427 11549
rect 37369 11509 37381 11543
rect 37415 11540 37427 11543
rect 37642 11540 37648 11552
rect 37415 11512 37648 11540
rect 37415 11509 37427 11512
rect 37369 11503 37427 11509
rect 37642 11500 37648 11512
rect 37700 11500 37706 11552
rect 38378 11540 38384 11552
rect 38339 11512 38384 11540
rect 38378 11500 38384 11512
rect 38436 11500 38442 11552
rect 42889 11543 42947 11549
rect 42889 11509 42901 11543
rect 42935 11540 42947 11543
rect 43070 11540 43076 11552
rect 42935 11512 43076 11540
rect 42935 11509 42947 11512
rect 42889 11503 42947 11509
rect 43070 11500 43076 11512
rect 43128 11500 43134 11552
rect 43441 11543 43499 11549
rect 43441 11509 43453 11543
rect 43487 11540 43499 11543
rect 43530 11540 43536 11552
rect 43487 11512 43536 11540
rect 43487 11509 43499 11512
rect 43441 11503 43499 11509
rect 43530 11500 43536 11512
rect 43588 11500 43594 11552
rect 1104 11450 58880 11472
rect 1104 11398 8174 11450
rect 8226 11398 8238 11450
rect 8290 11398 8302 11450
rect 8354 11398 8366 11450
rect 8418 11398 8430 11450
rect 8482 11398 22622 11450
rect 22674 11398 22686 11450
rect 22738 11398 22750 11450
rect 22802 11398 22814 11450
rect 22866 11398 22878 11450
rect 22930 11398 37070 11450
rect 37122 11398 37134 11450
rect 37186 11398 37198 11450
rect 37250 11398 37262 11450
rect 37314 11398 37326 11450
rect 37378 11398 51518 11450
rect 51570 11398 51582 11450
rect 51634 11398 51646 11450
rect 51698 11398 51710 11450
rect 51762 11398 51774 11450
rect 51826 11398 58880 11450
rect 1104 11376 58880 11398
rect 3878 11296 3884 11348
rect 3936 11336 3942 11348
rect 12710 11336 12716 11348
rect 3936 11308 12716 11336
rect 3936 11296 3942 11308
rect 12710 11296 12716 11308
rect 12768 11336 12774 11348
rect 13630 11336 13636 11348
rect 12768 11308 13636 11336
rect 12768 11296 12774 11308
rect 13630 11296 13636 11308
rect 13688 11336 13694 11348
rect 22462 11336 22468 11348
rect 13688 11308 22468 11336
rect 13688 11296 13694 11308
rect 22462 11296 22468 11308
rect 22520 11296 22526 11348
rect 25498 11336 25504 11348
rect 25459 11308 25504 11336
rect 25498 11296 25504 11308
rect 25556 11336 25562 11348
rect 26326 11336 26332 11348
rect 25556 11308 26332 11336
rect 25556 11296 25562 11308
rect 26326 11296 26332 11308
rect 26384 11296 26390 11348
rect 35713 11339 35771 11345
rect 35713 11305 35725 11339
rect 35759 11336 35771 11339
rect 38378 11336 38384 11348
rect 35759 11308 38384 11336
rect 35759 11305 35771 11308
rect 35713 11299 35771 11305
rect 38378 11296 38384 11308
rect 38436 11336 38442 11348
rect 39853 11339 39911 11345
rect 39853 11336 39865 11339
rect 38436 11308 39865 11336
rect 38436 11296 38442 11308
rect 39853 11305 39865 11308
rect 39899 11336 39911 11339
rect 41138 11336 41144 11348
rect 39899 11308 41144 11336
rect 39899 11305 39911 11308
rect 39853 11299 39911 11305
rect 41138 11296 41144 11308
rect 41196 11336 41202 11348
rect 43346 11336 43352 11348
rect 41196 11308 43352 11336
rect 41196 11296 41202 11308
rect 43346 11296 43352 11308
rect 43404 11296 43410 11348
rect 2038 11268 2044 11280
rect 1999 11240 2044 11268
rect 2038 11228 2044 11240
rect 2096 11228 2102 11280
rect 5902 11268 5908 11280
rect 5863 11240 5908 11268
rect 5902 11228 5908 11240
rect 5960 11268 5966 11280
rect 6362 11268 6368 11280
rect 5960 11240 6368 11268
rect 5960 11228 5966 11240
rect 6362 11228 6368 11240
rect 6420 11228 6426 11280
rect 6917 11271 6975 11277
rect 6917 11237 6929 11271
rect 6963 11237 6975 11271
rect 7742 11268 7748 11280
rect 7703 11240 7748 11268
rect 6917 11231 6975 11237
rect 3602 11160 3608 11212
rect 3660 11200 3666 11212
rect 6932 11200 6960 11231
rect 7742 11228 7748 11240
rect 7800 11228 7806 11280
rect 9030 11228 9036 11280
rect 9088 11268 9094 11280
rect 9401 11271 9459 11277
rect 9401 11268 9413 11271
rect 9088 11240 9413 11268
rect 9088 11228 9094 11240
rect 9401 11237 9413 11240
rect 9447 11237 9459 11271
rect 9401 11231 9459 11237
rect 10962 11228 10968 11280
rect 11020 11268 11026 11280
rect 11057 11271 11115 11277
rect 11057 11268 11069 11271
rect 11020 11240 11069 11268
rect 11020 11228 11026 11240
rect 11057 11237 11069 11240
rect 11103 11237 11115 11271
rect 15654 11268 15660 11280
rect 15615 11240 15660 11268
rect 11057 11231 11115 11237
rect 15654 11228 15660 11240
rect 15712 11228 15718 11280
rect 16022 11228 16028 11280
rect 16080 11268 16086 11280
rect 16117 11271 16175 11277
rect 16117 11268 16129 11271
rect 16080 11240 16129 11268
rect 16080 11228 16086 11240
rect 16117 11237 16129 11240
rect 16163 11237 16175 11271
rect 20162 11268 20168 11280
rect 20123 11240 20168 11268
rect 16117 11231 16175 11237
rect 20162 11228 20168 11240
rect 20220 11228 20226 11280
rect 21542 11268 21548 11280
rect 20916 11240 21548 11268
rect 10980 11200 11008 11228
rect 3660 11172 6960 11200
rect 7208 11172 11008 11200
rect 3660 11160 3666 11172
rect 3145 11135 3203 11141
rect 3145 11101 3157 11135
rect 3191 11132 3203 11135
rect 4430 11132 4436 11144
rect 3191 11104 4436 11132
rect 3191 11101 3203 11104
rect 3145 11095 3203 11101
rect 4430 11092 4436 11104
rect 4488 11092 4494 11144
rect 4801 11135 4859 11141
rect 4801 11101 4813 11135
rect 4847 11132 4859 11135
rect 4982 11132 4988 11144
rect 4847 11104 4988 11132
rect 4847 11101 4859 11104
rect 4801 11095 4859 11101
rect 4982 11092 4988 11104
rect 5040 11092 5046 11144
rect 6457 11135 6515 11141
rect 6457 11101 6469 11135
rect 6503 11132 6515 11135
rect 7098 11132 7104 11144
rect 6503 11104 7104 11132
rect 6503 11101 6515 11104
rect 6457 11095 6515 11101
rect 7098 11092 7104 11104
rect 7156 11092 7162 11144
rect 4154 11064 4160 11076
rect 4115 11036 4160 11064
rect 4154 11024 4160 11036
rect 4212 11024 4218 11076
rect 4890 11024 4896 11076
rect 4948 11064 4954 11076
rect 5810 11064 5816 11076
rect 4948 11036 5816 11064
rect 4948 11024 4954 11036
rect 5810 11024 5816 11036
rect 5868 11064 5874 11076
rect 7208 11064 7236 11172
rect 13630 11160 13636 11212
rect 13688 11200 13694 11212
rect 15013 11203 15071 11209
rect 15013 11200 15025 11203
rect 13688 11172 15025 11200
rect 13688 11160 13694 11172
rect 15013 11169 15025 11172
rect 15059 11169 15071 11203
rect 15013 11163 15071 11169
rect 15838 11160 15844 11212
rect 15896 11200 15902 11212
rect 17405 11203 17463 11209
rect 17405 11200 17417 11203
rect 15896 11172 17417 11200
rect 15896 11160 15902 11172
rect 17405 11169 17417 11172
rect 17451 11200 17463 11203
rect 20916 11200 20944 11240
rect 21542 11228 21548 11240
rect 21600 11228 21606 11280
rect 22094 11228 22100 11280
rect 22152 11268 22158 11280
rect 24762 11268 24768 11280
rect 22152 11240 24768 11268
rect 22152 11228 22158 11240
rect 24762 11228 24768 11240
rect 24820 11268 24826 11280
rect 24857 11271 24915 11277
rect 24857 11268 24869 11271
rect 24820 11240 24869 11268
rect 24820 11228 24826 11240
rect 24857 11237 24869 11240
rect 24903 11268 24915 11271
rect 38746 11268 38752 11280
rect 24903 11240 38752 11268
rect 24903 11237 24915 11240
rect 24857 11231 24915 11237
rect 38746 11228 38752 11240
rect 38804 11268 38810 11280
rect 39482 11268 39488 11280
rect 38804 11240 39488 11268
rect 38804 11228 38810 11240
rect 39482 11228 39488 11240
rect 39540 11228 39546 11280
rect 17451 11172 20944 11200
rect 17451 11169 17463 11172
rect 17405 11163 17463 11169
rect 20990 11160 20996 11212
rect 21048 11200 21054 11212
rect 36630 11200 36636 11212
rect 21048 11172 21093 11200
rect 26344 11172 36636 11200
rect 21048 11160 21054 11172
rect 7466 11092 7472 11144
rect 7524 11132 7530 11144
rect 7929 11135 7987 11141
rect 7929 11132 7941 11135
rect 7524 11104 7941 11132
rect 7524 11092 7530 11104
rect 7929 11101 7941 11104
rect 7975 11101 7987 11135
rect 7929 11095 7987 11101
rect 9585 11135 9643 11141
rect 9585 11101 9597 11135
rect 9631 11132 9643 11135
rect 12253 11135 12311 11141
rect 9631 11104 9996 11132
rect 9631 11101 9643 11104
rect 9585 11095 9643 11101
rect 9968 11076 9996 11104
rect 12253 11101 12265 11135
rect 12299 11132 12311 11135
rect 12342 11132 12348 11144
rect 12299 11104 12348 11132
rect 12299 11101 12311 11104
rect 12253 11095 12311 11101
rect 12342 11092 12348 11104
rect 12400 11092 12406 11144
rect 12897 11135 12955 11141
rect 12897 11101 12909 11135
rect 12943 11132 12955 11135
rect 13078 11132 13084 11144
rect 12943 11104 13084 11132
rect 12943 11101 12955 11104
rect 12897 11095 12955 11101
rect 13078 11092 13084 11104
rect 13136 11092 13142 11144
rect 13354 11132 13360 11144
rect 13315 11104 13360 11132
rect 13354 11092 13360 11104
rect 13412 11092 13418 11144
rect 13906 11092 13912 11144
rect 13964 11132 13970 11144
rect 14093 11135 14151 11141
rect 14093 11132 14105 11135
rect 13964 11104 14105 11132
rect 13964 11092 13970 11104
rect 14093 11101 14105 11104
rect 14139 11101 14151 11135
rect 14093 11095 14151 11101
rect 15473 11135 15531 11141
rect 15473 11101 15485 11135
rect 15519 11132 15531 11135
rect 15856 11132 15884 11160
rect 16298 11132 16304 11144
rect 15519 11104 15884 11132
rect 16259 11104 16304 11132
rect 15519 11101 15531 11104
rect 15473 11095 15531 11101
rect 5868 11036 7236 11064
rect 5868 11024 5874 11036
rect 8570 11024 8576 11076
rect 8628 11064 8634 11076
rect 9214 11064 9220 11076
rect 8628 11036 9220 11064
rect 8628 11024 8634 11036
rect 9214 11024 9220 11036
rect 9272 11064 9278 11076
rect 9272 11036 9904 11064
rect 9272 11024 9278 11036
rect 2590 10996 2596 11008
rect 2551 10968 2596 10996
rect 2590 10956 2596 10968
rect 2648 10956 2654 11008
rect 3786 10956 3792 11008
rect 3844 10996 3850 11008
rect 8478 10996 8484 11008
rect 3844 10968 8484 10996
rect 3844 10956 3850 10968
rect 8478 10956 8484 10968
rect 8536 10956 8542 11008
rect 9876 10996 9904 11036
rect 9950 11024 9956 11076
rect 10008 11064 10014 11076
rect 10045 11067 10103 11073
rect 10045 11064 10057 11067
rect 10008 11036 10057 11064
rect 10008 11024 10014 11036
rect 10045 11033 10057 11036
rect 10091 11033 10103 11067
rect 11517 11067 11575 11073
rect 11517 11064 11529 11067
rect 10045 11027 10103 11033
rect 10152 11036 11529 11064
rect 10152 10996 10180 11036
rect 11517 11033 11529 11036
rect 11563 11033 11575 11067
rect 11517 11027 11575 11033
rect 13262 11024 13268 11076
rect 13320 11064 13326 11076
rect 15488 11064 15516 11095
rect 16298 11092 16304 11104
rect 16356 11092 16362 11144
rect 16761 11135 16819 11141
rect 16761 11101 16773 11135
rect 16807 11132 16819 11135
rect 16850 11132 16856 11144
rect 16807 11104 16856 11132
rect 16807 11101 16819 11104
rect 16761 11095 16819 11101
rect 16850 11092 16856 11104
rect 16908 11092 16914 11144
rect 18598 11092 18604 11144
rect 18656 11132 18662 11144
rect 19242 11132 19248 11144
rect 18656 11104 19248 11132
rect 18656 11092 18662 11104
rect 19242 11092 19248 11104
rect 19300 11132 19306 11144
rect 22094 11132 22100 11144
rect 19300 11104 22100 11132
rect 19300 11092 19306 11104
rect 22094 11092 22100 11104
rect 22152 11092 22158 11144
rect 22186 11092 22192 11144
rect 22244 11132 22250 11144
rect 26344 11132 26372 11172
rect 36630 11160 36636 11172
rect 36688 11160 36694 11212
rect 27430 11132 27436 11144
rect 22244 11104 26372 11132
rect 27264 11104 27436 11132
rect 22244 11092 22250 11104
rect 13320 11036 15516 11064
rect 13320 11024 13326 11036
rect 15838 11024 15844 11076
rect 15896 11064 15902 11076
rect 17957 11067 18015 11073
rect 17957 11064 17969 11067
rect 15896 11036 17969 11064
rect 15896 11024 15902 11036
rect 17957 11033 17969 11036
rect 18003 11033 18015 11067
rect 17957 11027 18015 11033
rect 18693 11067 18751 11073
rect 18693 11033 18705 11067
rect 18739 11064 18751 11067
rect 18782 11064 18788 11076
rect 18739 11036 18788 11064
rect 18739 11033 18751 11036
rect 18693 11027 18751 11033
rect 18782 11024 18788 11036
rect 18840 11024 18846 11076
rect 19337 11067 19395 11073
rect 19337 11033 19349 11067
rect 19383 11064 19395 11067
rect 19518 11064 19524 11076
rect 19383 11036 19524 11064
rect 19383 11033 19395 11036
rect 19337 11027 19395 11033
rect 19518 11024 19524 11036
rect 19576 11024 19582 11076
rect 21450 11064 21456 11076
rect 21411 11036 21456 11064
rect 21450 11024 21456 11036
rect 21508 11024 21514 11076
rect 21542 11024 21548 11076
rect 21600 11064 21606 11076
rect 21600 11036 22416 11064
rect 21600 11024 21606 11036
rect 9876 10968 10180 10996
rect 22388 10996 22416 11036
rect 22462 11024 22468 11076
rect 22520 11064 22526 11076
rect 22649 11067 22707 11073
rect 22649 11064 22661 11067
rect 22520 11036 22661 11064
rect 22520 11024 22526 11036
rect 22649 11033 22661 11036
rect 22695 11033 22707 11067
rect 24118 11064 24124 11076
rect 22649 11027 22707 11033
rect 22756 11036 24124 11064
rect 22756 10996 22784 11036
rect 24118 11024 24124 11036
rect 24176 11024 24182 11076
rect 25866 11024 25872 11076
rect 25924 11064 25930 11076
rect 25961 11067 26019 11073
rect 25961 11064 25973 11067
rect 25924 11036 25973 11064
rect 25924 11024 25930 11036
rect 25961 11033 25973 11036
rect 26007 11033 26019 11067
rect 26602 11064 26608 11076
rect 26563 11036 26608 11064
rect 25961 11027 26019 11033
rect 26602 11024 26608 11036
rect 26660 11024 26666 11076
rect 26694 11024 26700 11076
rect 26752 11064 26758 11076
rect 27264 11073 27292 11104
rect 27430 11092 27436 11104
rect 27488 11132 27494 11144
rect 27801 11135 27859 11141
rect 27801 11132 27813 11135
rect 27488 11104 27813 11132
rect 27488 11092 27494 11104
rect 27801 11101 27813 11104
rect 27847 11101 27859 11135
rect 27801 11095 27859 11101
rect 27982 11092 27988 11144
rect 28040 11132 28046 11144
rect 38654 11132 38660 11144
rect 28040 11104 38660 11132
rect 28040 11092 28046 11104
rect 38654 11092 38660 11104
rect 38712 11092 38718 11144
rect 27249 11067 27307 11073
rect 27249 11064 27261 11067
rect 26752 11036 27261 11064
rect 26752 11024 26758 11036
rect 27249 11033 27261 11036
rect 27295 11033 27307 11067
rect 27249 11027 27307 11033
rect 27522 11024 27528 11076
rect 27580 11064 27586 11076
rect 28629 11067 28687 11073
rect 28629 11064 28641 11067
rect 27580 11036 28641 11064
rect 27580 11024 27586 11036
rect 28629 11033 28641 11036
rect 28675 11033 28687 11067
rect 28629 11027 28687 11033
rect 29362 11024 29368 11076
rect 29420 11064 29426 11076
rect 29549 11067 29607 11073
rect 29549 11064 29561 11067
rect 29420 11036 29561 11064
rect 29420 11024 29426 11036
rect 29549 11033 29561 11036
rect 29595 11033 29607 11067
rect 35158 11064 35164 11076
rect 35119 11036 35164 11064
rect 29549 11027 29607 11033
rect 35158 11024 35164 11036
rect 35216 11024 35222 11076
rect 36170 11064 36176 11076
rect 36131 11036 36176 11064
rect 36170 11024 36176 11036
rect 36228 11024 36234 11076
rect 36630 11024 36636 11076
rect 36688 11064 36694 11076
rect 36725 11067 36783 11073
rect 36725 11064 36737 11067
rect 36688 11036 36737 11064
rect 36688 11024 36694 11036
rect 36725 11033 36737 11036
rect 36771 11033 36783 11067
rect 36725 11027 36783 11033
rect 37461 11067 37519 11073
rect 37461 11033 37473 11067
rect 37507 11033 37519 11067
rect 39117 11067 39175 11073
rect 39117 11064 39129 11067
rect 37461 11027 37519 11033
rect 38212 11036 39129 11064
rect 22388 10968 22784 10996
rect 23293 10999 23351 11005
rect 23293 10965 23305 10999
rect 23339 10996 23351 10999
rect 23382 10996 23388 11008
rect 23339 10968 23388 10996
rect 23339 10965 23351 10968
rect 23293 10959 23351 10965
rect 23382 10956 23388 10968
rect 23440 10956 23446 11008
rect 23658 10956 23664 11008
rect 23716 10996 23722 11008
rect 23753 10999 23811 11005
rect 23753 10996 23765 10999
rect 23716 10968 23765 10996
rect 23716 10956 23722 10968
rect 23753 10965 23765 10968
rect 23799 10965 23811 10999
rect 23753 10959 23811 10965
rect 36906 10956 36912 11008
rect 36964 10996 36970 11008
rect 37476 10996 37504 11027
rect 38212 11008 38240 11036
rect 39117 11033 39129 11036
rect 39163 11033 39175 11067
rect 40402 11064 40408 11076
rect 40363 11036 40408 11064
rect 39117 11027 39175 11033
rect 40402 11024 40408 11036
rect 40460 11024 40466 11076
rect 41966 11064 41972 11076
rect 41927 11036 41972 11064
rect 41966 11024 41972 11036
rect 42024 11024 42030 11076
rect 42705 11067 42763 11073
rect 42705 11033 42717 11067
rect 42751 11064 42763 11067
rect 42886 11064 42892 11076
rect 42751 11036 42892 11064
rect 42751 11033 42763 11036
rect 42705 11027 42763 11033
rect 42886 11024 42892 11036
rect 42944 11024 42950 11076
rect 43806 11024 43812 11076
rect 43864 11064 43870 11076
rect 43901 11067 43959 11073
rect 43901 11064 43913 11067
rect 43864 11036 43913 11064
rect 43864 11024 43870 11036
rect 43901 11033 43913 11036
rect 43947 11033 43959 11067
rect 43901 11027 43959 11033
rect 36964 10968 37504 10996
rect 38105 10999 38163 11005
rect 36964 10956 36970 10968
rect 38105 10965 38117 10999
rect 38151 10996 38163 10999
rect 38194 10996 38200 11008
rect 38151 10968 38200 10996
rect 38151 10965 38163 10968
rect 38105 10959 38163 10965
rect 38194 10956 38200 10968
rect 38252 10956 38258 11008
rect 38562 10996 38568 11008
rect 38523 10968 38568 10996
rect 38562 10956 38568 10968
rect 38620 10956 38626 11008
rect 45002 10996 45008 11008
rect 44963 10968 45008 10996
rect 45002 10956 45008 10968
rect 45060 10956 45066 11008
rect 1104 10906 58880 10928
rect 1104 10854 15398 10906
rect 15450 10854 15462 10906
rect 15514 10854 15526 10906
rect 15578 10854 15590 10906
rect 15642 10854 15654 10906
rect 15706 10854 29846 10906
rect 29898 10854 29910 10906
rect 29962 10854 29974 10906
rect 30026 10854 30038 10906
rect 30090 10854 30102 10906
rect 30154 10854 44294 10906
rect 44346 10854 44358 10906
rect 44410 10854 44422 10906
rect 44474 10854 44486 10906
rect 44538 10854 44550 10906
rect 44602 10854 58880 10906
rect 1104 10832 58880 10854
rect 1762 10792 1768 10804
rect 1723 10764 1768 10792
rect 1762 10752 1768 10764
rect 1820 10752 1826 10804
rect 2590 10752 2596 10804
rect 2648 10792 2654 10804
rect 3786 10792 3792 10804
rect 2648 10764 3792 10792
rect 2648 10752 2654 10764
rect 3786 10752 3792 10764
rect 3844 10752 3850 10804
rect 3970 10792 3976 10804
rect 3931 10764 3976 10792
rect 3970 10752 3976 10764
rect 4028 10752 4034 10804
rect 5810 10792 5816 10804
rect 5771 10764 5816 10792
rect 5810 10752 5816 10764
rect 5868 10752 5874 10804
rect 8205 10795 8263 10801
rect 8205 10761 8217 10795
rect 8251 10761 8263 10795
rect 8205 10755 8263 10761
rect 1578 10656 1584 10668
rect 1539 10628 1584 10656
rect 1578 10616 1584 10628
rect 1636 10616 1642 10668
rect 2225 10659 2283 10665
rect 2225 10625 2237 10659
rect 2271 10656 2283 10659
rect 2608 10656 2636 10752
rect 2682 10684 2688 10736
rect 2740 10724 2746 10736
rect 8220 10724 8248 10755
rect 23290 10752 23296 10804
rect 23348 10792 23354 10804
rect 25777 10795 25835 10801
rect 25777 10792 25789 10795
rect 23348 10764 25789 10792
rect 23348 10752 23354 10764
rect 25777 10761 25789 10764
rect 25823 10792 25835 10795
rect 26234 10792 26240 10804
rect 25823 10764 26240 10792
rect 25823 10761 25835 10764
rect 25777 10755 25835 10761
rect 26234 10752 26240 10764
rect 26292 10752 26298 10804
rect 36538 10792 36544 10804
rect 36499 10764 36544 10792
rect 36538 10752 36544 10764
rect 36596 10752 36602 10804
rect 37458 10752 37464 10804
rect 37516 10792 37522 10804
rect 37921 10795 37979 10801
rect 37921 10792 37933 10795
rect 37516 10764 37933 10792
rect 37516 10752 37522 10764
rect 37921 10761 37933 10764
rect 37967 10792 37979 10795
rect 38562 10792 38568 10804
rect 37967 10764 38568 10792
rect 37967 10761 37979 10764
rect 37921 10755 37979 10761
rect 38562 10752 38568 10764
rect 38620 10752 38626 10804
rect 39482 10792 39488 10804
rect 39443 10764 39488 10792
rect 39482 10752 39488 10764
rect 39540 10752 39546 10804
rect 41138 10792 41144 10804
rect 41099 10764 41144 10792
rect 41138 10752 41144 10764
rect 41196 10752 41202 10804
rect 41782 10792 41788 10804
rect 41743 10764 41788 10792
rect 41782 10752 41788 10764
rect 41840 10752 41846 10804
rect 43346 10752 43352 10804
rect 43404 10792 43410 10804
rect 44082 10792 44088 10804
rect 43404 10764 44088 10792
rect 43404 10752 43410 10764
rect 44082 10752 44088 10764
rect 44140 10792 44146 10804
rect 44453 10795 44511 10801
rect 44453 10792 44465 10795
rect 44140 10764 44465 10792
rect 44140 10752 44146 10764
rect 44453 10761 44465 10764
rect 44499 10792 44511 10795
rect 48317 10795 48375 10801
rect 48317 10792 48329 10795
rect 44499 10764 48329 10792
rect 44499 10761 44511 10764
rect 44453 10755 44511 10761
rect 48317 10761 48329 10764
rect 48363 10792 48375 10795
rect 48777 10795 48835 10801
rect 48777 10792 48789 10795
rect 48363 10764 48789 10792
rect 48363 10761 48375 10764
rect 48317 10755 48375 10761
rect 48777 10761 48789 10764
rect 48823 10761 48835 10795
rect 48777 10755 48835 10761
rect 2740 10696 8248 10724
rect 2740 10684 2746 10696
rect 10042 10684 10048 10736
rect 10100 10724 10106 10736
rect 14182 10724 14188 10736
rect 10100 10696 14188 10724
rect 10100 10684 10106 10696
rect 14182 10684 14188 10696
rect 14240 10684 14246 10736
rect 23308 10724 23336 10752
rect 19904 10696 23336 10724
rect 2271 10628 2636 10656
rect 3789 10659 3847 10665
rect 2271 10625 2283 10628
rect 2225 10619 2283 10625
rect 3789 10625 3801 10659
rect 3835 10656 3847 10659
rect 4154 10656 4160 10668
rect 3835 10628 4160 10656
rect 3835 10625 3847 10628
rect 3789 10619 3847 10625
rect 4154 10616 4160 10628
rect 4212 10616 4218 10668
rect 4706 10656 4712 10668
rect 4667 10628 4712 10656
rect 4706 10616 4712 10628
rect 4764 10616 4770 10668
rect 7101 10659 7159 10665
rect 7101 10625 7113 10659
rect 7147 10656 7159 10659
rect 7374 10656 7380 10668
rect 7147 10628 7380 10656
rect 7147 10625 7159 10628
rect 7101 10619 7159 10625
rect 7374 10616 7380 10628
rect 7432 10616 7438 10668
rect 7745 10659 7803 10665
rect 7745 10656 7757 10659
rect 7484 10628 7757 10656
rect 2038 10548 2044 10600
rect 2096 10588 2102 10600
rect 6457 10591 6515 10597
rect 2096 10560 2774 10588
rect 2096 10548 2102 10560
rect 2746 10520 2774 10560
rect 6457 10557 6469 10591
rect 6503 10588 6515 10591
rect 7006 10588 7012 10600
rect 6503 10560 7012 10588
rect 6503 10557 6515 10560
rect 6457 10551 6515 10557
rect 7006 10548 7012 10560
rect 7064 10588 7070 10600
rect 7484 10588 7512 10628
rect 7745 10625 7757 10628
rect 7791 10625 7803 10659
rect 7745 10619 7803 10625
rect 8389 10659 8447 10665
rect 8389 10625 8401 10659
rect 8435 10625 8447 10659
rect 8389 10619 8447 10625
rect 8941 10659 8999 10665
rect 8941 10625 8953 10659
rect 8987 10656 8999 10659
rect 9306 10656 9312 10668
rect 8987 10628 9312 10656
rect 8987 10625 8999 10628
rect 8941 10619 8999 10625
rect 7064 10560 7512 10588
rect 7064 10548 7070 10560
rect 7650 10548 7656 10600
rect 7708 10588 7714 10600
rect 8404 10588 8432 10619
rect 9306 10616 9312 10628
rect 9364 10656 9370 10668
rect 9401 10659 9459 10665
rect 9401 10656 9413 10659
rect 9364 10628 9413 10656
rect 9364 10616 9370 10628
rect 9401 10625 9413 10628
rect 9447 10625 9459 10659
rect 9401 10619 9459 10625
rect 10134 10616 10140 10668
rect 10192 10656 10198 10668
rect 10413 10659 10471 10665
rect 10413 10656 10425 10659
rect 10192 10628 10425 10656
rect 10192 10616 10198 10628
rect 10413 10625 10425 10628
rect 10459 10656 10471 10659
rect 10873 10659 10931 10665
rect 10873 10656 10885 10659
rect 10459 10628 10885 10656
rect 10459 10625 10471 10628
rect 10413 10619 10471 10625
rect 10873 10625 10885 10628
rect 10919 10625 10931 10659
rect 11790 10656 11796 10668
rect 11751 10628 11796 10656
rect 10873 10619 10931 10625
rect 11790 10616 11796 10628
rect 11848 10616 11854 10668
rect 15838 10616 15844 10668
rect 15896 10656 15902 10668
rect 16117 10659 16175 10665
rect 16117 10656 16129 10659
rect 15896 10628 16129 10656
rect 15896 10616 15902 10628
rect 16117 10625 16129 10628
rect 16163 10625 16175 10659
rect 16117 10619 16175 10625
rect 16206 10616 16212 10668
rect 16264 10656 16270 10668
rect 16669 10659 16727 10665
rect 16669 10656 16681 10659
rect 16264 10628 16681 10656
rect 16264 10616 16270 10628
rect 16669 10625 16681 10628
rect 16715 10625 16727 10659
rect 17678 10656 17684 10668
rect 17639 10628 17684 10656
rect 16669 10619 16727 10625
rect 17678 10616 17684 10628
rect 17736 10616 17742 10668
rect 19904 10665 19932 10696
rect 28902 10684 28908 10736
rect 28960 10724 28966 10736
rect 34606 10724 34612 10736
rect 28960 10696 34612 10724
rect 28960 10684 28966 10696
rect 34606 10684 34612 10696
rect 34664 10724 34670 10736
rect 35250 10724 35256 10736
rect 34664 10696 35256 10724
rect 34664 10684 34670 10696
rect 35250 10684 35256 10696
rect 35308 10684 35314 10736
rect 36556 10724 36584 10752
rect 46934 10724 46940 10736
rect 36556 10696 46940 10724
rect 46934 10684 46940 10696
rect 46992 10684 46998 10736
rect 19889 10659 19947 10665
rect 19889 10625 19901 10659
rect 19935 10625 19947 10659
rect 19889 10619 19947 10625
rect 20073 10659 20131 10665
rect 20073 10625 20085 10659
rect 20119 10656 20131 10659
rect 20717 10659 20775 10665
rect 20717 10656 20729 10659
rect 20119 10628 20729 10656
rect 20119 10625 20131 10628
rect 20073 10619 20131 10625
rect 20717 10625 20729 10628
rect 20763 10625 20775 10659
rect 20717 10619 20775 10625
rect 22370 10616 22376 10668
rect 22428 10656 22434 10668
rect 22649 10659 22707 10665
rect 22649 10656 22661 10659
rect 22428 10628 22661 10656
rect 22428 10616 22434 10628
rect 22649 10625 22661 10628
rect 22695 10625 22707 10659
rect 23474 10656 23480 10668
rect 23435 10628 23480 10656
rect 22649 10619 22707 10625
rect 23474 10616 23480 10628
rect 23532 10616 23538 10668
rect 25222 10616 25228 10668
rect 25280 10656 25286 10668
rect 25593 10659 25651 10665
rect 25593 10656 25605 10659
rect 25280 10628 25605 10656
rect 25280 10616 25286 10628
rect 25593 10625 25605 10628
rect 25639 10625 25651 10659
rect 27154 10656 27160 10668
rect 27115 10628 27160 10656
rect 25593 10619 25651 10625
rect 27154 10616 27160 10628
rect 27212 10616 27218 10668
rect 28810 10616 28816 10668
rect 28868 10656 28874 10668
rect 29365 10659 29423 10665
rect 29365 10656 29377 10659
rect 28868 10628 29377 10656
rect 28868 10616 28874 10628
rect 29365 10625 29377 10628
rect 29411 10625 29423 10659
rect 29365 10619 29423 10625
rect 38654 10616 38660 10668
rect 38712 10656 38718 10668
rect 38712 10628 46704 10656
rect 38712 10616 38718 10628
rect 7708 10560 8432 10588
rect 7708 10548 7714 10560
rect 11422 10548 11428 10600
rect 11480 10588 11486 10600
rect 11517 10591 11575 10597
rect 11517 10588 11529 10591
rect 11480 10560 11529 10588
rect 11480 10548 11486 10560
rect 11517 10557 11529 10560
rect 11563 10557 11575 10591
rect 11517 10551 11575 10557
rect 17310 10548 17316 10600
rect 17368 10588 17374 10600
rect 17405 10591 17463 10597
rect 17405 10588 17417 10591
rect 17368 10560 17417 10588
rect 17368 10548 17374 10560
rect 17405 10557 17417 10560
rect 17451 10557 17463 10591
rect 17405 10551 17463 10557
rect 19705 10591 19763 10597
rect 19705 10557 19717 10591
rect 19751 10588 19763 10591
rect 20162 10588 20168 10600
rect 19751 10560 20168 10588
rect 19751 10557 19763 10560
rect 19705 10551 19763 10557
rect 20162 10548 20168 10560
rect 20220 10548 20226 10600
rect 23382 10548 23388 10600
rect 23440 10588 23446 10600
rect 26050 10588 26056 10600
rect 23440 10560 26056 10588
rect 23440 10548 23446 10560
rect 26050 10548 26056 10560
rect 26108 10588 26114 10600
rect 26237 10591 26295 10597
rect 26237 10588 26249 10591
rect 26108 10560 26249 10588
rect 26108 10548 26114 10560
rect 26237 10557 26249 10560
rect 26283 10588 26295 10591
rect 31202 10588 31208 10600
rect 26283 10560 31208 10588
rect 26283 10557 26295 10560
rect 26237 10551 26295 10557
rect 31202 10548 31208 10560
rect 31260 10548 31266 10600
rect 33965 10591 34023 10597
rect 33965 10557 33977 10591
rect 34011 10588 34023 10591
rect 34514 10588 34520 10600
rect 34011 10560 34520 10588
rect 34011 10557 34023 10560
rect 33965 10551 34023 10557
rect 34514 10548 34520 10560
rect 34572 10548 34578 10600
rect 36906 10548 36912 10600
rect 36964 10588 36970 10600
rect 38933 10591 38991 10597
rect 38933 10588 38945 10591
rect 36964 10560 38945 10588
rect 36964 10548 36970 10560
rect 38933 10557 38945 10560
rect 38979 10557 38991 10591
rect 43990 10588 43996 10600
rect 38933 10551 38991 10557
rect 39040 10560 43996 10588
rect 7561 10523 7619 10529
rect 7561 10520 7573 10523
rect 2746 10492 7573 10520
rect 7561 10489 7573 10492
rect 7607 10489 7619 10523
rect 7561 10483 7619 10489
rect 8938 10480 8944 10532
rect 8996 10520 9002 10532
rect 10229 10523 10287 10529
rect 10229 10520 10241 10523
rect 8996 10492 10241 10520
rect 8996 10480 9002 10492
rect 10229 10489 10241 10492
rect 10275 10489 10287 10523
rect 10229 10483 10287 10489
rect 13541 10523 13599 10529
rect 13541 10489 13553 10523
rect 13587 10520 13599 10523
rect 14274 10520 14280 10532
rect 13587 10492 14280 10520
rect 13587 10489 13599 10492
rect 13541 10483 13599 10489
rect 14274 10480 14280 10492
rect 14332 10480 14338 10532
rect 15473 10523 15531 10529
rect 15473 10489 15485 10523
rect 15519 10520 15531 10523
rect 16114 10520 16120 10532
rect 15519 10492 16120 10520
rect 15519 10489 15531 10492
rect 15473 10483 15531 10489
rect 16114 10480 16120 10492
rect 16172 10480 16178 10532
rect 19245 10523 19303 10529
rect 19245 10489 19257 10523
rect 19291 10520 19303 10523
rect 20254 10520 20260 10532
rect 19291 10492 20260 10520
rect 19291 10489 19303 10492
rect 19245 10483 19303 10489
rect 20254 10480 20260 10492
rect 20312 10520 20318 10532
rect 21177 10523 21235 10529
rect 21177 10520 21189 10523
rect 20312 10492 21189 10520
rect 20312 10480 20318 10492
rect 21177 10489 21189 10492
rect 21223 10489 21235 10523
rect 21177 10483 21235 10489
rect 23661 10523 23719 10529
rect 23661 10489 23673 10523
rect 23707 10520 23719 10523
rect 24670 10520 24676 10532
rect 23707 10492 24676 10520
rect 23707 10489 23719 10492
rect 23661 10483 23719 10489
rect 24670 10480 24676 10492
rect 24728 10480 24734 10532
rect 29086 10480 29092 10532
rect 29144 10520 29150 10532
rect 30561 10523 30619 10529
rect 30561 10520 30573 10523
rect 29144 10492 30573 10520
rect 29144 10480 29150 10492
rect 30561 10489 30573 10492
rect 30607 10489 30619 10523
rect 30561 10483 30619 10489
rect 38194 10480 38200 10532
rect 38252 10520 38258 10532
rect 38381 10523 38439 10529
rect 38381 10520 38393 10523
rect 38252 10492 38393 10520
rect 38252 10480 38258 10492
rect 38381 10489 38393 10492
rect 38427 10489 38439 10523
rect 38381 10483 38439 10489
rect 2409 10455 2467 10461
rect 2409 10421 2421 10455
rect 2455 10452 2467 10455
rect 2682 10452 2688 10464
rect 2455 10424 2688 10452
rect 2455 10421 2467 10424
rect 2409 10415 2467 10421
rect 2682 10412 2688 10424
rect 2740 10412 2746 10464
rect 3329 10455 3387 10461
rect 3329 10421 3341 10455
rect 3375 10452 3387 10455
rect 3786 10452 3792 10464
rect 3375 10424 3792 10452
rect 3375 10421 3387 10424
rect 3329 10415 3387 10421
rect 3786 10412 3792 10424
rect 3844 10412 3850 10464
rect 4890 10452 4896 10464
rect 4851 10424 4896 10452
rect 4890 10412 4896 10424
rect 4948 10412 4954 10464
rect 6914 10452 6920 10464
rect 6875 10424 6920 10452
rect 6914 10412 6920 10424
rect 6972 10412 6978 10464
rect 9582 10452 9588 10464
rect 9543 10424 9588 10452
rect 9582 10412 9588 10424
rect 9640 10412 9646 10464
rect 12250 10412 12256 10464
rect 12308 10452 12314 10464
rect 12529 10455 12587 10461
rect 12529 10452 12541 10455
rect 12308 10424 12541 10452
rect 12308 10412 12314 10424
rect 12529 10421 12541 10424
rect 12575 10452 12587 10455
rect 13446 10452 13452 10464
rect 12575 10424 13452 10452
rect 12575 10421 12587 10424
rect 12529 10415 12587 10421
rect 13446 10412 13452 10424
rect 13504 10412 13510 10464
rect 14185 10455 14243 10461
rect 14185 10421 14197 10455
rect 14231 10452 14243 10455
rect 14734 10452 14740 10464
rect 14231 10424 14740 10452
rect 14231 10421 14243 10424
rect 14185 10415 14243 10421
rect 14734 10412 14740 10424
rect 14792 10412 14798 10464
rect 14829 10455 14887 10461
rect 14829 10421 14841 10455
rect 14875 10452 14887 10455
rect 15286 10452 15292 10464
rect 14875 10424 15292 10452
rect 14875 10421 14887 10424
rect 14829 10415 14887 10421
rect 15286 10412 15292 10424
rect 15344 10412 15350 10464
rect 15930 10452 15936 10464
rect 15891 10424 15936 10452
rect 15930 10412 15936 10424
rect 15988 10412 15994 10464
rect 16853 10455 16911 10461
rect 16853 10421 16865 10455
rect 16899 10452 16911 10455
rect 17402 10452 17408 10464
rect 16899 10424 17408 10452
rect 16899 10421 16911 10424
rect 16853 10415 16911 10421
rect 17402 10412 17408 10424
rect 17460 10412 17466 10464
rect 18414 10452 18420 10464
rect 18375 10424 18420 10452
rect 18414 10412 18420 10424
rect 18472 10412 18478 10464
rect 20438 10412 20444 10464
rect 20496 10452 20502 10464
rect 20533 10455 20591 10461
rect 20533 10452 20545 10455
rect 20496 10424 20545 10452
rect 20496 10412 20502 10424
rect 20533 10421 20545 10424
rect 20579 10421 20591 10455
rect 20533 10415 20591 10421
rect 22094 10412 22100 10464
rect 22152 10452 22158 10464
rect 22833 10455 22891 10461
rect 22152 10424 22197 10452
rect 22152 10412 22158 10424
rect 22833 10421 22845 10455
rect 22879 10452 22891 10455
rect 23014 10452 23020 10464
rect 22879 10424 23020 10452
rect 22879 10421 22891 10424
rect 22833 10415 22891 10421
rect 23014 10412 23020 10424
rect 23072 10412 23078 10464
rect 24210 10412 24216 10464
rect 24268 10452 24274 10464
rect 24581 10455 24639 10461
rect 24581 10452 24593 10455
rect 24268 10424 24593 10452
rect 24268 10412 24274 10424
rect 24581 10421 24593 10424
rect 24627 10421 24639 10455
rect 24581 10415 24639 10421
rect 26418 10412 26424 10464
rect 26476 10452 26482 10464
rect 26973 10455 27031 10461
rect 26973 10452 26985 10455
rect 26476 10424 26985 10452
rect 26476 10412 26482 10424
rect 26973 10421 26985 10424
rect 27019 10421 27031 10455
rect 26973 10415 27031 10421
rect 27614 10412 27620 10464
rect 27672 10452 27678 10464
rect 27985 10455 28043 10461
rect 27985 10452 27997 10455
rect 27672 10424 27997 10452
rect 27672 10412 27678 10424
rect 27985 10421 27997 10424
rect 28031 10452 28043 10455
rect 28721 10455 28779 10461
rect 28721 10452 28733 10455
rect 28031 10424 28733 10452
rect 28031 10421 28043 10424
rect 27985 10415 28043 10421
rect 28721 10421 28733 10424
rect 28767 10421 28779 10455
rect 29546 10452 29552 10464
rect 29507 10424 29552 10452
rect 28721 10415 28779 10421
rect 29546 10412 29552 10424
rect 29604 10412 29610 10464
rect 30101 10455 30159 10461
rect 30101 10421 30113 10455
rect 30147 10452 30159 10455
rect 30190 10452 30196 10464
rect 30147 10424 30196 10452
rect 30147 10421 30159 10424
rect 30101 10415 30159 10421
rect 30190 10412 30196 10424
rect 30248 10412 30254 10464
rect 33134 10412 33140 10464
rect 33192 10452 33198 10464
rect 33321 10455 33379 10461
rect 33321 10452 33333 10455
rect 33192 10424 33333 10452
rect 33192 10412 33198 10424
rect 33321 10421 33333 10424
rect 33367 10421 33379 10455
rect 33321 10415 33379 10421
rect 34609 10455 34667 10461
rect 34609 10421 34621 10455
rect 34655 10452 34667 10455
rect 34790 10452 34796 10464
rect 34655 10424 34796 10452
rect 34655 10421 34667 10424
rect 34609 10415 34667 10421
rect 34790 10412 34796 10424
rect 34848 10412 34854 10464
rect 35529 10455 35587 10461
rect 35529 10421 35541 10455
rect 35575 10452 35587 10455
rect 36078 10452 36084 10464
rect 35575 10424 36084 10452
rect 35575 10421 35587 10424
rect 35529 10415 35587 10421
rect 36078 10412 36084 10424
rect 36136 10412 36142 10464
rect 37369 10455 37427 10461
rect 37369 10421 37381 10455
rect 37415 10452 37427 10455
rect 37550 10452 37556 10464
rect 37415 10424 37556 10452
rect 37415 10421 37427 10424
rect 37369 10415 37427 10421
rect 37550 10412 37556 10424
rect 37608 10452 37614 10464
rect 39040 10452 39068 10560
rect 43990 10548 43996 10560
rect 44048 10548 44054 10600
rect 46676 10588 46704 10628
rect 46750 10616 46756 10668
rect 46808 10656 46814 10668
rect 47581 10659 47639 10665
rect 47581 10656 47593 10659
rect 46808 10628 47593 10656
rect 46808 10616 46814 10628
rect 47581 10625 47593 10628
rect 47627 10625 47639 10659
rect 47581 10619 47639 10625
rect 50522 10588 50528 10600
rect 46676 10560 50528 10588
rect 50522 10548 50528 10560
rect 50580 10548 50586 10600
rect 41230 10480 41236 10532
rect 41288 10520 41294 10532
rect 45002 10520 45008 10532
rect 41288 10492 45008 10520
rect 41288 10480 41294 10492
rect 45002 10480 45008 10492
rect 45060 10520 45066 10532
rect 45281 10523 45339 10529
rect 45281 10520 45293 10523
rect 45060 10492 45293 10520
rect 45060 10480 45066 10492
rect 45281 10489 45293 10492
rect 45327 10489 45339 10523
rect 45281 10483 45339 10489
rect 37608 10424 39068 10452
rect 37608 10412 37614 10424
rect 39850 10412 39856 10464
rect 39908 10452 39914 10464
rect 40037 10455 40095 10461
rect 40037 10452 40049 10455
rect 39908 10424 40049 10452
rect 39908 10412 39914 10424
rect 40037 10421 40049 10424
rect 40083 10421 40095 10455
rect 40037 10415 40095 10421
rect 40494 10412 40500 10464
rect 40552 10452 40558 10464
rect 40589 10455 40647 10461
rect 40589 10452 40601 10455
rect 40552 10424 40601 10452
rect 40552 10412 40558 10424
rect 40589 10421 40601 10424
rect 40635 10421 40647 10455
rect 42518 10452 42524 10464
rect 42479 10424 42524 10452
rect 40589 10415 40647 10421
rect 42518 10412 42524 10424
rect 42576 10412 42582 10464
rect 42886 10412 42892 10464
rect 42944 10452 42950 10464
rect 42981 10455 43039 10461
rect 42981 10452 42993 10455
rect 42944 10424 42993 10452
rect 42944 10412 42950 10424
rect 42981 10421 42993 10424
rect 43027 10421 43039 10455
rect 43990 10452 43996 10464
rect 43951 10424 43996 10452
rect 42981 10415 43039 10421
rect 43990 10412 43996 10424
rect 44048 10412 44054 10464
rect 45462 10412 45468 10464
rect 45520 10452 45526 10464
rect 45833 10455 45891 10461
rect 45833 10452 45845 10455
rect 45520 10424 45845 10452
rect 45520 10412 45526 10424
rect 45833 10421 45845 10424
rect 45879 10421 45891 10455
rect 46382 10452 46388 10464
rect 46343 10424 46388 10452
rect 45833 10415 45891 10421
rect 46382 10412 46388 10424
rect 46440 10412 46446 10464
rect 47765 10455 47823 10461
rect 47765 10421 47777 10455
rect 47811 10452 47823 10455
rect 48958 10452 48964 10464
rect 47811 10424 48964 10452
rect 47811 10421 47823 10424
rect 47765 10415 47823 10421
rect 48958 10412 48964 10424
rect 49016 10412 49022 10464
rect 1104 10362 58880 10384
rect 1104 10310 8174 10362
rect 8226 10310 8238 10362
rect 8290 10310 8302 10362
rect 8354 10310 8366 10362
rect 8418 10310 8430 10362
rect 8482 10310 22622 10362
rect 22674 10310 22686 10362
rect 22738 10310 22750 10362
rect 22802 10310 22814 10362
rect 22866 10310 22878 10362
rect 22930 10310 37070 10362
rect 37122 10310 37134 10362
rect 37186 10310 37198 10362
rect 37250 10310 37262 10362
rect 37314 10310 37326 10362
rect 37378 10310 51518 10362
rect 51570 10310 51582 10362
rect 51634 10310 51646 10362
rect 51698 10310 51710 10362
rect 51762 10310 51774 10362
rect 51826 10310 58880 10362
rect 1104 10288 58880 10310
rect 4062 10248 4068 10260
rect 3804 10220 4068 10248
rect 3145 10183 3203 10189
rect 3145 10149 3157 10183
rect 3191 10149 3203 10183
rect 3145 10143 3203 10149
rect 1670 10044 1676 10056
rect 1631 10016 1676 10044
rect 1670 10004 1676 10016
rect 1728 10004 1734 10056
rect 2317 10047 2375 10053
rect 2317 10013 2329 10047
rect 2363 10044 2375 10047
rect 2958 10044 2964 10056
rect 2363 10016 2774 10044
rect 2919 10016 2964 10044
rect 2363 10013 2375 10016
rect 2317 10007 2375 10013
rect 2746 9976 2774 10016
rect 2958 10004 2964 10016
rect 3016 10004 3022 10056
rect 3160 10044 3188 10143
rect 3804 10121 3832 10220
rect 4062 10208 4068 10220
rect 4120 10248 4126 10260
rect 6914 10248 6920 10260
rect 4120 10220 6920 10248
rect 4120 10208 4126 10220
rect 5813 10183 5871 10189
rect 5813 10149 5825 10183
rect 5859 10149 5871 10183
rect 5813 10143 5871 10149
rect 3789 10115 3847 10121
rect 3789 10081 3801 10115
rect 3835 10081 3847 10115
rect 3789 10075 3847 10081
rect 4065 10047 4123 10053
rect 4065 10044 4077 10047
rect 3160 10016 4077 10044
rect 4065 10013 4077 10016
rect 4111 10013 4123 10047
rect 5626 10044 5632 10056
rect 5587 10016 5632 10044
rect 4065 10007 4123 10013
rect 5626 10004 5632 10016
rect 5684 10004 5690 10056
rect 5828 10044 5856 10143
rect 6288 10121 6316 10220
rect 6914 10208 6920 10220
rect 6972 10208 6978 10260
rect 10229 10251 10287 10257
rect 10229 10217 10241 10251
rect 10275 10248 10287 10251
rect 11790 10248 11796 10260
rect 10275 10220 11796 10248
rect 10275 10217 10287 10220
rect 10229 10211 10287 10217
rect 11790 10208 11796 10220
rect 11848 10208 11854 10260
rect 16669 10251 16727 10257
rect 11992 10220 15516 10248
rect 6273 10115 6331 10121
rect 6273 10081 6285 10115
rect 6319 10081 6331 10115
rect 6273 10075 6331 10081
rect 11422 10072 11428 10124
rect 11480 10112 11486 10124
rect 11992 10121 12020 10220
rect 14936 10121 14964 10220
rect 15488 10180 15516 10220
rect 16669 10217 16681 10251
rect 16715 10248 16727 10251
rect 17678 10248 17684 10260
rect 16715 10220 17684 10248
rect 16715 10217 16727 10220
rect 16669 10211 16727 10217
rect 17678 10208 17684 10220
rect 17736 10208 17742 10260
rect 17770 10208 17776 10260
rect 17828 10248 17834 10260
rect 46382 10248 46388 10260
rect 17828 10220 46388 10248
rect 17828 10208 17834 10220
rect 46382 10208 46388 10220
rect 46440 10248 46446 10260
rect 47210 10248 47216 10260
rect 46440 10220 47216 10248
rect 46440 10208 46446 10220
rect 47210 10208 47216 10220
rect 47268 10208 47274 10260
rect 17129 10183 17187 10189
rect 17129 10180 17141 10183
rect 15488 10152 17141 10180
rect 17129 10149 17141 10152
rect 17175 10149 17187 10183
rect 35250 10180 35256 10192
rect 35211 10152 35256 10180
rect 17129 10143 17187 10149
rect 35250 10140 35256 10152
rect 35308 10140 35314 10192
rect 38654 10140 38660 10192
rect 38712 10180 38718 10192
rect 38841 10183 38899 10189
rect 38841 10180 38853 10183
rect 38712 10152 38853 10180
rect 38712 10140 38718 10152
rect 38841 10149 38853 10152
rect 38887 10149 38899 10183
rect 42061 10183 42119 10189
rect 42061 10180 42073 10183
rect 38841 10143 38899 10149
rect 40236 10152 42073 10180
rect 11977 10115 12035 10121
rect 11977 10112 11989 10115
rect 11480 10084 11989 10112
rect 11480 10072 11486 10084
rect 11977 10081 11989 10084
rect 12023 10081 12035 10115
rect 11977 10075 12035 10081
rect 14921 10115 14979 10121
rect 14921 10081 14933 10115
rect 14967 10081 14979 10115
rect 14921 10075 14979 10081
rect 20717 10115 20775 10121
rect 20717 10081 20729 10115
rect 20763 10112 20775 10115
rect 20898 10112 20904 10124
rect 20763 10084 20904 10112
rect 20763 10081 20775 10084
rect 20717 10075 20775 10081
rect 20898 10072 20904 10084
rect 20956 10112 20962 10124
rect 22554 10112 22560 10124
rect 20956 10084 22560 10112
rect 20956 10072 20962 10084
rect 22554 10072 22560 10084
rect 22612 10072 22618 10124
rect 32306 10072 32312 10124
rect 32364 10112 32370 10124
rect 32364 10084 33088 10112
rect 32364 10072 32370 10084
rect 6549 10047 6607 10053
rect 6549 10044 6561 10047
rect 5828 10016 6561 10044
rect 6549 10013 6561 10016
rect 6595 10013 6607 10047
rect 6549 10007 6607 10013
rect 8389 10047 8447 10053
rect 8389 10013 8401 10047
rect 8435 10013 8447 10047
rect 8389 10007 8447 10013
rect 4430 9976 4436 9988
rect 2746 9948 4436 9976
rect 4430 9936 4436 9948
rect 4488 9936 4494 9988
rect 8404 9976 8432 10007
rect 9122 10004 9128 10056
rect 9180 10044 9186 10056
rect 9585 10047 9643 10053
rect 9585 10044 9597 10047
rect 9180 10016 9597 10044
rect 9180 10004 9186 10016
rect 9585 10013 9597 10016
rect 9631 10013 9643 10047
rect 10042 10044 10048 10056
rect 10003 10016 10048 10044
rect 9585 10007 9643 10013
rect 10042 10004 10048 10016
rect 10100 10004 10106 10056
rect 10689 10047 10747 10053
rect 10689 10013 10701 10047
rect 10735 10044 10747 10047
rect 11238 10044 11244 10056
rect 10735 10016 11244 10044
rect 10735 10013 10747 10016
rect 10689 10007 10747 10013
rect 11238 10004 11244 10016
rect 11296 10004 11302 10056
rect 11330 10004 11336 10056
rect 11388 10044 11394 10056
rect 12253 10047 12311 10053
rect 11388 10016 11433 10044
rect 11388 10004 11394 10016
rect 12253 10013 12265 10047
rect 12299 10013 12311 10047
rect 14090 10044 14096 10056
rect 14051 10016 14096 10044
rect 12253 10007 12311 10013
rect 10778 9976 10784 9988
rect 8404 9948 10784 9976
rect 10778 9936 10784 9948
rect 10836 9936 10842 9988
rect 12268 9976 12296 10007
rect 14090 10004 14096 10016
rect 14148 10004 14154 10056
rect 15197 10047 15255 10053
rect 15197 10044 15209 10047
rect 14292 10016 15209 10044
rect 10888 9948 12296 9976
rect 1854 9908 1860 9920
rect 1815 9880 1860 9908
rect 1854 9868 1860 9880
rect 1912 9868 1918 9920
rect 2498 9908 2504 9920
rect 2459 9880 2504 9908
rect 2498 9868 2504 9880
rect 2556 9868 2562 9920
rect 4798 9908 4804 9920
rect 4711 9880 4804 9908
rect 4798 9868 4804 9880
rect 4856 9908 4862 9920
rect 7285 9911 7343 9917
rect 7285 9908 7297 9911
rect 4856 9880 7297 9908
rect 4856 9868 4862 9880
rect 7285 9877 7297 9880
rect 7331 9908 7343 9911
rect 7558 9908 7564 9920
rect 7331 9880 7564 9908
rect 7331 9877 7343 9880
rect 7285 9871 7343 9877
rect 7558 9868 7564 9880
rect 7616 9868 7622 9920
rect 7834 9868 7840 9920
rect 7892 9908 7898 9920
rect 8205 9911 8263 9917
rect 8205 9908 8217 9911
rect 7892 9880 8217 9908
rect 7892 9868 7898 9880
rect 8205 9877 8217 9880
rect 8251 9877 8263 9911
rect 8205 9871 8263 9877
rect 9493 9911 9551 9917
rect 9493 9877 9505 9911
rect 9539 9908 9551 9911
rect 10226 9908 10232 9920
rect 9539 9880 10232 9908
rect 9539 9877 9551 9880
rect 9493 9871 9551 9877
rect 10226 9868 10232 9880
rect 10284 9868 10290 9920
rect 10888 9917 10916 9948
rect 10873 9911 10931 9917
rect 10873 9877 10885 9911
rect 10919 9877 10931 9911
rect 10873 9871 10931 9877
rect 11517 9911 11575 9917
rect 11517 9877 11529 9911
rect 11563 9908 11575 9911
rect 12618 9908 12624 9920
rect 11563 9880 12624 9908
rect 11563 9877 11575 9880
rect 11517 9871 11575 9877
rect 12618 9868 12624 9880
rect 12676 9868 12682 9920
rect 12989 9911 13047 9917
rect 12989 9877 13001 9911
rect 13035 9908 13047 9911
rect 13446 9908 13452 9920
rect 13035 9880 13452 9908
rect 13035 9877 13047 9880
rect 12989 9871 13047 9877
rect 13446 9868 13452 9880
rect 13504 9868 13510 9920
rect 13541 9911 13599 9917
rect 13541 9877 13553 9911
rect 13587 9908 13599 9911
rect 14182 9908 14188 9920
rect 13587 9880 14188 9908
rect 13587 9877 13599 9880
rect 13541 9871 13599 9877
rect 14182 9868 14188 9880
rect 14240 9868 14246 9920
rect 14292 9917 14320 10016
rect 15197 10013 15209 10016
rect 15243 10013 15255 10047
rect 16485 10047 16543 10053
rect 16485 10044 16497 10047
rect 15197 10007 15255 10013
rect 15396 10016 16497 10044
rect 14277 9911 14335 9917
rect 14277 9877 14289 9911
rect 14323 9877 14335 9911
rect 14277 9871 14335 9877
rect 14918 9868 14924 9920
rect 14976 9908 14982 9920
rect 15396 9908 15424 10016
rect 16485 10013 16497 10016
rect 16531 10013 16543 10047
rect 17310 10044 17316 10056
rect 17223 10016 17316 10044
rect 16485 10007 16543 10013
rect 17310 10004 17316 10016
rect 17368 10004 17374 10056
rect 18049 10047 18107 10053
rect 18049 10013 18061 10047
rect 18095 10044 18107 10047
rect 18138 10044 18144 10056
rect 18095 10016 18144 10044
rect 18095 10013 18107 10016
rect 18049 10007 18107 10013
rect 18138 10004 18144 10016
rect 18196 10004 18202 10056
rect 18506 10044 18512 10056
rect 18467 10016 18512 10044
rect 18506 10004 18512 10016
rect 18564 10004 18570 10056
rect 20438 10044 20444 10056
rect 20399 10016 20444 10044
rect 20438 10004 20444 10016
rect 20496 10004 20502 10056
rect 21361 10047 21419 10053
rect 21361 10013 21373 10047
rect 21407 10013 21419 10047
rect 21361 10007 21419 10013
rect 22097 10047 22155 10053
rect 22097 10013 22109 10047
rect 22143 10044 22155 10047
rect 22278 10044 22284 10056
rect 22143 10016 22284 10044
rect 22143 10013 22155 10016
rect 22097 10007 22155 10013
rect 17328 9976 17356 10004
rect 21376 9976 21404 10007
rect 22278 10004 22284 10016
rect 22336 10004 22342 10056
rect 22833 10047 22891 10053
rect 22833 10013 22845 10047
rect 22879 10044 22891 10047
rect 23014 10044 23020 10056
rect 22879 10016 23020 10044
rect 22879 10013 22891 10016
rect 22833 10007 22891 10013
rect 23014 10004 23020 10016
rect 23072 10004 23078 10056
rect 24394 10044 24400 10056
rect 24355 10016 24400 10044
rect 24394 10004 24400 10016
rect 24452 10004 24458 10056
rect 24670 10044 24676 10056
rect 24631 10016 24676 10044
rect 24670 10004 24676 10016
rect 24728 10004 24734 10056
rect 25682 10004 25688 10056
rect 25740 10044 25746 10056
rect 26145 10047 26203 10053
rect 26145 10044 26157 10047
rect 25740 10016 26157 10044
rect 25740 10004 25746 10016
rect 26145 10013 26157 10016
rect 26191 10013 26203 10047
rect 26418 10044 26424 10056
rect 26379 10016 26424 10044
rect 26145 10007 26203 10013
rect 26418 10004 26424 10016
rect 26476 10004 26482 10056
rect 30834 10044 30840 10056
rect 30795 10016 30840 10044
rect 30834 10004 30840 10016
rect 30892 10004 30898 10056
rect 31113 10047 31171 10053
rect 31113 10013 31125 10047
rect 31159 10013 31171 10047
rect 31113 10007 31171 10013
rect 24854 9976 24860 9988
rect 17328 9948 21220 9976
rect 21376 9948 24860 9976
rect 14976 9880 15424 9908
rect 14976 9868 14982 9880
rect 15470 9868 15476 9920
rect 15528 9908 15534 9920
rect 15933 9911 15991 9917
rect 15933 9908 15945 9911
rect 15528 9880 15945 9908
rect 15528 9868 15534 9880
rect 15933 9877 15945 9880
rect 15979 9908 15991 9911
rect 18414 9908 18420 9920
rect 15979 9880 18420 9908
rect 15979 9877 15991 9880
rect 15933 9871 15991 9877
rect 18414 9868 18420 9880
rect 18472 9868 18478 9920
rect 19702 9908 19708 9920
rect 19663 9880 19708 9908
rect 19702 9868 19708 9880
rect 19760 9868 19766 9920
rect 21192 9917 21220 9948
rect 24854 9936 24860 9948
rect 24912 9936 24918 9988
rect 27982 9976 27988 9988
rect 27172 9948 27988 9976
rect 21177 9911 21235 9917
rect 21177 9877 21189 9911
rect 21223 9877 21235 9911
rect 21910 9908 21916 9920
rect 21871 9880 21916 9908
rect 21177 9871 21235 9877
rect 21910 9868 21916 9880
rect 21968 9868 21974 9920
rect 22002 9868 22008 9920
rect 22060 9908 22066 9920
rect 27172 9917 27200 9948
rect 27982 9936 27988 9948
rect 28040 9936 28046 9988
rect 28074 9936 28080 9988
rect 28132 9976 28138 9988
rect 28813 9979 28871 9985
rect 28813 9976 28825 9979
rect 28132 9948 28825 9976
rect 28132 9936 28138 9948
rect 28813 9945 28825 9948
rect 28859 9976 28871 9979
rect 28902 9976 28908 9988
rect 28859 9948 28908 9976
rect 28859 9945 28871 9948
rect 28813 9939 28871 9945
rect 28902 9936 28908 9948
rect 28960 9936 28966 9988
rect 30558 9936 30564 9988
rect 30616 9976 30622 9988
rect 31128 9976 31156 10007
rect 31202 10004 31208 10056
rect 31260 10044 31266 10056
rect 31260 10016 32996 10044
rect 31260 10004 31266 10016
rect 30616 9948 31156 9976
rect 30616 9936 30622 9948
rect 23569 9911 23627 9917
rect 23569 9908 23581 9911
rect 22060 9880 23581 9908
rect 22060 9868 22066 9880
rect 23569 9877 23581 9880
rect 23615 9908 23627 9911
rect 25409 9911 25467 9917
rect 25409 9908 25421 9911
rect 23615 9880 25421 9908
rect 23615 9877 23627 9880
rect 23569 9871 23627 9877
rect 25409 9877 25421 9880
rect 25455 9908 25467 9911
rect 27157 9911 27215 9917
rect 27157 9908 27169 9911
rect 25455 9880 27169 9908
rect 25455 9877 25467 9880
rect 25409 9871 25467 9877
rect 27157 9877 27169 9880
rect 27203 9877 27215 9911
rect 27157 9871 27215 9877
rect 27338 9868 27344 9920
rect 27396 9908 27402 9920
rect 27617 9911 27675 9917
rect 27617 9908 27629 9911
rect 27396 9880 27629 9908
rect 27396 9868 27402 9880
rect 27617 9877 27629 9880
rect 27663 9877 27675 9911
rect 27617 9871 27675 9877
rect 28353 9911 28411 9917
rect 28353 9877 28365 9911
rect 28399 9908 28411 9911
rect 28442 9908 28448 9920
rect 28399 9880 28448 9908
rect 28399 9877 28411 9880
rect 28353 9871 28411 9877
rect 28442 9868 28448 9880
rect 28500 9868 28506 9920
rect 29454 9868 29460 9920
rect 29512 9908 29518 9920
rect 29549 9911 29607 9917
rect 29549 9908 29561 9911
rect 29512 9880 29561 9908
rect 29512 9868 29518 9880
rect 29549 9877 29561 9880
rect 29595 9877 29607 9911
rect 29549 9871 29607 9877
rect 30101 9911 30159 9917
rect 30101 9877 30113 9911
rect 30147 9908 30159 9911
rect 30282 9908 30288 9920
rect 30147 9880 30288 9908
rect 30147 9877 30159 9880
rect 30101 9871 30159 9877
rect 30282 9868 30288 9880
rect 30340 9908 30346 9920
rect 32490 9908 32496 9920
rect 30340 9880 32496 9908
rect 30340 9868 30346 9880
rect 32490 9868 32496 9880
rect 32548 9868 32554 9920
rect 32582 9868 32588 9920
rect 32640 9908 32646 9920
rect 32968 9908 32996 10016
rect 33060 9976 33088 10084
rect 40236 10056 40264 10152
rect 42061 10149 42073 10152
rect 42107 10180 42119 10183
rect 42107 10152 42748 10180
rect 42107 10149 42119 10152
rect 42061 10143 42119 10149
rect 42720 10121 42748 10152
rect 42705 10115 42763 10121
rect 42705 10081 42717 10115
rect 42751 10081 42763 10115
rect 42705 10075 42763 10081
rect 48958 10072 48964 10124
rect 49016 10112 49022 10124
rect 52270 10112 52276 10124
rect 49016 10084 52276 10112
rect 49016 10072 49022 10084
rect 52270 10072 52276 10084
rect 52328 10072 52334 10124
rect 33137 10047 33195 10053
rect 33137 10013 33149 10047
rect 33183 10044 33195 10047
rect 33318 10044 33324 10056
rect 33183 10016 33324 10044
rect 33183 10013 33195 10016
rect 33137 10007 33195 10013
rect 33318 10004 33324 10016
rect 33376 10004 33382 10056
rect 33413 10047 33471 10053
rect 33413 10013 33425 10047
rect 33459 10013 33471 10047
rect 33413 10007 33471 10013
rect 36265 10047 36323 10053
rect 36265 10013 36277 10047
rect 36311 10044 36323 10047
rect 36538 10044 36544 10056
rect 36311 10016 36544 10044
rect 36311 10013 36323 10016
rect 36265 10007 36323 10013
rect 33428 9976 33456 10007
rect 36538 10004 36544 10016
rect 36596 10004 36602 10056
rect 38102 10044 38108 10056
rect 36648 10016 37872 10044
rect 38063 10016 38108 10044
rect 36648 9976 36676 10016
rect 33060 9948 33456 9976
rect 33980 9948 36676 9976
rect 33980 9908 34008 9948
rect 34146 9908 34152 9920
rect 32640 9880 32685 9908
rect 32968 9880 34008 9908
rect 34107 9880 34152 9908
rect 32640 9868 32646 9880
rect 34146 9868 34152 9880
rect 34204 9868 34210 9920
rect 34793 9911 34851 9917
rect 34793 9877 34805 9911
rect 34839 9908 34851 9911
rect 36170 9908 36176 9920
rect 34839 9880 36176 9908
rect 34839 9877 34851 9880
rect 34793 9871 34851 9877
rect 36170 9868 36176 9880
rect 36228 9868 36234 9920
rect 36354 9908 36360 9920
rect 36315 9880 36360 9908
rect 36354 9868 36360 9880
rect 36412 9908 36418 9920
rect 36906 9908 36912 9920
rect 36412 9880 36912 9908
rect 36412 9868 36418 9880
rect 36906 9868 36912 9880
rect 36964 9868 36970 9920
rect 37366 9908 37372 9920
rect 37327 9880 37372 9908
rect 37366 9868 37372 9880
rect 37424 9868 37430 9920
rect 37844 9908 37872 10016
rect 38102 10004 38108 10016
rect 38160 10004 38166 10056
rect 38381 10047 38439 10053
rect 38381 10013 38393 10047
rect 38427 10044 38439 10047
rect 40218 10044 40224 10056
rect 38427 10016 40224 10044
rect 38427 10013 38439 10016
rect 38381 10007 38439 10013
rect 38010 9936 38016 9988
rect 38068 9976 38074 9988
rect 38396 9976 38424 10007
rect 40218 10004 40224 10016
rect 40276 10004 40282 10056
rect 42245 10047 42303 10053
rect 42245 10013 42257 10047
rect 42291 10044 42303 10047
rect 42426 10044 42432 10056
rect 42291 10016 42432 10044
rect 42291 10013 42303 10016
rect 42245 10007 42303 10013
rect 42426 10004 42432 10016
rect 42484 10004 42490 10056
rect 42978 10044 42984 10056
rect 42939 10016 42984 10044
rect 42978 10004 42984 10016
rect 43036 10004 43042 10056
rect 45646 10044 45652 10056
rect 45607 10016 45652 10044
rect 45646 10004 45652 10016
rect 45704 10004 45710 10056
rect 46474 10044 46480 10056
rect 46435 10016 46480 10044
rect 46474 10004 46480 10016
rect 46532 10004 46538 10056
rect 46750 10044 46756 10056
rect 46711 10016 46756 10044
rect 46750 10004 46756 10016
rect 46808 10044 46814 10056
rect 47397 10047 47455 10053
rect 47397 10044 47409 10047
rect 46808 10016 47409 10044
rect 46808 10004 46814 10016
rect 47397 10013 47409 10016
rect 47443 10013 47455 10047
rect 47670 10044 47676 10056
rect 47631 10016 47676 10044
rect 47397 10007 47455 10013
rect 47670 10004 47676 10016
rect 47728 10004 47734 10056
rect 48501 10047 48559 10053
rect 48501 10013 48513 10047
rect 48547 10013 48559 10047
rect 49234 10044 49240 10056
rect 49195 10016 49240 10044
rect 48501 10007 48559 10013
rect 41049 9979 41107 9985
rect 41049 9976 41061 9979
rect 38068 9948 38424 9976
rect 38856 9948 41061 9976
rect 38068 9936 38074 9948
rect 38856 9908 38884 9948
rect 41049 9945 41061 9948
rect 41095 9976 41107 9979
rect 41230 9976 41236 9988
rect 41095 9948 41236 9976
rect 41095 9945 41107 9948
rect 41049 9939 41107 9945
rect 41230 9936 41236 9948
rect 41288 9936 41294 9988
rect 45664 9976 45692 10004
rect 48516 9976 48544 10007
rect 49234 10004 49240 10016
rect 49292 10004 49298 10056
rect 52546 10044 52552 10056
rect 52507 10016 52552 10044
rect 52546 10004 52552 10016
rect 52604 10004 52610 10056
rect 53374 10044 53380 10056
rect 53335 10016 53380 10044
rect 53374 10004 53380 10016
rect 53432 10004 53438 10056
rect 50062 9976 50068 9988
rect 45664 9948 50068 9976
rect 50062 9936 50068 9948
rect 50120 9936 50126 9988
rect 37844 9880 38884 9908
rect 39758 9868 39764 9920
rect 39816 9908 39822 9920
rect 39853 9911 39911 9917
rect 39853 9908 39865 9911
rect 39816 9880 39865 9908
rect 39816 9868 39822 9880
rect 39853 9877 39865 9880
rect 39899 9908 39911 9911
rect 40405 9911 40463 9917
rect 40405 9908 40417 9911
rect 39899 9880 40417 9908
rect 39899 9877 39911 9880
rect 39853 9871 39911 9877
rect 40405 9877 40417 9880
rect 40451 9877 40463 9911
rect 43714 9908 43720 9920
rect 43675 9880 43720 9908
rect 40405 9871 40463 9877
rect 43714 9868 43720 9880
rect 43772 9868 43778 9920
rect 44174 9908 44180 9920
rect 44135 9880 44180 9908
rect 44174 9868 44180 9880
rect 44232 9868 44238 9920
rect 44634 9868 44640 9920
rect 44692 9908 44698 9920
rect 45005 9911 45063 9917
rect 45005 9908 45017 9911
rect 44692 9880 45017 9908
rect 44692 9868 44698 9880
rect 45005 9877 45017 9880
rect 45051 9877 45063 9911
rect 45005 9871 45063 9877
rect 48866 9868 48872 9920
rect 48924 9908 48930 9920
rect 49053 9911 49111 9917
rect 49053 9908 49065 9911
rect 48924 9880 49065 9908
rect 48924 9868 48930 9880
rect 49053 9877 49065 9880
rect 49099 9877 49111 9911
rect 49053 9871 49111 9877
rect 1104 9818 58880 9840
rect 1104 9766 15398 9818
rect 15450 9766 15462 9818
rect 15514 9766 15526 9818
rect 15578 9766 15590 9818
rect 15642 9766 15654 9818
rect 15706 9766 29846 9818
rect 29898 9766 29910 9818
rect 29962 9766 29974 9818
rect 30026 9766 30038 9818
rect 30090 9766 30102 9818
rect 30154 9766 44294 9818
rect 44346 9766 44358 9818
rect 44410 9766 44422 9818
rect 44474 9766 44486 9818
rect 44538 9766 44550 9818
rect 44602 9766 58880 9818
rect 1104 9744 58880 9766
rect 2777 9707 2835 9713
rect 2777 9673 2789 9707
rect 2823 9704 2835 9707
rect 2958 9704 2964 9716
rect 2823 9676 2964 9704
rect 2823 9673 2835 9676
rect 2777 9667 2835 9673
rect 2958 9664 2964 9676
rect 3016 9664 3022 9716
rect 4249 9707 4307 9713
rect 4249 9673 4261 9707
rect 4295 9704 4307 9707
rect 4798 9704 4804 9716
rect 4295 9676 4804 9704
rect 4295 9673 4307 9676
rect 4249 9667 4307 9673
rect 4798 9664 4804 9676
rect 4856 9664 4862 9716
rect 5626 9664 5632 9716
rect 5684 9704 5690 9716
rect 6365 9707 6423 9713
rect 6365 9704 6377 9707
rect 5684 9676 6377 9704
rect 5684 9664 5690 9676
rect 6365 9673 6377 9676
rect 6411 9673 6423 9707
rect 6365 9667 6423 9673
rect 10042 9664 10048 9716
rect 10100 9704 10106 9716
rect 10505 9707 10563 9713
rect 10505 9704 10517 9707
rect 10100 9676 10517 9704
rect 10100 9664 10106 9676
rect 10505 9673 10517 9676
rect 10551 9673 10563 9707
rect 12250 9704 12256 9716
rect 10505 9667 10563 9673
rect 11164 9676 12256 9704
rect 3142 9636 3148 9648
rect 2516 9608 3148 9636
rect 1762 9568 1768 9580
rect 1723 9540 1768 9568
rect 1762 9528 1768 9540
rect 1820 9528 1826 9580
rect 2516 9577 2544 9608
rect 3142 9596 3148 9608
rect 3200 9596 3206 9648
rect 4062 9636 4068 9648
rect 3252 9608 4068 9636
rect 2501 9571 2559 9577
rect 2501 9537 2513 9571
rect 2547 9537 2559 9571
rect 2501 9531 2559 9537
rect 2593 9571 2651 9577
rect 2593 9537 2605 9571
rect 2639 9568 2651 9571
rect 3050 9568 3056 9580
rect 2639 9540 3056 9568
rect 2639 9537 2651 9540
rect 2593 9531 2651 9537
rect 2516 9500 2544 9531
rect 3050 9528 3056 9540
rect 3108 9528 3114 9580
rect 3252 9577 3280 9608
rect 4062 9596 4068 9608
rect 4120 9596 4126 9648
rect 7282 9596 7288 9648
rect 7340 9636 7346 9648
rect 11164 9636 11192 9676
rect 12250 9664 12256 9676
rect 12308 9664 12314 9716
rect 13446 9664 13452 9716
rect 13504 9704 13510 9716
rect 17770 9704 17776 9716
rect 13504 9676 17776 9704
rect 13504 9664 13510 9676
rect 17770 9664 17776 9676
rect 17828 9664 17834 9716
rect 18141 9707 18199 9713
rect 18141 9673 18153 9707
rect 18187 9704 18199 9707
rect 18414 9704 18420 9716
rect 18187 9676 18420 9704
rect 18187 9673 18199 9676
rect 18141 9667 18199 9673
rect 18414 9664 18420 9676
rect 18472 9664 18478 9716
rect 19334 9664 19340 9716
rect 19392 9704 19398 9716
rect 19702 9704 19708 9716
rect 19392 9676 19708 9704
rect 19392 9664 19398 9676
rect 19702 9664 19708 9676
rect 19760 9704 19766 9716
rect 19889 9707 19947 9713
rect 19889 9704 19901 9707
rect 19760 9676 19901 9704
rect 19760 9664 19766 9676
rect 19889 9673 19901 9676
rect 19935 9704 19947 9707
rect 22002 9704 22008 9716
rect 19935 9676 22008 9704
rect 19935 9673 19947 9676
rect 19889 9667 19947 9673
rect 22002 9664 22008 9676
rect 22060 9664 22066 9716
rect 22370 9704 22376 9716
rect 22331 9676 22376 9704
rect 22370 9664 22376 9676
rect 22428 9664 22434 9716
rect 22554 9664 22560 9716
rect 22612 9704 22618 9716
rect 24213 9707 24271 9713
rect 24213 9704 24225 9707
rect 22612 9676 24225 9704
rect 22612 9664 22618 9676
rect 24213 9673 24225 9676
rect 24259 9704 24271 9707
rect 24394 9704 24400 9716
rect 24259 9676 24400 9704
rect 24259 9673 24271 9676
rect 24213 9667 24271 9673
rect 24394 9664 24400 9676
rect 24452 9664 24458 9716
rect 24854 9704 24860 9716
rect 24815 9676 24860 9704
rect 24854 9664 24860 9676
rect 24912 9664 24918 9716
rect 26421 9707 26479 9713
rect 26421 9673 26433 9707
rect 26467 9704 26479 9707
rect 27154 9704 27160 9716
rect 26467 9676 27160 9704
rect 26467 9673 26479 9676
rect 26421 9667 26479 9673
rect 27154 9664 27160 9676
rect 27212 9664 27218 9716
rect 27982 9704 27988 9716
rect 27943 9676 27988 9704
rect 27982 9664 27988 9676
rect 28040 9664 28046 9716
rect 30834 9664 30840 9716
rect 30892 9704 30898 9716
rect 30929 9707 30987 9713
rect 30929 9704 30941 9707
rect 30892 9676 30941 9704
rect 30892 9664 30898 9676
rect 30929 9673 30941 9676
rect 30975 9673 30987 9707
rect 32306 9704 32312 9716
rect 32267 9676 32312 9704
rect 30929 9667 30987 9673
rect 32306 9664 32312 9676
rect 32364 9664 32370 9716
rect 32490 9664 32496 9716
rect 32548 9704 32554 9716
rect 33781 9707 33839 9713
rect 33781 9704 33793 9707
rect 32548 9676 33793 9704
rect 32548 9664 32554 9676
rect 33781 9673 33793 9676
rect 33827 9704 33839 9707
rect 34146 9704 34152 9716
rect 33827 9676 34152 9704
rect 33827 9673 33839 9676
rect 33781 9667 33839 9673
rect 34146 9664 34152 9676
rect 34204 9704 34210 9716
rect 34241 9707 34299 9713
rect 34241 9704 34253 9707
rect 34204 9676 34253 9704
rect 34204 9664 34210 9676
rect 34241 9673 34253 9676
rect 34287 9673 34299 9707
rect 37366 9704 37372 9716
rect 34241 9667 34299 9673
rect 36280 9676 37372 9704
rect 7340 9608 11192 9636
rect 7340 9596 7346 9608
rect 11238 9596 11244 9648
rect 11296 9636 11302 9648
rect 11517 9639 11575 9645
rect 11517 9636 11529 9639
rect 11296 9608 11529 9636
rect 11296 9596 11302 9608
rect 11517 9605 11529 9608
rect 11563 9605 11575 9639
rect 11517 9599 11575 9605
rect 13081 9639 13139 9645
rect 13081 9605 13093 9639
rect 13127 9636 13139 9639
rect 14090 9636 14096 9648
rect 13127 9608 14096 9636
rect 13127 9605 13139 9608
rect 13081 9599 13139 9605
rect 14090 9596 14096 9608
rect 14148 9596 14154 9648
rect 14918 9636 14924 9648
rect 14879 9608 14924 9636
rect 14918 9596 14924 9608
rect 14976 9596 14982 9648
rect 15749 9639 15807 9645
rect 15749 9605 15761 9639
rect 15795 9636 15807 9639
rect 16206 9636 16212 9648
rect 15795 9608 16212 9636
rect 15795 9605 15807 9608
rect 15749 9599 15807 9605
rect 16206 9596 16212 9608
rect 16264 9596 16270 9648
rect 17310 9636 17316 9648
rect 17144 9608 17316 9636
rect 3237 9571 3295 9577
rect 3237 9537 3249 9571
rect 3283 9537 3295 9571
rect 3510 9568 3516 9580
rect 3471 9540 3516 9568
rect 3237 9531 3295 9537
rect 3510 9528 3516 9540
rect 3568 9528 3574 9580
rect 3878 9528 3884 9580
rect 3936 9568 3942 9580
rect 4985 9571 5043 9577
rect 4985 9568 4997 9571
rect 3936 9540 4997 9568
rect 3936 9528 3942 9540
rect 4985 9537 4997 9540
rect 5031 9537 5043 9571
rect 4985 9531 5043 9537
rect 5074 9528 5080 9580
rect 5132 9568 5138 9580
rect 5169 9571 5227 9577
rect 5169 9568 5181 9571
rect 5132 9540 5181 9568
rect 5132 9528 5138 9540
rect 5169 9537 5181 9540
rect 5215 9537 5227 9571
rect 5169 9531 5227 9537
rect 5629 9571 5687 9577
rect 5629 9537 5641 9571
rect 5675 9568 5687 9571
rect 6454 9568 6460 9580
rect 5675 9540 6460 9568
rect 5675 9537 5687 9540
rect 5629 9531 5687 9537
rect 6454 9528 6460 9540
rect 6512 9528 6518 9580
rect 6549 9571 6607 9577
rect 6549 9537 6561 9571
rect 6595 9568 6607 9571
rect 7834 9568 7840 9580
rect 6595 9540 7840 9568
rect 6595 9537 6607 9540
rect 6549 9531 6607 9537
rect 2774 9500 2780 9512
rect 2516 9472 2780 9500
rect 2774 9460 2780 9472
rect 2832 9460 2838 9512
rect 4522 9460 4528 9512
rect 4580 9500 4586 9512
rect 6564 9500 6592 9531
rect 7834 9528 7840 9540
rect 7892 9528 7898 9580
rect 8754 9568 8760 9580
rect 8715 9540 8760 9568
rect 8754 9528 8760 9540
rect 8812 9528 8818 9580
rect 9858 9528 9864 9580
rect 9916 9568 9922 9580
rect 9953 9571 10011 9577
rect 9953 9568 9965 9571
rect 9916 9540 9965 9568
rect 9916 9528 9922 9540
rect 9953 9537 9965 9540
rect 9999 9537 10011 9571
rect 10686 9568 10692 9580
rect 10647 9540 10692 9568
rect 9953 9531 10011 9537
rect 10686 9528 10692 9540
rect 10744 9568 10750 9580
rect 17144 9577 17172 9608
rect 17310 9596 17316 9608
rect 17368 9596 17374 9648
rect 23201 9639 23259 9645
rect 19260 9608 22094 9636
rect 11701 9571 11759 9577
rect 11701 9568 11713 9571
rect 10744 9540 11713 9568
rect 10744 9528 10750 9540
rect 11701 9537 11713 9540
rect 11747 9568 11759 9571
rect 12897 9571 12955 9577
rect 12897 9568 12909 9571
rect 11747 9540 12909 9568
rect 11747 9537 11759 9540
rect 11701 9531 11759 9537
rect 12897 9537 12909 9540
rect 12943 9568 12955 9571
rect 14737 9571 14795 9577
rect 14737 9568 14749 9571
rect 12943 9540 14749 9568
rect 12943 9537 12955 9540
rect 12897 9531 12955 9537
rect 14737 9537 14749 9540
rect 14783 9568 14795 9571
rect 15565 9571 15623 9577
rect 15565 9568 15577 9571
rect 14783 9540 15577 9568
rect 14783 9537 14795 9540
rect 14737 9531 14795 9537
rect 15565 9537 15577 9540
rect 15611 9537 15623 9571
rect 15565 9531 15623 9537
rect 17129 9571 17187 9577
rect 17129 9537 17141 9571
rect 17175 9537 17187 9571
rect 17402 9568 17408 9580
rect 17363 9540 17408 9568
rect 17129 9531 17187 9537
rect 17402 9528 17408 9540
rect 17460 9528 17466 9580
rect 19260 9577 19288 9608
rect 19245 9571 19303 9577
rect 19245 9537 19257 9571
rect 19291 9537 19303 9571
rect 19245 9531 19303 9537
rect 20070 9528 20076 9580
rect 20128 9568 20134 9580
rect 20625 9571 20683 9577
rect 20625 9568 20637 9571
rect 20128 9540 20637 9568
rect 20128 9528 20134 9540
rect 20625 9537 20637 9540
rect 20671 9537 20683 9571
rect 20898 9568 20904 9580
rect 20859 9540 20904 9568
rect 20625 9531 20683 9537
rect 20898 9528 20904 9540
rect 20956 9528 20962 9580
rect 22066 9568 22094 9608
rect 23201 9605 23213 9639
rect 23247 9636 23259 9639
rect 23474 9636 23480 9648
rect 23247 9608 23480 9636
rect 23247 9605 23259 9608
rect 23201 9599 23259 9605
rect 23474 9596 23480 9608
rect 23532 9596 23538 9648
rect 23753 9639 23811 9645
rect 23753 9605 23765 9639
rect 23799 9636 23811 9639
rect 30558 9636 30564 9648
rect 23799 9608 28764 9636
rect 23799 9605 23811 9608
rect 23753 9599 23811 9605
rect 22189 9571 22247 9577
rect 22189 9568 22201 9571
rect 22066 9540 22201 9568
rect 22189 9537 22201 9540
rect 22235 9568 22247 9571
rect 23017 9571 23075 9577
rect 23017 9568 23029 9571
rect 22235 9540 23029 9568
rect 22235 9537 22247 9540
rect 22189 9531 22247 9537
rect 23017 9537 23029 9540
rect 23063 9568 23075 9571
rect 23290 9568 23296 9580
rect 23063 9540 23296 9568
rect 23063 9537 23075 9540
rect 23017 9531 23075 9537
rect 23290 9528 23296 9540
rect 23348 9528 23354 9580
rect 25056 9577 25084 9608
rect 24397 9571 24455 9577
rect 24397 9537 24409 9571
rect 24443 9537 24455 9571
rect 24397 9531 24455 9537
rect 25041 9571 25099 9577
rect 25041 9537 25053 9571
rect 25087 9537 25099 9571
rect 25222 9568 25228 9580
rect 25183 9540 25228 9568
rect 25041 9531 25099 9537
rect 4580 9472 6592 9500
rect 6733 9503 6791 9509
rect 4580 9460 4586 9472
rect 6733 9469 6745 9503
rect 6779 9500 6791 9503
rect 6822 9500 6828 9512
rect 6779 9472 6828 9500
rect 6779 9469 6791 9472
rect 6733 9463 6791 9469
rect 6822 9460 6828 9472
rect 6880 9460 6886 9512
rect 7926 9460 7932 9512
rect 7984 9500 7990 9512
rect 8021 9503 8079 9509
rect 8021 9500 8033 9503
rect 7984 9472 8033 9500
rect 7984 9460 7990 9472
rect 8021 9469 8033 9472
rect 8067 9469 8079 9503
rect 8021 9463 8079 9469
rect 8481 9503 8539 9509
rect 8481 9469 8493 9503
rect 8527 9469 8539 9503
rect 8481 9463 8539 9469
rect 10873 9503 10931 9509
rect 10873 9469 10885 9503
rect 10919 9500 10931 9503
rect 10962 9500 10968 9512
rect 10919 9472 10968 9500
rect 10919 9469 10931 9472
rect 10873 9463 10931 9469
rect 5074 9432 5080 9444
rect 3988 9404 5080 9432
rect 1949 9367 2007 9373
rect 1949 9333 1961 9367
rect 1995 9364 2007 9367
rect 3988 9364 4016 9404
rect 5074 9392 5080 9404
rect 5132 9392 5138 9444
rect 5813 9435 5871 9441
rect 5813 9401 5825 9435
rect 5859 9432 5871 9435
rect 7374 9432 7380 9444
rect 5859 9404 7380 9432
rect 5859 9401 5871 9404
rect 5813 9395 5871 9401
rect 7374 9392 7380 9404
rect 7432 9432 7438 9444
rect 8496 9432 8524 9463
rect 10962 9460 10968 9472
rect 11020 9460 11026 9512
rect 11885 9503 11943 9509
rect 11885 9469 11897 9503
rect 11931 9469 11943 9503
rect 12710 9500 12716 9512
rect 12671 9472 12716 9500
rect 11885 9463 11943 9469
rect 11900 9432 11928 9463
rect 12710 9460 12716 9472
rect 12768 9460 12774 9512
rect 14550 9500 14556 9512
rect 14511 9472 14556 9500
rect 14550 9460 14556 9472
rect 14608 9460 14614 9512
rect 15378 9500 15384 9512
rect 15339 9472 15384 9500
rect 15378 9460 15384 9472
rect 15436 9460 15442 9512
rect 15470 9460 15476 9512
rect 15528 9500 15534 9512
rect 16942 9500 16948 9512
rect 15528 9472 16948 9500
rect 15528 9460 15534 9472
rect 16942 9460 16948 9472
rect 17000 9460 17006 9512
rect 18966 9460 18972 9512
rect 19024 9500 19030 9512
rect 19061 9503 19119 9509
rect 19061 9500 19073 9503
rect 19024 9472 19073 9500
rect 19024 9460 19030 9472
rect 19061 9469 19073 9472
rect 19107 9469 19119 9503
rect 22005 9503 22063 9509
rect 22005 9500 22017 9503
rect 19061 9463 19119 9469
rect 21376 9472 22017 9500
rect 14182 9432 14188 9444
rect 7432 9404 8524 9432
rect 9416 9404 14188 9432
rect 7432 9392 7438 9404
rect 1995 9336 4016 9364
rect 4985 9367 5043 9373
rect 1995 9333 2007 9336
rect 1949 9327 2007 9333
rect 4985 9333 4997 9367
rect 5031 9364 5043 9367
rect 5626 9364 5632 9376
rect 5031 9336 5632 9364
rect 5031 9333 5043 9336
rect 4985 9327 5043 9333
rect 5626 9324 5632 9336
rect 5684 9324 5690 9376
rect 6730 9324 6736 9376
rect 6788 9364 6794 9376
rect 7653 9367 7711 9373
rect 7653 9364 7665 9367
rect 6788 9336 7665 9364
rect 6788 9324 6794 9336
rect 7653 9333 7665 9336
rect 7699 9333 7711 9367
rect 7653 9327 7711 9333
rect 7926 9324 7932 9376
rect 7984 9364 7990 9376
rect 9416 9364 9444 9404
rect 14182 9392 14188 9404
rect 14240 9392 14246 9444
rect 7984 9336 9444 9364
rect 9493 9367 9551 9373
rect 7984 9324 7990 9336
rect 9493 9333 9505 9367
rect 9539 9364 9551 9367
rect 9766 9364 9772 9376
rect 9539 9336 9772 9364
rect 9539 9333 9551 9336
rect 9493 9327 9551 9333
rect 9766 9324 9772 9336
rect 9824 9364 9830 9376
rect 10594 9364 10600 9376
rect 9824 9336 10600 9364
rect 9824 9324 9830 9336
rect 10594 9324 10600 9336
rect 10652 9324 10658 9376
rect 14093 9367 14151 9373
rect 14093 9333 14105 9367
rect 14139 9364 14151 9367
rect 14366 9364 14372 9376
rect 14139 9336 14372 9364
rect 14139 9333 14151 9336
rect 14093 9327 14151 9333
rect 14366 9324 14372 9336
rect 14424 9324 14430 9376
rect 14568 9364 14596 9460
rect 15194 9392 15200 9444
rect 15252 9432 15258 9444
rect 16482 9432 16488 9444
rect 15252 9404 16488 9432
rect 15252 9392 15258 9404
rect 16482 9392 16488 9404
rect 16540 9432 16546 9444
rect 17126 9432 17132 9444
rect 16540 9404 17132 9432
rect 16540 9392 16546 9404
rect 17126 9392 17132 9404
rect 17184 9392 17190 9444
rect 19306 9404 20392 9432
rect 19306 9364 19334 9404
rect 14568 9336 19334 9364
rect 19429 9367 19487 9373
rect 19429 9333 19441 9367
rect 19475 9364 19487 9367
rect 19610 9364 19616 9376
rect 19475 9336 19616 9364
rect 19475 9333 19487 9336
rect 19429 9327 19487 9333
rect 19610 9324 19616 9336
rect 19668 9324 19674 9376
rect 19886 9324 19892 9376
rect 19944 9364 19950 9376
rect 20254 9364 20260 9376
rect 19944 9336 20260 9364
rect 19944 9324 19950 9336
rect 20254 9324 20260 9336
rect 20312 9324 20318 9376
rect 20364 9364 20392 9404
rect 21376 9364 21404 9472
rect 22005 9469 22017 9472
rect 22051 9500 22063 9503
rect 22094 9500 22100 9512
rect 22051 9472 22100 9500
rect 22051 9469 22063 9472
rect 22005 9463 22063 9469
rect 22094 9460 22100 9472
rect 22152 9460 22158 9512
rect 22462 9460 22468 9512
rect 22520 9500 22526 9512
rect 22833 9503 22891 9509
rect 22833 9500 22845 9503
rect 22520 9472 22845 9500
rect 22520 9460 22526 9472
rect 22833 9469 22845 9472
rect 22879 9469 22891 9503
rect 22833 9463 22891 9469
rect 22848 9432 22876 9463
rect 23014 9432 23020 9444
rect 22848 9404 23020 9432
rect 23014 9392 23020 9404
rect 23072 9392 23078 9444
rect 24412 9432 24440 9531
rect 25222 9528 25228 9540
rect 25280 9528 25286 9580
rect 26050 9568 26056 9580
rect 26011 9540 26056 9568
rect 26050 9528 26056 9540
rect 26108 9528 26114 9580
rect 26234 9568 26240 9580
rect 26195 9540 26240 9568
rect 26234 9528 26240 9540
rect 26292 9528 26298 9580
rect 26326 9528 26332 9580
rect 26384 9568 26390 9580
rect 27249 9571 27307 9577
rect 27249 9568 27261 9571
rect 26384 9540 27261 9568
rect 26384 9528 26390 9540
rect 27249 9537 27261 9540
rect 27295 9537 27307 9571
rect 28442 9568 28448 9580
rect 28403 9540 28448 9568
rect 27249 9531 27307 9537
rect 28442 9528 28448 9540
rect 28500 9528 28506 9580
rect 28629 9571 28687 9577
rect 28629 9537 28641 9571
rect 28675 9537 28687 9571
rect 28736 9568 28764 9608
rect 29288 9608 30564 9636
rect 28994 9568 29000 9580
rect 28736 9540 29000 9568
rect 28629 9531 28687 9537
rect 26970 9500 26976 9512
rect 26931 9472 26976 9500
rect 26970 9460 26976 9472
rect 27028 9460 27034 9512
rect 24412 9404 25268 9432
rect 20364 9336 21404 9364
rect 22278 9324 22284 9376
rect 22336 9364 22342 9376
rect 25038 9364 25044 9376
rect 22336 9336 25044 9364
rect 22336 9324 22342 9336
rect 25038 9324 25044 9336
rect 25096 9324 25102 9376
rect 25240 9373 25268 9404
rect 25225 9367 25283 9373
rect 25225 9333 25237 9367
rect 25271 9364 25283 9367
rect 25682 9364 25688 9376
rect 25271 9336 25688 9364
rect 25271 9333 25283 9336
rect 25225 9327 25283 9333
rect 25682 9324 25688 9336
rect 25740 9324 25746 9376
rect 28644 9364 28672 9531
rect 28994 9528 29000 9540
rect 29052 9528 29058 9580
rect 29288 9577 29316 9608
rect 30558 9596 30564 9608
rect 30616 9596 30622 9648
rect 31754 9596 31760 9648
rect 31812 9636 31818 9648
rect 31812 9608 35480 9636
rect 31812 9596 31818 9608
rect 29273 9571 29331 9577
rect 29273 9537 29285 9571
rect 29319 9537 29331 9571
rect 29546 9568 29552 9580
rect 29507 9540 29552 9568
rect 29273 9531 29331 9537
rect 29546 9528 29552 9540
rect 29604 9528 29610 9580
rect 29638 9528 29644 9580
rect 29696 9568 29702 9580
rect 30742 9568 30748 9580
rect 29696 9540 30512 9568
rect 30703 9540 30748 9568
rect 29696 9528 29702 9540
rect 28810 9500 28816 9512
rect 28771 9472 28816 9500
rect 28810 9460 28816 9472
rect 28868 9460 28874 9512
rect 30484 9500 30512 9540
rect 30742 9528 30748 9540
rect 30800 9528 30806 9580
rect 31570 9528 31576 9580
rect 31628 9568 31634 9580
rect 32125 9571 32183 9577
rect 32125 9568 32137 9571
rect 31628 9540 32137 9568
rect 31628 9528 31634 9540
rect 32125 9537 32137 9540
rect 32171 9537 32183 9571
rect 32125 9531 32183 9537
rect 32950 9528 32956 9580
rect 33008 9568 33014 9580
rect 33045 9571 33103 9577
rect 33045 9568 33057 9571
rect 33008 9540 33057 9568
rect 33008 9528 33014 9540
rect 33045 9537 33057 9540
rect 33091 9537 33103 9571
rect 34974 9568 34980 9580
rect 34935 9540 34980 9568
rect 33045 9531 33103 9537
rect 34974 9528 34980 9540
rect 35032 9528 35038 9580
rect 35066 9528 35072 9580
rect 35124 9568 35130 9580
rect 35253 9571 35311 9577
rect 35253 9568 35265 9571
rect 35124 9540 35265 9568
rect 35124 9528 35130 9540
rect 35253 9537 35265 9540
rect 35299 9537 35311 9571
rect 35253 9531 35311 9537
rect 35452 9568 35480 9608
rect 36280 9568 36308 9676
rect 37366 9664 37372 9676
rect 37424 9664 37430 9716
rect 38010 9704 38016 9716
rect 37660 9676 38016 9704
rect 36446 9568 36452 9580
rect 35452 9540 36308 9568
rect 36407 9540 36452 9568
rect 32766 9500 32772 9512
rect 30484 9472 31754 9500
rect 32727 9472 32772 9500
rect 31294 9432 31300 9444
rect 29840 9404 31300 9432
rect 28810 9364 28816 9376
rect 28644 9336 28816 9364
rect 28810 9324 28816 9336
rect 28868 9364 28874 9376
rect 29840 9364 29868 9404
rect 31294 9392 31300 9404
rect 31352 9392 31358 9444
rect 28868 9336 29868 9364
rect 28868 9324 28874 9336
rect 30006 9324 30012 9376
rect 30064 9364 30070 9376
rect 30282 9364 30288 9376
rect 30064 9336 30288 9364
rect 30064 9324 30070 9336
rect 30282 9324 30288 9336
rect 30340 9324 30346 9376
rect 31110 9324 31116 9376
rect 31168 9364 31174 9376
rect 31389 9367 31447 9373
rect 31389 9364 31401 9367
rect 31168 9336 31401 9364
rect 31168 9324 31174 9336
rect 31389 9333 31401 9336
rect 31435 9333 31447 9367
rect 31726 9364 31754 9472
rect 32766 9460 32772 9472
rect 32824 9460 32830 9512
rect 35452 9432 35480 9540
rect 36446 9528 36452 9540
rect 36504 9528 36510 9580
rect 36725 9571 36783 9577
rect 36725 9537 36737 9571
rect 36771 9568 36783 9571
rect 37660 9568 37688 9676
rect 38010 9664 38016 9676
rect 38068 9664 38074 9716
rect 38102 9664 38108 9716
rect 38160 9704 38166 9716
rect 38381 9707 38439 9713
rect 38381 9704 38393 9707
rect 38160 9676 38393 9704
rect 38160 9664 38166 9676
rect 38381 9673 38393 9676
rect 38427 9673 38439 9707
rect 38381 9667 38439 9673
rect 39209 9707 39267 9713
rect 39209 9673 39221 9707
rect 39255 9673 39267 9707
rect 39209 9667 39267 9673
rect 37737 9639 37795 9645
rect 37737 9605 37749 9639
rect 37783 9636 37795 9639
rect 38654 9636 38660 9648
rect 37783 9608 38660 9636
rect 37783 9605 37795 9608
rect 37737 9599 37795 9605
rect 38654 9596 38660 9608
rect 38712 9596 38718 9648
rect 39224 9636 39252 9667
rect 42978 9664 42984 9716
rect 43036 9704 43042 9716
rect 43901 9707 43959 9713
rect 43901 9704 43913 9707
rect 43036 9676 43913 9704
rect 43036 9664 43042 9676
rect 43901 9673 43913 9676
rect 43947 9673 43959 9707
rect 46474 9704 46480 9716
rect 46435 9676 46480 9704
rect 43901 9667 43959 9673
rect 46474 9664 46480 9676
rect 46532 9664 46538 9716
rect 47670 9664 47676 9716
rect 47728 9704 47734 9716
rect 47765 9707 47823 9713
rect 47765 9704 47777 9707
rect 47728 9676 47777 9704
rect 47728 9664 47734 9676
rect 47765 9673 47777 9676
rect 47811 9673 47823 9707
rect 47765 9667 47823 9673
rect 41601 9639 41659 9645
rect 39224 9608 41552 9636
rect 38562 9568 38568 9580
rect 36771 9540 37688 9568
rect 38523 9540 38568 9568
rect 36771 9537 36783 9540
rect 36725 9531 36783 9537
rect 38562 9528 38568 9540
rect 38620 9528 38626 9580
rect 37366 9460 37372 9512
rect 37424 9500 37430 9512
rect 39224 9500 39252 9608
rect 39942 9568 39948 9580
rect 39903 9540 39948 9568
rect 39942 9528 39948 9540
rect 40000 9528 40006 9580
rect 40218 9568 40224 9580
rect 40179 9540 40224 9568
rect 40218 9528 40224 9540
rect 40276 9528 40282 9580
rect 40310 9528 40316 9580
rect 40368 9568 40374 9580
rect 41417 9571 41475 9577
rect 41417 9568 41429 9571
rect 40368 9540 41429 9568
rect 40368 9528 40374 9540
rect 41417 9537 41429 9540
rect 41463 9537 41475 9571
rect 41417 9531 41475 9537
rect 41230 9500 41236 9512
rect 37424 9472 39252 9500
rect 41191 9472 41236 9500
rect 37424 9460 37430 9472
rect 41230 9460 41236 9472
rect 41288 9460 41294 9512
rect 35713 9435 35771 9441
rect 35713 9432 35725 9435
rect 35452 9404 35725 9432
rect 35713 9401 35725 9404
rect 35759 9401 35771 9435
rect 35713 9395 35771 9401
rect 38102 9392 38108 9444
rect 38160 9432 38166 9444
rect 38160 9404 39344 9432
rect 38160 9392 38166 9404
rect 37829 9367 37887 9373
rect 37829 9364 37841 9367
rect 31726 9336 37841 9364
rect 31389 9327 31447 9333
rect 37829 9333 37841 9336
rect 37875 9364 37887 9367
rect 38838 9364 38844 9376
rect 37875 9336 38844 9364
rect 37875 9333 37887 9336
rect 37829 9327 37887 9333
rect 38838 9324 38844 9336
rect 38896 9324 38902 9376
rect 39316 9364 39344 9404
rect 40681 9367 40739 9373
rect 40681 9364 40693 9367
rect 39316 9336 40693 9364
rect 40681 9333 40693 9336
rect 40727 9333 40739 9367
rect 41524 9364 41552 9608
rect 41601 9605 41613 9639
rect 41647 9636 41659 9639
rect 41647 9608 44128 9636
rect 41647 9605 41659 9608
rect 41601 9599 41659 9605
rect 42150 9528 42156 9580
rect 42208 9568 42214 9580
rect 44100 9577 44128 9608
rect 44174 9596 44180 9648
rect 44232 9636 44238 9648
rect 45462 9636 45468 9648
rect 44232 9608 45468 9636
rect 44232 9596 44238 9608
rect 45462 9596 45468 9608
rect 45520 9636 45526 9648
rect 50522 9636 50528 9648
rect 45520 9608 45876 9636
rect 50483 9608 50528 9636
rect 45520 9596 45526 9608
rect 42705 9571 42763 9577
rect 42705 9568 42717 9571
rect 42208 9540 42717 9568
rect 42208 9528 42214 9540
rect 42705 9537 42717 9540
rect 42751 9537 42763 9571
rect 42705 9531 42763 9537
rect 44085 9571 44143 9577
rect 44085 9537 44097 9571
rect 44131 9537 44143 9571
rect 44634 9568 44640 9580
rect 44595 9540 44640 9568
rect 44085 9531 44143 9537
rect 44634 9528 44640 9540
rect 44692 9528 44698 9580
rect 45002 9528 45008 9580
rect 45060 9568 45066 9580
rect 45848 9577 45876 9608
rect 50522 9596 50528 9608
rect 50580 9596 50586 9648
rect 53374 9636 53380 9648
rect 51046 9608 53380 9636
rect 45649 9571 45707 9577
rect 45649 9568 45661 9571
rect 45060 9540 45661 9568
rect 45060 9528 45066 9540
rect 45649 9537 45661 9540
rect 45695 9537 45707 9571
rect 45649 9531 45707 9537
rect 45833 9571 45891 9577
rect 45833 9537 45845 9571
rect 45879 9537 45891 9571
rect 46658 9568 46664 9580
rect 46619 9540 46664 9568
rect 45833 9531 45891 9537
rect 46658 9528 46664 9540
rect 46716 9528 46722 9580
rect 47581 9571 47639 9577
rect 47581 9537 47593 9571
rect 47627 9537 47639 9571
rect 47581 9531 47639 9537
rect 42426 9500 42432 9512
rect 42387 9472 42432 9500
rect 42426 9460 42432 9472
rect 42484 9460 42490 9512
rect 46017 9503 46075 9509
rect 46017 9469 46029 9503
rect 46063 9500 46075 9503
rect 47596 9500 47624 9531
rect 48130 9528 48136 9580
rect 48188 9568 48194 9580
rect 48317 9571 48375 9577
rect 48317 9568 48329 9571
rect 48188 9540 48329 9568
rect 48188 9528 48194 9540
rect 48317 9537 48329 9540
rect 48363 9537 48375 9571
rect 49237 9571 49295 9577
rect 49237 9568 49249 9571
rect 48317 9531 48375 9537
rect 48516 9540 49249 9568
rect 46063 9472 47624 9500
rect 46063 9469 46075 9472
rect 46017 9463 46075 9469
rect 44821 9435 44879 9441
rect 44821 9401 44833 9435
rect 44867 9432 44879 9435
rect 46750 9432 46756 9444
rect 44867 9404 46756 9432
rect 44867 9401 44879 9404
rect 44821 9395 44879 9401
rect 46750 9392 46756 9404
rect 46808 9392 46814 9444
rect 48516 9441 48544 9540
rect 49237 9537 49249 9540
rect 49283 9537 49295 9571
rect 50062 9568 50068 9580
rect 50023 9540 50068 9568
rect 49237 9531 49295 9537
rect 50062 9528 50068 9540
rect 50120 9568 50126 9580
rect 51046 9568 51074 9608
rect 53374 9596 53380 9608
rect 53432 9636 53438 9648
rect 53770 9639 53828 9645
rect 53770 9636 53782 9639
rect 53432 9608 53782 9636
rect 53432 9596 53438 9608
rect 53770 9605 53782 9608
rect 53816 9605 53828 9639
rect 53770 9599 53828 9605
rect 50120 9540 51074 9568
rect 50120 9528 50126 9540
rect 51258 9528 51264 9580
rect 51316 9568 51322 9580
rect 51353 9571 51411 9577
rect 51353 9568 51365 9571
rect 51316 9540 51365 9568
rect 51316 9528 51322 9540
rect 51353 9537 51365 9540
rect 51399 9537 51411 9571
rect 51994 9568 52000 9580
rect 51955 9540 52000 9568
rect 51353 9531 51411 9537
rect 51994 9528 52000 9540
rect 52052 9528 52058 9580
rect 53009 9571 53067 9577
rect 53009 9568 53021 9571
rect 52196 9540 53021 9568
rect 48958 9500 48964 9512
rect 48919 9472 48964 9500
rect 48958 9460 48964 9472
rect 49016 9460 49022 9512
rect 49694 9460 49700 9512
rect 49752 9500 49758 9512
rect 50522 9500 50528 9512
rect 49752 9472 50528 9500
rect 49752 9460 49758 9472
rect 50522 9460 50528 9472
rect 50580 9500 50586 9512
rect 51442 9500 51448 9512
rect 50580 9472 51448 9500
rect 50580 9460 50586 9472
rect 51442 9460 51448 9472
rect 51500 9460 51506 9512
rect 52196 9441 52224 9540
rect 53009 9537 53021 9540
rect 53055 9537 53067 9571
rect 53009 9531 53067 9537
rect 52270 9460 52276 9512
rect 52328 9500 52334 9512
rect 52733 9503 52791 9509
rect 52733 9500 52745 9503
rect 52328 9472 52745 9500
rect 52328 9460 52334 9472
rect 52733 9469 52745 9472
rect 52779 9469 52791 9503
rect 52733 9463 52791 9469
rect 48501 9435 48559 9441
rect 48501 9401 48513 9435
rect 48547 9401 48559 9435
rect 48501 9395 48559 9401
rect 52181 9435 52239 9441
rect 52181 9401 52193 9435
rect 52227 9401 52239 9435
rect 52181 9395 52239 9401
rect 42794 9364 42800 9376
rect 41524 9336 42800 9364
rect 40681 9327 40739 9333
rect 42794 9324 42800 9336
rect 42852 9364 42858 9376
rect 43441 9367 43499 9373
rect 43441 9364 43453 9367
rect 42852 9336 43453 9364
rect 42852 9324 42858 9336
rect 43441 9333 43453 9336
rect 43487 9364 43499 9367
rect 43714 9364 43720 9376
rect 43487 9336 43720 9364
rect 43487 9333 43499 9336
rect 43441 9327 43499 9333
rect 43714 9324 43720 9336
rect 43772 9324 43778 9376
rect 43990 9324 43996 9376
rect 44048 9364 44054 9376
rect 50522 9364 50528 9376
rect 44048 9336 50528 9364
rect 44048 9324 44054 9336
rect 50522 9324 50528 9336
rect 50580 9324 50586 9376
rect 51537 9367 51595 9373
rect 51537 9333 51549 9367
rect 51583 9364 51595 9367
rect 52546 9364 52552 9376
rect 51583 9336 52552 9364
rect 51583 9333 51595 9336
rect 51537 9327 51595 9333
rect 52546 9324 52552 9336
rect 52604 9324 52610 9376
rect 1104 9274 58880 9296
rect 1104 9222 8174 9274
rect 8226 9222 8238 9274
rect 8290 9222 8302 9274
rect 8354 9222 8366 9274
rect 8418 9222 8430 9274
rect 8482 9222 22622 9274
rect 22674 9222 22686 9274
rect 22738 9222 22750 9274
rect 22802 9222 22814 9274
rect 22866 9222 22878 9274
rect 22930 9222 37070 9274
rect 37122 9222 37134 9274
rect 37186 9222 37198 9274
rect 37250 9222 37262 9274
rect 37314 9222 37326 9274
rect 37378 9222 51518 9274
rect 51570 9222 51582 9274
rect 51634 9222 51646 9274
rect 51698 9222 51710 9274
rect 51762 9222 51774 9274
rect 51826 9222 58880 9274
rect 1104 9200 58880 9222
rect 2409 9163 2467 9169
rect 2409 9129 2421 9163
rect 2455 9160 2467 9163
rect 3510 9160 3516 9172
rect 2455 9132 3516 9160
rect 2455 9129 2467 9132
rect 2409 9123 2467 9129
rect 3510 9120 3516 9132
rect 3568 9120 3574 9172
rect 4157 9163 4215 9169
rect 4157 9129 4169 9163
rect 4203 9160 4215 9163
rect 4246 9160 4252 9172
rect 4203 9132 4252 9160
rect 4203 9129 4215 9132
rect 4157 9123 4215 9129
rect 4246 9120 4252 9132
rect 4304 9120 4310 9172
rect 6917 9163 6975 9169
rect 6917 9129 6929 9163
rect 6963 9160 6975 9163
rect 8754 9160 8760 9172
rect 6963 9132 8760 9160
rect 6963 9129 6975 9132
rect 6917 9123 6975 9129
rect 8754 9120 8760 9132
rect 8812 9120 8818 9172
rect 9309 9163 9367 9169
rect 9309 9129 9321 9163
rect 9355 9160 9367 9163
rect 10686 9160 10692 9172
rect 9355 9132 10692 9160
rect 9355 9129 9367 9132
rect 9309 9123 9367 9129
rect 10686 9120 10692 9132
rect 10744 9120 10750 9172
rect 12250 9160 12256 9172
rect 12211 9132 12256 9160
rect 12250 9120 12256 9132
rect 12308 9120 12314 9172
rect 12897 9163 12955 9169
rect 12897 9129 12909 9163
rect 12943 9160 12955 9163
rect 14550 9160 14556 9172
rect 12943 9132 14556 9160
rect 12943 9129 12955 9132
rect 12897 9123 12955 9129
rect 14550 9120 14556 9132
rect 14608 9120 14614 9172
rect 18230 9120 18236 9172
rect 18288 9160 18294 9172
rect 18601 9163 18659 9169
rect 18601 9160 18613 9163
rect 18288 9132 18613 9160
rect 18288 9120 18294 9132
rect 18601 9129 18613 9132
rect 18647 9129 18659 9163
rect 18601 9123 18659 9129
rect 19797 9163 19855 9169
rect 19797 9129 19809 9163
rect 19843 9129 19855 9163
rect 20257 9163 20315 9169
rect 20257 9160 20269 9163
rect 19797 9123 19855 9129
rect 20180 9132 20269 9160
rect 1673 9095 1731 9101
rect 1673 9061 1685 9095
rect 1719 9092 1731 9095
rect 3878 9092 3884 9104
rect 1719 9064 3884 9092
rect 1719 9061 1731 9064
rect 1673 9055 1731 9061
rect 2424 9036 2452 9064
rect 3878 9052 3884 9064
rect 3936 9052 3942 9104
rect 5629 9095 5687 9101
rect 5629 9061 5641 9095
rect 5675 9092 5687 9095
rect 5675 9064 7236 9092
rect 5675 9061 5687 9064
rect 5629 9055 5687 9061
rect 2406 8984 2412 9036
rect 2464 8984 2470 9036
rect 2958 8984 2964 9036
rect 3016 9024 3022 9036
rect 3237 9027 3295 9033
rect 3237 9024 3249 9027
rect 3016 8996 3249 9024
rect 3016 8984 3022 8996
rect 3237 8993 3249 8996
rect 3283 9024 3295 9027
rect 3418 9024 3424 9036
rect 3283 8996 3424 9024
rect 3283 8993 3295 8996
rect 3237 8987 3295 8993
rect 3418 8984 3424 8996
rect 3476 8984 3482 9036
rect 4062 8984 4068 9036
rect 4120 9024 4126 9036
rect 4617 9027 4675 9033
rect 4617 9024 4629 9027
rect 4120 8996 4629 9024
rect 4120 8984 4126 8996
rect 4617 8993 4629 8996
rect 4663 8993 4675 9027
rect 4617 8987 4675 8993
rect 1581 8959 1639 8965
rect 1581 8925 1593 8959
rect 1627 8925 1639 8959
rect 1581 8919 1639 8925
rect 1765 8959 1823 8965
rect 1765 8925 1777 8959
rect 1811 8956 1823 8959
rect 1946 8956 1952 8968
rect 1811 8928 1952 8956
rect 1811 8925 1823 8928
rect 1765 8919 1823 8925
rect 1596 8820 1624 8919
rect 1946 8916 1952 8928
rect 2004 8916 2010 8968
rect 2225 8959 2283 8965
rect 2225 8925 2237 8959
rect 2271 8956 2283 8959
rect 2869 8959 2927 8965
rect 2869 8956 2881 8959
rect 2271 8928 2881 8956
rect 2271 8925 2283 8928
rect 2225 8919 2283 8925
rect 2869 8925 2881 8928
rect 2915 8925 2927 8959
rect 2869 8919 2927 8925
rect 3050 8916 3056 8968
rect 3108 8956 3114 8968
rect 3108 8928 3201 8956
rect 3108 8916 3114 8928
rect 3786 8916 3792 8968
rect 3844 8956 3850 8968
rect 3973 8959 4031 8965
rect 3973 8956 3985 8959
rect 3844 8928 3985 8956
rect 3844 8916 3850 8928
rect 3973 8925 3985 8928
rect 4019 8925 4031 8959
rect 4890 8956 4896 8968
rect 4851 8928 4896 8956
rect 3973 8919 4031 8925
rect 4890 8916 4896 8928
rect 4948 8916 4954 8968
rect 6086 8956 6092 8968
rect 6047 8928 6092 8956
rect 6086 8916 6092 8928
rect 6144 8916 6150 8968
rect 6730 8956 6736 8968
rect 6691 8928 6736 8956
rect 6730 8916 6736 8928
rect 6788 8916 6794 8968
rect 7208 8956 7236 9064
rect 8018 9052 8024 9104
rect 8076 9092 8082 9104
rect 10413 9095 10471 9101
rect 10413 9092 10425 9095
rect 8076 9064 10425 9092
rect 8076 9052 8082 9064
rect 10413 9061 10425 9064
rect 10459 9061 10471 9095
rect 10413 9055 10471 9061
rect 15197 9095 15255 9101
rect 15197 9061 15209 9095
rect 15243 9092 15255 9095
rect 15562 9092 15568 9104
rect 15243 9064 15568 9092
rect 15243 9061 15255 9064
rect 15197 9055 15255 9061
rect 15562 9052 15568 9064
rect 15620 9052 15626 9104
rect 15841 9095 15899 9101
rect 15841 9061 15853 9095
rect 15887 9092 15899 9095
rect 16482 9092 16488 9104
rect 15887 9064 16488 9092
rect 15887 9061 15899 9064
rect 15841 9055 15899 9061
rect 16482 9052 16488 9064
rect 16540 9052 16546 9104
rect 19812 9092 19840 9123
rect 20070 9092 20076 9104
rect 16592 9064 17172 9092
rect 19812 9064 20076 9092
rect 7374 9024 7380 9036
rect 7335 8996 7380 9024
rect 7374 8984 7380 8996
rect 7432 8984 7438 9036
rect 16592 9024 16620 9064
rect 9784 8996 11100 9024
rect 7558 8956 7564 8968
rect 7208 8928 7564 8956
rect 7558 8916 7564 8928
rect 7616 8916 7622 8968
rect 9784 8965 9812 8996
rect 7653 8959 7711 8965
rect 7653 8925 7665 8959
rect 7699 8925 7711 8959
rect 7653 8919 7711 8925
rect 9125 8959 9183 8965
rect 9125 8925 9137 8959
rect 9171 8925 9183 8959
rect 9125 8919 9183 8925
rect 9769 8959 9827 8965
rect 9769 8925 9781 8959
rect 9815 8925 9827 8959
rect 10594 8956 10600 8968
rect 10555 8928 10600 8956
rect 9769 8919 9827 8925
rect 3068 8888 3096 8916
rect 4522 8888 4528 8900
rect 3068 8860 4528 8888
rect 4522 8848 4528 8860
rect 4580 8848 4586 8900
rect 7668 8888 7696 8919
rect 6288 8860 7696 8888
rect 9140 8888 9168 8919
rect 10594 8916 10600 8928
rect 10652 8916 10658 8968
rect 10781 8959 10839 8965
rect 10781 8925 10793 8959
rect 10827 8925 10839 8959
rect 10781 8919 10839 8925
rect 10612 8888 10640 8916
rect 9140 8860 10640 8888
rect 3326 8820 3332 8832
rect 1596 8792 3332 8820
rect 3326 8780 3332 8792
rect 3384 8780 3390 8832
rect 6288 8829 6316 8860
rect 6273 8823 6331 8829
rect 6273 8789 6285 8823
rect 6319 8789 6331 8823
rect 6273 8783 6331 8789
rect 7558 8780 7564 8832
rect 7616 8820 7622 8832
rect 8389 8823 8447 8829
rect 8389 8820 8401 8823
rect 7616 8792 8401 8820
rect 7616 8780 7622 8792
rect 8389 8789 8401 8792
rect 8435 8820 8447 8823
rect 9766 8820 9772 8832
rect 8435 8792 9772 8820
rect 8435 8789 8447 8792
rect 8389 8783 8447 8789
rect 9766 8780 9772 8792
rect 9824 8780 9830 8832
rect 9953 8823 10011 8829
rect 9953 8789 9965 8823
rect 9999 8820 10011 8823
rect 10594 8820 10600 8832
rect 9999 8792 10600 8820
rect 9999 8789 10011 8792
rect 9953 8783 10011 8789
rect 10594 8780 10600 8792
rect 10652 8780 10658 8832
rect 10796 8820 10824 8919
rect 11072 8888 11100 8996
rect 14844 8996 16620 9024
rect 14844 8968 14872 8996
rect 16666 8984 16672 9036
rect 16724 9024 16730 9036
rect 16724 8996 16769 9024
rect 16724 8984 16730 8996
rect 11241 8959 11299 8965
rect 11241 8925 11253 8959
rect 11287 8956 11299 8959
rect 11422 8956 11428 8968
rect 11287 8928 11428 8956
rect 11287 8925 11299 8928
rect 11241 8919 11299 8925
rect 11422 8916 11428 8928
rect 11480 8916 11486 8968
rect 11514 8916 11520 8968
rect 11572 8956 11578 8968
rect 12710 8956 12716 8968
rect 11572 8928 11617 8956
rect 12671 8928 12716 8956
rect 11572 8916 11578 8928
rect 12710 8916 12716 8928
rect 12768 8956 12774 8968
rect 13262 8956 13268 8968
rect 12768 8928 13268 8956
rect 12768 8916 12774 8928
rect 13262 8916 13268 8928
rect 13320 8916 13326 8968
rect 13357 8959 13415 8965
rect 13357 8925 13369 8959
rect 13403 8956 13415 8959
rect 13446 8956 13452 8968
rect 13403 8928 13452 8956
rect 13403 8925 13415 8928
rect 13357 8919 13415 8925
rect 13446 8916 13452 8928
rect 13504 8916 13510 8968
rect 14185 8959 14243 8965
rect 14185 8925 14197 8959
rect 14231 8925 14243 8959
rect 14458 8956 14464 8968
rect 14419 8928 14464 8956
rect 14185 8919 14243 8925
rect 13814 8888 13820 8900
rect 11072 8860 13820 8888
rect 13814 8848 13820 8860
rect 13872 8848 13878 8900
rect 14200 8888 14228 8919
rect 14458 8916 14464 8928
rect 14516 8916 14522 8968
rect 14826 8916 14832 8968
rect 14884 8916 14890 8968
rect 15657 8959 15715 8965
rect 15657 8925 15669 8959
rect 15703 8956 15715 8959
rect 16390 8956 16396 8968
rect 15703 8928 16396 8956
rect 15703 8925 15715 8928
rect 15657 8919 15715 8925
rect 16390 8916 16396 8928
rect 16448 8916 16454 8968
rect 16485 8959 16543 8965
rect 16485 8925 16497 8959
rect 16531 8956 16543 8959
rect 17034 8956 17040 8968
rect 16531 8928 17040 8956
rect 16531 8925 16543 8928
rect 16485 8919 16543 8925
rect 17034 8916 17040 8928
rect 17092 8916 17098 8968
rect 17144 8965 17172 9064
rect 20070 9052 20076 9064
rect 20128 9052 20134 9104
rect 17129 8959 17187 8965
rect 17129 8925 17141 8959
rect 17175 8925 17187 8959
rect 17402 8956 17408 8968
rect 17363 8928 17408 8956
rect 17129 8919 17187 8925
rect 14844 8888 14872 8916
rect 14200 8860 14872 8888
rect 14918 8848 14924 8900
rect 14976 8888 14982 8900
rect 16301 8891 16359 8897
rect 16301 8888 16313 8891
rect 14976 8860 16313 8888
rect 14976 8848 14982 8860
rect 16301 8857 16313 8860
rect 16347 8857 16359 8891
rect 17144 8888 17172 8919
rect 17402 8916 17408 8928
rect 17460 8916 17466 8968
rect 19610 8956 19616 8968
rect 19571 8928 19616 8956
rect 19610 8916 19616 8928
rect 19668 8916 19674 8968
rect 19702 8916 19708 8968
rect 19760 8956 19766 8968
rect 20180 8956 20208 9132
rect 20257 9129 20269 9132
rect 20303 9129 20315 9163
rect 20257 9123 20315 9129
rect 20714 9120 20720 9172
rect 20772 9160 20778 9172
rect 21910 9160 21916 9172
rect 20772 9132 21916 9160
rect 20772 9120 20778 9132
rect 21910 9120 21916 9132
rect 21968 9120 21974 9172
rect 26326 9160 26332 9172
rect 22066 9132 26188 9160
rect 26287 9132 26332 9160
rect 21818 9092 21824 9104
rect 21779 9064 21824 9092
rect 21818 9052 21824 9064
rect 21876 9052 21882 9104
rect 20254 8984 20260 9036
rect 20312 9024 20318 9036
rect 20625 9027 20683 9033
rect 20625 9024 20637 9027
rect 20312 8996 20637 9024
rect 20312 8984 20318 8996
rect 20625 8993 20637 8996
rect 20671 9024 20683 9027
rect 20671 8996 21772 9024
rect 20671 8993 20683 8996
rect 20625 8987 20683 8993
rect 20438 8956 20444 8968
rect 19760 8928 20208 8956
rect 20399 8928 20444 8956
rect 19760 8916 19766 8928
rect 20438 8916 20444 8928
rect 20496 8916 20502 8968
rect 21634 8956 21640 8968
rect 21595 8928 21640 8956
rect 21634 8916 21640 8928
rect 21692 8916 21698 8968
rect 21744 8956 21772 8996
rect 22066 8956 22094 9132
rect 25041 9095 25099 9101
rect 25041 9061 25053 9095
rect 25087 9061 25099 9095
rect 25682 9092 25688 9104
rect 25643 9064 25688 9092
rect 25041 9055 25099 9061
rect 22278 9024 22284 9036
rect 22239 8996 22284 9024
rect 22278 8984 22284 8996
rect 22336 8984 22342 9036
rect 24394 8984 24400 9036
rect 24452 9024 24458 9036
rect 24452 8996 24992 9024
rect 24452 8984 24458 8996
rect 22557 8959 22615 8965
rect 22557 8958 22569 8959
rect 21744 8928 22094 8956
rect 22388 8930 22569 8958
rect 20070 8888 20076 8900
rect 17144 8860 20076 8888
rect 16301 8851 16359 8857
rect 20070 8848 20076 8860
rect 20128 8888 20134 8900
rect 20714 8888 20720 8900
rect 20128 8860 20720 8888
rect 20128 8848 20134 8860
rect 20714 8848 20720 8860
rect 20772 8848 20778 8900
rect 20824 8860 21312 8888
rect 11790 8820 11796 8832
rect 10796 8792 11796 8820
rect 11790 8780 11796 8792
rect 11848 8780 11854 8832
rect 13446 8820 13452 8832
rect 13407 8792 13452 8820
rect 13446 8780 13452 8792
rect 13504 8780 13510 8832
rect 13538 8780 13544 8832
rect 13596 8820 13602 8832
rect 15470 8820 15476 8832
rect 13596 8792 15476 8820
rect 13596 8780 13602 8792
rect 15470 8780 15476 8792
rect 15528 8780 15534 8832
rect 15562 8780 15568 8832
rect 15620 8820 15626 8832
rect 16206 8820 16212 8832
rect 15620 8792 16212 8820
rect 15620 8780 15626 8792
rect 16206 8780 16212 8792
rect 16264 8820 16270 8832
rect 18141 8823 18199 8829
rect 18141 8820 18153 8823
rect 16264 8792 18153 8820
rect 16264 8780 16270 8792
rect 18141 8789 18153 8792
rect 18187 8820 18199 8823
rect 20824 8820 20852 8860
rect 21284 8832 21312 8860
rect 21818 8848 21824 8900
rect 21876 8888 21882 8900
rect 22388 8888 22416 8930
rect 22557 8925 22569 8930
rect 22603 8925 22615 8959
rect 24854 8956 24860 8968
rect 24815 8928 24860 8956
rect 22557 8919 22615 8925
rect 24854 8916 24860 8928
rect 24912 8916 24918 8968
rect 21876 8860 22416 8888
rect 21876 8848 21882 8860
rect 21174 8820 21180 8832
rect 18187 8792 20852 8820
rect 21135 8792 21180 8820
rect 18187 8789 18199 8792
rect 18141 8783 18199 8789
rect 21174 8780 21180 8792
rect 21232 8780 21238 8832
rect 21266 8780 21272 8832
rect 21324 8820 21330 8832
rect 23290 8820 23296 8832
rect 21324 8792 23296 8820
rect 21324 8780 21330 8792
rect 23290 8780 23296 8792
rect 23348 8780 23354 8832
rect 23474 8780 23480 8832
rect 23532 8820 23538 8832
rect 23658 8820 23664 8832
rect 23532 8792 23664 8820
rect 23532 8780 23538 8792
rect 23658 8780 23664 8792
rect 23716 8780 23722 8832
rect 23845 8823 23903 8829
rect 23845 8789 23857 8823
rect 23891 8820 23903 8823
rect 23934 8820 23940 8832
rect 23891 8792 23940 8820
rect 23891 8789 23903 8792
rect 23845 8783 23903 8789
rect 23934 8780 23940 8792
rect 23992 8780 23998 8832
rect 24964 8820 24992 8996
rect 25056 8956 25084 9055
rect 25682 9052 25688 9064
rect 25740 9052 25746 9104
rect 26160 9092 26188 9132
rect 26326 9120 26332 9132
rect 26384 9120 26390 9172
rect 28997 9163 29055 9169
rect 28997 9129 29009 9163
rect 29043 9160 29055 9163
rect 30742 9160 30748 9172
rect 29043 9132 30748 9160
rect 29043 9129 29055 9132
rect 28997 9123 29055 9129
rect 30742 9120 30748 9132
rect 30800 9120 30806 9172
rect 31570 9160 31576 9172
rect 31531 9132 31576 9160
rect 31570 9120 31576 9132
rect 31628 9120 31634 9172
rect 32950 9160 32956 9172
rect 32911 9132 32956 9160
rect 32950 9120 32956 9132
rect 33008 9120 33014 9172
rect 33042 9120 33048 9172
rect 33100 9160 33106 9172
rect 35253 9163 35311 9169
rect 35253 9160 35265 9163
rect 33100 9132 35265 9160
rect 33100 9120 33106 9132
rect 35253 9129 35265 9132
rect 35299 9129 35311 9163
rect 35253 9123 35311 9129
rect 35526 9120 35532 9172
rect 35584 9160 35590 9172
rect 37550 9160 37556 9172
rect 35584 9132 37556 9160
rect 35584 9120 35590 9132
rect 37550 9120 37556 9132
rect 37608 9120 37614 9172
rect 37737 9163 37795 9169
rect 37737 9129 37749 9163
rect 37783 9160 37795 9163
rect 38562 9160 38568 9172
rect 37783 9132 38568 9160
rect 37783 9129 37795 9132
rect 37737 9123 37795 9129
rect 38562 9120 38568 9132
rect 38620 9120 38626 9172
rect 38746 9120 38752 9172
rect 38804 9160 38810 9172
rect 42150 9160 42156 9172
rect 38804 9132 41414 9160
rect 42111 9132 42156 9160
rect 38804 9120 38810 9132
rect 32766 9092 32772 9104
rect 26160 9064 28994 9092
rect 26970 9024 26976 9036
rect 26068 8996 26976 9024
rect 25501 8959 25559 8965
rect 25501 8956 25513 8959
rect 25056 8928 25513 8956
rect 25501 8925 25513 8928
rect 25547 8956 25559 8959
rect 26068 8956 26096 8996
rect 26970 8984 26976 8996
rect 27028 8984 27034 9036
rect 25547 8928 26096 8956
rect 26145 8959 26203 8965
rect 25547 8925 25559 8928
rect 25501 8919 25559 8925
rect 26145 8925 26157 8959
rect 26191 8956 26203 8959
rect 27062 8956 27068 8968
rect 26191 8928 27068 8956
rect 26191 8925 26203 8928
rect 26145 8919 26203 8925
rect 27062 8916 27068 8928
rect 27120 8916 27126 8968
rect 27982 8956 27988 8968
rect 27943 8928 27988 8956
rect 27982 8916 27988 8928
rect 28040 8916 28046 8968
rect 28166 8956 28172 8968
rect 28127 8928 28172 8956
rect 28166 8916 28172 8928
rect 28224 8916 28230 8968
rect 28629 8959 28687 8965
rect 28629 8925 28641 8959
rect 28675 8956 28687 8959
rect 28810 8956 28816 8968
rect 28675 8928 28709 8956
rect 28771 8928 28816 8956
rect 28675 8925 28687 8928
rect 28629 8919 28687 8925
rect 25038 8848 25044 8900
rect 25096 8888 25102 8900
rect 25958 8888 25964 8900
rect 25096 8860 25964 8888
rect 25096 8848 25102 8860
rect 25958 8848 25964 8860
rect 26016 8848 26022 8900
rect 26234 8848 26240 8900
rect 26292 8888 26298 8900
rect 26789 8891 26847 8897
rect 26789 8888 26801 8891
rect 26292 8860 26801 8888
rect 26292 8848 26298 8860
rect 26789 8857 26801 8860
rect 26835 8857 26847 8891
rect 26970 8888 26976 8900
rect 26931 8860 26976 8888
rect 26789 8851 26847 8857
rect 26970 8848 26976 8860
rect 27028 8848 27034 8900
rect 27154 8888 27160 8900
rect 27115 8860 27160 8888
rect 27154 8848 27160 8860
rect 27212 8848 27218 8900
rect 28644 8888 28672 8919
rect 28810 8916 28816 8928
rect 28868 8916 28874 8968
rect 28966 8956 28994 9064
rect 30760 9064 32772 9092
rect 30469 8959 30527 8965
rect 28966 8928 30420 8956
rect 29454 8888 29460 8900
rect 27264 8860 29460 8888
rect 27264 8820 27292 8860
rect 29454 8848 29460 8860
rect 29512 8848 29518 8900
rect 24964 8792 27292 8820
rect 27430 8780 27436 8832
rect 27488 8820 27494 8832
rect 27985 8823 28043 8829
rect 27985 8820 27997 8823
rect 27488 8792 27997 8820
rect 27488 8780 27494 8792
rect 27985 8789 27997 8792
rect 28031 8820 28043 8823
rect 29178 8820 29184 8832
rect 28031 8792 29184 8820
rect 28031 8789 28043 8792
rect 27985 8783 28043 8789
rect 29178 8780 29184 8792
rect 29236 8780 29242 8832
rect 29546 8780 29552 8832
rect 29604 8820 29610 8832
rect 29733 8823 29791 8829
rect 29733 8820 29745 8823
rect 29604 8792 29745 8820
rect 29604 8780 29610 8792
rect 29733 8789 29745 8792
rect 29779 8820 29791 8823
rect 30006 8820 30012 8832
rect 29779 8792 30012 8820
rect 29779 8789 29791 8792
rect 29733 8783 29791 8789
rect 30006 8780 30012 8792
rect 30064 8780 30070 8832
rect 30392 8820 30420 8928
rect 30469 8925 30481 8959
rect 30515 8925 30527 8959
rect 30469 8919 30527 8925
rect 30484 8888 30512 8919
rect 30558 8916 30564 8968
rect 30616 8956 30622 8968
rect 30760 8965 30788 9064
rect 32766 9052 32772 9064
rect 32824 9092 32830 9104
rect 33413 9095 33471 9101
rect 33413 9092 33425 9095
rect 32824 9064 33425 9092
rect 32824 9052 32830 9064
rect 33413 9061 33425 9064
rect 33459 9061 33471 9095
rect 33413 9055 33471 9061
rect 33594 9052 33600 9104
rect 33652 9092 33658 9104
rect 34701 9095 34759 9101
rect 34701 9092 34713 9095
rect 33652 9064 34713 9092
rect 33652 9052 33658 9064
rect 34701 9061 34713 9064
rect 34747 9092 34759 9095
rect 36354 9092 36360 9104
rect 34747 9064 36360 9092
rect 34747 9061 34759 9064
rect 34701 9055 34759 9061
rect 36354 9052 36360 9064
rect 36412 9052 36418 9104
rect 36446 9052 36452 9104
rect 36504 9092 36510 9104
rect 38197 9095 38255 9101
rect 38197 9092 38209 9095
rect 36504 9064 38209 9092
rect 36504 9052 36510 9064
rect 38197 9061 38209 9064
rect 38243 9061 38255 9095
rect 38197 9055 38255 9061
rect 38838 9052 38844 9104
rect 38896 9092 38902 9104
rect 39758 9092 39764 9104
rect 38896 9064 39764 9092
rect 38896 9052 38902 9064
rect 39758 9052 39764 9064
rect 39816 9092 39822 9104
rect 41386 9092 41414 9132
rect 42150 9120 42156 9132
rect 42208 9120 42214 9172
rect 42613 9163 42671 9169
rect 42613 9129 42625 9163
rect 42659 9160 42671 9163
rect 42794 9160 42800 9172
rect 42659 9132 42800 9160
rect 42659 9129 42671 9132
rect 42613 9123 42671 9129
rect 42794 9120 42800 9132
rect 42852 9120 42858 9172
rect 44453 9163 44511 9169
rect 43088 9132 43668 9160
rect 43088 9092 43116 9132
rect 39816 9064 39896 9092
rect 41386 9064 43116 9092
rect 39816 9052 39822 9064
rect 34882 8984 34888 9036
rect 34940 9024 34946 9036
rect 39868 9033 39896 9064
rect 35345 9027 35403 9033
rect 35345 9024 35357 9027
rect 34940 8996 35357 9024
rect 34940 8984 34946 8996
rect 35345 8993 35357 8996
rect 35391 8993 35403 9027
rect 36817 9027 36875 9033
rect 35345 8987 35403 8993
rect 36188 8996 36768 9024
rect 30745 8959 30803 8965
rect 30745 8956 30757 8959
rect 30616 8928 30757 8956
rect 30616 8916 30622 8928
rect 30745 8925 30757 8928
rect 30791 8925 30803 8959
rect 31205 8959 31263 8965
rect 31205 8956 31217 8959
rect 30745 8919 30803 8925
rect 31131 8928 31217 8956
rect 30650 8888 30656 8900
rect 30484 8860 30656 8888
rect 30650 8848 30656 8860
rect 30708 8848 30714 8900
rect 31131 8820 31159 8928
rect 31205 8925 31217 8928
rect 31251 8925 31263 8959
rect 31386 8956 31392 8968
rect 31347 8928 31392 8956
rect 31205 8919 31263 8925
rect 31386 8916 31392 8928
rect 31444 8916 31450 8968
rect 32769 8959 32827 8965
rect 32769 8925 32781 8959
rect 32815 8956 32827 8959
rect 33226 8956 33232 8968
rect 32815 8928 33232 8956
rect 32815 8925 32827 8928
rect 32769 8919 32827 8925
rect 33226 8916 33232 8928
rect 33284 8916 33290 8968
rect 33318 8916 33324 8968
rect 33376 8956 33382 8968
rect 33597 8959 33655 8965
rect 33597 8956 33609 8959
rect 33376 8928 33609 8956
rect 33376 8916 33382 8928
rect 33597 8925 33609 8928
rect 33643 8925 33655 8959
rect 35250 8956 35256 8968
rect 35211 8928 35256 8956
rect 33597 8919 33655 8925
rect 35250 8916 35256 8928
rect 35308 8916 35314 8968
rect 36188 8900 36216 8996
rect 36262 8916 36268 8968
rect 36320 8956 36326 8968
rect 36449 8959 36507 8965
rect 36449 8956 36461 8959
rect 36320 8928 36461 8956
rect 36320 8916 36326 8928
rect 36449 8925 36461 8928
rect 36495 8925 36507 8959
rect 36449 8919 36507 8925
rect 36633 8959 36691 8965
rect 36633 8925 36645 8959
rect 36679 8925 36691 8959
rect 36740 8956 36768 8996
rect 36817 8993 36829 9027
rect 36863 9024 36875 9027
rect 39853 9027 39911 9033
rect 36863 8996 38424 9024
rect 36863 8993 36875 8996
rect 36817 8987 36875 8993
rect 37369 8959 37427 8965
rect 37369 8956 37381 8959
rect 36740 8928 37381 8956
rect 36633 8919 36691 8925
rect 37369 8925 37381 8928
rect 37415 8956 37427 8959
rect 37458 8956 37464 8968
rect 37415 8928 37464 8956
rect 37415 8925 37427 8928
rect 37369 8919 37427 8925
rect 36170 8888 36176 8900
rect 32048 8860 36176 8888
rect 32048 8829 32076 8860
rect 36170 8848 36176 8860
rect 36228 8848 36234 8900
rect 36648 8888 36676 8919
rect 37458 8916 37464 8928
rect 37516 8916 37522 8968
rect 38396 8965 38424 8996
rect 38488 8996 39160 9024
rect 37553 8959 37611 8965
rect 37553 8925 37565 8959
rect 37599 8925 37611 8959
rect 37553 8919 37611 8925
rect 38381 8959 38439 8965
rect 38381 8925 38393 8959
rect 38427 8925 38439 8959
rect 38381 8919 38439 8925
rect 37568 8888 37596 8919
rect 38488 8888 38516 8996
rect 39132 8965 39160 8996
rect 39853 8993 39865 9027
rect 39899 8993 39911 9027
rect 39853 8987 39911 8993
rect 40126 8984 40132 9036
rect 40184 9024 40190 9036
rect 43640 9024 43668 9132
rect 44453 9129 44465 9163
rect 44499 9160 44511 9163
rect 46658 9160 46664 9172
rect 44499 9132 46664 9160
rect 44499 9129 44511 9132
rect 44453 9123 44511 9129
rect 46658 9120 46664 9132
rect 46716 9120 46722 9172
rect 48130 9160 48136 9172
rect 48091 9132 48136 9160
rect 48130 9120 48136 9132
rect 48188 9120 48194 9172
rect 48222 9120 48228 9172
rect 48280 9160 48286 9172
rect 51258 9160 51264 9172
rect 48280 9132 51074 9160
rect 51219 9132 51264 9160
rect 48280 9120 48286 9132
rect 50522 9092 50528 9104
rect 50483 9064 50528 9092
rect 50522 9052 50528 9064
rect 50580 9052 50586 9104
rect 44085 9027 44143 9033
rect 44085 9024 44097 9027
rect 40184 8996 42012 9024
rect 43640 8996 44097 9024
rect 40184 8984 40190 8996
rect 38933 8959 38991 8965
rect 38933 8925 38945 8959
rect 38979 8925 38991 8959
rect 38933 8919 38991 8925
rect 39117 8959 39175 8965
rect 39117 8925 39129 8959
rect 39163 8956 39175 8959
rect 39666 8956 39672 8968
rect 39163 8928 39672 8956
rect 39163 8925 39175 8928
rect 39117 8919 39175 8925
rect 36648 8860 38516 8888
rect 32033 8823 32091 8829
rect 32033 8820 32045 8823
rect 30392 8792 32045 8820
rect 32033 8789 32045 8792
rect 32079 8789 32091 8823
rect 32033 8783 32091 8789
rect 33410 8780 33416 8832
rect 33468 8820 33474 8832
rect 34057 8823 34115 8829
rect 34057 8820 34069 8823
rect 33468 8792 34069 8820
rect 33468 8780 33474 8792
rect 34057 8789 34069 8792
rect 34103 8789 34115 8823
rect 34057 8783 34115 8789
rect 35621 8823 35679 8829
rect 35621 8789 35633 8823
rect 35667 8820 35679 8823
rect 36906 8820 36912 8832
rect 35667 8792 36912 8820
rect 35667 8789 35679 8792
rect 35621 8783 35679 8789
rect 36906 8780 36912 8792
rect 36964 8780 36970 8832
rect 37826 8780 37832 8832
rect 37884 8820 37890 8832
rect 38948 8820 38976 8919
rect 39666 8916 39672 8928
rect 39724 8956 39730 8968
rect 40037 8959 40095 8965
rect 39724 8952 39988 8956
rect 40037 8952 40049 8959
rect 39724 8928 40049 8952
rect 39724 8916 39730 8928
rect 39960 8925 40049 8928
rect 40083 8956 40095 8959
rect 40310 8956 40316 8968
rect 40083 8928 40316 8956
rect 40083 8925 40095 8928
rect 39960 8924 40095 8925
rect 40037 8919 40095 8924
rect 40310 8916 40316 8928
rect 40368 8916 40374 8968
rect 40681 8959 40739 8965
rect 40681 8925 40693 8959
rect 40727 8925 40739 8959
rect 41322 8956 41328 8968
rect 41283 8928 41328 8956
rect 40681 8919 40739 8925
rect 39022 8848 39028 8900
rect 39080 8888 39086 8900
rect 40696 8888 40724 8919
rect 41322 8916 41328 8928
rect 41380 8916 41386 8968
rect 41984 8965 42012 8996
rect 44085 8993 44097 8996
rect 44131 9024 44143 9027
rect 45005 9027 45063 9033
rect 45005 9024 45017 9027
rect 44131 8996 45017 9024
rect 44131 8993 44143 8996
rect 44085 8987 44143 8993
rect 45005 8993 45017 8996
rect 45051 8993 45063 9027
rect 48593 9027 48651 9033
rect 48593 9024 48605 9027
rect 45005 8987 45063 8993
rect 46676 8996 48605 9024
rect 46676 8968 46704 8996
rect 48593 8993 48605 8996
rect 48639 8993 48651 9027
rect 48593 8987 48651 8993
rect 41969 8959 42027 8965
rect 41969 8925 41981 8959
rect 42015 8925 42027 8959
rect 41969 8919 42027 8925
rect 43349 8959 43407 8965
rect 43349 8925 43361 8959
rect 43395 8956 43407 8959
rect 43438 8956 43444 8968
rect 43395 8928 43444 8956
rect 43395 8925 43407 8928
rect 43349 8919 43407 8925
rect 43438 8916 43444 8928
rect 43496 8916 43502 8968
rect 43622 8956 43628 8968
rect 43583 8928 43628 8956
rect 43622 8916 43628 8928
rect 43680 8916 43686 8968
rect 44266 8956 44272 8968
rect 44227 8928 44272 8956
rect 44266 8916 44272 8928
rect 44324 8916 44330 8968
rect 46382 8956 46388 8968
rect 46343 8928 46388 8956
rect 46382 8916 46388 8928
rect 46440 8916 46446 8968
rect 46658 8956 46664 8968
rect 46619 8928 46664 8956
rect 46658 8916 46664 8928
rect 46716 8916 46722 8968
rect 47857 8959 47915 8965
rect 47857 8925 47869 8959
rect 47903 8925 47915 8959
rect 47857 8919 47915 8925
rect 47949 8959 48007 8965
rect 47949 8925 47961 8959
rect 47995 8956 48007 8959
rect 48222 8956 48228 8968
rect 47995 8928 48228 8956
rect 47995 8925 48007 8928
rect 47949 8919 48007 8925
rect 39080 8860 40724 8888
rect 39080 8848 39086 8860
rect 42426 8848 42432 8900
rect 42484 8888 42490 8900
rect 43640 8888 43668 8916
rect 42484 8860 43668 8888
rect 42484 8848 42490 8860
rect 45462 8848 45468 8900
rect 45520 8888 45526 8900
rect 47121 8891 47179 8897
rect 47121 8888 47133 8891
rect 45520 8860 47133 8888
rect 45520 8848 45526 8860
rect 47121 8857 47133 8860
rect 47167 8857 47179 8891
rect 47872 8888 47900 8919
rect 48222 8916 48228 8928
rect 48280 8916 48286 8968
rect 48406 8888 48412 8900
rect 47872 8860 48412 8888
rect 47121 8851 47179 8857
rect 48406 8848 48412 8860
rect 48464 8848 48470 8900
rect 48608 8888 48636 8987
rect 48866 8956 48872 8968
rect 48827 8928 48872 8956
rect 48866 8916 48872 8928
rect 48924 8916 48930 8968
rect 51046 8956 51074 9132
rect 51258 9120 51264 9132
rect 51316 9120 51322 9172
rect 52270 8984 52276 9036
rect 52328 9024 52334 9036
rect 52365 9027 52423 9033
rect 52365 9024 52377 9027
rect 52328 8996 52377 9024
rect 52328 8984 52334 8996
rect 52365 8993 52377 8996
rect 52411 8993 52423 9027
rect 52365 8987 52423 8993
rect 51445 8959 51503 8965
rect 51445 8956 51457 8959
rect 50540 8928 50844 8956
rect 51046 8928 51457 8956
rect 50338 8888 50344 8900
rect 48608 8860 50344 8888
rect 50338 8848 50344 8860
rect 50396 8848 50402 8900
rect 37884 8792 38976 8820
rect 39301 8823 39359 8829
rect 37884 8780 37890 8792
rect 39301 8789 39313 8823
rect 39347 8820 39359 8823
rect 40126 8820 40132 8832
rect 39347 8792 40132 8820
rect 39347 8789 39359 8792
rect 39301 8783 39359 8789
rect 40126 8780 40132 8792
rect 40184 8780 40190 8832
rect 40221 8823 40279 8829
rect 40221 8789 40233 8823
rect 40267 8820 40279 8823
rect 40310 8820 40316 8832
rect 40267 8792 40316 8820
rect 40267 8789 40279 8792
rect 40221 8783 40279 8789
rect 40310 8780 40316 8792
rect 40368 8780 40374 8832
rect 40865 8823 40923 8829
rect 40865 8789 40877 8823
rect 40911 8820 40923 8823
rect 41138 8820 41144 8832
rect 40911 8792 41144 8820
rect 40911 8789 40923 8792
rect 40865 8783 40923 8789
rect 41138 8780 41144 8792
rect 41196 8780 41202 8832
rect 41509 8823 41567 8829
rect 41509 8789 41521 8823
rect 41555 8820 41567 8823
rect 41690 8820 41696 8832
rect 41555 8792 41696 8820
rect 41555 8789 41567 8792
rect 41509 8783 41567 8789
rect 41690 8780 41696 8792
rect 41748 8780 41754 8832
rect 41874 8780 41880 8832
rect 41932 8820 41938 8832
rect 45649 8823 45707 8829
rect 45649 8820 45661 8823
rect 41932 8792 45661 8820
rect 41932 8780 41938 8792
rect 45649 8789 45661 8792
rect 45695 8820 45707 8823
rect 46290 8820 46296 8832
rect 45695 8792 46296 8820
rect 45695 8789 45707 8792
rect 45649 8783 45707 8789
rect 46290 8780 46296 8792
rect 46348 8820 46354 8832
rect 49605 8823 49663 8829
rect 49605 8820 49617 8823
rect 46348 8792 49617 8820
rect 46348 8780 46354 8792
rect 49605 8789 49617 8792
rect 49651 8820 49663 8823
rect 50540 8820 50568 8928
rect 50706 8888 50712 8900
rect 50667 8860 50712 8888
rect 50706 8848 50712 8860
rect 50764 8848 50770 8900
rect 49651 8792 50568 8820
rect 50816 8820 50844 8928
rect 51445 8925 51457 8928
rect 51491 8956 51503 8959
rect 51534 8956 51540 8968
rect 51491 8928 51540 8956
rect 51491 8925 51503 8928
rect 51445 8919 51503 8925
rect 51534 8916 51540 8928
rect 51592 8916 51598 8968
rect 51629 8959 51687 8965
rect 51629 8925 51641 8959
rect 51675 8956 51687 8959
rect 52086 8956 52092 8968
rect 51675 8928 52092 8956
rect 51675 8925 51687 8928
rect 51629 8919 51687 8925
rect 52086 8916 52092 8928
rect 52144 8916 52150 8968
rect 52641 8959 52699 8965
rect 52641 8925 52653 8959
rect 52687 8925 52699 8959
rect 52641 8919 52699 8925
rect 52656 8888 52684 8919
rect 53374 8916 53380 8968
rect 53432 8956 53438 8968
rect 53469 8959 53527 8965
rect 53469 8956 53481 8959
rect 53432 8928 53481 8956
rect 53432 8916 53438 8928
rect 53469 8925 53481 8928
rect 53515 8925 53527 8959
rect 54110 8956 54116 8968
rect 54071 8928 54116 8956
rect 53469 8919 53527 8925
rect 54110 8916 54116 8928
rect 54168 8916 54174 8968
rect 52656 8860 53972 8888
rect 51166 8820 51172 8832
rect 50816 8792 51172 8820
rect 49651 8789 49663 8792
rect 49605 8783 49663 8789
rect 51166 8780 51172 8792
rect 51224 8780 51230 8832
rect 53944 8829 53972 8860
rect 53929 8823 53987 8829
rect 53929 8789 53941 8823
rect 53975 8789 53987 8823
rect 53929 8783 53987 8789
rect 1104 8730 58880 8752
rect 1104 8678 15398 8730
rect 15450 8678 15462 8730
rect 15514 8678 15526 8730
rect 15578 8678 15590 8730
rect 15642 8678 15654 8730
rect 15706 8678 29846 8730
rect 29898 8678 29910 8730
rect 29962 8678 29974 8730
rect 30026 8678 30038 8730
rect 30090 8678 30102 8730
rect 30154 8678 44294 8730
rect 44346 8678 44358 8730
rect 44410 8678 44422 8730
rect 44474 8678 44486 8730
rect 44538 8678 44550 8730
rect 44602 8678 58880 8730
rect 1104 8656 58880 8678
rect 4706 8616 4712 8628
rect 4667 8588 4712 8616
rect 4706 8576 4712 8588
rect 4764 8576 4770 8628
rect 6454 8576 6460 8628
rect 6512 8616 6518 8628
rect 7837 8619 7895 8625
rect 7837 8616 7849 8619
rect 6512 8588 7849 8616
rect 6512 8576 6518 8588
rect 7837 8585 7849 8588
rect 7883 8585 7895 8619
rect 7837 8579 7895 8585
rect 7926 8576 7932 8628
rect 7984 8616 7990 8628
rect 7984 8588 9260 8616
rect 7984 8576 7990 8588
rect 2314 8548 2320 8560
rect 1596 8520 2320 8548
rect 1596 8489 1624 8520
rect 2314 8508 2320 8520
rect 2372 8548 2378 8560
rect 2590 8548 2596 8560
rect 2372 8520 2596 8548
rect 2372 8508 2378 8520
rect 2590 8508 2596 8520
rect 2648 8508 2654 8560
rect 4982 8508 4988 8560
rect 5040 8548 5046 8560
rect 9033 8551 9091 8557
rect 9033 8548 9045 8551
rect 5040 8520 9045 8548
rect 5040 8508 5046 8520
rect 9033 8517 9045 8520
rect 9079 8517 9091 8551
rect 9232 8548 9260 8588
rect 10778 8576 10784 8628
rect 10836 8616 10842 8628
rect 10873 8619 10931 8625
rect 10873 8616 10885 8619
rect 10836 8588 10885 8616
rect 10836 8576 10842 8588
rect 10873 8585 10885 8588
rect 10919 8585 10931 8619
rect 10873 8579 10931 8585
rect 11330 8576 11336 8628
rect 11388 8616 11394 8628
rect 12437 8619 12495 8625
rect 12437 8616 12449 8619
rect 11388 8588 12449 8616
rect 11388 8576 11394 8588
rect 12437 8585 12449 8588
rect 12483 8585 12495 8619
rect 12437 8579 12495 8585
rect 13357 8619 13415 8625
rect 13357 8585 13369 8619
rect 13403 8616 13415 8619
rect 13538 8616 13544 8628
rect 13403 8588 13544 8616
rect 13403 8585 13415 8588
rect 13357 8579 13415 8585
rect 13538 8576 13544 8588
rect 13596 8576 13602 8628
rect 14001 8619 14059 8625
rect 14001 8585 14013 8619
rect 14047 8616 14059 8619
rect 14458 8616 14464 8628
rect 14047 8588 14464 8616
rect 14047 8585 14059 8588
rect 14001 8579 14059 8585
rect 14458 8576 14464 8588
rect 14516 8576 14522 8628
rect 14645 8619 14703 8625
rect 14645 8585 14657 8619
rect 14691 8616 14703 8619
rect 17402 8616 17408 8628
rect 14691 8588 17408 8616
rect 14691 8585 14703 8588
rect 14645 8579 14703 8585
rect 17402 8576 17408 8588
rect 17460 8576 17466 8628
rect 18785 8619 18843 8625
rect 18785 8585 18797 8619
rect 18831 8616 18843 8619
rect 21085 8619 21143 8625
rect 18831 8588 20484 8616
rect 18831 8585 18843 8588
rect 18785 8579 18843 8585
rect 9232 8520 9352 8548
rect 9033 8511 9091 8517
rect 1581 8483 1639 8489
rect 1581 8449 1593 8483
rect 1627 8449 1639 8483
rect 1581 8443 1639 8449
rect 1765 8483 1823 8489
rect 1765 8449 1777 8483
rect 1811 8480 1823 8483
rect 2038 8480 2044 8492
rect 1811 8452 2044 8480
rect 1811 8449 1823 8452
rect 1765 8443 1823 8449
rect 2038 8440 2044 8452
rect 2096 8440 2102 8492
rect 2409 8483 2467 8489
rect 2409 8449 2421 8483
rect 2455 8480 2467 8483
rect 3510 8480 3516 8492
rect 2455 8452 3516 8480
rect 2455 8449 2467 8452
rect 2409 8443 2467 8449
rect 3510 8440 3516 8452
rect 3568 8440 3574 8492
rect 3697 8483 3755 8489
rect 3697 8449 3709 8483
rect 3743 8480 3755 8483
rect 4338 8480 4344 8492
rect 3743 8452 4344 8480
rect 3743 8449 3755 8452
rect 3697 8443 3755 8449
rect 4338 8440 4344 8452
rect 4396 8440 4402 8492
rect 4522 8480 4528 8492
rect 4483 8452 4528 8480
rect 4522 8440 4528 8452
rect 4580 8440 4586 8492
rect 5810 8480 5816 8492
rect 5771 8452 5816 8480
rect 5810 8440 5816 8452
rect 5868 8440 5874 8492
rect 6641 8483 6699 8489
rect 6641 8480 6653 8483
rect 5920 8452 6653 8480
rect 2593 8415 2651 8421
rect 2593 8381 2605 8415
rect 2639 8412 2651 8415
rect 2774 8412 2780 8424
rect 2639 8384 2780 8412
rect 2639 8381 2651 8384
rect 2593 8375 2651 8381
rect 2774 8372 2780 8384
rect 2832 8412 2838 8424
rect 3418 8412 3424 8424
rect 2832 8384 3424 8412
rect 2832 8372 2838 8384
rect 3418 8372 3424 8384
rect 3476 8372 3482 8424
rect 4356 8412 4384 8440
rect 5442 8412 5448 8424
rect 4356 8384 5448 8412
rect 5442 8372 5448 8384
rect 5500 8372 5506 8424
rect 1394 8304 1400 8356
rect 1452 8344 1458 8356
rect 1673 8347 1731 8353
rect 1673 8344 1685 8347
rect 1452 8316 1685 8344
rect 1452 8304 1458 8316
rect 1673 8313 1685 8316
rect 1719 8313 1731 8347
rect 1673 8307 1731 8313
rect 1854 8304 1860 8356
rect 1912 8344 1918 8356
rect 3329 8347 3387 8353
rect 3329 8344 3341 8347
rect 1912 8316 3341 8344
rect 1912 8304 1918 8316
rect 3329 8313 3341 8316
rect 3375 8313 3387 8347
rect 3329 8307 3387 8313
rect 4246 8304 4252 8356
rect 4304 8344 4310 8356
rect 5920 8344 5948 8452
rect 6641 8449 6653 8452
rect 6687 8449 6699 8483
rect 6641 8443 6699 8449
rect 8021 8483 8079 8489
rect 8021 8449 8033 8483
rect 8067 8449 8079 8483
rect 8202 8480 8208 8492
rect 8163 8452 8208 8480
rect 8021 8443 8079 8449
rect 6365 8415 6423 8421
rect 6365 8381 6377 8415
rect 6411 8381 6423 8415
rect 6365 8375 6423 8381
rect 4304 8316 5948 8344
rect 4304 8304 4310 8316
rect 1578 8236 1584 8288
rect 1636 8276 1642 8288
rect 2225 8279 2283 8285
rect 2225 8276 2237 8279
rect 1636 8248 2237 8276
rect 1636 8236 1642 8248
rect 2225 8245 2237 8248
rect 2271 8245 2283 8279
rect 2225 8239 2283 8245
rect 5629 8279 5687 8285
rect 5629 8245 5641 8279
rect 5675 8276 5687 8279
rect 5718 8276 5724 8288
rect 5675 8248 5724 8276
rect 5675 8245 5687 8248
rect 5629 8239 5687 8245
rect 5718 8236 5724 8248
rect 5776 8236 5782 8288
rect 5810 8236 5816 8288
rect 5868 8276 5874 8288
rect 6380 8276 6408 8375
rect 8037 8344 8065 8443
rect 8202 8440 8208 8452
rect 8260 8440 8266 8492
rect 9324 8489 9352 8520
rect 9490 8508 9496 8560
rect 9548 8548 9554 8560
rect 11517 8551 11575 8557
rect 11517 8548 11529 8551
rect 9548 8520 11529 8548
rect 9548 8508 9554 8520
rect 11517 8517 11529 8520
rect 11563 8517 11575 8551
rect 14918 8548 14924 8560
rect 11517 8511 11575 8517
rect 11624 8520 12434 8548
rect 9217 8483 9275 8489
rect 9217 8449 9229 8483
rect 9263 8449 9275 8483
rect 9217 8443 9275 8449
rect 9309 8483 9367 8489
rect 9309 8449 9321 8483
rect 9355 8449 9367 8483
rect 9309 8443 9367 8449
rect 10137 8483 10195 8489
rect 10137 8449 10149 8483
rect 10183 8449 10195 8483
rect 10318 8480 10324 8492
rect 10279 8452 10324 8480
rect 10137 8443 10195 8449
rect 9232 8412 9260 8443
rect 6932 8316 8065 8344
rect 8128 8384 9260 8412
rect 10152 8412 10180 8443
rect 10318 8440 10324 8452
rect 10376 8440 10382 8492
rect 10410 8440 10416 8492
rect 10468 8480 10474 8492
rect 10781 8483 10839 8489
rect 10781 8480 10793 8483
rect 10468 8452 10793 8480
rect 10468 8440 10474 8452
rect 10781 8449 10793 8452
rect 10827 8449 10839 8483
rect 10781 8443 10839 8449
rect 10965 8483 11023 8489
rect 10965 8449 10977 8483
rect 11011 8480 11023 8483
rect 11146 8480 11152 8492
rect 11011 8452 11152 8480
rect 11011 8449 11023 8452
rect 10965 8443 11023 8449
rect 10428 8412 10456 8440
rect 10152 8384 10456 8412
rect 6932 8276 6960 8316
rect 7374 8276 7380 8288
rect 5868 8248 6960 8276
rect 7335 8248 7380 8276
rect 5868 8236 5874 8248
rect 7374 8236 7380 8248
rect 7432 8236 7438 8288
rect 7742 8236 7748 8288
rect 7800 8276 7806 8288
rect 8128 8276 8156 8384
rect 8386 8304 8392 8356
rect 8444 8344 8450 8356
rect 10321 8347 10379 8353
rect 10321 8344 10333 8347
rect 8444 8316 10333 8344
rect 8444 8304 8450 8316
rect 10321 8313 10333 8316
rect 10367 8344 10379 8347
rect 10796 8344 10824 8443
rect 11146 8440 11152 8452
rect 11204 8440 11210 8492
rect 11238 8440 11244 8492
rect 11296 8480 11302 8492
rect 11624 8480 11652 8520
rect 11296 8452 11652 8480
rect 11701 8483 11759 8489
rect 11296 8440 11302 8452
rect 11701 8449 11713 8483
rect 11747 8449 11759 8483
rect 11701 8443 11759 8449
rect 10870 8372 10876 8424
rect 10928 8412 10934 8424
rect 11716 8412 11744 8443
rect 11790 8440 11796 8492
rect 11848 8480 11854 8492
rect 12406 8480 12434 8520
rect 14568 8520 14924 8548
rect 12621 8483 12679 8489
rect 12621 8480 12633 8483
rect 11848 8452 11893 8480
rect 12406 8452 12633 8480
rect 11848 8440 11854 8452
rect 12621 8449 12633 8452
rect 12667 8449 12679 8483
rect 12621 8443 12679 8449
rect 13817 8483 13875 8489
rect 13817 8449 13829 8483
rect 13863 8449 13875 8483
rect 13817 8443 13875 8449
rect 14461 8483 14519 8489
rect 14461 8449 14473 8483
rect 14507 8480 14519 8483
rect 14568 8480 14596 8520
rect 14918 8508 14924 8520
rect 14976 8508 14982 8560
rect 16666 8508 16672 8560
rect 16724 8548 16730 8560
rect 17218 8548 17224 8560
rect 16724 8520 17224 8548
rect 16724 8508 16730 8520
rect 17218 8508 17224 8520
rect 17276 8548 17282 8560
rect 20254 8548 20260 8560
rect 17276 8520 20260 8548
rect 17276 8508 17282 8520
rect 20254 8508 20260 8520
rect 20312 8508 20318 8560
rect 14507 8452 14596 8480
rect 14507 8449 14519 8452
rect 14461 8443 14519 8449
rect 10928 8384 11744 8412
rect 12805 8415 12863 8421
rect 10928 8372 10934 8384
rect 12805 8381 12817 8415
rect 12851 8381 12863 8415
rect 12805 8375 12863 8381
rect 10962 8344 10968 8356
rect 10367 8316 10732 8344
rect 10796 8316 10968 8344
rect 10367 8313 10379 8316
rect 10321 8307 10379 8313
rect 7800 8248 8156 8276
rect 10704 8276 10732 8316
rect 10962 8304 10968 8316
rect 11020 8304 11026 8356
rect 11238 8276 11244 8288
rect 10704 8248 11244 8276
rect 7800 8236 7806 8248
rect 11238 8236 11244 8248
rect 11296 8236 11302 8288
rect 11790 8236 11796 8288
rect 11848 8276 11854 8288
rect 12434 8276 12440 8288
rect 11848 8248 12440 8276
rect 11848 8236 11854 8248
rect 12434 8236 12440 8248
rect 12492 8276 12498 8288
rect 12820 8276 12848 8375
rect 13832 8344 13860 8443
rect 14642 8440 14648 8492
rect 14700 8480 14706 8492
rect 15102 8480 15108 8492
rect 14700 8452 15108 8480
rect 14700 8440 14706 8452
rect 15102 8440 15108 8452
rect 15160 8440 15166 8492
rect 15194 8440 15200 8492
rect 15252 8480 15258 8492
rect 15289 8483 15347 8489
rect 15289 8480 15301 8483
rect 15252 8452 15301 8480
rect 15252 8440 15258 8452
rect 15289 8449 15301 8452
rect 15335 8449 15347 8483
rect 15289 8443 15347 8449
rect 15933 8483 15991 8489
rect 15933 8449 15945 8483
rect 15979 8480 15991 8483
rect 16390 8480 16396 8492
rect 15979 8452 16396 8480
rect 15979 8449 15991 8452
rect 15933 8443 15991 8449
rect 16390 8440 16396 8452
rect 16448 8440 16454 8492
rect 13998 8372 14004 8424
rect 14056 8412 14062 8424
rect 15749 8415 15807 8421
rect 15749 8412 15761 8415
rect 14056 8384 15761 8412
rect 14056 8372 14062 8384
rect 15749 8381 15761 8384
rect 15795 8381 15807 8415
rect 15749 8375 15807 8381
rect 16117 8415 16175 8421
rect 16117 8381 16129 8415
rect 16163 8412 16175 8415
rect 16684 8412 16712 8508
rect 17034 8480 17040 8492
rect 16947 8452 17040 8480
rect 17034 8440 17040 8452
rect 17092 8480 17098 8492
rect 17865 8483 17923 8489
rect 17865 8480 17877 8483
rect 17092 8452 17877 8480
rect 17092 8440 17098 8452
rect 17865 8449 17877 8452
rect 17911 8449 17923 8483
rect 17865 8443 17923 8449
rect 18601 8483 18659 8489
rect 18601 8449 18613 8483
rect 18647 8449 18659 8483
rect 19426 8480 19432 8492
rect 19387 8452 19432 8480
rect 18601 8443 18659 8449
rect 16163 8384 16712 8412
rect 16163 8381 16175 8384
rect 16117 8375 16175 8381
rect 16942 8372 16948 8424
rect 17000 8412 17006 8424
rect 17221 8415 17279 8421
rect 17221 8412 17233 8415
rect 17000 8384 17233 8412
rect 17000 8372 17006 8384
rect 17221 8381 17233 8384
rect 17267 8412 17279 8415
rect 17770 8412 17776 8424
rect 17267 8384 17776 8412
rect 17267 8381 17279 8384
rect 17221 8375 17279 8381
rect 17770 8372 17776 8384
rect 17828 8372 17834 8424
rect 16853 8347 16911 8353
rect 16853 8344 16865 8347
rect 13832 8316 16865 8344
rect 16853 8313 16865 8316
rect 16899 8313 16911 8347
rect 17880 8344 17908 8443
rect 18049 8415 18107 8421
rect 18049 8381 18061 8415
rect 18095 8412 18107 8415
rect 18230 8412 18236 8424
rect 18095 8384 18236 8412
rect 18095 8381 18107 8384
rect 18049 8375 18107 8381
rect 18230 8372 18236 8384
rect 18288 8372 18294 8424
rect 18616 8412 18644 8443
rect 19426 8440 19432 8452
rect 19484 8440 19490 8492
rect 19613 8483 19671 8489
rect 19613 8449 19625 8483
rect 19659 8480 19671 8483
rect 19886 8480 19892 8492
rect 19659 8452 19892 8480
rect 19659 8449 19671 8452
rect 19613 8443 19671 8449
rect 19886 8440 19892 8452
rect 19944 8440 19950 8492
rect 20349 8483 20407 8489
rect 20349 8449 20361 8483
rect 20395 8480 20407 8483
rect 20456 8480 20484 8588
rect 21085 8585 21097 8619
rect 21131 8616 21143 8619
rect 21266 8616 21272 8628
rect 21131 8588 21272 8616
rect 21131 8585 21143 8588
rect 21085 8579 21143 8585
rect 21266 8576 21272 8588
rect 21324 8576 21330 8628
rect 21634 8576 21640 8628
rect 21692 8616 21698 8628
rect 22833 8619 22891 8625
rect 22833 8616 22845 8619
rect 21692 8588 22845 8616
rect 21692 8576 21698 8588
rect 22833 8585 22845 8588
rect 22879 8585 22891 8619
rect 22833 8579 22891 8585
rect 23290 8576 23296 8628
rect 23348 8616 23354 8628
rect 24949 8619 25007 8625
rect 24949 8616 24961 8619
rect 23348 8588 24961 8616
rect 23348 8576 23354 8588
rect 24949 8585 24961 8588
rect 24995 8585 25007 8619
rect 24949 8579 25007 8585
rect 25222 8576 25228 8628
rect 25280 8616 25286 8628
rect 26142 8616 26148 8628
rect 25280 8588 26148 8616
rect 25280 8576 25286 8588
rect 26142 8576 26148 8588
rect 26200 8576 26206 8628
rect 27062 8616 27068 8628
rect 27023 8588 27068 8616
rect 27062 8576 27068 8588
rect 27120 8576 27126 8628
rect 28537 8619 28595 8625
rect 28537 8585 28549 8619
rect 28583 8616 28595 8619
rect 28994 8616 29000 8628
rect 28583 8588 29000 8616
rect 28583 8585 28595 8588
rect 28537 8579 28595 8585
rect 28994 8576 29000 8588
rect 29052 8576 29058 8628
rect 31478 8616 31484 8628
rect 30208 8588 31340 8616
rect 31439 8588 31484 8616
rect 22094 8508 22100 8560
rect 22152 8548 22158 8560
rect 30208 8548 30236 8588
rect 22152 8520 30236 8548
rect 31312 8548 31340 8588
rect 31478 8576 31484 8588
rect 31536 8576 31542 8628
rect 33226 8616 33232 8628
rect 33187 8588 33232 8616
rect 33226 8576 33232 8588
rect 33284 8576 33290 8628
rect 33318 8576 33324 8628
rect 33376 8616 33382 8628
rect 34885 8619 34943 8625
rect 34885 8616 34897 8619
rect 33376 8588 34897 8616
rect 33376 8576 33382 8588
rect 34885 8585 34897 8588
rect 34931 8616 34943 8619
rect 35066 8616 35072 8628
rect 34931 8588 35072 8616
rect 34931 8585 34943 8588
rect 34885 8579 34943 8585
rect 35066 8576 35072 8588
rect 35124 8576 35130 8628
rect 39022 8616 39028 8628
rect 38983 8588 39028 8616
rect 39022 8576 39028 8588
rect 39080 8576 39086 8628
rect 39666 8616 39672 8628
rect 39627 8588 39672 8616
rect 39666 8576 39672 8588
rect 39724 8576 39730 8628
rect 39942 8576 39948 8628
rect 40000 8616 40006 8628
rect 40129 8619 40187 8625
rect 40129 8616 40141 8619
rect 40000 8588 40141 8616
rect 40000 8576 40006 8588
rect 40129 8585 40141 8588
rect 40175 8585 40187 8619
rect 40129 8579 40187 8585
rect 40770 8576 40776 8628
rect 40828 8616 40834 8628
rect 43438 8616 43444 8628
rect 40828 8588 43300 8616
rect 43399 8588 43444 8616
rect 40828 8576 40834 8588
rect 31312 8520 35204 8548
rect 22152 8508 22158 8520
rect 20395 8452 20484 8480
rect 21928 8452 22232 8480
rect 20395 8449 20407 8452
rect 20349 8443 20407 8449
rect 19702 8412 19708 8424
rect 18616 8384 19708 8412
rect 19702 8372 19708 8384
rect 19760 8372 19766 8424
rect 20070 8412 20076 8424
rect 20031 8384 20076 8412
rect 20070 8372 20076 8384
rect 20128 8372 20134 8424
rect 21928 8356 21956 8452
rect 22204 8412 22232 8452
rect 22278 8440 22284 8492
rect 22336 8480 22342 8492
rect 23017 8483 23075 8489
rect 22336 8452 22381 8480
rect 22336 8440 22342 8452
rect 23017 8449 23029 8483
rect 23063 8449 23075 8483
rect 23658 8480 23664 8492
rect 23619 8452 23664 8480
rect 23017 8443 23075 8449
rect 23032 8412 23060 8443
rect 23658 8440 23664 8452
rect 23716 8440 23722 8492
rect 24210 8440 24216 8492
rect 24268 8480 24274 8492
rect 24305 8483 24363 8489
rect 24305 8480 24317 8483
rect 24268 8452 24317 8480
rect 24268 8440 24274 8452
rect 24305 8449 24317 8452
rect 24351 8449 24363 8483
rect 24305 8443 24363 8449
rect 24394 8440 24400 8492
rect 24452 8480 24458 8492
rect 24489 8483 24547 8489
rect 24489 8480 24501 8483
rect 24452 8452 24501 8480
rect 24452 8440 24458 8452
rect 24489 8449 24501 8452
rect 24535 8480 24547 8483
rect 24670 8480 24676 8492
rect 24535 8452 24676 8480
rect 24535 8449 24547 8452
rect 24489 8443 24547 8449
rect 24670 8440 24676 8452
rect 24728 8440 24734 8492
rect 25685 8483 25743 8489
rect 25685 8480 25697 8483
rect 24780 8452 25697 8480
rect 22204 8384 23060 8412
rect 23201 8415 23259 8421
rect 23201 8381 23213 8415
rect 23247 8412 23259 8415
rect 23290 8412 23296 8424
rect 23247 8384 23296 8412
rect 23247 8381 23259 8384
rect 23201 8375 23259 8381
rect 23290 8372 23296 8384
rect 23348 8372 23354 8424
rect 24780 8412 24808 8452
rect 25685 8449 25697 8452
rect 25731 8449 25743 8483
rect 25958 8480 25964 8492
rect 25919 8452 25964 8480
rect 25685 8443 25743 8449
rect 25958 8440 25964 8452
rect 26016 8440 26022 8492
rect 26142 8440 26148 8492
rect 26200 8480 26206 8492
rect 27249 8483 27307 8489
rect 27249 8480 27261 8483
rect 26200 8452 27261 8480
rect 26200 8440 26206 8452
rect 27249 8449 27261 8452
rect 27295 8449 27307 8483
rect 27249 8443 27307 8449
rect 27338 8440 27344 8492
rect 27396 8480 27402 8492
rect 28350 8480 28356 8492
rect 27396 8452 27441 8480
rect 27632 8452 28356 8480
rect 27396 8440 27402 8452
rect 23860 8384 24808 8412
rect 21910 8344 21916 8356
rect 17880 8316 20208 8344
rect 16853 8307 16911 8313
rect 12492 8248 12848 8276
rect 12492 8236 12498 8248
rect 14090 8236 14096 8288
rect 14148 8276 14154 8288
rect 15289 8279 15347 8285
rect 15289 8276 15301 8279
rect 14148 8248 15301 8276
rect 14148 8236 14154 8248
rect 15289 8245 15301 8248
rect 15335 8245 15347 8279
rect 17678 8276 17684 8288
rect 17639 8248 17684 8276
rect 15289 8239 15347 8245
rect 17678 8236 17684 8248
rect 17736 8236 17742 8288
rect 19242 8276 19248 8288
rect 19203 8248 19248 8276
rect 19242 8236 19248 8248
rect 19300 8236 19306 8288
rect 20180 8276 20208 8316
rect 21192 8316 21916 8344
rect 20438 8276 20444 8288
rect 20180 8248 20444 8276
rect 20438 8236 20444 8248
rect 20496 8276 20502 8288
rect 21192 8276 21220 8316
rect 21910 8304 21916 8316
rect 21968 8304 21974 8356
rect 22002 8304 22008 8356
rect 22060 8344 22066 8356
rect 23860 8353 23888 8384
rect 22097 8347 22155 8353
rect 22097 8344 22109 8347
rect 22060 8316 22109 8344
rect 22060 8304 22066 8316
rect 22097 8313 22109 8316
rect 22143 8313 22155 8347
rect 22097 8307 22155 8313
rect 23845 8347 23903 8353
rect 23845 8313 23857 8347
rect 23891 8313 23903 8347
rect 23845 8307 23903 8313
rect 24489 8347 24547 8353
rect 24489 8313 24501 8347
rect 24535 8344 24547 8347
rect 25222 8344 25228 8356
rect 24535 8316 25228 8344
rect 24535 8313 24547 8316
rect 24489 8307 24547 8313
rect 25222 8304 25228 8316
rect 25280 8304 25286 8356
rect 20496 8248 21220 8276
rect 20496 8236 20502 8248
rect 21266 8236 21272 8288
rect 21324 8276 21330 8288
rect 24578 8276 24584 8288
rect 21324 8248 24584 8276
rect 21324 8236 21330 8248
rect 24578 8236 24584 8248
rect 24636 8236 24642 8288
rect 24670 8236 24676 8288
rect 24728 8276 24734 8288
rect 27632 8276 27660 8452
rect 28350 8440 28356 8452
rect 28408 8440 28414 8492
rect 28537 8483 28595 8489
rect 28537 8449 28549 8483
rect 28583 8449 28595 8483
rect 28537 8443 28595 8449
rect 28442 8304 28448 8356
rect 28500 8344 28506 8356
rect 28552 8344 28580 8443
rect 28626 8440 28632 8492
rect 28684 8480 28690 8492
rect 29089 8483 29147 8489
rect 29089 8480 29101 8483
rect 28684 8452 29101 8480
rect 28684 8440 28690 8452
rect 29089 8449 29101 8452
rect 29135 8449 29147 8483
rect 30193 8483 30251 8489
rect 29089 8443 29147 8449
rect 29196 8452 30144 8480
rect 29196 8344 29224 8452
rect 29730 8372 29736 8424
rect 29788 8412 29794 8424
rect 30009 8415 30067 8421
rect 30009 8412 30021 8415
rect 29788 8384 30021 8412
rect 29788 8372 29794 8384
rect 30009 8381 30021 8384
rect 30055 8381 30067 8415
rect 30116 8412 30144 8452
rect 30193 8449 30205 8483
rect 30239 8480 30251 8483
rect 30282 8480 30288 8492
rect 30239 8452 30288 8480
rect 30239 8449 30251 8452
rect 30193 8443 30251 8449
rect 30282 8440 30288 8452
rect 30340 8440 30346 8492
rect 30834 8480 30840 8492
rect 30392 8452 30840 8480
rect 30392 8412 30420 8452
rect 30834 8440 30840 8452
rect 30892 8440 30898 8492
rect 31018 8480 31024 8492
rect 30979 8452 31024 8480
rect 31018 8440 31024 8452
rect 31076 8440 31082 8492
rect 31202 8440 31208 8492
rect 31260 8480 31266 8492
rect 32125 8483 32183 8489
rect 32125 8480 32137 8483
rect 31260 8452 32137 8480
rect 31260 8440 31266 8452
rect 32125 8449 32137 8452
rect 32171 8480 32183 8483
rect 33042 8480 33048 8492
rect 32171 8452 33048 8480
rect 32171 8449 32183 8452
rect 32125 8443 32183 8449
rect 33042 8440 33048 8452
rect 33100 8440 33106 8492
rect 34348 8489 34376 8520
rect 33413 8483 33471 8489
rect 33413 8449 33425 8483
rect 33459 8480 33471 8483
rect 34241 8483 34299 8489
rect 34241 8480 34253 8483
rect 33459 8452 34253 8480
rect 33459 8449 33471 8452
rect 33413 8443 33471 8449
rect 34241 8449 34253 8452
rect 34287 8449 34299 8483
rect 34241 8443 34299 8449
rect 34333 8483 34391 8489
rect 34333 8449 34345 8483
rect 34379 8449 34391 8483
rect 35066 8480 35072 8492
rect 35027 8452 35072 8480
rect 34333 8443 34391 8449
rect 32858 8412 32864 8424
rect 30116 8384 30420 8412
rect 30484 8384 32864 8412
rect 30009 8375 30067 8381
rect 28500 8316 28580 8344
rect 28644 8316 29224 8344
rect 29549 8347 29607 8353
rect 28500 8304 28506 8316
rect 24728 8248 27660 8276
rect 24728 8236 24734 8248
rect 27798 8236 27804 8288
rect 27856 8276 27862 8288
rect 28166 8276 28172 8288
rect 27856 8248 28172 8276
rect 27856 8236 27862 8248
rect 28166 8236 28172 8248
rect 28224 8276 28230 8288
rect 28644 8276 28672 8316
rect 29549 8313 29561 8347
rect 29595 8344 29607 8347
rect 30282 8344 30288 8356
rect 29595 8316 30288 8344
rect 29595 8313 29607 8316
rect 29549 8307 29607 8313
rect 30282 8304 30288 8316
rect 30340 8304 30346 8356
rect 29178 8276 29184 8288
rect 28224 8248 28672 8276
rect 29139 8248 29184 8276
rect 28224 8236 28230 8248
rect 29178 8236 29184 8248
rect 29236 8236 29242 8288
rect 30377 8279 30435 8285
rect 30377 8245 30389 8279
rect 30423 8276 30435 8279
rect 30484 8276 30512 8384
rect 32858 8372 32864 8384
rect 32916 8372 32922 8424
rect 30558 8304 30564 8356
rect 30616 8344 30622 8356
rect 31021 8347 31079 8353
rect 31021 8344 31033 8347
rect 30616 8316 31033 8344
rect 30616 8304 30622 8316
rect 31021 8313 31033 8316
rect 31067 8344 31079 8347
rect 31202 8344 31208 8356
rect 31067 8316 31208 8344
rect 31067 8313 31079 8316
rect 31021 8307 31079 8313
rect 31202 8304 31208 8316
rect 31260 8304 31266 8356
rect 31386 8304 31392 8356
rect 31444 8344 31450 8356
rect 32309 8347 32367 8353
rect 32309 8344 32321 8347
rect 31444 8316 32321 8344
rect 31444 8304 31450 8316
rect 32309 8313 32321 8316
rect 32355 8344 32367 8347
rect 33428 8344 33456 8443
rect 35066 8440 35072 8452
rect 35124 8440 35130 8492
rect 35176 8480 35204 8520
rect 35250 8508 35256 8560
rect 35308 8548 35314 8560
rect 43272 8548 43300 8588
rect 43438 8576 43444 8588
rect 43496 8576 43502 8628
rect 43622 8576 43628 8628
rect 43680 8616 43686 8628
rect 43901 8619 43959 8625
rect 43901 8616 43913 8619
rect 43680 8588 43913 8616
rect 43680 8576 43686 8588
rect 43901 8585 43913 8588
rect 43947 8585 43959 8619
rect 43901 8579 43959 8585
rect 44913 8619 44971 8625
rect 44913 8585 44925 8619
rect 44959 8616 44971 8619
rect 46658 8616 46664 8628
rect 44959 8588 46664 8616
rect 44959 8585 44971 8588
rect 44913 8579 44971 8585
rect 46658 8576 46664 8588
rect 46716 8576 46722 8628
rect 49053 8619 49111 8625
rect 49053 8585 49065 8619
rect 49099 8616 49111 8619
rect 49234 8616 49240 8628
rect 49099 8588 49240 8616
rect 49099 8585 49111 8588
rect 49053 8579 49111 8585
rect 49234 8576 49240 8588
rect 49292 8576 49298 8628
rect 51813 8619 51871 8625
rect 51813 8585 51825 8619
rect 51859 8616 51871 8619
rect 51994 8616 52000 8628
rect 51859 8588 52000 8616
rect 51859 8585 51871 8588
rect 51813 8579 51871 8585
rect 51994 8576 52000 8588
rect 52052 8576 52058 8628
rect 53101 8619 53159 8625
rect 53101 8585 53113 8619
rect 53147 8616 53159 8619
rect 54110 8616 54116 8628
rect 53147 8588 54116 8616
rect 53147 8585 53159 8588
rect 53101 8579 53159 8585
rect 54110 8576 54116 8588
rect 54168 8576 54174 8628
rect 48222 8548 48228 8560
rect 35308 8520 38884 8548
rect 35308 8508 35314 8520
rect 35805 8483 35863 8489
rect 35805 8480 35817 8483
rect 35176 8452 35817 8480
rect 35805 8449 35817 8452
rect 35851 8480 35863 8483
rect 36262 8480 36268 8492
rect 35851 8452 36268 8480
rect 35851 8449 35863 8452
rect 35805 8443 35863 8449
rect 36262 8440 36268 8452
rect 36320 8440 36326 8492
rect 36354 8440 36360 8492
rect 36412 8480 36418 8492
rect 37826 8480 37832 8492
rect 36412 8452 37832 8480
rect 36412 8440 36418 8452
rect 37826 8440 37832 8452
rect 37884 8440 37890 8492
rect 38013 8483 38071 8489
rect 38013 8449 38025 8483
rect 38059 8480 38071 8483
rect 38102 8480 38108 8492
rect 38059 8452 38108 8480
rect 38059 8449 38071 8452
rect 38013 8443 38071 8449
rect 38102 8440 38108 8452
rect 38160 8440 38166 8492
rect 38746 8480 38752 8492
rect 38707 8452 38752 8480
rect 38746 8440 38752 8452
rect 38804 8440 38810 8492
rect 38856 8489 38884 8520
rect 40420 8520 41414 8548
rect 43272 8520 44772 8548
rect 38841 8483 38899 8489
rect 38841 8449 38853 8483
rect 38887 8449 38899 8483
rect 39482 8480 39488 8492
rect 39443 8452 39488 8480
rect 38841 8443 38899 8449
rect 33594 8412 33600 8424
rect 33555 8384 33600 8412
rect 33594 8372 33600 8384
rect 33652 8372 33658 8424
rect 35526 8412 35532 8424
rect 35487 8384 35532 8412
rect 35526 8372 35532 8384
rect 35584 8372 35590 8424
rect 36280 8412 36308 8440
rect 37277 8415 37335 8421
rect 37277 8412 37289 8415
rect 36280 8384 37289 8412
rect 37277 8381 37289 8384
rect 37323 8412 37335 8415
rect 37550 8412 37556 8424
rect 37323 8384 37556 8412
rect 37323 8381 37335 8384
rect 37277 8375 37335 8381
rect 37550 8372 37556 8384
rect 37608 8372 37614 8424
rect 38197 8347 38255 8353
rect 32355 8316 33456 8344
rect 33888 8316 34192 8344
rect 32355 8313 32367 8316
rect 32309 8307 32367 8313
rect 30423 8248 30512 8276
rect 30423 8245 30435 8248
rect 30377 8239 30435 8245
rect 32214 8236 32220 8288
rect 32272 8276 32278 8288
rect 33888 8276 33916 8316
rect 32272 8248 33916 8276
rect 32272 8236 32278 8248
rect 33962 8236 33968 8288
rect 34020 8276 34026 8288
rect 34057 8279 34115 8285
rect 34057 8276 34069 8279
rect 34020 8248 34069 8276
rect 34020 8236 34026 8248
rect 34057 8245 34069 8248
rect 34103 8245 34115 8279
rect 34164 8276 34192 8316
rect 38197 8313 38209 8347
rect 38243 8344 38255 8347
rect 38378 8344 38384 8356
rect 38243 8316 38384 8344
rect 38243 8313 38255 8316
rect 38197 8307 38255 8313
rect 38378 8304 38384 8316
rect 38436 8304 38442 8356
rect 38856 8344 38884 8443
rect 39482 8440 39488 8452
rect 39540 8440 39546 8492
rect 40310 8480 40316 8492
rect 40271 8452 40316 8480
rect 40310 8440 40316 8452
rect 40368 8440 40374 8492
rect 39500 8412 39528 8440
rect 40420 8412 40448 8520
rect 41138 8480 41144 8492
rect 41099 8452 41144 8480
rect 41138 8440 41144 8452
rect 41196 8440 41202 8492
rect 41386 8480 41414 8520
rect 42613 8483 42671 8489
rect 42613 8480 42625 8483
rect 41386 8452 42625 8480
rect 42613 8449 42625 8452
rect 42659 8449 42671 8483
rect 42613 8443 42671 8449
rect 42797 8483 42855 8489
rect 42797 8449 42809 8483
rect 42843 8480 42855 8483
rect 43257 8483 43315 8489
rect 43257 8480 43269 8483
rect 42843 8452 43269 8480
rect 42843 8449 42855 8452
rect 42797 8443 42855 8449
rect 43257 8449 43269 8452
rect 43303 8449 43315 8483
rect 43257 8443 43315 8449
rect 43346 8440 43352 8492
rect 43404 8480 43410 8492
rect 44744 8489 44772 8520
rect 46492 8520 48228 8548
rect 44085 8483 44143 8489
rect 44085 8480 44097 8483
rect 43404 8452 44097 8480
rect 43404 8440 43410 8452
rect 44085 8449 44097 8452
rect 44131 8449 44143 8483
rect 44085 8443 44143 8449
rect 44729 8483 44787 8489
rect 44729 8449 44741 8483
rect 44775 8480 44787 8483
rect 45278 8480 45284 8492
rect 44775 8452 45284 8480
rect 44775 8449 44787 8452
rect 44729 8443 44787 8449
rect 45278 8440 45284 8452
rect 45336 8440 45342 8492
rect 45462 8440 45468 8492
rect 45520 8480 45526 8492
rect 46201 8483 46259 8489
rect 46201 8480 46213 8483
rect 45520 8452 46213 8480
rect 45520 8440 45526 8452
rect 46201 8449 46213 8452
rect 46247 8449 46259 8483
rect 46201 8443 46259 8449
rect 39500 8384 40448 8412
rect 40770 8372 40776 8424
rect 40828 8412 40834 8424
rect 40865 8415 40923 8421
rect 40865 8412 40877 8415
rect 40828 8384 40877 8412
rect 40828 8372 40834 8384
rect 40865 8381 40877 8384
rect 40911 8381 40923 8415
rect 40865 8375 40923 8381
rect 42429 8415 42487 8421
rect 42429 8381 42441 8415
rect 42475 8412 42487 8415
rect 42518 8412 42524 8424
rect 42475 8384 42524 8412
rect 42475 8381 42487 8384
rect 42429 8375 42487 8381
rect 42518 8372 42524 8384
rect 42576 8412 42582 8424
rect 44634 8412 44640 8424
rect 42576 8384 44640 8412
rect 42576 8372 42582 8384
rect 44634 8372 44640 8384
rect 44692 8372 44698 8424
rect 45094 8372 45100 8424
rect 45152 8412 45158 8424
rect 45925 8415 45983 8421
rect 45925 8412 45937 8415
rect 45152 8384 45937 8412
rect 45152 8372 45158 8384
rect 45925 8381 45937 8384
rect 45971 8412 45983 8415
rect 46492 8412 46520 8520
rect 48222 8508 48228 8520
rect 48280 8508 48286 8560
rect 48406 8548 48412 8560
rect 48319 8520 48412 8548
rect 48406 8508 48412 8520
rect 48464 8548 48470 8560
rect 49142 8548 49148 8560
rect 48464 8520 49148 8548
rect 48464 8508 48470 8520
rect 49142 8508 49148 8520
rect 49200 8508 49206 8560
rect 50080 8520 53052 8548
rect 50080 8492 50108 8520
rect 46750 8480 46756 8492
rect 46711 8452 46756 8480
rect 46750 8440 46756 8452
rect 46808 8440 46814 8492
rect 46842 8440 46848 8492
rect 46900 8480 46906 8492
rect 49237 8483 49295 8489
rect 46900 8452 46945 8480
rect 46900 8440 46906 8452
rect 49237 8449 49249 8483
rect 49283 8480 49295 8483
rect 49326 8480 49332 8492
rect 49283 8452 49332 8480
rect 49283 8449 49295 8452
rect 49237 8443 49295 8449
rect 49326 8440 49332 8452
rect 49384 8440 49390 8492
rect 50062 8480 50068 8492
rect 50023 8452 50068 8480
rect 50062 8440 50068 8452
rect 50120 8440 50126 8492
rect 50798 8480 50804 8492
rect 50759 8452 50804 8480
rect 50798 8440 50804 8452
rect 50856 8440 50862 8492
rect 51534 8440 51540 8492
rect 51592 8480 51598 8492
rect 51629 8483 51687 8489
rect 51629 8480 51641 8483
rect 51592 8452 51641 8480
rect 51592 8440 51598 8452
rect 51629 8449 51641 8452
rect 51675 8480 51687 8483
rect 52917 8483 52975 8489
rect 52917 8480 52929 8483
rect 51675 8452 52929 8480
rect 51675 8449 51687 8452
rect 51629 8443 51687 8449
rect 52917 8449 52929 8452
rect 52963 8449 52975 8483
rect 52917 8443 52975 8449
rect 45971 8384 46520 8412
rect 45971 8381 45983 8384
rect 45925 8375 45983 8381
rect 46934 8372 46940 8424
rect 46992 8412 46998 8424
rect 48225 8415 48283 8421
rect 48225 8412 48237 8415
rect 46992 8384 48237 8412
rect 46992 8372 46998 8384
rect 48225 8381 48237 8384
rect 48271 8381 48283 8415
rect 48225 8375 48283 8381
rect 49421 8415 49479 8421
rect 49421 8381 49433 8415
rect 49467 8412 49479 8415
rect 50706 8412 50712 8424
rect 49467 8384 50712 8412
rect 49467 8381 49479 8384
rect 49421 8375 49479 8381
rect 50706 8372 50712 8384
rect 50764 8412 50770 8424
rect 51445 8415 51503 8421
rect 51445 8412 51457 8415
rect 50764 8384 51457 8412
rect 50764 8372 50770 8384
rect 51445 8381 51457 8384
rect 51491 8381 51503 8415
rect 51445 8375 51503 8381
rect 52733 8415 52791 8421
rect 52733 8381 52745 8415
rect 52779 8412 52791 8415
rect 53024 8412 53052 8520
rect 55766 8480 55772 8492
rect 53208 8452 55772 8480
rect 53208 8412 53236 8452
rect 55766 8440 55772 8452
rect 55824 8440 55830 8492
rect 52779 8384 53052 8412
rect 53116 8384 53236 8412
rect 52779 8381 52791 8384
rect 52733 8375 52791 8381
rect 44174 8344 44180 8356
rect 38856 8316 41000 8344
rect 40218 8276 40224 8288
rect 34164 8248 40224 8276
rect 34057 8239 34115 8245
rect 40218 8236 40224 8248
rect 40276 8236 40282 8288
rect 40972 8276 41000 8316
rect 41432 8316 44180 8344
rect 41432 8276 41460 8316
rect 44174 8304 44180 8316
rect 44232 8304 44238 8356
rect 46842 8304 46848 8356
rect 46900 8344 46906 8356
rect 48314 8344 48320 8356
rect 46900 8316 48320 8344
rect 46900 8304 46906 8316
rect 48314 8304 48320 8316
rect 48372 8304 48378 8356
rect 49694 8344 49700 8356
rect 49620 8316 49700 8344
rect 41874 8276 41880 8288
rect 40972 8248 41460 8276
rect 41835 8248 41880 8276
rect 41874 8236 41880 8248
rect 41932 8236 41938 8288
rect 46934 8236 46940 8288
rect 46992 8276 46998 8288
rect 47029 8279 47087 8285
rect 47029 8276 47041 8279
rect 46992 8248 47041 8276
rect 46992 8236 46998 8248
rect 47029 8245 47041 8248
rect 47075 8245 47087 8279
rect 47578 8276 47584 8288
rect 47539 8248 47584 8276
rect 47029 8239 47087 8245
rect 47578 8236 47584 8248
rect 47636 8236 47642 8288
rect 49142 8236 49148 8288
rect 49200 8276 49206 8288
rect 49620 8276 49648 8316
rect 49694 8304 49700 8316
rect 49752 8304 49758 8356
rect 49878 8344 49884 8356
rect 49839 8316 49884 8344
rect 49878 8304 49884 8316
rect 49936 8344 49942 8356
rect 51350 8344 51356 8356
rect 49936 8316 51356 8344
rect 49936 8304 49942 8316
rect 51350 8304 51356 8316
rect 51408 8304 51414 8356
rect 51460 8344 51488 8375
rect 52932 8356 52960 8384
rect 51460 8316 52868 8344
rect 50614 8276 50620 8288
rect 49200 8248 49648 8276
rect 50575 8248 50620 8276
rect 49200 8236 49206 8248
rect 50614 8236 50620 8248
rect 50672 8236 50678 8288
rect 52840 8276 52868 8316
rect 52914 8304 52920 8356
rect 52972 8304 52978 8356
rect 53116 8276 53144 8384
rect 54386 8372 54392 8424
rect 54444 8412 54450 8424
rect 54665 8415 54723 8421
rect 54665 8412 54677 8415
rect 54444 8384 54677 8412
rect 54444 8372 54450 8384
rect 54665 8381 54677 8384
rect 54711 8381 54723 8415
rect 54665 8375 54723 8381
rect 53190 8304 53196 8356
rect 53248 8344 53254 8356
rect 53561 8347 53619 8353
rect 53561 8344 53573 8347
rect 53248 8316 53573 8344
rect 53248 8304 53254 8316
rect 53561 8313 53573 8316
rect 53607 8313 53619 8347
rect 53561 8307 53619 8313
rect 54205 8347 54263 8353
rect 54205 8313 54217 8347
rect 54251 8344 54263 8347
rect 55306 8344 55312 8356
rect 54251 8316 55312 8344
rect 54251 8313 54263 8316
rect 54205 8307 54263 8313
rect 55306 8304 55312 8316
rect 55364 8304 55370 8356
rect 52840 8248 53144 8276
rect 1104 8186 58880 8208
rect 1104 8134 8174 8186
rect 8226 8134 8238 8186
rect 8290 8134 8302 8186
rect 8354 8134 8366 8186
rect 8418 8134 8430 8186
rect 8482 8134 22622 8186
rect 22674 8134 22686 8186
rect 22738 8134 22750 8186
rect 22802 8134 22814 8186
rect 22866 8134 22878 8186
rect 22930 8134 37070 8186
rect 37122 8134 37134 8186
rect 37186 8134 37198 8186
rect 37250 8134 37262 8186
rect 37314 8134 37326 8186
rect 37378 8134 51518 8186
rect 51570 8134 51582 8186
rect 51634 8134 51646 8186
rect 51698 8134 51710 8186
rect 51762 8134 51774 8186
rect 51826 8134 58880 8186
rect 1104 8112 58880 8134
rect 1762 8032 1768 8084
rect 1820 8072 1826 8084
rect 2038 8072 2044 8084
rect 1820 8044 2044 8072
rect 1820 8032 1826 8044
rect 2038 8032 2044 8044
rect 2096 8032 2102 8084
rect 3510 8032 3516 8084
rect 3568 8072 3574 8084
rect 6178 8072 6184 8084
rect 3568 8044 6184 8072
rect 3568 8032 3574 8044
rect 6178 8032 6184 8044
rect 6236 8032 6242 8084
rect 7745 8075 7803 8081
rect 7745 8041 7757 8075
rect 7791 8072 7803 8075
rect 10502 8072 10508 8084
rect 7791 8044 10508 8072
rect 7791 8041 7803 8044
rect 7745 8035 7803 8041
rect 10502 8032 10508 8044
rect 10560 8032 10566 8084
rect 10962 8032 10968 8084
rect 11020 8072 11026 8084
rect 11698 8072 11704 8084
rect 11020 8044 11704 8072
rect 11020 8032 11026 8044
rect 11698 8032 11704 8044
rect 11756 8032 11762 8084
rect 15841 8075 15899 8081
rect 14200 8044 15424 8072
rect 4525 8007 4583 8013
rect 4525 7973 4537 8007
rect 4571 8004 4583 8007
rect 5534 8004 5540 8016
rect 4571 7976 5540 8004
rect 4571 7973 4583 7976
rect 4525 7967 4583 7973
rect 5534 7964 5540 7976
rect 5592 7964 5598 8016
rect 9214 7964 9220 8016
rect 9272 7964 9278 8016
rect 11425 8007 11483 8013
rect 11425 7973 11437 8007
rect 11471 8004 11483 8007
rect 11471 7976 11928 8004
rect 11471 7973 11483 7976
rect 11425 7967 11483 7973
rect 2869 7939 2927 7945
rect 2869 7905 2881 7939
rect 2915 7936 2927 7939
rect 2958 7936 2964 7948
rect 2915 7908 2964 7936
rect 2915 7905 2927 7908
rect 2869 7899 2927 7905
rect 2958 7896 2964 7908
rect 3016 7896 3022 7948
rect 8294 7896 8300 7948
rect 8352 7936 8358 7948
rect 9232 7936 9260 7964
rect 8352 7908 9720 7936
rect 8352 7896 8358 7908
rect 1854 7868 1860 7880
rect 1815 7840 1860 7868
rect 1854 7828 1860 7840
rect 1912 7828 1918 7880
rect 2685 7871 2743 7877
rect 2685 7837 2697 7871
rect 2731 7868 2743 7871
rect 3510 7868 3516 7880
rect 2731 7840 3516 7868
rect 2731 7837 2743 7840
rect 2685 7831 2743 7837
rect 3510 7828 3516 7840
rect 3568 7828 3574 7880
rect 4338 7868 4344 7880
rect 4299 7840 4344 7868
rect 4338 7828 4344 7840
rect 4396 7828 4402 7880
rect 4982 7868 4988 7880
rect 4943 7840 4988 7868
rect 4982 7828 4988 7840
rect 5040 7828 5046 7880
rect 5629 7871 5687 7877
rect 5629 7837 5641 7871
rect 5675 7868 5687 7871
rect 5810 7868 5816 7880
rect 5675 7840 5816 7868
rect 5675 7837 5687 7840
rect 5629 7831 5687 7837
rect 5810 7828 5816 7840
rect 5868 7828 5874 7880
rect 5902 7828 5908 7880
rect 5960 7868 5966 7880
rect 7558 7868 7564 7880
rect 5960 7840 6005 7868
rect 7519 7840 7564 7868
rect 5960 7828 5966 7840
rect 7558 7828 7564 7840
rect 7616 7828 7622 7880
rect 8018 7828 8024 7880
rect 8076 7868 8082 7880
rect 8205 7871 8263 7877
rect 8205 7868 8217 7871
rect 8076 7840 8217 7868
rect 8076 7828 8082 7840
rect 8205 7837 8217 7840
rect 8251 7837 8263 7871
rect 9214 7868 9220 7880
rect 9175 7840 9220 7868
rect 8205 7831 8263 7837
rect 9214 7828 9220 7840
rect 9272 7828 9278 7880
rect 9692 7877 9720 7908
rect 9677 7871 9735 7877
rect 9677 7837 9689 7871
rect 9723 7868 9735 7871
rect 9858 7868 9864 7880
rect 9723 7840 9864 7868
rect 9723 7837 9735 7840
rect 9677 7831 9735 7837
rect 9858 7828 9864 7840
rect 9916 7828 9922 7880
rect 9953 7871 10011 7877
rect 9953 7837 9965 7871
rect 9999 7868 10011 7871
rect 11900 7868 11928 7976
rect 12434 7868 12440 7880
rect 9999 7840 10088 7868
rect 11900 7840 12440 7868
rect 9999 7837 10011 7840
rect 9953 7831 10011 7837
rect 10060 7800 10088 7840
rect 12434 7828 12440 7840
rect 12492 7828 12498 7880
rect 12618 7868 12624 7880
rect 12579 7840 12624 7868
rect 12618 7828 12624 7840
rect 12676 7828 12682 7880
rect 12897 7871 12955 7877
rect 12897 7837 12909 7871
rect 12943 7837 12955 7871
rect 12897 7831 12955 7837
rect 13357 7871 13415 7877
rect 13357 7837 13369 7871
rect 13403 7868 13415 7871
rect 13538 7868 13544 7880
rect 13403 7840 13544 7868
rect 13403 7837 13415 7840
rect 13357 7831 13415 7837
rect 5184 7772 10088 7800
rect 2038 7732 2044 7744
rect 1999 7704 2044 7732
rect 2038 7692 2044 7704
rect 2096 7692 2102 7744
rect 2498 7732 2504 7744
rect 2459 7704 2504 7732
rect 2498 7692 2504 7704
rect 2556 7692 2562 7744
rect 3881 7735 3939 7741
rect 3881 7701 3893 7735
rect 3927 7732 3939 7735
rect 4706 7732 4712 7744
rect 3927 7704 4712 7732
rect 3927 7701 3939 7704
rect 3881 7695 3939 7701
rect 4706 7692 4712 7704
rect 4764 7692 4770 7744
rect 5184 7741 5212 7772
rect 11698 7760 11704 7812
rect 11756 7800 11762 7812
rect 12912 7800 12940 7831
rect 13538 7828 13544 7840
rect 13596 7828 13602 7880
rect 14200 7877 14228 8044
rect 14369 8007 14427 8013
rect 14369 7973 14381 8007
rect 14415 8004 14427 8007
rect 14642 8004 14648 8016
rect 14415 7976 14648 8004
rect 14415 7973 14427 7976
rect 14369 7967 14427 7973
rect 14642 7964 14648 7976
rect 14700 7964 14706 8016
rect 15396 8004 15424 8044
rect 15841 8041 15853 8075
rect 15887 8072 15899 8075
rect 16206 8072 16212 8084
rect 15887 8044 16212 8072
rect 15887 8041 15899 8044
rect 15841 8035 15899 8041
rect 16206 8032 16212 8044
rect 16264 8032 16270 8084
rect 16574 8072 16580 8084
rect 16535 8044 16580 8072
rect 16574 8032 16580 8044
rect 16632 8032 16638 8084
rect 17862 8032 17868 8084
rect 17920 8072 17926 8084
rect 18049 8075 18107 8081
rect 18049 8072 18061 8075
rect 17920 8044 18061 8072
rect 17920 8032 17926 8044
rect 18049 8041 18061 8044
rect 18095 8041 18107 8075
rect 18782 8072 18788 8084
rect 18049 8035 18107 8041
rect 18524 8044 18788 8072
rect 17678 8004 17684 8016
rect 15396 7976 17684 8004
rect 17678 7964 17684 7976
rect 17736 7964 17742 8016
rect 14826 7936 14832 7948
rect 14787 7908 14832 7936
rect 14826 7896 14832 7908
rect 14884 7896 14890 7948
rect 14185 7871 14243 7877
rect 14185 7837 14197 7871
rect 14231 7837 14243 7871
rect 15105 7871 15163 7877
rect 15105 7868 15117 7871
rect 14185 7831 14243 7837
rect 15028 7840 15117 7868
rect 11756 7772 13676 7800
rect 11756 7760 11762 7772
rect 5169 7735 5227 7741
rect 5169 7701 5181 7735
rect 5215 7701 5227 7735
rect 5169 7695 5227 7701
rect 5350 7692 5356 7744
rect 5408 7732 5414 7744
rect 6641 7735 6699 7741
rect 6641 7732 6653 7735
rect 5408 7704 6653 7732
rect 5408 7692 5414 7704
rect 6641 7701 6653 7704
rect 6687 7732 6699 7735
rect 7374 7732 7380 7744
rect 6687 7704 7380 7732
rect 6687 7701 6699 7704
rect 6641 7695 6699 7701
rect 7374 7692 7380 7704
rect 7432 7732 7438 7744
rect 8202 7732 8208 7744
rect 7432 7704 8208 7732
rect 7432 7692 7438 7704
rect 8202 7692 8208 7704
rect 8260 7692 8266 7744
rect 8389 7735 8447 7741
rect 8389 7701 8401 7735
rect 8435 7732 8447 7735
rect 10042 7732 10048 7744
rect 8435 7704 10048 7732
rect 8435 7701 8447 7704
rect 8389 7695 8447 7701
rect 10042 7692 10048 7704
rect 10100 7692 10106 7744
rect 10686 7732 10692 7744
rect 10647 7704 10692 7732
rect 10686 7692 10692 7704
rect 10744 7732 10750 7744
rect 11885 7735 11943 7741
rect 11885 7732 11897 7735
rect 10744 7704 11897 7732
rect 10744 7692 10750 7704
rect 11885 7701 11897 7704
rect 11931 7701 11943 7735
rect 11885 7695 11943 7701
rect 13262 7692 13268 7744
rect 13320 7732 13326 7744
rect 13541 7735 13599 7741
rect 13541 7732 13553 7735
rect 13320 7704 13553 7732
rect 13320 7692 13326 7704
rect 13541 7701 13553 7704
rect 13587 7701 13599 7735
rect 13648 7732 13676 7772
rect 14642 7760 14648 7812
rect 14700 7800 14706 7812
rect 15028 7800 15056 7840
rect 15105 7837 15117 7840
rect 15151 7837 15163 7871
rect 15105 7831 15163 7837
rect 16390 7828 16396 7880
rect 16448 7868 16454 7880
rect 16761 7871 16819 7877
rect 16761 7868 16773 7871
rect 16448 7840 16773 7868
rect 16448 7828 16454 7840
rect 16761 7837 16773 7840
rect 16807 7837 16819 7871
rect 16942 7868 16948 7880
rect 16903 7840 16948 7868
rect 16761 7831 16819 7837
rect 16942 7828 16948 7840
rect 17000 7828 17006 7880
rect 17126 7828 17132 7880
rect 17184 7868 17190 7880
rect 17865 7871 17923 7877
rect 17865 7868 17877 7871
rect 17184 7840 17877 7868
rect 17184 7828 17190 7840
rect 17865 7837 17877 7840
rect 17911 7837 17923 7871
rect 17865 7831 17923 7837
rect 18049 7871 18107 7877
rect 18049 7837 18061 7871
rect 18095 7868 18107 7871
rect 18414 7868 18420 7880
rect 18095 7840 18420 7868
rect 18095 7837 18107 7840
rect 18049 7831 18107 7837
rect 18414 7828 18420 7840
rect 18472 7828 18478 7880
rect 18524 7877 18552 8044
rect 18782 8032 18788 8044
rect 18840 8072 18846 8084
rect 18840 8044 19748 8072
rect 18840 8032 18846 8044
rect 19518 8004 19524 8016
rect 18708 7976 19524 8004
rect 18708 7877 18736 7976
rect 19518 7964 19524 7976
rect 19576 7964 19582 8016
rect 19720 8004 19748 8044
rect 19794 8032 19800 8084
rect 19852 8072 19858 8084
rect 21082 8072 21088 8084
rect 19852 8044 21088 8072
rect 19852 8032 19858 8044
rect 21082 8032 21088 8044
rect 21140 8032 21146 8084
rect 22741 8075 22799 8081
rect 22741 8041 22753 8075
rect 22787 8072 22799 8075
rect 23014 8072 23020 8084
rect 22787 8044 23020 8072
rect 22787 8041 22799 8044
rect 22741 8035 22799 8041
rect 23014 8032 23020 8044
rect 23072 8032 23078 8084
rect 23658 8032 23664 8084
rect 23716 8072 23722 8084
rect 24397 8075 24455 8081
rect 24397 8072 24409 8075
rect 23716 8044 24409 8072
rect 23716 8032 23722 8044
rect 24397 8041 24409 8044
rect 24443 8041 24455 8075
rect 24397 8035 24455 8041
rect 24854 8032 24860 8084
rect 24912 8072 24918 8084
rect 25501 8075 25559 8081
rect 25501 8072 25513 8075
rect 24912 8044 25513 8072
rect 24912 8032 24918 8044
rect 25501 8041 25513 8044
rect 25547 8041 25559 8075
rect 25501 8035 25559 8041
rect 25958 8032 25964 8084
rect 26016 8072 26022 8084
rect 26881 8075 26939 8081
rect 26881 8072 26893 8075
rect 26016 8044 26893 8072
rect 26016 8032 26022 8044
rect 26881 8041 26893 8044
rect 26927 8041 26939 8075
rect 26881 8035 26939 8041
rect 27614 8032 27620 8084
rect 27672 8072 27678 8084
rect 28442 8072 28448 8084
rect 27672 8044 28448 8072
rect 27672 8032 27678 8044
rect 28442 8032 28448 8044
rect 28500 8032 28506 8084
rect 28718 8072 28724 8084
rect 28679 8044 28724 8072
rect 28718 8032 28724 8044
rect 28776 8032 28782 8084
rect 30650 8032 30656 8084
rect 30708 8072 30714 8084
rect 32677 8075 32735 8081
rect 32677 8072 32689 8075
rect 30708 8044 32689 8072
rect 30708 8032 30714 8044
rect 32677 8041 32689 8044
rect 32723 8041 32735 8075
rect 35066 8072 35072 8084
rect 35027 8044 35072 8072
rect 32677 8035 32735 8041
rect 35066 8032 35072 8044
rect 35124 8032 35130 8084
rect 38381 8075 38439 8081
rect 38381 8041 38393 8075
rect 38427 8072 38439 8075
rect 41322 8072 41328 8084
rect 38427 8044 41328 8072
rect 38427 8041 38439 8044
rect 38381 8035 38439 8041
rect 41322 8032 41328 8044
rect 41380 8032 41386 8084
rect 42518 8072 42524 8084
rect 41524 8044 42524 8072
rect 25774 8004 25780 8016
rect 19720 7976 25780 8004
rect 25774 7964 25780 7976
rect 25832 7964 25838 8016
rect 26050 7964 26056 8016
rect 26108 8004 26114 8016
rect 33226 8004 33232 8016
rect 26108 7976 33232 8004
rect 26108 7964 26114 7976
rect 33226 7964 33232 7976
rect 33284 7964 33290 8016
rect 33505 8007 33563 8013
rect 33505 7973 33517 8007
rect 33551 8004 33563 8007
rect 39482 8004 39488 8016
rect 33551 7976 39488 8004
rect 33551 7973 33563 7976
rect 33505 7967 33563 7973
rect 39482 7964 39488 7976
rect 39540 7964 39546 8016
rect 40218 8004 40224 8016
rect 40131 7976 40224 8004
rect 40218 7964 40224 7976
rect 40276 8004 40282 8016
rect 41524 8004 41552 8044
rect 42518 8032 42524 8044
rect 42576 8032 42582 8084
rect 43257 8075 43315 8081
rect 43257 8041 43269 8075
rect 43303 8072 43315 8075
rect 43346 8072 43352 8084
rect 43303 8044 43352 8072
rect 43303 8041 43315 8044
rect 43257 8035 43315 8041
rect 43346 8032 43352 8044
rect 43404 8032 43410 8084
rect 46290 8072 46296 8084
rect 46251 8044 46296 8072
rect 46290 8032 46296 8044
rect 46348 8032 46354 8084
rect 46382 8032 46388 8084
rect 46440 8072 46446 8084
rect 46753 8075 46811 8081
rect 46753 8072 46765 8075
rect 46440 8044 46765 8072
rect 46440 8032 46446 8044
rect 46753 8041 46765 8044
rect 46799 8041 46811 8075
rect 46753 8035 46811 8041
rect 49605 8075 49663 8081
rect 49605 8041 49617 8075
rect 49651 8072 49663 8075
rect 50798 8072 50804 8084
rect 49651 8044 50804 8072
rect 49651 8041 49663 8044
rect 49605 8035 49663 8041
rect 50798 8032 50804 8044
rect 50856 8032 50862 8084
rect 51166 8072 51172 8084
rect 51127 8044 51172 8072
rect 51166 8032 51172 8044
rect 51224 8032 51230 8084
rect 51350 8032 51356 8084
rect 51408 8072 51414 8084
rect 51629 8075 51687 8081
rect 51629 8072 51641 8075
rect 51408 8044 51641 8072
rect 51408 8032 51414 8044
rect 51629 8041 51641 8044
rect 51675 8041 51687 8075
rect 51629 8035 51687 8041
rect 49326 8004 49332 8016
rect 40276 7976 41552 8004
rect 48700 7976 49332 8004
rect 40276 7964 40282 7976
rect 19702 7896 19708 7948
rect 19760 7936 19766 7948
rect 19760 7908 21496 7936
rect 19760 7896 19766 7908
rect 18509 7871 18567 7877
rect 18509 7837 18521 7871
rect 18555 7837 18567 7871
rect 18509 7831 18567 7837
rect 18693 7871 18751 7877
rect 18693 7837 18705 7871
rect 18739 7837 18751 7871
rect 19242 7868 19248 7880
rect 19203 7840 19248 7868
rect 18693 7831 18751 7837
rect 19242 7828 19248 7840
rect 19300 7828 19306 7880
rect 20162 7828 20168 7880
rect 20220 7868 20226 7880
rect 20533 7871 20591 7877
rect 20533 7868 20545 7871
rect 20220 7840 20545 7868
rect 20220 7828 20226 7840
rect 20533 7837 20545 7840
rect 20579 7837 20591 7871
rect 20533 7831 20591 7837
rect 20809 7871 20867 7877
rect 20809 7837 20821 7871
rect 20855 7868 20867 7871
rect 20898 7868 20904 7880
rect 20855 7840 20904 7868
rect 20855 7837 20867 7840
rect 20809 7831 20867 7837
rect 20898 7828 20904 7840
rect 20956 7828 20962 7880
rect 21266 7868 21272 7880
rect 21227 7840 21272 7868
rect 21266 7828 21272 7840
rect 21324 7828 21330 7880
rect 21468 7877 21496 7908
rect 23014 7896 23020 7948
rect 23072 7936 23078 7948
rect 23290 7936 23296 7948
rect 23072 7908 23296 7936
rect 23072 7896 23078 7908
rect 23290 7896 23296 7908
rect 23348 7896 23354 7948
rect 26068 7936 26096 7964
rect 26418 7936 26424 7948
rect 23676 7908 26096 7936
rect 26379 7908 26424 7936
rect 23676 7877 23704 7908
rect 26418 7896 26424 7908
rect 26476 7896 26482 7948
rect 26970 7896 26976 7948
rect 27028 7936 27034 7948
rect 34057 7939 34115 7945
rect 27028 7908 34008 7936
rect 27028 7896 27034 7908
rect 21453 7871 21511 7877
rect 21453 7837 21465 7871
rect 21499 7837 21511 7871
rect 21453 7831 21511 7837
rect 22189 7871 22247 7877
rect 22189 7837 22201 7871
rect 22235 7868 22247 7871
rect 23661 7871 23719 7877
rect 23661 7868 23673 7871
rect 22235 7840 23673 7868
rect 22235 7837 22247 7840
rect 22189 7831 22247 7837
rect 23661 7837 23673 7840
rect 23707 7837 23719 7871
rect 23661 7831 23719 7837
rect 23845 7871 23903 7877
rect 23845 7837 23857 7871
rect 23891 7837 23903 7871
rect 24578 7868 24584 7880
rect 24539 7840 24584 7868
rect 23845 7831 23903 7837
rect 14700 7772 15056 7800
rect 14700 7760 14706 7772
rect 17954 7760 17960 7812
rect 18012 7800 18018 7812
rect 18601 7803 18659 7809
rect 18601 7800 18613 7803
rect 18012 7772 18613 7800
rect 18012 7760 18018 7772
rect 18601 7769 18613 7772
rect 18647 7800 18659 7803
rect 20254 7800 20260 7812
rect 18647 7772 20260 7800
rect 18647 7769 18659 7772
rect 18601 7763 18659 7769
rect 20254 7760 20260 7772
rect 20312 7760 20318 7812
rect 21174 7760 21180 7812
rect 21232 7800 21238 7812
rect 22204 7800 22232 7831
rect 21232 7772 22232 7800
rect 21232 7760 21238 7772
rect 22370 7760 22376 7812
rect 22428 7800 22434 7812
rect 22833 7803 22891 7809
rect 22833 7800 22845 7803
rect 22428 7772 22845 7800
rect 22428 7760 22434 7772
rect 22833 7769 22845 7772
rect 22879 7800 22891 7803
rect 23474 7800 23480 7812
rect 22879 7772 23480 7800
rect 22879 7769 22891 7772
rect 22833 7763 22891 7769
rect 23474 7760 23480 7772
rect 23532 7760 23538 7812
rect 23750 7800 23756 7812
rect 23711 7772 23756 7800
rect 23750 7760 23756 7772
rect 23808 7760 23814 7812
rect 15194 7732 15200 7744
rect 13648 7704 15200 7732
rect 13541 7695 13599 7701
rect 15194 7692 15200 7704
rect 15252 7692 15258 7744
rect 19429 7735 19487 7741
rect 19429 7701 19441 7735
rect 19475 7732 19487 7735
rect 19518 7732 19524 7744
rect 19475 7704 19524 7732
rect 19475 7701 19487 7704
rect 19429 7695 19487 7701
rect 19518 7692 19524 7704
rect 19576 7692 19582 7744
rect 21634 7732 21640 7744
rect 21595 7704 21640 7732
rect 21634 7692 21640 7704
rect 21692 7692 21698 7744
rect 23860 7732 23888 7831
rect 24578 7828 24584 7840
rect 24636 7828 24642 7880
rect 24762 7868 24768 7880
rect 24723 7840 24768 7868
rect 24762 7828 24768 7840
rect 24820 7828 24826 7880
rect 25869 7871 25927 7877
rect 25869 7837 25881 7871
rect 25915 7868 25927 7871
rect 25958 7868 25964 7880
rect 25915 7840 25964 7868
rect 25915 7837 25927 7840
rect 25869 7831 25927 7837
rect 25958 7828 25964 7840
rect 26016 7828 26022 7880
rect 27065 7871 27123 7877
rect 27065 7837 27077 7871
rect 27111 7868 27123 7871
rect 27430 7868 27436 7880
rect 27111 7840 27436 7868
rect 27111 7837 27123 7840
rect 27065 7831 27123 7837
rect 27430 7828 27436 7840
rect 27488 7828 27494 7880
rect 27525 7871 27583 7877
rect 27525 7837 27537 7871
rect 27571 7868 27583 7871
rect 27614 7868 27620 7880
rect 27571 7840 27620 7868
rect 27571 7837 27583 7840
rect 27525 7831 27583 7837
rect 24596 7800 24624 7828
rect 25685 7803 25743 7809
rect 25685 7800 25697 7803
rect 24596 7772 25697 7800
rect 25685 7769 25697 7772
rect 25731 7769 25743 7803
rect 25685 7763 25743 7769
rect 26786 7760 26792 7812
rect 26844 7800 26850 7812
rect 27540 7800 27568 7831
rect 27614 7828 27620 7840
rect 27672 7828 27678 7880
rect 27798 7868 27804 7880
rect 27759 7840 27804 7868
rect 27798 7828 27804 7840
rect 27856 7828 27862 7880
rect 27890 7828 27896 7880
rect 27948 7868 27954 7880
rect 28902 7868 28908 7880
rect 27948 7840 27993 7868
rect 28863 7840 28908 7868
rect 27948 7828 27954 7840
rect 28902 7828 28908 7840
rect 28960 7828 28966 7880
rect 29730 7828 29736 7880
rect 29788 7868 29794 7880
rect 30653 7871 30711 7877
rect 30653 7868 30665 7871
rect 29788 7840 30665 7868
rect 29788 7828 29794 7840
rect 30653 7837 30665 7840
rect 30699 7837 30711 7871
rect 30653 7831 30711 7837
rect 31205 7871 31263 7877
rect 31205 7837 31217 7871
rect 31251 7837 31263 7871
rect 31205 7831 31263 7837
rect 26844 7772 27568 7800
rect 26844 7760 26850 7772
rect 28718 7760 28724 7812
rect 28776 7800 28782 7812
rect 30009 7803 30067 7809
rect 30009 7800 30021 7803
rect 28776 7772 30021 7800
rect 28776 7760 28782 7772
rect 30009 7769 30021 7772
rect 30055 7769 30067 7803
rect 30009 7763 30067 7769
rect 30374 7760 30380 7812
rect 30432 7800 30438 7812
rect 31220 7800 31248 7831
rect 31294 7828 31300 7880
rect 31352 7868 31358 7880
rect 32033 7871 32091 7877
rect 32033 7868 32045 7871
rect 31352 7840 32045 7868
rect 31352 7828 31358 7840
rect 32033 7837 32045 7840
rect 32079 7837 32091 7871
rect 32214 7868 32220 7880
rect 32175 7840 32220 7868
rect 32033 7831 32091 7837
rect 32214 7828 32220 7840
rect 32272 7828 32278 7880
rect 32858 7868 32864 7880
rect 32819 7840 32864 7868
rect 32858 7828 32864 7840
rect 32916 7828 32922 7880
rect 33321 7871 33379 7877
rect 33321 7837 33333 7871
rect 33367 7868 33379 7871
rect 33410 7868 33416 7880
rect 33367 7840 33416 7868
rect 33367 7837 33379 7840
rect 33321 7831 33379 7837
rect 33410 7828 33416 7840
rect 33468 7828 33474 7880
rect 33980 7877 34008 7908
rect 34057 7905 34069 7939
rect 34103 7936 34115 7939
rect 34103 7908 34744 7936
rect 34103 7905 34115 7908
rect 34057 7899 34115 7905
rect 34716 7877 34744 7908
rect 36170 7896 36176 7948
rect 36228 7936 36234 7948
rect 36357 7939 36415 7945
rect 36357 7936 36369 7939
rect 36228 7908 36369 7936
rect 36228 7896 36234 7908
rect 36357 7905 36369 7908
rect 36403 7936 36415 7939
rect 37369 7939 37427 7945
rect 36403 7908 37320 7936
rect 36403 7905 36415 7908
rect 36357 7899 36415 7905
rect 33505 7871 33563 7877
rect 33505 7837 33517 7871
rect 33551 7837 33563 7871
rect 33505 7831 33563 7837
rect 33965 7871 34023 7877
rect 33965 7837 33977 7871
rect 34011 7837 34023 7871
rect 33965 7831 34023 7837
rect 34149 7871 34207 7877
rect 34149 7837 34161 7871
rect 34195 7837 34207 7871
rect 34149 7831 34207 7837
rect 34701 7871 34759 7877
rect 34701 7837 34713 7871
rect 34747 7868 34759 7871
rect 35250 7868 35256 7880
rect 34747 7840 35256 7868
rect 34747 7837 34759 7840
rect 34701 7831 34759 7837
rect 33520 7800 33548 7831
rect 34164 7800 34192 7831
rect 35250 7828 35256 7840
rect 35308 7828 35314 7880
rect 36630 7868 36636 7880
rect 36591 7840 36636 7868
rect 36630 7828 36636 7840
rect 36688 7828 36694 7880
rect 36906 7828 36912 7880
rect 36964 7868 36970 7880
rect 37185 7871 37243 7877
rect 37185 7868 37197 7871
rect 36964 7840 37197 7868
rect 36964 7828 36970 7840
rect 37185 7837 37197 7840
rect 37231 7837 37243 7871
rect 37292 7868 37320 7908
rect 37369 7905 37381 7939
rect 37415 7936 37427 7939
rect 45278 7936 45284 7948
rect 37415 7908 40540 7936
rect 45239 7908 45284 7936
rect 37415 7905 37427 7908
rect 37369 7899 37427 7905
rect 38013 7871 38071 7877
rect 38013 7868 38025 7871
rect 37292 7840 38025 7868
rect 37185 7831 37243 7837
rect 38013 7837 38025 7840
rect 38059 7837 38071 7871
rect 38013 7831 38071 7837
rect 38197 7871 38255 7877
rect 38197 7837 38209 7871
rect 38243 7837 38255 7871
rect 38838 7868 38844 7880
rect 38799 7840 38844 7868
rect 38197 7831 38255 7837
rect 34882 7800 34888 7812
rect 30432 7772 31248 7800
rect 32048 7772 34192 7800
rect 34843 7772 34888 7800
rect 30432 7760 30438 7772
rect 32048 7744 32076 7772
rect 34882 7760 34888 7772
rect 34940 7760 34946 7812
rect 38102 7800 38108 7812
rect 37476 7772 38108 7800
rect 37476 7744 37504 7772
rect 38102 7760 38108 7772
rect 38160 7800 38166 7812
rect 38212 7800 38240 7831
rect 38838 7828 38844 7840
rect 38896 7828 38902 7880
rect 39025 7871 39083 7877
rect 39025 7837 39037 7871
rect 39071 7837 39083 7871
rect 39025 7831 39083 7837
rect 38160 7772 38240 7800
rect 38160 7760 38166 7772
rect 25222 7732 25228 7744
rect 23860 7704 25228 7732
rect 25222 7692 25228 7704
rect 25280 7692 25286 7744
rect 25774 7692 25780 7744
rect 25832 7732 25838 7744
rect 30101 7735 30159 7741
rect 30101 7732 30113 7735
rect 25832 7704 30113 7732
rect 25832 7692 25838 7704
rect 30101 7701 30113 7704
rect 30147 7732 30159 7735
rect 30742 7732 30748 7744
rect 30147 7704 30748 7732
rect 30147 7701 30159 7704
rect 30101 7695 30159 7701
rect 30742 7692 30748 7704
rect 30800 7692 30806 7744
rect 31389 7735 31447 7741
rect 31389 7701 31401 7735
rect 31435 7732 31447 7735
rect 31570 7732 31576 7744
rect 31435 7704 31576 7732
rect 31435 7701 31447 7704
rect 31389 7695 31447 7701
rect 31570 7692 31576 7704
rect 31628 7692 31634 7744
rect 31846 7732 31852 7744
rect 31807 7704 31852 7732
rect 31846 7692 31852 7704
rect 31904 7692 31910 7744
rect 32030 7692 32036 7744
rect 32088 7692 32094 7744
rect 32306 7692 32312 7744
rect 32364 7732 32370 7744
rect 37458 7732 37464 7744
rect 32364 7704 37464 7732
rect 32364 7692 32370 7704
rect 37458 7692 37464 7704
rect 37516 7692 37522 7744
rect 38212 7732 38240 7772
rect 39040 7732 39068 7831
rect 40402 7800 40408 7812
rect 40363 7772 40408 7800
rect 40402 7760 40408 7772
rect 40460 7760 40466 7812
rect 40512 7800 40540 7908
rect 45278 7896 45284 7908
rect 45336 7896 45342 7948
rect 48314 7936 48320 7948
rect 46124 7908 48320 7936
rect 40586 7828 40592 7880
rect 40644 7868 40650 7880
rect 41417 7871 41475 7877
rect 41417 7868 41429 7871
rect 40644 7840 41429 7868
rect 40644 7828 40650 7840
rect 41417 7837 41429 7840
rect 41463 7837 41475 7871
rect 41690 7868 41696 7880
rect 41651 7840 41696 7868
rect 41417 7831 41475 7837
rect 41690 7828 41696 7840
rect 41748 7828 41754 7880
rect 43070 7868 43076 7880
rect 42812 7840 43076 7868
rect 42812 7800 42840 7840
rect 43070 7828 43076 7840
rect 43128 7828 43134 7880
rect 44174 7868 44180 7880
rect 44135 7840 44180 7868
rect 44174 7828 44180 7840
rect 44232 7828 44238 7880
rect 45557 7871 45615 7877
rect 45557 7837 45569 7871
rect 45603 7868 45615 7871
rect 46014 7868 46020 7880
rect 45603 7840 46020 7868
rect 45603 7837 45615 7840
rect 45557 7831 45615 7837
rect 46014 7828 46020 7840
rect 46072 7828 46078 7880
rect 40512 7772 42840 7800
rect 42886 7760 42892 7812
rect 42944 7800 42950 7812
rect 45370 7800 45376 7812
rect 42944 7772 42989 7800
rect 44376 7772 45376 7800
rect 42944 7760 42950 7772
rect 38212 7704 39068 7732
rect 39209 7735 39267 7741
rect 39209 7701 39221 7735
rect 39255 7732 39267 7735
rect 40218 7732 40224 7744
rect 39255 7704 40224 7732
rect 39255 7701 39267 7704
rect 39209 7695 39267 7701
rect 40218 7692 40224 7704
rect 40276 7692 40282 7744
rect 41414 7692 41420 7744
rect 41472 7732 41478 7744
rect 44376 7741 44404 7772
rect 45370 7760 45376 7772
rect 45428 7800 45434 7812
rect 46124 7800 46152 7908
rect 48314 7896 48320 7908
rect 48372 7936 48378 7948
rect 48700 7936 48728 7976
rect 49326 7964 49332 7976
rect 49384 7964 49390 8016
rect 48372 7908 48728 7936
rect 48372 7896 48378 7908
rect 46934 7868 46940 7880
rect 46895 7840 46940 7868
rect 46934 7828 46940 7840
rect 46992 7828 46998 7880
rect 47765 7871 47823 7877
rect 47765 7837 47777 7871
rect 47811 7868 47823 7871
rect 48409 7871 48467 7877
rect 48409 7868 48421 7871
rect 47811 7840 48421 7868
rect 47811 7837 47823 7840
rect 47765 7831 47823 7837
rect 48409 7837 48421 7840
rect 48455 7837 48467 7871
rect 48409 7831 48467 7837
rect 48593 7871 48651 7877
rect 48593 7837 48605 7871
rect 48639 7868 48651 7871
rect 48700 7868 48728 7908
rect 48777 7939 48835 7945
rect 48777 7905 48789 7939
rect 48823 7936 48835 7939
rect 50062 7936 50068 7948
rect 48823 7908 50068 7936
rect 48823 7905 48835 7908
rect 48777 7899 48835 7905
rect 50062 7896 50068 7908
rect 50120 7896 50126 7948
rect 48639 7840 48728 7868
rect 48639 7837 48651 7840
rect 48593 7831 48651 7837
rect 49142 7828 49148 7880
rect 49200 7868 49206 7880
rect 49237 7871 49295 7877
rect 49237 7868 49249 7871
rect 49200 7840 49249 7868
rect 49200 7828 49206 7840
rect 49237 7837 49249 7840
rect 49283 7837 49295 7871
rect 49237 7831 49295 7837
rect 49326 7828 49332 7880
rect 49384 7868 49390 7880
rect 49421 7871 49479 7877
rect 49421 7868 49433 7871
rect 49384 7840 49433 7868
rect 49384 7828 49390 7840
rect 49421 7837 49433 7840
rect 49467 7837 49479 7871
rect 49421 7831 49479 7837
rect 50157 7871 50215 7877
rect 50157 7837 50169 7871
rect 50203 7868 50215 7871
rect 50338 7868 50344 7880
rect 50203 7840 50344 7868
rect 50203 7837 50215 7840
rect 50157 7831 50215 7837
rect 50338 7828 50344 7840
rect 50396 7828 50402 7880
rect 50433 7871 50491 7877
rect 50433 7837 50445 7871
rect 50479 7837 50491 7871
rect 50433 7831 50491 7837
rect 50448 7800 50476 7831
rect 53098 7828 53104 7880
rect 53156 7868 53162 7880
rect 53929 7871 53987 7877
rect 53929 7868 53941 7871
rect 53156 7840 53941 7868
rect 53156 7828 53162 7840
rect 53929 7837 53941 7840
rect 53975 7837 53987 7871
rect 53929 7831 53987 7837
rect 45428 7772 46152 7800
rect 47964 7772 50476 7800
rect 45428 7760 45434 7772
rect 42429 7735 42487 7741
rect 42429 7732 42441 7735
rect 41472 7704 42441 7732
rect 41472 7692 41478 7704
rect 42429 7701 42441 7704
rect 42475 7701 42487 7735
rect 42429 7695 42487 7701
rect 44361 7735 44419 7741
rect 44361 7701 44373 7735
rect 44407 7701 44419 7735
rect 44361 7695 44419 7701
rect 44634 7692 44640 7744
rect 44692 7732 44698 7744
rect 47578 7732 47584 7744
rect 44692 7704 47584 7732
rect 44692 7692 44698 7704
rect 47578 7692 47584 7704
rect 47636 7692 47642 7744
rect 47964 7741 47992 7772
rect 52454 7760 52460 7812
rect 52512 7800 52518 7812
rect 53377 7803 53435 7809
rect 53377 7800 53389 7803
rect 52512 7772 53389 7800
rect 52512 7760 52518 7772
rect 53377 7769 53389 7772
rect 53423 7800 53435 7803
rect 54573 7803 54631 7809
rect 54573 7800 54585 7803
rect 53423 7772 54585 7800
rect 53423 7769 53435 7772
rect 53377 7763 53435 7769
rect 54573 7769 54585 7772
rect 54619 7769 54631 7803
rect 54573 7763 54631 7769
rect 47949 7735 48007 7741
rect 47949 7701 47961 7735
rect 47995 7701 48007 7735
rect 52178 7732 52184 7744
rect 52139 7704 52184 7732
rect 47949 7695 48007 7701
rect 52178 7692 52184 7704
rect 52236 7692 52242 7744
rect 52730 7732 52736 7744
rect 52691 7704 52736 7732
rect 52730 7692 52736 7704
rect 52788 7692 52794 7744
rect 54113 7735 54171 7741
rect 54113 7701 54125 7735
rect 54159 7732 54171 7735
rect 54202 7732 54208 7744
rect 54159 7704 54208 7732
rect 54159 7701 54171 7704
rect 54113 7695 54171 7701
rect 54202 7692 54208 7704
rect 54260 7692 54266 7744
rect 55306 7732 55312 7744
rect 55267 7704 55312 7732
rect 55306 7692 55312 7704
rect 55364 7692 55370 7744
rect 1104 7642 58880 7664
rect 1104 7590 15398 7642
rect 15450 7590 15462 7642
rect 15514 7590 15526 7642
rect 15578 7590 15590 7642
rect 15642 7590 15654 7642
rect 15706 7590 29846 7642
rect 29898 7590 29910 7642
rect 29962 7590 29974 7642
rect 30026 7590 30038 7642
rect 30090 7590 30102 7642
rect 30154 7590 44294 7642
rect 44346 7590 44358 7642
rect 44410 7590 44422 7642
rect 44474 7590 44486 7642
rect 44538 7590 44550 7642
rect 44602 7590 58880 7642
rect 1104 7568 58880 7590
rect 1765 7531 1823 7537
rect 1765 7497 1777 7531
rect 1811 7528 1823 7531
rect 4246 7528 4252 7540
rect 1811 7500 4252 7528
rect 1811 7497 1823 7500
rect 1765 7491 1823 7497
rect 4246 7488 4252 7500
rect 4304 7488 4310 7540
rect 4338 7488 4344 7540
rect 4396 7528 4402 7540
rect 6365 7531 6423 7537
rect 6365 7528 6377 7531
rect 4396 7500 6377 7528
rect 4396 7488 4402 7500
rect 6365 7497 6377 7500
rect 6411 7497 6423 7531
rect 7742 7528 7748 7540
rect 6365 7491 6423 7497
rect 7392 7500 7748 7528
rect 2038 7420 2044 7472
rect 2096 7460 2102 7472
rect 2096 7432 4936 7460
rect 2096 7420 2102 7432
rect 1578 7392 1584 7404
rect 1539 7364 1584 7392
rect 1578 7352 1584 7364
rect 1636 7352 1642 7404
rect 2409 7395 2467 7401
rect 2409 7361 2421 7395
rect 2455 7392 2467 7395
rect 3237 7395 3295 7401
rect 3237 7392 3249 7395
rect 2455 7364 3249 7392
rect 2455 7361 2467 7364
rect 2409 7355 2467 7361
rect 3237 7361 3249 7364
rect 3283 7361 3295 7395
rect 3418 7392 3424 7404
rect 3379 7364 3424 7392
rect 3237 7355 3295 7361
rect 2593 7327 2651 7333
rect 2593 7293 2605 7327
rect 2639 7293 2651 7327
rect 3252 7324 3280 7355
rect 3418 7352 3424 7364
rect 3476 7352 3482 7404
rect 4908 7401 4936 7432
rect 5442 7420 5448 7472
rect 5500 7460 5506 7472
rect 5500 7432 6684 7460
rect 5500 7420 5506 7432
rect 4893 7395 4951 7401
rect 4893 7361 4905 7395
rect 4939 7361 4951 7395
rect 4893 7355 4951 7361
rect 5629 7395 5687 7401
rect 5629 7361 5641 7395
rect 5675 7392 5687 7395
rect 6270 7392 6276 7404
rect 5675 7364 6276 7392
rect 5675 7361 5687 7364
rect 5629 7355 5687 7361
rect 6270 7352 6276 7364
rect 6328 7352 6334 7404
rect 6362 7352 6368 7404
rect 6420 7392 6426 7404
rect 6656 7401 6684 7432
rect 7392 7404 7420 7500
rect 7742 7488 7748 7500
rect 7800 7488 7806 7540
rect 8202 7488 8208 7540
rect 8260 7528 8266 7540
rect 9033 7531 9091 7537
rect 9033 7528 9045 7531
rect 8260 7500 9045 7528
rect 8260 7488 8266 7500
rect 9033 7497 9045 7500
rect 9079 7528 9091 7531
rect 10686 7528 10692 7540
rect 9079 7500 10692 7528
rect 9079 7497 9091 7500
rect 9033 7491 9091 7497
rect 10686 7488 10692 7500
rect 10744 7488 10750 7540
rect 10965 7531 11023 7537
rect 10965 7497 10977 7531
rect 11011 7528 11023 7531
rect 15378 7528 15384 7540
rect 11011 7500 15384 7528
rect 11011 7497 11023 7500
rect 10965 7491 11023 7497
rect 15378 7488 15384 7500
rect 15436 7488 15442 7540
rect 16942 7488 16948 7540
rect 17000 7528 17006 7540
rect 17678 7528 17684 7540
rect 17000 7500 17684 7528
rect 17000 7488 17006 7500
rect 17678 7488 17684 7500
rect 17736 7488 17742 7540
rect 18414 7488 18420 7540
rect 18472 7528 18478 7540
rect 24302 7528 24308 7540
rect 18472 7500 24308 7528
rect 18472 7488 18478 7500
rect 24302 7488 24308 7500
rect 24360 7488 24366 7540
rect 26234 7528 26240 7540
rect 25148 7500 26240 7528
rect 7558 7420 7564 7472
rect 7616 7460 7622 7472
rect 11517 7463 11575 7469
rect 11517 7460 11529 7463
rect 7616 7432 11529 7460
rect 7616 7420 7622 7432
rect 11517 7429 11529 7432
rect 11563 7429 11575 7463
rect 13998 7460 14004 7472
rect 11517 7423 11575 7429
rect 11624 7432 14004 7460
rect 6549 7395 6607 7401
rect 6549 7392 6561 7395
rect 6420 7364 6561 7392
rect 6420 7352 6426 7364
rect 6549 7361 6561 7364
rect 6595 7361 6607 7395
rect 6549 7355 6607 7361
rect 6641 7395 6699 7401
rect 6641 7361 6653 7395
rect 6687 7361 6699 7395
rect 7374 7392 7380 7404
rect 7287 7364 7380 7392
rect 6641 7355 6699 7361
rect 7374 7352 7380 7364
rect 7432 7352 7438 7404
rect 8297 7395 8355 7401
rect 8297 7392 8309 7395
rect 7484 7364 8309 7392
rect 4154 7324 4160 7336
rect 3252 7296 4160 7324
rect 2593 7287 2651 7293
rect 2608 7256 2636 7287
rect 4154 7284 4160 7296
rect 4212 7284 4218 7336
rect 5169 7327 5227 7333
rect 5169 7293 5181 7327
rect 5215 7324 5227 7327
rect 5810 7324 5816 7336
rect 5215 7296 5816 7324
rect 5215 7293 5227 7296
rect 5169 7287 5227 7293
rect 5810 7284 5816 7296
rect 5868 7284 5874 7336
rect 5994 7284 6000 7336
rect 6052 7324 6058 7336
rect 7484 7324 7512 7364
rect 8297 7361 8309 7364
rect 8343 7361 8355 7395
rect 8297 7355 8355 7361
rect 9677 7395 9735 7401
rect 9677 7361 9689 7395
rect 9723 7392 9735 7395
rect 10781 7395 10839 7401
rect 9723 7364 10732 7392
rect 9723 7361 9735 7364
rect 9677 7355 9735 7361
rect 6052 7296 7512 7324
rect 7561 7327 7619 7333
rect 6052 7284 6058 7296
rect 7561 7293 7573 7327
rect 7607 7293 7619 7327
rect 8018 7324 8024 7336
rect 7979 7296 8024 7324
rect 7561 7287 7619 7293
rect 2958 7256 2964 7268
rect 2608 7228 2964 7256
rect 2958 7216 2964 7228
rect 3016 7216 3022 7268
rect 5442 7216 5448 7268
rect 5500 7256 5506 7268
rect 7193 7259 7251 7265
rect 7193 7256 7205 7259
rect 5500 7228 7205 7256
rect 5500 7216 5506 7228
rect 7193 7225 7205 7228
rect 7239 7225 7251 7259
rect 7193 7219 7251 7225
rect 2222 7188 2228 7200
rect 2183 7160 2228 7188
rect 2222 7148 2228 7160
rect 2280 7148 2286 7200
rect 3050 7188 3056 7200
rect 3011 7160 3056 7188
rect 3050 7148 3056 7160
rect 3108 7148 3114 7200
rect 4154 7188 4160 7200
rect 4115 7160 4160 7188
rect 4154 7148 4160 7160
rect 4212 7188 4218 7200
rect 5350 7188 5356 7200
rect 4212 7160 5356 7188
rect 4212 7148 4218 7160
rect 5350 7148 5356 7160
rect 5408 7148 5414 7200
rect 5813 7191 5871 7197
rect 5813 7157 5825 7191
rect 5859 7188 5871 7191
rect 6730 7188 6736 7200
rect 5859 7160 6736 7188
rect 5859 7157 5871 7160
rect 5813 7151 5871 7157
rect 6730 7148 6736 7160
rect 6788 7148 6794 7200
rect 6914 7148 6920 7200
rect 6972 7188 6978 7200
rect 7576 7188 7604 7287
rect 8018 7284 8024 7296
rect 8076 7284 8082 7336
rect 9490 7324 9496 7336
rect 9451 7296 9496 7324
rect 9490 7284 9496 7296
rect 9548 7284 9554 7336
rect 9861 7327 9919 7333
rect 9861 7293 9873 7327
rect 9907 7293 9919 7327
rect 10704 7324 10732 7364
rect 10781 7361 10793 7395
rect 10827 7392 10839 7395
rect 11624 7392 11652 7432
rect 13998 7420 14004 7432
rect 14056 7420 14062 7472
rect 19242 7460 19248 7472
rect 17236 7432 19248 7460
rect 10827 7364 11652 7392
rect 11701 7395 11759 7401
rect 10827 7361 10839 7364
rect 10781 7355 10839 7361
rect 11701 7361 11713 7395
rect 11747 7392 11759 7395
rect 12437 7395 12495 7401
rect 12437 7392 12449 7395
rect 11747 7364 12449 7392
rect 11747 7361 11759 7364
rect 11701 7355 11759 7361
rect 12437 7361 12449 7364
rect 12483 7361 12495 7395
rect 12437 7355 12495 7361
rect 11716 7324 11744 7355
rect 10704 7296 11744 7324
rect 9861 7287 9919 7293
rect 9876 7256 9904 7287
rect 11790 7284 11796 7336
rect 11848 7324 11854 7336
rect 11885 7327 11943 7333
rect 11885 7324 11897 7327
rect 11848 7296 11897 7324
rect 11848 7284 11854 7296
rect 11885 7293 11897 7296
rect 11931 7293 11943 7327
rect 12452 7324 12480 7355
rect 12986 7352 12992 7404
rect 13044 7392 13050 7404
rect 13081 7395 13139 7401
rect 13081 7392 13093 7395
rect 13044 7364 13093 7392
rect 13044 7352 13050 7364
rect 13081 7361 13093 7364
rect 13127 7361 13139 7395
rect 13081 7355 13139 7361
rect 13814 7352 13820 7404
rect 13872 7392 13878 7404
rect 13909 7395 13967 7401
rect 13909 7392 13921 7395
rect 13872 7364 13921 7392
rect 13872 7352 13878 7364
rect 13909 7361 13921 7364
rect 13955 7361 13967 7395
rect 14090 7392 14096 7404
rect 14051 7364 14096 7392
rect 13909 7355 13967 7361
rect 14090 7352 14096 7364
rect 14148 7352 14154 7404
rect 14182 7352 14188 7404
rect 14240 7392 14246 7404
rect 15378 7392 15384 7404
rect 14240 7364 14285 7392
rect 15339 7364 15384 7392
rect 14240 7352 14246 7364
rect 15378 7352 15384 7364
rect 15436 7352 15442 7404
rect 16206 7352 16212 7404
rect 16264 7392 16270 7404
rect 17034 7392 17040 7404
rect 16264 7364 17040 7392
rect 16264 7352 16270 7364
rect 17034 7352 17040 7364
rect 17092 7352 17098 7404
rect 17236 7401 17264 7432
rect 19242 7420 19248 7432
rect 19300 7420 19306 7472
rect 24397 7463 24455 7469
rect 24397 7460 24409 7463
rect 22112 7432 24409 7460
rect 17221 7395 17279 7401
rect 17221 7361 17233 7395
rect 17267 7361 17279 7395
rect 17221 7355 17279 7361
rect 17865 7395 17923 7401
rect 17865 7361 17877 7395
rect 17911 7392 17923 7395
rect 17954 7392 17960 7404
rect 17911 7364 17960 7392
rect 17911 7361 17923 7364
rect 17865 7355 17923 7361
rect 17954 7352 17960 7364
rect 18012 7352 18018 7404
rect 18322 7392 18328 7404
rect 18283 7364 18328 7392
rect 18322 7352 18328 7364
rect 18380 7352 18386 7404
rect 18414 7352 18420 7404
rect 18472 7392 18478 7404
rect 19426 7392 19432 7404
rect 18472 7364 19432 7392
rect 18472 7352 18478 7364
rect 19426 7352 19432 7364
rect 19484 7352 19490 7404
rect 19610 7392 19616 7404
rect 19571 7364 19616 7392
rect 19610 7352 19616 7364
rect 19668 7352 19674 7404
rect 19702 7352 19708 7404
rect 19760 7392 19766 7404
rect 21085 7395 21143 7401
rect 21085 7392 21097 7395
rect 19760 7364 21097 7392
rect 19760 7352 19766 7364
rect 21085 7361 21097 7364
rect 21131 7361 21143 7395
rect 21085 7355 21143 7361
rect 21269 7395 21327 7401
rect 21269 7361 21281 7395
rect 21315 7392 21327 7395
rect 21450 7392 21456 7404
rect 21315 7364 21456 7392
rect 21315 7361 21327 7364
rect 21269 7355 21327 7361
rect 21450 7352 21456 7364
rect 21508 7352 21514 7404
rect 22112 7401 22140 7432
rect 24397 7429 24409 7432
rect 24443 7460 24455 7463
rect 24578 7460 24584 7472
rect 24443 7432 24584 7460
rect 24443 7429 24455 7432
rect 24397 7423 24455 7429
rect 24578 7420 24584 7432
rect 24636 7420 24642 7472
rect 22097 7395 22155 7401
rect 22097 7361 22109 7395
rect 22143 7361 22155 7395
rect 22833 7395 22891 7401
rect 22833 7392 22845 7395
rect 22097 7355 22155 7361
rect 22480 7364 22845 7392
rect 14108 7324 14136 7352
rect 12452 7296 14136 7324
rect 11885 7287 11943 7293
rect 14918 7284 14924 7336
rect 14976 7324 14982 7336
rect 15105 7327 15163 7333
rect 15105 7324 15117 7327
rect 14976 7296 15117 7324
rect 14976 7284 14982 7296
rect 15105 7293 15117 7296
rect 15151 7293 15163 7327
rect 15105 7287 15163 7293
rect 18966 7284 18972 7336
rect 19024 7324 19030 7336
rect 19889 7327 19947 7333
rect 19889 7324 19901 7327
rect 19024 7296 19901 7324
rect 19024 7284 19030 7296
rect 19889 7293 19901 7296
rect 19935 7293 19947 7327
rect 19889 7287 19947 7293
rect 21818 7284 21824 7336
rect 21876 7324 21882 7336
rect 22480 7324 22508 7364
rect 22833 7361 22845 7364
rect 22879 7361 22891 7395
rect 24302 7392 24308 7404
rect 24263 7364 24308 7392
rect 22833 7355 22891 7361
rect 24302 7352 24308 7364
rect 24360 7352 24366 7404
rect 24489 7395 24547 7401
rect 24489 7361 24501 7395
rect 24535 7392 24547 7395
rect 25148 7392 25176 7500
rect 26234 7488 26240 7500
rect 26292 7488 26298 7540
rect 31573 7531 31631 7537
rect 31573 7497 31585 7531
rect 31619 7528 31631 7531
rect 34149 7531 34207 7537
rect 31619 7500 31754 7528
rect 31619 7497 31631 7500
rect 31573 7491 31631 7497
rect 31726 7460 31754 7500
rect 34149 7497 34161 7531
rect 34195 7528 34207 7531
rect 34974 7528 34980 7540
rect 34195 7500 34980 7528
rect 34195 7497 34207 7500
rect 34149 7491 34207 7497
rect 34974 7488 34980 7500
rect 35032 7488 35038 7540
rect 42426 7528 42432 7540
rect 38304 7500 42432 7528
rect 35986 7460 35992 7472
rect 25700 7432 28764 7460
rect 31726 7432 32720 7460
rect 24535 7364 25176 7392
rect 24535 7361 24547 7364
rect 24489 7355 24547 7361
rect 25222 7352 25228 7404
rect 25280 7392 25286 7404
rect 25700 7401 25728 7432
rect 25685 7395 25743 7401
rect 25685 7392 25697 7395
rect 25280 7364 25697 7392
rect 25280 7352 25286 7364
rect 25685 7361 25697 7364
rect 25731 7361 25743 7395
rect 26050 7392 26056 7404
rect 26011 7364 26056 7392
rect 25685 7355 25743 7361
rect 26050 7352 26056 7364
rect 26108 7352 26114 7404
rect 26234 7352 26240 7404
rect 26292 7392 26298 7404
rect 26421 7395 26479 7401
rect 26421 7392 26433 7395
rect 26292 7364 26433 7392
rect 26292 7352 26298 7364
rect 26421 7361 26433 7364
rect 26467 7392 26479 7395
rect 26878 7392 26884 7404
rect 26467 7364 26884 7392
rect 26467 7361 26479 7364
rect 26421 7355 26479 7361
rect 26878 7352 26884 7364
rect 26936 7352 26942 7404
rect 21876 7296 22508 7324
rect 22557 7327 22615 7333
rect 21876 7284 21882 7296
rect 22557 7293 22569 7327
rect 22603 7293 22615 7327
rect 25038 7324 25044 7336
rect 24999 7296 25044 7324
rect 22557 7287 22615 7293
rect 9508 7228 9904 7256
rect 9508 7188 9536 7228
rect 12066 7216 12072 7268
rect 12124 7256 12130 7268
rect 13265 7259 13323 7265
rect 13265 7256 13277 7259
rect 12124 7228 13277 7256
rect 12124 7216 12130 7228
rect 13265 7225 13277 7228
rect 13311 7225 13323 7259
rect 13265 7219 13323 7225
rect 13722 7216 13728 7268
rect 13780 7256 13786 7268
rect 13780 7228 14044 7256
rect 13780 7216 13786 7228
rect 12526 7188 12532 7200
rect 6972 7160 9536 7188
rect 12487 7160 12532 7188
rect 6972 7148 6978 7160
rect 12526 7148 12532 7160
rect 12584 7188 12590 7200
rect 12894 7188 12900 7200
rect 12584 7160 12900 7188
rect 12584 7148 12590 7160
rect 12894 7148 12900 7160
rect 12952 7148 12958 7200
rect 14016 7188 14044 7228
rect 15672 7228 22094 7256
rect 15672 7188 15700 7228
rect 14016 7160 15700 7188
rect 16117 7191 16175 7197
rect 16117 7157 16129 7191
rect 16163 7188 16175 7191
rect 16298 7188 16304 7200
rect 16163 7160 16304 7188
rect 16163 7157 16175 7160
rect 16117 7151 16175 7157
rect 16298 7148 16304 7160
rect 16356 7148 16362 7200
rect 16390 7148 16396 7200
rect 16448 7188 16454 7200
rect 17037 7191 17095 7197
rect 17037 7188 17049 7191
rect 16448 7160 17049 7188
rect 16448 7148 16454 7160
rect 17037 7157 17049 7160
rect 17083 7188 17095 7191
rect 18414 7188 18420 7200
rect 17083 7160 18420 7188
rect 17083 7157 17095 7160
rect 17037 7151 17095 7157
rect 18414 7148 18420 7160
rect 18472 7148 18478 7200
rect 18509 7191 18567 7197
rect 18509 7157 18521 7191
rect 18555 7188 18567 7191
rect 19058 7188 19064 7200
rect 18555 7160 19064 7188
rect 18555 7157 18567 7160
rect 18509 7151 18567 7157
rect 19058 7148 19064 7160
rect 19116 7148 19122 7200
rect 19150 7148 19156 7200
rect 19208 7188 19214 7200
rect 19208 7160 19253 7188
rect 19208 7148 19214 7160
rect 19610 7148 19616 7200
rect 19668 7188 19674 7200
rect 20901 7191 20959 7197
rect 20901 7188 20913 7191
rect 19668 7160 20913 7188
rect 19668 7148 19674 7160
rect 20901 7157 20913 7160
rect 20947 7157 20959 7191
rect 21910 7188 21916 7200
rect 21871 7160 21916 7188
rect 20901 7151 20959 7157
rect 21910 7148 21916 7160
rect 21968 7148 21974 7200
rect 22066 7188 22094 7228
rect 22278 7216 22284 7268
rect 22336 7256 22342 7268
rect 22572 7256 22600 7287
rect 25038 7284 25044 7296
rect 25096 7284 25102 7336
rect 25130 7284 25136 7336
rect 25188 7324 25194 7336
rect 25188 7296 25233 7324
rect 25188 7284 25194 7296
rect 26786 7284 26792 7336
rect 26844 7324 26850 7336
rect 26973 7327 27031 7333
rect 26973 7324 26985 7327
rect 26844 7296 26985 7324
rect 26844 7284 26850 7296
rect 26973 7293 26985 7296
rect 27019 7293 27031 7327
rect 26973 7287 27031 7293
rect 27249 7327 27307 7333
rect 27249 7293 27261 7327
rect 27295 7293 27307 7327
rect 27249 7287 27307 7293
rect 27264 7256 27292 7287
rect 28350 7284 28356 7336
rect 28408 7324 28414 7336
rect 28736 7333 28764 7432
rect 28994 7392 29000 7404
rect 28955 7364 29000 7392
rect 28994 7352 29000 7364
rect 29052 7352 29058 7404
rect 29638 7352 29644 7404
rect 29696 7392 29702 7404
rect 30193 7395 30251 7401
rect 30193 7392 30205 7395
rect 29696 7364 30205 7392
rect 29696 7352 29702 7364
rect 30193 7361 30205 7364
rect 30239 7361 30251 7395
rect 30193 7355 30251 7361
rect 31389 7395 31447 7401
rect 31389 7361 31401 7395
rect 31435 7392 31447 7395
rect 31846 7392 31852 7404
rect 31435 7364 31852 7392
rect 31435 7361 31447 7364
rect 31389 7355 31447 7361
rect 28629 7327 28687 7333
rect 28629 7324 28641 7327
rect 28408 7296 28641 7324
rect 28408 7284 28414 7296
rect 28629 7293 28641 7296
rect 28675 7293 28687 7327
rect 28629 7287 28687 7293
rect 28721 7327 28779 7333
rect 28721 7293 28733 7327
rect 28767 7324 28779 7327
rect 29822 7324 29828 7336
rect 28767 7296 29828 7324
rect 28767 7293 28779 7296
rect 28721 7287 28779 7293
rect 29822 7284 29828 7296
rect 29880 7284 29886 7336
rect 29917 7327 29975 7333
rect 29917 7293 29929 7327
rect 29963 7293 29975 7327
rect 29917 7287 29975 7293
rect 29730 7256 29736 7268
rect 22336 7228 22600 7256
rect 23216 7228 29736 7256
rect 22336 7216 22342 7228
rect 23216 7188 23244 7228
rect 29730 7216 29736 7228
rect 29788 7216 29794 7268
rect 29932 7256 29960 7287
rect 29840 7228 29960 7256
rect 30208 7256 30236 7355
rect 31846 7352 31852 7364
rect 31904 7352 31910 7404
rect 32692 7401 32720 7432
rect 34624 7432 35992 7460
rect 34624 7404 34652 7432
rect 35986 7420 35992 7432
rect 36044 7420 36050 7472
rect 36354 7420 36360 7472
rect 36412 7460 36418 7472
rect 38304 7469 38332 7500
rect 42426 7488 42432 7500
rect 42484 7488 42490 7540
rect 46014 7528 46020 7540
rect 45975 7500 46020 7528
rect 46014 7488 46020 7500
rect 46072 7488 46078 7540
rect 51166 7488 51172 7540
rect 51224 7528 51230 7540
rect 51353 7531 51411 7537
rect 51353 7528 51365 7531
rect 51224 7500 51365 7528
rect 51224 7488 51230 7500
rect 51353 7497 51365 7500
rect 51399 7497 51411 7531
rect 51353 7491 51411 7497
rect 51442 7488 51448 7540
rect 51500 7528 51506 7540
rect 51997 7531 52055 7537
rect 51997 7528 52009 7531
rect 51500 7500 52009 7528
rect 51500 7488 51506 7500
rect 51997 7497 52009 7500
rect 52043 7497 52055 7531
rect 53098 7528 53104 7540
rect 53059 7500 53104 7528
rect 51997 7491 52055 7497
rect 53098 7488 53104 7500
rect 53156 7488 53162 7540
rect 38289 7463 38347 7469
rect 38289 7460 38301 7463
rect 36412 7432 38301 7460
rect 36412 7420 36418 7432
rect 38289 7429 38301 7432
rect 38335 7429 38347 7463
rect 38289 7423 38347 7429
rect 38930 7420 38936 7472
rect 38988 7460 38994 7472
rect 40586 7460 40592 7472
rect 38988 7432 40592 7460
rect 38988 7420 38994 7432
rect 32677 7395 32735 7401
rect 32677 7361 32689 7395
rect 32723 7361 32735 7395
rect 33962 7392 33968 7404
rect 33923 7364 33968 7392
rect 32677 7355 32735 7361
rect 33962 7352 33968 7364
rect 34020 7352 34026 7404
rect 34606 7392 34612 7404
rect 34567 7364 34612 7392
rect 34606 7352 34612 7364
rect 34664 7352 34670 7404
rect 34698 7352 34704 7404
rect 34756 7392 34762 7404
rect 35529 7395 35587 7401
rect 35529 7392 35541 7395
rect 34756 7364 35541 7392
rect 34756 7352 34762 7364
rect 35529 7361 35541 7364
rect 35575 7361 35587 7395
rect 37458 7392 37464 7404
rect 37419 7364 37464 7392
rect 35529 7355 35587 7361
rect 37458 7352 37464 7364
rect 37516 7352 37522 7404
rect 37550 7352 37556 7404
rect 37608 7392 37614 7404
rect 37608 7364 37653 7392
rect 37608 7352 37614 7364
rect 38654 7352 38660 7404
rect 38712 7392 38718 7404
rect 40420 7401 40448 7432
rect 40586 7420 40592 7432
rect 40644 7420 40650 7472
rect 43990 7460 43996 7472
rect 43548 7432 43996 7460
rect 39209 7395 39267 7401
rect 39209 7392 39221 7395
rect 38712 7364 39221 7392
rect 38712 7352 38718 7364
rect 39209 7361 39221 7364
rect 39255 7361 39267 7395
rect 39209 7355 39267 7361
rect 40405 7395 40463 7401
rect 40405 7361 40417 7395
rect 40451 7361 40463 7395
rect 40678 7392 40684 7404
rect 40639 7364 40684 7392
rect 40405 7355 40463 7361
rect 40678 7352 40684 7364
rect 40736 7352 40742 7404
rect 42797 7395 42855 7401
rect 42797 7361 42809 7395
rect 42843 7392 42855 7395
rect 42886 7392 42892 7404
rect 42843 7364 42892 7392
rect 42843 7361 42855 7364
rect 42797 7355 42855 7361
rect 42886 7352 42892 7364
rect 42944 7352 42950 7404
rect 43548 7401 43576 7432
rect 43990 7420 43996 7432
rect 44048 7420 44054 7472
rect 44637 7463 44695 7469
rect 44637 7429 44649 7463
rect 44683 7460 44695 7463
rect 44683 7432 46704 7460
rect 44683 7429 44695 7432
rect 44637 7423 44695 7429
rect 43533 7395 43591 7401
rect 43533 7361 43545 7395
rect 43579 7361 43591 7395
rect 43533 7355 43591 7361
rect 43625 7395 43683 7401
rect 43625 7361 43637 7395
rect 43671 7392 43683 7395
rect 44453 7395 44511 7401
rect 44453 7392 44465 7395
rect 43671 7364 44465 7392
rect 43671 7361 43683 7364
rect 43625 7355 43683 7361
rect 44453 7361 44465 7364
rect 44499 7392 44511 7395
rect 44499 7364 45324 7392
rect 44499 7361 44511 7364
rect 44453 7355 44511 7361
rect 31570 7284 31576 7336
rect 31628 7324 31634 7336
rect 32401 7327 32459 7333
rect 32401 7324 32413 7327
rect 31628 7296 32413 7324
rect 31628 7284 31634 7296
rect 32401 7293 32413 7296
rect 32447 7293 32459 7327
rect 35250 7324 35256 7336
rect 35211 7296 35256 7324
rect 32401 7287 32459 7293
rect 32306 7256 32312 7268
rect 30208 7228 32312 7256
rect 22066 7160 23244 7188
rect 23290 7148 23296 7200
rect 23348 7188 23354 7200
rect 23569 7191 23627 7197
rect 23569 7188 23581 7191
rect 23348 7160 23581 7188
rect 23348 7148 23354 7160
rect 23569 7157 23581 7160
rect 23615 7157 23627 7191
rect 23569 7151 23627 7157
rect 23934 7148 23940 7200
rect 23992 7188 23998 7200
rect 26326 7188 26332 7200
rect 23992 7160 26332 7188
rect 23992 7148 23998 7160
rect 26326 7148 26332 7160
rect 26384 7148 26390 7200
rect 27246 7148 27252 7200
rect 27304 7188 27310 7200
rect 29840 7188 29868 7228
rect 32306 7216 32312 7228
rect 32364 7216 32370 7268
rect 31294 7188 31300 7200
rect 27304 7160 31300 7188
rect 27304 7148 27310 7160
rect 31294 7148 31300 7160
rect 31352 7148 31358 7200
rect 32416 7188 32444 7287
rect 35250 7284 35256 7296
rect 35308 7284 35314 7336
rect 36814 7284 36820 7336
rect 36872 7324 36878 7336
rect 37918 7324 37924 7336
rect 36872 7296 37924 7324
rect 36872 7284 36878 7296
rect 37918 7284 37924 7296
rect 37976 7284 37982 7336
rect 38930 7324 38936 7336
rect 38891 7296 38936 7324
rect 38930 7284 38936 7296
rect 38988 7284 38994 7336
rect 35268 7256 35296 7284
rect 32968 7228 35296 7256
rect 32968 7188 32996 7228
rect 36630 7216 36636 7268
rect 36688 7256 36694 7268
rect 37734 7256 37740 7268
rect 36688 7228 37740 7256
rect 36688 7216 36694 7228
rect 37734 7216 37740 7228
rect 37792 7216 37798 7268
rect 38102 7256 38108 7268
rect 38063 7228 38108 7256
rect 38102 7216 38108 7228
rect 38160 7216 38166 7268
rect 41414 7256 41420 7268
rect 41386 7216 41420 7256
rect 41472 7256 41478 7268
rect 42981 7259 43039 7265
rect 41472 7228 41517 7256
rect 41472 7216 41478 7228
rect 42981 7225 42993 7259
rect 43027 7256 43039 7259
rect 43640 7256 43668 7355
rect 44269 7327 44327 7333
rect 44269 7293 44281 7327
rect 44315 7324 44327 7327
rect 44634 7324 44640 7336
rect 44315 7296 44640 7324
rect 44315 7293 44327 7296
rect 44269 7287 44327 7293
rect 44634 7284 44640 7296
rect 44692 7284 44698 7336
rect 45002 7284 45008 7336
rect 45060 7324 45066 7336
rect 45189 7327 45247 7333
rect 45189 7324 45201 7327
rect 45060 7296 45201 7324
rect 45060 7284 45066 7296
rect 45189 7293 45201 7296
rect 45235 7293 45247 7327
rect 45296 7324 45324 7364
rect 45370 7352 45376 7404
rect 45428 7392 45434 7404
rect 46676 7401 46704 7432
rect 49344 7432 52960 7460
rect 49344 7401 49372 7432
rect 45557 7395 45615 7401
rect 45428 7364 45473 7392
rect 45428 7352 45434 7364
rect 45557 7361 45569 7395
rect 45603 7392 45615 7395
rect 46201 7395 46259 7401
rect 46201 7392 46213 7395
rect 45603 7364 46213 7392
rect 45603 7361 45615 7364
rect 45557 7355 45615 7361
rect 46201 7361 46213 7364
rect 46247 7361 46259 7395
rect 46201 7355 46259 7361
rect 46661 7395 46719 7401
rect 46661 7361 46673 7395
rect 46707 7361 46719 7395
rect 48225 7395 48283 7401
rect 48225 7392 48237 7395
rect 46661 7355 46719 7361
rect 46768 7364 48237 7392
rect 46768 7324 46796 7364
rect 48225 7361 48237 7364
rect 48271 7392 48283 7395
rect 49329 7395 49387 7401
rect 49329 7392 49341 7395
rect 48271 7364 49341 7392
rect 48271 7361 48283 7364
rect 48225 7355 48283 7361
rect 49329 7361 49341 7364
rect 49375 7361 49387 7395
rect 50338 7392 50344 7404
rect 50299 7364 50344 7392
rect 49329 7355 49387 7361
rect 50338 7352 50344 7364
rect 50396 7352 50402 7404
rect 50614 7392 50620 7404
rect 50575 7364 50620 7392
rect 50614 7352 50620 7364
rect 50672 7352 50678 7404
rect 52086 7392 52092 7404
rect 51999 7364 52092 7392
rect 52086 7352 52092 7364
rect 52144 7352 52150 7404
rect 52932 7401 52960 7432
rect 55858 7420 55864 7472
rect 55916 7460 55922 7472
rect 55916 7432 56548 7460
rect 55916 7420 55922 7432
rect 52917 7395 52975 7401
rect 52917 7361 52929 7395
rect 52963 7361 52975 7395
rect 54202 7392 54208 7404
rect 54163 7364 54208 7392
rect 52917 7355 52975 7361
rect 54202 7352 54208 7364
rect 54260 7352 54266 7404
rect 55677 7395 55735 7401
rect 55677 7361 55689 7395
rect 55723 7392 55735 7395
rect 56226 7392 56232 7404
rect 55723 7364 56232 7392
rect 55723 7361 55735 7364
rect 55677 7355 55735 7361
rect 56226 7352 56232 7364
rect 56284 7352 56290 7404
rect 56520 7401 56548 7432
rect 56321 7395 56379 7401
rect 56321 7361 56333 7395
rect 56367 7361 56379 7395
rect 56321 7355 56379 7361
rect 56505 7395 56563 7401
rect 56505 7361 56517 7395
rect 56551 7361 56563 7395
rect 56505 7355 56563 7361
rect 57885 7395 57943 7401
rect 57885 7361 57897 7395
rect 57931 7361 57943 7395
rect 57885 7355 57943 7361
rect 48038 7324 48044 7336
rect 45296 7296 46796 7324
rect 47951 7296 48044 7324
rect 45189 7287 45247 7293
rect 48038 7284 48044 7296
rect 48096 7284 48102 7336
rect 49145 7327 49203 7333
rect 49145 7293 49157 7327
rect 49191 7324 49203 7327
rect 49234 7324 49240 7336
rect 49191 7296 49240 7324
rect 49191 7293 49203 7296
rect 49145 7287 49203 7293
rect 49234 7284 49240 7296
rect 49292 7284 49298 7336
rect 52104 7324 52132 7352
rect 52362 7324 52368 7336
rect 52104 7296 52368 7324
rect 52362 7284 52368 7296
rect 52420 7324 52426 7336
rect 52733 7327 52791 7333
rect 52733 7324 52745 7327
rect 52420 7296 52745 7324
rect 52420 7284 52426 7296
rect 52733 7293 52745 7296
rect 52779 7293 52791 7327
rect 52733 7287 52791 7293
rect 52822 7284 52828 7336
rect 52880 7324 52886 7336
rect 53929 7327 53987 7333
rect 53929 7324 53941 7327
rect 52880 7296 53941 7324
rect 52880 7284 52886 7296
rect 53929 7293 53941 7296
rect 53975 7293 53987 7327
rect 53929 7287 53987 7293
rect 55582 7284 55588 7336
rect 55640 7324 55646 7336
rect 56336 7324 56364 7355
rect 55640 7296 56364 7324
rect 56413 7327 56471 7333
rect 55640 7284 55646 7296
rect 56413 7293 56425 7327
rect 56459 7324 56471 7327
rect 57514 7324 57520 7336
rect 56459 7296 57520 7324
rect 56459 7293 56471 7296
rect 56413 7287 56471 7293
rect 57514 7284 57520 7296
rect 57572 7324 57578 7336
rect 57900 7324 57928 7355
rect 57572 7296 57928 7324
rect 57572 7284 57578 7296
rect 48056 7256 48084 7284
rect 43027 7228 43668 7256
rect 43732 7228 48084 7256
rect 48409 7259 48467 7265
rect 43027 7225 43039 7228
rect 42981 7219 43039 7225
rect 32416 7160 32996 7188
rect 33413 7191 33471 7197
rect 33413 7157 33425 7191
rect 33459 7188 33471 7191
rect 33594 7188 33600 7200
rect 33459 7160 33600 7188
rect 33459 7157 33471 7160
rect 33413 7151 33471 7157
rect 33594 7148 33600 7160
rect 33652 7148 33658 7200
rect 34701 7191 34759 7197
rect 34701 7157 34713 7191
rect 34747 7188 34759 7191
rect 34882 7188 34888 7200
rect 34747 7160 34888 7188
rect 34747 7157 34759 7160
rect 34701 7151 34759 7157
rect 34882 7148 34888 7160
rect 34940 7188 34946 7200
rect 35894 7188 35900 7200
rect 34940 7160 35900 7188
rect 34940 7148 34946 7160
rect 35894 7148 35900 7160
rect 35952 7148 35958 7200
rect 36170 7148 36176 7200
rect 36228 7188 36234 7200
rect 36265 7191 36323 7197
rect 36265 7188 36277 7191
rect 36228 7160 36277 7188
rect 36228 7148 36234 7160
rect 36265 7157 36277 7160
rect 36311 7188 36323 7191
rect 36906 7188 36912 7200
rect 36311 7160 36912 7188
rect 36311 7157 36323 7160
rect 36265 7151 36323 7157
rect 36906 7148 36912 7160
rect 36964 7148 36970 7200
rect 37277 7191 37335 7197
rect 37277 7157 37289 7191
rect 37323 7188 37335 7191
rect 37458 7188 37464 7200
rect 37323 7160 37464 7188
rect 37323 7157 37335 7160
rect 37277 7151 37335 7157
rect 37458 7148 37464 7160
rect 37516 7148 37522 7200
rect 38746 7148 38752 7200
rect 38804 7188 38810 7200
rect 39945 7191 40003 7197
rect 39945 7188 39957 7191
rect 38804 7160 39957 7188
rect 38804 7148 38810 7160
rect 39945 7157 39957 7160
rect 39991 7188 40003 7191
rect 41386 7188 41414 7216
rect 39991 7160 41414 7188
rect 39991 7157 40003 7160
rect 39945 7151 40003 7157
rect 42886 7148 42892 7200
rect 42944 7188 42950 7200
rect 43732 7188 43760 7228
rect 48409 7225 48421 7259
rect 48455 7256 48467 7259
rect 50062 7256 50068 7268
rect 48455 7228 50068 7256
rect 48455 7225 48467 7228
rect 48409 7219 48467 7225
rect 50062 7216 50068 7228
rect 50120 7216 50126 7268
rect 42944 7160 43760 7188
rect 43809 7191 43867 7197
rect 42944 7148 42950 7160
rect 43809 7157 43821 7191
rect 43855 7188 43867 7191
rect 44174 7188 44180 7200
rect 43855 7160 44180 7188
rect 43855 7157 43867 7160
rect 43809 7151 43867 7157
rect 44174 7148 44180 7160
rect 44232 7148 44238 7200
rect 46842 7188 46848 7200
rect 46803 7160 46848 7188
rect 46842 7148 46848 7160
rect 46900 7148 46906 7200
rect 49513 7191 49571 7197
rect 49513 7157 49525 7191
rect 49559 7188 49571 7191
rect 50706 7188 50712 7200
rect 49559 7160 50712 7188
rect 49559 7157 49571 7160
rect 49513 7151 49571 7157
rect 50706 7148 50712 7160
rect 50764 7148 50770 7200
rect 51258 7148 51264 7200
rect 51316 7188 51322 7200
rect 54941 7191 54999 7197
rect 54941 7188 54953 7191
rect 51316 7160 54953 7188
rect 51316 7148 51322 7160
rect 54941 7157 54953 7160
rect 54987 7157 54999 7191
rect 54941 7151 54999 7157
rect 55861 7191 55919 7197
rect 55861 7157 55873 7191
rect 55907 7188 55919 7191
rect 57790 7188 57796 7200
rect 55907 7160 57796 7188
rect 55907 7157 55919 7160
rect 55861 7151 55919 7157
rect 57790 7148 57796 7160
rect 57848 7148 57854 7200
rect 57974 7188 57980 7200
rect 57935 7160 57980 7188
rect 57974 7148 57980 7160
rect 58032 7148 58038 7200
rect 1104 7098 58880 7120
rect 1104 7046 8174 7098
rect 8226 7046 8238 7098
rect 8290 7046 8302 7098
rect 8354 7046 8366 7098
rect 8418 7046 8430 7098
rect 8482 7046 22622 7098
rect 22674 7046 22686 7098
rect 22738 7046 22750 7098
rect 22802 7046 22814 7098
rect 22866 7046 22878 7098
rect 22930 7046 37070 7098
rect 37122 7046 37134 7098
rect 37186 7046 37198 7098
rect 37250 7046 37262 7098
rect 37314 7046 37326 7098
rect 37378 7046 51518 7098
rect 51570 7046 51582 7098
rect 51634 7046 51646 7098
rect 51698 7046 51710 7098
rect 51762 7046 51774 7098
rect 51826 7046 58880 7098
rect 1104 7024 58880 7046
rect 5629 6987 5687 6993
rect 5629 6953 5641 6987
rect 5675 6984 5687 6987
rect 5810 6984 5816 6996
rect 5675 6956 5816 6984
rect 5675 6953 5687 6956
rect 5629 6947 5687 6953
rect 5810 6944 5816 6956
rect 5868 6944 5874 6996
rect 6089 6987 6147 6993
rect 6089 6953 6101 6987
rect 6135 6984 6147 6987
rect 6178 6984 6184 6996
rect 6135 6956 6184 6984
rect 6135 6953 6147 6956
rect 6089 6947 6147 6953
rect 6178 6944 6184 6956
rect 6236 6984 6242 6996
rect 7374 6984 7380 6996
rect 6236 6956 7380 6984
rect 6236 6944 6242 6956
rect 7374 6944 7380 6956
rect 7432 6944 7438 6996
rect 10594 6944 10600 6996
rect 10652 6984 10658 6996
rect 10652 6956 11744 6984
rect 10652 6944 10658 6956
rect 1949 6919 2007 6925
rect 1949 6885 1961 6919
rect 1995 6914 2007 6919
rect 1995 6886 2029 6914
rect 1995 6885 2007 6886
rect 1949 6879 2007 6885
rect 1964 6848 1992 6879
rect 4706 6876 4712 6928
rect 4764 6916 4770 6928
rect 5350 6916 5356 6928
rect 4764 6888 5356 6916
rect 4764 6876 4770 6888
rect 5350 6876 5356 6888
rect 5408 6916 5414 6928
rect 8018 6916 8024 6928
rect 5408 6888 8024 6916
rect 5408 6876 5414 6888
rect 8018 6876 8024 6888
rect 8076 6876 8082 6928
rect 3694 6848 3700 6860
rect 1964 6820 3700 6848
rect 3694 6808 3700 6820
rect 3752 6808 3758 6860
rect 10870 6808 10876 6860
rect 10928 6848 10934 6860
rect 11057 6851 11115 6857
rect 11057 6848 11069 6851
rect 10928 6820 11069 6848
rect 10928 6808 10934 6820
rect 11057 6817 11069 6820
rect 11103 6817 11115 6851
rect 11716 6848 11744 6956
rect 11790 6944 11796 6996
rect 11848 6984 11854 6996
rect 13722 6984 13728 6996
rect 11848 6956 13728 6984
rect 11848 6944 11854 6956
rect 13722 6944 13728 6956
rect 13780 6944 13786 6996
rect 16298 6944 16304 6996
rect 16356 6984 16362 6996
rect 17957 6987 18015 6993
rect 17957 6984 17969 6987
rect 16356 6956 17969 6984
rect 16356 6944 16362 6956
rect 17957 6953 17969 6956
rect 18003 6984 18015 6987
rect 18414 6984 18420 6996
rect 18003 6956 18420 6984
rect 18003 6953 18015 6956
rect 17957 6947 18015 6953
rect 18414 6944 18420 6956
rect 18472 6944 18478 6996
rect 21818 6984 21824 6996
rect 21779 6956 21824 6984
rect 21818 6944 21824 6956
rect 21876 6944 21882 6996
rect 23290 6984 23296 6996
rect 23251 6956 23296 6984
rect 23290 6944 23296 6956
rect 23348 6944 23354 6996
rect 24026 6944 24032 6996
rect 24084 6984 24090 6996
rect 24394 6984 24400 6996
rect 24084 6956 24400 6984
rect 24084 6944 24090 6956
rect 24394 6944 24400 6956
rect 24452 6944 24458 6996
rect 28810 6984 28816 6996
rect 25884 6956 28816 6984
rect 14366 6876 14372 6928
rect 14424 6916 14430 6928
rect 15657 6919 15715 6925
rect 15657 6916 15669 6919
rect 14424 6888 15669 6916
rect 14424 6876 14430 6888
rect 15657 6885 15669 6888
rect 15703 6916 15715 6919
rect 16390 6916 16396 6928
rect 15703 6888 16396 6916
rect 15703 6885 15715 6888
rect 15657 6879 15715 6885
rect 16390 6876 16396 6888
rect 16448 6876 16454 6928
rect 23845 6919 23903 6925
rect 23845 6885 23857 6919
rect 23891 6916 23903 6919
rect 25884 6916 25912 6956
rect 28810 6944 28816 6956
rect 28868 6944 28874 6996
rect 29730 6984 29736 6996
rect 29691 6956 29736 6984
rect 29730 6944 29736 6956
rect 29788 6944 29794 6996
rect 30561 6987 30619 6993
rect 30561 6953 30573 6987
rect 30607 6984 30619 6987
rect 33410 6984 33416 6996
rect 30607 6956 33416 6984
rect 30607 6953 30619 6956
rect 30561 6947 30619 6953
rect 26050 6916 26056 6928
rect 23891 6888 25912 6916
rect 25963 6888 26056 6916
rect 23891 6885 23903 6888
rect 23845 6879 23903 6885
rect 11716 6820 12940 6848
rect 11057 6811 11115 6817
rect 1765 6783 1823 6789
rect 1765 6749 1777 6783
rect 1811 6780 1823 6783
rect 2130 6780 2136 6792
rect 1811 6752 2136 6780
rect 1811 6749 1823 6752
rect 1765 6743 1823 6749
rect 2130 6740 2136 6752
rect 2188 6740 2194 6792
rect 2409 6783 2467 6789
rect 2409 6749 2421 6783
rect 2455 6780 2467 6783
rect 3142 6780 3148 6792
rect 2455 6752 3148 6780
rect 2455 6749 2467 6752
rect 2409 6743 2467 6749
rect 3142 6740 3148 6752
rect 3200 6740 3206 6792
rect 3237 6783 3295 6789
rect 3237 6749 3249 6783
rect 3283 6780 3295 6783
rect 3510 6780 3516 6792
rect 3283 6752 3516 6780
rect 3283 6749 3295 6752
rect 3237 6743 3295 6749
rect 3510 6740 3516 6752
rect 3568 6740 3574 6792
rect 3789 6783 3847 6789
rect 3789 6749 3801 6783
rect 3835 6780 3847 6783
rect 3970 6780 3976 6792
rect 3835 6752 3976 6780
rect 3835 6749 3847 6752
rect 3789 6743 3847 6749
rect 3970 6740 3976 6752
rect 4028 6740 4034 6792
rect 4065 6783 4123 6789
rect 4065 6749 4077 6783
rect 4111 6749 4123 6783
rect 4065 6743 4123 6749
rect 1854 6672 1860 6724
rect 1912 6712 1918 6724
rect 4080 6712 4108 6743
rect 5350 6740 5356 6792
rect 5408 6780 5414 6792
rect 5445 6783 5503 6789
rect 5445 6780 5457 6783
rect 5408 6752 5457 6780
rect 5408 6740 5414 6752
rect 5445 6749 5457 6752
rect 5491 6749 5503 6783
rect 5445 6743 5503 6749
rect 6273 6783 6331 6789
rect 6273 6749 6285 6783
rect 6319 6780 6331 6783
rect 6546 6780 6552 6792
rect 6319 6752 6552 6780
rect 6319 6749 6331 6752
rect 6273 6743 6331 6749
rect 6546 6740 6552 6752
rect 6604 6740 6610 6792
rect 6730 6780 6736 6792
rect 6691 6752 6736 6780
rect 6730 6740 6736 6752
rect 6788 6740 6794 6792
rect 6917 6783 6975 6789
rect 6917 6749 6929 6783
rect 6963 6749 6975 6783
rect 6917 6743 6975 6749
rect 7009 6783 7067 6789
rect 7009 6749 7021 6783
rect 7055 6749 7067 6783
rect 7009 6743 7067 6749
rect 7101 6783 7159 6789
rect 7101 6749 7113 6783
rect 7147 6780 7159 6783
rect 7282 6780 7288 6792
rect 7147 6752 7288 6780
rect 7147 6749 7159 6752
rect 7101 6743 7159 6749
rect 6932 6712 6960 6743
rect 1912 6684 4108 6712
rect 4172 6684 6960 6712
rect 7024 6712 7052 6743
rect 7282 6740 7288 6752
rect 7340 6740 7346 6792
rect 7926 6740 7932 6792
rect 7984 6780 7990 6792
rect 8389 6783 8447 6789
rect 8389 6780 8401 6783
rect 7984 6752 8401 6780
rect 7984 6740 7990 6752
rect 8389 6749 8401 6752
rect 8435 6749 8447 6783
rect 9490 6780 9496 6792
rect 9451 6752 9496 6780
rect 8389 6743 8447 6749
rect 9490 6740 9496 6752
rect 9548 6740 9554 6792
rect 9674 6740 9680 6792
rect 9732 6780 9738 6792
rect 10137 6783 10195 6789
rect 10137 6780 10149 6783
rect 9732 6752 10149 6780
rect 9732 6740 9738 6752
rect 10137 6749 10149 6752
rect 10183 6780 10195 6783
rect 10183 6752 10456 6780
rect 10183 6749 10195 6752
rect 10137 6743 10195 6749
rect 10318 6712 10324 6724
rect 7024 6684 10180 6712
rect 10279 6684 10324 6712
rect 1912 6672 1918 6684
rect 2590 6644 2596 6656
rect 2551 6616 2596 6644
rect 2590 6604 2596 6616
rect 2648 6604 2654 6656
rect 3142 6604 3148 6656
rect 3200 6644 3206 6656
rect 4172 6644 4200 6684
rect 3200 6616 4200 6644
rect 3200 6604 3206 6616
rect 4706 6604 4712 6656
rect 4764 6644 4770 6656
rect 4801 6647 4859 6653
rect 4801 6644 4813 6647
rect 4764 6616 4813 6644
rect 4764 6604 4770 6616
rect 4801 6613 4813 6616
rect 4847 6613 4859 6647
rect 4801 6607 4859 6613
rect 5994 6604 6000 6656
rect 6052 6644 6058 6656
rect 7024 6644 7052 6684
rect 7374 6644 7380 6656
rect 6052 6616 7052 6644
rect 7335 6616 7380 6644
rect 6052 6604 6058 6616
rect 7374 6604 7380 6616
rect 7432 6604 7438 6656
rect 8018 6604 8024 6656
rect 8076 6644 8082 6656
rect 8205 6647 8263 6653
rect 8205 6644 8217 6647
rect 8076 6616 8217 6644
rect 8076 6604 8082 6616
rect 8205 6613 8217 6616
rect 8251 6613 8263 6647
rect 8205 6607 8263 6613
rect 8754 6604 8760 6656
rect 8812 6644 8818 6656
rect 9122 6644 9128 6656
rect 8812 6616 9128 6644
rect 8812 6604 8818 6616
rect 9122 6604 9128 6616
rect 9180 6604 9186 6656
rect 9214 6604 9220 6656
rect 9272 6644 9278 6656
rect 9309 6647 9367 6653
rect 9309 6644 9321 6647
rect 9272 6616 9321 6644
rect 9272 6604 9278 6616
rect 9309 6613 9321 6616
rect 9355 6613 9367 6647
rect 10152 6644 10180 6684
rect 10318 6672 10324 6684
rect 10376 6672 10382 6724
rect 10428 6712 10456 6752
rect 10502 6740 10508 6792
rect 10560 6780 10566 6792
rect 12912 6780 12940 6820
rect 14918 6808 14924 6860
rect 14976 6848 14982 6860
rect 16942 6848 16948 6860
rect 14976 6820 16948 6848
rect 14976 6808 14982 6820
rect 16942 6808 16948 6820
rect 17000 6808 17006 6860
rect 17678 6808 17684 6860
rect 17736 6848 17742 6860
rect 19245 6851 19303 6857
rect 19245 6848 19257 6851
rect 17736 6820 19257 6848
rect 17736 6808 17742 6820
rect 19245 6817 19257 6820
rect 19291 6817 19303 6851
rect 19245 6811 19303 6817
rect 20254 6808 20260 6860
rect 20312 6848 20318 6860
rect 22278 6848 22284 6860
rect 20312 6820 22284 6848
rect 20312 6808 20318 6820
rect 22278 6808 22284 6820
rect 22336 6808 22342 6860
rect 23382 6808 23388 6860
rect 23440 6848 23446 6860
rect 23566 6848 23572 6860
rect 23440 6820 23572 6848
rect 23440 6808 23446 6820
rect 23566 6808 23572 6820
rect 23624 6848 23630 6860
rect 24026 6848 24032 6860
rect 23624 6820 24032 6848
rect 23624 6808 23630 6820
rect 24026 6808 24032 6820
rect 24084 6808 24090 6860
rect 24118 6808 24124 6860
rect 24176 6848 24182 6860
rect 24397 6851 24455 6857
rect 24397 6848 24409 6851
rect 24176 6820 24409 6848
rect 24176 6808 24182 6820
rect 24397 6817 24409 6820
rect 24443 6817 24455 6851
rect 24397 6811 24455 6817
rect 25130 6808 25136 6860
rect 25188 6848 25194 6860
rect 25777 6851 25835 6857
rect 25777 6848 25789 6851
rect 25188 6820 25789 6848
rect 25188 6808 25194 6820
rect 25777 6817 25789 6820
rect 25823 6817 25835 6851
rect 25777 6811 25835 6817
rect 13265 6783 13323 6789
rect 13265 6780 13277 6783
rect 10560 6759 11374 6780
rect 10560 6753 11391 6759
rect 10560 6752 11345 6753
rect 10560 6740 10566 6752
rect 10686 6712 10692 6724
rect 10428 6684 10692 6712
rect 10686 6672 10692 6684
rect 10744 6672 10750 6724
rect 11333 6719 11345 6752
rect 11379 6719 11391 6753
rect 12912 6752 13277 6780
rect 13265 6749 13277 6752
rect 13311 6749 13323 6783
rect 13538 6780 13544 6792
rect 13499 6752 13544 6780
rect 13265 6743 13323 6749
rect 13538 6740 13544 6752
rect 13596 6740 13602 6792
rect 14090 6780 14096 6792
rect 14051 6752 14096 6780
rect 14090 6740 14096 6752
rect 14148 6740 14154 6792
rect 14642 6740 14648 6792
rect 14700 6780 14706 6792
rect 15013 6783 15071 6789
rect 15013 6780 15025 6783
rect 14700 6752 15025 6780
rect 14700 6740 14706 6752
rect 15013 6749 15025 6752
rect 15059 6749 15071 6783
rect 15841 6783 15899 6789
rect 15841 6780 15853 6783
rect 15013 6743 15071 6749
rect 15212 6752 15853 6780
rect 11333 6713 11391 6719
rect 12250 6672 12256 6724
rect 12308 6712 12314 6724
rect 12308 6684 12664 6712
rect 12308 6672 12314 6684
rect 10594 6644 10600 6656
rect 10152 6616 10600 6644
rect 9309 6607 9367 6613
rect 10594 6604 10600 6616
rect 10652 6644 10658 6656
rect 11422 6644 11428 6656
rect 10652 6616 11428 6644
rect 10652 6604 10658 6616
rect 11422 6604 11428 6616
rect 11480 6604 11486 6656
rect 11514 6604 11520 6656
rect 11572 6644 11578 6656
rect 12069 6647 12127 6653
rect 12069 6644 12081 6647
rect 11572 6616 12081 6644
rect 11572 6604 11578 6616
rect 12069 6613 12081 6616
rect 12115 6644 12127 6647
rect 12529 6647 12587 6653
rect 12529 6644 12541 6647
rect 12115 6616 12541 6644
rect 12115 6613 12127 6616
rect 12069 6607 12127 6613
rect 12529 6613 12541 6616
rect 12575 6613 12587 6647
rect 12636 6644 12664 6684
rect 15212 6653 15240 6752
rect 15841 6749 15853 6752
rect 15887 6749 15899 6783
rect 15841 6743 15899 6749
rect 16485 6783 16543 6789
rect 16485 6749 16497 6783
rect 16531 6780 16543 6783
rect 17126 6780 17132 6792
rect 16531 6752 17132 6780
rect 16531 6749 16543 6752
rect 16485 6743 16543 6749
rect 14277 6647 14335 6653
rect 14277 6644 14289 6647
rect 12636 6616 14289 6644
rect 12529 6607 12587 6613
rect 14277 6613 14289 6616
rect 14323 6613 14335 6647
rect 14277 6607 14335 6613
rect 15197 6647 15255 6653
rect 15197 6613 15209 6647
rect 15243 6613 15255 6647
rect 15856 6644 15884 6743
rect 17126 6740 17132 6752
rect 17184 6740 17190 6792
rect 17221 6783 17279 6789
rect 17221 6749 17233 6783
rect 17267 6749 17279 6783
rect 17221 6743 17279 6749
rect 18693 6783 18751 6789
rect 18693 6749 18705 6783
rect 18739 6749 18751 6783
rect 19518 6780 19524 6792
rect 19479 6752 19524 6780
rect 18693 6743 18751 6749
rect 16574 6672 16580 6724
rect 16632 6712 16638 6724
rect 17236 6712 17264 6743
rect 16632 6684 17264 6712
rect 18708 6712 18736 6743
rect 19518 6740 19524 6752
rect 19576 6740 19582 6792
rect 21177 6783 21235 6789
rect 21177 6749 21189 6783
rect 21223 6749 21235 6783
rect 21634 6780 21640 6792
rect 21595 6752 21640 6780
rect 21177 6743 21235 6749
rect 20070 6712 20076 6724
rect 18708 6684 20076 6712
rect 16632 6672 16638 6684
rect 20070 6672 20076 6684
rect 20128 6672 20134 6724
rect 21192 6712 21220 6743
rect 21634 6740 21640 6752
rect 21692 6740 21698 6792
rect 22554 6780 22560 6792
rect 22515 6752 22560 6780
rect 22554 6740 22560 6752
rect 22612 6740 22618 6792
rect 24854 6780 24860 6792
rect 23492 6752 24860 6780
rect 23492 6712 23520 6752
rect 24854 6740 24860 6752
rect 24912 6740 24918 6792
rect 25869 6783 25927 6789
rect 25869 6780 25881 6783
rect 24964 6752 25881 6780
rect 21192 6684 23520 6712
rect 23566 6672 23572 6724
rect 23624 6712 23630 6724
rect 24964 6721 24992 6752
rect 25869 6749 25881 6752
rect 25915 6749 25927 6783
rect 25869 6743 25927 6749
rect 24949 6715 25007 6721
rect 24949 6712 24961 6715
rect 23624 6684 24961 6712
rect 23624 6672 23630 6684
rect 24949 6681 24961 6684
rect 24995 6681 25007 6715
rect 24949 6675 25007 6681
rect 25133 6715 25191 6721
rect 25133 6681 25145 6715
rect 25179 6712 25191 6715
rect 25222 6712 25228 6724
rect 25179 6684 25228 6712
rect 25179 6681 25191 6684
rect 25133 6675 25191 6681
rect 25222 6672 25228 6684
rect 25280 6672 25286 6724
rect 25317 6715 25375 6721
rect 25317 6681 25329 6715
rect 25363 6712 25375 6715
rect 25976 6712 26004 6888
rect 26050 6876 26056 6888
rect 26108 6916 26114 6928
rect 26418 6916 26424 6928
rect 26108 6888 26424 6916
rect 26108 6876 26114 6888
rect 26418 6876 26424 6888
rect 26476 6876 26482 6928
rect 26970 6916 26976 6928
rect 26931 6888 26976 6916
rect 26970 6876 26976 6888
rect 27028 6876 27034 6928
rect 30576 6916 30604 6947
rect 33410 6944 33416 6956
rect 33468 6944 33474 6996
rect 33594 6944 33600 6996
rect 33652 6984 33658 6996
rect 36170 6984 36176 6996
rect 33652 6956 36176 6984
rect 33652 6944 33658 6956
rect 36170 6944 36176 6956
rect 36228 6944 36234 6996
rect 36354 6984 36360 6996
rect 36315 6956 36360 6984
rect 36354 6944 36360 6956
rect 36412 6944 36418 6996
rect 37642 6984 37648 6996
rect 36924 6956 37648 6984
rect 32214 6916 32220 6928
rect 28552 6888 30604 6916
rect 31726 6888 32220 6916
rect 28552 6848 28580 6888
rect 28718 6848 28724 6860
rect 25363 6684 26004 6712
rect 26068 6820 28580 6848
rect 28679 6820 28724 6848
rect 25363 6681 25375 6684
rect 25317 6675 25375 6681
rect 18230 6644 18236 6656
rect 15856 6616 18236 6644
rect 15197 6607 15255 6613
rect 18230 6604 18236 6616
rect 18288 6604 18294 6656
rect 18414 6604 18420 6656
rect 18472 6644 18478 6656
rect 20257 6647 20315 6653
rect 20257 6644 20269 6647
rect 18472 6616 20269 6644
rect 18472 6604 18478 6616
rect 20257 6613 20269 6616
rect 20303 6644 20315 6647
rect 22094 6644 22100 6656
rect 20303 6616 22100 6644
rect 20303 6613 20315 6616
rect 20257 6607 20315 6613
rect 22094 6604 22100 6616
rect 22152 6644 22158 6656
rect 23290 6644 23296 6656
rect 22152 6616 23296 6644
rect 22152 6604 22158 6616
rect 23290 6604 23296 6616
rect 23348 6604 23354 6656
rect 24026 6604 24032 6656
rect 24084 6644 24090 6656
rect 26068 6644 26096 6820
rect 28718 6808 28724 6820
rect 28776 6848 28782 6860
rect 31481 6851 31539 6857
rect 28776 6820 30052 6848
rect 28776 6808 28782 6820
rect 26145 6783 26203 6789
rect 26145 6749 26157 6783
rect 26191 6780 26203 6783
rect 28994 6780 29000 6792
rect 26191 6752 27752 6780
rect 28955 6752 29000 6780
rect 26191 6749 26203 6752
rect 26145 6743 26203 6749
rect 26418 6672 26424 6724
rect 26476 6712 26482 6724
rect 26605 6715 26663 6721
rect 26605 6712 26617 6715
rect 26476 6684 26617 6712
rect 26476 6672 26482 6684
rect 26605 6681 26617 6684
rect 26651 6681 26663 6715
rect 26605 6675 26663 6681
rect 24084 6616 26096 6644
rect 26620 6644 26648 6675
rect 26694 6672 26700 6724
rect 26752 6712 26758 6724
rect 26789 6715 26847 6721
rect 26789 6712 26801 6715
rect 26752 6684 26801 6712
rect 26752 6672 26758 6684
rect 26789 6681 26801 6684
rect 26835 6712 26847 6715
rect 27430 6712 27436 6724
rect 26835 6684 27436 6712
rect 26835 6681 26847 6684
rect 26789 6675 26847 6681
rect 27430 6672 27436 6684
rect 27488 6712 27494 6724
rect 27724 6721 27752 6752
rect 28994 6740 29000 6752
rect 29052 6740 29058 6792
rect 30024 6789 30052 6820
rect 31481 6817 31493 6851
rect 31527 6848 31539 6851
rect 31726 6848 31754 6888
rect 32214 6876 32220 6888
rect 32272 6876 32278 6928
rect 32582 6916 32588 6928
rect 32324 6888 32588 6916
rect 32030 6848 32036 6860
rect 31527 6820 31754 6848
rect 31991 6820 32036 6848
rect 31527 6817 31539 6820
rect 31481 6811 31539 6817
rect 32030 6808 32036 6820
rect 32088 6808 32094 6860
rect 30009 6783 30067 6789
rect 30009 6749 30021 6783
rect 30055 6780 30067 6783
rect 30469 6783 30527 6789
rect 30469 6780 30481 6783
rect 30055 6752 30481 6780
rect 30055 6749 30067 6752
rect 30009 6743 30067 6749
rect 30469 6749 30481 6752
rect 30515 6780 30527 6783
rect 30558 6780 30564 6792
rect 30515 6752 30564 6780
rect 30515 6749 30527 6752
rect 30469 6743 30527 6749
rect 30558 6740 30564 6752
rect 30616 6740 30622 6792
rect 30653 6783 30711 6789
rect 30653 6749 30665 6783
rect 30699 6749 30711 6783
rect 30653 6743 30711 6749
rect 27525 6715 27583 6721
rect 27525 6712 27537 6715
rect 27488 6684 27537 6712
rect 27488 6672 27494 6684
rect 27525 6681 27537 6684
rect 27571 6681 27583 6715
rect 27525 6675 27583 6681
rect 27709 6715 27767 6721
rect 27709 6681 27721 6715
rect 27755 6712 27767 6715
rect 28902 6712 28908 6724
rect 27755 6684 28908 6712
rect 27755 6681 27767 6684
rect 27709 6675 27767 6681
rect 28902 6672 28908 6684
rect 28960 6712 28966 6724
rect 30374 6712 30380 6724
rect 28960 6684 30380 6712
rect 28960 6672 28966 6684
rect 30374 6672 30380 6684
rect 30432 6712 30438 6724
rect 30668 6712 30696 6743
rect 31846 6740 31852 6792
rect 31904 6780 31910 6792
rect 31941 6783 31999 6789
rect 31941 6780 31953 6783
rect 31904 6752 31953 6780
rect 31904 6740 31910 6752
rect 31941 6749 31953 6752
rect 31987 6749 31999 6783
rect 32324 6780 32352 6888
rect 32582 6876 32588 6888
rect 32640 6916 32646 6928
rect 33134 6916 33140 6928
rect 32640 6888 33140 6916
rect 32640 6876 32646 6888
rect 33134 6876 33140 6888
rect 33192 6916 33198 6928
rect 36924 6916 36952 6956
rect 37642 6944 37648 6956
rect 37700 6944 37706 6996
rect 37734 6944 37740 6996
rect 37792 6984 37798 6996
rect 42886 6984 42892 6996
rect 37792 6956 42892 6984
rect 37792 6944 37798 6956
rect 42886 6944 42892 6956
rect 42944 6944 42950 6996
rect 43070 6944 43076 6996
rect 43128 6984 43134 6996
rect 48590 6984 48596 6996
rect 43128 6956 44404 6984
rect 48551 6956 48596 6984
rect 43128 6944 43134 6956
rect 33192 6888 36952 6916
rect 37829 6919 37887 6925
rect 33192 6876 33198 6888
rect 35802 6848 35808 6860
rect 35763 6820 35808 6848
rect 35802 6808 35808 6820
rect 35860 6808 35866 6860
rect 36188 6857 36216 6888
rect 37829 6885 37841 6919
rect 37875 6885 37887 6919
rect 41598 6916 41604 6928
rect 41559 6888 41604 6916
rect 37829 6879 37887 6885
rect 36173 6851 36231 6857
rect 36173 6817 36185 6851
rect 36219 6817 36231 6851
rect 36173 6811 36231 6817
rect 37844 6848 37872 6879
rect 41598 6876 41604 6888
rect 41656 6876 41662 6928
rect 44376 6916 44404 6956
rect 48590 6944 48596 6956
rect 48648 6944 48654 6996
rect 49234 6944 49240 6996
rect 49292 6984 49298 6996
rect 51258 6984 51264 6996
rect 49292 6956 51074 6984
rect 51219 6956 51264 6984
rect 49292 6944 49298 6956
rect 51046 6916 51074 6956
rect 51258 6944 51264 6956
rect 51316 6944 51322 6996
rect 52362 6944 52368 6996
rect 52420 6984 52426 6996
rect 55858 6984 55864 6996
rect 52420 6956 53788 6984
rect 55819 6956 55864 6984
rect 52420 6944 52426 6956
rect 52270 6916 52276 6928
rect 44376 6888 44496 6916
rect 51046 6888 52276 6916
rect 38746 6848 38752 6860
rect 37844 6820 38752 6848
rect 32401 6783 32459 6789
rect 32401 6780 32413 6783
rect 31941 6743 31999 6749
rect 32232 6752 32413 6780
rect 30432 6684 30696 6712
rect 30432 6672 30438 6684
rect 31386 6672 31392 6724
rect 31444 6712 31450 6724
rect 32232 6712 32260 6752
rect 32401 6749 32413 6752
rect 32447 6749 32459 6783
rect 32401 6743 32459 6749
rect 32490 6740 32496 6792
rect 32548 6780 32554 6792
rect 33229 6783 33287 6789
rect 33229 6780 33241 6783
rect 32548 6752 33241 6780
rect 32548 6740 32554 6752
rect 33229 6749 33241 6752
rect 33275 6780 33287 6783
rect 33870 6780 33876 6792
rect 33275 6752 33876 6780
rect 33275 6749 33287 6752
rect 33229 6743 33287 6749
rect 33870 6740 33876 6752
rect 33928 6740 33934 6792
rect 33965 6783 34023 6789
rect 33965 6749 33977 6783
rect 34011 6780 34023 6783
rect 36814 6780 36820 6792
rect 34011 6752 35664 6780
rect 36775 6752 36820 6780
rect 34011 6749 34023 6752
rect 33965 6743 34023 6749
rect 32950 6712 32956 6724
rect 31444 6684 32260 6712
rect 32324 6684 32956 6712
rect 31444 6672 31450 6684
rect 28994 6644 29000 6656
rect 26620 6616 29000 6644
rect 24084 6604 24090 6616
rect 28994 6604 29000 6616
rect 29052 6604 29058 6656
rect 29454 6604 29460 6656
rect 29512 6644 29518 6656
rect 29549 6647 29607 6653
rect 29549 6644 29561 6647
rect 29512 6616 29561 6644
rect 29512 6604 29518 6616
rect 29549 6613 29561 6616
rect 29595 6613 29607 6647
rect 29549 6607 29607 6613
rect 29822 6604 29828 6656
rect 29880 6644 29886 6656
rect 32324 6644 32352 6684
rect 32950 6672 32956 6684
rect 33008 6672 33014 6724
rect 34422 6672 34428 6724
rect 34480 6712 34486 6724
rect 35069 6715 35127 6721
rect 35069 6712 35081 6715
rect 34480 6684 35081 6712
rect 34480 6672 34486 6684
rect 35069 6681 35081 6684
rect 35115 6681 35127 6715
rect 35069 6675 35127 6681
rect 35253 6715 35311 6721
rect 35253 6681 35265 6715
rect 35299 6681 35311 6715
rect 35636 6712 35664 6752
rect 36814 6740 36820 6752
rect 36872 6740 36878 6792
rect 37090 6780 37096 6792
rect 37051 6752 37096 6780
rect 37090 6740 37096 6752
rect 37148 6740 37154 6792
rect 37274 6740 37280 6792
rect 37332 6780 37338 6792
rect 37844 6780 37872 6820
rect 38746 6808 38752 6820
rect 38804 6808 38810 6860
rect 38838 6808 38844 6860
rect 38896 6848 38902 6860
rect 39025 6851 39083 6857
rect 39025 6848 39037 6851
rect 38896 6820 39037 6848
rect 38896 6808 38902 6820
rect 39025 6817 39037 6820
rect 39071 6817 39083 6851
rect 39025 6811 39083 6817
rect 40034 6808 40040 6860
rect 40092 6848 40098 6860
rect 44468 6857 44496 6888
rect 52270 6876 52276 6888
rect 52328 6876 52334 6928
rect 53760 6916 53788 6956
rect 55858 6944 55864 6956
rect 55916 6944 55922 6996
rect 56781 6919 56839 6925
rect 56781 6916 56793 6919
rect 53760 6888 56793 6916
rect 56781 6885 56793 6888
rect 56827 6885 56839 6919
rect 56781 6879 56839 6885
rect 40221 6851 40279 6857
rect 40221 6848 40233 6851
rect 40092 6820 40233 6848
rect 40092 6808 40098 6820
rect 40221 6817 40233 6820
rect 40267 6817 40279 6851
rect 40221 6811 40279 6817
rect 44453 6851 44511 6857
rect 44453 6817 44465 6851
rect 44499 6848 44511 6851
rect 45002 6848 45008 6860
rect 44499 6820 45008 6848
rect 44499 6817 44511 6820
rect 44453 6811 44511 6817
rect 45002 6808 45008 6820
rect 45060 6808 45066 6860
rect 51997 6851 52055 6857
rect 51997 6817 52009 6851
rect 52043 6848 52055 6851
rect 52454 6848 52460 6860
rect 52043 6820 52460 6848
rect 52043 6817 52055 6820
rect 51997 6811 52055 6817
rect 52454 6808 52460 6820
rect 52512 6808 52518 6860
rect 53837 6851 53895 6857
rect 53837 6817 53849 6851
rect 53883 6848 53895 6851
rect 54110 6848 54116 6860
rect 53883 6820 54116 6848
rect 53883 6817 53895 6820
rect 53837 6811 53895 6817
rect 54110 6808 54116 6820
rect 54168 6808 54174 6860
rect 57790 6808 57796 6860
rect 57848 6848 57854 6860
rect 57848 6820 57893 6848
rect 57848 6808 57854 6820
rect 38378 6780 38384 6792
rect 37332 6752 37872 6780
rect 38339 6752 38384 6780
rect 37332 6740 37338 6752
rect 38378 6740 38384 6752
rect 38436 6740 38442 6792
rect 38470 6740 38476 6792
rect 38528 6780 38534 6792
rect 41325 6783 41383 6789
rect 41325 6780 41337 6783
rect 38528 6752 41337 6780
rect 38528 6740 38534 6752
rect 41325 6749 41337 6752
rect 41371 6780 41383 6783
rect 41690 6780 41696 6792
rect 41371 6752 41696 6780
rect 41371 6749 41383 6752
rect 41325 6743 41383 6749
rect 41690 6740 41696 6752
rect 41748 6740 41754 6792
rect 42426 6780 42432 6792
rect 42387 6752 42432 6780
rect 42426 6740 42432 6752
rect 42484 6740 42490 6792
rect 43990 6740 43996 6792
rect 44048 6780 44054 6792
rect 44177 6783 44235 6789
rect 44177 6780 44189 6783
rect 44048 6752 44189 6780
rect 44048 6740 44054 6752
rect 44177 6749 44189 6752
rect 44223 6749 44235 6783
rect 44177 6743 44235 6749
rect 45281 6783 45339 6789
rect 45281 6749 45293 6783
rect 45327 6749 45339 6783
rect 46566 6780 46572 6792
rect 46527 6752 46572 6780
rect 45281 6743 45339 6749
rect 37458 6712 37464 6724
rect 35636 6684 37464 6712
rect 35253 6675 35311 6681
rect 29880 6616 32352 6644
rect 29880 6604 29886 6616
rect 32398 6604 32404 6656
rect 32456 6644 32462 6656
rect 33051 6647 33109 6653
rect 33051 6644 33063 6647
rect 32456 6616 33063 6644
rect 32456 6604 32462 6616
rect 33051 6613 33063 6616
rect 33097 6613 33109 6647
rect 33051 6607 33109 6613
rect 33137 6647 33195 6653
rect 33137 6613 33149 6647
rect 33183 6644 33195 6647
rect 33226 6644 33232 6656
rect 33183 6616 33232 6644
rect 33183 6613 33195 6616
rect 33137 6607 33195 6613
rect 33226 6604 33232 6616
rect 33284 6604 33290 6656
rect 34149 6647 34207 6653
rect 34149 6613 34161 6647
rect 34195 6644 34207 6647
rect 34698 6644 34704 6656
rect 34195 6616 34704 6644
rect 34195 6613 34207 6616
rect 34149 6607 34207 6613
rect 34698 6604 34704 6616
rect 34756 6604 34762 6656
rect 35268 6644 35296 6675
rect 37458 6672 37464 6684
rect 37516 6672 37522 6724
rect 38930 6712 38936 6724
rect 37752 6684 38936 6712
rect 35802 6644 35808 6656
rect 35268 6616 35808 6644
rect 35802 6604 35808 6616
rect 35860 6604 35866 6656
rect 35986 6644 35992 6656
rect 35947 6616 35992 6644
rect 35986 6604 35992 6616
rect 36044 6604 36050 6656
rect 36814 6604 36820 6656
rect 36872 6644 36878 6656
rect 37752 6644 37780 6684
rect 38930 6672 38936 6684
rect 38988 6672 38994 6724
rect 39209 6715 39267 6721
rect 39209 6681 39221 6715
rect 39255 6712 39267 6715
rect 40402 6712 40408 6724
rect 39255 6684 40408 6712
rect 39255 6681 39267 6684
rect 39209 6675 39267 6681
rect 40402 6672 40408 6684
rect 40460 6712 40466 6724
rect 40862 6712 40868 6724
rect 40460 6684 40868 6712
rect 40460 6672 40466 6684
rect 40862 6672 40868 6684
rect 40920 6672 40926 6724
rect 41601 6715 41659 6721
rect 41601 6712 41613 6715
rect 40972 6684 41613 6712
rect 36872 6616 37780 6644
rect 38565 6647 38623 6653
rect 36872 6604 36878 6616
rect 38565 6613 38577 6647
rect 38611 6644 38623 6647
rect 38654 6644 38660 6656
rect 38611 6616 38660 6644
rect 38611 6613 38623 6616
rect 38565 6607 38623 6613
rect 38654 6604 38660 6616
rect 38712 6604 38718 6656
rect 39298 6604 39304 6656
rect 39356 6644 39362 6656
rect 40972 6644 41000 6684
rect 41601 6681 41613 6684
rect 41647 6712 41659 6715
rect 41782 6712 41788 6724
rect 41647 6684 41788 6712
rect 41647 6681 41659 6684
rect 41601 6675 41659 6681
rect 41782 6672 41788 6684
rect 41840 6672 41846 6724
rect 42610 6712 42616 6724
rect 42571 6684 42616 6712
rect 42610 6672 42616 6684
rect 42668 6672 42674 6724
rect 43346 6672 43352 6724
rect 43404 6712 43410 6724
rect 45296 6712 45324 6743
rect 46566 6740 46572 6752
rect 46624 6740 46630 6792
rect 46842 6780 46848 6792
rect 46803 6752 46848 6780
rect 46842 6740 46848 6752
rect 46900 6740 46906 6792
rect 47504 6752 49280 6780
rect 43404 6684 45324 6712
rect 46584 6712 46612 6740
rect 47504 6712 47532 6752
rect 48590 6712 48596 6724
rect 46584 6684 47532 6712
rect 47596 6684 48596 6712
rect 43404 6672 43410 6684
rect 39356 6616 41000 6644
rect 41417 6647 41475 6653
rect 39356 6604 39362 6616
rect 41417 6613 41429 6647
rect 41463 6644 41475 6647
rect 41966 6644 41972 6656
rect 41463 6616 41972 6644
rect 41463 6613 41475 6616
rect 41417 6607 41475 6613
rect 41966 6604 41972 6616
rect 42024 6644 42030 6656
rect 42628 6644 42656 6672
rect 42024 6616 42656 6644
rect 42024 6604 42030 6616
rect 42702 6604 42708 6656
rect 42760 6644 42766 6656
rect 47596 6653 47624 6684
rect 48590 6672 48596 6684
rect 48648 6672 48654 6724
rect 43441 6647 43499 6653
rect 43441 6644 43453 6647
rect 42760 6616 43453 6644
rect 42760 6604 42766 6616
rect 43441 6613 43453 6616
rect 43487 6644 43499 6647
rect 46017 6647 46075 6653
rect 46017 6644 46029 6647
rect 43487 6616 46029 6644
rect 43487 6613 43499 6616
rect 43441 6607 43499 6613
rect 46017 6613 46029 6616
rect 46063 6644 46075 6647
rect 47581 6647 47639 6653
rect 47581 6644 47593 6647
rect 46063 6616 47593 6644
rect 46063 6613 46075 6616
rect 46017 6607 46075 6613
rect 47581 6613 47593 6616
rect 47627 6613 47639 6647
rect 48038 6644 48044 6656
rect 47999 6616 48044 6644
rect 47581 6607 47639 6613
rect 48038 6604 48044 6616
rect 48096 6604 48102 6656
rect 49252 6644 49280 6752
rect 49326 6740 49332 6792
rect 49384 6780 49390 6792
rect 49605 6783 49663 6789
rect 49384 6752 49429 6780
rect 49384 6740 49390 6752
rect 49605 6749 49617 6783
rect 49651 6780 49663 6783
rect 50249 6783 50307 6789
rect 50249 6780 50261 6783
rect 49651 6752 50261 6780
rect 49651 6749 49663 6752
rect 49605 6743 49663 6749
rect 49988 6644 50016 6752
rect 50249 6749 50261 6752
rect 50295 6749 50307 6783
rect 50522 6780 50528 6792
rect 50483 6752 50528 6780
rect 50249 6743 50307 6749
rect 50264 6712 50292 6743
rect 50522 6740 50528 6752
rect 50580 6740 50586 6792
rect 52822 6780 52828 6792
rect 51046 6752 52828 6780
rect 51046 6712 51074 6752
rect 52822 6740 52828 6752
rect 52880 6740 52886 6792
rect 53561 6783 53619 6789
rect 53561 6749 53573 6783
rect 53607 6780 53619 6783
rect 57514 6780 57520 6792
rect 53607 6752 55812 6780
rect 57475 6752 57520 6780
rect 53607 6749 53619 6752
rect 53561 6743 53619 6749
rect 50264 6684 51074 6712
rect 51813 6715 51871 6721
rect 51813 6681 51825 6715
rect 51859 6712 51871 6715
rect 52178 6712 52184 6724
rect 51859 6684 52184 6712
rect 51859 6681 51871 6684
rect 51813 6675 51871 6681
rect 52178 6672 52184 6684
rect 52236 6672 52242 6724
rect 54297 6715 54355 6721
rect 54297 6712 54309 6715
rect 52748 6684 54309 6712
rect 52748 6656 52776 6684
rect 54297 6681 54309 6684
rect 54343 6681 54355 6715
rect 55674 6712 55680 6724
rect 55635 6684 55680 6712
rect 54297 6675 54355 6681
rect 55674 6672 55680 6684
rect 55732 6672 55738 6724
rect 55784 6712 55812 6752
rect 57514 6740 57520 6752
rect 57572 6740 57578 6792
rect 57974 6712 57980 6724
rect 55784 6684 57980 6712
rect 57974 6672 57980 6684
rect 58032 6672 58038 6724
rect 49252 6616 50016 6644
rect 51442 6604 51448 6656
rect 51500 6644 51506 6656
rect 52730 6644 52736 6656
rect 51500 6616 52736 6644
rect 51500 6604 51506 6616
rect 52730 6604 52736 6616
rect 52788 6604 52794 6656
rect 52825 6647 52883 6653
rect 52825 6613 52837 6647
rect 52871 6644 52883 6647
rect 52914 6644 52920 6656
rect 52871 6616 52920 6644
rect 52871 6613 52883 6616
rect 52825 6607 52883 6613
rect 52914 6604 52920 6616
rect 52972 6604 52978 6656
rect 55582 6604 55588 6656
rect 55640 6644 55646 6656
rect 55877 6647 55935 6653
rect 55877 6644 55889 6647
rect 55640 6616 55889 6644
rect 55640 6604 55646 6616
rect 55877 6613 55889 6616
rect 55923 6613 55935 6647
rect 56042 6644 56048 6656
rect 56003 6616 56048 6644
rect 55877 6607 55935 6613
rect 56042 6604 56048 6616
rect 56100 6604 56106 6656
rect 1104 6554 58880 6576
rect 1104 6502 15398 6554
rect 15450 6502 15462 6554
rect 15514 6502 15526 6554
rect 15578 6502 15590 6554
rect 15642 6502 15654 6554
rect 15706 6502 29846 6554
rect 29898 6502 29910 6554
rect 29962 6502 29974 6554
rect 30026 6502 30038 6554
rect 30090 6502 30102 6554
rect 30154 6502 44294 6554
rect 44346 6502 44358 6554
rect 44410 6502 44422 6554
rect 44474 6502 44486 6554
rect 44538 6502 44550 6554
rect 44602 6502 58880 6554
rect 1104 6480 58880 6502
rect 2130 6400 2136 6452
rect 2188 6440 2194 6452
rect 5442 6440 5448 6452
rect 2188 6412 5448 6440
rect 2188 6400 2194 6412
rect 5442 6400 5448 6412
rect 5500 6400 5506 6452
rect 7834 6400 7840 6452
rect 7892 6440 7898 6452
rect 8297 6443 8355 6449
rect 8297 6440 8309 6443
rect 7892 6412 8309 6440
rect 7892 6400 7898 6412
rect 8297 6409 8309 6412
rect 8343 6440 8355 6443
rect 9766 6440 9772 6452
rect 8343 6412 9772 6440
rect 8343 6409 8355 6412
rect 8297 6403 8355 6409
rect 9766 6400 9772 6412
rect 9824 6440 9830 6452
rect 9861 6443 9919 6449
rect 9861 6440 9873 6443
rect 9824 6412 9873 6440
rect 9824 6400 9830 6412
rect 9861 6409 9873 6412
rect 9907 6409 9919 6443
rect 9861 6403 9919 6409
rect 10042 6400 10048 6452
rect 10100 6440 10106 6452
rect 11146 6440 11152 6452
rect 10100 6412 11152 6440
rect 10100 6400 10106 6412
rect 11146 6400 11152 6412
rect 11204 6400 11210 6452
rect 19334 6440 19340 6452
rect 13924 6412 19340 6440
rect 5902 6372 5908 6384
rect 2700 6344 5908 6372
rect 2041 6307 2099 6313
rect 2041 6273 2053 6307
rect 2087 6304 2099 6307
rect 2130 6304 2136 6316
rect 2087 6276 2136 6304
rect 2087 6273 2099 6276
rect 2041 6267 2099 6273
rect 2130 6264 2136 6276
rect 2188 6264 2194 6316
rect 2498 6304 2504 6316
rect 2459 6276 2504 6304
rect 2498 6264 2504 6276
rect 2556 6264 2562 6316
rect 2700 6177 2728 6344
rect 5902 6332 5908 6344
rect 5960 6332 5966 6384
rect 6730 6332 6736 6384
rect 6788 6372 6794 6384
rect 6788 6344 9812 6372
rect 6788 6332 6794 6344
rect 3878 6304 3884 6316
rect 3839 6276 3884 6304
rect 3878 6264 3884 6276
rect 3936 6264 3942 6316
rect 3970 6264 3976 6316
rect 4028 6304 4034 6316
rect 4028 6276 4200 6304
rect 4028 6264 4034 6276
rect 4172 6245 4200 6276
rect 4246 6264 4252 6316
rect 4304 6304 4310 6316
rect 4617 6307 4675 6313
rect 4617 6304 4629 6307
rect 4304 6276 4629 6304
rect 4304 6264 4310 6276
rect 4617 6273 4629 6276
rect 4663 6273 4675 6307
rect 4617 6267 4675 6273
rect 4801 6307 4859 6313
rect 4801 6273 4813 6307
rect 4847 6273 4859 6307
rect 4801 6267 4859 6273
rect 4896 6310 4954 6316
rect 4896 6276 4908 6310
rect 4942 6276 4954 6310
rect 4896 6270 4954 6276
rect 4985 6310 5043 6313
rect 5166 6310 5172 6316
rect 4985 6307 5172 6310
rect 4985 6273 4997 6307
rect 5031 6282 5172 6307
rect 5031 6273 5043 6282
rect 4157 6239 4215 6245
rect 4157 6205 4169 6239
rect 4203 6236 4215 6239
rect 4338 6236 4344 6248
rect 4203 6208 4344 6236
rect 4203 6205 4215 6208
rect 4157 6199 4215 6205
rect 4338 6196 4344 6208
rect 4396 6196 4402 6248
rect 4816 6236 4844 6267
rect 4724 6208 4844 6236
rect 4908 6236 4936 6270
rect 4985 6267 5043 6273
rect 5166 6264 5172 6282
rect 5224 6264 5230 6316
rect 5534 6264 5540 6316
rect 5592 6304 5598 6316
rect 7561 6307 7619 6313
rect 7561 6304 7573 6307
rect 5592 6276 7573 6304
rect 5592 6264 5598 6276
rect 7561 6273 7573 6276
rect 7607 6273 7619 6307
rect 9122 6304 9128 6316
rect 9083 6276 9128 6304
rect 7561 6267 7619 6273
rect 9122 6264 9128 6276
rect 9180 6264 9186 6316
rect 4908 6208 5028 6236
rect 2685 6171 2743 6177
rect 2685 6137 2697 6171
rect 2731 6137 2743 6171
rect 2685 6131 2743 6137
rect 4246 6128 4252 6180
rect 4304 6168 4310 6180
rect 4724 6168 4752 6208
rect 4304 6140 4752 6168
rect 4304 6128 4310 6140
rect 4798 6128 4804 6180
rect 4856 6168 4862 6180
rect 5000 6168 5028 6208
rect 5350 6196 5356 6248
rect 5408 6236 5414 6248
rect 5718 6236 5724 6248
rect 5408 6208 5724 6236
rect 5408 6196 5414 6208
rect 5718 6196 5724 6208
rect 5776 6236 5782 6248
rect 7285 6239 7343 6245
rect 7285 6236 7297 6239
rect 5776 6208 7297 6236
rect 5776 6196 5782 6208
rect 7285 6205 7297 6208
rect 7331 6205 7343 6239
rect 7285 6199 7343 6205
rect 8849 6239 8907 6245
rect 8849 6205 8861 6239
rect 8895 6205 8907 6239
rect 9784 6236 9812 6344
rect 9876 6344 10456 6372
rect 9876 6316 9904 6344
rect 9858 6264 9864 6316
rect 9916 6264 9922 6316
rect 10309 6307 10367 6313
rect 10244 6279 10321 6307
rect 10244 6236 10272 6279
rect 10309 6273 10321 6279
rect 10355 6273 10367 6307
rect 10428 6304 10456 6344
rect 11422 6332 11428 6384
rect 11480 6372 11486 6384
rect 13924 6372 13952 6412
rect 19334 6400 19340 6412
rect 19392 6400 19398 6452
rect 19797 6443 19855 6449
rect 19797 6409 19809 6443
rect 19843 6440 19855 6443
rect 22554 6440 22560 6452
rect 19843 6412 22560 6440
rect 19843 6409 19855 6412
rect 19797 6403 19855 6409
rect 22554 6400 22560 6412
rect 22612 6400 22618 6452
rect 23474 6440 23480 6452
rect 23435 6412 23480 6440
rect 23474 6400 23480 6412
rect 23532 6400 23538 6452
rect 25240 6412 28764 6440
rect 15933 6375 15991 6381
rect 15933 6372 15945 6375
rect 11480 6344 13768 6372
rect 11480 6332 11486 6344
rect 10484 6310 10542 6316
rect 10484 6304 10496 6310
rect 10428 6276 10496 6304
rect 10530 6276 10542 6310
rect 10597 6307 10655 6313
rect 10597 6282 10609 6307
rect 10643 6282 10655 6307
rect 10689 6307 10747 6313
rect 10309 6267 10367 6273
rect 10484 6270 10542 6276
rect 9784 6208 10272 6236
rect 10594 6230 10600 6282
rect 10652 6230 10658 6282
rect 10689 6273 10701 6307
rect 10735 6304 10747 6307
rect 10962 6304 10968 6316
rect 10735 6276 10968 6304
rect 10735 6273 10747 6276
rect 10689 6267 10747 6273
rect 10962 6264 10968 6276
rect 11020 6264 11026 6316
rect 11146 6264 11152 6316
rect 11204 6304 11210 6316
rect 11517 6307 11575 6313
rect 11517 6304 11529 6307
rect 11204 6276 11529 6304
rect 11204 6264 11210 6276
rect 11517 6273 11529 6276
rect 11563 6273 11575 6307
rect 12710 6304 12716 6316
rect 12671 6276 12716 6304
rect 11517 6267 11575 6273
rect 12710 6264 12716 6276
rect 12768 6264 12774 6316
rect 13740 6313 13768 6344
rect 13832 6344 13952 6372
rect 14660 6344 15945 6372
rect 13832 6313 13860 6344
rect 13449 6307 13507 6313
rect 13449 6273 13461 6307
rect 13495 6273 13507 6307
rect 13449 6267 13507 6273
rect 13628 6307 13686 6313
rect 13628 6273 13640 6307
rect 13674 6273 13686 6307
rect 13628 6267 13686 6273
rect 13725 6307 13783 6313
rect 13725 6273 13737 6307
rect 13771 6273 13783 6307
rect 13725 6267 13783 6273
rect 13817 6307 13875 6313
rect 13817 6273 13829 6307
rect 13863 6273 13875 6307
rect 13817 6267 13875 6273
rect 8849 6199 8907 6205
rect 4856 6140 5028 6168
rect 5261 6171 5319 6177
rect 4856 6128 4862 6140
rect 5261 6137 5273 6171
rect 5307 6168 5319 6171
rect 5534 6168 5540 6180
rect 5307 6140 5540 6168
rect 5307 6137 5319 6140
rect 5261 6131 5319 6137
rect 5534 6128 5540 6140
rect 5592 6128 5598 6180
rect 1857 6103 1915 6109
rect 1857 6069 1869 6103
rect 1903 6100 1915 6103
rect 1946 6100 1952 6112
rect 1903 6072 1952 6100
rect 1903 6069 1915 6072
rect 1857 6063 1915 6069
rect 1946 6060 1952 6072
rect 2004 6060 2010 6112
rect 2958 6060 2964 6112
rect 3016 6100 3022 6112
rect 3145 6103 3203 6109
rect 3145 6100 3157 6103
rect 3016 6072 3157 6100
rect 3016 6060 3022 6072
rect 3145 6069 3157 6072
rect 3191 6100 3203 6103
rect 4706 6100 4712 6112
rect 3191 6072 4712 6100
rect 3191 6069 3203 6072
rect 3145 6063 3203 6069
rect 4706 6060 4712 6072
rect 4764 6060 4770 6112
rect 5442 6060 5448 6112
rect 5500 6100 5506 6112
rect 5721 6103 5779 6109
rect 5721 6100 5733 6103
rect 5500 6072 5733 6100
rect 5500 6060 5506 6072
rect 5721 6069 5733 6072
rect 5767 6069 5779 6103
rect 5721 6063 5779 6069
rect 6730 6060 6736 6112
rect 6788 6100 6794 6112
rect 6825 6103 6883 6109
rect 6825 6100 6837 6103
rect 6788 6072 6837 6100
rect 6788 6060 6794 6072
rect 6825 6069 6837 6072
rect 6871 6069 6883 6103
rect 7300 6100 7328 6199
rect 8864 6168 8892 6199
rect 7852 6140 8892 6168
rect 10244 6168 10272 6208
rect 12894 6196 12900 6248
rect 12952 6196 12958 6248
rect 12912 6168 12940 6196
rect 13464 6168 13492 6267
rect 10244 6140 13492 6168
rect 7852 6100 7880 6140
rect 7300 6072 7880 6100
rect 6825 6063 6883 6069
rect 8570 6060 8576 6112
rect 8628 6100 8634 6112
rect 9766 6100 9772 6112
rect 8628 6072 9772 6100
rect 8628 6060 8634 6072
rect 9766 6060 9772 6072
rect 9824 6060 9830 6112
rect 10962 6100 10968 6112
rect 10923 6072 10968 6100
rect 10962 6060 10968 6072
rect 11020 6060 11026 6112
rect 11146 6060 11152 6112
rect 11204 6100 11210 6112
rect 11701 6103 11759 6109
rect 11701 6100 11713 6103
rect 11204 6072 11713 6100
rect 11204 6060 11210 6072
rect 11701 6069 11713 6072
rect 11747 6069 11759 6103
rect 11701 6063 11759 6069
rect 11790 6060 11796 6112
rect 11848 6100 11854 6112
rect 12897 6103 12955 6109
rect 12897 6100 12909 6103
rect 11848 6072 12909 6100
rect 11848 6060 11854 6072
rect 12897 6069 12909 6072
rect 12943 6069 12955 6103
rect 13648 6100 13676 6267
rect 13740 6236 13768 6267
rect 14090 6264 14096 6316
rect 14148 6304 14154 6316
rect 14660 6304 14688 6344
rect 15933 6341 15945 6344
rect 15979 6341 15991 6375
rect 15933 6335 15991 6341
rect 18322 6332 18328 6384
rect 18380 6372 18386 6384
rect 18569 6375 18627 6381
rect 18569 6372 18581 6375
rect 18380 6344 18581 6372
rect 18380 6332 18386 6344
rect 18569 6341 18581 6344
rect 18615 6341 18627 6375
rect 18782 6372 18788 6384
rect 18743 6344 18788 6372
rect 18569 6335 18627 6341
rect 18782 6332 18788 6344
rect 18840 6332 18846 6384
rect 19058 6332 19064 6384
rect 19116 6372 19122 6384
rect 19116 6344 20576 6372
rect 19116 6332 19122 6344
rect 14148 6276 14688 6304
rect 14737 6307 14795 6313
rect 14148 6264 14154 6276
rect 14737 6273 14749 6307
rect 14783 6304 14795 6307
rect 14826 6304 14832 6316
rect 14783 6276 14832 6304
rect 14783 6273 14795 6276
rect 14737 6267 14795 6273
rect 14826 6264 14832 6276
rect 14884 6264 14890 6316
rect 14921 6307 14979 6313
rect 14921 6273 14933 6307
rect 14967 6304 14979 6307
rect 15102 6304 15108 6316
rect 14967 6276 15108 6304
rect 14967 6273 14979 6276
rect 14921 6267 14979 6273
rect 15102 6264 15108 6276
rect 15160 6264 15166 6316
rect 16942 6264 16948 6316
rect 17000 6304 17006 6316
rect 17405 6307 17463 6313
rect 17405 6304 17417 6307
rect 17000 6276 17417 6304
rect 17000 6264 17006 6276
rect 17405 6273 17417 6276
rect 17451 6273 17463 6307
rect 17405 6267 17463 6273
rect 17497 6307 17555 6313
rect 17497 6273 17509 6307
rect 17543 6304 17555 6307
rect 18690 6304 18696 6316
rect 17543 6276 18696 6304
rect 17543 6273 17555 6276
rect 17497 6267 17555 6273
rect 18690 6264 18696 6276
rect 18748 6264 18754 6316
rect 19610 6304 19616 6316
rect 19571 6276 19616 6304
rect 19610 6264 19616 6276
rect 19668 6264 19674 6316
rect 20254 6304 20260 6316
rect 20215 6276 20260 6304
rect 20254 6264 20260 6276
rect 20312 6264 20318 6316
rect 20548 6313 20576 6344
rect 21634 6332 21640 6384
rect 21692 6372 21698 6384
rect 25240 6372 25268 6412
rect 21692 6344 25268 6372
rect 21692 6332 21698 6344
rect 20533 6307 20591 6313
rect 20533 6273 20545 6307
rect 20579 6273 20591 6307
rect 21821 6307 21879 6313
rect 21821 6304 21833 6307
rect 20533 6267 20591 6273
rect 20916 6276 21833 6304
rect 16666 6236 16672 6248
rect 13740 6208 16672 6236
rect 16666 6196 16672 6208
rect 16724 6196 16730 6248
rect 17862 6236 17868 6248
rect 17823 6208 17868 6236
rect 17862 6196 17868 6208
rect 17920 6196 17926 6248
rect 14093 6171 14151 6177
rect 14093 6137 14105 6171
rect 14139 6168 14151 6171
rect 14182 6168 14188 6180
rect 14139 6140 14188 6168
rect 14139 6137 14151 6140
rect 14093 6131 14151 6137
rect 14182 6128 14188 6140
rect 14240 6128 14246 6180
rect 16408 6140 19334 6168
rect 16408 6112 16436 6140
rect 14553 6103 14611 6109
rect 14553 6100 14565 6103
rect 13648 6072 14565 6100
rect 12897 6063 12955 6069
rect 14553 6069 14565 6072
rect 14599 6069 14611 6103
rect 14553 6063 14611 6069
rect 16025 6103 16083 6109
rect 16025 6069 16037 6103
rect 16071 6100 16083 6103
rect 16390 6100 16396 6112
rect 16071 6072 16396 6100
rect 16071 6069 16083 6072
rect 16025 6063 16083 6069
rect 16390 6060 16396 6072
rect 16448 6060 16454 6112
rect 16758 6100 16764 6112
rect 16719 6072 16764 6100
rect 16758 6060 16764 6072
rect 16816 6060 16822 6112
rect 17218 6100 17224 6112
rect 17179 6072 17224 6100
rect 17218 6060 17224 6072
rect 17276 6060 17282 6112
rect 17402 6060 17408 6112
rect 17460 6100 17466 6112
rect 18417 6103 18475 6109
rect 18417 6100 18429 6103
rect 17460 6072 18429 6100
rect 17460 6060 17466 6072
rect 18417 6069 18429 6072
rect 18463 6069 18475 6103
rect 18598 6100 18604 6112
rect 18559 6072 18604 6100
rect 18417 6063 18475 6069
rect 18598 6060 18604 6072
rect 18656 6060 18662 6112
rect 19306 6100 19334 6140
rect 20916 6100 20944 6276
rect 21821 6273 21833 6276
rect 21867 6273 21879 6307
rect 22002 6304 22008 6316
rect 21963 6276 22008 6304
rect 21821 6267 21879 6273
rect 21836 6236 21864 6267
rect 22002 6264 22008 6276
rect 22060 6264 22066 6316
rect 22112 6313 22140 6344
rect 22097 6307 22155 6313
rect 22097 6273 22109 6307
rect 22143 6273 22155 6307
rect 22097 6267 22155 6273
rect 22186 6264 22192 6316
rect 22244 6304 22250 6316
rect 23382 6304 23388 6316
rect 22244 6276 22289 6304
rect 23343 6276 23388 6304
rect 22244 6264 22250 6276
rect 23382 6264 23388 6276
rect 23440 6264 23446 6316
rect 23566 6304 23572 6316
rect 23527 6276 23572 6304
rect 23566 6264 23572 6276
rect 23624 6264 23630 6316
rect 24026 6304 24032 6316
rect 23987 6276 24032 6304
rect 24026 6264 24032 6276
rect 24084 6264 24090 6316
rect 24210 6304 24216 6316
rect 24171 6276 24216 6304
rect 24210 6264 24216 6276
rect 24268 6264 24274 6316
rect 24670 6264 24676 6316
rect 24728 6304 24734 6316
rect 25240 6313 25268 6344
rect 25516 6344 27936 6372
rect 25516 6316 25544 6344
rect 25087 6307 25145 6313
rect 25087 6304 25099 6307
rect 24728 6276 25099 6304
rect 24728 6264 24734 6276
rect 25087 6273 25099 6276
rect 25133 6273 25145 6307
rect 25087 6267 25145 6273
rect 25225 6307 25283 6313
rect 25225 6273 25237 6307
rect 25271 6273 25283 6307
rect 25225 6267 25283 6273
rect 25317 6307 25375 6313
rect 25317 6273 25329 6307
rect 25363 6279 25452 6307
rect 25363 6273 25375 6279
rect 25317 6267 25375 6273
rect 24762 6236 24768 6248
rect 21836 6208 24768 6236
rect 24762 6196 24768 6208
rect 24820 6196 24826 6248
rect 20990 6128 20996 6180
rect 21048 6168 21054 6180
rect 24026 6168 24032 6180
rect 21048 6140 24032 6168
rect 21048 6128 21054 6140
rect 24026 6128 24032 6140
rect 24084 6128 24090 6180
rect 24397 6171 24455 6177
rect 24397 6137 24409 6171
rect 24443 6168 24455 6171
rect 24443 6140 25084 6168
rect 24443 6137 24455 6140
rect 24397 6131 24455 6137
rect 19306 6072 20944 6100
rect 21269 6103 21327 6109
rect 21269 6069 21281 6103
rect 21315 6100 21327 6103
rect 22094 6100 22100 6112
rect 21315 6072 22100 6100
rect 21315 6069 21327 6072
rect 21269 6063 21327 6069
rect 22094 6060 22100 6072
rect 22152 6060 22158 6112
rect 22462 6100 22468 6112
rect 22423 6072 22468 6100
rect 22462 6060 22468 6072
rect 22520 6060 22526 6112
rect 24857 6103 24915 6109
rect 24857 6069 24869 6103
rect 24903 6100 24915 6103
rect 24946 6100 24952 6112
rect 24903 6072 24952 6100
rect 24903 6069 24915 6072
rect 24857 6063 24915 6069
rect 24946 6060 24952 6072
rect 25004 6060 25010 6112
rect 25056 6100 25084 6140
rect 25424 6100 25452 6279
rect 25498 6264 25504 6316
rect 25556 6304 25562 6316
rect 25556 6276 25601 6304
rect 25556 6264 25562 6276
rect 25866 6264 25872 6316
rect 25924 6304 25930 6316
rect 25961 6307 26019 6313
rect 25961 6304 25973 6307
rect 25924 6276 25973 6304
rect 25924 6264 25930 6276
rect 25961 6273 25973 6276
rect 26007 6273 26019 6307
rect 26142 6304 26148 6316
rect 26103 6276 26148 6304
rect 25961 6267 26019 6273
rect 26142 6264 26148 6276
rect 26200 6264 26206 6316
rect 26234 6264 26240 6316
rect 26292 6304 26298 6316
rect 27908 6313 27936 6344
rect 27249 6307 27307 6313
rect 27249 6304 27261 6307
rect 26292 6276 27261 6304
rect 26292 6264 26298 6276
rect 27249 6273 27261 6276
rect 27295 6273 27307 6307
rect 27249 6267 27307 6273
rect 27893 6307 27951 6313
rect 27893 6273 27905 6307
rect 27939 6273 27951 6307
rect 28074 6304 28080 6316
rect 28035 6276 28080 6304
rect 27893 6267 27951 6273
rect 27908 6236 27936 6267
rect 28074 6264 28080 6276
rect 28132 6264 28138 6316
rect 28184 6313 28212 6412
rect 28736 6372 28764 6412
rect 28810 6400 28816 6452
rect 28868 6440 28874 6452
rect 30745 6443 30803 6449
rect 28868 6412 30696 6440
rect 28868 6400 28874 6412
rect 30374 6372 30380 6384
rect 28736 6344 29592 6372
rect 30287 6344 30380 6372
rect 28169 6307 28227 6313
rect 28169 6273 28181 6307
rect 28215 6273 28227 6307
rect 28169 6267 28227 6273
rect 28281 6307 28339 6313
rect 28281 6273 28293 6307
rect 28327 6304 28396 6307
rect 28810 6304 28816 6316
rect 28327 6279 28816 6304
rect 28327 6273 28339 6279
rect 28368 6276 28816 6279
rect 28281 6267 28339 6273
rect 28810 6264 28816 6276
rect 28868 6264 28874 6316
rect 29273 6307 29331 6313
rect 29273 6273 29285 6307
rect 29319 6273 29331 6307
rect 29454 6304 29460 6316
rect 29415 6276 29460 6304
rect 29273 6267 29331 6273
rect 29288 6236 29316 6267
rect 29454 6264 29460 6276
rect 29512 6264 29518 6316
rect 29564 6313 29592 6344
rect 30374 6332 30380 6344
rect 30432 6332 30438 6384
rect 30466 6332 30472 6384
rect 30524 6372 30530 6384
rect 30577 6375 30635 6381
rect 30577 6372 30589 6375
rect 30524 6344 30589 6372
rect 30524 6332 30530 6344
rect 30577 6341 30589 6344
rect 30623 6341 30635 6375
rect 30668 6372 30696 6412
rect 30745 6409 30757 6443
rect 30791 6440 30803 6443
rect 31938 6440 31944 6452
rect 30791 6412 31944 6440
rect 30791 6409 30803 6412
rect 30745 6403 30803 6409
rect 31938 6400 31944 6412
rect 31996 6400 32002 6452
rect 34422 6440 34428 6452
rect 32048 6412 34428 6440
rect 31662 6372 31668 6384
rect 30668 6344 31668 6372
rect 30577 6335 30635 6341
rect 29549 6307 29607 6313
rect 29549 6273 29561 6307
rect 29595 6273 29607 6307
rect 29549 6267 29607 6273
rect 29638 6264 29644 6316
rect 29696 6304 29702 6316
rect 29696 6276 29741 6304
rect 29696 6264 29702 6276
rect 27908 6208 29316 6236
rect 26145 6171 26203 6177
rect 26145 6137 26157 6171
rect 26191 6168 26203 6171
rect 27246 6168 27252 6180
rect 26191 6140 27252 6168
rect 26191 6137 26203 6140
rect 26145 6131 26203 6137
rect 27246 6128 27252 6140
rect 27304 6128 27310 6180
rect 27430 6168 27436 6180
rect 27391 6140 27436 6168
rect 27430 6128 27436 6140
rect 27488 6128 27494 6180
rect 30392 6168 30420 6332
rect 30592 6304 30620 6335
rect 31662 6332 31668 6344
rect 31720 6332 31726 6384
rect 32048 6304 32076 6412
rect 34422 6400 34428 6412
rect 34480 6400 34486 6452
rect 34882 6400 34888 6452
rect 34940 6440 34946 6452
rect 35437 6443 35495 6449
rect 35437 6440 35449 6443
rect 34940 6412 35449 6440
rect 34940 6400 34946 6412
rect 35437 6409 35449 6412
rect 35483 6440 35495 6443
rect 36998 6440 37004 6452
rect 35483 6412 37004 6440
rect 35483 6409 35495 6412
rect 35437 6403 35495 6409
rect 36998 6400 37004 6412
rect 37056 6400 37062 6452
rect 37461 6443 37519 6449
rect 37461 6409 37473 6443
rect 37507 6440 37519 6443
rect 37507 6412 39804 6440
rect 37507 6409 37519 6412
rect 37461 6403 37519 6409
rect 32125 6375 32183 6381
rect 32125 6341 32137 6375
rect 32171 6372 32183 6375
rect 32306 6372 32312 6384
rect 32171 6344 32312 6372
rect 32171 6341 32183 6344
rect 32125 6335 32183 6341
rect 32306 6332 32312 6344
rect 32364 6332 32370 6384
rect 32950 6332 32956 6384
rect 33008 6372 33014 6384
rect 33045 6375 33103 6381
rect 33045 6372 33057 6375
rect 33008 6344 33057 6372
rect 33008 6332 33014 6344
rect 33045 6341 33057 6344
rect 33091 6341 33103 6375
rect 33045 6335 33103 6341
rect 33134 6332 33140 6384
rect 33192 6372 33198 6384
rect 33229 6375 33287 6381
rect 33229 6372 33241 6375
rect 33192 6344 33241 6372
rect 33192 6332 33198 6344
rect 33229 6341 33241 6344
rect 33275 6372 33287 6375
rect 33781 6375 33839 6381
rect 33781 6372 33793 6375
rect 33275 6344 33793 6372
rect 33275 6341 33287 6344
rect 33229 6335 33287 6341
rect 33781 6341 33793 6344
rect 33827 6341 33839 6375
rect 33781 6335 33839 6341
rect 33870 6332 33876 6384
rect 33928 6372 33934 6384
rect 38470 6372 38476 6384
rect 33928 6344 38476 6372
rect 33928 6332 33934 6344
rect 32217 6307 32275 6313
rect 32217 6304 32229 6307
rect 30592 6276 32229 6304
rect 32217 6273 32229 6276
rect 32263 6273 32275 6307
rect 32398 6304 32404 6316
rect 32359 6276 32404 6304
rect 32217 6267 32275 6273
rect 32398 6264 32404 6276
rect 32456 6264 32462 6316
rect 34422 6304 34428 6316
rect 34383 6276 34428 6304
rect 34422 6264 34428 6276
rect 34480 6264 34486 6316
rect 34606 6304 34612 6316
rect 34567 6276 34612 6304
rect 34606 6264 34612 6276
rect 34664 6264 34670 6316
rect 35253 6307 35311 6313
rect 35253 6304 35265 6307
rect 34992 6276 35265 6304
rect 32493 6239 32551 6245
rect 32493 6205 32505 6239
rect 32539 6236 32551 6239
rect 32582 6236 32588 6248
rect 32539 6208 32588 6236
rect 32539 6205 32551 6208
rect 32493 6199 32551 6205
rect 32582 6196 32588 6208
rect 32640 6196 32646 6248
rect 34333 6239 34391 6245
rect 34333 6205 34345 6239
rect 34379 6236 34391 6239
rect 34882 6236 34888 6248
rect 34379 6208 34888 6236
rect 34379 6205 34391 6208
rect 34333 6199 34391 6205
rect 34882 6196 34888 6208
rect 34940 6196 34946 6248
rect 34992 6168 35020 6276
rect 35253 6273 35265 6276
rect 35299 6273 35311 6307
rect 35253 6267 35311 6273
rect 35529 6307 35587 6313
rect 35529 6273 35541 6307
rect 35575 6304 35587 6307
rect 35802 6304 35808 6316
rect 35575 6276 35808 6304
rect 35575 6273 35587 6276
rect 35529 6267 35587 6273
rect 35802 6264 35808 6276
rect 35860 6264 35866 6316
rect 35894 6264 35900 6316
rect 35952 6304 35958 6316
rect 37568 6313 37596 6344
rect 38470 6332 38476 6344
rect 38528 6332 38534 6384
rect 39776 6381 39804 6412
rect 40678 6400 40684 6452
rect 40736 6440 40742 6452
rect 40773 6443 40831 6449
rect 40773 6440 40785 6443
rect 40736 6412 40785 6440
rect 40736 6400 40742 6412
rect 40773 6409 40785 6412
rect 40819 6409 40831 6443
rect 40773 6403 40831 6409
rect 40862 6400 40868 6452
rect 40920 6440 40926 6452
rect 46198 6440 46204 6452
rect 40920 6412 46204 6440
rect 40920 6400 40926 6412
rect 46198 6400 46204 6412
rect 46256 6400 46262 6452
rect 47673 6443 47731 6449
rect 47673 6409 47685 6443
rect 47719 6440 47731 6443
rect 49970 6440 49976 6452
rect 47719 6412 49976 6440
rect 47719 6409 47731 6412
rect 47673 6403 47731 6409
rect 49970 6400 49976 6412
rect 50028 6400 50034 6452
rect 50522 6440 50528 6452
rect 50483 6412 50528 6440
rect 50522 6400 50528 6412
rect 50580 6400 50586 6452
rect 57885 6443 57943 6449
rect 57885 6440 57897 6443
rect 51552 6412 55444 6440
rect 39761 6375 39819 6381
rect 39761 6341 39773 6375
rect 39807 6341 39819 6375
rect 39761 6335 39819 6341
rect 41782 6332 41788 6384
rect 41840 6372 41846 6384
rect 42981 6375 43039 6381
rect 42981 6372 42993 6375
rect 41840 6344 42993 6372
rect 41840 6332 41846 6344
rect 42981 6341 42993 6344
rect 43027 6341 43039 6375
rect 42981 6335 43039 6341
rect 36357 6307 36415 6313
rect 36357 6304 36369 6307
rect 35952 6276 36369 6304
rect 35952 6264 35958 6276
rect 36357 6273 36369 6276
rect 36403 6273 36415 6307
rect 36357 6267 36415 6273
rect 37461 6307 37519 6313
rect 37461 6273 37473 6307
rect 37507 6273 37519 6307
rect 37461 6267 37519 6273
rect 37553 6307 37611 6313
rect 37553 6273 37565 6307
rect 37599 6273 37611 6307
rect 37553 6267 37611 6273
rect 37476 6236 37504 6267
rect 37734 6264 37740 6316
rect 37792 6304 37798 6316
rect 37792 6276 38424 6304
rect 37792 6264 37798 6276
rect 38286 6236 38292 6248
rect 35268 6208 37504 6236
rect 38247 6208 38292 6236
rect 35268 6177 35296 6208
rect 38286 6196 38292 6208
rect 38344 6196 38350 6248
rect 38396 6236 38424 6276
rect 38654 6264 38660 6316
rect 38712 6264 38718 6316
rect 40218 6264 40224 6316
rect 40276 6304 40282 6316
rect 40589 6307 40647 6313
rect 40589 6304 40601 6307
rect 40276 6276 40601 6304
rect 40276 6264 40282 6276
rect 40589 6273 40601 6276
rect 40635 6273 40647 6307
rect 40589 6267 40647 6273
rect 41509 6307 41567 6313
rect 41509 6273 41521 6307
rect 41555 6304 41567 6307
rect 41598 6304 41604 6316
rect 41555 6276 41604 6304
rect 41555 6273 41567 6276
rect 41509 6267 41567 6273
rect 41598 6264 41604 6276
rect 41656 6264 41662 6316
rect 41690 6264 41696 6316
rect 41748 6304 41754 6316
rect 41748 6276 41793 6304
rect 41748 6264 41754 6276
rect 39298 6236 39304 6248
rect 38396 6208 39304 6236
rect 39298 6196 39304 6208
rect 39356 6196 39362 6248
rect 40034 6236 40040 6248
rect 39995 6208 40040 6236
rect 40034 6196 40040 6208
rect 40092 6196 40098 6248
rect 41414 6196 41420 6248
rect 41472 6236 41478 6248
rect 41785 6239 41843 6245
rect 41785 6236 41797 6239
rect 41472 6208 41797 6236
rect 41472 6196 41478 6208
rect 41785 6205 41797 6208
rect 41831 6236 41843 6239
rect 42610 6236 42616 6248
rect 41831 6208 42616 6236
rect 41831 6205 41843 6208
rect 41785 6199 41843 6205
rect 42610 6196 42616 6208
rect 42668 6196 42674 6248
rect 30392 6140 35020 6168
rect 35253 6171 35311 6177
rect 35253 6137 35265 6171
rect 35299 6137 35311 6171
rect 35253 6131 35311 6137
rect 35894 6128 35900 6180
rect 35952 6168 35958 6180
rect 36078 6168 36084 6180
rect 35952 6140 36084 6168
rect 35952 6128 35958 6140
rect 36078 6128 36084 6140
rect 36136 6168 36142 6180
rect 36906 6168 36912 6180
rect 36136 6140 36912 6168
rect 36136 6128 36142 6140
rect 36906 6128 36912 6140
rect 36964 6128 36970 6180
rect 36998 6128 37004 6180
rect 37056 6168 37062 6180
rect 38010 6168 38016 6180
rect 37056 6140 38016 6168
rect 37056 6128 37062 6140
rect 38010 6128 38016 6140
rect 38068 6128 38074 6180
rect 40126 6128 40132 6180
rect 40184 6168 40190 6180
rect 42429 6171 42487 6177
rect 42429 6168 42441 6171
rect 40184 6140 42441 6168
rect 40184 6128 40190 6140
rect 42429 6137 42441 6140
rect 42475 6137 42487 6171
rect 42996 6168 43024 6335
rect 44082 6332 44088 6384
rect 44140 6372 44146 6384
rect 46937 6375 46995 6381
rect 44140 6344 45416 6372
rect 44140 6332 44146 6344
rect 45388 6316 45416 6344
rect 46937 6341 46949 6375
rect 46983 6372 46995 6375
rect 51442 6372 51448 6384
rect 46983 6344 47978 6372
rect 51046 6344 51448 6372
rect 46983 6341 46995 6344
rect 46937 6335 46995 6341
rect 45094 6264 45100 6316
rect 45152 6313 45158 6316
rect 45152 6304 45164 6313
rect 45152 6276 45197 6304
rect 45152 6267 45164 6276
rect 45152 6264 45158 6267
rect 45370 6264 45376 6316
rect 45428 6304 45434 6316
rect 46842 6304 46848 6316
rect 45428 6276 45521 6304
rect 46803 6276 46848 6304
rect 45428 6264 45434 6276
rect 46842 6264 46848 6276
rect 46900 6264 46906 6316
rect 50062 6304 50068 6316
rect 50023 6276 50068 6304
rect 50062 6264 50068 6276
rect 50120 6264 50126 6316
rect 50706 6304 50712 6316
rect 50667 6276 50712 6304
rect 50706 6264 50712 6276
rect 50764 6264 50770 6316
rect 49145 6239 49203 6245
rect 49145 6205 49157 6239
rect 49191 6236 49203 6239
rect 49191 6208 49372 6236
rect 49191 6205 49203 6208
rect 49145 6199 49203 6205
rect 43993 6171 44051 6177
rect 43993 6168 44005 6171
rect 42996 6140 44005 6168
rect 42429 6131 42487 6137
rect 43993 6137 44005 6140
rect 44039 6137 44051 6171
rect 45830 6168 45836 6180
rect 45791 6140 45836 6168
rect 43993 6131 44051 6137
rect 45830 6128 45836 6140
rect 45888 6128 45894 6180
rect 49344 6168 49372 6208
rect 49418 6196 49424 6248
rect 49476 6236 49482 6248
rect 51046 6236 51074 6344
rect 51442 6332 51448 6344
rect 51500 6332 51506 6384
rect 49476 6208 51074 6236
rect 49476 6196 49482 6208
rect 51169 6171 51227 6177
rect 51169 6168 51181 6171
rect 49344 6140 51181 6168
rect 51169 6137 51181 6140
rect 51215 6137 51227 6171
rect 51169 6131 51227 6137
rect 25056 6072 25452 6100
rect 28537 6103 28595 6109
rect 28537 6069 28549 6103
rect 28583 6100 28595 6103
rect 28718 6100 28724 6112
rect 28583 6072 28724 6100
rect 28583 6069 28595 6072
rect 28537 6063 28595 6069
rect 28718 6060 28724 6072
rect 28776 6060 28782 6112
rect 29914 6100 29920 6112
rect 29875 6072 29920 6100
rect 29914 6060 29920 6072
rect 29972 6060 29978 6112
rect 30558 6100 30564 6112
rect 30519 6072 30564 6100
rect 30558 6060 30564 6072
rect 30616 6060 30622 6112
rect 31202 6100 31208 6112
rect 31163 6072 31208 6100
rect 31202 6060 31208 6072
rect 31260 6060 31266 6112
rect 32585 6103 32643 6109
rect 32585 6069 32597 6103
rect 32631 6100 32643 6103
rect 33042 6100 33048 6112
rect 32631 6072 33048 6100
rect 32631 6069 32643 6072
rect 32585 6063 32643 6069
rect 33042 6060 33048 6072
rect 33100 6060 33106 6112
rect 34793 6103 34851 6109
rect 34793 6069 34805 6103
rect 34839 6100 34851 6103
rect 35158 6100 35164 6112
rect 34839 6072 35164 6100
rect 34839 6069 34851 6072
rect 34793 6063 34851 6069
rect 35158 6060 35164 6072
rect 35216 6060 35222 6112
rect 36541 6103 36599 6109
rect 36541 6069 36553 6103
rect 36587 6100 36599 6103
rect 40770 6100 40776 6112
rect 36587 6072 40776 6100
rect 36587 6069 36599 6072
rect 36541 6063 36599 6069
rect 40770 6060 40776 6072
rect 40828 6060 40834 6112
rect 41322 6100 41328 6112
rect 41283 6072 41328 6100
rect 41322 6060 41328 6072
rect 41380 6060 41386 6112
rect 42610 6060 42616 6112
rect 42668 6100 42674 6112
rect 48038 6100 48044 6112
rect 42668 6072 48044 6100
rect 42668 6060 42674 6072
rect 48038 6060 48044 6072
rect 48096 6060 48102 6112
rect 49326 6060 49332 6112
rect 49384 6100 49390 6112
rect 49881 6103 49939 6109
rect 49881 6100 49893 6103
rect 49384 6072 49893 6100
rect 49384 6060 49390 6072
rect 49881 6069 49893 6072
rect 49927 6069 49939 6103
rect 49881 6063 49939 6069
rect 49970 6060 49976 6112
rect 50028 6100 50034 6112
rect 51552 6100 51580 6412
rect 55416 6316 55444 6412
rect 55508 6412 57897 6440
rect 51905 6307 51963 6313
rect 51905 6273 51917 6307
rect 51951 6304 51963 6307
rect 52638 6304 52644 6316
rect 51951 6276 52644 6304
rect 51951 6273 51963 6276
rect 51905 6267 51963 6273
rect 52638 6264 52644 6276
rect 52696 6264 52702 6316
rect 53837 6308 53895 6313
rect 53837 6307 53972 6308
rect 53837 6273 53849 6307
rect 53883 6304 53972 6307
rect 55398 6304 55404 6316
rect 53883 6280 55260 6304
rect 53883 6273 53895 6280
rect 53944 6276 55260 6280
rect 55311 6276 55404 6304
rect 53837 6267 53895 6273
rect 52178 6196 52184 6248
rect 52236 6236 52242 6248
rect 52236 6208 53512 6236
rect 52236 6196 52242 6208
rect 53098 6100 53104 6112
rect 50028 6072 51580 6100
rect 53059 6072 53104 6100
rect 50028 6060 50034 6072
rect 53098 6060 53104 6072
rect 53156 6060 53162 6112
rect 53484 6100 53512 6208
rect 54110 6196 54116 6248
rect 54168 6236 54174 6248
rect 55122 6236 55128 6248
rect 54168 6208 54261 6236
rect 55083 6208 55128 6236
rect 54168 6196 54174 6208
rect 55122 6196 55128 6208
rect 55180 6196 55186 6248
rect 55232 6236 55260 6276
rect 55398 6264 55404 6276
rect 55456 6264 55462 6316
rect 55508 6236 55536 6412
rect 57885 6409 57897 6412
rect 57931 6409 57943 6443
rect 57885 6403 57943 6409
rect 56042 6332 56048 6384
rect 56100 6372 56106 6384
rect 56100 6344 58112 6372
rect 56100 6332 56106 6344
rect 55582 6264 55588 6316
rect 55640 6304 55646 6316
rect 56137 6307 56195 6313
rect 56137 6304 56149 6307
rect 55640 6276 56149 6304
rect 55640 6264 55646 6276
rect 56137 6273 56149 6276
rect 56183 6273 56195 6307
rect 56137 6267 56195 6273
rect 56318 6264 56324 6316
rect 56376 6304 56382 6316
rect 58084 6313 58112 6344
rect 56965 6307 57023 6313
rect 56965 6304 56977 6307
rect 56376 6276 56977 6304
rect 56376 6264 56382 6276
rect 56965 6273 56977 6276
rect 57011 6273 57023 6307
rect 56965 6267 57023 6273
rect 58069 6307 58127 6313
rect 58069 6273 58081 6307
rect 58115 6273 58127 6307
rect 58069 6267 58127 6273
rect 55232 6208 55536 6236
rect 55861 6239 55919 6245
rect 55861 6205 55873 6239
rect 55907 6236 55919 6239
rect 55950 6236 55956 6248
rect 55907 6208 55956 6236
rect 55907 6205 55919 6208
rect 55861 6199 55919 6205
rect 55950 6196 55956 6208
rect 56008 6196 56014 6248
rect 54128 6168 54156 6196
rect 56781 6171 56839 6177
rect 56781 6168 56793 6171
rect 54128 6140 56793 6168
rect 54128 6100 54156 6140
rect 56781 6137 56793 6140
rect 56827 6137 56839 6171
rect 56781 6131 56839 6137
rect 53484 6072 54156 6100
rect 55398 6060 55404 6112
rect 55456 6100 55462 6112
rect 55953 6103 56011 6109
rect 55953 6100 55965 6103
rect 55456 6072 55965 6100
rect 55456 6060 55462 6072
rect 55953 6069 55965 6072
rect 55999 6100 56011 6103
rect 56134 6100 56140 6112
rect 55999 6072 56140 6100
rect 55999 6069 56011 6072
rect 55953 6063 56011 6069
rect 56134 6060 56140 6072
rect 56192 6060 56198 6112
rect 56318 6100 56324 6112
rect 56279 6072 56324 6100
rect 56318 6060 56324 6072
rect 56376 6060 56382 6112
rect 1104 6010 58880 6032
rect 1104 5958 8174 6010
rect 8226 5958 8238 6010
rect 8290 5958 8302 6010
rect 8354 5958 8366 6010
rect 8418 5958 8430 6010
rect 8482 5958 22622 6010
rect 22674 5958 22686 6010
rect 22738 5958 22750 6010
rect 22802 5958 22814 6010
rect 22866 5958 22878 6010
rect 22930 5958 37070 6010
rect 37122 5958 37134 6010
rect 37186 5958 37198 6010
rect 37250 5958 37262 6010
rect 37314 5958 37326 6010
rect 37378 5958 51518 6010
rect 51570 5958 51582 6010
rect 51634 5958 51646 6010
rect 51698 5958 51710 6010
rect 51762 5958 51774 6010
rect 51826 5958 58880 6010
rect 1104 5936 58880 5958
rect 1765 5899 1823 5905
rect 1765 5865 1777 5899
rect 1811 5896 1823 5899
rect 1854 5896 1860 5908
rect 1811 5868 1860 5896
rect 1811 5865 1823 5868
rect 1765 5859 1823 5865
rect 1854 5856 1860 5868
rect 1912 5856 1918 5908
rect 2409 5899 2467 5905
rect 2409 5865 2421 5899
rect 2455 5896 2467 5899
rect 3878 5896 3884 5908
rect 2455 5868 3884 5896
rect 2455 5865 2467 5868
rect 2409 5859 2467 5865
rect 3878 5856 3884 5868
rect 3936 5856 3942 5908
rect 4706 5856 4712 5908
rect 4764 5896 4770 5908
rect 7834 5896 7840 5908
rect 4764 5868 7840 5896
rect 4764 5856 4770 5868
rect 7834 5856 7840 5868
rect 7892 5856 7898 5908
rect 8205 5899 8263 5905
rect 8205 5865 8217 5899
rect 8251 5896 8263 5899
rect 9766 5896 9772 5908
rect 8251 5868 9772 5896
rect 8251 5865 8263 5868
rect 8205 5859 8263 5865
rect 9766 5856 9772 5868
rect 9824 5856 9830 5908
rect 9858 5856 9864 5908
rect 9916 5896 9922 5908
rect 10045 5899 10103 5905
rect 10045 5896 10057 5899
rect 9916 5868 10057 5896
rect 9916 5856 9922 5868
rect 10045 5865 10057 5868
rect 10091 5865 10103 5899
rect 13722 5896 13728 5908
rect 10045 5859 10103 5865
rect 10704 5868 13728 5896
rect 3237 5831 3295 5837
rect 3237 5797 3249 5831
rect 3283 5828 3295 5831
rect 4246 5828 4252 5840
rect 3283 5800 4252 5828
rect 3283 5797 3295 5800
rect 3237 5791 3295 5797
rect 4246 5788 4252 5800
rect 4304 5788 4310 5840
rect 6638 5828 6644 5840
rect 6551 5800 6644 5828
rect 6638 5788 6644 5800
rect 6696 5828 6702 5840
rect 8570 5828 8576 5840
rect 6696 5800 8576 5828
rect 6696 5788 6702 5800
rect 8570 5788 8576 5800
rect 8628 5788 8634 5840
rect 9122 5788 9128 5840
rect 9180 5828 9186 5840
rect 10704 5828 10732 5868
rect 13722 5856 13728 5868
rect 13780 5856 13786 5908
rect 16758 5896 16764 5908
rect 14108 5868 16764 5896
rect 9180 5800 10732 5828
rect 9180 5788 9186 5800
rect 3050 5760 3056 5772
rect 1596 5732 3056 5760
rect 1596 5701 1624 5732
rect 3050 5720 3056 5732
rect 3108 5720 3114 5772
rect 6362 5720 6368 5772
rect 6420 5760 6426 5772
rect 6420 5732 6914 5760
rect 6420 5720 6426 5732
rect 1581 5695 1639 5701
rect 1581 5661 1593 5695
rect 1627 5661 1639 5695
rect 2222 5692 2228 5704
rect 2183 5664 2228 5692
rect 1581 5655 1639 5661
rect 2222 5652 2228 5664
rect 2280 5652 2286 5704
rect 2774 5652 2780 5704
rect 2832 5692 2838 5704
rect 2869 5695 2927 5701
rect 2869 5692 2881 5695
rect 2832 5664 2881 5692
rect 2832 5652 2838 5664
rect 2869 5661 2881 5664
rect 2915 5692 2927 5695
rect 3418 5692 3424 5704
rect 2915 5664 3424 5692
rect 2915 5661 2927 5664
rect 2869 5655 2927 5661
rect 3418 5652 3424 5664
rect 3476 5652 3482 5704
rect 3694 5652 3700 5704
rect 3752 5692 3758 5704
rect 3970 5701 3976 5704
rect 3789 5695 3847 5701
rect 3789 5692 3801 5695
rect 3752 5664 3801 5692
rect 3752 5652 3758 5664
rect 3789 5661 3801 5664
rect 3835 5661 3847 5695
rect 3968 5692 3976 5701
rect 3931 5664 3976 5692
rect 3789 5655 3847 5661
rect 3968 5655 3976 5664
rect 3970 5652 3976 5655
rect 4028 5652 4034 5704
rect 4068 5689 4126 5695
rect 4068 5655 4080 5689
rect 4114 5655 4126 5689
rect 4068 5649 4126 5655
rect 4154 5652 4160 5704
rect 4212 5692 4218 5704
rect 5261 5695 5319 5701
rect 4212 5664 4257 5692
rect 4212 5652 4218 5664
rect 5261 5661 5273 5695
rect 5307 5692 5319 5695
rect 5350 5692 5356 5704
rect 5307 5664 5356 5692
rect 5307 5661 5319 5664
rect 5261 5655 5319 5661
rect 5350 5652 5356 5664
rect 5408 5652 5414 5704
rect 5534 5701 5540 5704
rect 5528 5692 5540 5701
rect 5495 5664 5540 5692
rect 5528 5655 5540 5664
rect 5534 5652 5540 5655
rect 5592 5652 5598 5704
rect 3050 5624 3056 5636
rect 3011 5596 3056 5624
rect 3050 5584 3056 5596
rect 3108 5584 3114 5636
rect 4080 5568 4108 5649
rect 5166 5584 5172 5636
rect 5224 5624 5230 5636
rect 5902 5624 5908 5636
rect 5224 5596 5908 5624
rect 5224 5584 5230 5596
rect 5902 5584 5908 5596
rect 5960 5584 5966 5636
rect 6886 5624 6914 5732
rect 10226 5720 10232 5772
rect 10284 5760 10290 5772
rect 14108 5769 14136 5868
rect 16758 5856 16764 5868
rect 16816 5856 16822 5908
rect 17494 5896 17500 5908
rect 17455 5868 17500 5896
rect 17494 5856 17500 5868
rect 17552 5856 17558 5908
rect 18230 5856 18236 5908
rect 18288 5896 18294 5908
rect 18782 5896 18788 5908
rect 18288 5868 18788 5896
rect 18288 5856 18294 5868
rect 18782 5856 18788 5868
rect 18840 5856 18846 5908
rect 19613 5899 19671 5905
rect 19613 5865 19625 5899
rect 19659 5896 19671 5899
rect 22002 5896 22008 5908
rect 19659 5868 22008 5896
rect 19659 5865 19671 5868
rect 19613 5859 19671 5865
rect 22002 5856 22008 5868
rect 22060 5856 22066 5908
rect 24210 5856 24216 5908
rect 24268 5896 24274 5908
rect 26053 5899 26111 5905
rect 26053 5896 26065 5899
rect 24268 5868 26065 5896
rect 24268 5856 24274 5868
rect 26053 5865 26065 5868
rect 26099 5865 26111 5899
rect 26053 5859 26111 5865
rect 27157 5899 27215 5905
rect 27157 5865 27169 5899
rect 27203 5896 27215 5899
rect 28074 5896 28080 5908
rect 27203 5868 28080 5896
rect 27203 5865 27215 5868
rect 27157 5859 27215 5865
rect 28074 5856 28080 5868
rect 28132 5856 28138 5908
rect 29454 5856 29460 5908
rect 29512 5896 29518 5908
rect 29917 5899 29975 5905
rect 29917 5896 29929 5899
rect 29512 5868 29929 5896
rect 29512 5856 29518 5868
rect 29917 5865 29929 5868
rect 29963 5865 29975 5899
rect 29917 5859 29975 5865
rect 32306 5856 32312 5908
rect 32364 5896 32370 5908
rect 33137 5899 33195 5905
rect 33137 5896 33149 5899
rect 32364 5868 33149 5896
rect 32364 5856 32370 5868
rect 33137 5865 33149 5868
rect 33183 5865 33195 5899
rect 33778 5896 33784 5908
rect 33739 5868 33784 5896
rect 33137 5859 33195 5865
rect 33778 5856 33784 5868
rect 33836 5856 33842 5908
rect 34606 5856 34612 5908
rect 34664 5896 34670 5908
rect 34701 5899 34759 5905
rect 34701 5896 34713 5899
rect 34664 5868 34713 5896
rect 34664 5856 34670 5868
rect 34701 5865 34713 5868
rect 34747 5865 34759 5899
rect 34701 5859 34759 5865
rect 35621 5899 35679 5905
rect 35621 5865 35633 5899
rect 35667 5896 35679 5899
rect 36814 5896 36820 5908
rect 35667 5868 36820 5896
rect 35667 5865 35679 5868
rect 35621 5859 35679 5865
rect 36814 5856 36820 5868
rect 36872 5856 36878 5908
rect 36906 5856 36912 5908
rect 36964 5896 36970 5908
rect 41322 5905 41328 5908
rect 41312 5899 41328 5905
rect 36964 5868 41184 5896
rect 36964 5856 36970 5868
rect 15102 5788 15108 5840
rect 15160 5828 15166 5840
rect 20990 5828 20996 5840
rect 15160 5800 20996 5828
rect 15160 5788 15166 5800
rect 20990 5788 20996 5800
rect 21048 5788 21054 5840
rect 29730 5788 29736 5840
rect 29788 5828 29794 5840
rect 30466 5828 30472 5840
rect 29788 5800 30472 5828
rect 29788 5788 29794 5800
rect 30466 5788 30472 5800
rect 30524 5828 30530 5840
rect 31297 5831 31355 5837
rect 31297 5828 31309 5831
rect 30524 5800 31309 5828
rect 30524 5788 30530 5800
rect 31297 5797 31309 5800
rect 31343 5797 31355 5831
rect 31297 5791 31355 5797
rect 33226 5788 33232 5840
rect 33284 5828 33290 5840
rect 36078 5828 36084 5840
rect 33284 5800 36084 5828
rect 33284 5788 33290 5800
rect 36078 5788 36084 5800
rect 36136 5788 36142 5840
rect 37642 5788 37648 5840
rect 37700 5828 37706 5840
rect 37829 5831 37887 5837
rect 37829 5828 37841 5831
rect 37700 5800 37841 5828
rect 37700 5788 37706 5800
rect 37829 5797 37841 5800
rect 37875 5797 37887 5831
rect 37829 5791 37887 5797
rect 38010 5788 38016 5840
rect 38068 5828 38074 5840
rect 39945 5831 40003 5837
rect 39945 5828 39957 5831
rect 38068 5800 39957 5828
rect 38068 5788 38074 5800
rect 39945 5797 39957 5800
rect 39991 5828 40003 5831
rect 40126 5828 40132 5840
rect 39991 5800 40132 5828
rect 39991 5797 40003 5800
rect 39945 5791 40003 5797
rect 40126 5788 40132 5800
rect 40184 5788 40190 5840
rect 14093 5763 14151 5769
rect 14093 5760 14105 5763
rect 10284 5732 10732 5760
rect 10284 5720 10290 5732
rect 7650 5692 7656 5704
rect 7611 5664 7656 5692
rect 7650 5652 7656 5664
rect 7708 5652 7714 5704
rect 8389 5695 8447 5701
rect 8389 5661 8401 5695
rect 8435 5692 8447 5695
rect 8662 5692 8668 5704
rect 8435 5664 8668 5692
rect 8435 5661 8447 5664
rect 8389 5655 8447 5661
rect 8662 5652 8668 5664
rect 8720 5652 8726 5704
rect 9122 5652 9128 5704
rect 9180 5692 9186 5704
rect 10704 5701 10732 5732
rect 11716 5732 14105 5760
rect 11716 5704 11744 5732
rect 14093 5729 14105 5732
rect 14139 5729 14151 5763
rect 14093 5723 14151 5729
rect 17862 5720 17868 5772
rect 17920 5760 17926 5772
rect 21634 5760 21640 5772
rect 17920 5732 21640 5760
rect 17920 5720 17926 5732
rect 9217 5695 9275 5701
rect 9217 5692 9229 5695
rect 9180 5664 9229 5692
rect 9180 5652 9186 5664
rect 9217 5661 9229 5664
rect 9263 5661 9275 5695
rect 9217 5655 9275 5661
rect 9861 5695 9919 5701
rect 9861 5661 9873 5695
rect 9907 5692 9919 5695
rect 10689 5695 10747 5701
rect 9907 5664 10640 5692
rect 9907 5661 9919 5664
rect 9861 5655 9919 5661
rect 9490 5624 9496 5636
rect 6886 5596 9496 5624
rect 9490 5584 9496 5596
rect 9548 5624 9554 5636
rect 9677 5627 9735 5633
rect 9677 5624 9689 5627
rect 9548 5596 9689 5624
rect 9548 5584 9554 5596
rect 9677 5593 9689 5596
rect 9723 5593 9735 5627
rect 9677 5587 9735 5593
rect 4062 5516 4068 5568
rect 4120 5516 4126 5568
rect 4433 5559 4491 5565
rect 4433 5525 4445 5559
rect 4479 5556 4491 5559
rect 4522 5556 4528 5568
rect 4479 5528 4528 5556
rect 4479 5525 4491 5528
rect 4433 5519 4491 5525
rect 4522 5516 4528 5528
rect 4580 5516 4586 5568
rect 7469 5559 7527 5565
rect 7469 5525 7481 5559
rect 7515 5556 7527 5559
rect 7834 5556 7840 5568
rect 7515 5528 7840 5556
rect 7515 5525 7527 5528
rect 7469 5519 7527 5525
rect 7834 5516 7840 5528
rect 7892 5516 7898 5568
rect 9033 5559 9091 5565
rect 9033 5525 9045 5559
rect 9079 5556 9091 5559
rect 10226 5556 10232 5568
rect 9079 5528 10232 5556
rect 9079 5525 9091 5528
rect 9033 5519 9091 5525
rect 10226 5516 10232 5528
rect 10284 5516 10290 5568
rect 10612 5556 10640 5664
rect 10689 5661 10701 5695
rect 10735 5692 10747 5695
rect 11698 5692 11704 5704
rect 10735 5664 11704 5692
rect 10735 5661 10747 5664
rect 10689 5655 10747 5661
rect 11698 5652 11704 5664
rect 11756 5652 11762 5704
rect 12529 5695 12587 5701
rect 12529 5692 12541 5695
rect 12084 5664 12541 5692
rect 10962 5633 10968 5636
rect 10956 5624 10968 5633
rect 10923 5596 10968 5624
rect 10956 5587 10968 5596
rect 10962 5584 10968 5587
rect 11020 5584 11026 5636
rect 12084 5565 12112 5664
rect 12529 5661 12541 5664
rect 12575 5661 12587 5695
rect 13446 5692 13452 5704
rect 13407 5664 13452 5692
rect 12529 5655 12587 5661
rect 13446 5652 13452 5664
rect 13504 5692 13510 5704
rect 13998 5692 14004 5704
rect 13504 5664 14004 5692
rect 13504 5652 13510 5664
rect 13998 5652 14004 5664
rect 14056 5652 14062 5704
rect 14182 5652 14188 5704
rect 14240 5692 14246 5704
rect 14349 5695 14407 5701
rect 14349 5692 14361 5695
rect 14240 5664 14361 5692
rect 14240 5652 14246 5664
rect 14349 5661 14361 5664
rect 14395 5661 14407 5695
rect 16390 5692 16396 5704
rect 16351 5664 16396 5692
rect 14349 5655 14407 5661
rect 16390 5652 16396 5664
rect 16448 5652 16454 5704
rect 16482 5652 16488 5704
rect 16540 5692 16546 5704
rect 16577 5695 16635 5701
rect 16577 5692 16589 5695
rect 16540 5664 16589 5692
rect 16540 5652 16546 5664
rect 16577 5661 16589 5664
rect 16623 5661 16635 5695
rect 16577 5655 16635 5661
rect 16666 5652 16672 5704
rect 16724 5692 16730 5704
rect 16807 5695 16865 5701
rect 16724 5664 16769 5692
rect 16724 5652 16730 5664
rect 16807 5661 16819 5695
rect 16853 5692 16865 5695
rect 17034 5692 17040 5704
rect 16853 5664 17040 5692
rect 16853 5661 16865 5664
rect 16807 5655 16865 5661
rect 17034 5652 17040 5664
rect 17092 5652 17098 5704
rect 18049 5695 18107 5701
rect 18049 5661 18061 5695
rect 18095 5661 18107 5695
rect 18230 5692 18236 5704
rect 18191 5664 18236 5692
rect 18049 5655 18107 5661
rect 13170 5584 13176 5636
rect 13228 5624 13234 5636
rect 13265 5627 13323 5633
rect 13265 5624 13277 5627
rect 13228 5596 13277 5624
rect 13228 5584 13234 5596
rect 13265 5593 13277 5596
rect 13311 5624 13323 5627
rect 18064 5624 18092 5655
rect 18230 5652 18236 5664
rect 18288 5652 18294 5704
rect 18340 5701 18368 5732
rect 21634 5720 21640 5732
rect 21692 5720 21698 5772
rect 23106 5760 23112 5772
rect 23067 5732 23112 5760
rect 23106 5720 23112 5732
rect 23164 5720 23170 5772
rect 23290 5720 23296 5772
rect 23348 5760 23354 5772
rect 24673 5763 24731 5769
rect 24673 5760 24685 5763
rect 23348 5732 24685 5760
rect 23348 5720 23354 5732
rect 24673 5729 24685 5732
rect 24719 5729 24731 5763
rect 24673 5723 24731 5729
rect 33042 5720 33048 5772
rect 33100 5760 33106 5772
rect 36357 5763 36415 5769
rect 36357 5760 36369 5763
rect 33100 5732 36369 5760
rect 33100 5720 33106 5732
rect 36357 5729 36369 5732
rect 36403 5729 36415 5763
rect 36357 5723 36415 5729
rect 36446 5720 36452 5772
rect 36504 5760 36510 5772
rect 36504 5732 38700 5760
rect 36504 5720 36510 5732
rect 18325 5695 18383 5701
rect 18325 5661 18337 5695
rect 18371 5661 18383 5695
rect 18325 5655 18383 5661
rect 18414 5652 18420 5704
rect 18472 5692 18478 5704
rect 18472 5664 18517 5692
rect 18472 5652 18478 5664
rect 18690 5652 18696 5704
rect 18748 5692 18754 5704
rect 19610 5692 19616 5704
rect 18748 5664 19616 5692
rect 18748 5652 18754 5664
rect 19610 5652 19616 5664
rect 19668 5652 19674 5704
rect 20625 5695 20683 5701
rect 20625 5661 20637 5695
rect 20671 5692 20683 5695
rect 21082 5692 21088 5704
rect 20671 5664 21088 5692
rect 20671 5661 20683 5664
rect 20625 5655 20683 5661
rect 21082 5652 21088 5664
rect 21140 5652 21146 5704
rect 21266 5692 21272 5704
rect 21227 5664 21272 5692
rect 21266 5652 21272 5664
rect 21324 5652 21330 5704
rect 22462 5652 22468 5704
rect 22520 5692 22526 5704
rect 22842 5695 22900 5701
rect 22842 5692 22854 5695
rect 22520 5664 22854 5692
rect 22520 5652 22526 5664
rect 22842 5661 22854 5664
rect 22888 5661 22900 5695
rect 23842 5692 23848 5704
rect 23803 5664 23848 5692
rect 22842 5655 22900 5661
rect 23842 5652 23848 5664
rect 23900 5652 23906 5704
rect 24946 5701 24952 5704
rect 24940 5692 24952 5701
rect 24907 5664 24952 5692
rect 24940 5655 24952 5664
rect 24946 5652 24952 5655
rect 25004 5652 25010 5704
rect 26789 5695 26847 5701
rect 26789 5661 26801 5695
rect 26835 5692 26847 5695
rect 26835 5664 27752 5692
rect 26835 5661 26847 5664
rect 26789 5655 26847 5661
rect 18708 5624 18736 5652
rect 13311 5596 18736 5624
rect 13311 5593 13323 5596
rect 13265 5587 13323 5593
rect 18874 5584 18880 5636
rect 18932 5624 18938 5636
rect 19245 5627 19303 5633
rect 19245 5624 19257 5627
rect 18932 5596 19257 5624
rect 18932 5584 18938 5596
rect 19245 5593 19257 5596
rect 19291 5593 19303 5627
rect 19426 5624 19432 5636
rect 19387 5596 19432 5624
rect 19245 5587 19303 5593
rect 19426 5584 19432 5596
rect 19484 5624 19490 5636
rect 19484 5596 21772 5624
rect 19484 5584 19490 5596
rect 12069 5559 12127 5565
rect 12069 5556 12081 5559
rect 10612 5528 12081 5556
rect 12069 5525 12081 5528
rect 12115 5525 12127 5559
rect 12710 5556 12716 5568
rect 12671 5528 12716 5556
rect 12069 5519 12127 5525
rect 12710 5516 12716 5528
rect 12768 5516 12774 5568
rect 13814 5516 13820 5568
rect 13872 5556 13878 5568
rect 14826 5556 14832 5568
rect 13872 5528 14832 5556
rect 13872 5516 13878 5528
rect 14826 5516 14832 5528
rect 14884 5556 14890 5568
rect 15473 5559 15531 5565
rect 15473 5556 15485 5559
rect 14884 5528 15485 5556
rect 14884 5516 14890 5528
rect 15473 5525 15485 5528
rect 15519 5525 15531 5559
rect 17034 5556 17040 5568
rect 16995 5528 17040 5556
rect 15473 5519 15531 5525
rect 17034 5516 17040 5528
rect 17092 5516 17098 5568
rect 18693 5559 18751 5565
rect 18693 5525 18705 5559
rect 18739 5556 18751 5559
rect 19518 5556 19524 5568
rect 18739 5528 19524 5556
rect 18739 5525 18751 5528
rect 18693 5519 18751 5525
rect 19518 5516 19524 5528
rect 19576 5516 19582 5568
rect 21744 5565 21772 5596
rect 24026 5584 24032 5636
rect 24084 5624 24090 5636
rect 26804 5624 26832 5655
rect 26970 5624 26976 5636
rect 24084 5596 26832 5624
rect 26931 5596 26976 5624
rect 24084 5584 24090 5596
rect 26970 5584 26976 5596
rect 27028 5624 27034 5636
rect 27724 5624 27752 5664
rect 28718 5652 28724 5704
rect 28776 5701 28782 5704
rect 28776 5692 28788 5701
rect 28994 5692 29000 5704
rect 28776 5664 28821 5692
rect 28955 5664 29000 5692
rect 28776 5655 28788 5664
rect 28776 5652 28782 5655
rect 28994 5652 29000 5664
rect 29052 5652 29058 5704
rect 29730 5692 29736 5704
rect 29691 5664 29736 5692
rect 29730 5652 29736 5664
rect 29788 5652 29794 5704
rect 30374 5692 30380 5704
rect 30335 5664 30380 5692
rect 30374 5652 30380 5664
rect 30432 5652 30438 5704
rect 32674 5692 32680 5704
rect 32635 5664 32680 5692
rect 32674 5652 32680 5664
rect 32732 5652 32738 5704
rect 34882 5692 34888 5704
rect 34843 5664 34888 5692
rect 34882 5652 34888 5664
rect 34940 5652 34946 5704
rect 34977 5695 35035 5701
rect 34977 5661 34989 5695
rect 35023 5661 35035 5695
rect 34977 5655 35035 5661
rect 29549 5627 29607 5633
rect 29549 5624 29561 5627
rect 27028 5596 27660 5624
rect 27724 5596 29561 5624
rect 27028 5584 27034 5596
rect 21729 5559 21787 5565
rect 21729 5525 21741 5559
rect 21775 5525 21787 5559
rect 21729 5519 21787 5525
rect 22186 5516 22192 5568
rect 22244 5556 22250 5568
rect 26234 5556 26240 5568
rect 22244 5528 26240 5556
rect 22244 5516 22250 5528
rect 26234 5516 26240 5528
rect 26292 5516 26298 5568
rect 27632 5565 27660 5596
rect 29549 5593 29561 5596
rect 29595 5593 29607 5627
rect 29549 5587 29607 5593
rect 29914 5584 29920 5636
rect 29972 5624 29978 5636
rect 32410 5627 32468 5633
rect 32410 5624 32422 5627
rect 29972 5596 32422 5624
rect 29972 5584 29978 5596
rect 32410 5593 32422 5596
rect 32456 5593 32468 5627
rect 32410 5587 32468 5593
rect 32582 5584 32588 5636
rect 32640 5624 32646 5636
rect 33318 5624 33324 5636
rect 32640 5596 33324 5624
rect 32640 5584 32646 5596
rect 33318 5584 33324 5596
rect 33376 5624 33382 5636
rect 34701 5627 34759 5633
rect 34701 5624 34713 5627
rect 33376 5596 34713 5624
rect 33376 5584 33382 5596
rect 34701 5593 34713 5596
rect 34747 5624 34759 5627
rect 34992 5624 35020 5655
rect 35342 5652 35348 5704
rect 35400 5692 35406 5704
rect 35437 5695 35495 5701
rect 35437 5692 35449 5695
rect 35400 5664 35449 5692
rect 35400 5652 35406 5664
rect 35437 5661 35449 5664
rect 35483 5661 35495 5695
rect 36078 5692 36084 5704
rect 36039 5664 36084 5692
rect 35437 5655 35495 5661
rect 36078 5652 36084 5664
rect 36136 5652 36142 5704
rect 38562 5692 38568 5704
rect 38523 5664 38568 5692
rect 38562 5652 38568 5664
rect 38620 5652 38626 5704
rect 35894 5624 35900 5636
rect 34747 5596 34928 5624
rect 34992 5596 35900 5624
rect 34747 5593 34759 5596
rect 34701 5587 34759 5593
rect 27617 5559 27675 5565
rect 27617 5525 27629 5559
rect 27663 5525 27675 5559
rect 27617 5519 27675 5525
rect 30742 5516 30748 5568
rect 30800 5556 30806 5568
rect 34790 5556 34796 5568
rect 30800 5528 34796 5556
rect 30800 5516 30806 5528
rect 34790 5516 34796 5528
rect 34848 5516 34854 5568
rect 34900 5556 34928 5596
rect 35894 5584 35900 5596
rect 35952 5584 35958 5636
rect 38473 5627 38531 5633
rect 38473 5624 38485 5627
rect 37582 5596 38485 5624
rect 38473 5593 38485 5596
rect 38519 5593 38531 5627
rect 38672 5624 38700 5732
rect 40034 5720 40040 5772
rect 40092 5760 40098 5772
rect 41049 5763 41107 5769
rect 41049 5760 41061 5763
rect 40092 5732 41061 5760
rect 40092 5720 40098 5732
rect 41049 5729 41061 5732
rect 41095 5729 41107 5763
rect 41156 5760 41184 5868
rect 41312 5865 41324 5899
rect 41312 5859 41328 5865
rect 41322 5856 41328 5859
rect 41380 5856 41386 5908
rect 42426 5856 42432 5908
rect 42484 5896 42490 5908
rect 42797 5899 42855 5905
rect 42797 5896 42809 5899
rect 42484 5868 42809 5896
rect 42484 5856 42490 5868
rect 42797 5865 42809 5868
rect 42843 5865 42855 5899
rect 43990 5896 43996 5908
rect 43951 5868 43996 5896
rect 42797 5859 42855 5865
rect 43990 5856 43996 5868
rect 44048 5856 44054 5908
rect 45646 5896 45652 5908
rect 45204 5868 45652 5896
rect 43349 5831 43407 5837
rect 43349 5797 43361 5831
rect 43395 5828 43407 5831
rect 45204 5828 45232 5868
rect 45646 5856 45652 5868
rect 45704 5856 45710 5908
rect 51537 5899 51595 5905
rect 51537 5896 51549 5899
rect 50356 5868 51549 5896
rect 43395 5800 45232 5828
rect 43395 5797 43407 5800
rect 43349 5791 43407 5797
rect 43364 5760 43392 5791
rect 45554 5788 45560 5840
rect 45612 5828 45618 5840
rect 46293 5831 46351 5837
rect 46293 5828 46305 5831
rect 45612 5800 46305 5828
rect 45612 5788 45618 5800
rect 46293 5797 46305 5800
rect 46339 5797 46351 5831
rect 46293 5791 46351 5797
rect 49234 5788 49240 5840
rect 49292 5828 49298 5840
rect 50249 5831 50307 5837
rect 50249 5828 50261 5831
rect 49292 5800 50261 5828
rect 49292 5788 49298 5800
rect 50249 5797 50261 5800
rect 50295 5797 50307 5831
rect 50249 5791 50307 5797
rect 41156 5732 43392 5760
rect 41049 5723 41107 5729
rect 45370 5720 45376 5772
rect 45428 5760 45434 5772
rect 47578 5760 47584 5772
rect 45428 5732 47584 5760
rect 45428 5720 45434 5732
rect 47578 5720 47584 5732
rect 47636 5760 47642 5772
rect 47857 5763 47915 5769
rect 47857 5760 47869 5763
rect 47636 5732 47869 5760
rect 47636 5720 47642 5732
rect 47857 5729 47869 5732
rect 47903 5729 47915 5763
rect 47857 5723 47915 5729
rect 48133 5763 48191 5769
rect 48133 5729 48145 5763
rect 48179 5760 48191 5763
rect 50356 5760 50384 5868
rect 51537 5865 51549 5868
rect 51583 5865 51595 5899
rect 53561 5899 53619 5905
rect 53561 5896 53573 5899
rect 51537 5859 51595 5865
rect 52012 5868 53573 5896
rect 50798 5828 50804 5840
rect 50759 5800 50804 5828
rect 50798 5788 50804 5800
rect 50856 5828 50862 5840
rect 52012 5828 52040 5868
rect 53561 5865 53573 5868
rect 53607 5865 53619 5899
rect 53561 5859 53619 5865
rect 50856 5800 52040 5828
rect 50856 5788 50862 5800
rect 53190 5788 53196 5840
rect 53248 5828 53254 5840
rect 56597 5831 56655 5837
rect 56597 5828 56609 5831
rect 53248 5800 56609 5828
rect 53248 5788 53254 5800
rect 56597 5797 56609 5800
rect 56643 5797 56655 5831
rect 56597 5791 56655 5797
rect 48179 5732 50384 5760
rect 48179 5729 48191 5732
rect 48133 5723 48191 5729
rect 52546 5720 52552 5772
rect 52604 5760 52610 5772
rect 57609 5763 57667 5769
rect 52604 5732 52649 5760
rect 52604 5720 52610 5732
rect 57609 5729 57621 5763
rect 57655 5760 57667 5763
rect 57790 5760 57796 5772
rect 57655 5732 57796 5760
rect 57655 5729 57667 5732
rect 57609 5723 57667 5729
rect 57790 5720 57796 5732
rect 57848 5720 57854 5772
rect 40402 5692 40408 5704
rect 40363 5664 40408 5692
rect 40402 5652 40408 5664
rect 40460 5652 40466 5704
rect 42426 5652 42432 5704
rect 42484 5652 42490 5704
rect 44174 5692 44180 5704
rect 44135 5664 44180 5692
rect 44174 5652 44180 5664
rect 44232 5652 44238 5704
rect 45002 5692 45008 5704
rect 44963 5664 45008 5692
rect 45002 5652 45008 5664
rect 45060 5652 45066 5704
rect 45278 5652 45284 5704
rect 45336 5692 45342 5704
rect 45649 5695 45707 5701
rect 45649 5692 45661 5695
rect 45336 5664 45661 5692
rect 45336 5652 45342 5664
rect 45649 5661 45661 5664
rect 45695 5661 45707 5695
rect 47210 5692 47216 5704
rect 47171 5664 47216 5692
rect 45649 5655 45707 5661
rect 47210 5652 47216 5664
rect 47268 5652 47274 5704
rect 49234 5652 49240 5704
rect 49292 5652 49298 5704
rect 50157 5695 50215 5701
rect 50157 5661 50169 5695
rect 50203 5661 50215 5695
rect 50157 5655 50215 5661
rect 41414 5624 41420 5636
rect 38672 5596 41420 5624
rect 38473 5587 38531 5593
rect 41414 5584 41420 5596
rect 41472 5584 41478 5636
rect 46842 5584 46848 5636
rect 46900 5624 46906 5636
rect 50172 5624 50200 5655
rect 52178 5652 52184 5704
rect 52236 5692 52242 5704
rect 52273 5695 52331 5701
rect 52273 5692 52285 5695
rect 52236 5664 52285 5692
rect 52236 5652 52242 5664
rect 52273 5661 52285 5664
rect 52319 5661 52331 5695
rect 52273 5655 52331 5661
rect 54113 5695 54171 5701
rect 54113 5661 54125 5695
rect 54159 5661 54171 5695
rect 54113 5655 54171 5661
rect 54128 5624 54156 5655
rect 55214 5652 55220 5704
rect 55272 5692 55278 5704
rect 55309 5695 55367 5701
rect 55309 5692 55321 5695
rect 55272 5664 55321 5692
rect 55272 5652 55278 5664
rect 55309 5661 55321 5664
rect 55355 5661 55367 5695
rect 55582 5692 55588 5704
rect 55543 5664 55588 5692
rect 55309 5655 55367 5661
rect 55582 5652 55588 5664
rect 55640 5652 55646 5704
rect 57330 5692 57336 5704
rect 57291 5664 57336 5692
rect 57330 5652 57336 5664
rect 57388 5652 57394 5704
rect 55950 5624 55956 5636
rect 46900 5596 48544 5624
rect 46900 5584 46906 5596
rect 37734 5556 37740 5568
rect 34900 5528 37740 5556
rect 37734 5516 37740 5528
rect 37792 5516 37798 5568
rect 39114 5556 39120 5568
rect 39075 5528 39120 5556
rect 39114 5516 39120 5528
rect 39172 5516 39178 5568
rect 40589 5559 40647 5565
rect 40589 5525 40601 5559
rect 40635 5556 40647 5559
rect 43346 5556 43352 5568
rect 40635 5528 43352 5556
rect 40635 5525 40647 5528
rect 40589 5519 40647 5525
rect 43346 5516 43352 5528
rect 43404 5516 43410 5568
rect 45189 5559 45247 5565
rect 45189 5525 45201 5559
rect 45235 5556 45247 5559
rect 46566 5556 46572 5568
rect 45235 5528 46572 5556
rect 45235 5525 45247 5528
rect 45189 5519 45247 5525
rect 46566 5516 46572 5528
rect 46624 5516 46630 5568
rect 47305 5559 47363 5565
rect 47305 5525 47317 5559
rect 47351 5556 47363 5559
rect 48314 5556 48320 5568
rect 47351 5528 48320 5556
rect 47351 5525 47363 5528
rect 47305 5519 47363 5525
rect 48314 5516 48320 5528
rect 48372 5516 48378 5568
rect 48516 5556 48544 5596
rect 49528 5596 50200 5624
rect 50356 5596 55956 5624
rect 49528 5556 49556 5596
rect 48516 5528 49556 5556
rect 49605 5559 49663 5565
rect 49605 5525 49617 5559
rect 49651 5556 49663 5559
rect 50356 5556 50384 5596
rect 55950 5584 55956 5596
rect 56008 5584 56014 5636
rect 49651 5528 50384 5556
rect 53101 5559 53159 5565
rect 49651 5525 49663 5528
rect 49605 5519 49663 5525
rect 53101 5525 53113 5559
rect 53147 5556 53159 5559
rect 53834 5556 53840 5568
rect 53147 5528 53840 5556
rect 53147 5525 53159 5528
rect 53101 5519 53159 5525
rect 53834 5516 53840 5528
rect 53892 5516 53898 5568
rect 54202 5556 54208 5568
rect 54115 5528 54208 5556
rect 54202 5516 54208 5528
rect 54260 5556 54266 5568
rect 55674 5556 55680 5568
rect 54260 5528 55680 5556
rect 54260 5516 54266 5528
rect 55674 5516 55680 5528
rect 55732 5516 55738 5568
rect 57974 5516 57980 5568
rect 58032 5556 58038 5568
rect 58069 5559 58127 5565
rect 58069 5556 58081 5559
rect 58032 5528 58081 5556
rect 58032 5516 58038 5528
rect 58069 5525 58081 5528
rect 58115 5525 58127 5559
rect 58069 5519 58127 5525
rect 1104 5466 58880 5488
rect 1104 5414 15398 5466
rect 15450 5414 15462 5466
rect 15514 5414 15526 5466
rect 15578 5414 15590 5466
rect 15642 5414 15654 5466
rect 15706 5414 29846 5466
rect 29898 5414 29910 5466
rect 29962 5414 29974 5466
rect 30026 5414 30038 5466
rect 30090 5414 30102 5466
rect 30154 5414 44294 5466
rect 44346 5414 44358 5466
rect 44410 5414 44422 5466
rect 44474 5414 44486 5466
rect 44538 5414 44550 5466
rect 44602 5414 58880 5466
rect 1104 5392 58880 5414
rect 2317 5355 2375 5361
rect 2317 5321 2329 5355
rect 2363 5352 2375 5355
rect 3970 5352 3976 5364
rect 2363 5324 3976 5352
rect 2363 5321 2375 5324
rect 2317 5315 2375 5321
rect 3970 5312 3976 5324
rect 4028 5312 4034 5364
rect 9033 5355 9091 5361
rect 9033 5352 9045 5355
rect 4356 5324 9045 5352
rect 1946 5284 1952 5296
rect 1859 5256 1952 5284
rect 1946 5244 1952 5256
rect 2004 5284 2010 5296
rect 2774 5284 2780 5296
rect 2004 5256 2780 5284
rect 2004 5244 2010 5256
rect 2774 5244 2780 5256
rect 2832 5244 2838 5296
rect 3142 5284 3148 5296
rect 3103 5256 3148 5284
rect 3142 5244 3148 5256
rect 3200 5244 3206 5296
rect 4356 5284 4384 5324
rect 9033 5321 9045 5324
rect 9079 5352 9091 5355
rect 10042 5352 10048 5364
rect 9079 5324 10048 5352
rect 9079 5321 9091 5324
rect 9033 5315 9091 5321
rect 10042 5312 10048 5324
rect 10100 5312 10106 5364
rect 10633 5324 11836 5352
rect 5442 5284 5448 5296
rect 3712 5256 4384 5284
rect 4448 5256 5448 5284
rect 2130 5216 2136 5228
rect 2091 5188 2136 5216
rect 2130 5176 2136 5188
rect 2188 5176 2194 5228
rect 2961 5219 3019 5225
rect 2961 5185 2973 5219
rect 3007 5216 3019 5219
rect 3712 5216 3740 5256
rect 3007 5188 3740 5216
rect 3789 5219 3847 5225
rect 3007 5185 3019 5188
rect 2961 5179 3019 5185
rect 3789 5185 3801 5219
rect 3835 5216 3847 5219
rect 4246 5216 4252 5228
rect 3835 5188 4252 5216
rect 3835 5185 3847 5188
rect 3789 5179 3847 5185
rect 4246 5176 4252 5188
rect 4304 5176 4310 5228
rect 4448 5225 4476 5256
rect 5442 5244 5448 5256
rect 5500 5244 5506 5296
rect 7374 5244 7380 5296
rect 7432 5284 7438 5296
rect 7898 5287 7956 5293
rect 7898 5284 7910 5287
rect 7432 5256 7910 5284
rect 7432 5244 7438 5256
rect 7898 5253 7910 5256
rect 7944 5253 7956 5287
rect 7898 5247 7956 5253
rect 9493 5287 9551 5293
rect 9493 5253 9505 5287
rect 9539 5284 9551 5287
rect 9861 5287 9919 5293
rect 9539 5256 9812 5284
rect 9539 5253 9551 5256
rect 9493 5247 9551 5253
rect 4433 5219 4491 5225
rect 4433 5185 4445 5219
rect 4479 5185 4491 5219
rect 4433 5179 4491 5185
rect 1489 5151 1547 5157
rect 1489 5117 1501 5151
rect 1535 5148 1547 5151
rect 4448 5148 4476 5179
rect 4522 5176 4528 5228
rect 4580 5216 4586 5228
rect 4689 5219 4747 5225
rect 4689 5216 4701 5219
rect 4580 5188 4701 5216
rect 4580 5176 4586 5188
rect 4689 5185 4701 5188
rect 4735 5185 4747 5219
rect 4689 5179 4747 5185
rect 7193 5219 7251 5225
rect 7193 5185 7205 5219
rect 7239 5216 7251 5219
rect 7282 5216 7288 5228
rect 7239 5188 7288 5216
rect 7239 5185 7251 5188
rect 7193 5179 7251 5185
rect 7282 5176 7288 5188
rect 7340 5176 7346 5228
rect 7653 5219 7711 5225
rect 7653 5185 7665 5219
rect 7699 5216 7711 5219
rect 8202 5216 8208 5228
rect 7699 5188 8208 5216
rect 7699 5185 7711 5188
rect 7653 5179 7711 5185
rect 1535 5120 4476 5148
rect 1535 5117 1547 5120
rect 1489 5111 1547 5117
rect 5442 5108 5448 5160
rect 5500 5148 5506 5160
rect 6457 5151 6515 5157
rect 6457 5148 6469 5151
rect 5500 5120 6469 5148
rect 5500 5108 5506 5120
rect 6457 5117 6469 5120
rect 6503 5148 6515 5151
rect 6822 5148 6828 5160
rect 6503 5120 6828 5148
rect 6503 5117 6515 5120
rect 6457 5111 6515 5117
rect 6822 5108 6828 5120
rect 6880 5148 6886 5160
rect 7668 5148 7696 5179
rect 8202 5176 8208 5188
rect 8260 5176 8266 5228
rect 9677 5219 9735 5225
rect 9677 5216 9689 5219
rect 8772 5188 9689 5216
rect 6880 5120 7696 5148
rect 6880 5108 6886 5120
rect 3973 5083 4031 5089
rect 3973 5049 3985 5083
rect 4019 5049 4031 5083
rect 5810 5080 5816 5092
rect 5771 5052 5816 5080
rect 3973 5043 4031 5049
rect 3988 5012 4016 5043
rect 5810 5040 5816 5052
rect 5868 5040 5874 5092
rect 4798 5012 4804 5024
rect 3988 4984 4804 5012
rect 4798 4972 4804 4984
rect 4856 5012 4862 5024
rect 5994 5012 6000 5024
rect 4856 4984 6000 5012
rect 4856 4972 4862 4984
rect 5994 4972 6000 4984
rect 6052 4972 6058 5024
rect 7009 5015 7067 5021
rect 7009 4981 7021 5015
rect 7055 5012 7067 5015
rect 7374 5012 7380 5024
rect 7055 4984 7380 5012
rect 7055 4981 7067 4984
rect 7009 4975 7067 4981
rect 7374 4972 7380 4984
rect 7432 4972 7438 5024
rect 7926 4972 7932 5024
rect 7984 5012 7990 5024
rect 8772 5012 8800 5188
rect 9677 5185 9689 5188
rect 9723 5185 9735 5219
rect 9677 5179 9735 5185
rect 9784 5148 9812 5256
rect 9861 5253 9873 5287
rect 9907 5284 9919 5287
rect 10502 5284 10508 5296
rect 9907 5256 10508 5284
rect 9907 5253 9919 5256
rect 9861 5247 9919 5253
rect 10502 5244 10508 5256
rect 10560 5284 10566 5296
rect 10633 5284 10661 5324
rect 10560 5256 10661 5284
rect 10704 5256 11192 5284
rect 10560 5244 10566 5256
rect 10244 5216 10364 5219
rect 10594 5216 10600 5228
rect 9966 5191 10456 5216
rect 9966 5188 10272 5191
rect 10336 5188 10456 5191
rect 10555 5188 10600 5216
rect 9966 5148 9994 5188
rect 9784 5120 9994 5148
rect 9490 5040 9496 5092
rect 9548 5080 9554 5092
rect 9858 5080 9864 5092
rect 9548 5052 9864 5080
rect 9548 5040 9554 5052
rect 9858 5040 9864 5052
rect 9916 5040 9922 5092
rect 10428 5080 10456 5188
rect 10594 5176 10600 5188
rect 10652 5176 10658 5228
rect 10704 5225 10732 5256
rect 10689 5219 10747 5225
rect 10689 5185 10701 5219
rect 10735 5185 10747 5219
rect 10689 5179 10747 5185
rect 10781 5219 10839 5225
rect 10781 5185 10793 5219
rect 10827 5185 10839 5219
rect 10781 5179 10839 5185
rect 10977 5219 11035 5225
rect 10977 5185 10989 5219
rect 11023 5185 11035 5219
rect 10977 5179 11035 5185
rect 10796 5080 10824 5179
rect 10980 5092 11008 5179
rect 10428 5052 10824 5080
rect 10962 5040 10968 5092
rect 11020 5040 11026 5092
rect 11164 5080 11192 5256
rect 11808 5225 11836 5324
rect 13722 5312 13728 5364
rect 13780 5352 13786 5364
rect 16117 5355 16175 5361
rect 13780 5324 15976 5352
rect 13780 5312 13786 5324
rect 12894 5244 12900 5296
rect 12952 5284 12958 5296
rect 12952 5256 14412 5284
rect 12952 5244 12958 5256
rect 11793 5219 11851 5225
rect 11793 5185 11805 5219
rect 11839 5216 11851 5219
rect 11882 5216 11888 5228
rect 11839 5188 11888 5216
rect 11839 5185 11851 5188
rect 11793 5179 11851 5185
rect 11882 5176 11888 5188
rect 11940 5176 11946 5228
rect 13998 5176 14004 5228
rect 14056 5216 14062 5228
rect 14384 5225 14412 5256
rect 14918 5244 14924 5296
rect 14976 5284 14982 5296
rect 15948 5293 15976 5324
rect 16117 5321 16129 5355
rect 16163 5352 16175 5355
rect 16482 5352 16488 5364
rect 16163 5324 16488 5352
rect 16163 5321 16175 5324
rect 16117 5315 16175 5321
rect 16482 5312 16488 5324
rect 16540 5312 16546 5364
rect 16669 5355 16727 5361
rect 16669 5321 16681 5355
rect 16715 5321 16727 5355
rect 16669 5315 16727 5321
rect 15933 5287 15991 5293
rect 14976 5256 15884 5284
rect 14976 5244 14982 5256
rect 14093 5219 14151 5225
rect 14093 5216 14105 5219
rect 14056 5188 14105 5216
rect 14056 5176 14062 5188
rect 14093 5185 14105 5188
rect 14139 5185 14151 5219
rect 14093 5179 14151 5185
rect 14369 5219 14427 5225
rect 14369 5185 14381 5219
rect 14415 5185 14427 5219
rect 14369 5179 14427 5185
rect 15102 5176 15108 5228
rect 15160 5216 15166 5228
rect 15749 5219 15807 5225
rect 15749 5216 15761 5219
rect 15160 5188 15761 5216
rect 15160 5176 15166 5188
rect 15749 5185 15761 5188
rect 15795 5185 15807 5219
rect 15856 5216 15884 5256
rect 15933 5253 15945 5287
rect 15979 5284 15991 5287
rect 16684 5284 16712 5315
rect 16942 5312 16948 5364
rect 17000 5352 17006 5364
rect 17402 5352 17408 5364
rect 17000 5324 17408 5352
rect 17000 5312 17006 5324
rect 17402 5312 17408 5324
rect 17460 5312 17466 5364
rect 18230 5312 18236 5364
rect 18288 5352 18294 5364
rect 18509 5355 18567 5361
rect 18509 5352 18521 5355
rect 18288 5324 18521 5352
rect 18288 5312 18294 5324
rect 18509 5321 18521 5324
rect 18555 5321 18567 5355
rect 19889 5355 19947 5361
rect 19889 5352 19901 5355
rect 18509 5315 18567 5321
rect 19306 5324 19901 5352
rect 15979 5256 16712 5284
rect 15979 5253 15991 5256
rect 15933 5247 15991 5253
rect 17034 5244 17040 5296
rect 17092 5284 17098 5296
rect 17782 5287 17840 5293
rect 17782 5284 17794 5287
rect 17092 5256 17794 5284
rect 17092 5244 17098 5256
rect 17782 5253 17794 5256
rect 17828 5253 17840 5287
rect 17782 5247 17840 5253
rect 17954 5244 17960 5296
rect 18012 5284 18018 5296
rect 18874 5284 18880 5296
rect 18012 5256 18880 5284
rect 18012 5244 18018 5256
rect 18874 5244 18880 5256
rect 18932 5244 18938 5296
rect 18693 5219 18751 5225
rect 18693 5216 18705 5219
rect 15856 5188 18705 5216
rect 15749 5179 15807 5185
rect 18693 5185 18705 5188
rect 18739 5216 18751 5219
rect 19306 5216 19334 5324
rect 19889 5321 19901 5324
rect 19935 5321 19947 5355
rect 19889 5315 19947 5321
rect 21174 5312 21180 5364
rect 21232 5352 21238 5364
rect 22370 5352 22376 5364
rect 21232 5324 22376 5352
rect 21232 5312 21238 5324
rect 22370 5312 22376 5324
rect 22428 5312 22434 5364
rect 24673 5355 24731 5361
rect 24673 5321 24685 5355
rect 24719 5321 24731 5355
rect 24673 5315 24731 5321
rect 19518 5244 19524 5296
rect 19576 5284 19582 5296
rect 21002 5287 21060 5293
rect 21002 5284 21014 5287
rect 19576 5256 21014 5284
rect 19576 5244 19582 5256
rect 21002 5253 21014 5256
rect 21048 5253 21060 5287
rect 21002 5247 21060 5253
rect 21450 5244 21456 5296
rect 21508 5284 21514 5296
rect 24578 5284 24584 5296
rect 21508 5256 24584 5284
rect 21508 5244 21514 5256
rect 24578 5244 24584 5256
rect 24636 5244 24642 5296
rect 24688 5284 24716 5315
rect 25958 5312 25964 5364
rect 26016 5352 26022 5364
rect 27982 5352 27988 5364
rect 26016 5324 27988 5352
rect 26016 5312 26022 5324
rect 27982 5312 27988 5324
rect 28040 5312 28046 5364
rect 31294 5312 31300 5364
rect 31352 5352 31358 5364
rect 32493 5355 32551 5361
rect 32493 5352 32505 5355
rect 31352 5324 32505 5352
rect 31352 5312 31358 5324
rect 32493 5321 32505 5324
rect 32539 5321 32551 5355
rect 34790 5352 34796 5364
rect 32493 5315 32551 5321
rect 33244 5324 34796 5352
rect 24688 5256 26372 5284
rect 18739 5188 19334 5216
rect 18739 5185 18751 5188
rect 18693 5179 18751 5185
rect 21726 5176 21732 5228
rect 21784 5216 21790 5228
rect 21821 5219 21879 5225
rect 21821 5216 21833 5219
rect 21784 5188 21833 5216
rect 21784 5176 21790 5188
rect 21821 5185 21833 5188
rect 21867 5185 21879 5219
rect 21821 5179 21879 5185
rect 22278 5176 22284 5228
rect 22336 5216 22342 5228
rect 23290 5216 23296 5228
rect 22336 5188 23296 5216
rect 22336 5176 22342 5188
rect 23290 5176 23296 5188
rect 23348 5176 23354 5228
rect 23382 5176 23388 5228
rect 23440 5216 23446 5228
rect 25700 5225 25728 5256
rect 23549 5219 23607 5225
rect 23549 5216 23561 5219
rect 23440 5188 23561 5216
rect 23440 5176 23446 5188
rect 23549 5185 23561 5188
rect 23595 5185 23607 5219
rect 23549 5179 23607 5185
rect 25685 5219 25743 5225
rect 25685 5185 25697 5219
rect 25731 5185 25743 5219
rect 25685 5179 25743 5185
rect 25869 5219 25927 5225
rect 25869 5185 25881 5219
rect 25915 5185 25927 5219
rect 25869 5179 25927 5185
rect 11514 5148 11520 5160
rect 11475 5120 11520 5148
rect 11514 5108 11520 5120
rect 11572 5148 11578 5160
rect 12805 5151 12863 5157
rect 12805 5148 12817 5151
rect 11572 5120 12817 5148
rect 11572 5108 11578 5120
rect 12805 5117 12817 5120
rect 12851 5117 12863 5151
rect 12805 5111 12863 5117
rect 13081 5151 13139 5157
rect 13081 5117 13093 5151
rect 13127 5148 13139 5151
rect 15120 5148 15148 5176
rect 13127 5120 15148 5148
rect 13127 5117 13139 5120
rect 13081 5111 13139 5117
rect 15838 5108 15844 5160
rect 15896 5148 15902 5160
rect 16482 5148 16488 5160
rect 15896 5120 16488 5148
rect 15896 5108 15902 5120
rect 16482 5108 16488 5120
rect 16540 5108 16546 5160
rect 18049 5151 18107 5157
rect 18049 5117 18061 5151
rect 18095 5148 18107 5151
rect 19518 5148 19524 5160
rect 18095 5120 19524 5148
rect 18095 5117 18107 5120
rect 18049 5111 18107 5117
rect 16942 5080 16948 5092
rect 11164 5052 16948 5080
rect 16942 5040 16948 5052
rect 17000 5040 17006 5092
rect 7984 4984 8800 5012
rect 10321 5015 10379 5021
rect 7984 4972 7990 4984
rect 10321 4981 10333 5015
rect 10367 5012 10379 5015
rect 10410 5012 10416 5024
rect 10367 4984 10416 5012
rect 10367 4981 10379 4984
rect 10321 4975 10379 4981
rect 10410 4972 10416 4984
rect 10468 4972 10474 5024
rect 11974 4972 11980 5024
rect 12032 5012 12038 5024
rect 15194 5012 15200 5024
rect 12032 4984 15200 5012
rect 12032 4972 12038 4984
rect 15194 4972 15200 4984
rect 15252 4972 15258 5024
rect 16758 4972 16764 5024
rect 16816 5012 16822 5024
rect 18064 5012 18092 5111
rect 19518 5108 19524 5120
rect 19576 5108 19582 5160
rect 21269 5151 21327 5157
rect 21269 5117 21281 5151
rect 21315 5148 21327 5151
rect 21634 5148 21640 5160
rect 21315 5120 21640 5148
rect 21315 5117 21327 5120
rect 21269 5111 21327 5117
rect 21634 5108 21640 5120
rect 21692 5148 21698 5160
rect 23106 5148 23112 5160
rect 21692 5120 23112 5148
rect 21692 5108 21698 5120
rect 23106 5108 23112 5120
rect 23164 5108 23170 5160
rect 25498 5108 25504 5160
rect 25556 5148 25562 5160
rect 25884 5148 25912 5179
rect 25958 5176 25964 5228
rect 26016 5216 26022 5228
rect 26016 5188 26061 5216
rect 26016 5176 26022 5188
rect 26344 5148 26372 5256
rect 27522 5244 27528 5296
rect 27580 5284 27586 5296
rect 32674 5284 32680 5296
rect 27580 5256 32680 5284
rect 27580 5244 27586 5256
rect 26418 5176 26424 5228
rect 26476 5216 26482 5228
rect 26973 5219 27031 5225
rect 26973 5216 26985 5219
rect 26476 5188 26985 5216
rect 26476 5176 26482 5188
rect 26973 5185 26985 5188
rect 27019 5185 27031 5219
rect 27706 5216 27712 5228
rect 27667 5188 27712 5216
rect 26973 5179 27031 5185
rect 27706 5176 27712 5188
rect 27764 5176 27770 5228
rect 27798 5176 27804 5228
rect 27856 5216 27862 5228
rect 27893 5219 27951 5225
rect 27893 5216 27905 5219
rect 27856 5188 27905 5216
rect 27856 5176 27862 5188
rect 27893 5185 27905 5188
rect 27939 5185 27951 5219
rect 27893 5179 27951 5185
rect 27982 5176 27988 5228
rect 28040 5216 28046 5228
rect 28442 5216 28448 5228
rect 28040 5188 28085 5216
rect 28403 5188 28448 5216
rect 28040 5176 28046 5188
rect 28442 5176 28448 5188
rect 28500 5176 28506 5228
rect 28718 5216 28724 5228
rect 28679 5188 28724 5216
rect 28718 5176 28724 5188
rect 28776 5176 28782 5228
rect 30208 5225 30236 5256
rect 32674 5244 32680 5256
rect 32732 5244 32738 5296
rect 33244 5293 33272 5324
rect 34790 5312 34796 5324
rect 34848 5312 34854 5364
rect 37553 5355 37611 5361
rect 37553 5321 37565 5355
rect 37599 5352 37611 5355
rect 38654 5352 38660 5364
rect 37599 5324 38660 5352
rect 37599 5321 37611 5324
rect 37553 5315 37611 5321
rect 38654 5312 38660 5324
rect 38712 5312 38718 5364
rect 38764 5324 41414 5352
rect 33229 5287 33287 5293
rect 33229 5253 33241 5287
rect 33275 5253 33287 5287
rect 33229 5247 33287 5253
rect 34514 5244 34520 5296
rect 34572 5244 34578 5296
rect 38562 5244 38568 5296
rect 38620 5284 38626 5296
rect 38764 5284 38792 5324
rect 40034 5284 40040 5296
rect 38620 5256 38792 5284
rect 38856 5256 40040 5284
rect 38620 5244 38626 5256
rect 30193 5219 30251 5225
rect 30193 5185 30205 5219
rect 30239 5185 30251 5219
rect 30193 5179 30251 5185
rect 30282 5176 30288 5228
rect 30340 5216 30346 5228
rect 30449 5219 30507 5225
rect 30449 5216 30461 5219
rect 30340 5188 30461 5216
rect 30340 5176 30346 5188
rect 30449 5185 30461 5188
rect 30495 5185 30507 5219
rect 32309 5219 32367 5225
rect 32309 5216 32321 5219
rect 30449 5179 30507 5185
rect 31588 5188 32321 5216
rect 28537 5151 28595 5157
rect 28537 5148 28549 5151
rect 25556 5120 26096 5148
rect 26344 5120 28549 5148
rect 25556 5108 25562 5120
rect 26068 5080 26096 5120
rect 28537 5117 28549 5120
rect 28583 5117 28595 5151
rect 28537 5111 28595 5117
rect 24780 5052 25728 5080
rect 26068 5052 27660 5080
rect 19334 5012 19340 5024
rect 16816 4984 18092 5012
rect 19295 4984 19340 5012
rect 16816 4972 16822 4984
rect 19334 4972 19340 4984
rect 19392 4972 19398 5024
rect 20898 4972 20904 5024
rect 20956 5012 20962 5024
rect 22005 5015 22063 5021
rect 22005 5012 22017 5015
rect 20956 4984 22017 5012
rect 20956 4972 20962 4984
rect 22005 4981 22017 4984
rect 22051 4981 22063 5015
rect 22005 4975 22063 4981
rect 22833 5015 22891 5021
rect 22833 4981 22845 5015
rect 22879 5012 22891 5015
rect 24780 5012 24808 5052
rect 22879 4984 24808 5012
rect 22879 4981 22891 4984
rect 22833 4975 22891 4981
rect 24946 4972 24952 5024
rect 25004 5012 25010 5024
rect 25501 5015 25559 5021
rect 25501 5012 25513 5015
rect 25004 4984 25513 5012
rect 25004 4972 25010 4984
rect 25501 4981 25513 4984
rect 25547 4981 25559 5015
rect 25700 5012 25728 5052
rect 26786 5012 26792 5024
rect 25700 4984 26792 5012
rect 25501 4975 25559 4981
rect 26786 4972 26792 4984
rect 26844 4972 26850 5024
rect 26878 4972 26884 5024
rect 26936 5012 26942 5024
rect 27525 5015 27583 5021
rect 27525 5012 27537 5015
rect 26936 4984 27537 5012
rect 26936 4972 26942 4984
rect 27525 4981 27537 4984
rect 27571 4981 27583 5015
rect 27632 5012 27660 5052
rect 27706 5040 27712 5092
rect 27764 5080 27770 5092
rect 28718 5080 28724 5092
rect 27764 5052 28724 5080
rect 27764 5040 27770 5052
rect 28718 5040 28724 5052
rect 28776 5040 28782 5092
rect 28902 5080 28908 5092
rect 28863 5052 28908 5080
rect 28902 5040 28908 5052
rect 28960 5040 28966 5092
rect 29288 5052 30236 5080
rect 27798 5012 27804 5024
rect 27632 4984 27804 5012
rect 27525 4975 27583 4981
rect 27798 4972 27804 4984
rect 27856 4972 27862 5024
rect 28629 5015 28687 5021
rect 28629 4981 28641 5015
rect 28675 5012 28687 5015
rect 29288 5012 29316 5052
rect 29454 5012 29460 5024
rect 28675 4984 29316 5012
rect 29415 4984 29460 5012
rect 28675 4981 28687 4984
rect 28629 4975 28687 4981
rect 29454 4972 29460 4984
rect 29512 4972 29518 5024
rect 30208 5012 30236 5052
rect 31588 5021 31616 5188
rect 32309 5185 32321 5188
rect 32355 5185 32367 5219
rect 32309 5179 32367 5185
rect 32585 5219 32643 5225
rect 32585 5185 32597 5219
rect 32631 5216 32643 5219
rect 32766 5216 32772 5228
rect 32631 5188 32772 5216
rect 32631 5185 32643 5188
rect 32585 5179 32643 5185
rect 32766 5176 32772 5188
rect 32824 5176 32830 5228
rect 35621 5219 35679 5225
rect 35621 5216 35633 5219
rect 35176 5188 35633 5216
rect 33778 5108 33784 5160
rect 33836 5148 33842 5160
rect 35176 5148 35204 5188
rect 35621 5185 35633 5188
rect 35667 5216 35679 5219
rect 36078 5216 36084 5228
rect 35667 5188 36084 5216
rect 35667 5185 35679 5188
rect 35621 5179 35679 5185
rect 36078 5176 36084 5188
rect 36136 5176 36142 5228
rect 37645 5219 37703 5225
rect 37645 5185 37657 5219
rect 37691 5216 37703 5219
rect 38580 5216 38608 5244
rect 38746 5216 38752 5228
rect 37691 5188 38608 5216
rect 38707 5188 38752 5216
rect 37691 5185 37703 5188
rect 37645 5179 37703 5185
rect 38746 5176 38752 5188
rect 38804 5176 38810 5228
rect 33836 5120 35204 5148
rect 33836 5108 33842 5120
rect 35250 5108 35256 5160
rect 35308 5148 35314 5160
rect 35308 5120 35353 5148
rect 35308 5108 35314 5120
rect 36906 5108 36912 5160
rect 36964 5148 36970 5160
rect 38856 5148 38884 5256
rect 38933 5219 38991 5225
rect 38933 5185 38945 5219
rect 38979 5185 38991 5219
rect 38933 5179 38991 5185
rect 36964 5120 38884 5148
rect 36964 5108 36970 5120
rect 31754 5040 31760 5092
rect 31812 5080 31818 5092
rect 33045 5083 33103 5089
rect 33045 5080 33057 5083
rect 31812 5052 33057 5080
rect 31812 5040 31818 5052
rect 33045 5049 33057 5052
rect 33091 5049 33103 5083
rect 33045 5043 33103 5049
rect 31573 5015 31631 5021
rect 31573 5012 31585 5015
rect 30208 4984 31585 5012
rect 31573 4981 31585 4984
rect 31619 4981 31631 5015
rect 31573 4975 31631 4981
rect 31662 4972 31668 5024
rect 31720 5012 31726 5024
rect 32125 5015 32183 5021
rect 32125 5012 32137 5015
rect 31720 4984 32137 5012
rect 31720 4972 31726 4984
rect 32125 4981 32137 4984
rect 32171 4981 32183 5015
rect 32125 4975 32183 4981
rect 33686 4972 33692 5024
rect 33744 5012 33750 5024
rect 33827 5015 33885 5021
rect 33827 5012 33839 5015
rect 33744 4984 33839 5012
rect 33744 4972 33750 4984
rect 33827 4981 33839 4984
rect 33873 4981 33885 5015
rect 33827 4975 33885 4981
rect 35618 4972 35624 5024
rect 35676 5012 35682 5024
rect 36541 5015 36599 5021
rect 36541 5012 36553 5015
rect 35676 4984 36553 5012
rect 35676 4972 35682 4984
rect 36541 4981 36553 4984
rect 36587 4981 36599 5015
rect 36541 4975 36599 4981
rect 37734 4972 37740 5024
rect 37792 5012 37798 5024
rect 38565 5015 38623 5021
rect 38565 5012 38577 5015
rect 37792 4984 38577 5012
rect 37792 4972 37798 4984
rect 38565 4981 38577 4984
rect 38611 4981 38623 5015
rect 38948 5012 38976 5179
rect 39022 5176 39028 5228
rect 39080 5216 39086 5228
rect 39080 5188 39125 5216
rect 39080 5176 39086 5188
rect 39592 5157 39620 5256
rect 40034 5244 40040 5256
rect 40092 5244 40098 5296
rect 41386 5284 41414 5324
rect 42426 5312 42432 5364
rect 42484 5352 42490 5364
rect 42521 5355 42579 5361
rect 42521 5352 42533 5355
rect 42484 5324 42533 5352
rect 42484 5312 42490 5324
rect 42521 5321 42533 5324
rect 42567 5321 42579 5355
rect 46842 5352 46848 5364
rect 42521 5315 42579 5321
rect 42628 5324 46848 5352
rect 42628 5284 42656 5324
rect 46842 5312 46848 5324
rect 46900 5312 46906 5364
rect 47578 5352 47584 5364
rect 47539 5324 47584 5352
rect 47578 5312 47584 5324
rect 47636 5352 47642 5364
rect 48682 5352 48688 5364
rect 47636 5324 48688 5352
rect 47636 5312 47642 5324
rect 48682 5312 48688 5324
rect 48740 5352 48746 5364
rect 49418 5352 49424 5364
rect 48740 5324 49424 5352
rect 48740 5312 48746 5324
rect 49418 5312 49424 5324
rect 49476 5312 49482 5364
rect 49510 5312 49516 5364
rect 49568 5352 49574 5364
rect 51442 5352 51448 5364
rect 49568 5324 51448 5352
rect 49568 5312 49574 5324
rect 51442 5312 51448 5324
rect 51500 5312 51506 5364
rect 52638 5312 52644 5364
rect 52696 5352 52702 5364
rect 52733 5355 52791 5361
rect 52733 5352 52745 5355
rect 52696 5324 52745 5352
rect 52696 5312 52702 5324
rect 52733 5321 52745 5324
rect 52779 5321 52791 5355
rect 52733 5315 52791 5321
rect 52917 5355 52975 5361
rect 52917 5321 52929 5355
rect 52963 5321 52975 5355
rect 52917 5315 52975 5321
rect 54941 5355 54999 5361
rect 54941 5321 54953 5355
rect 54987 5352 54999 5355
rect 55674 5352 55680 5364
rect 54987 5324 55680 5352
rect 54987 5321 54999 5324
rect 54941 5315 54999 5321
rect 44082 5284 44088 5296
rect 41386 5256 42656 5284
rect 39666 5176 39672 5228
rect 39724 5216 39730 5228
rect 39833 5219 39891 5225
rect 39833 5216 39845 5219
rect 39724 5188 39845 5216
rect 39724 5176 39730 5188
rect 39833 5185 39845 5188
rect 39879 5185 39891 5219
rect 40052 5216 40080 5244
rect 42628 5225 42656 5256
rect 43732 5256 44088 5284
rect 42613 5219 42671 5225
rect 40052 5188 41414 5216
rect 39833 5179 39891 5185
rect 39577 5151 39635 5157
rect 39577 5117 39589 5151
rect 39623 5117 39635 5151
rect 41386 5148 41414 5188
rect 42613 5185 42625 5219
rect 42659 5185 42671 5219
rect 43533 5219 43591 5225
rect 43533 5216 43545 5219
rect 42613 5179 42671 5185
rect 42720 5188 43545 5216
rect 42720 5148 42748 5188
rect 43533 5185 43545 5188
rect 43579 5216 43591 5219
rect 43732 5216 43760 5256
rect 44082 5244 44088 5256
rect 44140 5244 44146 5296
rect 44450 5244 44456 5296
rect 44508 5284 44514 5296
rect 44508 5256 45876 5284
rect 44508 5244 44514 5256
rect 43806 5225 43812 5228
rect 43579 5188 43760 5216
rect 43579 5185 43591 5188
rect 43533 5179 43591 5185
rect 43800 5179 43812 5225
rect 43864 5216 43870 5228
rect 45186 5216 45192 5228
rect 43864 5188 43900 5216
rect 44928 5188 45192 5216
rect 43806 5176 43812 5179
rect 43864 5176 43870 5188
rect 41386 5120 42748 5148
rect 39577 5111 39635 5117
rect 40586 5040 40592 5092
rect 40644 5080 40650 5092
rect 44928 5089 44956 5188
rect 45186 5176 45192 5188
rect 45244 5216 45250 5228
rect 45848 5225 45876 5256
rect 48314 5244 48320 5296
rect 48372 5284 48378 5296
rect 49436 5284 49464 5312
rect 52932 5284 52960 5315
rect 55674 5312 55680 5324
rect 55732 5312 55738 5364
rect 57330 5312 57336 5364
rect 57388 5352 57394 5364
rect 57885 5355 57943 5361
rect 57885 5352 57897 5355
rect 57388 5324 57897 5352
rect 57388 5312 57394 5324
rect 57885 5321 57897 5324
rect 57931 5321 57943 5355
rect 57885 5315 57943 5321
rect 55309 5287 55367 5293
rect 55309 5284 55321 5287
rect 48372 5256 48438 5284
rect 49436 5256 49924 5284
rect 52932 5256 55321 5284
rect 48372 5244 48378 5256
rect 45557 5219 45615 5225
rect 45557 5216 45569 5219
rect 45244 5188 45569 5216
rect 45244 5176 45250 5188
rect 45557 5185 45569 5188
rect 45603 5185 45615 5219
rect 45557 5179 45615 5185
rect 45741 5219 45799 5225
rect 45741 5185 45753 5219
rect 45787 5185 45799 5219
rect 45741 5179 45799 5185
rect 45833 5219 45891 5225
rect 45833 5185 45845 5219
rect 45879 5216 45891 5219
rect 45922 5216 45928 5228
rect 45879 5188 45928 5216
rect 45879 5185 45891 5188
rect 45833 5179 45891 5185
rect 45756 5148 45784 5179
rect 45922 5176 45928 5188
rect 45980 5176 45986 5228
rect 47029 5219 47087 5225
rect 47029 5185 47041 5219
rect 47075 5216 47087 5219
rect 47210 5216 47216 5228
rect 47075 5188 47216 5216
rect 47075 5185 47087 5188
rect 47029 5179 47087 5185
rect 47210 5176 47216 5188
rect 47268 5176 47274 5228
rect 49896 5225 49924 5256
rect 49881 5219 49939 5225
rect 49881 5185 49893 5219
rect 49927 5185 49939 5219
rect 52086 5216 52092 5228
rect 52047 5188 52092 5216
rect 49881 5179 49939 5185
rect 52086 5176 52092 5188
rect 52144 5176 52150 5228
rect 52914 5219 52972 5225
rect 52914 5185 52926 5219
rect 52960 5216 52972 5219
rect 53282 5216 53288 5228
rect 52960 5188 53288 5216
rect 52960 5185 52972 5188
rect 52914 5179 52972 5185
rect 53282 5176 53288 5188
rect 53340 5176 53346 5228
rect 54202 5216 54208 5228
rect 54163 5188 54208 5216
rect 54202 5176 54208 5188
rect 54260 5176 54266 5228
rect 54312 5225 54340 5256
rect 55309 5253 55321 5256
rect 55355 5253 55367 5287
rect 56318 5284 56324 5296
rect 55309 5247 55367 5253
rect 55876 5256 56324 5284
rect 54297 5219 54355 5225
rect 54297 5185 54309 5219
rect 54343 5185 54355 5219
rect 54297 5179 54355 5185
rect 54754 5176 54760 5228
rect 54812 5216 54818 5228
rect 54849 5219 54907 5225
rect 54849 5216 54861 5219
rect 54812 5188 54861 5216
rect 54812 5176 54818 5188
rect 54849 5185 54861 5188
rect 54895 5185 54907 5219
rect 54849 5179 54907 5185
rect 55125 5219 55183 5225
rect 55125 5185 55137 5219
rect 55171 5216 55183 5219
rect 55876 5216 55904 5256
rect 56318 5244 56324 5256
rect 56376 5244 56382 5296
rect 55171 5188 55904 5216
rect 55953 5219 56011 5225
rect 55171 5185 55183 5188
rect 55125 5179 55183 5185
rect 55953 5185 55965 5219
rect 55999 5185 56011 5219
rect 55953 5179 56011 5185
rect 46014 5148 46020 5160
rect 45756 5120 46020 5148
rect 46014 5108 46020 5120
rect 46072 5108 46078 5160
rect 46198 5108 46204 5160
rect 46256 5148 46262 5160
rect 49510 5148 49516 5160
rect 46256 5120 49516 5148
rect 46256 5108 46262 5120
rect 49510 5108 49516 5120
rect 49568 5108 49574 5160
rect 49605 5151 49663 5157
rect 49605 5117 49617 5151
rect 49651 5148 49663 5151
rect 53190 5148 53196 5160
rect 49651 5120 53196 5148
rect 49651 5117 49663 5120
rect 49605 5111 49663 5117
rect 53190 5108 53196 5120
rect 53248 5108 53254 5160
rect 53377 5151 53435 5157
rect 53377 5117 53389 5151
rect 53423 5148 53435 5151
rect 53466 5148 53472 5160
rect 53423 5120 53472 5148
rect 53423 5117 53435 5120
rect 53377 5111 53435 5117
rect 53466 5108 53472 5120
rect 53524 5108 53530 5160
rect 54021 5151 54079 5157
rect 54021 5117 54033 5151
rect 54067 5117 54079 5151
rect 54021 5111 54079 5117
rect 54113 5151 54171 5157
rect 54113 5117 54125 5151
rect 54159 5117 54171 5151
rect 54113 5111 54171 5117
rect 41417 5083 41475 5089
rect 41417 5080 41429 5083
rect 40644 5052 41429 5080
rect 40644 5040 40650 5052
rect 41417 5049 41429 5052
rect 41463 5049 41475 5083
rect 41417 5043 41475 5049
rect 44913 5083 44971 5089
rect 44913 5049 44925 5083
rect 44959 5049 44971 5083
rect 44913 5043 44971 5049
rect 52086 5040 52092 5092
rect 52144 5080 52150 5092
rect 54036 5080 54064 5111
rect 52144 5052 54064 5080
rect 54128 5080 54156 5111
rect 55214 5108 55220 5160
rect 55272 5148 55278 5160
rect 55968 5148 55996 5179
rect 56134 5176 56140 5228
rect 56192 5216 56198 5228
rect 56781 5219 56839 5225
rect 56781 5216 56793 5219
rect 56192 5188 56793 5216
rect 56192 5176 56198 5188
rect 56781 5185 56793 5188
rect 56827 5185 56839 5219
rect 58066 5216 58072 5228
rect 58027 5188 58072 5216
rect 56781 5179 56839 5185
rect 58066 5176 58072 5188
rect 58124 5176 58130 5228
rect 55272 5120 55996 5148
rect 55272 5108 55278 5120
rect 56042 5108 56048 5160
rect 56100 5148 56106 5160
rect 56100 5120 56145 5148
rect 56100 5108 56106 5120
rect 55122 5080 55128 5092
rect 54128 5052 55128 5080
rect 52144 5040 52150 5052
rect 55122 5040 55128 5052
rect 55180 5040 55186 5092
rect 56321 5083 56379 5089
rect 56321 5049 56333 5083
rect 56367 5080 56379 5083
rect 57698 5080 57704 5092
rect 56367 5052 57704 5080
rect 56367 5049 56379 5052
rect 56321 5043 56379 5049
rect 57698 5040 57704 5052
rect 57756 5040 57762 5092
rect 40310 5012 40316 5024
rect 38948 4984 40316 5012
rect 38565 4975 38623 4981
rect 40310 4972 40316 4984
rect 40368 4972 40374 5024
rect 40957 5015 41015 5021
rect 40957 4981 40969 5015
rect 41003 5012 41015 5015
rect 41046 5012 41052 5024
rect 41003 4984 41052 5012
rect 41003 4981 41015 4984
rect 40957 4975 41015 4981
rect 41046 4972 41052 4984
rect 41104 4972 41110 5024
rect 42978 4972 42984 5024
rect 43036 5012 43042 5024
rect 45373 5015 45431 5021
rect 45373 5012 45385 5015
rect 43036 4984 45385 5012
rect 43036 4972 43042 4984
rect 45373 4981 45385 4984
rect 45419 4981 45431 5015
rect 48130 5012 48136 5024
rect 48091 4984 48136 5012
rect 45373 4975 45431 4981
rect 48130 4972 48136 4984
rect 48188 4972 48194 5024
rect 50246 4972 50252 5024
rect 50304 5012 50310 5024
rect 50341 5015 50399 5021
rect 50341 5012 50353 5015
rect 50304 4984 50353 5012
rect 50304 4972 50310 4984
rect 50341 4981 50353 4984
rect 50387 4981 50399 5015
rect 50341 4975 50399 4981
rect 51074 4972 51080 5024
rect 51132 5012 51138 5024
rect 51902 5012 51908 5024
rect 51132 4984 51908 5012
rect 51132 4972 51138 4984
rect 51902 4972 51908 4984
rect 51960 4972 51966 5024
rect 51994 4972 52000 5024
rect 52052 5012 52058 5024
rect 53006 5012 53012 5024
rect 52052 4984 53012 5012
rect 52052 4972 52058 4984
rect 53006 4972 53012 4984
rect 53064 4972 53070 5024
rect 53285 5015 53343 5021
rect 53285 4981 53297 5015
rect 53331 5012 53343 5015
rect 53837 5015 53895 5021
rect 53837 5012 53849 5015
rect 53331 4984 53849 5012
rect 53331 4981 53343 4984
rect 53285 4975 53343 4981
rect 53837 4981 53849 4984
rect 53883 4981 53895 5015
rect 53837 4975 53895 4981
rect 55858 4972 55864 5024
rect 55916 5012 55922 5024
rect 56137 5015 56195 5021
rect 56137 5012 56149 5015
rect 55916 4984 56149 5012
rect 55916 4972 55922 4984
rect 56137 4981 56149 4984
rect 56183 5012 56195 5015
rect 56873 5015 56931 5021
rect 56873 5012 56885 5015
rect 56183 4984 56885 5012
rect 56183 4981 56195 4984
rect 56137 4975 56195 4981
rect 56873 4981 56885 4984
rect 56919 4981 56931 5015
rect 56873 4975 56931 4981
rect 1104 4922 58880 4944
rect 1104 4870 8174 4922
rect 8226 4870 8238 4922
rect 8290 4870 8302 4922
rect 8354 4870 8366 4922
rect 8418 4870 8430 4922
rect 8482 4870 22622 4922
rect 22674 4870 22686 4922
rect 22738 4870 22750 4922
rect 22802 4870 22814 4922
rect 22866 4870 22878 4922
rect 22930 4870 37070 4922
rect 37122 4870 37134 4922
rect 37186 4870 37198 4922
rect 37250 4870 37262 4922
rect 37314 4870 37326 4922
rect 37378 4870 51518 4922
rect 51570 4870 51582 4922
rect 51634 4870 51646 4922
rect 51698 4870 51710 4922
rect 51762 4870 51774 4922
rect 51826 4870 58880 4922
rect 1104 4848 58880 4870
rect 4341 4811 4399 4817
rect 4341 4777 4353 4811
rect 4387 4808 4399 4811
rect 4387 4780 7788 4808
rect 4387 4777 4399 4780
rect 4341 4771 4399 4777
rect 1673 4675 1731 4681
rect 1673 4641 1685 4675
rect 1719 4672 1731 4675
rect 4062 4672 4068 4684
rect 1719 4644 2728 4672
rect 1719 4641 1731 4644
rect 1673 4635 1731 4641
rect 2498 4604 2504 4616
rect 2459 4576 2504 4604
rect 2498 4564 2504 4576
rect 2556 4564 2562 4616
rect 2700 4613 2728 4644
rect 2792 4644 4068 4672
rect 2792 4613 2820 4644
rect 4062 4632 4068 4644
rect 4120 4672 4126 4684
rect 4356 4672 4384 4771
rect 6178 4700 6184 4752
rect 6236 4740 6242 4752
rect 6273 4743 6331 4749
rect 6273 4740 6285 4743
rect 6236 4712 6285 4740
rect 6236 4700 6242 4712
rect 6273 4709 6285 4712
rect 6319 4709 6331 4743
rect 7760 4740 7788 4780
rect 7926 4768 7932 4820
rect 7984 4808 7990 4820
rect 8205 4811 8263 4817
rect 8205 4808 8217 4811
rect 7984 4780 8217 4808
rect 7984 4768 7990 4780
rect 8205 4777 8217 4780
rect 8251 4777 8263 4811
rect 8205 4771 8263 4777
rect 8386 4768 8392 4820
rect 8444 4808 8450 4820
rect 10410 4808 10416 4820
rect 8444 4780 10416 4808
rect 8444 4768 8450 4780
rect 10410 4768 10416 4780
rect 10468 4768 10474 4820
rect 10778 4768 10784 4820
rect 10836 4808 10842 4820
rect 10836 4780 11008 4808
rect 10836 4768 10842 4780
rect 10594 4740 10600 4752
rect 7760 4712 10600 4740
rect 6273 4703 6331 4709
rect 10594 4700 10600 4712
rect 10652 4740 10658 4752
rect 10652 4712 10916 4740
rect 10652 4700 10658 4712
rect 6822 4672 6828 4684
rect 4120 4644 4384 4672
rect 6783 4644 6828 4672
rect 4120 4632 4126 4644
rect 6822 4632 6828 4644
rect 6880 4632 6886 4684
rect 10042 4632 10048 4684
rect 10100 4632 10106 4684
rect 10137 4675 10195 4681
rect 10137 4641 10149 4675
rect 10183 4672 10195 4675
rect 10183 4644 10824 4672
rect 10183 4641 10195 4644
rect 10137 4635 10195 4641
rect 2685 4607 2743 4613
rect 2685 4573 2697 4607
rect 2731 4573 2743 4607
rect 2685 4567 2743 4573
rect 2777 4607 2835 4613
rect 2777 4573 2789 4607
rect 2823 4573 2835 4607
rect 2777 4567 2835 4573
rect 2869 4607 2927 4613
rect 2869 4573 2881 4607
rect 2915 4604 2927 4607
rect 2958 4604 2964 4616
rect 2915 4576 2964 4604
rect 2915 4573 2927 4576
rect 2869 4567 2927 4573
rect 2958 4564 2964 4576
rect 3016 4564 3022 4616
rect 4246 4604 4252 4616
rect 4207 4576 4252 4604
rect 4246 4564 4252 4576
rect 4304 4564 4310 4616
rect 4893 4607 4951 4613
rect 4893 4573 4905 4607
rect 4939 4604 4951 4607
rect 5442 4604 5448 4616
rect 4939 4576 5448 4604
rect 4939 4573 4951 4576
rect 4893 4567 4951 4573
rect 5442 4564 5448 4576
rect 5500 4564 5506 4616
rect 7092 4607 7150 4613
rect 7092 4573 7104 4607
rect 7138 4604 7150 4607
rect 8386 4604 8392 4616
rect 7138 4576 8392 4604
rect 7138 4573 7150 4576
rect 7092 4567 7150 4573
rect 8386 4564 8392 4576
rect 8444 4564 8450 4616
rect 8570 4564 8576 4616
rect 8628 4604 8634 4616
rect 9125 4607 9183 4613
rect 9125 4604 9137 4607
rect 8628 4576 9137 4604
rect 8628 4564 8634 4576
rect 9125 4573 9137 4576
rect 9171 4573 9183 4607
rect 9125 4567 9183 4573
rect 9674 4564 9680 4616
rect 9732 4604 9738 4616
rect 9769 4607 9827 4613
rect 9769 4604 9781 4607
rect 9732 4576 9781 4604
rect 9732 4564 9738 4576
rect 9769 4573 9781 4576
rect 9815 4573 9827 4607
rect 9769 4567 9827 4573
rect 1854 4536 1860 4548
rect 1815 4508 1860 4536
rect 1854 4496 1860 4508
rect 1912 4496 1918 4548
rect 2041 4539 2099 4545
rect 2041 4505 2053 4539
rect 2087 4536 2099 4539
rect 2130 4536 2136 4548
rect 2087 4508 2136 4536
rect 2087 4505 2099 4508
rect 2041 4499 2099 4505
rect 2130 4496 2136 4508
rect 2188 4496 2194 4548
rect 5166 4545 5172 4548
rect 3145 4539 3203 4545
rect 3145 4505 3157 4539
rect 3191 4536 3203 4539
rect 3191 4508 5120 4536
rect 3191 4505 3203 4508
rect 3145 4499 3203 4505
rect 5092 4468 5120 4508
rect 5160 4499 5172 4545
rect 5224 4536 5230 4548
rect 5224 4508 5260 4536
rect 5166 4496 5172 4499
rect 5224 4496 5230 4508
rect 7558 4496 7564 4548
rect 7616 4536 7622 4548
rect 7926 4536 7932 4548
rect 7616 4508 7932 4536
rect 7616 4496 7622 4508
rect 7926 4496 7932 4508
rect 7984 4496 7990 4548
rect 8110 4496 8116 4548
rect 8168 4536 8174 4548
rect 8662 4536 8668 4548
rect 8168 4508 8668 4536
rect 8168 4496 8174 4508
rect 8662 4496 8668 4508
rect 8720 4536 8726 4548
rect 8941 4539 8999 4545
rect 8941 4536 8953 4539
rect 8720 4508 8953 4536
rect 8720 4496 8726 4508
rect 8941 4505 8953 4508
rect 8987 4505 8999 4539
rect 9490 4536 9496 4548
rect 8941 4499 8999 4505
rect 9232 4508 9496 4536
rect 5534 4468 5540 4480
rect 5092 4440 5540 4468
rect 5534 4428 5540 4440
rect 5592 4428 5598 4480
rect 6362 4428 6368 4480
rect 6420 4468 6426 4480
rect 9232 4468 9260 4508
rect 9490 4496 9496 4508
rect 9548 4496 9554 4548
rect 9953 4539 10011 4545
rect 9953 4505 9965 4539
rect 9999 4505 10011 4539
rect 10060 4536 10088 4632
rect 10796 4613 10824 4644
rect 10888 4613 10916 4712
rect 10980 4613 11008 4780
rect 12986 4768 12992 4820
rect 13044 4808 13050 4820
rect 13081 4811 13139 4817
rect 13081 4808 13093 4811
rect 13044 4780 13093 4808
rect 13044 4768 13050 4780
rect 13081 4777 13093 4780
rect 13127 4777 13139 4811
rect 13081 4771 13139 4777
rect 14090 4768 14096 4820
rect 14148 4808 14154 4820
rect 14826 4808 14832 4820
rect 14148 4780 14832 4808
rect 14148 4768 14154 4780
rect 14826 4768 14832 4780
rect 14884 4768 14890 4820
rect 17494 4768 17500 4820
rect 17552 4808 17558 4820
rect 21450 4808 21456 4820
rect 17552 4780 21456 4808
rect 17552 4768 17558 4780
rect 21450 4768 21456 4780
rect 21508 4768 21514 4820
rect 22646 4768 22652 4820
rect 22704 4808 22710 4820
rect 23106 4808 23112 4820
rect 22704 4780 23112 4808
rect 22704 4768 22710 4780
rect 23106 4768 23112 4780
rect 23164 4768 23170 4820
rect 23201 4811 23259 4817
rect 23201 4777 23213 4811
rect 23247 4808 23259 4811
rect 23382 4808 23388 4820
rect 23247 4780 23388 4808
rect 23247 4777 23259 4780
rect 23201 4771 23259 4777
rect 23382 4768 23388 4780
rect 23440 4768 23446 4820
rect 24486 4768 24492 4820
rect 24544 4808 24550 4820
rect 24581 4811 24639 4817
rect 24581 4808 24593 4811
rect 24544 4780 24593 4808
rect 24544 4768 24550 4780
rect 24581 4777 24593 4780
rect 24627 4777 24639 4811
rect 24581 4771 24639 4777
rect 25682 4768 25688 4820
rect 25740 4808 25746 4820
rect 26053 4811 26111 4817
rect 26053 4808 26065 4811
rect 25740 4780 26065 4808
rect 25740 4768 25746 4780
rect 26053 4777 26065 4780
rect 26099 4777 26111 4811
rect 26053 4771 26111 4777
rect 27798 4768 27804 4820
rect 27856 4808 27862 4820
rect 29362 4808 29368 4820
rect 27856 4780 29368 4808
rect 27856 4768 27862 4780
rect 29362 4768 29368 4780
rect 29420 4768 29426 4820
rect 30193 4811 30251 4817
rect 30193 4777 30205 4811
rect 30239 4808 30251 4811
rect 30282 4808 30288 4820
rect 30239 4780 30288 4808
rect 30239 4777 30251 4780
rect 30193 4771 30251 4777
rect 30282 4768 30288 4780
rect 30340 4768 30346 4820
rect 30745 4811 30803 4817
rect 30745 4777 30757 4811
rect 30791 4808 30803 4811
rect 30834 4808 30840 4820
rect 30791 4780 30840 4808
rect 30791 4777 30803 4780
rect 30745 4771 30803 4777
rect 30834 4768 30840 4780
rect 30892 4768 30898 4820
rect 33410 4768 33416 4820
rect 33468 4808 33474 4820
rect 35253 4811 35311 4817
rect 35253 4808 35265 4811
rect 33468 4780 35265 4808
rect 33468 4768 33474 4780
rect 35253 4777 35265 4780
rect 35299 4777 35311 4811
rect 35253 4771 35311 4777
rect 36078 4768 36084 4820
rect 36136 4808 36142 4820
rect 36633 4811 36691 4817
rect 36136 4780 36584 4808
rect 36136 4768 36142 4780
rect 17862 4740 17868 4752
rect 17823 4712 17868 4740
rect 17862 4700 17868 4712
rect 17920 4700 17926 4752
rect 20714 4700 20720 4752
rect 20772 4740 20778 4752
rect 25133 4743 25191 4749
rect 25133 4740 25145 4743
rect 20772 4712 25145 4740
rect 20772 4700 20778 4712
rect 25133 4709 25145 4712
rect 25179 4709 25191 4743
rect 25133 4703 25191 4709
rect 25406 4700 25412 4752
rect 25464 4740 25470 4752
rect 34146 4740 34152 4752
rect 25464 4712 29868 4740
rect 34107 4712 34152 4740
rect 25464 4700 25470 4712
rect 11698 4672 11704 4684
rect 11659 4644 11704 4672
rect 11698 4632 11704 4644
rect 11756 4632 11762 4684
rect 14182 4672 14188 4684
rect 14095 4644 14188 4672
rect 14182 4632 14188 4644
rect 14240 4672 14246 4684
rect 14826 4672 14832 4684
rect 14240 4644 14832 4672
rect 14240 4632 14246 4644
rect 14826 4632 14832 4644
rect 14884 4632 14890 4684
rect 16758 4672 16764 4684
rect 16719 4644 16764 4672
rect 16758 4632 16764 4644
rect 16816 4632 16822 4684
rect 20622 4632 20628 4684
rect 20680 4672 20686 4684
rect 22278 4672 22284 4684
rect 20680 4644 22284 4672
rect 20680 4632 20686 4644
rect 22278 4632 22284 4644
rect 22336 4632 22342 4684
rect 22646 4632 22652 4684
rect 22704 4672 22710 4684
rect 23290 4672 23296 4684
rect 22704 4644 22784 4672
rect 22704 4632 22710 4644
rect 10597 4607 10655 4613
rect 10597 4573 10609 4607
rect 10643 4573 10655 4607
rect 10597 4567 10655 4573
rect 10781 4607 10839 4613
rect 10781 4573 10793 4607
rect 10827 4573 10839 4607
rect 10781 4567 10839 4573
rect 10873 4607 10931 4613
rect 10873 4573 10885 4607
rect 10919 4573 10931 4607
rect 10873 4567 10931 4573
rect 10965 4607 11023 4613
rect 10965 4573 10977 4607
rect 11011 4573 11023 4607
rect 10965 4567 11023 4573
rect 11072 4576 12112 4604
rect 10612 4536 10640 4567
rect 10060 4508 10640 4536
rect 10888 4536 10916 4567
rect 11072 4536 11100 4576
rect 10888 4508 11100 4536
rect 11241 4539 11299 4545
rect 9953 4499 10011 4505
rect 11241 4505 11253 4539
rect 11287 4536 11299 4539
rect 11946 4539 12004 4545
rect 11946 4536 11958 4539
rect 11287 4508 11958 4536
rect 11287 4505 11299 4508
rect 11241 4499 11299 4505
rect 11946 4505 11958 4508
rect 11992 4505 12004 4539
rect 12084 4536 12112 4576
rect 13998 4564 14004 4616
rect 14056 4604 14062 4616
rect 14645 4607 14703 4613
rect 14645 4604 14657 4607
rect 14056 4576 14657 4604
rect 14056 4564 14062 4576
rect 14645 4573 14657 4576
rect 14691 4604 14703 4607
rect 14918 4604 14924 4616
rect 14691 4576 14924 4604
rect 14691 4573 14703 4576
rect 14645 4567 14703 4573
rect 14918 4564 14924 4576
rect 14976 4564 14982 4616
rect 17681 4607 17739 4613
rect 17681 4604 17693 4607
rect 15028 4576 17693 4604
rect 15028 4536 15056 4576
rect 17681 4573 17693 4576
rect 17727 4573 17739 4607
rect 17681 4567 17739 4573
rect 18601 4607 18659 4613
rect 18601 4573 18613 4607
rect 18647 4573 18659 4607
rect 19518 4604 19524 4616
rect 19431 4576 19524 4604
rect 18601 4567 18659 4573
rect 16516 4539 16574 4545
rect 12084 4508 15056 4536
rect 15304 4508 16436 4536
rect 11946 4499 12004 4505
rect 6420 4440 9260 4468
rect 9309 4471 9367 4477
rect 6420 4428 6426 4440
rect 9309 4437 9321 4471
rect 9355 4468 9367 4471
rect 9858 4468 9864 4480
rect 9355 4440 9864 4468
rect 9355 4437 9367 4440
rect 9309 4431 9367 4437
rect 9858 4428 9864 4440
rect 9916 4428 9922 4480
rect 9968 4468 9996 4499
rect 12986 4468 12992 4480
rect 9968 4440 12992 4468
rect 12986 4428 12992 4440
rect 13044 4428 13050 4480
rect 13722 4428 13728 4480
rect 13780 4468 13786 4480
rect 15304 4468 15332 4508
rect 13780 4440 15332 4468
rect 15381 4471 15439 4477
rect 13780 4428 13786 4440
rect 15381 4437 15393 4471
rect 15427 4468 15439 4471
rect 15838 4468 15844 4480
rect 15427 4440 15844 4468
rect 15427 4437 15439 4440
rect 15381 4431 15439 4437
rect 15838 4428 15844 4440
rect 15896 4428 15902 4480
rect 16408 4468 16436 4508
rect 16516 4505 16528 4539
rect 16562 4536 16574 4539
rect 16666 4536 16672 4548
rect 16562 4508 16672 4536
rect 16562 4505 16574 4508
rect 16516 4499 16574 4505
rect 16666 4496 16672 4508
rect 16724 4496 16730 4548
rect 18322 4536 18328 4548
rect 18248 4508 18328 4536
rect 18248 4468 18276 4508
rect 18322 4496 18328 4508
rect 18380 4496 18386 4548
rect 18414 4468 18420 4480
rect 16408 4440 18276 4468
rect 18375 4440 18420 4468
rect 18414 4428 18420 4440
rect 18472 4428 18478 4480
rect 18616 4468 18644 4567
rect 19518 4564 19524 4576
rect 19576 4604 19582 4616
rect 20640 4604 20668 4632
rect 21358 4604 21364 4616
rect 19576 4576 20668 4604
rect 21319 4576 21364 4604
rect 19576 4564 19582 4576
rect 21358 4564 21364 4576
rect 21416 4564 21422 4616
rect 21450 4564 21456 4616
rect 21508 4604 21514 4616
rect 21634 4604 21640 4616
rect 21508 4576 21553 4604
rect 21595 4576 21640 4604
rect 21508 4564 21514 4576
rect 21634 4564 21640 4576
rect 21692 4564 21698 4616
rect 22554 4604 22560 4616
rect 22515 4576 22560 4604
rect 22554 4564 22560 4576
rect 22612 4564 22618 4616
rect 22756 4610 22784 4644
rect 22857 4644 23296 4672
rect 22857 4610 22885 4644
rect 23290 4632 23296 4644
rect 23348 4632 23354 4684
rect 23845 4675 23903 4681
rect 23845 4641 23857 4675
rect 23891 4672 23903 4675
rect 25222 4672 25228 4684
rect 23891 4644 25228 4672
rect 23891 4641 23903 4644
rect 23845 4635 23903 4641
rect 25222 4632 25228 4644
rect 25280 4632 25286 4684
rect 28442 4672 28448 4684
rect 25332 4644 28448 4672
rect 22736 4604 22794 4610
rect 22736 4570 22748 4604
rect 22782 4570 22794 4604
rect 22736 4564 22794 4570
rect 22836 4604 22894 4610
rect 22836 4570 22848 4604
rect 22882 4570 22894 4604
rect 22836 4564 22894 4570
rect 22925 4607 22983 4613
rect 22925 4573 22937 4607
rect 22971 4573 22983 4607
rect 22925 4567 22983 4573
rect 19426 4496 19432 4548
rect 19484 4536 19490 4548
rect 19766 4539 19824 4545
rect 19766 4536 19778 4539
rect 19484 4508 19778 4536
rect 19484 4496 19490 4508
rect 19766 4505 19778 4508
rect 19812 4505 19824 4539
rect 22940 4536 22968 4567
rect 23106 4564 23112 4616
rect 23164 4604 23170 4616
rect 24946 4604 24952 4616
rect 23164 4576 24952 4604
rect 23164 4564 23170 4576
rect 24946 4564 24952 4576
rect 25004 4564 25010 4616
rect 25332 4613 25360 4644
rect 28442 4632 28448 4644
rect 28500 4632 28506 4684
rect 29840 4672 29868 4712
rect 34146 4700 34152 4712
rect 34204 4700 34210 4752
rect 35710 4700 35716 4752
rect 35768 4740 35774 4752
rect 35768 4712 36400 4740
rect 35768 4700 35774 4712
rect 29840 4644 31524 4672
rect 25317 4607 25375 4613
rect 25317 4573 25329 4607
rect 25363 4573 25375 4607
rect 25317 4567 25375 4573
rect 25593 4607 25651 4613
rect 25593 4573 25605 4607
rect 25639 4604 25651 4607
rect 25958 4604 25964 4616
rect 25639 4576 25964 4604
rect 25639 4573 25651 4576
rect 25593 4567 25651 4573
rect 23198 4536 23204 4548
rect 19766 4499 19824 4505
rect 20916 4508 22600 4536
rect 22940 4508 23204 4536
rect 20162 4468 20168 4480
rect 18616 4440 20168 4468
rect 20162 4428 20168 4440
rect 20220 4428 20226 4480
rect 20916 4477 20944 4508
rect 22572 4480 22600 4508
rect 23198 4496 23204 4508
rect 23256 4496 23262 4548
rect 24026 4496 24032 4548
rect 24084 4536 24090 4548
rect 24489 4539 24547 4545
rect 24489 4536 24501 4539
rect 24084 4508 24501 4536
rect 24084 4496 24090 4508
rect 24489 4505 24501 4508
rect 24535 4505 24547 4539
rect 25332 4536 25360 4567
rect 25958 4564 25964 4576
rect 26016 4564 26022 4616
rect 26602 4604 26608 4616
rect 26563 4576 26608 4604
rect 26602 4564 26608 4576
rect 26660 4564 26666 4616
rect 28813 4607 28871 4613
rect 28813 4573 28825 4607
rect 28859 4573 28871 4607
rect 28813 4567 28871 4573
rect 29549 4607 29607 4613
rect 29549 4573 29561 4607
rect 29595 4604 29607 4607
rect 29638 4604 29644 4616
rect 29595 4576 29644 4604
rect 29595 4573 29607 4576
rect 29549 4567 29607 4573
rect 25498 4536 25504 4548
rect 24489 4499 24547 4505
rect 24596 4508 25360 4536
rect 25459 4508 25504 4536
rect 20901 4471 20959 4477
rect 20901 4437 20913 4471
rect 20947 4437 20959 4471
rect 20901 4431 20959 4437
rect 21821 4471 21879 4477
rect 21821 4437 21833 4471
rect 21867 4468 21879 4471
rect 22278 4468 22284 4480
rect 21867 4440 22284 4468
rect 21867 4437 21879 4440
rect 21821 4431 21879 4437
rect 22278 4428 22284 4440
rect 22336 4428 22342 4480
rect 22554 4428 22560 4480
rect 22612 4428 22618 4480
rect 22646 4428 22652 4480
rect 22704 4468 22710 4480
rect 24596 4468 24624 4508
rect 25498 4496 25504 4508
rect 25556 4496 25562 4548
rect 28828 4536 28856 4567
rect 29638 4564 29644 4576
rect 29696 4564 29702 4616
rect 29840 4613 29868 4644
rect 29733 4607 29791 4613
rect 29733 4573 29745 4607
rect 29779 4573 29791 4607
rect 29733 4567 29791 4573
rect 29825 4607 29883 4613
rect 29825 4573 29837 4607
rect 29871 4573 29883 4607
rect 29825 4567 29883 4573
rect 25976 4508 28856 4536
rect 22704 4440 24624 4468
rect 22704 4428 22710 4440
rect 24670 4428 24676 4480
rect 24728 4468 24734 4480
rect 25976 4468 26004 4508
rect 27890 4468 27896 4480
rect 24728 4440 26004 4468
rect 27851 4440 27896 4468
rect 24728 4428 24734 4440
rect 27890 4428 27896 4440
rect 27948 4428 27954 4480
rect 29748 4468 29776 4567
rect 29914 4564 29920 4616
rect 29972 4604 29978 4616
rect 30190 4604 30196 4616
rect 29972 4576 30196 4604
rect 29972 4564 29978 4576
rect 30190 4564 30196 4576
rect 30248 4564 30254 4616
rect 31018 4564 31024 4616
rect 31076 4604 31082 4616
rect 31496 4613 31524 4644
rect 36078 4632 36084 4684
rect 36136 4672 36142 4684
rect 36136 4644 36308 4672
rect 36136 4632 36142 4644
rect 31205 4607 31263 4613
rect 31205 4604 31217 4607
rect 31076 4576 31217 4604
rect 31076 4564 31082 4576
rect 31205 4573 31217 4576
rect 31251 4573 31263 4607
rect 31205 4567 31263 4573
rect 31389 4607 31447 4613
rect 31389 4573 31401 4607
rect 31435 4573 31447 4607
rect 31389 4567 31447 4573
rect 31481 4607 31539 4613
rect 31481 4573 31493 4607
rect 31527 4573 31539 4607
rect 31481 4567 31539 4573
rect 30282 4496 30288 4548
rect 30340 4536 30346 4548
rect 31404 4536 31432 4567
rect 30340 4508 31432 4536
rect 31496 4536 31524 4567
rect 31570 4564 31576 4616
rect 31628 4604 31634 4616
rect 31628 4576 31673 4604
rect 31628 4564 31634 4576
rect 32674 4564 32680 4616
rect 32732 4604 32738 4616
rect 32769 4607 32827 4613
rect 32769 4604 32781 4607
rect 32732 4576 32781 4604
rect 32732 4564 32738 4576
rect 32769 4573 32781 4576
rect 32815 4604 32827 4607
rect 32815 4576 34836 4604
rect 32815 4573 32827 4576
rect 32769 4567 32827 4573
rect 31754 4536 31760 4548
rect 31496 4508 31760 4536
rect 30340 4496 30346 4508
rect 31754 4496 31760 4508
rect 31812 4496 31818 4548
rect 31849 4539 31907 4545
rect 31849 4505 31861 4539
rect 31895 4536 31907 4539
rect 33014 4539 33072 4545
rect 33014 4536 33026 4539
rect 31895 4508 33026 4536
rect 31895 4505 31907 4508
rect 31849 4499 31907 4505
rect 33014 4505 33026 4508
rect 33060 4505 33072 4539
rect 33014 4499 33072 4505
rect 31662 4468 31668 4480
rect 29748 4440 31668 4468
rect 31662 4428 31668 4440
rect 31720 4428 31726 4480
rect 34808 4477 34836 4576
rect 35434 4564 35440 4616
rect 35492 4604 35498 4616
rect 36280 4613 36308 4644
rect 36372 4613 36400 4712
rect 36556 4672 36584 4780
rect 36633 4777 36645 4811
rect 36679 4808 36691 4811
rect 39666 4808 39672 4820
rect 36679 4780 39672 4808
rect 36679 4777 36691 4780
rect 36633 4771 36691 4777
rect 39666 4768 39672 4780
rect 39724 4768 39730 4820
rect 40405 4811 40463 4817
rect 40405 4777 40417 4811
rect 40451 4808 40463 4811
rect 41046 4808 41052 4820
rect 40451 4780 41052 4808
rect 40451 4777 40463 4780
rect 40405 4771 40463 4777
rect 41046 4768 41052 4780
rect 41104 4768 41110 4820
rect 43441 4811 43499 4817
rect 43441 4777 43453 4811
rect 43487 4808 43499 4811
rect 43806 4808 43812 4820
rect 43487 4780 43812 4808
rect 43487 4777 43499 4780
rect 43441 4771 43499 4777
rect 43806 4768 43812 4780
rect 43864 4768 43870 4820
rect 45186 4808 45192 4820
rect 45147 4780 45192 4808
rect 45186 4768 45192 4780
rect 45244 4768 45250 4820
rect 46934 4768 46940 4820
rect 46992 4808 46998 4820
rect 50157 4811 50215 4817
rect 50157 4808 50169 4811
rect 46992 4780 50169 4808
rect 46992 4768 46998 4780
rect 50157 4777 50169 4780
rect 50203 4777 50215 4811
rect 50157 4771 50215 4777
rect 51442 4768 51448 4820
rect 51500 4808 51506 4820
rect 51721 4811 51779 4817
rect 51721 4808 51733 4811
rect 51500 4780 51733 4808
rect 51500 4768 51506 4780
rect 51721 4777 51733 4780
rect 51767 4777 51779 4811
rect 51721 4771 51779 4777
rect 51902 4768 51908 4820
rect 51960 4808 51966 4820
rect 53282 4808 53288 4820
rect 51960 4780 52684 4808
rect 53243 4780 53288 4808
rect 51960 4768 51966 4780
rect 38657 4743 38715 4749
rect 38657 4709 38669 4743
rect 38703 4740 38715 4743
rect 38746 4740 38752 4752
rect 38703 4712 38752 4740
rect 38703 4709 38715 4712
rect 38657 4703 38715 4709
rect 38746 4700 38752 4712
rect 38804 4740 38810 4752
rect 38804 4712 40172 4740
rect 38804 4700 38810 4712
rect 36906 4672 36912 4684
rect 36556 4644 36912 4672
rect 36906 4632 36912 4644
rect 36964 4672 36970 4684
rect 37277 4675 37335 4681
rect 37277 4672 37289 4675
rect 36964 4644 37289 4672
rect 36964 4632 36970 4644
rect 37277 4641 37289 4644
rect 37323 4641 37335 4675
rect 37277 4635 37335 4641
rect 35989 4607 36047 4613
rect 35989 4604 36001 4607
rect 35492 4576 36001 4604
rect 35492 4564 35498 4576
rect 35989 4573 36001 4576
rect 36035 4573 36047 4607
rect 35989 4567 36047 4573
rect 36173 4607 36231 4613
rect 36173 4573 36185 4607
rect 36219 4573 36231 4607
rect 36173 4567 36231 4573
rect 36265 4607 36323 4613
rect 36265 4573 36277 4607
rect 36311 4573 36323 4607
rect 36265 4567 36323 4573
rect 36357 4607 36415 4613
rect 36357 4573 36369 4607
rect 36403 4573 36415 4607
rect 36357 4567 36415 4573
rect 36464 4576 38516 4604
rect 34793 4471 34851 4477
rect 34793 4437 34805 4471
rect 34839 4468 34851 4471
rect 35526 4468 35532 4480
rect 34839 4440 35532 4468
rect 34839 4437 34851 4440
rect 34793 4431 34851 4437
rect 35526 4428 35532 4440
rect 35584 4428 35590 4480
rect 36004 4468 36032 4567
rect 36188 4536 36216 4567
rect 36464 4536 36492 4576
rect 36188 4508 36492 4536
rect 37274 4496 37280 4548
rect 37332 4536 37338 4548
rect 37522 4539 37580 4545
rect 37522 4536 37534 4539
rect 37332 4508 37534 4536
rect 37332 4496 37338 4508
rect 37522 4505 37534 4508
rect 37568 4505 37580 4539
rect 38488 4536 38516 4576
rect 38654 4564 38660 4616
rect 38712 4604 38718 4616
rect 40144 4613 40172 4712
rect 41322 4700 41328 4752
rect 41380 4740 41386 4752
rect 44450 4740 44456 4752
rect 41380 4712 44456 4740
rect 41380 4700 41386 4712
rect 44450 4700 44456 4712
rect 44508 4700 44514 4752
rect 47305 4743 47363 4749
rect 47305 4740 47317 4743
rect 45204 4712 47317 4740
rect 40218 4632 40224 4684
rect 40276 4672 40282 4684
rect 40276 4644 40321 4672
rect 40276 4632 40282 4644
rect 41230 4632 41236 4684
rect 41288 4672 41294 4684
rect 41785 4675 41843 4681
rect 41785 4672 41797 4675
rect 41288 4644 41797 4672
rect 41288 4632 41294 4644
rect 41785 4641 41797 4644
rect 41831 4641 41843 4675
rect 41785 4635 41843 4641
rect 42886 4632 42892 4684
rect 42944 4672 42950 4684
rect 45204 4672 45232 4712
rect 47305 4709 47317 4712
rect 47351 4709 47363 4743
rect 52656 4740 52684 4780
rect 53282 4768 53288 4780
rect 53340 4768 53346 4820
rect 54754 4808 54760 4820
rect 54715 4780 54760 4808
rect 54754 4768 54760 4780
rect 54812 4768 54818 4820
rect 55490 4808 55496 4820
rect 55451 4780 55496 4808
rect 55490 4768 55496 4780
rect 55548 4768 55554 4820
rect 55677 4811 55735 4817
rect 55677 4777 55689 4811
rect 55723 4808 55735 4811
rect 58066 4808 58072 4820
rect 55723 4780 58072 4808
rect 55723 4777 55735 4780
rect 55677 4771 55735 4777
rect 58066 4768 58072 4780
rect 58124 4768 58130 4820
rect 53929 4743 53987 4749
rect 53929 4740 53941 4743
rect 52656 4712 53941 4740
rect 47305 4703 47363 4709
rect 53929 4709 53941 4712
rect 53975 4709 53987 4743
rect 53929 4703 53987 4709
rect 55766 4700 55772 4752
rect 55824 4740 55830 4752
rect 56229 4743 56287 4749
rect 56229 4740 56241 4743
rect 55824 4712 56241 4740
rect 55824 4700 55830 4712
rect 56229 4709 56241 4712
rect 56275 4709 56287 4743
rect 56229 4703 56287 4709
rect 42944 4644 43116 4672
rect 42944 4632 42950 4644
rect 39117 4607 39175 4613
rect 39117 4604 39129 4607
rect 38712 4576 39129 4604
rect 38712 4564 38718 4576
rect 39117 4573 39129 4576
rect 39163 4573 39175 4607
rect 39117 4567 39175 4573
rect 40129 4607 40187 4613
rect 40129 4573 40141 4607
rect 40175 4573 40187 4607
rect 41046 4604 41052 4616
rect 41007 4576 41052 4604
rect 40129 4567 40187 4573
rect 41046 4564 41052 4576
rect 41104 4564 41110 4616
rect 41322 4604 41328 4616
rect 41283 4576 41328 4604
rect 41322 4564 41328 4576
rect 41380 4564 41386 4616
rect 42794 4564 42800 4616
rect 42852 4604 42858 4616
rect 42978 4604 42984 4616
rect 42852 4576 42897 4604
rect 42939 4576 42984 4604
rect 42852 4564 42858 4576
rect 42978 4564 42984 4576
rect 43036 4564 43042 4616
rect 43088 4613 43116 4644
rect 44192 4644 45232 4672
rect 43073 4607 43131 4613
rect 43073 4573 43085 4607
rect 43119 4573 43131 4607
rect 43073 4567 43131 4573
rect 43162 4564 43168 4616
rect 43220 4604 43226 4616
rect 44192 4613 44220 4644
rect 44177 4607 44235 4613
rect 43220 4576 43265 4604
rect 43220 4564 43226 4576
rect 44177 4573 44189 4607
rect 44223 4573 44235 4607
rect 44450 4604 44456 4616
rect 44411 4576 44456 4604
rect 44177 4567 44235 4573
rect 44450 4564 44456 4576
rect 44508 4564 44514 4616
rect 45204 4613 45232 4644
rect 45370 4632 45376 4684
rect 45428 4672 45434 4684
rect 46385 4675 46443 4681
rect 46385 4672 46397 4675
rect 45428 4644 46397 4672
rect 45428 4632 45434 4644
rect 46385 4641 46397 4644
rect 46431 4641 46443 4675
rect 48682 4672 48688 4684
rect 48643 4644 48688 4672
rect 46385 4635 46443 4641
rect 48682 4632 48688 4644
rect 48740 4632 48746 4684
rect 57241 4675 57299 4681
rect 57241 4641 57253 4675
rect 57287 4672 57299 4675
rect 57790 4672 57796 4684
rect 57287 4644 57796 4672
rect 57287 4641 57299 4644
rect 57241 4635 57299 4641
rect 57790 4632 57796 4644
rect 57848 4632 57854 4684
rect 45189 4607 45247 4613
rect 45189 4573 45201 4607
rect 45235 4573 45247 4607
rect 45189 4567 45247 4573
rect 45281 4607 45339 4613
rect 45281 4573 45293 4607
rect 45327 4604 45339 4607
rect 45327 4576 45876 4604
rect 45327 4573 45339 4576
rect 45281 4567 45339 4573
rect 40405 4539 40463 4545
rect 38488 4508 40080 4536
rect 37522 4499 37580 4505
rect 37918 4468 37924 4480
rect 36004 4440 37924 4468
rect 37918 4428 37924 4440
rect 37976 4428 37982 4480
rect 39942 4468 39948 4480
rect 39903 4440 39948 4468
rect 39942 4428 39948 4440
rect 40000 4428 40006 4480
rect 40052 4468 40080 4508
rect 40405 4505 40417 4539
rect 40451 4536 40463 4539
rect 45462 4536 45468 4548
rect 40451 4508 45048 4536
rect 45423 4508 45468 4536
rect 40451 4505 40463 4508
rect 40405 4499 40463 4505
rect 40865 4471 40923 4477
rect 40865 4468 40877 4471
rect 40052 4440 40877 4468
rect 40865 4437 40877 4440
rect 40911 4437 40923 4471
rect 41230 4468 41236 4480
rect 41191 4440 41236 4468
rect 40865 4431 40923 4437
rect 41230 4428 41236 4440
rect 41288 4428 41294 4480
rect 43162 4428 43168 4480
rect 43220 4468 43226 4480
rect 43993 4471 44051 4477
rect 43993 4468 44005 4471
rect 43220 4440 44005 4468
rect 43220 4428 43226 4440
rect 43993 4437 44005 4440
rect 44039 4437 44051 4471
rect 43993 4431 44051 4437
rect 44082 4428 44088 4480
rect 44140 4468 44146 4480
rect 45020 4477 45048 4508
rect 45462 4496 45468 4508
rect 45520 4496 45526 4548
rect 45848 4536 45876 4576
rect 45922 4564 45928 4616
rect 45980 4604 45986 4616
rect 46201 4607 46259 4613
rect 45980 4576 46025 4604
rect 45980 4564 45986 4576
rect 46201 4573 46213 4607
rect 46247 4573 46259 4607
rect 48406 4604 48412 4616
rect 48464 4613 48470 4616
rect 48376 4576 48412 4604
rect 46201 4567 46259 4573
rect 46216 4536 46244 4567
rect 48406 4564 48412 4576
rect 48464 4567 48476 4613
rect 49145 4607 49203 4613
rect 49145 4604 49157 4607
rect 48516 4576 49157 4604
rect 48464 4564 48470 4567
rect 48516 4548 48544 4576
rect 49145 4573 49157 4576
rect 49191 4573 49203 4607
rect 49145 4567 49203 4573
rect 50801 4607 50859 4613
rect 50801 4573 50813 4607
rect 50847 4573 50859 4607
rect 52454 4604 52460 4616
rect 52415 4576 52460 4604
rect 50801 4567 50859 4573
rect 48314 4536 48320 4548
rect 45848 4508 48320 4536
rect 48314 4496 48320 4508
rect 48372 4496 48378 4548
rect 48498 4496 48504 4548
rect 48556 4496 48562 4548
rect 48590 4496 48596 4548
rect 48648 4536 48654 4548
rect 50816 4536 50844 4567
rect 52454 4564 52460 4576
rect 52512 4564 52518 4616
rect 52546 4564 52552 4616
rect 52604 4604 52610 4616
rect 52733 4607 52791 4613
rect 52733 4604 52745 4607
rect 52604 4576 52745 4604
rect 52604 4564 52610 4576
rect 52733 4573 52745 4576
rect 52779 4604 52791 4607
rect 53282 4604 53288 4616
rect 52779 4576 53288 4604
rect 52779 4573 52791 4576
rect 52733 4567 52791 4573
rect 53282 4564 53288 4576
rect 53340 4564 53346 4616
rect 53469 4607 53527 4613
rect 53469 4573 53481 4607
rect 53515 4604 53527 4607
rect 53558 4604 53564 4616
rect 53515 4576 53564 4604
rect 53515 4573 53527 4576
rect 53469 4567 53527 4573
rect 53558 4564 53564 4576
rect 53616 4564 53622 4616
rect 54573 4607 54631 4613
rect 54573 4573 54585 4607
rect 54619 4573 54631 4607
rect 54573 4567 54631 4573
rect 54757 4607 54815 4613
rect 54757 4573 54769 4607
rect 54803 4604 54815 4607
rect 55582 4604 55588 4616
rect 54803 4576 55588 4604
rect 54803 4573 54815 4576
rect 54757 4567 54815 4573
rect 48648 4508 50844 4536
rect 54588 4536 54616 4567
rect 55582 4564 55588 4576
rect 55640 4604 55646 4616
rect 55950 4604 55956 4616
rect 55640 4576 55956 4604
rect 55640 4564 55646 4576
rect 55950 4564 55956 4576
rect 56008 4564 56014 4616
rect 56965 4607 57023 4613
rect 56965 4573 56977 4607
rect 57011 4573 57023 4607
rect 57698 4604 57704 4616
rect 57659 4576 57704 4604
rect 56965 4567 57023 4573
rect 55122 4536 55128 4548
rect 54588 4508 55128 4536
rect 48648 4496 48654 4508
rect 55122 4496 55128 4508
rect 55180 4536 55186 4548
rect 55309 4539 55367 4545
rect 55309 4536 55321 4539
rect 55180 4508 55321 4536
rect 55180 4496 55186 4508
rect 55309 4505 55321 4508
rect 55355 4505 55367 4539
rect 55309 4499 55367 4505
rect 44361 4471 44419 4477
rect 44361 4468 44373 4471
rect 44140 4440 44373 4468
rect 44140 4428 44146 4440
rect 44361 4437 44373 4440
rect 44407 4437 44419 4471
rect 44361 4431 44419 4437
rect 45005 4471 45063 4477
rect 45005 4437 45017 4471
rect 45051 4437 45063 4471
rect 45005 4431 45063 4437
rect 46014 4428 46020 4480
rect 46072 4468 46078 4480
rect 46072 4440 46117 4468
rect 46072 4428 46078 4440
rect 48130 4428 48136 4480
rect 48188 4468 48194 4480
rect 55214 4468 55220 4480
rect 48188 4440 55220 4468
rect 48188 4428 48194 4440
rect 55214 4428 55220 4440
rect 55272 4428 55278 4480
rect 55398 4428 55404 4480
rect 55456 4468 55462 4480
rect 55509 4471 55567 4477
rect 55509 4468 55521 4471
rect 55456 4440 55521 4468
rect 55456 4428 55462 4440
rect 55509 4437 55521 4440
rect 55555 4437 55567 4471
rect 56980 4468 57008 4567
rect 57698 4564 57704 4576
rect 57756 4564 57762 4616
rect 57882 4468 57888 4480
rect 56980 4440 57888 4468
rect 55509 4431 55567 4437
rect 57882 4428 57888 4440
rect 57940 4428 57946 4480
rect 1104 4378 58880 4400
rect 1104 4326 15398 4378
rect 15450 4326 15462 4378
rect 15514 4326 15526 4378
rect 15578 4326 15590 4378
rect 15642 4326 15654 4378
rect 15706 4326 29846 4378
rect 29898 4326 29910 4378
rect 29962 4326 29974 4378
rect 30026 4326 30038 4378
rect 30090 4326 30102 4378
rect 30154 4326 44294 4378
rect 44346 4326 44358 4378
rect 44410 4326 44422 4378
rect 44474 4326 44486 4378
rect 44538 4326 44550 4378
rect 44602 4326 58880 4378
rect 1104 4304 58880 4326
rect 2130 4224 2136 4276
rect 2188 4264 2194 4276
rect 4430 4264 4436 4276
rect 2188 4236 4436 4264
rect 2188 4224 2194 4236
rect 4430 4224 4436 4236
rect 4488 4264 4494 4276
rect 6362 4264 6368 4276
rect 4488 4236 6368 4264
rect 4488 4224 4494 4236
rect 6362 4224 6368 4236
rect 6420 4224 6426 4276
rect 7466 4264 7472 4276
rect 7427 4236 7472 4264
rect 7466 4224 7472 4236
rect 7524 4224 7530 4276
rect 7742 4224 7748 4276
rect 7800 4264 7806 4276
rect 8021 4267 8079 4273
rect 8021 4264 8033 4267
rect 7800 4236 8033 4264
rect 7800 4224 7806 4236
rect 8021 4233 8033 4236
rect 8067 4264 8079 4267
rect 17218 4264 17224 4276
rect 8067 4236 10272 4264
rect 8067 4233 8079 4236
rect 8021 4227 8079 4233
rect 5629 4199 5687 4205
rect 5629 4165 5641 4199
rect 5675 4196 5687 4199
rect 6270 4196 6276 4208
rect 5675 4168 6276 4196
rect 5675 4165 5687 4168
rect 5629 4159 5687 4165
rect 6270 4156 6276 4168
rect 6328 4156 6334 4208
rect 7098 4156 7104 4208
rect 7156 4196 7162 4208
rect 7558 4196 7564 4208
rect 7156 4168 7564 4196
rect 7156 4156 7162 4168
rect 7558 4156 7564 4168
rect 7616 4156 7622 4208
rect 10137 4199 10195 4205
rect 10137 4165 10149 4199
rect 10183 4165 10195 4199
rect 10137 4159 10195 4165
rect 1762 4088 1768 4140
rect 1820 4128 1826 4140
rect 1857 4131 1915 4137
rect 1857 4128 1869 4131
rect 1820 4100 1869 4128
rect 1820 4088 1826 4100
rect 1857 4097 1869 4100
rect 1903 4097 1915 4131
rect 1857 4091 1915 4097
rect 2682 4088 2688 4140
rect 2740 4132 2746 4140
rect 2777 4132 2835 4137
rect 2740 4131 2835 4132
rect 2740 4104 2789 4131
rect 2740 4088 2746 4104
rect 2777 4097 2789 4104
rect 2823 4097 2835 4131
rect 2777 4091 2835 4097
rect 2869 4134 2927 4140
rect 2869 4100 2881 4134
rect 2915 4100 2927 4134
rect 2869 4094 2927 4100
rect 2038 4020 2044 4072
rect 2096 4060 2102 4072
rect 2884 4060 2912 4094
rect 2958 4088 2964 4140
rect 3016 4128 3022 4140
rect 3145 4131 3203 4137
rect 3016 4100 3061 4128
rect 3016 4088 3022 4100
rect 3145 4097 3157 4131
rect 3191 4128 3203 4131
rect 3234 4128 3240 4140
rect 3191 4100 3240 4128
rect 3191 4097 3203 4100
rect 3145 4091 3203 4097
rect 3234 4088 3240 4100
rect 3292 4088 3298 4140
rect 4338 4128 4344 4140
rect 4299 4100 4344 4128
rect 4338 4088 4344 4100
rect 4396 4088 4402 4140
rect 4890 4088 4896 4140
rect 4948 4128 4954 4140
rect 5077 4131 5135 4137
rect 5077 4128 5089 4131
rect 4948 4100 5089 4128
rect 4948 4088 4954 4100
rect 5077 4097 5089 4100
rect 5123 4097 5135 4131
rect 5077 4091 5135 4097
rect 5166 4088 5172 4140
rect 5224 4088 5230 4140
rect 6638 4088 6644 4140
rect 6696 4128 6702 4140
rect 6733 4131 6791 4137
rect 6733 4128 6745 4131
rect 6696 4100 6745 4128
rect 6696 4088 6702 4100
rect 6733 4097 6745 4100
rect 6779 4097 6791 4131
rect 7282 4128 7288 4140
rect 7243 4100 7288 4128
rect 6733 4091 6791 4097
rect 7282 4088 7288 4100
rect 7340 4088 7346 4140
rect 7469 4131 7527 4137
rect 7469 4097 7481 4131
rect 7515 4128 7527 4131
rect 8754 4128 8760 4140
rect 7515 4100 8760 4128
rect 7515 4097 7527 4100
rect 7469 4091 7527 4097
rect 8754 4088 8760 4100
rect 8812 4088 8818 4140
rect 9145 4131 9203 4137
rect 9145 4097 9157 4131
rect 9191 4128 9203 4131
rect 10152 4128 10180 4159
rect 9191 4100 10180 4128
rect 10244 4128 10272 4236
rect 10704 4236 17224 4264
rect 10367 4131 10425 4137
rect 10367 4128 10379 4131
rect 10244 4100 10379 4128
rect 9191 4097 9203 4100
rect 9145 4091 9203 4097
rect 10367 4097 10379 4100
rect 10413 4097 10425 4131
rect 10502 4128 10508 4140
rect 10463 4100 10508 4128
rect 10367 4091 10425 4097
rect 10502 4088 10508 4100
rect 10560 4088 10566 4140
rect 10618 4131 10676 4137
rect 10618 4097 10630 4131
rect 10664 4128 10676 4131
rect 10704 4128 10732 4236
rect 17218 4224 17224 4236
rect 17276 4224 17282 4276
rect 19426 4264 19432 4276
rect 19387 4236 19432 4264
rect 19426 4224 19432 4236
rect 19484 4224 19490 4276
rect 21358 4224 21364 4276
rect 21416 4264 21422 4276
rect 24210 4264 24216 4276
rect 21416 4236 24216 4264
rect 21416 4224 21422 4236
rect 24210 4224 24216 4236
rect 24268 4224 24274 4276
rect 24578 4224 24584 4276
rect 24636 4264 24642 4276
rect 25869 4267 25927 4273
rect 25869 4264 25881 4267
rect 24636 4236 25881 4264
rect 24636 4224 24642 4236
rect 25869 4233 25881 4236
rect 25915 4264 25927 4267
rect 28537 4267 28595 4273
rect 25915 4236 27660 4264
rect 25915 4233 25927 4236
rect 25869 4227 25927 4233
rect 10962 4196 10968 4208
rect 10796 4168 10968 4196
rect 10796 4137 10824 4168
rect 10962 4156 10968 4168
rect 11020 4196 11026 4208
rect 13170 4196 13176 4208
rect 11020 4168 13176 4196
rect 11020 4156 11026 4168
rect 13170 4156 13176 4168
rect 13228 4156 13234 4208
rect 13725 4199 13783 4205
rect 13725 4196 13737 4199
rect 13280 4168 13737 4196
rect 10664 4100 10732 4128
rect 10781 4131 10839 4137
rect 10664 4097 10676 4100
rect 10618 4091 10676 4097
rect 10781 4097 10793 4131
rect 10827 4097 10839 4131
rect 10781 4091 10839 4097
rect 11784 4131 11842 4137
rect 11784 4097 11796 4131
rect 11830 4128 11842 4131
rect 13280 4128 13308 4168
rect 13725 4165 13737 4168
rect 13771 4165 13783 4199
rect 14826 4196 14832 4208
rect 14787 4168 14832 4196
rect 13725 4159 13783 4165
rect 14826 4156 14832 4168
rect 14884 4156 14890 4208
rect 14918 4156 14924 4208
rect 14976 4196 14982 4208
rect 15013 4199 15071 4205
rect 15013 4196 15025 4199
rect 14976 4168 15025 4196
rect 14976 4156 14982 4168
rect 15013 4165 15025 4168
rect 15059 4165 15071 4199
rect 15013 4159 15071 4165
rect 15102 4156 15108 4208
rect 15160 4196 15166 4208
rect 16758 4196 16764 4208
rect 15160 4168 16764 4196
rect 15160 4156 15166 4168
rect 16758 4156 16764 4168
rect 16816 4196 16822 4208
rect 18138 4196 18144 4208
rect 16816 4168 16896 4196
rect 18099 4168 18144 4196
rect 16816 4156 16822 4168
rect 11830 4100 13308 4128
rect 11830 4097 11842 4100
rect 11784 4091 11842 4097
rect 13814 4088 13820 4140
rect 13872 4128 13878 4140
rect 14087 4137 14093 4140
rect 13955 4131 14013 4137
rect 13955 4128 13967 4131
rect 13872 4100 13967 4128
rect 13872 4088 13878 4100
rect 13955 4097 13967 4100
rect 14001 4097 14013 4131
rect 13955 4091 14013 4097
rect 14074 4131 14093 4137
rect 14074 4097 14086 4131
rect 14074 4091 14093 4097
rect 14087 4088 14093 4091
rect 14145 4088 14151 4140
rect 14182 4088 14188 4140
rect 14240 4137 14246 4140
rect 14240 4128 14248 4137
rect 14240 4100 14285 4128
rect 14240 4091 14248 4100
rect 14240 4088 14246 4091
rect 14366 4088 14372 4140
rect 14424 4128 14430 4140
rect 15838 4128 15844 4140
rect 14424 4100 14469 4128
rect 15799 4100 15844 4128
rect 14424 4088 14430 4100
rect 15838 4088 15844 4100
rect 15896 4088 15902 4140
rect 16025 4131 16083 4137
rect 16025 4097 16037 4131
rect 16071 4097 16083 4131
rect 16025 4091 16083 4097
rect 16117 4131 16175 4137
rect 16117 4097 16129 4131
rect 16163 4128 16175 4131
rect 16298 4128 16304 4140
rect 16163 4100 16304 4128
rect 16163 4097 16175 4100
rect 16117 4091 16175 4097
rect 2096 4032 2912 4060
rect 2096 4020 2102 4032
rect 2501 3995 2559 4001
rect 2501 3961 2513 3995
rect 2547 3992 2559 3995
rect 5184 3992 5212 4088
rect 5258 4020 5264 4072
rect 5316 4060 5322 4072
rect 9401 4063 9459 4069
rect 5316 4032 8432 4060
rect 5316 4020 5322 4032
rect 5810 3992 5816 4004
rect 2547 3964 2774 3992
rect 2547 3961 2559 3964
rect 2501 3955 2559 3961
rect 2041 3927 2099 3933
rect 2041 3893 2053 3927
rect 2087 3924 2099 3927
rect 2130 3924 2136 3936
rect 2087 3896 2136 3924
rect 2087 3893 2099 3896
rect 2041 3887 2099 3893
rect 2130 3884 2136 3896
rect 2188 3884 2194 3936
rect 2746 3924 2774 3964
rect 3804 3964 5212 3992
rect 5771 3964 5816 3992
rect 3804 3924 3832 3964
rect 5810 3952 5816 3964
rect 5868 3952 5874 4004
rect 7466 3952 7472 4004
rect 7524 3992 7530 4004
rect 8110 3992 8116 4004
rect 7524 3964 8116 3992
rect 7524 3952 7530 3964
rect 8110 3952 8116 3964
rect 8168 3952 8174 4004
rect 2746 3896 3832 3924
rect 4157 3927 4215 3933
rect 4157 3893 4169 3927
rect 4203 3924 4215 3927
rect 4798 3924 4804 3936
rect 4203 3896 4804 3924
rect 4203 3893 4215 3896
rect 4157 3887 4215 3893
rect 4798 3884 4804 3896
rect 4856 3884 4862 3936
rect 4890 3884 4896 3936
rect 4948 3924 4954 3936
rect 6549 3927 6607 3933
rect 4948 3896 4993 3924
rect 4948 3884 4954 3896
rect 6549 3893 6561 3927
rect 6595 3924 6607 3927
rect 7742 3924 7748 3936
rect 6595 3896 7748 3924
rect 6595 3893 6607 3896
rect 6549 3887 6607 3893
rect 7742 3884 7748 3896
rect 7800 3884 7806 3936
rect 8404 3924 8432 4032
rect 9401 4029 9413 4063
rect 9447 4060 9459 4063
rect 11514 4060 11520 4072
rect 9447 4032 11520 4060
rect 9447 4029 9459 4032
rect 9401 4023 9459 4029
rect 9416 3924 9444 4023
rect 11514 4020 11520 4032
rect 11572 4020 11578 4072
rect 16040 4060 16068 4091
rect 16298 4088 16304 4100
rect 16356 4088 16362 4140
rect 16868 4118 16896 4168
rect 18138 4156 18144 4168
rect 18196 4156 18202 4208
rect 23290 4196 23296 4208
rect 19076 4168 23296 4196
rect 17031 4137 17037 4140
rect 16925 4131 16983 4137
rect 16925 4118 16937 4131
rect 16868 4097 16937 4118
rect 16971 4128 16983 4131
rect 17018 4131 17037 4137
rect 16971 4097 16988 4128
rect 16868 4090 16988 4097
rect 17018 4097 17030 4131
rect 17018 4091 17037 4097
rect 17031 4088 17037 4091
rect 17089 4088 17095 4140
rect 17134 4131 17192 4137
rect 17134 4097 17146 4131
rect 17180 4097 17192 4131
rect 17134 4091 17192 4097
rect 17313 4131 17371 4137
rect 17313 4097 17325 4131
rect 17359 4097 17371 4131
rect 17313 4091 17371 4097
rect 16390 4060 16396 4072
rect 16040 4032 16396 4060
rect 16390 4020 16396 4032
rect 16448 4020 16454 4072
rect 16666 4060 16672 4072
rect 16627 4032 16672 4060
rect 16666 4020 16672 4032
rect 16724 4020 16730 4072
rect 12897 3995 12955 4001
rect 12897 3961 12909 3995
rect 12943 3992 12955 3995
rect 15657 3995 15715 4001
rect 12943 3964 15608 3992
rect 12943 3961 12955 3964
rect 12897 3955 12955 3961
rect 8404 3896 9444 3924
rect 13814 3884 13820 3936
rect 13872 3924 13878 3936
rect 14918 3924 14924 3936
rect 13872 3896 14924 3924
rect 13872 3884 13878 3896
rect 14918 3884 14924 3896
rect 14976 3884 14982 3936
rect 15580 3924 15608 3964
rect 15657 3961 15669 3995
rect 15703 3992 15715 3995
rect 17144 3992 17172 4091
rect 17328 4060 17356 4091
rect 17954 4088 17960 4140
rect 18012 4128 18018 4140
rect 19076 4137 19104 4168
rect 23290 4156 23296 4168
rect 23348 4196 23354 4208
rect 25406 4196 25412 4208
rect 23348 4168 25412 4196
rect 23348 4156 23354 4168
rect 18785 4131 18843 4137
rect 18785 4128 18797 4131
rect 18012 4100 18797 4128
rect 18012 4088 18018 4100
rect 18785 4097 18797 4100
rect 18831 4097 18843 4131
rect 18785 4091 18843 4097
rect 18969 4131 19027 4137
rect 18969 4097 18981 4131
rect 19015 4097 19027 4131
rect 18969 4091 19027 4097
rect 19061 4131 19119 4137
rect 19061 4097 19073 4131
rect 19107 4097 19119 4131
rect 19061 4091 19119 4097
rect 17586 4060 17592 4072
rect 17328 4032 17592 4060
rect 17586 4020 17592 4032
rect 17644 4060 17650 4072
rect 18325 4063 18383 4069
rect 18325 4060 18337 4063
rect 17644 4032 18337 4060
rect 17644 4020 17650 4032
rect 18325 4029 18337 4032
rect 18371 4029 18383 4063
rect 18984 4060 19012 4091
rect 19150 4088 19156 4140
rect 19208 4128 19214 4140
rect 20714 4128 20720 4140
rect 19208 4100 19253 4128
rect 19306 4100 20720 4128
rect 19208 4088 19214 4100
rect 19306 4060 19334 4100
rect 20714 4088 20720 4100
rect 20772 4088 20778 4140
rect 21013 4131 21071 4137
rect 21013 4097 21025 4131
rect 21059 4128 21071 4131
rect 21269 4131 21327 4137
rect 21059 4100 21220 4128
rect 21059 4097 21071 4100
rect 21013 4091 21071 4097
rect 18984 4032 19334 4060
rect 21192 4060 21220 4100
rect 21269 4097 21281 4131
rect 21315 4128 21327 4131
rect 21726 4128 21732 4140
rect 21315 4100 21732 4128
rect 21315 4097 21327 4100
rect 21269 4091 21327 4097
rect 21726 4088 21732 4100
rect 21784 4088 21790 4140
rect 22097 4131 22155 4137
rect 22097 4097 22109 4131
rect 22143 4097 22155 4131
rect 22097 4091 22155 4097
rect 22189 4131 22247 4137
rect 22189 4097 22201 4131
rect 22235 4097 22247 4131
rect 22189 4091 22247 4097
rect 21821 4063 21879 4069
rect 21821 4060 21833 4063
rect 21192 4032 21833 4060
rect 18325 4023 18383 4029
rect 21821 4029 21833 4032
rect 21867 4029 21879 4063
rect 21821 4023 21879 4029
rect 15703 3964 17172 3992
rect 15703 3961 15715 3964
rect 15657 3955 15715 3961
rect 16574 3924 16580 3936
rect 15580 3896 16580 3924
rect 16574 3884 16580 3896
rect 16632 3884 16638 3936
rect 18340 3924 18368 4023
rect 22112 3992 22140 4091
rect 22204 4060 22232 4091
rect 22278 4088 22284 4140
rect 22336 4128 22342 4140
rect 22465 4131 22523 4137
rect 22336 4100 22381 4128
rect 22336 4088 22342 4100
rect 22465 4097 22477 4131
rect 22511 4128 22523 4131
rect 23658 4128 23664 4140
rect 22511 4100 23664 4128
rect 22511 4097 22523 4100
rect 22465 4091 22523 4097
rect 23658 4088 23664 4100
rect 23716 4088 23722 4140
rect 23845 4131 23903 4137
rect 23845 4097 23857 4131
rect 23891 4128 23903 4131
rect 23934 4128 23940 4140
rect 23891 4100 23940 4128
rect 23891 4097 23903 4100
rect 23845 4091 23903 4097
rect 23934 4088 23940 4100
rect 23992 4088 23998 4140
rect 24486 4088 24492 4140
rect 24544 4128 24550 4140
rect 24673 4131 24731 4137
rect 24673 4128 24685 4131
rect 24544 4100 24685 4128
rect 24544 4088 24550 4100
rect 24673 4097 24685 4100
rect 24719 4097 24731 4131
rect 24673 4091 24731 4097
rect 24762 4088 24768 4140
rect 24820 4134 24826 4140
rect 24964 4137 24992 4168
rect 25406 4156 25412 4168
rect 25464 4156 25470 4208
rect 27522 4196 27528 4208
rect 27172 4168 27528 4196
rect 24857 4134 24915 4137
rect 24820 4131 24915 4134
rect 24820 4106 24869 4131
rect 24820 4088 24826 4106
rect 24857 4097 24869 4106
rect 24903 4097 24915 4131
rect 24857 4091 24915 4097
rect 24949 4131 25007 4137
rect 24949 4097 24961 4131
rect 24995 4097 25007 4131
rect 24949 4091 25007 4097
rect 25038 4088 25044 4140
rect 25096 4128 25102 4140
rect 25774 4128 25780 4140
rect 25096 4100 25141 4128
rect 25735 4100 25780 4128
rect 25096 4088 25102 4100
rect 25774 4088 25780 4100
rect 25832 4088 25838 4140
rect 26050 4128 26056 4140
rect 26011 4100 26056 4128
rect 26050 4088 26056 4100
rect 26108 4088 26114 4140
rect 27172 4137 27200 4168
rect 27522 4156 27528 4168
rect 27580 4156 27586 4208
rect 27157 4131 27215 4137
rect 27157 4097 27169 4131
rect 27203 4097 27215 4131
rect 27413 4131 27471 4137
rect 27413 4128 27425 4131
rect 27157 4091 27215 4097
rect 27264 4100 27425 4128
rect 22370 4060 22376 4072
rect 22204 4032 22376 4060
rect 22370 4020 22376 4032
rect 22428 4060 22434 4072
rect 23106 4060 23112 4072
rect 22428 4032 23112 4060
rect 22428 4020 22434 4032
rect 23106 4020 23112 4032
rect 23164 4020 23170 4072
rect 25056 3992 25084 4088
rect 25317 4063 25375 4069
rect 25317 4029 25329 4063
rect 25363 4060 25375 4063
rect 27264 4060 27292 4100
rect 27413 4097 27425 4100
rect 27459 4097 27471 4131
rect 27632 4128 27660 4236
rect 28537 4233 28549 4267
rect 28583 4264 28595 4267
rect 28718 4264 28724 4276
rect 28583 4236 28724 4264
rect 28583 4233 28595 4236
rect 28537 4227 28595 4233
rect 28718 4224 28724 4236
rect 28776 4224 28782 4276
rect 31018 4224 31024 4276
rect 31076 4264 31082 4276
rect 31938 4264 31944 4276
rect 31076 4236 31944 4264
rect 31076 4224 31082 4236
rect 31938 4224 31944 4236
rect 31996 4224 32002 4276
rect 32766 4264 32772 4276
rect 32048 4236 32772 4264
rect 27982 4156 27988 4208
rect 28040 4196 28046 4208
rect 28040 4168 29316 4196
rect 28040 4156 28046 4168
rect 28997 4131 29055 4137
rect 28997 4128 29009 4131
rect 27632 4100 29009 4128
rect 27413 4091 27471 4097
rect 28997 4097 29009 4100
rect 29043 4097 29055 4131
rect 28997 4091 29055 4097
rect 29181 4131 29239 4137
rect 29181 4097 29193 4131
rect 29227 4097 29239 4131
rect 29288 4128 29316 4168
rect 29362 4156 29368 4208
rect 29420 4196 29426 4208
rect 31294 4196 31300 4208
rect 29420 4168 31300 4196
rect 29420 4156 29426 4168
rect 29932 4137 29960 4168
rect 31294 4156 31300 4168
rect 31352 4156 31358 4208
rect 29825 4131 29883 4137
rect 29825 4128 29837 4131
rect 29288 4100 29837 4128
rect 29181 4091 29239 4097
rect 29825 4097 29837 4100
rect 29871 4097 29883 4131
rect 29825 4091 29883 4097
rect 29917 4131 29975 4137
rect 29917 4097 29929 4131
rect 29963 4097 29975 4131
rect 30098 4128 30104 4140
rect 30059 4100 30104 4128
rect 29917 4091 29975 4097
rect 25363 4032 27292 4060
rect 25363 4029 25375 4032
rect 25317 4023 25375 4029
rect 29196 3992 29224 4091
rect 29840 4060 29868 4091
rect 30098 4088 30104 4100
rect 30156 4088 30162 4140
rect 30282 4128 30288 4140
rect 30243 4100 30288 4128
rect 30282 4088 30288 4100
rect 30340 4088 30346 4140
rect 32048 4128 32076 4236
rect 32766 4224 32772 4236
rect 32824 4224 32830 4276
rect 37274 4264 37280 4276
rect 37235 4236 37280 4264
rect 37274 4224 37280 4236
rect 37332 4224 37338 4276
rect 40310 4224 40316 4276
rect 40368 4264 40374 4276
rect 41230 4264 41236 4276
rect 40368 4236 41236 4264
rect 40368 4224 40374 4236
rect 41230 4224 41236 4236
rect 41288 4264 41294 4276
rect 43990 4264 43996 4276
rect 41288 4236 43996 4264
rect 41288 4224 41294 4236
rect 43990 4224 43996 4236
rect 44048 4264 44054 4276
rect 46014 4264 46020 4276
rect 44048 4236 46020 4264
rect 44048 4224 44054 4236
rect 46014 4224 46020 4236
rect 46072 4224 46078 4276
rect 48314 4264 48320 4276
rect 48275 4236 48320 4264
rect 48314 4224 48320 4236
rect 48372 4224 48378 4276
rect 51994 4224 52000 4276
rect 52052 4224 52058 4276
rect 53558 4224 53564 4276
rect 53616 4264 53622 4276
rect 57974 4264 57980 4276
rect 53616 4236 57980 4264
rect 53616 4224 53622 4236
rect 57974 4224 57980 4236
rect 58032 4224 58038 4276
rect 32674 4196 32680 4208
rect 32140 4168 32680 4196
rect 32140 4137 32168 4168
rect 32674 4156 32680 4168
rect 32732 4156 32738 4208
rect 32858 4156 32864 4208
rect 32916 4196 32922 4208
rect 35802 4196 35808 4208
rect 32916 4168 35808 4196
rect 32916 4156 32922 4168
rect 30392 4100 32076 4128
rect 32125 4131 32183 4137
rect 30392 4060 30420 4100
rect 32125 4097 32137 4131
rect 32171 4097 32183 4131
rect 32125 4091 32183 4097
rect 32214 4088 32220 4140
rect 32272 4128 32278 4140
rect 32381 4131 32439 4137
rect 32381 4128 32393 4131
rect 32272 4100 32393 4128
rect 32272 4088 32278 4100
rect 32381 4097 32393 4100
rect 32427 4097 32439 4131
rect 32381 4091 32439 4097
rect 32766 4088 32772 4140
rect 32824 4128 32830 4140
rect 34241 4131 34299 4137
rect 34241 4128 34253 4131
rect 32824 4100 34253 4128
rect 32824 4088 32830 4100
rect 34241 4097 34253 4100
rect 34287 4097 34299 4131
rect 34241 4091 34299 4097
rect 34606 4088 34612 4140
rect 34664 4128 34670 4140
rect 35066 4128 35072 4140
rect 34664 4100 35072 4128
rect 34664 4088 34670 4100
rect 35066 4088 35072 4100
rect 35124 4128 35130 4140
rect 35544 4137 35572 4168
rect 35802 4156 35808 4168
rect 35860 4156 35866 4208
rect 40034 4156 40040 4208
rect 40092 4196 40098 4208
rect 40954 4196 40960 4208
rect 40092 4168 40960 4196
rect 40092 4156 40098 4168
rect 40954 4156 40960 4168
rect 41012 4156 41018 4208
rect 45370 4196 45376 4208
rect 42996 4168 44128 4196
rect 35253 4131 35311 4137
rect 35253 4128 35265 4131
rect 35124 4100 35265 4128
rect 35124 4088 35130 4100
rect 35253 4097 35265 4100
rect 35299 4097 35311 4131
rect 35253 4091 35311 4097
rect 35437 4131 35495 4137
rect 35437 4097 35449 4131
rect 35483 4097 35495 4131
rect 35437 4091 35495 4097
rect 35529 4131 35587 4137
rect 35529 4097 35541 4131
rect 35575 4097 35587 4131
rect 35529 4091 35587 4097
rect 35621 4131 35679 4137
rect 35621 4097 35633 4131
rect 35667 4128 35679 4131
rect 35710 4128 35716 4140
rect 35667 4100 35716 4128
rect 35667 4097 35679 4100
rect 35621 4091 35679 4097
rect 31294 4060 31300 4072
rect 29840 4032 30420 4060
rect 31255 4032 31300 4060
rect 31294 4020 31300 4032
rect 31352 4020 31358 4072
rect 31570 4060 31576 4072
rect 31531 4032 31576 4060
rect 31570 4020 31576 4032
rect 31628 4020 31634 4072
rect 33594 4060 33600 4072
rect 33336 4032 33600 4060
rect 29270 3992 29276 4004
rect 22112 3964 25084 3992
rect 29183 3964 29276 3992
rect 29270 3952 29276 3964
rect 29328 3992 29334 4004
rect 29328 3964 31754 3992
rect 29328 3952 29334 3964
rect 18874 3924 18880 3936
rect 18340 3896 18880 3924
rect 18874 3884 18880 3896
rect 18932 3884 18938 3936
rect 19886 3924 19892 3936
rect 19847 3896 19892 3924
rect 19886 3884 19892 3896
rect 19944 3924 19950 3936
rect 21634 3924 21640 3936
rect 19944 3896 21640 3924
rect 19944 3884 19950 3896
rect 21634 3884 21640 3896
rect 21692 3884 21698 3936
rect 23293 3927 23351 3933
rect 23293 3893 23305 3927
rect 23339 3924 23351 3927
rect 23566 3924 23572 3936
rect 23339 3896 23572 3924
rect 23339 3893 23351 3896
rect 23293 3887 23351 3893
rect 23566 3884 23572 3896
rect 23624 3884 23630 3936
rect 23658 3884 23664 3936
rect 23716 3924 23722 3936
rect 23937 3927 23995 3933
rect 23937 3924 23949 3927
rect 23716 3896 23949 3924
rect 23716 3884 23722 3896
rect 23937 3893 23949 3896
rect 23983 3924 23995 3927
rect 25314 3924 25320 3936
rect 23983 3896 25320 3924
rect 23983 3893 23995 3896
rect 23937 3887 23995 3893
rect 25314 3884 25320 3896
rect 25372 3884 25378 3936
rect 25682 3884 25688 3936
rect 25740 3924 25746 3936
rect 26237 3927 26295 3933
rect 26237 3924 26249 3927
rect 25740 3896 26249 3924
rect 25740 3884 25746 3896
rect 26237 3893 26249 3896
rect 26283 3893 26295 3927
rect 26237 3887 26295 3893
rect 26786 3884 26792 3936
rect 26844 3924 26850 3936
rect 28442 3924 28448 3936
rect 26844 3896 28448 3924
rect 26844 3884 26850 3896
rect 28442 3884 28448 3896
rect 28500 3884 28506 3936
rect 31726 3924 31754 3964
rect 33336 3924 33364 4032
rect 33594 4020 33600 4032
rect 33652 4060 33658 4072
rect 33965 4063 34023 4069
rect 33965 4060 33977 4063
rect 33652 4032 33977 4060
rect 33652 4020 33658 4032
rect 33965 4029 33977 4032
rect 34011 4060 34023 4063
rect 34422 4060 34428 4072
rect 34011 4032 34428 4060
rect 34011 4029 34023 4032
rect 33965 4023 34023 4029
rect 34422 4020 34428 4032
rect 34480 4020 34486 4072
rect 35452 4060 35480 4091
rect 35710 4088 35716 4100
rect 35768 4088 35774 4140
rect 37458 4088 37464 4140
rect 37516 4128 37522 4140
rect 37553 4131 37611 4137
rect 37553 4128 37565 4131
rect 37516 4100 37565 4128
rect 37516 4088 37522 4100
rect 37553 4097 37565 4100
rect 37599 4097 37611 4131
rect 37553 4091 37611 4097
rect 37645 4131 37703 4137
rect 37645 4097 37657 4131
rect 37691 4097 37703 4131
rect 37645 4091 37703 4097
rect 36814 4060 36820 4072
rect 35452 4032 36820 4060
rect 36814 4020 36820 4032
rect 36872 4020 36878 4072
rect 34054 3952 34060 4004
rect 34112 3992 34118 4004
rect 36357 3995 36415 4001
rect 36357 3992 36369 3995
rect 34112 3964 36369 3992
rect 34112 3952 34118 3964
rect 36357 3961 36369 3964
rect 36403 3961 36415 3995
rect 36357 3955 36415 3961
rect 33502 3924 33508 3936
rect 31726 3896 33364 3924
rect 33463 3896 33508 3924
rect 33502 3884 33508 3896
rect 33560 3884 33566 3936
rect 35894 3924 35900 3936
rect 35855 3896 35900 3924
rect 35894 3884 35900 3896
rect 35952 3884 35958 3936
rect 35986 3884 35992 3936
rect 36044 3924 36050 3936
rect 36170 3924 36176 3936
rect 36044 3896 36176 3924
rect 36044 3884 36050 3896
rect 36170 3884 36176 3896
rect 36228 3924 36234 3936
rect 37660 3924 37688 4091
rect 37734 4088 37740 4140
rect 37792 4128 37798 4140
rect 37918 4137 37924 4140
rect 37792 4100 37837 4128
rect 37792 4088 37798 4100
rect 37915 4091 37924 4137
rect 37976 4128 37982 4140
rect 39022 4128 39028 4140
rect 37976 4100 38015 4128
rect 38983 4100 39028 4128
rect 37918 4088 37924 4091
rect 37976 4088 37982 4100
rect 39022 4088 39028 4100
rect 39080 4088 39086 4140
rect 39298 4128 39304 4140
rect 39211 4100 39304 4128
rect 39298 4088 39304 4100
rect 39356 4128 39362 4140
rect 39850 4128 39856 4140
rect 39356 4100 39856 4128
rect 39356 4088 39362 4100
rect 39850 4088 39856 4100
rect 39908 4088 39914 4140
rect 40310 4128 40316 4140
rect 40271 4100 40316 4128
rect 40310 4088 40316 4100
rect 40368 4088 40374 4140
rect 40494 4088 40500 4140
rect 40552 4128 40558 4140
rect 40589 4131 40647 4137
rect 40589 4128 40601 4131
rect 40552 4100 40601 4128
rect 40552 4088 40558 4100
rect 40589 4097 40601 4100
rect 40635 4128 40647 4131
rect 40678 4128 40684 4140
rect 40635 4100 40684 4128
rect 40635 4097 40647 4100
rect 40589 4091 40647 4097
rect 40678 4088 40684 4100
rect 40736 4088 40742 4140
rect 40862 4088 40868 4140
rect 40920 4128 40926 4140
rect 41049 4131 41107 4137
rect 41049 4128 41061 4131
rect 40920 4100 41061 4128
rect 40920 4088 40926 4100
rect 41049 4097 41061 4100
rect 41095 4097 41107 4131
rect 41049 4091 41107 4097
rect 41141 4131 41199 4137
rect 41141 4097 41153 4131
rect 41187 4097 41199 4131
rect 41322 4128 41328 4140
rect 41283 4100 41328 4128
rect 41141 4091 41199 4097
rect 41156 4060 41184 4091
rect 41322 4088 41328 4100
rect 41380 4088 41386 4140
rect 42794 4088 42800 4140
rect 42852 4128 42858 4140
rect 42996 4137 43024 4168
rect 42981 4131 43039 4137
rect 42981 4128 42993 4131
rect 42852 4100 42993 4128
rect 42852 4088 42858 4100
rect 42981 4097 42993 4100
rect 43027 4097 43039 4131
rect 43162 4128 43168 4140
rect 43123 4100 43168 4128
rect 42981 4091 43039 4097
rect 43162 4088 43168 4100
rect 43220 4088 43226 4140
rect 43257 4131 43315 4137
rect 43257 4097 43269 4131
rect 43303 4097 43315 4131
rect 43257 4091 43315 4097
rect 43349 4131 43407 4137
rect 43349 4097 43361 4131
rect 43395 4128 43407 4131
rect 43530 4128 43536 4140
rect 43395 4100 43536 4128
rect 43395 4097 43407 4100
rect 43349 4091 43407 4097
rect 42886 4060 42892 4072
rect 41064 4032 41184 4060
rect 41386 4032 42892 4060
rect 41064 4004 41092 4032
rect 41046 3952 41052 4004
rect 41104 3952 41110 4004
rect 41386 3924 41414 4032
rect 42886 4020 42892 4032
rect 42944 4060 42950 4072
rect 43272 4060 43300 4091
rect 43530 4088 43536 4100
rect 43588 4128 43594 4140
rect 43990 4128 43996 4140
rect 43588 4100 43996 4128
rect 43588 4088 43594 4100
rect 43990 4088 43996 4100
rect 44048 4088 44054 4140
rect 44100 4137 44128 4168
rect 44284 4168 45376 4196
rect 44284 4137 44312 4168
rect 45370 4156 45376 4168
rect 45428 4156 45434 4208
rect 52012 4196 52040 4224
rect 55490 4196 55496 4208
rect 51736 4168 52040 4196
rect 55232 4168 55496 4196
rect 44085 4131 44143 4137
rect 44085 4097 44097 4131
rect 44131 4097 44143 4131
rect 44085 4091 44143 4097
rect 44269 4131 44327 4137
rect 44269 4097 44281 4131
rect 44315 4097 44327 4131
rect 44269 4091 44327 4097
rect 44361 4131 44419 4137
rect 44361 4097 44373 4131
rect 44407 4097 44419 4131
rect 44361 4091 44419 4097
rect 43622 4060 43628 4072
rect 42944 4032 43300 4060
rect 43583 4032 43628 4060
rect 42944 4020 42950 4032
rect 43272 3992 43300 4032
rect 43622 4020 43628 4032
rect 43680 4020 43686 4072
rect 44376 3992 44404 4091
rect 44450 4088 44456 4140
rect 44508 4128 44514 4140
rect 49430 4131 49488 4137
rect 49430 4128 49442 4131
rect 44508 4100 44553 4128
rect 44744 4100 49442 4128
rect 44508 4088 44514 4100
rect 44744 4069 44772 4100
rect 49430 4097 49442 4100
rect 49476 4097 49488 4131
rect 49430 4091 49488 4097
rect 49602 4088 49608 4140
rect 49660 4128 49666 4140
rect 49697 4131 49755 4137
rect 49697 4128 49709 4131
rect 49660 4100 49709 4128
rect 49660 4088 49666 4100
rect 49697 4097 49709 4100
rect 49743 4097 49755 4131
rect 49697 4091 49755 4097
rect 51258 4088 51264 4140
rect 51316 4128 51322 4140
rect 51736 4137 51764 4168
rect 51721 4131 51779 4137
rect 51721 4128 51733 4131
rect 51316 4100 51733 4128
rect 51316 4088 51322 4100
rect 51721 4097 51733 4100
rect 51767 4097 51779 4131
rect 51721 4091 51779 4097
rect 51810 4088 51816 4140
rect 51868 4128 51874 4140
rect 51997 4131 52055 4137
rect 51868 4100 51913 4128
rect 51868 4088 51874 4100
rect 51997 4097 52009 4131
rect 52043 4097 52055 4131
rect 52178 4128 52184 4140
rect 52139 4100 52184 4128
rect 51997 4091 52055 4097
rect 44729 4063 44787 4069
rect 44729 4029 44741 4063
rect 44775 4029 44787 4063
rect 45833 4063 45891 4069
rect 45833 4060 45845 4063
rect 44729 4023 44787 4029
rect 44836 4032 45845 4060
rect 43272 3964 44404 3992
rect 41506 3924 41512 3936
rect 36228 3896 41414 3924
rect 41467 3896 41512 3924
rect 36228 3884 36234 3896
rect 41506 3884 41512 3896
rect 41564 3884 41570 3936
rect 42426 3924 42432 3936
rect 42387 3896 42432 3924
rect 42426 3884 42432 3896
rect 42484 3884 42490 3936
rect 43162 3884 43168 3936
rect 43220 3924 43226 3936
rect 44836 3924 44864 4032
rect 45833 4029 45845 4032
rect 45879 4029 45891 4063
rect 52012 4060 52040 4091
rect 52178 4088 52184 4100
rect 52236 4088 52242 4140
rect 54018 4128 54024 4140
rect 53979 4100 54024 4128
rect 54018 4088 54024 4100
rect 54076 4088 54082 4140
rect 54113 4131 54171 4137
rect 54113 4097 54125 4131
rect 54159 4097 54171 4131
rect 54113 4091 54171 4097
rect 54481 4131 54539 4137
rect 54481 4097 54493 4131
rect 54527 4128 54539 4131
rect 55125 4131 55183 4137
rect 55125 4128 55137 4131
rect 54527 4100 55137 4128
rect 54527 4097 54539 4100
rect 54481 4091 54539 4097
rect 55125 4097 55137 4100
rect 55171 4128 55183 4131
rect 55232 4128 55260 4168
rect 55490 4156 55496 4168
rect 55548 4196 55554 4208
rect 55861 4199 55919 4205
rect 55861 4196 55873 4199
rect 55548 4168 55873 4196
rect 55548 4156 55554 4168
rect 55861 4165 55873 4168
rect 55907 4165 55919 4199
rect 55861 4159 55919 4165
rect 55171 4100 55260 4128
rect 55171 4097 55183 4100
rect 55125 4091 55183 4097
rect 54128 4060 54156 4091
rect 55674 4088 55680 4140
rect 55732 4128 55738 4140
rect 55769 4131 55827 4137
rect 55769 4128 55781 4131
rect 55732 4100 55781 4128
rect 55732 4088 55738 4100
rect 55769 4097 55781 4100
rect 55815 4097 55827 4131
rect 55950 4128 55956 4140
rect 55911 4100 55956 4128
rect 55769 4091 55827 4097
rect 55950 4088 55956 4100
rect 56008 4088 56014 4140
rect 57882 4128 57888 4140
rect 57843 4100 57888 4128
rect 57882 4088 57888 4100
rect 57940 4088 57946 4140
rect 55309 4063 55367 4069
rect 55309 4060 55321 4063
rect 52012 4032 53512 4060
rect 54128 4032 55321 4060
rect 45833 4023 45891 4029
rect 53484 4004 53512 4032
rect 55140 4004 55168 4032
rect 55309 4029 55321 4032
rect 55355 4029 55367 4063
rect 55309 4023 55367 4029
rect 45002 3952 45008 4004
rect 45060 3992 45066 4004
rect 46477 3995 46535 4001
rect 46477 3992 46489 3995
rect 45060 3964 46489 3992
rect 45060 3952 45066 3964
rect 46477 3961 46489 3964
rect 46523 3961 46535 3995
rect 46477 3955 46535 3961
rect 49694 3952 49700 4004
rect 49752 3992 49758 4004
rect 50801 3995 50859 4001
rect 50801 3992 50813 3995
rect 49752 3964 50813 3992
rect 49752 3952 49758 3964
rect 50801 3961 50813 3964
rect 50847 3961 50859 3995
rect 50801 3955 50859 3961
rect 51902 3952 51908 4004
rect 51960 3992 51966 4004
rect 53377 3995 53435 4001
rect 53377 3992 53389 3995
rect 51960 3964 53389 3992
rect 51960 3952 51966 3964
rect 53377 3961 53389 3964
rect 53423 3961 53435 3995
rect 53377 3955 53435 3961
rect 53466 3952 53472 4004
rect 53524 3992 53530 4004
rect 54297 3995 54355 4001
rect 54297 3992 54309 3995
rect 53524 3964 54309 3992
rect 53524 3952 53530 3964
rect 54297 3961 54309 3964
rect 54343 3961 54355 3995
rect 54297 3955 54355 3961
rect 55122 3952 55128 4004
rect 55180 3952 55186 4004
rect 55214 3952 55220 4004
rect 55272 3992 55278 4004
rect 57977 3995 58035 4001
rect 57977 3992 57989 3995
rect 55272 3964 57989 3992
rect 55272 3952 55278 3964
rect 57977 3961 57989 3964
rect 58023 3961 58035 3995
rect 57977 3955 58035 3961
rect 43220 3896 44864 3924
rect 43220 3884 43226 3896
rect 44910 3884 44916 3936
rect 44968 3924 44974 3936
rect 45189 3927 45247 3933
rect 45189 3924 45201 3927
rect 44968 3896 45201 3924
rect 44968 3884 44974 3896
rect 45189 3893 45201 3896
rect 45235 3893 45247 3927
rect 45189 3887 45247 3893
rect 45278 3884 45284 3936
rect 45336 3924 45342 3936
rect 47581 3927 47639 3933
rect 47581 3924 47593 3927
rect 45336 3896 47593 3924
rect 45336 3884 45342 3896
rect 47581 3893 47593 3896
rect 47627 3893 47639 3927
rect 47581 3887 47639 3893
rect 47762 3884 47768 3936
rect 47820 3924 47826 3936
rect 50157 3927 50215 3933
rect 50157 3924 50169 3927
rect 47820 3896 50169 3924
rect 47820 3884 47826 3896
rect 50157 3893 50169 3896
rect 50203 3893 50215 3927
rect 50157 3887 50215 3893
rect 51074 3884 51080 3936
rect 51132 3924 51138 3936
rect 52733 3927 52791 3933
rect 52733 3924 52745 3927
rect 51132 3896 52745 3924
rect 51132 3884 51138 3896
rect 52733 3893 52745 3896
rect 52779 3893 52791 3927
rect 52733 3887 52791 3893
rect 54570 3884 54576 3936
rect 54628 3924 54634 3936
rect 54941 3927 54999 3933
rect 54941 3924 54953 3927
rect 54628 3896 54953 3924
rect 54628 3884 54634 3896
rect 54941 3893 54953 3896
rect 54987 3893 54999 3927
rect 56502 3924 56508 3936
rect 56463 3896 56508 3924
rect 54941 3887 54999 3893
rect 56502 3884 56508 3896
rect 56560 3884 56566 3936
rect 57057 3927 57115 3933
rect 57057 3893 57069 3927
rect 57103 3924 57115 3927
rect 57790 3924 57796 3936
rect 57103 3896 57796 3924
rect 57103 3893 57115 3896
rect 57057 3887 57115 3893
rect 57790 3884 57796 3896
rect 57848 3884 57854 3936
rect 1104 3834 58880 3856
rect 1104 3782 8174 3834
rect 8226 3782 8238 3834
rect 8290 3782 8302 3834
rect 8354 3782 8366 3834
rect 8418 3782 8430 3834
rect 8482 3782 22622 3834
rect 22674 3782 22686 3834
rect 22738 3782 22750 3834
rect 22802 3782 22814 3834
rect 22866 3782 22878 3834
rect 22930 3782 37070 3834
rect 37122 3782 37134 3834
rect 37186 3782 37198 3834
rect 37250 3782 37262 3834
rect 37314 3782 37326 3834
rect 37378 3782 51518 3834
rect 51570 3782 51582 3834
rect 51634 3782 51646 3834
rect 51698 3782 51710 3834
rect 51762 3782 51774 3834
rect 51826 3782 58880 3834
rect 1104 3760 58880 3782
rect 2038 3720 2044 3732
rect 1999 3692 2044 3720
rect 2038 3680 2044 3692
rect 2096 3680 2102 3732
rect 2406 3680 2412 3732
rect 2464 3720 2470 3732
rect 2501 3723 2559 3729
rect 2501 3720 2513 3723
rect 2464 3692 2513 3720
rect 2464 3680 2470 3692
rect 2501 3689 2513 3692
rect 2547 3720 2559 3723
rect 3881 3723 3939 3729
rect 3881 3720 3893 3723
rect 2547 3692 3893 3720
rect 2547 3689 2559 3692
rect 2501 3683 2559 3689
rect 3881 3689 3893 3692
rect 3927 3689 3939 3723
rect 3881 3683 3939 3689
rect 4246 3680 4252 3732
rect 4304 3720 4310 3732
rect 4433 3723 4491 3729
rect 4433 3720 4445 3723
rect 4304 3692 4445 3720
rect 4304 3680 4310 3692
rect 4433 3689 4445 3692
rect 4479 3689 4491 3723
rect 4433 3683 4491 3689
rect 4798 3680 4804 3732
rect 4856 3720 4862 3732
rect 7006 3720 7012 3732
rect 4856 3692 7012 3720
rect 4856 3680 4862 3692
rect 7006 3680 7012 3692
rect 7064 3680 7070 3732
rect 7466 3680 7472 3732
rect 7524 3720 7530 3732
rect 7561 3723 7619 3729
rect 7561 3720 7573 3723
rect 7524 3692 7573 3720
rect 7524 3680 7530 3692
rect 7561 3689 7573 3692
rect 7607 3689 7619 3723
rect 7561 3683 7619 3689
rect 7742 3680 7748 3732
rect 7800 3720 7806 3732
rect 10042 3720 10048 3732
rect 7800 3692 10048 3720
rect 7800 3680 7806 3692
rect 10042 3680 10048 3692
rect 10100 3680 10106 3732
rect 13538 3720 13544 3732
rect 11348 3692 13400 3720
rect 13499 3692 13544 3720
rect 1394 3612 1400 3664
rect 1452 3652 1458 3664
rect 1949 3655 2007 3661
rect 1949 3652 1961 3655
rect 1452 3624 1961 3652
rect 1452 3612 1458 3624
rect 1949 3621 1961 3624
rect 1995 3652 2007 3655
rect 1995 3624 2636 3652
rect 1995 3621 2007 3624
rect 1949 3615 2007 3621
rect 1765 3587 1823 3593
rect 1765 3553 1777 3587
rect 1811 3584 1823 3587
rect 2406 3584 2412 3596
rect 1811 3556 2412 3584
rect 1811 3553 1823 3556
rect 1765 3547 1823 3553
rect 2406 3544 2412 3556
rect 2464 3544 2470 3596
rect 2608 3593 2636 3624
rect 2774 3612 2780 3664
rect 2832 3612 2838 3664
rect 2958 3652 2964 3664
rect 2919 3624 2964 3652
rect 2958 3612 2964 3624
rect 3016 3612 3022 3664
rect 6546 3612 6552 3664
rect 6604 3652 6610 3664
rect 6641 3655 6699 3661
rect 6641 3652 6653 3655
rect 6604 3624 6653 3652
rect 6604 3612 6610 3624
rect 6641 3621 6653 3624
rect 6687 3621 6699 3655
rect 6641 3615 6699 3621
rect 7374 3612 7380 3664
rect 7432 3652 7438 3664
rect 8478 3652 8484 3664
rect 7432 3624 8484 3652
rect 7432 3612 7438 3624
rect 8478 3612 8484 3624
rect 8536 3612 8542 3664
rect 10502 3612 10508 3664
rect 10560 3652 10566 3664
rect 10870 3652 10876 3664
rect 10560 3624 10876 3652
rect 10560 3612 10566 3624
rect 10870 3612 10876 3624
rect 10928 3612 10934 3664
rect 2593 3587 2651 3593
rect 2593 3553 2605 3587
rect 2639 3553 2651 3587
rect 2792 3584 2820 3612
rect 4706 3584 4712 3596
rect 2792 3556 4712 3584
rect 2593 3547 2651 3553
rect 4706 3544 4712 3556
rect 4764 3544 4770 3596
rect 5258 3584 5264 3596
rect 5219 3556 5264 3584
rect 5258 3544 5264 3556
rect 5316 3544 5322 3596
rect 7098 3544 7104 3596
rect 7156 3584 7162 3596
rect 7742 3584 7748 3596
rect 7156 3556 7748 3584
rect 7156 3544 7162 3556
rect 7742 3544 7748 3556
rect 7800 3544 7806 3596
rect 8110 3584 8116 3596
rect 7852 3556 8116 3584
rect 2041 3519 2099 3525
rect 2041 3485 2053 3519
rect 2087 3516 2099 3519
rect 2777 3519 2835 3525
rect 2087 3488 2544 3516
rect 2087 3485 2099 3488
rect 2041 3479 2099 3485
rect 2516 3457 2544 3488
rect 2777 3485 2789 3519
rect 2823 3516 2835 3519
rect 2866 3516 2872 3528
rect 2823 3488 2872 3516
rect 2823 3485 2835 3488
rect 2777 3479 2835 3485
rect 2866 3476 2872 3488
rect 2924 3476 2930 3528
rect 4157 3519 4215 3525
rect 4157 3485 4169 3519
rect 4203 3485 4215 3519
rect 4157 3479 4215 3485
rect 2501 3451 2559 3457
rect 2501 3417 2513 3451
rect 2547 3417 2559 3451
rect 3786 3448 3792 3460
rect 3747 3420 3792 3448
rect 2501 3411 2559 3417
rect 2516 3380 2544 3411
rect 3786 3408 3792 3420
rect 3844 3408 3850 3460
rect 4172 3448 4200 3479
rect 4246 3476 4252 3528
rect 4304 3516 4310 3528
rect 5534 3525 5540 3528
rect 5528 3516 5540 3525
rect 4304 3488 4349 3516
rect 5495 3488 5540 3516
rect 4304 3476 4310 3488
rect 5528 3479 5540 3488
rect 5534 3476 5540 3479
rect 5592 3476 5598 3528
rect 6914 3476 6920 3528
rect 6972 3516 6978 3528
rect 7374 3516 7380 3528
rect 6972 3488 7380 3516
rect 6972 3476 6978 3488
rect 7374 3476 7380 3488
rect 7432 3476 7438 3528
rect 7653 3519 7711 3525
rect 7653 3485 7665 3519
rect 7699 3516 7711 3519
rect 7852 3516 7880 3556
rect 8110 3544 8116 3556
rect 8168 3584 8174 3596
rect 8570 3584 8576 3596
rect 8168 3556 8576 3584
rect 8168 3544 8174 3556
rect 8570 3544 8576 3556
rect 8628 3544 8634 3596
rect 8846 3544 8852 3596
rect 8904 3584 8910 3596
rect 9033 3587 9091 3593
rect 9033 3584 9045 3587
rect 8904 3556 9045 3584
rect 8904 3544 8910 3556
rect 9033 3553 9045 3556
rect 9079 3553 9091 3587
rect 9033 3547 9091 3553
rect 9858 3544 9864 3596
rect 9916 3584 9922 3596
rect 10778 3584 10784 3596
rect 9916 3556 10784 3584
rect 9916 3544 9922 3556
rect 10778 3544 10784 3556
rect 10836 3544 10842 3596
rect 10965 3587 11023 3593
rect 10965 3553 10977 3587
rect 11011 3584 11023 3587
rect 11348 3584 11376 3692
rect 13372 3652 13400 3692
rect 13538 3680 13544 3692
rect 13596 3680 13602 3732
rect 15378 3720 15384 3732
rect 13648 3692 15384 3720
rect 13648 3652 13676 3692
rect 15378 3680 15384 3692
rect 15436 3680 15442 3732
rect 15838 3680 15844 3732
rect 15896 3720 15902 3732
rect 16761 3723 16819 3729
rect 16761 3720 16773 3723
rect 15896 3692 16773 3720
rect 15896 3680 15902 3692
rect 16761 3689 16773 3692
rect 16807 3689 16819 3723
rect 17034 3720 17040 3732
rect 16761 3683 16819 3689
rect 16868 3692 17040 3720
rect 13372 3624 13676 3652
rect 14090 3612 14096 3664
rect 14148 3652 14154 3664
rect 16868 3652 16896 3692
rect 17034 3680 17040 3692
rect 17092 3720 17098 3732
rect 22370 3720 22376 3732
rect 17092 3692 22376 3720
rect 17092 3680 17098 3692
rect 22370 3680 22376 3692
rect 22428 3680 22434 3732
rect 22462 3680 22468 3732
rect 22520 3720 22526 3732
rect 23753 3723 23811 3729
rect 23753 3720 23765 3723
rect 22520 3692 23765 3720
rect 22520 3680 22526 3692
rect 23753 3689 23765 3692
rect 23799 3689 23811 3723
rect 23753 3683 23811 3689
rect 23842 3680 23848 3732
rect 23900 3720 23906 3732
rect 25130 3720 25136 3732
rect 23900 3692 25136 3720
rect 23900 3680 23906 3692
rect 25130 3680 25136 3692
rect 25188 3680 25194 3732
rect 26050 3680 26056 3732
rect 26108 3720 26114 3732
rect 26789 3723 26847 3729
rect 26789 3720 26801 3723
rect 26108 3692 26801 3720
rect 26108 3680 26114 3692
rect 26789 3689 26801 3692
rect 26835 3720 26847 3723
rect 26878 3720 26884 3732
rect 26835 3692 26884 3720
rect 26835 3689 26847 3692
rect 26789 3683 26847 3689
rect 26878 3680 26884 3692
rect 26936 3680 26942 3732
rect 27062 3680 27068 3732
rect 27120 3720 27126 3732
rect 31202 3720 31208 3732
rect 27120 3692 31208 3720
rect 27120 3680 27126 3692
rect 31202 3680 31208 3692
rect 31260 3680 31266 3732
rect 32674 3720 32680 3732
rect 32635 3692 32680 3720
rect 32674 3680 32680 3692
rect 32732 3680 32738 3732
rect 33318 3680 33324 3732
rect 33376 3720 33382 3732
rect 33413 3723 33471 3729
rect 33413 3720 33425 3723
rect 33376 3692 33425 3720
rect 33376 3680 33382 3692
rect 33413 3689 33425 3692
rect 33459 3689 33471 3723
rect 34790 3720 34796 3732
rect 34751 3692 34796 3720
rect 33413 3683 33471 3689
rect 34790 3680 34796 3692
rect 34848 3680 34854 3732
rect 35250 3680 35256 3732
rect 35308 3720 35314 3732
rect 35308 3692 36492 3720
rect 35308 3680 35314 3692
rect 14148 3624 16896 3652
rect 14148 3612 14154 3624
rect 11514 3584 11520 3596
rect 11011 3556 11376 3584
rect 11475 3556 11520 3584
rect 11011 3553 11023 3556
rect 10965 3547 11023 3553
rect 11514 3544 11520 3556
rect 11572 3544 11578 3596
rect 7699 3488 7880 3516
rect 7929 3519 7987 3525
rect 7699 3485 7711 3488
rect 7653 3479 7711 3485
rect 7929 3485 7941 3519
rect 7975 3485 7987 3519
rect 7929 3479 7987 3485
rect 7282 3448 7288 3460
rect 4172 3420 7288 3448
rect 7282 3408 7288 3420
rect 7340 3448 7346 3460
rect 7340 3420 7420 3448
rect 7340 3408 7346 3420
rect 5442 3380 5448 3392
rect 2516 3352 5448 3380
rect 5442 3340 5448 3352
rect 5500 3340 5506 3392
rect 7392 3389 7420 3420
rect 7466 3408 7472 3460
rect 7524 3448 7530 3460
rect 7944 3448 7972 3479
rect 8754 3476 8760 3528
rect 8812 3516 8818 3528
rect 9309 3519 9367 3525
rect 9309 3516 9321 3519
rect 8812 3488 9321 3516
rect 8812 3476 8818 3488
rect 9309 3485 9321 3488
rect 9355 3516 9367 3519
rect 9490 3516 9496 3528
rect 9355 3488 9496 3516
rect 9355 3485 9367 3488
rect 9309 3479 9367 3485
rect 9490 3476 9496 3488
rect 9548 3476 9554 3528
rect 10413 3519 10471 3525
rect 10413 3485 10425 3519
rect 10459 3516 10471 3519
rect 10502 3516 10508 3528
rect 10459 3488 10508 3516
rect 10459 3485 10471 3488
rect 10413 3479 10471 3485
rect 10502 3476 10508 3488
rect 10560 3476 10566 3528
rect 10597 3519 10655 3525
rect 10597 3485 10609 3519
rect 10643 3485 10655 3519
rect 10597 3479 10655 3485
rect 10612 3448 10640 3479
rect 12526 3476 12532 3528
rect 12584 3516 12590 3528
rect 13357 3519 13415 3525
rect 13357 3516 13369 3519
rect 12584 3488 13369 3516
rect 12584 3476 12590 3488
rect 13357 3485 13369 3488
rect 13403 3485 13415 3519
rect 13357 3479 13415 3485
rect 13541 3519 13599 3525
rect 13541 3485 13553 3519
rect 13587 3516 13599 3519
rect 13722 3516 13728 3528
rect 13587 3488 13728 3516
rect 13587 3485 13599 3488
rect 13541 3479 13599 3485
rect 13722 3476 13728 3488
rect 13780 3476 13786 3528
rect 14366 3476 14372 3528
rect 14424 3516 14430 3528
rect 14568 3525 14596 3624
rect 17402 3612 17408 3664
rect 17460 3652 17466 3664
rect 18414 3652 18420 3664
rect 17460 3624 18420 3652
rect 17460 3612 17466 3624
rect 18414 3612 18420 3624
rect 18472 3612 18478 3664
rect 21082 3612 21088 3664
rect 21140 3652 21146 3664
rect 25314 3652 25320 3664
rect 21140 3624 25320 3652
rect 21140 3612 21146 3624
rect 25314 3612 25320 3624
rect 25372 3612 25378 3664
rect 28258 3652 28264 3664
rect 27356 3624 28264 3652
rect 16853 3587 16911 3593
rect 16853 3584 16865 3587
rect 16040 3556 16865 3584
rect 14461 3519 14519 3525
rect 14461 3516 14473 3519
rect 14424 3488 14473 3516
rect 14424 3476 14430 3488
rect 14461 3485 14473 3488
rect 14507 3485 14519 3519
rect 14461 3479 14519 3485
rect 14553 3519 14611 3525
rect 14553 3485 14565 3519
rect 14599 3485 14611 3519
rect 14553 3479 14611 3485
rect 14645 3519 14703 3525
rect 14645 3485 14657 3519
rect 14691 3485 14703 3519
rect 14826 3516 14832 3528
rect 14787 3488 14832 3516
rect 14645 3479 14703 3485
rect 7524 3420 10640 3448
rect 11784 3451 11842 3457
rect 7524 3408 7530 3420
rect 11784 3417 11796 3451
rect 11830 3448 11842 3451
rect 14185 3451 14243 3457
rect 14185 3448 14197 3451
rect 11830 3420 14197 3448
rect 11830 3417 11842 3420
rect 11784 3411 11842 3417
rect 14185 3417 14197 3420
rect 14231 3417 14243 3451
rect 14660 3448 14688 3479
rect 14826 3476 14832 3488
rect 14884 3476 14890 3528
rect 15286 3476 15292 3528
rect 15344 3516 15350 3528
rect 15746 3516 15752 3528
rect 15344 3488 15752 3516
rect 15344 3476 15350 3488
rect 15746 3476 15752 3488
rect 15804 3476 15810 3528
rect 16040 3525 16068 3556
rect 16853 3553 16865 3556
rect 16899 3553 16911 3587
rect 19886 3584 19892 3596
rect 16853 3547 16911 3553
rect 17052 3556 19892 3584
rect 16025 3519 16083 3525
rect 16025 3485 16037 3519
rect 16071 3485 16083 3519
rect 16298 3516 16304 3528
rect 16211 3488 16304 3516
rect 16025 3479 16083 3485
rect 15841 3451 15899 3457
rect 15841 3448 15853 3451
rect 14660 3420 15853 3448
rect 14185 3411 14243 3417
rect 15841 3417 15853 3420
rect 15887 3417 15899 3451
rect 15841 3411 15899 3417
rect 7377 3383 7435 3389
rect 7377 3349 7389 3383
rect 7423 3349 7435 3383
rect 7377 3343 7435 3349
rect 8202 3340 8208 3392
rect 8260 3380 8266 3392
rect 9674 3380 9680 3392
rect 8260 3352 9680 3380
rect 8260 3340 8266 3352
rect 9674 3340 9680 3352
rect 9732 3340 9738 3392
rect 9950 3340 9956 3392
rect 10008 3380 10014 3392
rect 10686 3380 10692 3392
rect 10008 3352 10692 3380
rect 10008 3340 10014 3352
rect 10686 3340 10692 3352
rect 10744 3340 10750 3392
rect 10870 3340 10876 3392
rect 10928 3380 10934 3392
rect 12710 3380 12716 3392
rect 10928 3352 12716 3380
rect 10928 3340 10934 3352
rect 12710 3340 12716 3352
rect 12768 3340 12774 3392
rect 12897 3383 12955 3389
rect 12897 3349 12909 3383
rect 12943 3380 12955 3383
rect 16040 3380 16068 3479
rect 16298 3476 16304 3488
rect 16356 3476 16362 3528
rect 16574 3476 16580 3528
rect 16632 3516 16638 3528
rect 17052 3525 17080 3556
rect 19886 3544 19892 3556
rect 19944 3544 19950 3596
rect 21358 3584 21364 3596
rect 20732 3556 21364 3584
rect 16761 3519 16819 3525
rect 16761 3516 16773 3519
rect 16632 3488 16773 3516
rect 16632 3476 16638 3488
rect 16761 3485 16773 3488
rect 16807 3485 16819 3519
rect 16761 3479 16819 3485
rect 17037 3519 17095 3525
rect 17037 3485 17049 3519
rect 17083 3485 17095 3519
rect 17954 3516 17960 3528
rect 17915 3488 17960 3516
rect 17037 3479 17095 3485
rect 17954 3476 17960 3488
rect 18012 3476 18018 3528
rect 18322 3476 18328 3528
rect 18380 3516 18386 3528
rect 18417 3519 18475 3525
rect 18417 3516 18429 3519
rect 18380 3488 18429 3516
rect 18380 3476 18386 3488
rect 18417 3485 18429 3488
rect 18463 3485 18475 3519
rect 19242 3516 19248 3528
rect 19203 3488 19248 3516
rect 18417 3479 18475 3485
rect 19242 3476 19248 3488
rect 19300 3476 19306 3528
rect 19521 3519 19579 3525
rect 19521 3485 19533 3519
rect 19567 3516 19579 3519
rect 20732 3516 20760 3556
rect 21358 3544 21364 3556
rect 21416 3544 21422 3596
rect 25409 3587 25467 3593
rect 25409 3584 25421 3587
rect 22756 3556 25421 3584
rect 19567 3488 20760 3516
rect 20809 3519 20867 3525
rect 19567 3485 19579 3488
rect 19521 3479 19579 3485
rect 20809 3485 20821 3519
rect 20855 3516 20867 3519
rect 22094 3516 22100 3528
rect 20855 3488 22100 3516
rect 20855 3485 20867 3488
rect 20809 3479 20867 3485
rect 16316 3448 16344 3476
rect 17310 3448 17316 3460
rect 16316 3420 17316 3448
rect 17310 3408 17316 3420
rect 17368 3448 17374 3460
rect 19536 3448 19564 3479
rect 22094 3476 22100 3488
rect 22152 3476 22158 3528
rect 22756 3448 22784 3556
rect 25409 3553 25421 3556
rect 25455 3553 25467 3587
rect 25409 3547 25467 3553
rect 23293 3519 23351 3525
rect 23293 3485 23305 3519
rect 23339 3516 23351 3519
rect 23382 3516 23388 3528
rect 23339 3488 23388 3516
rect 23339 3485 23351 3488
rect 23293 3479 23351 3485
rect 23382 3476 23388 3488
rect 23440 3476 23446 3528
rect 24949 3519 25007 3525
rect 24949 3485 24961 3519
rect 24995 3516 25007 3519
rect 27356 3516 27384 3624
rect 28258 3612 28264 3624
rect 28316 3612 28322 3664
rect 30834 3612 30840 3664
rect 30892 3652 30898 3664
rect 34606 3652 34612 3664
rect 30892 3624 34612 3652
rect 30892 3612 30898 3624
rect 34606 3612 34612 3624
rect 34664 3612 34670 3664
rect 36464 3652 36492 3692
rect 37550 3680 37556 3732
rect 37608 3720 37614 3732
rect 38654 3720 38660 3732
rect 37608 3692 38660 3720
rect 37608 3680 37614 3692
rect 38654 3680 38660 3692
rect 38712 3680 38718 3732
rect 40497 3723 40555 3729
rect 40497 3689 40509 3723
rect 40543 3689 40555 3723
rect 40497 3683 40555 3689
rect 39482 3652 39488 3664
rect 36464 3624 39488 3652
rect 39482 3612 39488 3624
rect 39540 3612 39546 3664
rect 40037 3655 40095 3661
rect 40037 3621 40049 3655
rect 40083 3621 40095 3655
rect 40512 3652 40540 3683
rect 41966 3680 41972 3732
rect 42024 3720 42030 3732
rect 44910 3720 44916 3732
rect 42024 3692 44916 3720
rect 42024 3680 42030 3692
rect 44910 3680 44916 3692
rect 44968 3680 44974 3732
rect 48038 3680 48044 3732
rect 48096 3720 48102 3732
rect 50801 3723 50859 3729
rect 50801 3720 50813 3723
rect 48096 3692 50813 3720
rect 48096 3680 48102 3692
rect 50801 3689 50813 3692
rect 50847 3689 50859 3723
rect 52270 3720 52276 3732
rect 52231 3692 52276 3720
rect 50801 3683 50859 3689
rect 52270 3680 52276 3692
rect 52328 3680 52334 3732
rect 52546 3680 52552 3732
rect 52604 3720 52610 3732
rect 55953 3723 56011 3729
rect 55953 3720 55965 3723
rect 52604 3692 55965 3720
rect 52604 3680 52610 3692
rect 55953 3689 55965 3692
rect 55999 3689 56011 3723
rect 55953 3683 56011 3689
rect 56502 3680 56508 3732
rect 56560 3720 56566 3732
rect 57241 3723 57299 3729
rect 57241 3720 57253 3723
rect 56560 3692 57253 3720
rect 56560 3680 56566 3692
rect 57241 3689 57253 3692
rect 57287 3689 57299 3723
rect 57790 3720 57796 3732
rect 57751 3692 57796 3720
rect 57241 3683 57299 3689
rect 57790 3680 57796 3692
rect 57848 3680 57854 3732
rect 41322 3652 41328 3664
rect 40512 3624 41328 3652
rect 40037 3615 40095 3621
rect 27890 3544 27896 3596
rect 27948 3584 27954 3596
rect 27948 3556 31248 3584
rect 27948 3544 27954 3556
rect 24995 3488 27384 3516
rect 27433 3519 27491 3525
rect 24995 3485 25007 3488
rect 24949 3479 25007 3485
rect 27433 3485 27445 3519
rect 27479 3516 27491 3519
rect 27614 3516 27620 3528
rect 27479 3488 27620 3516
rect 27479 3485 27491 3488
rect 27433 3479 27491 3485
rect 27614 3476 27620 3488
rect 27672 3476 27678 3528
rect 27706 3476 27712 3528
rect 27764 3516 27770 3528
rect 29546 3516 29552 3528
rect 27764 3488 29552 3516
rect 27764 3476 27770 3488
rect 29546 3476 29552 3488
rect 29604 3476 29610 3528
rect 31220 3525 31248 3556
rect 37642 3544 37648 3596
rect 37700 3584 37706 3596
rect 39942 3584 39948 3596
rect 37700 3556 39948 3584
rect 37700 3544 37706 3556
rect 39942 3544 39948 3556
rect 40000 3544 40006 3596
rect 31205 3519 31263 3525
rect 31205 3485 31217 3519
rect 31251 3516 31263 3519
rect 32490 3516 32496 3528
rect 31251 3488 32496 3516
rect 31251 3485 31263 3488
rect 31205 3479 31263 3485
rect 32490 3476 32496 3488
rect 32548 3476 32554 3528
rect 33134 3476 33140 3528
rect 33192 3516 33198 3528
rect 33965 3519 34023 3525
rect 33965 3516 33977 3519
rect 33192 3488 33977 3516
rect 33192 3476 33198 3488
rect 33965 3485 33977 3488
rect 34011 3485 34023 3519
rect 33965 3479 34023 3485
rect 34422 3476 34428 3528
rect 34480 3516 34486 3528
rect 34701 3519 34759 3525
rect 34701 3516 34713 3519
rect 34480 3488 34713 3516
rect 34480 3476 34486 3488
rect 34701 3485 34713 3488
rect 34747 3485 34759 3519
rect 34882 3516 34888 3528
rect 34843 3488 34888 3516
rect 34701 3479 34759 3485
rect 34882 3476 34888 3488
rect 34940 3476 34946 3528
rect 35526 3516 35532 3528
rect 35439 3488 35532 3516
rect 35526 3476 35532 3488
rect 35584 3516 35590 3528
rect 36722 3516 36728 3528
rect 35584 3488 36728 3516
rect 35584 3476 35590 3488
rect 36722 3476 36728 3488
rect 36780 3476 36786 3528
rect 37461 3519 37519 3525
rect 37461 3516 37473 3519
rect 36832 3488 37473 3516
rect 17368 3420 19564 3448
rect 22112 3420 22784 3448
rect 17368 3408 17374 3420
rect 12943 3352 16068 3380
rect 16209 3383 16267 3389
rect 12943 3349 12955 3352
rect 12897 3343 12955 3349
rect 16209 3349 16221 3383
rect 16255 3380 16267 3383
rect 16390 3380 16396 3392
rect 16255 3352 16396 3380
rect 16255 3349 16267 3352
rect 16209 3343 16267 3349
rect 16390 3340 16396 3352
rect 16448 3380 16454 3392
rect 16942 3380 16948 3392
rect 16448 3352 16948 3380
rect 16448 3340 16454 3352
rect 16942 3340 16948 3352
rect 17000 3340 17006 3392
rect 17218 3380 17224 3392
rect 17179 3352 17224 3380
rect 17218 3340 17224 3352
rect 17276 3340 17282 3392
rect 18601 3383 18659 3389
rect 18601 3349 18613 3383
rect 18647 3380 18659 3383
rect 19886 3380 19892 3392
rect 18647 3352 19892 3380
rect 18647 3349 18659 3352
rect 18601 3343 18659 3349
rect 19886 3340 19892 3352
rect 19944 3340 19950 3392
rect 21726 3340 21732 3392
rect 21784 3380 21790 3392
rect 22112 3389 22140 3420
rect 23566 3408 23572 3460
rect 23624 3448 23630 3460
rect 23624 3420 25176 3448
rect 23624 3408 23630 3420
rect 22097 3383 22155 3389
rect 22097 3380 22109 3383
rect 21784 3352 22109 3380
rect 21784 3340 21790 3352
rect 22097 3349 22109 3352
rect 22143 3349 22155 3383
rect 22097 3343 22155 3349
rect 22370 3340 22376 3392
rect 22428 3380 22434 3392
rect 23109 3383 23167 3389
rect 23109 3380 23121 3383
rect 22428 3352 23121 3380
rect 22428 3340 22434 3352
rect 23109 3349 23121 3352
rect 23155 3349 23167 3383
rect 25148 3380 25176 3420
rect 25222 3408 25228 3460
rect 25280 3448 25286 3460
rect 25654 3451 25712 3457
rect 25654 3448 25666 3451
rect 25280 3420 25666 3448
rect 25280 3408 25286 3420
rect 25654 3417 25666 3420
rect 25700 3417 25712 3451
rect 25654 3411 25712 3417
rect 27522 3408 27528 3460
rect 27580 3448 27586 3460
rect 27985 3451 28043 3457
rect 27985 3448 27997 3451
rect 27580 3420 27997 3448
rect 27580 3408 27586 3420
rect 27985 3417 27997 3420
rect 28031 3417 28043 3451
rect 28166 3448 28172 3460
rect 28127 3420 28172 3448
rect 27985 3411 28043 3417
rect 28166 3408 28172 3420
rect 28224 3448 28230 3460
rect 28813 3451 28871 3457
rect 28813 3448 28825 3451
rect 28224 3420 28825 3448
rect 28224 3408 28230 3420
rect 28813 3417 28825 3420
rect 28859 3417 28871 3451
rect 28813 3411 28871 3417
rect 28997 3451 29055 3457
rect 28997 3417 29009 3451
rect 29043 3448 29055 3451
rect 31294 3448 31300 3460
rect 29043 3420 31300 3448
rect 29043 3417 29055 3420
rect 28997 3411 29055 3417
rect 31294 3408 31300 3420
rect 31352 3448 31358 3460
rect 32858 3448 32864 3460
rect 31352 3420 32864 3448
rect 31352 3408 31358 3420
rect 32858 3408 32864 3420
rect 32916 3408 32922 3460
rect 35796 3451 35854 3457
rect 35796 3417 35808 3451
rect 35842 3448 35854 3451
rect 35894 3448 35900 3460
rect 35842 3420 35900 3448
rect 35842 3417 35854 3420
rect 35796 3411 35854 3417
rect 35894 3408 35900 3420
rect 35952 3408 35958 3460
rect 27338 3380 27344 3392
rect 25148 3352 27344 3380
rect 23109 3343 23167 3349
rect 27338 3340 27344 3352
rect 27396 3340 27402 3392
rect 29779 3383 29837 3389
rect 29779 3349 29791 3383
rect 29825 3380 29837 3383
rect 31478 3380 31484 3392
rect 29825 3352 31484 3380
rect 29825 3349 29837 3352
rect 29779 3343 29837 3349
rect 31478 3340 31484 3352
rect 31536 3340 31542 3392
rect 33502 3340 33508 3392
rect 33560 3380 33566 3392
rect 36832 3380 36860 3488
rect 37461 3485 37473 3488
rect 37507 3485 37519 3519
rect 37461 3479 37519 3485
rect 37921 3519 37979 3525
rect 37921 3485 37933 3519
rect 37967 3485 37979 3519
rect 38286 3516 38292 3528
rect 38247 3488 38292 3516
rect 37921 3479 37979 3485
rect 33560 3352 36860 3380
rect 36909 3383 36967 3389
rect 33560 3340 33566 3352
rect 36909 3349 36921 3383
rect 36955 3380 36967 3383
rect 37458 3380 37464 3392
rect 36955 3352 37464 3380
rect 36955 3349 36967 3352
rect 36909 3343 36967 3349
rect 37458 3340 37464 3352
rect 37516 3380 37522 3392
rect 37936 3380 37964 3479
rect 38286 3476 38292 3488
rect 38344 3516 38350 3528
rect 38470 3516 38476 3528
rect 38344 3488 38476 3516
rect 38344 3476 38350 3488
rect 38470 3476 38476 3488
rect 38528 3476 38534 3528
rect 38841 3519 38899 3525
rect 38841 3485 38853 3519
rect 38887 3516 38899 3519
rect 40052 3516 40080 3615
rect 41322 3612 41328 3624
rect 41380 3652 41386 3664
rect 45189 3655 45247 3661
rect 45189 3652 45201 3655
rect 41380 3624 45201 3652
rect 41380 3612 41386 3624
rect 45189 3621 45201 3624
rect 45235 3621 45247 3655
rect 51445 3655 51503 3661
rect 51445 3652 51457 3655
rect 45189 3615 45247 3621
rect 51046 3624 51457 3652
rect 40405 3587 40463 3593
rect 40405 3553 40417 3587
rect 40451 3584 40463 3587
rect 40451 3556 41276 3584
rect 40451 3553 40463 3556
rect 40405 3547 40463 3553
rect 38887 3488 40080 3516
rect 40221 3519 40279 3525
rect 38887 3485 38899 3488
rect 38841 3479 38899 3485
rect 40221 3485 40233 3519
rect 40267 3516 40279 3519
rect 40862 3516 40868 3528
rect 40267 3488 40868 3516
rect 40267 3485 40279 3488
rect 40221 3479 40279 3485
rect 40862 3476 40868 3488
rect 40920 3476 40926 3528
rect 40954 3476 40960 3528
rect 41012 3516 41018 3528
rect 41248 3525 41276 3556
rect 41506 3544 41512 3596
rect 41564 3584 41570 3596
rect 46566 3584 46572 3596
rect 41564 3556 42840 3584
rect 41564 3544 41570 3556
rect 41233 3519 41291 3525
rect 41012 3488 41057 3516
rect 41012 3476 41018 3488
rect 41233 3485 41245 3519
rect 41279 3516 41291 3519
rect 41782 3516 41788 3528
rect 41279 3488 41788 3516
rect 41279 3485 41291 3488
rect 41233 3479 41291 3485
rect 41782 3476 41788 3488
rect 41840 3476 41846 3528
rect 41877 3519 41935 3525
rect 41877 3485 41889 3519
rect 41923 3485 41935 3519
rect 42610 3516 42616 3528
rect 42571 3488 42616 3516
rect 41877 3479 41935 3485
rect 38378 3408 38384 3460
rect 38436 3448 38442 3460
rect 38436 3420 38792 3448
rect 38436 3408 38442 3420
rect 37516 3352 37964 3380
rect 37516 3340 37522 3352
rect 38562 3340 38568 3392
rect 38620 3380 38626 3392
rect 38657 3383 38715 3389
rect 38657 3380 38669 3383
rect 38620 3352 38669 3380
rect 38620 3340 38626 3352
rect 38657 3349 38669 3352
rect 38703 3349 38715 3383
rect 38764 3380 38792 3420
rect 40126 3408 40132 3460
rect 40184 3448 40190 3460
rect 40497 3451 40555 3457
rect 40497 3448 40509 3451
rect 40184 3420 40509 3448
rect 40184 3408 40190 3420
rect 40497 3417 40509 3420
rect 40543 3417 40555 3451
rect 41892 3448 41920 3479
rect 42610 3476 42616 3488
rect 42668 3476 42674 3528
rect 42812 3525 42840 3556
rect 42904 3556 44036 3584
rect 46527 3556 46572 3584
rect 42904 3525 42932 3556
rect 42797 3519 42855 3525
rect 42797 3485 42809 3519
rect 42843 3485 42855 3519
rect 42797 3479 42855 3485
rect 42889 3519 42947 3525
rect 42889 3485 42901 3519
rect 42935 3485 42947 3519
rect 42889 3479 42947 3485
rect 42981 3519 43039 3525
rect 42981 3485 42993 3519
rect 43027 3510 43039 3519
rect 43070 3510 43076 3528
rect 43027 3485 43076 3510
rect 42981 3482 43076 3485
rect 42981 3479 43039 3482
rect 40497 3411 40555 3417
rect 40604 3420 41920 3448
rect 40604 3380 40632 3420
rect 42702 3408 42708 3460
rect 42760 3448 42766 3460
rect 42904 3448 42932 3479
rect 43070 3476 43076 3482
rect 43128 3476 43134 3528
rect 43714 3516 43720 3528
rect 43675 3488 43720 3516
rect 43714 3476 43720 3488
rect 43772 3476 43778 3528
rect 43898 3516 43904 3528
rect 43859 3488 43904 3516
rect 43898 3476 43904 3488
rect 43956 3476 43962 3528
rect 44008 3525 44036 3556
rect 46566 3544 46572 3556
rect 46624 3544 46630 3596
rect 49421 3587 49479 3593
rect 49421 3553 49433 3587
rect 49467 3584 49479 3587
rect 49602 3584 49608 3596
rect 49467 3556 49608 3584
rect 49467 3553 49479 3556
rect 49421 3547 49479 3553
rect 49602 3544 49608 3556
rect 49660 3544 49666 3596
rect 43993 3519 44051 3525
rect 43993 3485 44005 3519
rect 44039 3485 44051 3519
rect 43993 3479 44051 3485
rect 44082 3476 44088 3528
rect 44140 3516 44146 3528
rect 44140 3488 44185 3516
rect 44140 3476 44146 3488
rect 44634 3476 44640 3528
rect 44692 3516 44698 3528
rect 47029 3519 47087 3525
rect 47029 3516 47041 3519
rect 44692 3488 47041 3516
rect 44692 3476 44698 3488
rect 47029 3485 47041 3488
rect 47075 3485 47087 3519
rect 50157 3519 50215 3525
rect 50157 3516 50169 3519
rect 47029 3479 47087 3485
rect 47136 3488 50169 3516
rect 42760 3420 42932 3448
rect 43257 3451 43315 3457
rect 42760 3408 42766 3420
rect 43257 3417 43269 3451
rect 43303 3448 43315 3451
rect 46302 3451 46360 3457
rect 46302 3448 46314 3451
rect 43303 3420 46314 3448
rect 43303 3417 43315 3420
rect 43257 3411 43315 3417
rect 46302 3417 46314 3420
rect 46348 3417 46360 3451
rect 46302 3411 46360 3417
rect 46474 3408 46480 3460
rect 46532 3448 46538 3460
rect 47136 3448 47164 3488
rect 50157 3485 50169 3488
rect 50203 3485 50215 3519
rect 50157 3479 50215 3485
rect 46532 3420 47164 3448
rect 46532 3408 46538 3420
rect 47210 3408 47216 3460
rect 47268 3448 47274 3460
rect 47268 3420 48176 3448
rect 47268 3408 47274 3420
rect 41046 3380 41052 3392
rect 38764 3352 40632 3380
rect 41007 3352 41052 3380
rect 38657 3343 38715 3349
rect 41046 3340 41052 3352
rect 41104 3340 41110 3392
rect 41417 3383 41475 3389
rect 41417 3349 41429 3383
rect 41463 3380 41475 3383
rect 42886 3380 42892 3392
rect 41463 3352 42892 3380
rect 41463 3349 41475 3352
rect 41417 3343 41475 3349
rect 42886 3340 42892 3352
rect 42944 3340 42950 3392
rect 44361 3383 44419 3389
rect 44361 3349 44373 3383
rect 44407 3380 44419 3383
rect 45094 3380 45100 3392
rect 44407 3352 45100 3380
rect 44407 3349 44419 3352
rect 44361 3343 44419 3349
rect 45094 3340 45100 3352
rect 45152 3340 45158 3392
rect 45646 3340 45652 3392
rect 45704 3380 45710 3392
rect 48041 3383 48099 3389
rect 48041 3380 48053 3383
rect 45704 3352 48053 3380
rect 45704 3340 45710 3352
rect 48041 3349 48053 3352
rect 48087 3349 48099 3383
rect 48148 3380 48176 3420
rect 48314 3408 48320 3460
rect 48372 3448 48378 3460
rect 49154 3451 49212 3457
rect 49154 3448 49166 3451
rect 48372 3420 49166 3448
rect 48372 3408 48378 3420
rect 49154 3417 49166 3420
rect 49200 3417 49212 3451
rect 49154 3411 49212 3417
rect 51046 3380 51074 3624
rect 51445 3621 51457 3624
rect 51491 3621 51503 3655
rect 51445 3615 51503 3621
rect 54018 3612 54024 3664
rect 54076 3652 54082 3664
rect 55398 3652 55404 3664
rect 54076 3624 55404 3652
rect 54076 3612 54082 3624
rect 55398 3612 55404 3624
rect 55456 3612 55462 3664
rect 53282 3544 53288 3596
rect 53340 3584 53346 3596
rect 56597 3587 56655 3593
rect 56597 3584 56609 3587
rect 53340 3556 53385 3584
rect 53484 3556 56609 3584
rect 53340 3544 53346 3556
rect 52822 3476 52828 3528
rect 52880 3516 52886 3528
rect 53009 3519 53067 3525
rect 53009 3516 53021 3519
rect 52880 3488 53021 3516
rect 52880 3476 52886 3488
rect 53009 3485 53021 3488
rect 53055 3485 53067 3519
rect 53009 3479 53067 3485
rect 53098 3476 53104 3528
rect 53156 3516 53162 3528
rect 53484 3516 53512 3556
rect 56597 3553 56609 3556
rect 56643 3553 56655 3587
rect 56597 3547 56655 3553
rect 53156 3488 53512 3516
rect 53745 3519 53803 3525
rect 53156 3476 53162 3488
rect 53745 3485 53757 3519
rect 53791 3485 53803 3519
rect 53745 3479 53803 3485
rect 51350 3408 51356 3460
rect 51408 3448 51414 3460
rect 53760 3448 53788 3479
rect 53926 3476 53932 3528
rect 53984 3516 53990 3528
rect 54386 3516 54392 3528
rect 53984 3488 54392 3516
rect 53984 3476 53990 3488
rect 54386 3476 54392 3488
rect 54444 3476 54450 3528
rect 54570 3516 54576 3528
rect 54531 3488 54576 3516
rect 54570 3476 54576 3488
rect 54628 3476 54634 3528
rect 55309 3519 55367 3525
rect 55309 3485 55321 3519
rect 55355 3485 55367 3519
rect 55309 3479 55367 3485
rect 55324 3448 55352 3479
rect 51408 3420 53788 3448
rect 53852 3420 55352 3448
rect 51408 3408 51414 3420
rect 48148 3352 51074 3380
rect 48041 3343 48099 3349
rect 52362 3340 52368 3392
rect 52420 3380 52426 3392
rect 53852 3380 53880 3420
rect 52420 3352 53880 3380
rect 52420 3340 52426 3352
rect 1104 3290 58880 3312
rect 1104 3238 15398 3290
rect 15450 3238 15462 3290
rect 15514 3238 15526 3290
rect 15578 3238 15590 3290
rect 15642 3238 15654 3290
rect 15706 3238 29846 3290
rect 29898 3238 29910 3290
rect 29962 3238 29974 3290
rect 30026 3238 30038 3290
rect 30090 3238 30102 3290
rect 30154 3238 44294 3290
rect 44346 3238 44358 3290
rect 44410 3238 44422 3290
rect 44474 3238 44486 3290
rect 44538 3238 44550 3290
rect 44602 3238 58880 3290
rect 1104 3216 58880 3238
rect 1489 3179 1547 3185
rect 1489 3145 1501 3179
rect 1535 3176 1547 3179
rect 1762 3176 1768 3188
rect 1535 3148 1768 3176
rect 1535 3145 1547 3148
rect 1489 3139 1547 3145
rect 1762 3136 1768 3148
rect 1820 3136 1826 3188
rect 3053 3179 3111 3185
rect 3053 3145 3065 3179
rect 3099 3176 3111 3179
rect 3786 3176 3792 3188
rect 3099 3148 3792 3176
rect 3099 3145 3111 3148
rect 3053 3139 3111 3145
rect 3786 3136 3792 3148
rect 3844 3176 3850 3188
rect 3973 3179 4031 3185
rect 3973 3176 3985 3179
rect 3844 3148 3985 3176
rect 3844 3136 3850 3148
rect 3973 3145 3985 3148
rect 4019 3176 4031 3179
rect 5810 3176 5816 3188
rect 4019 3148 5816 3176
rect 4019 3145 4031 3148
rect 3973 3139 4031 3145
rect 5810 3136 5816 3148
rect 5868 3136 5874 3188
rect 6454 3176 6460 3188
rect 6415 3148 6460 3176
rect 6454 3136 6460 3148
rect 6512 3136 6518 3188
rect 7098 3176 7104 3188
rect 7011 3148 7104 3176
rect 7098 3136 7104 3148
rect 7156 3176 7162 3188
rect 7466 3176 7472 3188
rect 7156 3148 7472 3176
rect 7156 3136 7162 3148
rect 7466 3136 7472 3148
rect 7524 3136 7530 3188
rect 9490 3176 9496 3188
rect 7760 3148 9496 3176
rect 1946 3068 1952 3120
rect 2004 3108 2010 3120
rect 2685 3111 2743 3117
rect 2685 3108 2697 3111
rect 2004 3080 2697 3108
rect 2004 3068 2010 3080
rect 2685 3077 2697 3080
rect 2731 3108 2743 3111
rect 3697 3111 3755 3117
rect 3697 3108 3709 3111
rect 2731 3080 3709 3108
rect 2731 3077 2743 3080
rect 2685 3071 2743 3077
rect 3697 3077 3709 3080
rect 3743 3077 3755 3111
rect 3697 3071 3755 3077
rect 4065 3111 4123 3117
rect 4065 3077 4077 3111
rect 4111 3108 4123 3111
rect 6917 3111 6975 3117
rect 6917 3108 6929 3111
rect 4111 3080 6929 3108
rect 4111 3077 4123 3080
rect 4065 3071 4123 3077
rect 6917 3077 6929 3080
rect 6963 3077 6975 3111
rect 6917 3071 6975 3077
rect 7374 3068 7380 3120
rect 7432 3108 7438 3120
rect 7653 3111 7711 3117
rect 7653 3108 7665 3111
rect 7432 3080 7665 3108
rect 7432 3068 7438 3080
rect 7653 3077 7665 3080
rect 7699 3077 7711 3111
rect 7653 3071 7711 3077
rect 1486 3000 1492 3052
rect 1544 3040 1550 3052
rect 2225 3043 2283 3049
rect 2225 3040 2237 3043
rect 1544 3012 2237 3040
rect 1544 3000 1550 3012
rect 1964 2836 1992 3012
rect 2225 3009 2237 3012
rect 2271 3009 2283 3043
rect 2225 3003 2283 3009
rect 2869 3043 2927 3049
rect 2869 3009 2881 3043
rect 2915 3009 2927 3043
rect 2869 3003 2927 3009
rect 2884 2972 2912 3003
rect 2958 3000 2964 3052
rect 3016 3040 3022 3052
rect 3326 3040 3332 3052
rect 3016 3012 3061 3040
rect 3160 3012 3332 3040
rect 3016 3000 3022 3012
rect 3160 2972 3188 3012
rect 3326 3000 3332 3012
rect 3384 3040 3390 3052
rect 3878 3040 3884 3052
rect 3384 3012 3884 3040
rect 3384 3000 3390 3012
rect 3878 3000 3884 3012
rect 3936 3000 3942 3052
rect 4249 3043 4307 3049
rect 4249 3009 4261 3043
rect 4295 3040 4307 3043
rect 4430 3040 4436 3052
rect 4295 3012 4436 3040
rect 4295 3009 4307 3012
rect 4249 3003 4307 3009
rect 4430 3000 4436 3012
rect 4488 3000 4494 3052
rect 4614 3000 4620 3052
rect 4672 3040 4678 3052
rect 4893 3043 4951 3049
rect 4893 3040 4905 3043
rect 4672 3012 4905 3040
rect 4672 3000 4678 3012
rect 4893 3009 4905 3012
rect 4939 3009 4951 3043
rect 5074 3040 5080 3052
rect 5035 3012 5080 3040
rect 4893 3003 4951 3009
rect 5074 3000 5080 3012
rect 5132 3000 5138 3052
rect 5813 3043 5871 3049
rect 5813 3009 5825 3043
rect 5859 3040 5871 3043
rect 6822 3040 6828 3052
rect 5859 3012 6828 3040
rect 5859 3009 5871 3012
rect 5813 3003 5871 3009
rect 6822 3000 6828 3012
rect 6880 3000 6886 3052
rect 7193 3043 7251 3049
rect 7193 3009 7205 3043
rect 7239 3040 7251 3043
rect 7760 3040 7788 3148
rect 9490 3136 9496 3148
rect 9548 3176 9554 3188
rect 10686 3176 10692 3188
rect 9548 3148 10692 3176
rect 9548 3136 9554 3148
rect 10686 3136 10692 3148
rect 10744 3136 10750 3188
rect 11514 3136 11520 3188
rect 11572 3176 11578 3188
rect 12437 3179 12495 3185
rect 12437 3176 12449 3179
rect 11572 3148 12449 3176
rect 11572 3136 11578 3148
rect 12437 3145 12449 3148
rect 12483 3145 12495 3179
rect 12437 3139 12495 3145
rect 12618 3136 12624 3188
rect 12676 3176 12682 3188
rect 12676 3148 13952 3176
rect 12676 3136 12682 3148
rect 8110 3108 8116 3120
rect 7239 3012 7788 3040
rect 7852 3080 8116 3108
rect 7239 3009 7251 3012
rect 7193 3003 7251 3009
rect 2884 2944 3188 2972
rect 2041 2907 2099 2913
rect 2041 2873 2053 2907
rect 2087 2904 2099 2907
rect 2774 2904 2780 2916
rect 2087 2876 2780 2904
rect 2087 2873 2099 2876
rect 2041 2867 2099 2873
rect 2774 2864 2780 2876
rect 2832 2864 2838 2916
rect 7374 2904 7380 2916
rect 3068 2876 7380 2904
rect 3068 2836 3096 2876
rect 7374 2864 7380 2876
rect 7432 2864 7438 2916
rect 7653 2907 7711 2913
rect 7653 2873 7665 2907
rect 7699 2904 7711 2907
rect 7852 2904 7880 3080
rect 8110 3068 8116 3080
rect 8168 3068 8174 3120
rect 8662 3068 8668 3120
rect 8720 3108 8726 3120
rect 8720 3080 9076 3108
rect 8720 3068 8726 3080
rect 8754 3040 8760 3052
rect 8715 3012 8760 3040
rect 8754 3000 8760 3012
rect 8812 3000 8818 3052
rect 9048 3049 9076 3080
rect 9214 3068 9220 3120
rect 9272 3108 9278 3120
rect 13924 3108 13952 3148
rect 14182 3136 14188 3188
rect 14240 3176 14246 3188
rect 16853 3179 16911 3185
rect 16853 3176 16865 3179
rect 14240 3148 16865 3176
rect 14240 3136 14246 3148
rect 16853 3145 16865 3148
rect 16899 3145 16911 3179
rect 16853 3139 16911 3145
rect 16942 3136 16948 3188
rect 17000 3176 17006 3188
rect 17221 3179 17279 3185
rect 17221 3176 17233 3179
rect 17000 3148 17233 3176
rect 17000 3136 17006 3148
rect 17221 3145 17233 3148
rect 17267 3176 17279 3179
rect 17494 3176 17500 3188
rect 17267 3148 17500 3176
rect 17267 3145 17279 3148
rect 17221 3139 17279 3145
rect 17494 3136 17500 3148
rect 17552 3136 17558 3188
rect 22186 3176 22192 3188
rect 22147 3148 22192 3176
rect 22186 3136 22192 3148
rect 22244 3136 22250 3188
rect 25222 3176 25228 3188
rect 25183 3148 25228 3176
rect 25222 3136 25228 3148
rect 25280 3136 25286 3188
rect 25498 3136 25504 3188
rect 25556 3176 25562 3188
rect 25866 3176 25872 3188
rect 25556 3148 25872 3176
rect 25556 3136 25562 3148
rect 25866 3136 25872 3148
rect 25924 3136 25930 3188
rect 26421 3179 26479 3185
rect 26421 3145 26433 3179
rect 26467 3176 26479 3179
rect 28994 3176 29000 3188
rect 26467 3148 29000 3176
rect 26467 3145 26479 3148
rect 26421 3139 26479 3145
rect 28994 3136 29000 3148
rect 29052 3176 29058 3188
rect 33778 3176 33784 3188
rect 29052 3148 33784 3176
rect 29052 3136 29058 3148
rect 33778 3136 33784 3148
rect 33836 3136 33842 3188
rect 34882 3176 34888 3188
rect 34440 3148 34888 3176
rect 14366 3108 14372 3120
rect 9272 3080 12020 3108
rect 13924 3080 14372 3108
rect 9272 3068 9278 3080
rect 9033 3043 9091 3049
rect 9033 3009 9045 3043
rect 9079 3009 9091 3043
rect 9033 3003 9091 3009
rect 9398 3000 9404 3052
rect 9456 3040 9462 3052
rect 9493 3043 9551 3049
rect 11517 3046 11575 3049
rect 9493 3040 9505 3043
rect 9456 3012 9505 3040
rect 9456 3000 9462 3012
rect 9493 3009 9505 3012
rect 9539 3009 9551 3043
rect 11348 3043 11575 3046
rect 11348 3040 11529 3043
rect 9493 3003 9551 3009
rect 9600 3018 11529 3040
rect 9600 3012 11376 3018
rect 9214 2932 9220 2984
rect 9272 2972 9278 2984
rect 9600 2972 9628 3012
rect 11517 3009 11529 3018
rect 11563 3009 11575 3043
rect 11517 3003 11575 3009
rect 11698 3000 11704 3052
rect 11756 3040 11762 3052
rect 11793 3043 11851 3049
rect 11793 3040 11805 3043
rect 11756 3012 11805 3040
rect 11756 3000 11762 3012
rect 11793 3009 11805 3012
rect 11839 3009 11851 3043
rect 11793 3003 11851 3009
rect 9272 2944 9628 2972
rect 9769 2975 9827 2981
rect 9272 2932 9278 2944
rect 9769 2941 9781 2975
rect 9815 2972 9827 2975
rect 10594 2972 10600 2984
rect 9815 2944 10600 2972
rect 9815 2941 9827 2944
rect 9769 2935 9827 2941
rect 10594 2932 10600 2944
rect 10652 2932 10658 2984
rect 10778 2932 10784 2984
rect 10836 2972 10842 2984
rect 11609 2975 11667 2981
rect 11609 2972 11621 2975
rect 10836 2944 11621 2972
rect 10836 2932 10842 2944
rect 11609 2941 11621 2944
rect 11655 2941 11667 2975
rect 11609 2935 11667 2941
rect 7699 2876 7880 2904
rect 7699 2873 7711 2876
rect 7653 2867 7711 2873
rect 8478 2864 8484 2916
rect 8536 2904 8542 2916
rect 8754 2904 8760 2916
rect 8536 2876 8760 2904
rect 8536 2864 8542 2876
rect 8754 2864 8760 2876
rect 8812 2864 8818 2916
rect 8846 2864 8852 2916
rect 8904 2904 8910 2916
rect 9582 2904 9588 2916
rect 8904 2876 9588 2904
rect 8904 2864 8910 2876
rect 9582 2864 9588 2876
rect 9640 2864 9646 2916
rect 11422 2864 11428 2916
rect 11480 2904 11486 2916
rect 11992 2913 12020 3080
rect 14366 3068 14372 3080
rect 14424 3068 14430 3120
rect 15102 3068 15108 3120
rect 15160 3108 15166 3120
rect 15197 3111 15255 3117
rect 15197 3108 15209 3111
rect 15160 3080 15209 3108
rect 15160 3068 15166 3080
rect 15197 3077 15209 3080
rect 15243 3077 15255 3111
rect 15473 3111 15531 3117
rect 15473 3108 15485 3111
rect 15197 3071 15255 3077
rect 15304 3080 15485 3108
rect 15304 3052 15332 3080
rect 15473 3077 15485 3080
rect 15519 3077 15531 3111
rect 15930 3108 15936 3120
rect 15891 3080 15936 3108
rect 15473 3071 15531 3077
rect 15930 3068 15936 3080
rect 15988 3068 15994 3120
rect 18782 3068 18788 3120
rect 18840 3108 18846 3120
rect 18877 3111 18935 3117
rect 18877 3108 18889 3111
rect 18840 3080 18889 3108
rect 18840 3068 18846 3080
rect 18877 3077 18889 3080
rect 18923 3077 18935 3111
rect 19058 3108 19064 3120
rect 19019 3080 19064 3108
rect 18877 3071 18935 3077
rect 13170 3000 13176 3052
rect 13228 3040 13234 3052
rect 13265 3043 13323 3049
rect 13265 3040 13277 3043
rect 13228 3012 13277 3040
rect 13228 3000 13234 3012
rect 13265 3009 13277 3012
rect 13311 3009 13323 3043
rect 13722 3040 13728 3052
rect 13683 3012 13728 3040
rect 13265 3003 13323 3009
rect 13722 3000 13728 3012
rect 13780 3000 13786 3052
rect 14461 3043 14519 3049
rect 14461 3009 14473 3043
rect 14507 3040 14519 3043
rect 14550 3040 14556 3052
rect 14507 3012 14556 3040
rect 14507 3009 14519 3012
rect 14461 3003 14519 3009
rect 14550 3000 14556 3012
rect 14608 3000 14614 3052
rect 15286 3000 15292 3052
rect 15344 3000 15350 3052
rect 15381 3043 15439 3049
rect 15381 3009 15393 3043
rect 15427 3040 15439 3043
rect 16022 3040 16028 3052
rect 15427 3012 16028 3040
rect 15427 3009 15439 3012
rect 15381 3003 15439 3009
rect 16022 3000 16028 3012
rect 16080 3000 16086 3052
rect 16574 3000 16580 3052
rect 16632 3040 16638 3052
rect 17037 3043 17095 3049
rect 17037 3040 17049 3043
rect 16632 3012 17049 3040
rect 16632 3000 16638 3012
rect 17037 3009 17049 3012
rect 17083 3009 17095 3043
rect 17037 3003 17095 3009
rect 17310 3000 17316 3052
rect 17368 3040 17374 3052
rect 17368 3012 17413 3040
rect 17368 3000 17374 3012
rect 18046 3000 18052 3052
rect 18104 3040 18110 3052
rect 18141 3043 18199 3049
rect 18141 3040 18153 3043
rect 18104 3012 18153 3040
rect 18104 3000 18110 3012
rect 18141 3009 18153 3012
rect 18187 3009 18199 3043
rect 18892 3040 18920 3071
rect 19058 3068 19064 3080
rect 19116 3068 19122 3120
rect 19518 3108 19524 3120
rect 19479 3080 19524 3108
rect 19518 3068 19524 3080
rect 19576 3068 19582 3120
rect 21269 3111 21327 3117
rect 21269 3077 21281 3111
rect 21315 3108 21327 3111
rect 22094 3108 22100 3120
rect 21315 3080 22100 3108
rect 21315 3077 21327 3080
rect 21269 3071 21327 3077
rect 22094 3068 22100 3080
rect 22152 3068 22158 3120
rect 23106 3068 23112 3120
rect 23164 3108 23170 3120
rect 27522 3108 27528 3120
rect 23164 3080 27528 3108
rect 23164 3068 23170 3080
rect 21818 3040 21824 3052
rect 18892 3012 21824 3040
rect 18141 3003 18199 3009
rect 21818 3000 21824 3012
rect 21876 3000 21882 3052
rect 21910 3000 21916 3052
rect 21968 3040 21974 3052
rect 22005 3043 22063 3049
rect 22005 3040 22017 3043
rect 21968 3012 22017 3040
rect 21968 3000 21974 3012
rect 22005 3009 22017 3012
rect 22051 3009 22063 3043
rect 23014 3040 23020 3052
rect 22975 3012 23020 3040
rect 22005 3003 22063 3009
rect 23014 3000 23020 3012
rect 23072 3000 23078 3052
rect 23753 3043 23811 3049
rect 23753 3009 23765 3043
rect 23799 3040 23811 3043
rect 24578 3040 24584 3052
rect 23799 3012 24584 3040
rect 23799 3009 23811 3012
rect 23753 3003 23811 3009
rect 24578 3000 24584 3012
rect 24636 3000 24642 3052
rect 25498 3040 25504 3052
rect 25459 3012 25504 3040
rect 25498 3000 25504 3012
rect 25556 3000 25562 3052
rect 25608 3049 25636 3080
rect 27522 3068 27528 3080
rect 27580 3068 27586 3120
rect 27801 3111 27859 3117
rect 27801 3077 27813 3111
rect 27847 3108 27859 3111
rect 28166 3108 28172 3120
rect 27847 3080 28172 3108
rect 27847 3077 27859 3080
rect 27801 3071 27859 3077
rect 28166 3068 28172 3080
rect 28224 3068 28230 3120
rect 30377 3111 30435 3117
rect 30377 3077 30389 3111
rect 30423 3108 30435 3111
rect 30466 3108 30472 3120
rect 30423 3080 30472 3108
rect 30423 3077 30435 3080
rect 30377 3071 30435 3077
rect 30466 3068 30472 3080
rect 30524 3068 30530 3120
rect 31294 3108 31300 3120
rect 31131 3080 31300 3108
rect 25593 3043 25651 3049
rect 25593 3009 25605 3043
rect 25639 3009 25651 3043
rect 25593 3003 25651 3009
rect 25682 3000 25688 3052
rect 25740 3040 25746 3052
rect 25740 3012 25785 3040
rect 25740 3000 25746 3012
rect 25866 3000 25872 3052
rect 25924 3040 25930 3052
rect 27706 3040 27712 3052
rect 25924 3012 25969 3040
rect 27667 3012 27712 3040
rect 25924 3000 25930 3012
rect 27706 3000 27712 3012
rect 27764 3000 27770 3052
rect 27893 3043 27951 3049
rect 27893 3009 27905 3043
rect 27939 3040 27951 3043
rect 29270 3040 29276 3052
rect 27939 3012 29276 3040
rect 27939 3009 27951 3012
rect 27893 3003 27951 3009
rect 29270 3000 29276 3012
rect 29328 3000 29334 3052
rect 30834 3040 30840 3052
rect 30795 3012 30840 3040
rect 30834 3000 30840 3012
rect 30892 3000 30898 3052
rect 31018 3043 31024 3055
rect 30979 3015 31024 3043
rect 31018 3003 31024 3015
rect 31076 3003 31082 3055
rect 31131 3052 31159 3080
rect 31294 3068 31300 3080
rect 31352 3068 31358 3120
rect 31481 3111 31539 3117
rect 31481 3077 31493 3111
rect 31527 3108 31539 3111
rect 32214 3108 32220 3120
rect 31527 3080 32220 3108
rect 31527 3077 31539 3080
rect 31481 3071 31539 3077
rect 32214 3068 32220 3080
rect 32272 3068 32278 3120
rect 32490 3108 32496 3120
rect 32451 3080 32496 3108
rect 32490 3068 32496 3080
rect 32548 3068 32554 3120
rect 31116 3046 31174 3052
rect 31116 3012 31128 3046
rect 31162 3012 31174 3046
rect 31116 3006 31174 3012
rect 31202 3000 31208 3052
rect 31260 3040 31266 3052
rect 31260 3012 31305 3040
rect 31260 3000 31266 3012
rect 31570 3000 31576 3052
rect 31628 3040 31634 3052
rect 34440 3040 34468 3148
rect 34882 3136 34888 3148
rect 34940 3136 34946 3188
rect 36722 3176 36728 3188
rect 36683 3148 36728 3176
rect 36722 3136 36728 3148
rect 36780 3136 36786 3188
rect 36814 3136 36820 3188
rect 36872 3176 36878 3188
rect 37277 3179 37335 3185
rect 37277 3176 37289 3179
rect 36872 3148 37289 3176
rect 36872 3136 36878 3148
rect 37277 3145 37289 3148
rect 37323 3145 37335 3179
rect 37277 3139 37335 3145
rect 37384 3148 37596 3176
rect 34514 3068 34520 3120
rect 34572 3108 34578 3120
rect 35526 3108 35532 3120
rect 34572 3080 35532 3108
rect 34572 3068 34578 3080
rect 35526 3068 35532 3080
rect 35584 3068 35590 3120
rect 31628 3012 34468 3040
rect 34701 3043 34759 3049
rect 31628 3000 31634 3012
rect 34701 3009 34713 3043
rect 34747 3040 34759 3043
rect 34790 3040 34796 3052
rect 34747 3012 34796 3040
rect 34747 3009 34759 3012
rect 34701 3003 34759 3009
rect 34790 3000 34796 3012
rect 34848 3000 34854 3052
rect 35989 3043 36047 3049
rect 35989 3040 36001 3043
rect 34900 3012 36001 3040
rect 13630 2932 13636 2984
rect 13688 2972 13694 2984
rect 14918 2972 14924 2984
rect 13688 2944 14924 2972
rect 13688 2932 13694 2944
rect 14918 2932 14924 2944
rect 14976 2932 14982 2984
rect 19334 2972 19340 2984
rect 15856 2944 19340 2972
rect 11977 2907 12035 2913
rect 11480 2876 11652 2904
rect 11480 2864 11486 2876
rect 3234 2836 3240 2848
rect 1964 2808 3096 2836
rect 3195 2808 3240 2836
rect 3234 2796 3240 2808
rect 3292 2796 3298 2848
rect 5629 2839 5687 2845
rect 5629 2805 5641 2839
rect 5675 2836 5687 2839
rect 10410 2836 10416 2848
rect 5675 2808 10416 2836
rect 5675 2805 5687 2808
rect 5629 2799 5687 2805
rect 10410 2796 10416 2808
rect 10468 2796 10474 2848
rect 10962 2836 10968 2848
rect 10923 2808 10968 2836
rect 10962 2796 10968 2808
rect 11020 2796 11026 2848
rect 11330 2796 11336 2848
rect 11388 2836 11394 2848
rect 11517 2839 11575 2845
rect 11517 2836 11529 2839
rect 11388 2808 11529 2836
rect 11388 2796 11394 2808
rect 11517 2805 11529 2808
rect 11563 2805 11575 2839
rect 11624 2836 11652 2876
rect 11977 2873 11989 2907
rect 12023 2873 12035 2907
rect 13909 2907 13967 2913
rect 13909 2904 13921 2907
rect 11977 2867 12035 2873
rect 12084 2876 13921 2904
rect 12084 2836 12112 2876
rect 13909 2873 13921 2876
rect 13955 2873 13967 2907
rect 13909 2867 13967 2873
rect 14645 2907 14703 2913
rect 14645 2873 14657 2907
rect 14691 2904 14703 2907
rect 15856 2904 15884 2944
rect 19334 2932 19340 2944
rect 19392 2932 19398 2984
rect 24302 2972 24308 2984
rect 22066 2944 24308 2972
rect 14691 2876 15884 2904
rect 14691 2873 14703 2876
rect 14645 2867 14703 2873
rect 15930 2864 15936 2916
rect 15988 2904 15994 2916
rect 15988 2876 16033 2904
rect 15988 2864 15994 2876
rect 17770 2864 17776 2916
rect 17828 2904 17834 2916
rect 22066 2904 22094 2944
rect 24302 2932 24308 2944
rect 24360 2932 24366 2984
rect 24765 2975 24823 2981
rect 24765 2941 24777 2975
rect 24811 2972 24823 2975
rect 28718 2972 28724 2984
rect 24811 2944 28724 2972
rect 24811 2941 24823 2944
rect 24765 2935 24823 2941
rect 28718 2932 28724 2944
rect 28776 2932 28782 2984
rect 28997 2975 29055 2981
rect 28997 2941 29009 2975
rect 29043 2972 29055 2975
rect 29086 2972 29092 2984
rect 29043 2944 29092 2972
rect 29043 2941 29055 2944
rect 28997 2935 29055 2941
rect 29086 2932 29092 2944
rect 29144 2972 29150 2984
rect 29362 2972 29368 2984
rect 29144 2944 29368 2972
rect 29144 2932 29150 2944
rect 29362 2932 29368 2944
rect 29420 2932 29426 2984
rect 30742 2932 30748 2984
rect 30800 2972 30806 2984
rect 31220 2972 31248 3000
rect 30800 2944 31248 2972
rect 30800 2932 30806 2944
rect 31294 2932 31300 2984
rect 31352 2972 31358 2984
rect 31588 2972 31616 3000
rect 31352 2944 31616 2972
rect 31352 2932 31358 2944
rect 32306 2932 32312 2984
rect 32364 2972 32370 2984
rect 34900 2972 34928 3012
rect 35989 3009 36001 3012
rect 36035 3009 36047 3043
rect 35989 3003 36047 3009
rect 36814 3000 36820 3052
rect 36872 3040 36878 3052
rect 37384 3040 37412 3148
rect 37568 3108 37596 3148
rect 39942 3136 39948 3188
rect 40000 3176 40006 3188
rect 40865 3179 40923 3185
rect 40865 3176 40877 3179
rect 40000 3148 40877 3176
rect 40000 3136 40006 3148
rect 40865 3145 40877 3148
rect 40911 3176 40923 3179
rect 41046 3176 41052 3188
rect 40911 3148 41052 3176
rect 40911 3145 40923 3148
rect 40865 3139 40923 3145
rect 41046 3136 41052 3148
rect 41104 3136 41110 3188
rect 41233 3179 41291 3185
rect 41233 3145 41245 3179
rect 41279 3176 41291 3179
rect 43898 3176 43904 3188
rect 41279 3148 43904 3176
rect 41279 3145 41291 3148
rect 41233 3139 41291 3145
rect 43898 3136 43904 3148
rect 43956 3136 43962 3188
rect 43990 3136 43996 3188
rect 44048 3176 44054 3188
rect 45002 3176 45008 3188
rect 44048 3148 45008 3176
rect 44048 3136 44054 3148
rect 45002 3136 45008 3148
rect 45060 3136 45066 3188
rect 45830 3136 45836 3188
rect 45888 3176 45894 3188
rect 45888 3148 51304 3176
rect 45888 3136 45894 3148
rect 37568 3080 41736 3108
rect 36872 3012 37412 3040
rect 36872 3000 36878 3012
rect 37458 3000 37464 3052
rect 37516 3040 37522 3052
rect 37642 3040 37648 3052
rect 37516 3012 37561 3040
rect 37603 3012 37648 3040
rect 37516 3000 37522 3012
rect 37642 3000 37648 3012
rect 37700 3000 37706 3052
rect 37734 3000 37740 3052
rect 37792 3040 37798 3052
rect 40129 3043 40187 3049
rect 40129 3040 40141 3043
rect 37792 3012 37837 3040
rect 37936 3012 40141 3040
rect 37792 3000 37798 3012
rect 32364 2944 34928 2972
rect 34977 2975 35035 2981
rect 32364 2932 32370 2944
rect 34977 2941 34989 2975
rect 35023 2972 35035 2975
rect 35802 2972 35808 2984
rect 35023 2944 35808 2972
rect 35023 2941 35035 2944
rect 34977 2935 35035 2941
rect 35802 2932 35808 2944
rect 35860 2932 35866 2984
rect 35894 2932 35900 2984
rect 35952 2972 35958 2984
rect 37936 2972 37964 3012
rect 40129 3009 40141 3012
rect 40175 3009 40187 3043
rect 40770 3040 40776 3052
rect 40731 3012 40776 3040
rect 40129 3003 40187 3009
rect 40770 3000 40776 3012
rect 40828 3000 40834 3052
rect 41046 3040 41052 3052
rect 41007 3012 41052 3040
rect 41046 3000 41052 3012
rect 41104 3000 41110 3052
rect 41708 3049 41736 3080
rect 42886 3068 42892 3120
rect 42944 3108 42950 3120
rect 43806 3108 43812 3120
rect 42944 3080 43300 3108
rect 43767 3080 43812 3108
rect 42944 3068 42950 3080
rect 41693 3043 41751 3049
rect 41693 3009 41705 3043
rect 41739 3009 41751 3043
rect 41693 3003 41751 3009
rect 42610 3000 42616 3052
rect 42668 3040 42674 3052
rect 43165 3043 43223 3049
rect 42996 3040 43177 3043
rect 42668 3015 43177 3040
rect 42668 3012 43024 3015
rect 42668 3000 42674 3012
rect 43165 3009 43177 3015
rect 43211 3009 43223 3043
rect 43272 3040 43300 3080
rect 43806 3068 43812 3080
rect 43864 3068 43870 3120
rect 45094 3068 45100 3120
rect 45152 3108 45158 3120
rect 49246 3111 49304 3117
rect 49246 3108 49258 3111
rect 45152 3080 49258 3108
rect 45152 3068 45158 3080
rect 49246 3077 49258 3080
rect 49292 3077 49304 3111
rect 49246 3071 49304 3077
rect 49418 3068 49424 3120
rect 49476 3108 49482 3120
rect 49476 3080 49740 3108
rect 49476 3068 49482 3080
rect 43622 3049 43628 3052
rect 43344 3043 43402 3049
rect 43344 3040 43356 3043
rect 43272 3012 43356 3040
rect 43165 3003 43223 3009
rect 43344 3009 43356 3012
rect 43390 3009 43402 3043
rect 43444 3043 43502 3049
rect 43444 3040 43456 3043
rect 43344 3003 43402 3009
rect 43443 3009 43456 3040
rect 43490 3009 43502 3043
rect 43443 3003 43502 3009
rect 43579 3043 43628 3049
rect 43579 3009 43591 3043
rect 43625 3009 43628 3043
rect 43579 3003 43628 3009
rect 35952 2944 37964 2972
rect 35952 2932 35958 2944
rect 38286 2932 38292 2984
rect 38344 2972 38350 2984
rect 39666 2972 39672 2984
rect 38344 2944 39672 2972
rect 38344 2932 38350 2944
rect 39666 2932 39672 2944
rect 39724 2932 39730 2984
rect 42702 2932 42708 2984
rect 42760 2972 42766 2984
rect 43443 2972 43471 3003
rect 43622 3000 43628 3003
rect 43680 3000 43686 3052
rect 44174 3000 44180 3052
rect 44232 3040 44238 3052
rect 44269 3043 44327 3049
rect 44269 3040 44281 3043
rect 44232 3012 44281 3040
rect 44232 3000 44238 3012
rect 44269 3009 44281 3012
rect 44315 3009 44327 3043
rect 44269 3003 44327 3009
rect 45002 3000 45008 3052
rect 45060 3040 45066 3052
rect 49513 3043 49571 3049
rect 45060 3012 49464 3040
rect 45060 3000 45066 3012
rect 47578 2972 47584 2984
rect 42760 2944 43471 2972
rect 47539 2944 47584 2972
rect 42760 2932 42766 2944
rect 47578 2932 47584 2944
rect 47636 2932 47642 2984
rect 49436 2972 49464 3012
rect 49513 3009 49525 3043
rect 49559 3040 49571 3043
rect 49602 3040 49608 3052
rect 49559 3012 49608 3040
rect 49559 3009 49571 3012
rect 49513 3003 49571 3009
rect 49602 3000 49608 3012
rect 49660 3000 49666 3052
rect 49712 3040 49740 3080
rect 51276 3049 51304 3148
rect 52822 3136 52828 3188
rect 52880 3176 52886 3188
rect 52917 3179 52975 3185
rect 52917 3176 52929 3179
rect 52880 3148 52929 3176
rect 52880 3136 52886 3148
rect 52917 3145 52929 3148
rect 52963 3145 52975 3179
rect 52917 3139 52975 3145
rect 57790 3136 57796 3188
rect 57848 3176 57854 3188
rect 57885 3179 57943 3185
rect 57885 3176 57897 3179
rect 57848 3148 57897 3176
rect 57848 3136 57854 3148
rect 57885 3145 57897 3148
rect 57931 3145 57943 3179
rect 57885 3139 57943 3145
rect 51261 3043 51319 3049
rect 49712 3012 50936 3040
rect 50617 2975 50675 2981
rect 50617 2972 50629 2975
rect 49436 2944 49556 2972
rect 17828 2876 22094 2904
rect 17828 2864 17834 2876
rect 22278 2864 22284 2916
rect 22336 2904 22342 2916
rect 23569 2907 23627 2913
rect 23569 2904 23581 2907
rect 22336 2876 23581 2904
rect 22336 2864 22342 2876
rect 23569 2873 23581 2876
rect 23615 2873 23627 2907
rect 23569 2867 23627 2873
rect 25314 2864 25320 2916
rect 25372 2904 25378 2916
rect 25498 2904 25504 2916
rect 25372 2876 25504 2904
rect 25372 2864 25378 2876
rect 25498 2864 25504 2876
rect 25556 2904 25562 2916
rect 25774 2904 25780 2916
rect 25556 2876 25780 2904
rect 25556 2864 25562 2876
rect 25774 2864 25780 2876
rect 25832 2864 25838 2916
rect 25958 2864 25964 2916
rect 26016 2904 26022 2916
rect 28353 2907 28411 2913
rect 28353 2904 28365 2907
rect 26016 2876 28365 2904
rect 26016 2864 26022 2876
rect 28353 2873 28365 2876
rect 28399 2873 28411 2907
rect 28353 2867 28411 2873
rect 31202 2864 31208 2916
rect 31260 2904 31266 2916
rect 31260 2876 31616 2904
rect 31260 2864 31266 2876
rect 11624 2808 12112 2836
rect 13081 2839 13139 2845
rect 11517 2799 11575 2805
rect 13081 2805 13093 2839
rect 13127 2836 13139 2839
rect 13446 2836 13452 2848
rect 13127 2808 13452 2836
rect 13127 2805 13139 2808
rect 13081 2799 13139 2805
rect 13446 2796 13452 2808
rect 13504 2796 13510 2848
rect 16022 2796 16028 2848
rect 16080 2836 16086 2848
rect 16206 2836 16212 2848
rect 16080 2808 16212 2836
rect 16080 2796 16086 2808
rect 16206 2796 16212 2808
rect 16264 2796 16270 2848
rect 17954 2836 17960 2848
rect 17915 2808 17960 2836
rect 17954 2796 17960 2808
rect 18012 2796 18018 2848
rect 21542 2796 21548 2848
rect 21600 2836 21606 2848
rect 22002 2836 22008 2848
rect 21600 2808 22008 2836
rect 21600 2796 21606 2808
rect 22002 2796 22008 2808
rect 22060 2796 22066 2848
rect 22462 2796 22468 2848
rect 22520 2836 22526 2848
rect 22833 2839 22891 2845
rect 22833 2836 22845 2839
rect 22520 2808 22845 2836
rect 22520 2796 22526 2808
rect 22833 2805 22845 2808
rect 22879 2805 22891 2839
rect 22833 2799 22891 2805
rect 26786 2796 26792 2848
rect 26844 2836 26850 2848
rect 26973 2839 27031 2845
rect 26973 2836 26985 2839
rect 26844 2808 26985 2836
rect 26844 2796 26850 2808
rect 26973 2805 26985 2808
rect 27019 2805 27031 2839
rect 31588 2836 31616 2876
rect 31754 2864 31760 2916
rect 31812 2904 31818 2916
rect 35342 2904 35348 2916
rect 31812 2876 35348 2904
rect 31812 2864 31818 2876
rect 35342 2864 35348 2876
rect 35400 2864 35406 2916
rect 38197 2907 38255 2913
rect 38197 2904 38209 2907
rect 35452 2876 38209 2904
rect 33962 2836 33968 2848
rect 31588 2808 33968 2836
rect 26973 2799 27031 2805
rect 33962 2796 33968 2808
rect 34020 2796 34026 2848
rect 34238 2796 34244 2848
rect 34296 2836 34302 2848
rect 35452 2836 35480 2876
rect 38197 2873 38209 2876
rect 38243 2873 38255 2907
rect 42429 2907 42487 2913
rect 42429 2904 42441 2907
rect 38197 2867 38255 2873
rect 41524 2876 42441 2904
rect 34296 2808 35480 2836
rect 34296 2796 34302 2808
rect 35526 2796 35532 2848
rect 35584 2836 35590 2848
rect 38841 2839 38899 2845
rect 38841 2836 38853 2839
rect 35584 2808 38853 2836
rect 35584 2796 35590 2808
rect 38841 2805 38853 2808
rect 38887 2805 38899 2839
rect 39482 2836 39488 2848
rect 39443 2808 39488 2836
rect 38841 2799 38899 2805
rect 39482 2796 39488 2808
rect 39540 2796 39546 2848
rect 39666 2796 39672 2848
rect 39724 2836 39730 2848
rect 41524 2836 41552 2876
rect 42429 2873 42441 2876
rect 42475 2873 42487 2907
rect 42429 2867 42487 2873
rect 43254 2864 43260 2916
rect 43312 2904 43318 2916
rect 45278 2904 45284 2916
rect 43312 2876 45284 2904
rect 43312 2864 43318 2876
rect 45278 2864 45284 2876
rect 45336 2864 45342 2916
rect 45738 2864 45744 2916
rect 45796 2904 45802 2916
rect 48133 2907 48191 2913
rect 48133 2904 48145 2907
rect 45796 2876 48145 2904
rect 45796 2864 45802 2876
rect 48133 2873 48145 2876
rect 48179 2873 48191 2907
rect 49528 2904 49556 2944
rect 49896 2944 50629 2972
rect 49896 2904 49924 2944
rect 50617 2941 50629 2944
rect 50663 2941 50675 2975
rect 50617 2935 50675 2941
rect 49528 2876 49924 2904
rect 48133 2867 48191 2873
rect 50154 2864 50160 2916
rect 50212 2904 50218 2916
rect 50908 2904 50936 3012
rect 51261 3009 51273 3043
rect 51307 3009 51319 3043
rect 51261 3003 51319 3009
rect 52362 3000 52368 3052
rect 52420 3040 52426 3052
rect 52822 3040 52828 3052
rect 52420 3012 52828 3040
rect 52420 3000 52426 3012
rect 52822 3000 52828 3012
rect 52880 3000 52886 3052
rect 52917 3043 52975 3049
rect 52917 3009 52929 3043
rect 52963 3040 52975 3043
rect 53098 3040 53104 3052
rect 52963 3012 53104 3040
rect 52963 3009 52975 3012
rect 52917 3003 52975 3009
rect 53098 3000 53104 3012
rect 53156 3040 53162 3052
rect 53926 3040 53932 3052
rect 53156 3012 53932 3040
rect 53156 3000 53162 3012
rect 53926 3000 53932 3012
rect 53984 3000 53990 3052
rect 54110 3040 54116 3052
rect 54071 3012 54116 3040
rect 54110 3000 54116 3012
rect 54168 3000 54174 3052
rect 54754 3040 54760 3052
rect 54715 3012 54760 3040
rect 54754 3000 54760 3012
rect 54812 3000 54818 3052
rect 53469 2975 53527 2981
rect 53469 2972 53481 2975
rect 52104 2944 53481 2972
rect 51905 2907 51963 2913
rect 51905 2904 51917 2907
rect 50212 2876 50752 2904
rect 50908 2876 51917 2904
rect 50212 2864 50218 2876
rect 39724 2808 41552 2836
rect 39724 2796 39730 2808
rect 41690 2796 41696 2848
rect 41748 2836 41754 2848
rect 44542 2836 44548 2848
rect 41748 2808 44548 2836
rect 41748 2796 41754 2808
rect 44542 2796 44548 2808
rect 44600 2796 44606 2848
rect 44910 2836 44916 2848
rect 44871 2808 44916 2836
rect 44910 2796 44916 2808
rect 44968 2796 44974 2848
rect 45557 2839 45615 2845
rect 45557 2805 45569 2839
rect 45603 2836 45615 2839
rect 45646 2836 45652 2848
rect 45603 2808 45652 2836
rect 45603 2805 45615 2808
rect 45557 2799 45615 2805
rect 45646 2796 45652 2808
rect 45704 2796 45710 2848
rect 46198 2836 46204 2848
rect 46159 2808 46204 2836
rect 46198 2796 46204 2808
rect 46256 2796 46262 2848
rect 46842 2836 46848 2848
rect 46803 2808 46848 2836
rect 46842 2796 46848 2808
rect 46900 2796 46906 2848
rect 48774 2796 48780 2848
rect 48832 2836 48838 2848
rect 49326 2836 49332 2848
rect 48832 2808 49332 2836
rect 48832 2796 48838 2808
rect 49326 2796 49332 2808
rect 49384 2796 49390 2848
rect 49970 2836 49976 2848
rect 49931 2808 49976 2836
rect 49970 2796 49976 2808
rect 50028 2796 50034 2848
rect 50724 2836 50752 2876
rect 51905 2873 51917 2876
rect 51951 2873 51963 2907
rect 51905 2867 51963 2873
rect 52104 2836 52132 2944
rect 53469 2941 53481 2944
rect 53515 2941 53527 2975
rect 56689 2975 56747 2981
rect 56689 2972 56701 2975
rect 53469 2935 53527 2941
rect 53576 2944 56701 2972
rect 52454 2864 52460 2916
rect 52512 2904 52518 2916
rect 53576 2904 53604 2944
rect 56689 2941 56701 2944
rect 56735 2941 56747 2975
rect 56689 2935 56747 2941
rect 52512 2876 53604 2904
rect 52512 2864 52518 2876
rect 53834 2864 53840 2916
rect 53892 2904 53898 2916
rect 55401 2907 55459 2913
rect 55401 2904 55413 2907
rect 53892 2876 55413 2904
rect 53892 2864 53898 2876
rect 55401 2873 55413 2876
rect 55447 2873 55459 2907
rect 55401 2867 55459 2873
rect 50724 2808 52132 2836
rect 52178 2796 52184 2848
rect 52236 2836 52242 2848
rect 56045 2839 56103 2845
rect 56045 2836 56057 2839
rect 52236 2808 56057 2836
rect 52236 2796 52242 2808
rect 56045 2805 56057 2808
rect 56091 2805 56103 2839
rect 56045 2799 56103 2805
rect 1104 2746 58880 2768
rect 1104 2694 8174 2746
rect 8226 2694 8238 2746
rect 8290 2694 8302 2746
rect 8354 2694 8366 2746
rect 8418 2694 8430 2746
rect 8482 2694 22622 2746
rect 22674 2694 22686 2746
rect 22738 2694 22750 2746
rect 22802 2694 22814 2746
rect 22866 2694 22878 2746
rect 22930 2694 37070 2746
rect 37122 2694 37134 2746
rect 37186 2694 37198 2746
rect 37250 2694 37262 2746
rect 37314 2694 37326 2746
rect 37378 2694 51518 2746
rect 51570 2694 51582 2746
rect 51634 2694 51646 2746
rect 51698 2694 51710 2746
rect 51762 2694 51774 2746
rect 51826 2694 58880 2746
rect 1104 2672 58880 2694
rect 1857 2635 1915 2641
rect 1857 2601 1869 2635
rect 1903 2632 1915 2635
rect 1946 2632 1952 2644
rect 1903 2604 1952 2632
rect 1903 2601 1915 2604
rect 1857 2595 1915 2601
rect 1946 2592 1952 2604
rect 2004 2592 2010 2644
rect 2958 2592 2964 2644
rect 3016 2632 3022 2644
rect 3053 2635 3111 2641
rect 3053 2632 3065 2635
rect 3016 2604 3065 2632
rect 3016 2592 3022 2604
rect 3053 2601 3065 2604
rect 3099 2601 3111 2635
rect 3053 2595 3111 2601
rect 4338 2592 4344 2644
rect 4396 2632 4402 2644
rect 4433 2635 4491 2641
rect 4433 2632 4445 2635
rect 4396 2604 4445 2632
rect 4396 2592 4402 2604
rect 4433 2601 4445 2604
rect 4479 2601 4491 2635
rect 4433 2595 4491 2601
rect 5810 2592 5816 2644
rect 5868 2632 5874 2644
rect 6730 2632 6736 2644
rect 5868 2604 6736 2632
rect 5868 2592 5874 2604
rect 6730 2592 6736 2604
rect 6788 2592 6794 2644
rect 6825 2635 6883 2641
rect 6825 2601 6837 2635
rect 6871 2632 6883 2635
rect 6871 2604 7236 2632
rect 6871 2601 6883 2604
rect 6825 2595 6883 2601
rect 3602 2564 3608 2576
rect 2056 2536 3608 2564
rect 2056 2437 2084 2536
rect 3602 2524 3608 2536
rect 3660 2524 3666 2576
rect 6546 2524 6552 2576
rect 6604 2564 6610 2576
rect 6641 2567 6699 2573
rect 6641 2564 6653 2567
rect 6604 2536 6653 2564
rect 6604 2524 6610 2536
rect 6641 2533 6653 2536
rect 6687 2533 6699 2567
rect 6641 2527 6699 2533
rect 2222 2496 2228 2508
rect 2183 2468 2228 2496
rect 2222 2456 2228 2468
rect 2280 2456 2286 2508
rect 2314 2456 2320 2508
rect 2372 2496 2378 2508
rect 6840 2496 6868 2595
rect 6914 2524 6920 2576
rect 6972 2564 6978 2576
rect 6972 2536 7052 2564
rect 6972 2524 6978 2536
rect 7024 2505 7052 2536
rect 2372 2468 2912 2496
rect 2372 2456 2378 2468
rect 2884 2437 2912 2468
rect 6380 2468 6868 2496
rect 7009 2499 7067 2505
rect 2041 2431 2099 2437
rect 2041 2397 2053 2431
rect 2087 2397 2099 2431
rect 2041 2391 2099 2397
rect 2685 2431 2743 2437
rect 2685 2397 2697 2431
rect 2731 2397 2743 2431
rect 2685 2391 2743 2397
rect 2869 2431 2927 2437
rect 2869 2397 2881 2431
rect 2915 2397 2927 2431
rect 3970 2428 3976 2440
rect 3931 2400 3976 2428
rect 2869 2391 2927 2397
rect 1670 2320 1676 2372
rect 1728 2360 1734 2372
rect 2700 2360 2728 2391
rect 3970 2388 3976 2400
rect 4028 2388 4034 2440
rect 5258 2388 5264 2440
rect 5316 2428 5322 2440
rect 5813 2431 5871 2437
rect 5813 2428 5825 2431
rect 5316 2400 5825 2428
rect 5316 2388 5322 2400
rect 5813 2397 5825 2400
rect 5859 2397 5871 2431
rect 5813 2391 5871 2397
rect 5534 2360 5540 2372
rect 5592 2369 5598 2372
rect 1728 2332 2728 2360
rect 5504 2332 5540 2360
rect 1728 2320 1734 2332
rect 5534 2320 5540 2332
rect 5592 2323 5604 2369
rect 5592 2320 5598 2323
rect 2590 2252 2596 2304
rect 2648 2292 2654 2304
rect 6380 2292 6408 2468
rect 7009 2465 7021 2499
rect 7055 2465 7067 2499
rect 7009 2459 7067 2465
rect 7098 2456 7104 2508
rect 7156 2456 7162 2508
rect 7208 2496 7236 2604
rect 8110 2592 8116 2644
rect 8168 2632 8174 2644
rect 8168 2604 10916 2632
rect 8168 2592 8174 2604
rect 8294 2524 8300 2576
rect 8352 2564 8358 2576
rect 9214 2564 9220 2576
rect 8352 2536 9220 2564
rect 8352 2524 8358 2536
rect 9214 2524 9220 2536
rect 9272 2524 9278 2576
rect 10888 2564 10916 2604
rect 10962 2592 10968 2644
rect 11020 2632 11026 2644
rect 17770 2632 17776 2644
rect 11020 2604 17776 2632
rect 11020 2592 11026 2604
rect 17770 2592 17776 2604
rect 17828 2592 17834 2644
rect 17865 2635 17923 2641
rect 17865 2601 17877 2635
rect 17911 2632 17923 2635
rect 21542 2632 21548 2644
rect 17911 2604 21548 2632
rect 17911 2601 17923 2604
rect 17865 2595 17923 2601
rect 21542 2592 21548 2604
rect 21600 2592 21606 2644
rect 22094 2592 22100 2644
rect 22152 2632 22158 2644
rect 27890 2632 27896 2644
rect 22152 2604 27896 2632
rect 22152 2592 22158 2604
rect 27890 2592 27896 2604
rect 27948 2592 27954 2644
rect 29546 2632 29552 2644
rect 28920 2604 29552 2632
rect 13814 2564 13820 2576
rect 10888 2536 13820 2564
rect 13814 2524 13820 2536
rect 13872 2524 13878 2576
rect 15654 2524 15660 2576
rect 15712 2564 15718 2576
rect 16206 2564 16212 2576
rect 15712 2536 16212 2564
rect 15712 2524 15718 2536
rect 16206 2524 16212 2536
rect 16264 2524 16270 2576
rect 17037 2567 17095 2573
rect 17037 2533 17049 2567
rect 17083 2564 17095 2567
rect 17083 2536 19932 2564
rect 17083 2533 17095 2536
rect 17037 2527 17095 2533
rect 9309 2499 9367 2505
rect 9309 2496 9321 2499
rect 7208 2468 9321 2496
rect 9309 2465 9321 2468
rect 9355 2465 9367 2499
rect 9309 2459 9367 2465
rect 9401 2499 9459 2505
rect 9401 2465 9413 2499
rect 9447 2496 9459 2499
rect 9490 2496 9496 2508
rect 9447 2468 9496 2496
rect 9447 2465 9459 2468
rect 9401 2459 9459 2465
rect 9490 2456 9496 2468
rect 9548 2456 9554 2508
rect 13262 2456 13268 2508
rect 13320 2496 13326 2508
rect 13320 2468 15884 2496
rect 13320 2456 13326 2468
rect 6825 2431 6883 2437
rect 6825 2397 6837 2431
rect 6871 2397 6883 2431
rect 7116 2428 7144 2456
rect 6825 2391 6883 2397
rect 7024 2400 7144 2428
rect 6840 2360 6868 2391
rect 7024 2360 7052 2400
rect 7190 2388 7196 2440
rect 7248 2428 7254 2440
rect 7466 2428 7472 2440
rect 7248 2400 7472 2428
rect 7248 2388 7254 2400
rect 7466 2388 7472 2400
rect 7524 2428 7530 2440
rect 7561 2431 7619 2437
rect 7561 2428 7573 2431
rect 7524 2400 7573 2428
rect 7524 2388 7530 2400
rect 7561 2397 7573 2400
rect 7607 2397 7619 2431
rect 7561 2391 7619 2397
rect 7837 2431 7895 2437
rect 7837 2397 7849 2431
rect 7883 2428 7895 2431
rect 8110 2428 8116 2440
rect 7883 2400 8116 2428
rect 7883 2397 7895 2400
rect 7837 2391 7895 2397
rect 8110 2388 8116 2400
rect 8168 2388 8174 2440
rect 9030 2428 9036 2440
rect 8404 2400 9036 2428
rect 6840 2332 7052 2360
rect 7101 2363 7159 2369
rect 7101 2329 7113 2363
rect 7147 2360 7159 2363
rect 8404 2360 8432 2400
rect 9030 2388 9036 2400
rect 9088 2428 9094 2440
rect 9125 2431 9183 2437
rect 9125 2428 9137 2431
rect 9088 2400 9137 2428
rect 9088 2388 9094 2400
rect 9125 2397 9137 2400
rect 9171 2397 9183 2431
rect 9125 2391 9183 2397
rect 9214 2388 9220 2440
rect 9272 2428 9278 2440
rect 9272 2400 9317 2428
rect 9272 2388 9278 2400
rect 7147 2332 8432 2360
rect 8941 2363 8999 2369
rect 7147 2329 7159 2332
rect 7101 2323 7159 2329
rect 8941 2329 8953 2363
rect 8987 2329 8999 2363
rect 8941 2323 8999 2329
rect 2648 2264 6408 2292
rect 2648 2252 2654 2264
rect 6730 2252 6736 2304
rect 6788 2292 6794 2304
rect 8956 2292 8984 2323
rect 9232 2304 9260 2388
rect 9508 2360 9536 2456
rect 10686 2428 10692 2440
rect 10647 2400 10692 2428
rect 10686 2388 10692 2400
rect 10744 2388 10750 2440
rect 10962 2428 10968 2440
rect 10923 2400 10968 2428
rect 10962 2388 10968 2400
rect 11020 2388 11026 2440
rect 11517 2431 11575 2437
rect 11517 2397 11529 2431
rect 11563 2428 11575 2431
rect 11606 2428 11612 2440
rect 11563 2400 11612 2428
rect 11563 2397 11575 2400
rect 11517 2391 11575 2397
rect 11606 2388 11612 2400
rect 11664 2388 11670 2440
rect 11790 2428 11796 2440
rect 11751 2400 11796 2428
rect 11790 2388 11796 2400
rect 11848 2388 11854 2440
rect 13538 2428 13544 2440
rect 13499 2400 13544 2428
rect 13538 2388 13544 2400
rect 13596 2388 13602 2440
rect 14366 2428 14372 2440
rect 14327 2400 14372 2428
rect 14366 2388 14372 2400
rect 14424 2388 14430 2440
rect 14550 2388 14556 2440
rect 14608 2428 14614 2440
rect 15856 2437 15884 2468
rect 17586 2456 17592 2508
rect 17644 2496 17650 2508
rect 18417 2499 18475 2505
rect 18417 2496 18429 2499
rect 17644 2468 18429 2496
rect 17644 2456 17650 2468
rect 18417 2465 18429 2468
rect 18463 2465 18475 2499
rect 18417 2459 18475 2465
rect 15105 2431 15163 2437
rect 15105 2428 15117 2431
rect 14608 2400 15117 2428
rect 14608 2388 14614 2400
rect 15105 2397 15117 2400
rect 15151 2397 15163 2431
rect 15105 2391 15163 2397
rect 15841 2431 15899 2437
rect 15841 2397 15853 2431
rect 15887 2397 15899 2431
rect 17218 2428 17224 2440
rect 17179 2400 17224 2428
rect 15841 2391 15899 2397
rect 17218 2388 17224 2400
rect 17276 2388 17282 2440
rect 17678 2428 17684 2440
rect 17639 2400 17684 2428
rect 17678 2388 17684 2400
rect 17736 2388 17742 2440
rect 18601 2431 18659 2437
rect 18601 2397 18613 2431
rect 18647 2428 18659 2431
rect 18690 2428 18696 2440
rect 18647 2400 18696 2428
rect 18647 2397 18659 2400
rect 18601 2391 18659 2397
rect 18690 2388 18696 2400
rect 18748 2388 18754 2440
rect 11330 2360 11336 2372
rect 9508 2332 11336 2360
rect 11330 2320 11336 2332
rect 11388 2320 11394 2372
rect 19904 2360 19932 2536
rect 21266 2524 21272 2576
rect 21324 2564 21330 2576
rect 24489 2567 24547 2573
rect 24489 2564 24501 2567
rect 21324 2536 22508 2564
rect 21324 2524 21330 2536
rect 22480 2496 22508 2536
rect 22756 2536 24501 2564
rect 22756 2496 22784 2536
rect 24489 2533 24501 2536
rect 24535 2533 24547 2567
rect 24489 2527 24547 2533
rect 25777 2567 25835 2573
rect 25777 2533 25789 2567
rect 25823 2564 25835 2567
rect 28920 2564 28948 2604
rect 29546 2592 29552 2604
rect 29604 2592 29610 2644
rect 31018 2592 31024 2644
rect 31076 2632 31082 2644
rect 31113 2635 31171 2641
rect 31113 2632 31125 2635
rect 31076 2604 31125 2632
rect 31076 2592 31082 2604
rect 31113 2601 31125 2604
rect 31159 2601 31171 2635
rect 33502 2632 33508 2644
rect 31113 2595 31171 2601
rect 31312 2604 33508 2632
rect 25823 2536 28948 2564
rect 28997 2567 29055 2573
rect 25823 2533 25835 2536
rect 25777 2527 25835 2533
rect 28997 2533 29009 2567
rect 29043 2564 29055 2567
rect 30650 2564 30656 2576
rect 29043 2536 30656 2564
rect 29043 2533 29055 2536
rect 28997 2527 29055 2533
rect 30650 2524 30656 2536
rect 30708 2524 30714 2576
rect 23566 2496 23572 2508
rect 22480 2468 22784 2496
rect 22848 2468 23572 2496
rect 20254 2428 20260 2440
rect 20215 2400 20260 2428
rect 20254 2388 20260 2400
rect 20312 2388 20318 2440
rect 20530 2428 20536 2440
rect 20491 2400 20536 2428
rect 20530 2388 20536 2400
rect 20588 2388 20594 2440
rect 21174 2388 21180 2440
rect 21232 2428 21238 2440
rect 21269 2431 21327 2437
rect 21269 2428 21281 2431
rect 21232 2400 21281 2428
rect 21232 2388 21238 2400
rect 21269 2397 21281 2400
rect 21315 2397 21327 2431
rect 21818 2428 21824 2440
rect 21779 2400 21824 2428
rect 21269 2391 21327 2397
rect 21818 2388 21824 2400
rect 21876 2388 21882 2440
rect 22002 2428 22008 2440
rect 21963 2400 22008 2428
rect 22002 2388 22008 2400
rect 22060 2388 22066 2440
rect 22094 2388 22100 2440
rect 22152 2428 22158 2440
rect 22848 2437 22876 2468
rect 23566 2456 23572 2468
rect 23624 2456 23630 2508
rect 27709 2499 27767 2505
rect 27709 2465 27721 2499
rect 27755 2496 27767 2499
rect 29730 2496 29736 2508
rect 27755 2468 29736 2496
rect 27755 2465 27767 2468
rect 27709 2459 27767 2465
rect 29730 2456 29736 2468
rect 29788 2456 29794 2508
rect 30009 2499 30067 2505
rect 30009 2465 30021 2499
rect 30055 2496 30067 2499
rect 30926 2496 30932 2508
rect 30055 2468 30932 2496
rect 30055 2465 30067 2468
rect 30009 2459 30067 2465
rect 30926 2456 30932 2468
rect 30984 2456 30990 2508
rect 22649 2431 22707 2437
rect 22649 2428 22661 2431
rect 22152 2400 22661 2428
rect 22152 2388 22158 2400
rect 22649 2397 22661 2400
rect 22695 2397 22707 2431
rect 22649 2391 22707 2397
rect 22833 2431 22891 2437
rect 22833 2397 22845 2431
rect 22879 2397 22891 2431
rect 22833 2391 22891 2397
rect 22925 2431 22983 2437
rect 22925 2397 22937 2431
rect 22971 2397 22983 2431
rect 22925 2391 22983 2397
rect 23753 2431 23811 2437
rect 23753 2397 23765 2431
rect 23799 2428 23811 2431
rect 24394 2428 24400 2440
rect 23799 2400 24400 2428
rect 23799 2397 23811 2400
rect 23753 2391 23811 2397
rect 20898 2360 20904 2372
rect 13372 2332 17724 2360
rect 19904 2332 20904 2360
rect 6788 2264 8984 2292
rect 6788 2252 6794 2264
rect 9214 2252 9220 2304
rect 9272 2252 9278 2304
rect 13372 2301 13400 2332
rect 17696 2304 17724 2332
rect 20898 2320 20904 2332
rect 20956 2320 20962 2372
rect 22940 2360 22968 2391
rect 24394 2388 24400 2400
rect 24452 2388 24458 2440
rect 24670 2428 24676 2440
rect 24631 2400 24676 2428
rect 24670 2388 24676 2400
rect 24728 2388 24734 2440
rect 26421 2431 26479 2437
rect 26421 2397 26433 2431
rect 26467 2397 26479 2431
rect 26970 2428 26976 2440
rect 26931 2400 26976 2428
rect 26421 2391 26479 2397
rect 21008 2332 22968 2360
rect 26436 2360 26464 2391
rect 26970 2388 26976 2400
rect 27028 2388 27034 2440
rect 28353 2431 28411 2437
rect 28353 2397 28365 2431
rect 28399 2428 28411 2431
rect 30190 2428 30196 2440
rect 28399 2400 30196 2428
rect 28399 2397 28411 2400
rect 28353 2391 28411 2397
rect 30190 2388 30196 2400
rect 30248 2388 30254 2440
rect 30374 2388 30380 2440
rect 30432 2428 30438 2440
rect 31312 2437 31340 2604
rect 33502 2592 33508 2604
rect 33560 2592 33566 2644
rect 33962 2632 33968 2644
rect 33923 2604 33968 2632
rect 33962 2592 33968 2604
rect 34020 2592 34026 2644
rect 35342 2632 35348 2644
rect 35303 2604 35348 2632
rect 35342 2592 35348 2604
rect 35400 2592 35406 2644
rect 36725 2635 36783 2641
rect 36725 2601 36737 2635
rect 36771 2632 36783 2635
rect 36906 2632 36912 2644
rect 36771 2604 36912 2632
rect 36771 2601 36783 2604
rect 36725 2595 36783 2601
rect 36906 2592 36912 2604
rect 36964 2592 36970 2644
rect 37090 2592 37096 2644
rect 37148 2632 37154 2644
rect 37148 2604 41276 2632
rect 37148 2592 37154 2604
rect 32030 2524 32036 2576
rect 32088 2564 32094 2576
rect 32125 2567 32183 2573
rect 32125 2564 32137 2567
rect 32088 2536 32137 2564
rect 32088 2524 32094 2536
rect 32125 2533 32137 2536
rect 32171 2533 32183 2567
rect 32125 2527 32183 2533
rect 32858 2524 32864 2576
rect 32916 2564 32922 2576
rect 32916 2536 35894 2564
rect 32916 2524 32922 2536
rect 31478 2456 31484 2508
rect 31536 2496 31542 2508
rect 34701 2499 34759 2505
rect 34701 2496 34713 2499
rect 31536 2468 34713 2496
rect 31536 2456 31542 2468
rect 34701 2465 34713 2468
rect 34747 2465 34759 2499
rect 35866 2496 35894 2536
rect 36446 2524 36452 2576
rect 36504 2564 36510 2576
rect 41141 2567 41199 2573
rect 41141 2564 41153 2567
rect 36504 2536 41153 2564
rect 36504 2524 36510 2536
rect 41141 2533 41153 2536
rect 41187 2533 41199 2567
rect 41248 2564 41276 2604
rect 43714 2592 43720 2644
rect 43772 2632 43778 2644
rect 43772 2604 46520 2632
rect 43772 2592 43778 2604
rect 42429 2567 42487 2573
rect 42429 2564 42441 2567
rect 41248 2536 42441 2564
rect 41141 2527 41199 2533
rect 42429 2533 42441 2536
rect 42475 2533 42487 2567
rect 46293 2567 46351 2573
rect 46293 2564 46305 2567
rect 42429 2527 42487 2533
rect 42536 2536 46305 2564
rect 35989 2499 36047 2505
rect 35989 2496 36001 2499
rect 35866 2468 36001 2496
rect 34701 2459 34759 2465
rect 35989 2465 36001 2468
rect 36035 2465 36047 2499
rect 38565 2499 38623 2505
rect 38565 2496 38577 2499
rect 35989 2459 36047 2465
rect 37200 2468 38577 2496
rect 30469 2431 30527 2437
rect 30469 2428 30481 2431
rect 30432 2400 30481 2428
rect 30432 2388 30438 2400
rect 30469 2397 30481 2400
rect 30515 2397 30527 2431
rect 30469 2391 30527 2397
rect 31297 2431 31355 2437
rect 31297 2397 31309 2431
rect 31343 2397 31355 2431
rect 31570 2428 31576 2440
rect 31531 2400 31576 2428
rect 31297 2391 31355 2397
rect 31570 2388 31576 2400
rect 31628 2388 31634 2440
rect 33226 2428 33232 2440
rect 33187 2400 33232 2428
rect 33226 2388 33232 2400
rect 33284 2388 33290 2440
rect 33505 2431 33563 2437
rect 33505 2397 33517 2431
rect 33551 2428 33563 2431
rect 33594 2428 33600 2440
rect 33551 2400 33600 2428
rect 33551 2397 33563 2400
rect 33505 2391 33563 2397
rect 33594 2388 33600 2400
rect 33652 2388 33658 2440
rect 33686 2388 33692 2440
rect 33744 2428 33750 2440
rect 37200 2428 37228 2468
rect 38565 2465 38577 2468
rect 38611 2465 38623 2499
rect 39206 2496 39212 2508
rect 39167 2468 39212 2496
rect 38565 2459 38623 2465
rect 39206 2456 39212 2468
rect 39264 2456 39270 2508
rect 39482 2456 39488 2508
rect 39540 2496 39546 2508
rect 42536 2496 42564 2536
rect 46293 2533 46305 2536
rect 46339 2533 46351 2567
rect 46492 2564 46520 2604
rect 46566 2592 46572 2644
rect 46624 2632 46630 2644
rect 47029 2635 47087 2641
rect 47029 2632 47041 2635
rect 46624 2604 47041 2632
rect 46624 2592 46630 2604
rect 47029 2601 47041 2604
rect 47075 2632 47087 2635
rect 49510 2632 49516 2644
rect 47075 2604 49516 2632
rect 47075 2601 47087 2604
rect 47029 2595 47087 2601
rect 49510 2592 49516 2604
rect 49568 2632 49574 2644
rect 57241 2635 57299 2641
rect 57241 2632 57253 2635
rect 49568 2604 57253 2632
rect 49568 2592 49574 2604
rect 57241 2601 57253 2604
rect 57287 2632 57299 2635
rect 57882 2632 57888 2644
rect 57287 2604 57888 2632
rect 57287 2601 57299 2604
rect 57241 2595 57299 2601
rect 57882 2592 57888 2604
rect 57940 2592 57946 2644
rect 50338 2564 50344 2576
rect 46492 2536 50344 2564
rect 46293 2527 46351 2533
rect 50338 2524 50344 2536
rect 50396 2524 50402 2576
rect 50890 2524 50896 2576
rect 50948 2564 50954 2576
rect 56597 2567 56655 2573
rect 56597 2564 56609 2567
rect 50948 2536 56609 2564
rect 50948 2524 50954 2536
rect 56597 2533 56609 2536
rect 56643 2533 56655 2567
rect 56597 2527 56655 2533
rect 39540 2468 42564 2496
rect 39540 2456 39546 2468
rect 42702 2456 42708 2508
rect 42760 2496 42766 2508
rect 47581 2499 47639 2505
rect 47581 2496 47593 2499
rect 42760 2468 47593 2496
rect 42760 2456 42766 2468
rect 47581 2465 47593 2468
rect 47627 2465 47639 2499
rect 52086 2496 52092 2508
rect 52047 2468 52092 2496
rect 47581 2459 47639 2465
rect 52086 2456 52092 2468
rect 52144 2456 52150 2508
rect 55953 2499 56011 2505
rect 55953 2496 55965 2499
rect 52196 2468 55965 2496
rect 33744 2400 37228 2428
rect 37277 2431 37335 2437
rect 33744 2388 33750 2400
rect 37277 2397 37289 2431
rect 37323 2397 37335 2431
rect 37277 2391 37335 2397
rect 37921 2431 37979 2437
rect 37921 2397 37933 2431
rect 37967 2397 37979 2431
rect 39850 2428 39856 2440
rect 39811 2400 39856 2428
rect 37921 2391 37979 2397
rect 28994 2360 29000 2372
rect 26436 2332 29000 2360
rect 13357 2295 13415 2301
rect 13357 2261 13369 2295
rect 13403 2261 13415 2295
rect 14550 2292 14556 2304
rect 14511 2264 14556 2292
rect 13357 2255 13415 2261
rect 14550 2252 14556 2264
rect 14608 2252 14614 2304
rect 15286 2292 15292 2304
rect 15247 2264 15292 2292
rect 15286 2252 15292 2264
rect 15344 2252 15350 2304
rect 16022 2292 16028 2304
rect 15983 2264 16028 2292
rect 16022 2252 16028 2264
rect 16080 2252 16086 2304
rect 17678 2252 17684 2304
rect 17736 2252 17742 2304
rect 19518 2292 19524 2304
rect 19431 2264 19524 2292
rect 19518 2252 19524 2264
rect 19576 2292 19582 2304
rect 21008 2292 21036 2332
rect 28994 2320 29000 2332
rect 29052 2320 29058 2372
rect 31481 2363 31539 2369
rect 31481 2329 31493 2363
rect 31527 2360 31539 2363
rect 33244 2360 33272 2388
rect 31527 2332 33272 2360
rect 31527 2329 31539 2332
rect 31481 2323 31539 2329
rect 33318 2320 33324 2372
rect 33376 2360 33382 2372
rect 37292 2360 37320 2391
rect 33376 2332 37320 2360
rect 33376 2320 33382 2332
rect 19576 2264 21036 2292
rect 21085 2295 21143 2301
rect 19576 2252 19582 2264
rect 21085 2261 21097 2295
rect 21131 2292 21143 2295
rect 21818 2292 21824 2304
rect 21131 2264 21824 2292
rect 21131 2261 21143 2264
rect 21085 2255 21143 2261
rect 21818 2252 21824 2264
rect 21876 2252 21882 2304
rect 22189 2295 22247 2301
rect 22189 2261 22201 2295
rect 22235 2292 22247 2295
rect 22830 2292 22836 2304
rect 22235 2264 22836 2292
rect 22235 2261 22247 2264
rect 22189 2255 22247 2261
rect 22830 2252 22836 2264
rect 22888 2252 22894 2304
rect 22922 2252 22928 2304
rect 22980 2292 22986 2304
rect 23569 2295 23627 2301
rect 23569 2292 23581 2295
rect 22980 2264 23581 2292
rect 22980 2252 22986 2264
rect 23569 2261 23581 2264
rect 23615 2261 23627 2295
rect 23569 2255 23627 2261
rect 26970 2252 26976 2304
rect 27028 2292 27034 2304
rect 31294 2292 31300 2304
rect 27028 2264 31300 2292
rect 27028 2252 27034 2264
rect 31294 2252 31300 2264
rect 31352 2252 31358 2304
rect 32582 2252 32588 2304
rect 32640 2292 32646 2304
rect 37936 2292 37964 2391
rect 39850 2388 39856 2400
rect 39908 2388 39914 2440
rect 40494 2428 40500 2440
rect 40455 2400 40500 2428
rect 40494 2388 40500 2400
rect 40552 2388 40558 2440
rect 43070 2428 43076 2440
rect 43031 2400 43076 2428
rect 43070 2388 43076 2400
rect 43128 2388 43134 2440
rect 43714 2428 43720 2440
rect 43675 2400 43720 2428
rect 43714 2388 43720 2400
rect 43772 2388 43778 2440
rect 43898 2388 43904 2440
rect 43956 2428 43962 2440
rect 44361 2431 44419 2437
rect 44361 2428 44373 2431
rect 43956 2400 44373 2428
rect 43956 2388 43962 2400
rect 44361 2397 44373 2400
rect 44407 2397 44419 2431
rect 44361 2391 44419 2397
rect 45005 2431 45063 2437
rect 45005 2397 45017 2431
rect 45051 2397 45063 2431
rect 45649 2431 45707 2437
rect 45649 2428 45661 2431
rect 45005 2391 45063 2397
rect 45526 2400 45661 2428
rect 38010 2320 38016 2372
rect 38068 2360 38074 2372
rect 45020 2360 45048 2391
rect 38068 2332 45048 2360
rect 38068 2320 38074 2332
rect 45094 2320 45100 2372
rect 45152 2360 45158 2372
rect 45526 2360 45554 2400
rect 45649 2397 45661 2400
rect 45695 2397 45707 2431
rect 48222 2428 48228 2440
rect 48183 2400 48228 2428
rect 45649 2391 45707 2397
rect 48222 2388 48228 2400
rect 48280 2388 48286 2440
rect 48866 2428 48872 2440
rect 48827 2400 48872 2428
rect 48866 2388 48872 2400
rect 48924 2388 48930 2440
rect 49510 2428 49516 2440
rect 49471 2400 49516 2428
rect 49510 2388 49516 2400
rect 49568 2388 49574 2440
rect 50154 2428 50160 2440
rect 50115 2400 50160 2428
rect 50154 2388 50160 2400
rect 50212 2388 50218 2440
rect 50798 2428 50804 2440
rect 50759 2400 50804 2428
rect 50798 2388 50804 2400
rect 50856 2388 50862 2440
rect 51442 2428 51448 2440
rect 51403 2400 51448 2428
rect 51442 2388 51448 2400
rect 51500 2388 51506 2440
rect 52196 2428 52224 2468
rect 55953 2465 55965 2468
rect 55999 2465 56011 2499
rect 55953 2459 56011 2465
rect 51552 2400 52224 2428
rect 45152 2332 45554 2360
rect 45152 2320 45158 2332
rect 49418 2320 49424 2372
rect 49476 2360 49482 2372
rect 51552 2360 51580 2400
rect 52270 2388 52276 2440
rect 52328 2428 52334 2440
rect 52733 2431 52791 2437
rect 52733 2428 52745 2431
rect 52328 2400 52745 2428
rect 52328 2388 52334 2400
rect 52733 2397 52745 2400
rect 52779 2397 52791 2431
rect 53374 2428 53380 2440
rect 53335 2400 53380 2428
rect 52733 2391 52791 2397
rect 53374 2388 53380 2400
rect 53432 2388 53438 2440
rect 54018 2428 54024 2440
rect 53979 2400 54024 2428
rect 54018 2388 54024 2400
rect 54076 2388 54082 2440
rect 55309 2431 55367 2437
rect 55309 2428 55321 2431
rect 55186 2400 55321 2428
rect 55186 2360 55214 2400
rect 55309 2397 55321 2400
rect 55355 2397 55367 2431
rect 55309 2391 55367 2397
rect 49476 2332 51580 2360
rect 52288 2332 55214 2360
rect 49476 2320 49482 2332
rect 41782 2292 41788 2304
rect 32640 2264 37964 2292
rect 41743 2264 41788 2292
rect 32640 2252 32646 2264
rect 41782 2252 41788 2264
rect 41840 2252 41846 2304
rect 46750 2252 46756 2304
rect 46808 2292 46814 2304
rect 49050 2292 49056 2304
rect 46808 2264 49056 2292
rect 46808 2252 46814 2264
rect 49050 2252 49056 2264
rect 49108 2252 49114 2304
rect 49142 2252 49148 2304
rect 49200 2292 49206 2304
rect 52288 2292 52316 2332
rect 54662 2292 54668 2304
rect 49200 2264 52316 2292
rect 54623 2264 54668 2292
rect 49200 2252 49206 2264
rect 54662 2252 54668 2264
rect 54720 2252 54726 2304
rect 57882 2292 57888 2304
rect 57843 2264 57888 2292
rect 57882 2252 57888 2264
rect 57940 2252 57946 2304
rect 1104 2202 58880 2224
rect 1104 2150 15398 2202
rect 15450 2150 15462 2202
rect 15514 2150 15526 2202
rect 15578 2150 15590 2202
rect 15642 2150 15654 2202
rect 15706 2150 29846 2202
rect 29898 2150 29910 2202
rect 29962 2150 29974 2202
rect 30026 2150 30038 2202
rect 30090 2150 30102 2202
rect 30154 2150 44294 2202
rect 44346 2150 44358 2202
rect 44410 2150 44422 2202
rect 44474 2150 44486 2202
rect 44538 2150 44550 2202
rect 44602 2150 58880 2202
rect 1104 2128 58880 2150
rect 6914 2048 6920 2100
rect 6972 2088 6978 2100
rect 9214 2088 9220 2100
rect 6972 2060 9220 2088
rect 6972 2048 6978 2060
rect 9214 2048 9220 2060
rect 9272 2048 9278 2100
rect 20070 2048 20076 2100
rect 20128 2088 20134 2100
rect 20128 2060 21036 2088
rect 20128 2048 20134 2060
rect 2130 1980 2136 2032
rect 2188 2020 2194 2032
rect 14366 2020 14372 2032
rect 2188 1992 14372 2020
rect 2188 1980 2194 1992
rect 14366 1980 14372 1992
rect 14424 1980 14430 2032
rect 15286 1980 15292 2032
rect 15344 2020 15350 2032
rect 20438 2020 20444 2032
rect 15344 1992 20444 2020
rect 15344 1980 15350 1992
rect 20438 1980 20444 1992
rect 20496 1980 20502 2032
rect 21008 2020 21036 2060
rect 21082 2048 21088 2100
rect 21140 2088 21146 2100
rect 24670 2088 24676 2100
rect 21140 2060 24676 2088
rect 21140 2048 21146 2060
rect 24670 2048 24676 2060
rect 24728 2048 24734 2100
rect 32030 2048 32036 2100
rect 32088 2088 32094 2100
rect 33318 2088 33324 2100
rect 32088 2060 33324 2088
rect 32088 2048 32094 2060
rect 33318 2048 33324 2060
rect 33376 2048 33382 2100
rect 35066 2048 35072 2100
rect 35124 2088 35130 2100
rect 40494 2088 40500 2100
rect 35124 2060 40500 2088
rect 35124 2048 35130 2060
rect 40494 2048 40500 2060
rect 40552 2048 40558 2100
rect 40862 2048 40868 2100
rect 40920 2088 40926 2100
rect 42702 2088 42708 2100
rect 40920 2060 42708 2088
rect 40920 2048 40926 2060
rect 42702 2048 42708 2060
rect 42760 2048 42766 2100
rect 44726 2048 44732 2100
rect 44784 2088 44790 2100
rect 45186 2088 45192 2100
rect 44784 2060 45192 2088
rect 44784 2048 44790 2060
rect 45186 2048 45192 2060
rect 45244 2048 45250 2100
rect 45278 2048 45284 2100
rect 45336 2088 45342 2100
rect 53374 2088 53380 2100
rect 45336 2060 53380 2088
rect 45336 2048 45342 2060
rect 53374 2048 53380 2060
rect 53432 2048 53438 2100
rect 26234 2020 26240 2032
rect 21008 1992 26240 2020
rect 26234 1980 26240 1992
rect 26292 1980 26298 2032
rect 33226 1980 33232 2032
rect 33284 2020 33290 2032
rect 33284 1992 36676 2020
rect 33284 1980 33290 1992
rect 6546 1912 6552 1964
rect 6604 1952 6610 1964
rect 8294 1952 8300 1964
rect 6604 1924 8300 1952
rect 6604 1912 6610 1924
rect 8294 1912 8300 1924
rect 8352 1912 8358 1964
rect 8754 1912 8760 1964
rect 8812 1952 8818 1964
rect 9490 1952 9496 1964
rect 8812 1924 9496 1952
rect 8812 1912 8818 1924
rect 9490 1912 9496 1924
rect 9548 1912 9554 1964
rect 14458 1952 14464 1964
rect 12406 1924 14464 1952
rect 2774 1844 2780 1896
rect 2832 1884 2838 1896
rect 8110 1884 8116 1896
rect 2832 1856 8116 1884
rect 2832 1844 2838 1856
rect 8110 1844 8116 1856
rect 8168 1844 8174 1896
rect 3510 1776 3516 1828
rect 3568 1816 3574 1828
rect 12406 1816 12434 1924
rect 14458 1912 14464 1924
rect 14516 1912 14522 1964
rect 14550 1912 14556 1964
rect 14608 1952 14614 1964
rect 19610 1952 19616 1964
rect 14608 1924 19616 1952
rect 14608 1912 14614 1924
rect 19610 1912 19616 1924
rect 19668 1912 19674 1964
rect 34790 1912 34796 1964
rect 34848 1952 34854 1964
rect 36648 1952 36676 1992
rect 36722 1980 36728 2032
rect 36780 2020 36786 2032
rect 43070 2020 43076 2032
rect 36780 1992 43076 2020
rect 36780 1980 36786 1992
rect 43070 1980 43076 1992
rect 43128 1980 43134 2032
rect 44450 1980 44456 2032
rect 44508 2020 44514 2032
rect 51442 2020 51448 2032
rect 44508 1992 51448 2020
rect 44508 1980 44514 1992
rect 51442 1980 51448 1992
rect 51500 1980 51506 2032
rect 53282 1980 53288 2032
rect 53340 2020 53346 2032
rect 57882 2020 57888 2032
rect 53340 1992 57888 2020
rect 53340 1980 53346 1992
rect 57882 1980 57888 1992
rect 57940 1980 57946 2032
rect 37642 1952 37648 1964
rect 34848 1924 35940 1952
rect 36648 1924 37648 1952
rect 34848 1912 34854 1924
rect 13538 1844 13544 1896
rect 13596 1884 13602 1896
rect 26142 1884 26148 1896
rect 13596 1856 26148 1884
rect 13596 1844 13602 1856
rect 26142 1844 26148 1856
rect 26200 1844 26206 1896
rect 3568 1788 12434 1816
rect 3568 1776 3574 1788
rect 14918 1776 14924 1828
rect 14976 1816 14982 1828
rect 15286 1816 15292 1828
rect 14976 1788 15292 1816
rect 14976 1776 14982 1788
rect 15286 1776 15292 1788
rect 15344 1776 15350 1828
rect 19518 1816 19524 1828
rect 16546 1788 19524 1816
rect 5166 1708 5172 1760
rect 5224 1748 5230 1760
rect 7098 1748 7104 1760
rect 5224 1720 7104 1748
rect 5224 1708 5230 1720
rect 7098 1708 7104 1720
rect 7156 1708 7162 1760
rect 7834 1708 7840 1760
rect 7892 1748 7898 1760
rect 8754 1748 8760 1760
rect 7892 1720 8760 1748
rect 7892 1708 7898 1720
rect 8754 1708 8760 1720
rect 8812 1708 8818 1760
rect 10778 1708 10784 1760
rect 10836 1748 10842 1760
rect 11606 1748 11612 1760
rect 10836 1720 11612 1748
rect 10836 1708 10842 1720
rect 11606 1708 11612 1720
rect 11664 1708 11670 1760
rect 14090 1748 14096 1760
rect 12406 1720 14096 1748
rect 3142 1640 3148 1692
rect 3200 1680 3206 1692
rect 12406 1680 12434 1720
rect 14090 1708 14096 1720
rect 14148 1708 14154 1760
rect 14642 1708 14648 1760
rect 14700 1748 14706 1760
rect 16546 1748 16574 1788
rect 19518 1776 19524 1788
rect 19576 1776 19582 1828
rect 35912 1816 35940 1924
rect 37642 1912 37648 1924
rect 37700 1912 37706 1964
rect 41414 1912 41420 1964
rect 41472 1952 41478 1964
rect 48222 1952 48228 1964
rect 41472 1924 48228 1952
rect 41472 1912 41478 1924
rect 48222 1912 48228 1924
rect 48280 1912 48286 1964
rect 50338 1912 50344 1964
rect 50396 1952 50402 1964
rect 56410 1952 56416 1964
rect 50396 1924 56416 1952
rect 50396 1912 50402 1924
rect 56410 1912 56416 1924
rect 56468 1912 56474 1964
rect 38654 1844 38660 1896
rect 38712 1884 38718 1896
rect 45094 1884 45100 1896
rect 38712 1856 45100 1884
rect 38712 1844 38718 1856
rect 45094 1844 45100 1856
rect 45152 1844 45158 1896
rect 46106 1844 46112 1896
rect 46164 1884 46170 1896
rect 54018 1884 54024 1896
rect 46164 1856 54024 1884
rect 46164 1844 46170 1856
rect 54018 1844 54024 1856
rect 54076 1844 54082 1896
rect 39850 1816 39856 1828
rect 35912 1788 39856 1816
rect 39850 1776 39856 1788
rect 39908 1776 39914 1828
rect 43622 1776 43628 1828
rect 43680 1816 43686 1828
rect 50798 1816 50804 1828
rect 43680 1788 50804 1816
rect 43680 1776 43686 1788
rect 50798 1776 50804 1788
rect 50856 1776 50862 1828
rect 14700 1720 16574 1748
rect 14700 1708 14706 1720
rect 49050 1708 49056 1760
rect 49108 1748 49114 1760
rect 53834 1748 53840 1760
rect 49108 1720 53840 1748
rect 49108 1708 49114 1720
rect 53834 1708 53840 1720
rect 53892 1748 53898 1760
rect 54662 1748 54668 1760
rect 53892 1720 54668 1748
rect 53892 1708 53898 1720
rect 54662 1708 54668 1720
rect 54720 1708 54726 1760
rect 3200 1652 12434 1680
rect 3200 1640 3206 1652
rect 18138 1640 18144 1692
rect 18196 1680 18202 1692
rect 31386 1680 31392 1692
rect 18196 1652 31392 1680
rect 18196 1640 18202 1652
rect 31386 1640 31392 1652
rect 31444 1640 31450 1692
rect 44174 1640 44180 1692
rect 44232 1680 44238 1692
rect 44818 1680 44824 1692
rect 44232 1652 44824 1680
rect 44232 1640 44238 1652
rect 44818 1640 44824 1652
rect 44876 1640 44882 1692
rect 46658 1640 46664 1692
rect 46716 1680 46722 1692
rect 52270 1680 52276 1692
rect 46716 1652 52276 1680
rect 46716 1640 46722 1652
rect 52270 1640 52276 1652
rect 52328 1640 52334 1692
rect 19242 1572 19248 1624
rect 19300 1612 19306 1624
rect 27706 1612 27712 1624
rect 19300 1584 27712 1612
rect 19300 1572 19306 1584
rect 27706 1572 27712 1584
rect 27764 1572 27770 1624
rect 7466 1504 7472 1556
rect 7524 1504 7530 1556
rect 8202 1544 8208 1556
rect 8036 1516 8208 1544
rect 7484 1476 7512 1504
rect 8036 1488 8064 1516
rect 8202 1504 8208 1516
rect 8260 1504 8266 1556
rect 9674 1504 9680 1556
rect 9732 1544 9738 1556
rect 10502 1544 10508 1556
rect 9732 1516 10508 1544
rect 9732 1504 9738 1516
rect 10502 1504 10508 1516
rect 10560 1504 10566 1556
rect 10594 1504 10600 1556
rect 10652 1504 10658 1556
rect 39758 1504 39764 1556
rect 39816 1544 39822 1556
rect 45646 1544 45652 1556
rect 39816 1516 45652 1544
rect 39816 1504 39822 1516
rect 45646 1504 45652 1516
rect 45704 1504 45710 1556
rect 7484 1448 7604 1476
rect 7006 1368 7012 1420
rect 7064 1408 7070 1420
rect 7466 1408 7472 1420
rect 7064 1380 7472 1408
rect 7064 1368 7070 1380
rect 7466 1368 7472 1380
rect 7524 1368 7530 1420
rect 7576 1408 7604 1448
rect 8018 1436 8024 1488
rect 8076 1436 8082 1488
rect 8846 1436 8852 1488
rect 8904 1476 8910 1488
rect 9582 1476 9588 1488
rect 8904 1448 9588 1476
rect 8904 1436 8910 1448
rect 9582 1436 9588 1448
rect 9640 1436 9646 1488
rect 10612 1476 10640 1504
rect 10428 1448 10640 1476
rect 7576 1380 7788 1408
rect 7760 1340 7788 1380
rect 10428 1352 10456 1448
rect 16022 1436 16028 1488
rect 16080 1476 16086 1488
rect 20162 1476 20168 1488
rect 16080 1448 20168 1476
rect 16080 1436 16086 1448
rect 20162 1436 20168 1448
rect 20220 1436 20226 1488
rect 37274 1436 37280 1488
rect 37332 1476 37338 1488
rect 38286 1476 38292 1488
rect 37332 1448 38292 1476
rect 37332 1436 37338 1448
rect 38286 1436 38292 1448
rect 38344 1436 38350 1488
rect 39206 1436 39212 1488
rect 39264 1476 39270 1488
rect 44910 1476 44916 1488
rect 39264 1448 44916 1476
rect 39264 1436 39270 1448
rect 44910 1436 44916 1448
rect 44968 1436 44974 1488
rect 49970 1436 49976 1488
rect 50028 1476 50034 1488
rect 54754 1476 54760 1488
rect 50028 1448 54760 1476
rect 50028 1436 50034 1448
rect 54754 1436 54760 1448
rect 54812 1436 54818 1488
rect 10962 1408 10968 1420
rect 10520 1380 10968 1408
rect 10520 1352 10548 1380
rect 10962 1368 10968 1380
rect 11020 1368 11026 1420
rect 13446 1368 13452 1420
rect 13504 1408 13510 1420
rect 17126 1408 17132 1420
rect 13504 1380 17132 1408
rect 13504 1368 13510 1380
rect 17126 1368 17132 1380
rect 17184 1368 17190 1420
rect 24026 1368 24032 1420
rect 24084 1408 24090 1420
rect 29454 1408 29460 1420
rect 24084 1380 29460 1408
rect 24084 1368 24090 1380
rect 29454 1368 29460 1380
rect 29512 1368 29518 1420
rect 36170 1368 36176 1420
rect 36228 1408 36234 1420
rect 37090 1408 37096 1420
rect 36228 1380 37096 1408
rect 36228 1368 36234 1380
rect 37090 1368 37096 1380
rect 37148 1368 37154 1420
rect 41138 1368 41144 1420
rect 41196 1408 41202 1420
rect 46842 1408 46848 1420
rect 41196 1380 46848 1408
rect 41196 1368 41202 1380
rect 46842 1368 46848 1380
rect 46900 1368 46906 1420
rect 7926 1340 7932 1352
rect 7760 1312 7932 1340
rect 7926 1300 7932 1312
rect 7984 1300 7990 1352
rect 10410 1300 10416 1352
rect 10468 1300 10474 1352
rect 10502 1300 10508 1352
rect 10560 1300 10566 1352
rect 20530 1300 20536 1352
rect 20588 1340 20594 1352
rect 53282 1340 53288 1352
rect 20588 1312 53288 1340
rect 20588 1300 20594 1312
rect 53282 1300 53288 1312
rect 53340 1300 53346 1352
rect 7282 1232 7288 1284
rect 7340 1272 7346 1284
rect 7834 1272 7840 1284
rect 7340 1244 7840 1272
rect 7340 1232 7346 1244
rect 7834 1232 7840 1244
rect 7892 1232 7898 1284
rect 20254 1232 20260 1284
rect 20312 1272 20318 1284
rect 52638 1272 52644 1284
rect 20312 1244 52644 1272
rect 20312 1232 20318 1244
rect 52638 1232 52644 1244
rect 52696 1232 52702 1284
rect 6086 1164 6092 1216
rect 6144 1204 6150 1216
rect 8570 1204 8576 1216
rect 6144 1176 8576 1204
rect 6144 1164 6150 1176
rect 8570 1164 8576 1176
rect 8628 1164 8634 1216
rect 33778 1204 33784 1216
rect 9646 1176 33784 1204
rect 5902 1096 5908 1148
rect 5960 1136 5966 1148
rect 9646 1136 9674 1176
rect 33778 1164 33784 1176
rect 33836 1164 33842 1216
rect 38930 1164 38936 1216
rect 38988 1204 38994 1216
rect 43714 1204 43720 1216
rect 38988 1176 43720 1204
rect 38988 1164 38994 1176
rect 43714 1164 43720 1176
rect 43772 1164 43778 1216
rect 5960 1108 9674 1136
rect 5960 1096 5966 1108
rect 10410 1096 10416 1148
rect 10468 1136 10474 1148
rect 25314 1136 25320 1148
rect 10468 1108 25320 1136
rect 10468 1096 10474 1108
rect 25314 1096 25320 1108
rect 25372 1096 25378 1148
rect 26878 1096 26884 1148
rect 26936 1136 26942 1148
rect 40126 1136 40132 1148
rect 26936 1108 40132 1136
rect 26936 1096 26942 1108
rect 40126 1096 40132 1108
rect 40184 1096 40190 1148
rect 4890 1028 4896 1080
rect 4948 1068 4954 1080
rect 8386 1068 8392 1080
rect 4948 1040 8392 1068
rect 4948 1028 4954 1040
rect 8386 1028 8392 1040
rect 8444 1028 8450 1080
rect 18874 1028 18880 1080
rect 18932 1068 18938 1080
rect 35434 1068 35440 1080
rect 18932 1040 35440 1068
rect 18932 1028 18938 1040
rect 35434 1028 35440 1040
rect 35492 1028 35498 1080
rect 4522 960 4528 1012
rect 4580 1000 4586 1012
rect 8202 1000 8208 1012
rect 4580 972 8208 1000
rect 4580 960 4586 972
rect 8202 960 8208 972
rect 8260 960 8266 1012
rect 14826 960 14832 1012
rect 14884 1000 14890 1012
rect 29638 1000 29644 1012
rect 14884 972 29644 1000
rect 14884 960 14890 972
rect 29638 960 29644 972
rect 29696 960 29702 1012
rect 13170 892 13176 944
rect 13228 932 13234 944
rect 26326 932 26332 944
rect 13228 904 26332 932
rect 13228 892 13234 904
rect 26326 892 26332 904
rect 26384 892 26390 944
rect 26418 892 26424 944
rect 26476 892 26482 944
rect 26602 892 26608 944
rect 26660 892 26666 944
rect 3234 756 3240 808
rect 3292 796 3298 808
rect 3292 768 22508 796
rect 3292 756 3298 768
rect 7190 688 7196 740
rect 7248 728 7254 740
rect 7248 700 16574 728
rect 7248 688 7254 700
rect 16546 524 16574 700
rect 22480 592 22508 768
rect 26436 728 26464 892
rect 26206 700 26464 728
rect 26206 592 26234 700
rect 22480 564 26234 592
rect 26620 524 26648 892
rect 16546 496 26648 524
<< via1 >>
rect 15398 17382 15450 17434
rect 15462 17382 15514 17434
rect 15526 17382 15578 17434
rect 15590 17382 15642 17434
rect 15654 17382 15706 17434
rect 29846 17382 29898 17434
rect 29910 17382 29962 17434
rect 29974 17382 30026 17434
rect 30038 17382 30090 17434
rect 30102 17382 30154 17434
rect 44294 17382 44346 17434
rect 44358 17382 44410 17434
rect 44422 17382 44474 17434
rect 44486 17382 44538 17434
rect 44550 17382 44602 17434
rect 4436 17144 4488 17196
rect 4896 17144 4948 17196
rect 5816 17187 5868 17196
rect 5816 17153 5825 17187
rect 5825 17153 5859 17187
rect 5859 17153 5868 17187
rect 5816 17144 5868 17153
rect 7196 17144 7248 17196
rect 7656 17144 7708 17196
rect 8576 17144 8628 17196
rect 9036 17144 9088 17196
rect 9956 17144 10008 17196
rect 10416 17144 10468 17196
rect 11796 17144 11848 17196
rect 12716 17144 12768 17196
rect 13176 17144 13228 17196
rect 14556 17144 14608 17196
rect 15292 17144 15344 17196
rect 15936 17187 15988 17196
rect 15936 17153 15945 17187
rect 15945 17153 15979 17187
rect 15979 17153 15988 17187
rect 15936 17144 15988 17153
rect 17316 17144 17368 17196
rect 18236 17144 18288 17196
rect 18696 17187 18748 17196
rect 18696 17153 18705 17187
rect 18705 17153 18739 17187
rect 18739 17153 18748 17187
rect 18696 17144 18748 17153
rect 19616 17144 19668 17196
rect 20076 17144 20128 17196
rect 21456 17144 21508 17196
rect 22376 17144 22428 17196
rect 22836 17144 22888 17196
rect 23756 17144 23808 17196
rect 25136 17187 25188 17196
rect 25136 17153 25145 17187
rect 25145 17153 25179 17187
rect 25179 17153 25188 17187
rect 25136 17144 25188 17153
rect 25596 17187 25648 17196
rect 25596 17153 25605 17187
rect 25605 17153 25639 17187
rect 25639 17153 25648 17187
rect 25596 17144 25648 17153
rect 26516 17144 26568 17196
rect 27896 17144 27948 17196
rect 28356 17187 28408 17196
rect 28356 17153 28365 17187
rect 28365 17153 28399 17187
rect 28399 17153 28408 17187
rect 28356 17144 28408 17153
rect 29276 17144 29328 17196
rect 29736 17144 29788 17196
rect 30656 17144 30708 17196
rect 31116 17144 31168 17196
rect 32036 17144 32088 17196
rect 32496 17144 32548 17196
rect 33416 17144 33468 17196
rect 33876 17144 33928 17196
rect 34796 17144 34848 17196
rect 36636 17144 36688 17196
rect 37556 17144 37608 17196
rect 38016 17144 38068 17196
rect 38936 17144 38988 17196
rect 40316 17144 40368 17196
rect 40776 17144 40828 17196
rect 41696 17144 41748 17196
rect 43076 17144 43128 17196
rect 44640 17144 44692 17196
rect 45836 17144 45888 17196
rect 47216 17144 47268 17196
rect 47676 17144 47728 17196
rect 48596 17144 48648 17196
rect 49976 17144 50028 17196
rect 50436 17144 50488 17196
rect 51356 17144 51408 17196
rect 51816 17144 51868 17196
rect 53196 17144 53248 17196
rect 54576 17144 54628 17196
rect 55496 17144 55548 17196
rect 56048 17144 56100 17196
rect 35256 17076 35308 17128
rect 44916 17076 44968 17128
rect 42156 17008 42208 17060
rect 52736 17008 52788 17060
rect 8174 16838 8226 16890
rect 8238 16838 8290 16890
rect 8302 16838 8354 16890
rect 8366 16838 8418 16890
rect 8430 16838 8482 16890
rect 22622 16838 22674 16890
rect 22686 16838 22738 16890
rect 22750 16838 22802 16890
rect 22814 16838 22866 16890
rect 22878 16838 22930 16890
rect 37070 16838 37122 16890
rect 37134 16838 37186 16890
rect 37198 16838 37250 16890
rect 37262 16838 37314 16890
rect 37326 16838 37378 16890
rect 51518 16838 51570 16890
rect 51582 16838 51634 16890
rect 51646 16838 51698 16890
rect 51710 16838 51762 16890
rect 51774 16838 51826 16890
rect 6276 16736 6328 16788
rect 11336 16736 11388 16788
rect 14096 16736 14148 16788
rect 16856 16736 16908 16788
rect 20996 16736 21048 16788
rect 24216 16736 24268 16788
rect 26976 16736 27028 16788
rect 36176 16736 36228 16788
rect 39396 16736 39448 16788
rect 43536 16736 43588 16788
rect 46296 16736 46348 16788
rect 49056 16736 49108 16788
rect 54116 16736 54168 16788
rect 15398 16294 15450 16346
rect 15462 16294 15514 16346
rect 15526 16294 15578 16346
rect 15590 16294 15642 16346
rect 15654 16294 15706 16346
rect 29846 16294 29898 16346
rect 29910 16294 29962 16346
rect 29974 16294 30026 16346
rect 30038 16294 30090 16346
rect 30102 16294 30154 16346
rect 44294 16294 44346 16346
rect 44358 16294 44410 16346
rect 44422 16294 44474 16346
rect 44486 16294 44538 16346
rect 44550 16294 44602 16346
rect 8174 15750 8226 15802
rect 8238 15750 8290 15802
rect 8302 15750 8354 15802
rect 8366 15750 8418 15802
rect 8430 15750 8482 15802
rect 22622 15750 22674 15802
rect 22686 15750 22738 15802
rect 22750 15750 22802 15802
rect 22814 15750 22866 15802
rect 22878 15750 22930 15802
rect 37070 15750 37122 15802
rect 37134 15750 37186 15802
rect 37198 15750 37250 15802
rect 37262 15750 37314 15802
rect 37326 15750 37378 15802
rect 51518 15750 51570 15802
rect 51582 15750 51634 15802
rect 51646 15750 51698 15802
rect 51710 15750 51762 15802
rect 51774 15750 51826 15802
rect 15398 15206 15450 15258
rect 15462 15206 15514 15258
rect 15526 15206 15578 15258
rect 15590 15206 15642 15258
rect 15654 15206 15706 15258
rect 29846 15206 29898 15258
rect 29910 15206 29962 15258
rect 29974 15206 30026 15258
rect 30038 15206 30090 15258
rect 30102 15206 30154 15258
rect 44294 15206 44346 15258
rect 44358 15206 44410 15258
rect 44422 15206 44474 15258
rect 44486 15206 44538 15258
rect 44550 15206 44602 15258
rect 8174 14662 8226 14714
rect 8238 14662 8290 14714
rect 8302 14662 8354 14714
rect 8366 14662 8418 14714
rect 8430 14662 8482 14714
rect 22622 14662 22674 14714
rect 22686 14662 22738 14714
rect 22750 14662 22802 14714
rect 22814 14662 22866 14714
rect 22878 14662 22930 14714
rect 37070 14662 37122 14714
rect 37134 14662 37186 14714
rect 37198 14662 37250 14714
rect 37262 14662 37314 14714
rect 37326 14662 37378 14714
rect 51518 14662 51570 14714
rect 51582 14662 51634 14714
rect 51646 14662 51698 14714
rect 51710 14662 51762 14714
rect 51774 14662 51826 14714
rect 15398 14118 15450 14170
rect 15462 14118 15514 14170
rect 15526 14118 15578 14170
rect 15590 14118 15642 14170
rect 15654 14118 15706 14170
rect 29846 14118 29898 14170
rect 29910 14118 29962 14170
rect 29974 14118 30026 14170
rect 30038 14118 30090 14170
rect 30102 14118 30154 14170
rect 44294 14118 44346 14170
rect 44358 14118 44410 14170
rect 44422 14118 44474 14170
rect 44486 14118 44538 14170
rect 44550 14118 44602 14170
rect 20260 13880 20312 13932
rect 3148 13812 3200 13864
rect 13360 13855 13412 13864
rect 13360 13821 13369 13855
rect 13369 13821 13403 13855
rect 13403 13821 13412 13855
rect 13360 13812 13412 13821
rect 25412 13812 25464 13864
rect 8174 13574 8226 13626
rect 8238 13574 8290 13626
rect 8302 13574 8354 13626
rect 8366 13574 8418 13626
rect 8430 13574 8482 13626
rect 22622 13574 22674 13626
rect 22686 13574 22738 13626
rect 22750 13574 22802 13626
rect 22814 13574 22866 13626
rect 22878 13574 22930 13626
rect 37070 13574 37122 13626
rect 37134 13574 37186 13626
rect 37198 13574 37250 13626
rect 37262 13574 37314 13626
rect 37326 13574 37378 13626
rect 51518 13574 51570 13626
rect 51582 13574 51634 13626
rect 51646 13574 51698 13626
rect 51710 13574 51762 13626
rect 51774 13574 51826 13626
rect 11428 13311 11480 13320
rect 11428 13277 11437 13311
rect 11437 13277 11471 13311
rect 11471 13277 11480 13311
rect 11428 13268 11480 13277
rect 15200 13268 15252 13320
rect 5264 13200 5316 13252
rect 9496 13200 9548 13252
rect 12992 13200 13044 13252
rect 22284 13268 22336 13320
rect 16948 13243 17000 13252
rect 16948 13209 16957 13243
rect 16957 13209 16991 13243
rect 16991 13209 17000 13243
rect 16948 13200 17000 13209
rect 19708 13200 19760 13252
rect 1492 13132 1544 13184
rect 2688 13175 2740 13184
rect 2688 13141 2697 13175
rect 2697 13141 2731 13175
rect 2731 13141 2740 13175
rect 2688 13132 2740 13141
rect 3240 13175 3292 13184
rect 3240 13141 3249 13175
rect 3249 13141 3283 13175
rect 3283 13141 3292 13175
rect 3240 13132 3292 13141
rect 3792 13175 3844 13184
rect 3792 13141 3801 13175
rect 3801 13141 3835 13175
rect 3835 13141 3844 13175
rect 3792 13132 3844 13141
rect 4988 13132 5040 13184
rect 6276 13132 6328 13184
rect 9588 13132 9640 13184
rect 9680 13132 9732 13184
rect 11060 13132 11112 13184
rect 11612 13132 11664 13184
rect 12900 13132 12952 13184
rect 14188 13175 14240 13184
rect 14188 13141 14197 13175
rect 14197 13141 14231 13175
rect 14231 13141 14240 13175
rect 14188 13132 14240 13141
rect 15108 13175 15160 13184
rect 15108 13141 15117 13175
rect 15117 13141 15151 13175
rect 15151 13141 15160 13175
rect 15108 13132 15160 13141
rect 15844 13132 15896 13184
rect 17776 13175 17828 13184
rect 17776 13141 17785 13175
rect 17785 13141 17819 13175
rect 17819 13141 17828 13175
rect 17776 13132 17828 13141
rect 18052 13132 18104 13184
rect 27804 13132 27856 13184
rect 15398 13030 15450 13082
rect 15462 13030 15514 13082
rect 15526 13030 15578 13082
rect 15590 13030 15642 13082
rect 15654 13030 15706 13082
rect 29846 13030 29898 13082
rect 29910 13030 29962 13082
rect 29974 13030 30026 13082
rect 30038 13030 30090 13082
rect 30102 13030 30154 13082
rect 44294 13030 44346 13082
rect 44358 13030 44410 13082
rect 44422 13030 44474 13082
rect 44486 13030 44538 13082
rect 44550 13030 44602 13082
rect 9496 12971 9548 12980
rect 9496 12937 9505 12971
rect 9505 12937 9539 12971
rect 9539 12937 9548 12971
rect 9496 12928 9548 12937
rect 12992 12971 13044 12980
rect 12992 12937 13001 12971
rect 13001 12937 13035 12971
rect 13035 12937 13044 12971
rect 12992 12928 13044 12937
rect 3976 12860 4028 12912
rect 15108 12928 15160 12980
rect 15200 12928 15252 12980
rect 18236 12860 18288 12912
rect 21916 12903 21968 12912
rect 21916 12869 21925 12903
rect 21925 12869 21959 12903
rect 21959 12869 21968 12903
rect 21916 12860 21968 12869
rect 25044 12860 25096 12912
rect 5908 12792 5960 12844
rect 12900 12792 12952 12844
rect 17224 12792 17276 12844
rect 22100 12792 22152 12844
rect 11428 12724 11480 12776
rect 3148 12656 3200 12708
rect 1952 12631 2004 12640
rect 1952 12597 1961 12631
rect 1961 12597 1995 12631
rect 1995 12597 2004 12631
rect 1952 12588 2004 12597
rect 3608 12631 3660 12640
rect 3608 12597 3617 12631
rect 3617 12597 3651 12631
rect 3651 12597 3660 12631
rect 3608 12588 3660 12597
rect 5264 12631 5316 12640
rect 5264 12597 5273 12631
rect 5273 12597 5307 12631
rect 5307 12597 5316 12631
rect 5264 12588 5316 12597
rect 6552 12588 6604 12640
rect 9220 12656 9272 12708
rect 7012 12631 7064 12640
rect 7012 12597 7021 12631
rect 7021 12597 7055 12631
rect 7055 12597 7064 12631
rect 7012 12588 7064 12597
rect 7932 12588 7984 12640
rect 8852 12631 8904 12640
rect 8852 12597 8861 12631
rect 8861 12597 8895 12631
rect 8895 12597 8904 12631
rect 8852 12588 8904 12597
rect 10968 12631 11020 12640
rect 10968 12597 10977 12631
rect 10977 12597 11011 12631
rect 11011 12597 11020 12631
rect 10968 12588 11020 12597
rect 11704 12588 11756 12640
rect 16948 12724 17000 12776
rect 19064 12724 19116 12776
rect 23664 12724 23716 12776
rect 13176 12656 13228 12708
rect 20076 12656 20128 12708
rect 25136 12656 25188 12708
rect 16120 12631 16172 12640
rect 16120 12597 16129 12631
rect 16129 12597 16163 12631
rect 16163 12597 16172 12631
rect 16120 12588 16172 12597
rect 17224 12588 17276 12640
rect 18236 12631 18288 12640
rect 18236 12597 18245 12631
rect 18245 12597 18279 12631
rect 18279 12597 18288 12631
rect 18236 12588 18288 12597
rect 19984 12588 20036 12640
rect 20720 12631 20772 12640
rect 20720 12597 20729 12631
rect 20729 12597 20763 12631
rect 20763 12597 20772 12631
rect 20720 12588 20772 12597
rect 23480 12631 23532 12640
rect 23480 12597 23489 12631
rect 23489 12597 23523 12631
rect 23523 12597 23532 12631
rect 23480 12588 23532 12597
rect 23940 12631 23992 12640
rect 23940 12597 23949 12631
rect 23949 12597 23983 12631
rect 23983 12597 23992 12631
rect 23940 12588 23992 12597
rect 8174 12486 8226 12538
rect 8238 12486 8290 12538
rect 8302 12486 8354 12538
rect 8366 12486 8418 12538
rect 8430 12486 8482 12538
rect 22622 12486 22674 12538
rect 22686 12486 22738 12538
rect 22750 12486 22802 12538
rect 22814 12486 22866 12538
rect 22878 12486 22930 12538
rect 37070 12486 37122 12538
rect 37134 12486 37186 12538
rect 37198 12486 37250 12538
rect 37262 12486 37314 12538
rect 37326 12486 37378 12538
rect 51518 12486 51570 12538
rect 51582 12486 51634 12538
rect 51646 12486 51698 12538
rect 51710 12486 51762 12538
rect 51774 12486 51826 12538
rect 6552 12427 6604 12436
rect 6552 12393 6561 12427
rect 6561 12393 6595 12427
rect 6595 12393 6604 12427
rect 6552 12384 6604 12393
rect 9220 12427 9272 12436
rect 9220 12393 9229 12427
rect 9229 12393 9263 12427
rect 9263 12393 9272 12427
rect 9220 12384 9272 12393
rect 25136 12427 25188 12436
rect 25136 12393 25145 12427
rect 25145 12393 25179 12427
rect 25179 12393 25188 12427
rect 25136 12384 25188 12393
rect 10968 12316 11020 12368
rect 20168 12316 20220 12368
rect 1860 12180 1912 12232
rect 3148 12180 3200 12232
rect 3332 12180 3384 12232
rect 8576 12180 8628 12232
rect 19248 12180 19300 12232
rect 20536 12180 20588 12232
rect 5908 12112 5960 12164
rect 6920 12112 6972 12164
rect 17224 12112 17276 12164
rect 20076 12112 20128 12164
rect 22468 12180 22520 12232
rect 1676 12044 1728 12096
rect 2964 12044 3016 12096
rect 3884 12087 3936 12096
rect 3884 12053 3893 12087
rect 3893 12053 3927 12087
rect 3927 12053 3936 12087
rect 3884 12044 3936 12053
rect 5172 12087 5224 12096
rect 5172 12053 5181 12087
rect 5181 12053 5215 12087
rect 5215 12053 5224 12087
rect 5172 12044 5224 12053
rect 7840 12044 7892 12096
rect 8668 12044 8720 12096
rect 10048 12087 10100 12096
rect 10048 12053 10057 12087
rect 10057 12053 10091 12087
rect 10091 12053 10100 12087
rect 10048 12044 10100 12053
rect 10324 12044 10376 12096
rect 11152 12044 11204 12096
rect 12440 12044 12492 12096
rect 13268 12044 13320 12096
rect 14188 12087 14240 12096
rect 14188 12053 14197 12087
rect 14197 12053 14231 12087
rect 14231 12053 14240 12087
rect 14188 12044 14240 12053
rect 14648 12044 14700 12096
rect 16580 12044 16632 12096
rect 16948 12044 17000 12096
rect 18604 12087 18656 12096
rect 18604 12053 18613 12087
rect 18613 12053 18647 12087
rect 18647 12053 18656 12087
rect 18604 12044 18656 12053
rect 18788 12044 18840 12096
rect 19708 12044 19760 12096
rect 20628 12044 20680 12096
rect 22284 12087 22336 12096
rect 22284 12053 22293 12087
rect 22293 12053 22327 12087
rect 22327 12053 22336 12087
rect 22284 12044 22336 12053
rect 23848 12044 23900 12096
rect 24032 12044 24084 12096
rect 25596 12087 25648 12096
rect 25596 12053 25605 12087
rect 25605 12053 25639 12087
rect 25639 12053 25648 12087
rect 25596 12044 25648 12053
rect 36820 12044 36872 12096
rect 15398 11942 15450 11994
rect 15462 11942 15514 11994
rect 15526 11942 15578 11994
rect 15590 11942 15642 11994
rect 15654 11942 15706 11994
rect 29846 11942 29898 11994
rect 29910 11942 29962 11994
rect 29974 11942 30026 11994
rect 30038 11942 30090 11994
rect 30102 11942 30154 11994
rect 44294 11942 44346 11994
rect 44358 11942 44410 11994
rect 44422 11942 44474 11994
rect 44486 11942 44538 11994
rect 44550 11942 44602 11994
rect 2964 11883 3016 11892
rect 2964 11849 2973 11883
rect 2973 11849 3007 11883
rect 3007 11849 3016 11883
rect 2964 11840 3016 11849
rect 6920 11883 6972 11892
rect 6920 11849 6929 11883
rect 6929 11849 6963 11883
rect 6963 11849 6972 11883
rect 6920 11840 6972 11849
rect 8576 11840 8628 11892
rect 20076 11883 20128 11892
rect 20076 11849 20085 11883
rect 20085 11849 20119 11883
rect 20119 11849 20128 11883
rect 20076 11840 20128 11849
rect 22468 11840 22520 11892
rect 23112 11883 23164 11892
rect 23112 11849 23121 11883
rect 23121 11849 23155 11883
rect 23155 11849 23164 11883
rect 23112 11840 23164 11849
rect 4252 11772 4304 11824
rect 21916 11772 21968 11824
rect 11704 11704 11756 11756
rect 45652 11704 45704 11756
rect 20996 11636 21048 11688
rect 36544 11636 36596 11688
rect 3424 11568 3476 11620
rect 3608 11568 3660 11620
rect 14556 11611 14608 11620
rect 14556 11577 14565 11611
rect 14565 11577 14599 11611
rect 14599 11577 14608 11611
rect 14556 11568 14608 11577
rect 16580 11568 16632 11620
rect 23572 11568 23624 11620
rect 23756 11568 23808 11620
rect 1584 11500 1636 11552
rect 4344 11500 4396 11552
rect 4896 11543 4948 11552
rect 4896 11509 4905 11543
rect 4905 11509 4939 11543
rect 4939 11509 4948 11543
rect 4896 11500 4948 11509
rect 5816 11543 5868 11552
rect 5816 11509 5825 11543
rect 5825 11509 5859 11543
rect 5859 11509 5868 11543
rect 5816 11500 5868 11509
rect 7472 11500 7524 11552
rect 7656 11500 7708 11552
rect 9680 11500 9732 11552
rect 10416 11543 10468 11552
rect 10416 11509 10425 11543
rect 10425 11509 10459 11543
rect 10459 11509 10468 11543
rect 10416 11500 10468 11509
rect 12440 11543 12492 11552
rect 12440 11509 12449 11543
rect 12449 11509 12483 11543
rect 12483 11509 12492 11543
rect 12440 11500 12492 11509
rect 12808 11500 12860 11552
rect 13636 11543 13688 11552
rect 13636 11509 13645 11543
rect 13645 11509 13679 11543
rect 13679 11509 13688 11543
rect 13636 11500 13688 11509
rect 15016 11500 15068 11552
rect 15752 11500 15804 11552
rect 16304 11500 16356 11552
rect 17224 11543 17276 11552
rect 17224 11509 17233 11543
rect 17233 11509 17267 11543
rect 17267 11509 17276 11543
rect 17224 11500 17276 11509
rect 18236 11543 18288 11552
rect 18236 11509 18245 11543
rect 18245 11509 18279 11543
rect 18279 11509 18288 11543
rect 18236 11500 18288 11509
rect 19248 11543 19300 11552
rect 19248 11509 19257 11543
rect 19257 11509 19291 11543
rect 19291 11509 19300 11543
rect 19248 11500 19300 11509
rect 19800 11500 19852 11552
rect 20260 11500 20312 11552
rect 21732 11500 21784 11552
rect 22100 11543 22152 11552
rect 22100 11509 22109 11543
rect 22109 11509 22143 11543
rect 22143 11509 22152 11543
rect 22100 11500 22152 11509
rect 23204 11500 23256 11552
rect 24492 11543 24544 11552
rect 24492 11509 24501 11543
rect 24501 11509 24535 11543
rect 24535 11509 24544 11543
rect 24492 11500 24544 11509
rect 24952 11500 25004 11552
rect 25412 11500 25464 11552
rect 27436 11568 27488 11620
rect 41788 11568 41840 11620
rect 27988 11500 28040 11552
rect 35716 11543 35768 11552
rect 35716 11509 35725 11543
rect 35725 11509 35759 11543
rect 35759 11509 35768 11543
rect 35716 11500 35768 11509
rect 37648 11500 37700 11552
rect 38384 11543 38436 11552
rect 38384 11509 38393 11543
rect 38393 11509 38427 11543
rect 38427 11509 38436 11543
rect 38384 11500 38436 11509
rect 43076 11500 43128 11552
rect 43536 11500 43588 11552
rect 8174 11398 8226 11450
rect 8238 11398 8290 11450
rect 8302 11398 8354 11450
rect 8366 11398 8418 11450
rect 8430 11398 8482 11450
rect 22622 11398 22674 11450
rect 22686 11398 22738 11450
rect 22750 11398 22802 11450
rect 22814 11398 22866 11450
rect 22878 11398 22930 11450
rect 37070 11398 37122 11450
rect 37134 11398 37186 11450
rect 37198 11398 37250 11450
rect 37262 11398 37314 11450
rect 37326 11398 37378 11450
rect 51518 11398 51570 11450
rect 51582 11398 51634 11450
rect 51646 11398 51698 11450
rect 51710 11398 51762 11450
rect 51774 11398 51826 11450
rect 3884 11296 3936 11348
rect 12716 11296 12768 11348
rect 13636 11296 13688 11348
rect 22468 11296 22520 11348
rect 25504 11339 25556 11348
rect 25504 11305 25513 11339
rect 25513 11305 25547 11339
rect 25547 11305 25556 11339
rect 25504 11296 25556 11305
rect 26332 11296 26384 11348
rect 38384 11296 38436 11348
rect 41144 11296 41196 11348
rect 43352 11339 43404 11348
rect 43352 11305 43361 11339
rect 43361 11305 43395 11339
rect 43395 11305 43404 11339
rect 43352 11296 43404 11305
rect 2044 11271 2096 11280
rect 2044 11237 2053 11271
rect 2053 11237 2087 11271
rect 2087 11237 2096 11271
rect 2044 11228 2096 11237
rect 5908 11271 5960 11280
rect 5908 11237 5917 11271
rect 5917 11237 5951 11271
rect 5951 11237 5960 11271
rect 5908 11228 5960 11237
rect 6368 11228 6420 11280
rect 7748 11271 7800 11280
rect 3608 11160 3660 11212
rect 7748 11237 7757 11271
rect 7757 11237 7791 11271
rect 7791 11237 7800 11271
rect 7748 11228 7800 11237
rect 9036 11228 9088 11280
rect 10968 11228 11020 11280
rect 15660 11271 15712 11280
rect 15660 11237 15669 11271
rect 15669 11237 15703 11271
rect 15703 11237 15712 11271
rect 15660 11228 15712 11237
rect 16028 11228 16080 11280
rect 20168 11271 20220 11280
rect 20168 11237 20177 11271
rect 20177 11237 20211 11271
rect 20211 11237 20220 11271
rect 20168 11228 20220 11237
rect 4436 11092 4488 11144
rect 4988 11092 5040 11144
rect 7104 11135 7156 11144
rect 7104 11101 7113 11135
rect 7113 11101 7147 11135
rect 7147 11101 7156 11135
rect 7104 11092 7156 11101
rect 4160 11067 4212 11076
rect 4160 11033 4169 11067
rect 4169 11033 4203 11067
rect 4203 11033 4212 11067
rect 4160 11024 4212 11033
rect 4896 11024 4948 11076
rect 5816 11024 5868 11076
rect 13636 11160 13688 11212
rect 15844 11160 15896 11212
rect 21548 11228 21600 11280
rect 22100 11228 22152 11280
rect 24768 11228 24820 11280
rect 38752 11228 38804 11280
rect 39488 11228 39540 11280
rect 20996 11203 21048 11212
rect 20996 11169 21005 11203
rect 21005 11169 21039 11203
rect 21039 11169 21048 11203
rect 20996 11160 21048 11169
rect 7472 11092 7524 11144
rect 12348 11092 12400 11144
rect 13084 11092 13136 11144
rect 13360 11135 13412 11144
rect 13360 11101 13369 11135
rect 13369 11101 13403 11135
rect 13403 11101 13412 11135
rect 13360 11092 13412 11101
rect 13912 11092 13964 11144
rect 16304 11135 16356 11144
rect 8576 11024 8628 11076
rect 9220 11024 9272 11076
rect 2596 10999 2648 11008
rect 2596 10965 2605 10999
rect 2605 10965 2639 10999
rect 2639 10965 2648 10999
rect 2596 10956 2648 10965
rect 3792 10956 3844 11008
rect 8484 10956 8536 11008
rect 9956 11024 10008 11076
rect 13268 11024 13320 11076
rect 16304 11101 16313 11135
rect 16313 11101 16347 11135
rect 16347 11101 16356 11135
rect 16304 11092 16356 11101
rect 16856 11092 16908 11144
rect 18604 11092 18656 11144
rect 19248 11092 19300 11144
rect 22100 11092 22152 11144
rect 22192 11135 22244 11144
rect 22192 11101 22201 11135
rect 22201 11101 22235 11135
rect 22235 11101 22244 11135
rect 36636 11160 36688 11212
rect 22192 11092 22244 11101
rect 15844 11024 15896 11076
rect 18788 11024 18840 11076
rect 19524 11024 19576 11076
rect 21456 11067 21508 11076
rect 21456 11033 21465 11067
rect 21465 11033 21499 11067
rect 21499 11033 21508 11067
rect 21456 11024 21508 11033
rect 21548 11024 21600 11076
rect 22468 11024 22520 11076
rect 24124 11024 24176 11076
rect 25872 11024 25924 11076
rect 26608 11067 26660 11076
rect 26608 11033 26617 11067
rect 26617 11033 26651 11067
rect 26651 11033 26660 11067
rect 26608 11024 26660 11033
rect 26700 11024 26752 11076
rect 27436 11092 27488 11144
rect 27988 11092 28040 11144
rect 38660 11092 38712 11144
rect 27528 11024 27580 11076
rect 29368 11024 29420 11076
rect 35164 11067 35216 11076
rect 35164 11033 35173 11067
rect 35173 11033 35207 11067
rect 35207 11033 35216 11067
rect 35164 11024 35216 11033
rect 36176 11067 36228 11076
rect 36176 11033 36185 11067
rect 36185 11033 36219 11067
rect 36219 11033 36228 11067
rect 36176 11024 36228 11033
rect 36636 11024 36688 11076
rect 23388 10956 23440 11008
rect 23664 10956 23716 11008
rect 36912 10956 36964 11008
rect 40408 11067 40460 11076
rect 40408 11033 40417 11067
rect 40417 11033 40451 11067
rect 40451 11033 40460 11067
rect 40408 11024 40460 11033
rect 41972 11067 42024 11076
rect 41972 11033 41981 11067
rect 41981 11033 42015 11067
rect 42015 11033 42024 11067
rect 41972 11024 42024 11033
rect 42892 11024 42944 11076
rect 43812 11024 43864 11076
rect 38200 10956 38252 11008
rect 38568 10999 38620 11008
rect 38568 10965 38577 10999
rect 38577 10965 38611 10999
rect 38611 10965 38620 10999
rect 38568 10956 38620 10965
rect 45008 10999 45060 11008
rect 45008 10965 45017 10999
rect 45017 10965 45051 10999
rect 45051 10965 45060 10999
rect 45008 10956 45060 10965
rect 15398 10854 15450 10906
rect 15462 10854 15514 10906
rect 15526 10854 15578 10906
rect 15590 10854 15642 10906
rect 15654 10854 15706 10906
rect 29846 10854 29898 10906
rect 29910 10854 29962 10906
rect 29974 10854 30026 10906
rect 30038 10854 30090 10906
rect 30102 10854 30154 10906
rect 44294 10854 44346 10906
rect 44358 10854 44410 10906
rect 44422 10854 44474 10906
rect 44486 10854 44538 10906
rect 44550 10854 44602 10906
rect 1768 10795 1820 10804
rect 1768 10761 1777 10795
rect 1777 10761 1811 10795
rect 1811 10761 1820 10795
rect 1768 10752 1820 10761
rect 2596 10752 2648 10804
rect 3792 10752 3844 10804
rect 3976 10795 4028 10804
rect 3976 10761 3985 10795
rect 3985 10761 4019 10795
rect 4019 10761 4028 10795
rect 3976 10752 4028 10761
rect 5816 10795 5868 10804
rect 5816 10761 5825 10795
rect 5825 10761 5859 10795
rect 5859 10761 5868 10795
rect 5816 10752 5868 10761
rect 1584 10659 1636 10668
rect 1584 10625 1593 10659
rect 1593 10625 1627 10659
rect 1627 10625 1636 10659
rect 1584 10616 1636 10625
rect 2688 10684 2740 10736
rect 23296 10752 23348 10804
rect 26240 10752 26292 10804
rect 36544 10795 36596 10804
rect 36544 10761 36553 10795
rect 36553 10761 36587 10795
rect 36587 10761 36596 10795
rect 36544 10752 36596 10761
rect 37464 10752 37516 10804
rect 38568 10752 38620 10804
rect 39488 10795 39540 10804
rect 39488 10761 39497 10795
rect 39497 10761 39531 10795
rect 39531 10761 39540 10795
rect 39488 10752 39540 10761
rect 41144 10795 41196 10804
rect 41144 10761 41153 10795
rect 41153 10761 41187 10795
rect 41187 10761 41196 10795
rect 41144 10752 41196 10761
rect 41788 10795 41840 10804
rect 41788 10761 41797 10795
rect 41797 10761 41831 10795
rect 41831 10761 41840 10795
rect 41788 10752 41840 10761
rect 43352 10752 43404 10804
rect 44088 10752 44140 10804
rect 10048 10684 10100 10736
rect 14188 10684 14240 10736
rect 4160 10616 4212 10668
rect 4712 10659 4764 10668
rect 4712 10625 4721 10659
rect 4721 10625 4755 10659
rect 4755 10625 4764 10659
rect 4712 10616 4764 10625
rect 7380 10616 7432 10668
rect 2044 10548 2096 10600
rect 7012 10548 7064 10600
rect 7656 10548 7708 10600
rect 9312 10616 9364 10668
rect 10140 10616 10192 10668
rect 11796 10659 11848 10668
rect 11796 10625 11805 10659
rect 11805 10625 11839 10659
rect 11839 10625 11848 10659
rect 11796 10616 11848 10625
rect 15844 10616 15896 10668
rect 16212 10616 16264 10668
rect 17684 10659 17736 10668
rect 17684 10625 17693 10659
rect 17693 10625 17727 10659
rect 17727 10625 17736 10659
rect 17684 10616 17736 10625
rect 28908 10684 28960 10736
rect 34612 10684 34664 10736
rect 35256 10684 35308 10736
rect 46940 10727 46992 10736
rect 46940 10693 46949 10727
rect 46949 10693 46983 10727
rect 46983 10693 46992 10727
rect 46940 10684 46992 10693
rect 22376 10616 22428 10668
rect 23480 10659 23532 10668
rect 23480 10625 23489 10659
rect 23489 10625 23523 10659
rect 23523 10625 23532 10659
rect 23480 10616 23532 10625
rect 25228 10616 25280 10668
rect 27160 10659 27212 10668
rect 27160 10625 27169 10659
rect 27169 10625 27203 10659
rect 27203 10625 27212 10659
rect 27160 10616 27212 10625
rect 28816 10616 28868 10668
rect 38660 10616 38712 10668
rect 11428 10548 11480 10600
rect 17316 10548 17368 10600
rect 20168 10548 20220 10600
rect 23388 10548 23440 10600
rect 26056 10548 26108 10600
rect 31208 10548 31260 10600
rect 34520 10548 34572 10600
rect 36912 10548 36964 10600
rect 8944 10480 8996 10532
rect 14280 10480 14332 10532
rect 16120 10480 16172 10532
rect 20260 10480 20312 10532
rect 24676 10480 24728 10532
rect 29092 10480 29144 10532
rect 38200 10480 38252 10532
rect 2688 10412 2740 10464
rect 3792 10412 3844 10464
rect 4896 10455 4948 10464
rect 4896 10421 4905 10455
rect 4905 10421 4939 10455
rect 4939 10421 4948 10455
rect 4896 10412 4948 10421
rect 6920 10455 6972 10464
rect 6920 10421 6929 10455
rect 6929 10421 6963 10455
rect 6963 10421 6972 10455
rect 6920 10412 6972 10421
rect 9588 10455 9640 10464
rect 9588 10421 9597 10455
rect 9597 10421 9631 10455
rect 9631 10421 9640 10455
rect 9588 10412 9640 10421
rect 12256 10412 12308 10464
rect 13452 10412 13504 10464
rect 14740 10412 14792 10464
rect 15292 10412 15344 10464
rect 15936 10455 15988 10464
rect 15936 10421 15945 10455
rect 15945 10421 15979 10455
rect 15979 10421 15988 10455
rect 15936 10412 15988 10421
rect 17408 10412 17460 10464
rect 18420 10455 18472 10464
rect 18420 10421 18429 10455
rect 18429 10421 18463 10455
rect 18463 10421 18472 10455
rect 18420 10412 18472 10421
rect 20444 10412 20496 10464
rect 22100 10455 22152 10464
rect 22100 10421 22109 10455
rect 22109 10421 22143 10455
rect 22143 10421 22152 10455
rect 22100 10412 22152 10421
rect 23020 10412 23072 10464
rect 24216 10412 24268 10464
rect 26424 10412 26476 10464
rect 27620 10412 27672 10464
rect 29552 10455 29604 10464
rect 29552 10421 29561 10455
rect 29561 10421 29595 10455
rect 29595 10421 29604 10455
rect 29552 10412 29604 10421
rect 30196 10412 30248 10464
rect 33140 10412 33192 10464
rect 34796 10412 34848 10464
rect 36084 10455 36136 10464
rect 36084 10421 36093 10455
rect 36093 10421 36127 10455
rect 36127 10421 36136 10455
rect 36084 10412 36136 10421
rect 37556 10412 37608 10464
rect 43996 10548 44048 10600
rect 46756 10616 46808 10668
rect 50528 10548 50580 10600
rect 41236 10480 41288 10532
rect 45008 10480 45060 10532
rect 39856 10412 39908 10464
rect 40500 10412 40552 10464
rect 42524 10455 42576 10464
rect 42524 10421 42533 10455
rect 42533 10421 42567 10455
rect 42567 10421 42576 10455
rect 42524 10412 42576 10421
rect 42892 10412 42944 10464
rect 43996 10455 44048 10464
rect 43996 10421 44005 10455
rect 44005 10421 44039 10455
rect 44039 10421 44048 10455
rect 43996 10412 44048 10421
rect 45468 10412 45520 10464
rect 46388 10455 46440 10464
rect 46388 10421 46397 10455
rect 46397 10421 46431 10455
rect 46431 10421 46440 10455
rect 46388 10412 46440 10421
rect 48964 10412 49016 10464
rect 8174 10310 8226 10362
rect 8238 10310 8290 10362
rect 8302 10310 8354 10362
rect 8366 10310 8418 10362
rect 8430 10310 8482 10362
rect 22622 10310 22674 10362
rect 22686 10310 22738 10362
rect 22750 10310 22802 10362
rect 22814 10310 22866 10362
rect 22878 10310 22930 10362
rect 37070 10310 37122 10362
rect 37134 10310 37186 10362
rect 37198 10310 37250 10362
rect 37262 10310 37314 10362
rect 37326 10310 37378 10362
rect 51518 10310 51570 10362
rect 51582 10310 51634 10362
rect 51646 10310 51698 10362
rect 51710 10310 51762 10362
rect 51774 10310 51826 10362
rect 1676 10047 1728 10056
rect 1676 10013 1685 10047
rect 1685 10013 1719 10047
rect 1719 10013 1728 10047
rect 1676 10004 1728 10013
rect 2964 10047 3016 10056
rect 2964 10013 2973 10047
rect 2973 10013 3007 10047
rect 3007 10013 3016 10047
rect 2964 10004 3016 10013
rect 4068 10208 4120 10260
rect 5632 10047 5684 10056
rect 5632 10013 5641 10047
rect 5641 10013 5675 10047
rect 5675 10013 5684 10047
rect 5632 10004 5684 10013
rect 6920 10208 6972 10260
rect 11796 10208 11848 10260
rect 11428 10072 11480 10124
rect 17684 10208 17736 10260
rect 17776 10208 17828 10260
rect 46388 10208 46440 10260
rect 47216 10208 47268 10260
rect 35256 10183 35308 10192
rect 35256 10149 35265 10183
rect 35265 10149 35299 10183
rect 35299 10149 35308 10183
rect 35256 10140 35308 10149
rect 38660 10140 38712 10192
rect 20904 10072 20956 10124
rect 22560 10115 22612 10124
rect 22560 10081 22569 10115
rect 22569 10081 22603 10115
rect 22603 10081 22612 10115
rect 22560 10072 22612 10081
rect 32312 10072 32364 10124
rect 4436 9936 4488 9988
rect 9128 10004 9180 10056
rect 10048 10047 10100 10056
rect 10048 10013 10057 10047
rect 10057 10013 10091 10047
rect 10091 10013 10100 10047
rect 10048 10004 10100 10013
rect 11244 10004 11296 10056
rect 11336 10047 11388 10056
rect 11336 10013 11345 10047
rect 11345 10013 11379 10047
rect 11379 10013 11388 10047
rect 11336 10004 11388 10013
rect 14096 10047 14148 10056
rect 10784 9936 10836 9988
rect 14096 10013 14105 10047
rect 14105 10013 14139 10047
rect 14139 10013 14148 10047
rect 14096 10004 14148 10013
rect 1860 9911 1912 9920
rect 1860 9877 1869 9911
rect 1869 9877 1903 9911
rect 1903 9877 1912 9911
rect 1860 9868 1912 9877
rect 2504 9911 2556 9920
rect 2504 9877 2513 9911
rect 2513 9877 2547 9911
rect 2547 9877 2556 9911
rect 2504 9868 2556 9877
rect 4804 9911 4856 9920
rect 4804 9877 4813 9911
rect 4813 9877 4847 9911
rect 4847 9877 4856 9911
rect 4804 9868 4856 9877
rect 7564 9868 7616 9920
rect 7840 9868 7892 9920
rect 10232 9868 10284 9920
rect 12624 9868 12676 9920
rect 13452 9868 13504 9920
rect 14188 9868 14240 9920
rect 14924 9868 14976 9920
rect 17316 10047 17368 10056
rect 17316 10013 17325 10047
rect 17325 10013 17359 10047
rect 17359 10013 17368 10047
rect 17316 10004 17368 10013
rect 18144 10004 18196 10056
rect 18512 10047 18564 10056
rect 18512 10013 18521 10047
rect 18521 10013 18555 10047
rect 18555 10013 18564 10047
rect 18512 10004 18564 10013
rect 20444 10047 20496 10056
rect 20444 10013 20453 10047
rect 20453 10013 20487 10047
rect 20487 10013 20496 10047
rect 20444 10004 20496 10013
rect 22284 10004 22336 10056
rect 23020 10004 23072 10056
rect 24400 10047 24452 10056
rect 24400 10013 24409 10047
rect 24409 10013 24443 10047
rect 24443 10013 24452 10047
rect 24400 10004 24452 10013
rect 24676 10047 24728 10056
rect 24676 10013 24685 10047
rect 24685 10013 24719 10047
rect 24719 10013 24728 10047
rect 24676 10004 24728 10013
rect 25688 10004 25740 10056
rect 26424 10047 26476 10056
rect 26424 10013 26433 10047
rect 26433 10013 26467 10047
rect 26467 10013 26476 10047
rect 26424 10004 26476 10013
rect 30840 10047 30892 10056
rect 30840 10013 30849 10047
rect 30849 10013 30883 10047
rect 30883 10013 30892 10047
rect 30840 10004 30892 10013
rect 15476 9868 15528 9920
rect 18420 9868 18472 9920
rect 19708 9911 19760 9920
rect 19708 9877 19717 9911
rect 19717 9877 19751 9911
rect 19751 9877 19760 9911
rect 19708 9868 19760 9877
rect 24860 9936 24912 9988
rect 21916 9911 21968 9920
rect 21916 9877 21925 9911
rect 21925 9877 21959 9911
rect 21959 9877 21968 9911
rect 21916 9868 21968 9877
rect 22008 9868 22060 9920
rect 27988 9936 28040 9988
rect 28080 9936 28132 9988
rect 28908 9936 28960 9988
rect 30564 9936 30616 9988
rect 31208 10004 31260 10056
rect 27344 9868 27396 9920
rect 28448 9868 28500 9920
rect 29460 9868 29512 9920
rect 30288 9868 30340 9920
rect 32496 9868 32548 9920
rect 32588 9911 32640 9920
rect 32588 9877 32597 9911
rect 32597 9877 32631 9911
rect 32631 9877 32640 9911
rect 48964 10072 49016 10124
rect 52276 10115 52328 10124
rect 52276 10081 52285 10115
rect 52285 10081 52319 10115
rect 52319 10081 52328 10115
rect 52276 10072 52328 10081
rect 33324 10004 33376 10056
rect 36544 10004 36596 10056
rect 38108 10047 38160 10056
rect 34152 9911 34204 9920
rect 32588 9868 32640 9877
rect 34152 9877 34161 9911
rect 34161 9877 34195 9911
rect 34195 9877 34204 9911
rect 34152 9868 34204 9877
rect 36176 9868 36228 9920
rect 36360 9911 36412 9920
rect 36360 9877 36369 9911
rect 36369 9877 36403 9911
rect 36403 9877 36412 9911
rect 36360 9868 36412 9877
rect 36912 9868 36964 9920
rect 37372 9911 37424 9920
rect 37372 9877 37381 9911
rect 37381 9877 37415 9911
rect 37415 9877 37424 9911
rect 37372 9868 37424 9877
rect 38108 10013 38117 10047
rect 38117 10013 38151 10047
rect 38151 10013 38160 10047
rect 38108 10004 38160 10013
rect 38016 9936 38068 9988
rect 40224 10004 40276 10056
rect 42432 10004 42484 10056
rect 42984 10047 43036 10056
rect 42984 10013 42993 10047
rect 42993 10013 43027 10047
rect 43027 10013 43036 10047
rect 42984 10004 43036 10013
rect 45652 10047 45704 10056
rect 45652 10013 45661 10047
rect 45661 10013 45695 10047
rect 45695 10013 45704 10047
rect 45652 10004 45704 10013
rect 46480 10047 46532 10056
rect 46480 10013 46489 10047
rect 46489 10013 46523 10047
rect 46523 10013 46532 10047
rect 46480 10004 46532 10013
rect 46756 10047 46808 10056
rect 46756 10013 46765 10047
rect 46765 10013 46799 10047
rect 46799 10013 46808 10047
rect 46756 10004 46808 10013
rect 47676 10047 47728 10056
rect 47676 10013 47685 10047
rect 47685 10013 47719 10047
rect 47719 10013 47728 10047
rect 47676 10004 47728 10013
rect 49240 10047 49292 10056
rect 41236 9936 41288 9988
rect 49240 10013 49249 10047
rect 49249 10013 49283 10047
rect 49283 10013 49292 10047
rect 49240 10004 49292 10013
rect 52552 10047 52604 10056
rect 52552 10013 52561 10047
rect 52561 10013 52595 10047
rect 52595 10013 52604 10047
rect 52552 10004 52604 10013
rect 53380 10047 53432 10056
rect 53380 10013 53389 10047
rect 53389 10013 53423 10047
rect 53423 10013 53432 10047
rect 53380 10004 53432 10013
rect 50068 9936 50120 9988
rect 39764 9868 39816 9920
rect 43720 9911 43772 9920
rect 43720 9877 43729 9911
rect 43729 9877 43763 9911
rect 43763 9877 43772 9911
rect 43720 9868 43772 9877
rect 44180 9911 44232 9920
rect 44180 9877 44189 9911
rect 44189 9877 44223 9911
rect 44223 9877 44232 9911
rect 44180 9868 44232 9877
rect 44640 9868 44692 9920
rect 48872 9868 48924 9920
rect 15398 9766 15450 9818
rect 15462 9766 15514 9818
rect 15526 9766 15578 9818
rect 15590 9766 15642 9818
rect 15654 9766 15706 9818
rect 29846 9766 29898 9818
rect 29910 9766 29962 9818
rect 29974 9766 30026 9818
rect 30038 9766 30090 9818
rect 30102 9766 30154 9818
rect 44294 9766 44346 9818
rect 44358 9766 44410 9818
rect 44422 9766 44474 9818
rect 44486 9766 44538 9818
rect 44550 9766 44602 9818
rect 2964 9664 3016 9716
rect 4804 9664 4856 9716
rect 5632 9664 5684 9716
rect 10048 9664 10100 9716
rect 1768 9571 1820 9580
rect 1768 9537 1777 9571
rect 1777 9537 1811 9571
rect 1811 9537 1820 9571
rect 1768 9528 1820 9537
rect 3148 9596 3200 9648
rect 3056 9528 3108 9580
rect 4068 9596 4120 9648
rect 7288 9596 7340 9648
rect 12256 9664 12308 9716
rect 13452 9664 13504 9716
rect 17776 9664 17828 9716
rect 18420 9664 18472 9716
rect 19340 9664 19392 9716
rect 19708 9664 19760 9716
rect 22008 9664 22060 9716
rect 22376 9707 22428 9716
rect 22376 9673 22385 9707
rect 22385 9673 22419 9707
rect 22419 9673 22428 9707
rect 22376 9664 22428 9673
rect 22560 9664 22612 9716
rect 24400 9664 24452 9716
rect 24860 9707 24912 9716
rect 24860 9673 24869 9707
rect 24869 9673 24903 9707
rect 24903 9673 24912 9707
rect 24860 9664 24912 9673
rect 27160 9664 27212 9716
rect 27988 9707 28040 9716
rect 27988 9673 27997 9707
rect 27997 9673 28031 9707
rect 28031 9673 28040 9707
rect 27988 9664 28040 9673
rect 30840 9664 30892 9716
rect 32312 9707 32364 9716
rect 32312 9673 32321 9707
rect 32321 9673 32355 9707
rect 32355 9673 32364 9707
rect 32312 9664 32364 9673
rect 32496 9664 32548 9716
rect 34152 9664 34204 9716
rect 11244 9596 11296 9648
rect 14096 9596 14148 9648
rect 14924 9639 14976 9648
rect 14924 9605 14933 9639
rect 14933 9605 14967 9639
rect 14967 9605 14976 9639
rect 14924 9596 14976 9605
rect 16212 9596 16264 9648
rect 3516 9571 3568 9580
rect 3516 9537 3525 9571
rect 3525 9537 3559 9571
rect 3559 9537 3568 9571
rect 3516 9528 3568 9537
rect 3884 9528 3936 9580
rect 5080 9528 5132 9580
rect 6460 9528 6512 9580
rect 7840 9571 7892 9580
rect 2780 9460 2832 9512
rect 4528 9460 4580 9512
rect 7840 9537 7849 9571
rect 7849 9537 7883 9571
rect 7883 9537 7892 9571
rect 7840 9528 7892 9537
rect 8760 9571 8812 9580
rect 8760 9537 8769 9571
rect 8769 9537 8803 9571
rect 8803 9537 8812 9571
rect 8760 9528 8812 9537
rect 9864 9528 9916 9580
rect 10692 9571 10744 9580
rect 10692 9537 10701 9571
rect 10701 9537 10735 9571
rect 10735 9537 10744 9571
rect 17316 9596 17368 9648
rect 10692 9528 10744 9537
rect 17408 9571 17460 9580
rect 17408 9537 17417 9571
rect 17417 9537 17451 9571
rect 17451 9537 17460 9571
rect 17408 9528 17460 9537
rect 20076 9528 20128 9580
rect 20904 9571 20956 9580
rect 20904 9537 20913 9571
rect 20913 9537 20947 9571
rect 20947 9537 20956 9571
rect 20904 9528 20956 9537
rect 23480 9596 23532 9648
rect 23296 9528 23348 9580
rect 25228 9571 25280 9580
rect 6828 9460 6880 9512
rect 7932 9460 7984 9512
rect 5080 9392 5132 9444
rect 7380 9392 7432 9444
rect 10968 9460 11020 9512
rect 12716 9503 12768 9512
rect 12716 9469 12725 9503
rect 12725 9469 12759 9503
rect 12759 9469 12768 9503
rect 12716 9460 12768 9469
rect 14556 9503 14608 9512
rect 14556 9469 14565 9503
rect 14565 9469 14599 9503
rect 14599 9469 14608 9503
rect 14556 9460 14608 9469
rect 15384 9503 15436 9512
rect 15384 9469 15393 9503
rect 15393 9469 15427 9503
rect 15427 9469 15436 9503
rect 15384 9460 15436 9469
rect 15476 9460 15528 9512
rect 16948 9460 17000 9512
rect 18972 9460 19024 9512
rect 5632 9324 5684 9376
rect 6736 9324 6788 9376
rect 7932 9324 7984 9376
rect 14188 9392 14240 9444
rect 9772 9324 9824 9376
rect 10600 9324 10652 9376
rect 14372 9324 14424 9376
rect 15200 9392 15252 9444
rect 16488 9392 16540 9444
rect 17132 9392 17184 9444
rect 19616 9324 19668 9376
rect 19892 9324 19944 9376
rect 20260 9324 20312 9376
rect 22100 9460 22152 9512
rect 22468 9460 22520 9512
rect 23020 9392 23072 9444
rect 25228 9537 25237 9571
rect 25237 9537 25271 9571
rect 25271 9537 25280 9571
rect 25228 9528 25280 9537
rect 26056 9571 26108 9580
rect 26056 9537 26065 9571
rect 26065 9537 26099 9571
rect 26099 9537 26108 9571
rect 26056 9528 26108 9537
rect 26240 9571 26292 9580
rect 26240 9537 26249 9571
rect 26249 9537 26283 9571
rect 26283 9537 26292 9571
rect 26240 9528 26292 9537
rect 26332 9528 26384 9580
rect 28448 9571 28500 9580
rect 28448 9537 28457 9571
rect 28457 9537 28491 9571
rect 28491 9537 28500 9571
rect 28448 9528 28500 9537
rect 26976 9503 27028 9512
rect 26976 9469 26985 9503
rect 26985 9469 27019 9503
rect 27019 9469 27028 9503
rect 26976 9460 27028 9469
rect 22284 9324 22336 9376
rect 25044 9324 25096 9376
rect 25688 9324 25740 9376
rect 29000 9528 29052 9580
rect 30564 9596 30616 9648
rect 31760 9596 31812 9648
rect 29552 9571 29604 9580
rect 29552 9537 29561 9571
rect 29561 9537 29595 9571
rect 29595 9537 29604 9571
rect 29552 9528 29604 9537
rect 29644 9528 29696 9580
rect 30748 9571 30800 9580
rect 28816 9503 28868 9512
rect 28816 9469 28825 9503
rect 28825 9469 28859 9503
rect 28859 9469 28868 9503
rect 28816 9460 28868 9469
rect 30748 9537 30757 9571
rect 30757 9537 30791 9571
rect 30791 9537 30800 9571
rect 30748 9528 30800 9537
rect 31576 9528 31628 9580
rect 32956 9528 33008 9580
rect 34980 9571 35032 9580
rect 34980 9537 34989 9571
rect 34989 9537 35023 9571
rect 35023 9537 35032 9571
rect 34980 9528 35032 9537
rect 35072 9528 35124 9580
rect 37372 9664 37424 9716
rect 36452 9571 36504 9580
rect 32772 9503 32824 9512
rect 28816 9324 28868 9376
rect 31300 9392 31352 9444
rect 30012 9324 30064 9376
rect 30288 9367 30340 9376
rect 30288 9333 30297 9367
rect 30297 9333 30331 9367
rect 30331 9333 30340 9367
rect 30288 9324 30340 9333
rect 31116 9324 31168 9376
rect 32772 9469 32781 9503
rect 32781 9469 32815 9503
rect 32815 9469 32824 9503
rect 32772 9460 32824 9469
rect 36452 9537 36461 9571
rect 36461 9537 36495 9571
rect 36495 9537 36504 9571
rect 36452 9528 36504 9537
rect 38016 9664 38068 9716
rect 38108 9664 38160 9716
rect 38660 9596 38712 9648
rect 42984 9664 43036 9716
rect 46480 9707 46532 9716
rect 46480 9673 46489 9707
rect 46489 9673 46523 9707
rect 46523 9673 46532 9707
rect 46480 9664 46532 9673
rect 47676 9664 47728 9716
rect 38568 9571 38620 9580
rect 38568 9537 38577 9571
rect 38577 9537 38611 9571
rect 38611 9537 38620 9571
rect 38568 9528 38620 9537
rect 37372 9460 37424 9512
rect 39948 9571 40000 9580
rect 39948 9537 39957 9571
rect 39957 9537 39991 9571
rect 39991 9537 40000 9571
rect 39948 9528 40000 9537
rect 40224 9571 40276 9580
rect 40224 9537 40233 9571
rect 40233 9537 40267 9571
rect 40267 9537 40276 9571
rect 40224 9528 40276 9537
rect 40316 9528 40368 9580
rect 41236 9503 41288 9512
rect 41236 9469 41245 9503
rect 41245 9469 41279 9503
rect 41279 9469 41288 9503
rect 41236 9460 41288 9469
rect 38108 9392 38160 9444
rect 38844 9324 38896 9376
rect 42156 9528 42208 9580
rect 44180 9596 44232 9648
rect 45468 9596 45520 9648
rect 50528 9639 50580 9648
rect 44640 9571 44692 9580
rect 44640 9537 44649 9571
rect 44649 9537 44683 9571
rect 44683 9537 44692 9571
rect 44640 9528 44692 9537
rect 45008 9528 45060 9580
rect 50528 9605 50537 9639
rect 50537 9605 50571 9639
rect 50571 9605 50580 9639
rect 50528 9596 50580 9605
rect 46664 9571 46716 9580
rect 46664 9537 46673 9571
rect 46673 9537 46707 9571
rect 46707 9537 46716 9571
rect 46664 9528 46716 9537
rect 42432 9503 42484 9512
rect 42432 9469 42441 9503
rect 42441 9469 42475 9503
rect 42475 9469 42484 9503
rect 42432 9460 42484 9469
rect 48136 9528 48188 9580
rect 46756 9392 46808 9444
rect 50068 9571 50120 9580
rect 50068 9537 50077 9571
rect 50077 9537 50111 9571
rect 50111 9537 50120 9571
rect 53380 9596 53432 9648
rect 50068 9528 50120 9537
rect 51264 9528 51316 9580
rect 52000 9571 52052 9580
rect 52000 9537 52009 9571
rect 52009 9537 52043 9571
rect 52043 9537 52052 9571
rect 52000 9528 52052 9537
rect 48964 9503 49016 9512
rect 48964 9469 48973 9503
rect 48973 9469 49007 9503
rect 49007 9469 49016 9503
rect 48964 9460 49016 9469
rect 49700 9460 49752 9512
rect 50528 9460 50580 9512
rect 51448 9460 51500 9512
rect 52276 9460 52328 9512
rect 42800 9324 42852 9376
rect 43720 9324 43772 9376
rect 43996 9324 44048 9376
rect 50528 9324 50580 9376
rect 52552 9324 52604 9376
rect 8174 9222 8226 9274
rect 8238 9222 8290 9274
rect 8302 9222 8354 9274
rect 8366 9222 8418 9274
rect 8430 9222 8482 9274
rect 22622 9222 22674 9274
rect 22686 9222 22738 9274
rect 22750 9222 22802 9274
rect 22814 9222 22866 9274
rect 22878 9222 22930 9274
rect 37070 9222 37122 9274
rect 37134 9222 37186 9274
rect 37198 9222 37250 9274
rect 37262 9222 37314 9274
rect 37326 9222 37378 9274
rect 51518 9222 51570 9274
rect 51582 9222 51634 9274
rect 51646 9222 51698 9274
rect 51710 9222 51762 9274
rect 51774 9222 51826 9274
rect 3516 9120 3568 9172
rect 4252 9120 4304 9172
rect 8760 9120 8812 9172
rect 10692 9120 10744 9172
rect 12256 9163 12308 9172
rect 12256 9129 12265 9163
rect 12265 9129 12299 9163
rect 12299 9129 12308 9163
rect 12256 9120 12308 9129
rect 14556 9120 14608 9172
rect 18236 9120 18288 9172
rect 3884 9052 3936 9104
rect 2412 8984 2464 9036
rect 2964 8984 3016 9036
rect 3424 8984 3476 9036
rect 4068 8984 4120 9036
rect 1952 8916 2004 8968
rect 3056 8959 3108 8968
rect 3056 8925 3065 8959
rect 3065 8925 3099 8959
rect 3099 8925 3108 8959
rect 3056 8916 3108 8925
rect 3792 8916 3844 8968
rect 4896 8959 4948 8968
rect 4896 8925 4905 8959
rect 4905 8925 4939 8959
rect 4939 8925 4948 8959
rect 4896 8916 4948 8925
rect 6092 8959 6144 8968
rect 6092 8925 6101 8959
rect 6101 8925 6135 8959
rect 6135 8925 6144 8959
rect 6092 8916 6144 8925
rect 6736 8959 6788 8968
rect 6736 8925 6745 8959
rect 6745 8925 6779 8959
rect 6779 8925 6788 8959
rect 6736 8916 6788 8925
rect 8024 9052 8076 9104
rect 15568 9052 15620 9104
rect 16488 9052 16540 9104
rect 7380 9027 7432 9036
rect 7380 8993 7389 9027
rect 7389 8993 7423 9027
rect 7423 8993 7432 9027
rect 7380 8984 7432 8993
rect 7564 8916 7616 8968
rect 10600 8959 10652 8968
rect 4528 8848 4580 8900
rect 10600 8925 10609 8959
rect 10609 8925 10643 8959
rect 10643 8925 10652 8959
rect 10600 8916 10652 8925
rect 3332 8780 3384 8832
rect 7564 8780 7616 8832
rect 9772 8780 9824 8832
rect 10600 8780 10652 8832
rect 16672 9027 16724 9036
rect 16672 8993 16681 9027
rect 16681 8993 16715 9027
rect 16715 8993 16724 9027
rect 16672 8984 16724 8993
rect 11428 8916 11480 8968
rect 11520 8959 11572 8968
rect 11520 8925 11529 8959
rect 11529 8925 11563 8959
rect 11563 8925 11572 8959
rect 12716 8959 12768 8968
rect 11520 8916 11572 8925
rect 12716 8925 12725 8959
rect 12725 8925 12759 8959
rect 12759 8925 12768 8959
rect 12716 8916 12768 8925
rect 13268 8916 13320 8968
rect 13452 8916 13504 8968
rect 14464 8959 14516 8968
rect 13820 8848 13872 8900
rect 14464 8925 14473 8959
rect 14473 8925 14507 8959
rect 14507 8925 14516 8959
rect 14464 8916 14516 8925
rect 14832 8916 14884 8968
rect 16396 8916 16448 8968
rect 17040 8916 17092 8968
rect 20076 9052 20128 9104
rect 17408 8959 17460 8968
rect 14924 8848 14976 8900
rect 17408 8925 17417 8959
rect 17417 8925 17451 8959
rect 17451 8925 17460 8959
rect 17408 8916 17460 8925
rect 19616 8959 19668 8968
rect 19616 8925 19625 8959
rect 19625 8925 19659 8959
rect 19659 8925 19668 8959
rect 19616 8916 19668 8925
rect 19708 8916 19760 8968
rect 20720 9120 20772 9172
rect 21916 9120 21968 9172
rect 26332 9163 26384 9172
rect 21824 9095 21876 9104
rect 21824 9061 21833 9095
rect 21833 9061 21867 9095
rect 21867 9061 21876 9095
rect 21824 9052 21876 9061
rect 20260 8984 20312 9036
rect 20444 8959 20496 8968
rect 20444 8925 20453 8959
rect 20453 8925 20487 8959
rect 20487 8925 20496 8959
rect 20444 8916 20496 8925
rect 21640 8959 21692 8968
rect 21640 8925 21649 8959
rect 21649 8925 21683 8959
rect 21683 8925 21692 8959
rect 21640 8916 21692 8925
rect 25688 9095 25740 9104
rect 22284 9027 22336 9036
rect 22284 8993 22293 9027
rect 22293 8993 22327 9027
rect 22327 8993 22336 9027
rect 22284 8984 22336 8993
rect 24400 8984 24452 9036
rect 20076 8848 20128 8900
rect 20720 8848 20772 8900
rect 11796 8780 11848 8832
rect 13452 8823 13504 8832
rect 13452 8789 13461 8823
rect 13461 8789 13495 8823
rect 13495 8789 13504 8823
rect 13452 8780 13504 8789
rect 13544 8780 13596 8832
rect 15476 8780 15528 8832
rect 15568 8780 15620 8832
rect 16212 8780 16264 8832
rect 21824 8848 21876 8900
rect 24860 8959 24912 8968
rect 24860 8925 24869 8959
rect 24869 8925 24903 8959
rect 24903 8925 24912 8959
rect 24860 8916 24912 8925
rect 21180 8823 21232 8832
rect 21180 8789 21189 8823
rect 21189 8789 21223 8823
rect 21223 8789 21232 8823
rect 21180 8780 21232 8789
rect 21272 8780 21324 8832
rect 23296 8823 23348 8832
rect 23296 8789 23305 8823
rect 23305 8789 23339 8823
rect 23339 8789 23348 8823
rect 23296 8780 23348 8789
rect 23480 8780 23532 8832
rect 23664 8780 23716 8832
rect 23940 8780 23992 8832
rect 25688 9061 25697 9095
rect 25697 9061 25731 9095
rect 25731 9061 25740 9095
rect 25688 9052 25740 9061
rect 26332 9129 26341 9163
rect 26341 9129 26375 9163
rect 26375 9129 26384 9163
rect 26332 9120 26384 9129
rect 30748 9120 30800 9172
rect 31576 9163 31628 9172
rect 31576 9129 31585 9163
rect 31585 9129 31619 9163
rect 31619 9129 31628 9163
rect 31576 9120 31628 9129
rect 32956 9163 33008 9172
rect 32956 9129 32965 9163
rect 32965 9129 32999 9163
rect 32999 9129 33008 9163
rect 32956 9120 33008 9129
rect 33048 9120 33100 9172
rect 35532 9120 35584 9172
rect 37556 9120 37608 9172
rect 38568 9120 38620 9172
rect 38752 9120 38804 9172
rect 42156 9163 42208 9172
rect 26976 8984 27028 9036
rect 27068 8916 27120 8968
rect 27988 8959 28040 8968
rect 27988 8925 27997 8959
rect 27997 8925 28031 8959
rect 28031 8925 28040 8959
rect 27988 8916 28040 8925
rect 28172 8959 28224 8968
rect 28172 8925 28181 8959
rect 28181 8925 28215 8959
rect 28215 8925 28224 8959
rect 28172 8916 28224 8925
rect 28816 8959 28868 8968
rect 25044 8848 25096 8900
rect 25964 8848 26016 8900
rect 26240 8848 26292 8900
rect 26976 8891 27028 8900
rect 26976 8857 26985 8891
rect 26985 8857 27019 8891
rect 27019 8857 27028 8891
rect 26976 8848 27028 8857
rect 27160 8891 27212 8900
rect 27160 8857 27169 8891
rect 27169 8857 27203 8891
rect 27203 8857 27212 8891
rect 27160 8848 27212 8857
rect 28816 8925 28825 8959
rect 28825 8925 28859 8959
rect 28859 8925 28868 8959
rect 28816 8916 28868 8925
rect 29460 8848 29512 8900
rect 27436 8780 27488 8832
rect 29184 8780 29236 8832
rect 29552 8780 29604 8832
rect 30012 8780 30064 8832
rect 30564 8916 30616 8968
rect 32772 9052 32824 9104
rect 33600 9052 33652 9104
rect 36360 9052 36412 9104
rect 36452 9052 36504 9104
rect 38844 9052 38896 9104
rect 39764 9052 39816 9104
rect 42156 9129 42165 9163
rect 42165 9129 42199 9163
rect 42199 9129 42208 9163
rect 42156 9120 42208 9129
rect 42800 9120 42852 9172
rect 34888 8984 34940 9036
rect 30656 8848 30708 8900
rect 31392 8959 31444 8968
rect 31392 8925 31401 8959
rect 31401 8925 31435 8959
rect 31435 8925 31444 8959
rect 31392 8916 31444 8925
rect 33232 8916 33284 8968
rect 33324 8916 33376 8968
rect 35256 8959 35308 8968
rect 35256 8925 35265 8959
rect 35265 8925 35299 8959
rect 35299 8925 35308 8959
rect 35256 8916 35308 8925
rect 36268 8916 36320 8968
rect 36176 8848 36228 8900
rect 37464 8916 37516 8968
rect 40132 8984 40184 9036
rect 46664 9120 46716 9172
rect 48136 9163 48188 9172
rect 48136 9129 48145 9163
rect 48145 9129 48179 9163
rect 48179 9129 48188 9163
rect 48136 9120 48188 9129
rect 48228 9120 48280 9172
rect 51264 9163 51316 9172
rect 50528 9095 50580 9104
rect 50528 9061 50537 9095
rect 50537 9061 50571 9095
rect 50571 9061 50580 9095
rect 50528 9052 50580 9061
rect 33416 8780 33468 8832
rect 36912 8780 36964 8832
rect 37832 8780 37884 8832
rect 39672 8916 39724 8968
rect 40316 8916 40368 8968
rect 41328 8959 41380 8968
rect 39028 8848 39080 8900
rect 41328 8925 41337 8959
rect 41337 8925 41371 8959
rect 41371 8925 41380 8959
rect 41328 8916 41380 8925
rect 43444 8916 43496 8968
rect 43628 8959 43680 8968
rect 43628 8925 43637 8959
rect 43637 8925 43671 8959
rect 43671 8925 43680 8959
rect 43628 8916 43680 8925
rect 44272 8959 44324 8968
rect 44272 8925 44281 8959
rect 44281 8925 44315 8959
rect 44315 8925 44324 8959
rect 44272 8916 44324 8925
rect 46388 8959 46440 8968
rect 46388 8925 46397 8959
rect 46397 8925 46431 8959
rect 46431 8925 46440 8959
rect 46388 8916 46440 8925
rect 46664 8959 46716 8968
rect 46664 8925 46673 8959
rect 46673 8925 46707 8959
rect 46707 8925 46716 8959
rect 46664 8916 46716 8925
rect 42432 8848 42484 8900
rect 45468 8848 45520 8900
rect 48228 8916 48280 8968
rect 48412 8848 48464 8900
rect 48872 8959 48924 8968
rect 48872 8925 48881 8959
rect 48881 8925 48915 8959
rect 48915 8925 48924 8959
rect 48872 8916 48924 8925
rect 51264 9129 51273 9163
rect 51273 9129 51307 9163
rect 51307 9129 51316 9163
rect 51264 9120 51316 9129
rect 52276 8984 52328 9036
rect 50344 8848 50396 8900
rect 40132 8780 40184 8832
rect 40316 8780 40368 8832
rect 41144 8780 41196 8832
rect 41696 8780 41748 8832
rect 41880 8780 41932 8832
rect 46296 8780 46348 8832
rect 50712 8891 50764 8900
rect 50712 8857 50721 8891
rect 50721 8857 50755 8891
rect 50755 8857 50764 8891
rect 50712 8848 50764 8857
rect 51540 8916 51592 8968
rect 52092 8916 52144 8968
rect 53380 8916 53432 8968
rect 54116 8959 54168 8968
rect 54116 8925 54125 8959
rect 54125 8925 54159 8959
rect 54159 8925 54168 8959
rect 54116 8916 54168 8925
rect 51172 8780 51224 8832
rect 15398 8678 15450 8730
rect 15462 8678 15514 8730
rect 15526 8678 15578 8730
rect 15590 8678 15642 8730
rect 15654 8678 15706 8730
rect 29846 8678 29898 8730
rect 29910 8678 29962 8730
rect 29974 8678 30026 8730
rect 30038 8678 30090 8730
rect 30102 8678 30154 8730
rect 44294 8678 44346 8730
rect 44358 8678 44410 8730
rect 44422 8678 44474 8730
rect 44486 8678 44538 8730
rect 44550 8678 44602 8730
rect 4712 8619 4764 8628
rect 4712 8585 4721 8619
rect 4721 8585 4755 8619
rect 4755 8585 4764 8619
rect 4712 8576 4764 8585
rect 6460 8576 6512 8628
rect 7932 8576 7984 8628
rect 2320 8508 2372 8560
rect 2596 8508 2648 8560
rect 4988 8508 5040 8560
rect 10784 8576 10836 8628
rect 11336 8576 11388 8628
rect 13544 8576 13596 8628
rect 14464 8576 14516 8628
rect 17408 8576 17460 8628
rect 2044 8440 2096 8492
rect 3516 8483 3568 8492
rect 3516 8449 3525 8483
rect 3525 8449 3559 8483
rect 3559 8449 3568 8483
rect 3516 8440 3568 8449
rect 4344 8483 4396 8492
rect 4344 8449 4353 8483
rect 4353 8449 4387 8483
rect 4387 8449 4396 8483
rect 4344 8440 4396 8449
rect 4528 8483 4580 8492
rect 4528 8449 4537 8483
rect 4537 8449 4571 8483
rect 4571 8449 4580 8483
rect 4528 8440 4580 8449
rect 5816 8483 5868 8492
rect 5816 8449 5825 8483
rect 5825 8449 5859 8483
rect 5859 8449 5868 8483
rect 5816 8440 5868 8449
rect 2780 8372 2832 8424
rect 3424 8372 3476 8424
rect 5448 8372 5500 8424
rect 1400 8304 1452 8356
rect 1860 8304 1912 8356
rect 4252 8304 4304 8356
rect 8208 8483 8260 8492
rect 1584 8236 1636 8288
rect 5724 8236 5776 8288
rect 5816 8236 5868 8288
rect 8208 8449 8217 8483
rect 8217 8449 8251 8483
rect 8251 8449 8260 8483
rect 8208 8440 8260 8449
rect 9496 8508 9548 8560
rect 10324 8483 10376 8492
rect 10324 8449 10333 8483
rect 10333 8449 10367 8483
rect 10367 8449 10376 8483
rect 10324 8440 10376 8449
rect 10416 8440 10468 8492
rect 7380 8279 7432 8288
rect 7380 8245 7389 8279
rect 7389 8245 7423 8279
rect 7423 8245 7432 8279
rect 7380 8236 7432 8245
rect 7748 8236 7800 8288
rect 8392 8304 8444 8356
rect 11152 8440 11204 8492
rect 11244 8440 11296 8492
rect 10876 8372 10928 8424
rect 11796 8483 11848 8492
rect 11796 8449 11805 8483
rect 11805 8449 11839 8483
rect 11839 8449 11848 8483
rect 11796 8440 11848 8449
rect 14924 8508 14976 8560
rect 16672 8508 16724 8560
rect 17224 8508 17276 8560
rect 20260 8508 20312 8560
rect 10968 8304 11020 8356
rect 11244 8236 11296 8288
rect 11796 8236 11848 8288
rect 12440 8236 12492 8288
rect 14648 8440 14700 8492
rect 15108 8483 15160 8492
rect 15108 8449 15117 8483
rect 15117 8449 15151 8483
rect 15151 8449 15160 8483
rect 15108 8440 15160 8449
rect 15200 8440 15252 8492
rect 16396 8440 16448 8492
rect 14004 8372 14056 8424
rect 17040 8483 17092 8492
rect 17040 8449 17049 8483
rect 17049 8449 17083 8483
rect 17083 8449 17092 8483
rect 17040 8440 17092 8449
rect 19432 8483 19484 8492
rect 16948 8372 17000 8424
rect 17776 8372 17828 8424
rect 18236 8372 18288 8424
rect 19432 8449 19441 8483
rect 19441 8449 19475 8483
rect 19475 8449 19484 8483
rect 19432 8440 19484 8449
rect 19892 8440 19944 8492
rect 21272 8576 21324 8628
rect 21640 8576 21692 8628
rect 23296 8576 23348 8628
rect 25228 8576 25280 8628
rect 26148 8576 26200 8628
rect 27068 8619 27120 8628
rect 27068 8585 27077 8619
rect 27077 8585 27111 8619
rect 27111 8585 27120 8619
rect 27068 8576 27120 8585
rect 29000 8576 29052 8628
rect 31484 8619 31536 8628
rect 22100 8508 22152 8560
rect 31484 8585 31493 8619
rect 31493 8585 31527 8619
rect 31527 8585 31536 8619
rect 31484 8576 31536 8585
rect 33232 8619 33284 8628
rect 33232 8585 33241 8619
rect 33241 8585 33275 8619
rect 33275 8585 33284 8619
rect 33232 8576 33284 8585
rect 33324 8576 33376 8628
rect 35072 8576 35124 8628
rect 39028 8619 39080 8628
rect 39028 8585 39037 8619
rect 39037 8585 39071 8619
rect 39071 8585 39080 8619
rect 39028 8576 39080 8585
rect 39672 8619 39724 8628
rect 39672 8585 39681 8619
rect 39681 8585 39715 8619
rect 39715 8585 39724 8619
rect 39672 8576 39724 8585
rect 39948 8576 40000 8628
rect 40776 8576 40828 8628
rect 43444 8619 43496 8628
rect 19708 8372 19760 8424
rect 20076 8415 20128 8424
rect 20076 8381 20085 8415
rect 20085 8381 20119 8415
rect 20119 8381 20128 8415
rect 20076 8372 20128 8381
rect 22284 8483 22336 8492
rect 22284 8449 22293 8483
rect 22293 8449 22327 8483
rect 22327 8449 22336 8483
rect 22284 8440 22336 8449
rect 23664 8483 23716 8492
rect 23664 8449 23673 8483
rect 23673 8449 23707 8483
rect 23707 8449 23716 8483
rect 23664 8440 23716 8449
rect 24216 8440 24268 8492
rect 24400 8440 24452 8492
rect 24676 8440 24728 8492
rect 23296 8372 23348 8424
rect 25964 8483 26016 8492
rect 25964 8449 25973 8483
rect 25973 8449 26007 8483
rect 26007 8449 26016 8483
rect 25964 8440 26016 8449
rect 26148 8440 26200 8492
rect 27344 8483 27396 8492
rect 27344 8449 27353 8483
rect 27353 8449 27387 8483
rect 27387 8449 27396 8483
rect 28356 8483 28408 8492
rect 27344 8440 27396 8449
rect 14096 8236 14148 8288
rect 17684 8279 17736 8288
rect 17684 8245 17693 8279
rect 17693 8245 17727 8279
rect 17727 8245 17736 8279
rect 17684 8236 17736 8245
rect 19248 8279 19300 8288
rect 19248 8245 19257 8279
rect 19257 8245 19291 8279
rect 19291 8245 19300 8279
rect 19248 8236 19300 8245
rect 20444 8236 20496 8288
rect 21916 8304 21968 8356
rect 22008 8304 22060 8356
rect 25228 8304 25280 8356
rect 21272 8236 21324 8288
rect 24584 8236 24636 8288
rect 24676 8236 24728 8288
rect 28356 8449 28365 8483
rect 28365 8449 28399 8483
rect 28399 8449 28408 8483
rect 28356 8440 28408 8449
rect 28448 8304 28500 8356
rect 28632 8440 28684 8492
rect 29736 8372 29788 8424
rect 30288 8440 30340 8492
rect 30840 8483 30892 8492
rect 30840 8449 30849 8483
rect 30849 8449 30883 8483
rect 30883 8449 30892 8483
rect 30840 8440 30892 8449
rect 31024 8483 31076 8492
rect 31024 8449 31033 8483
rect 31033 8449 31067 8483
rect 31067 8449 31076 8483
rect 31024 8440 31076 8449
rect 31208 8440 31260 8492
rect 33048 8440 33100 8492
rect 35072 8483 35124 8492
rect 27804 8236 27856 8288
rect 28172 8236 28224 8288
rect 30288 8304 30340 8356
rect 29184 8279 29236 8288
rect 29184 8245 29193 8279
rect 29193 8245 29227 8279
rect 29227 8245 29236 8279
rect 29184 8236 29236 8245
rect 32864 8372 32916 8424
rect 30564 8304 30616 8356
rect 31208 8304 31260 8356
rect 31392 8304 31444 8356
rect 35072 8449 35081 8483
rect 35081 8449 35115 8483
rect 35115 8449 35124 8483
rect 35072 8440 35124 8449
rect 35256 8508 35308 8560
rect 43444 8585 43453 8619
rect 43453 8585 43487 8619
rect 43487 8585 43496 8619
rect 43444 8576 43496 8585
rect 43628 8576 43680 8628
rect 46664 8576 46716 8628
rect 49240 8576 49292 8628
rect 52000 8576 52052 8628
rect 54116 8576 54168 8628
rect 36268 8440 36320 8492
rect 36360 8440 36412 8492
rect 37832 8483 37884 8492
rect 37832 8449 37841 8483
rect 37841 8449 37875 8483
rect 37875 8449 37884 8483
rect 37832 8440 37884 8449
rect 38108 8440 38160 8492
rect 38752 8483 38804 8492
rect 38752 8449 38761 8483
rect 38761 8449 38795 8483
rect 38795 8449 38804 8483
rect 38752 8440 38804 8449
rect 39488 8483 39540 8492
rect 33600 8415 33652 8424
rect 33600 8381 33609 8415
rect 33609 8381 33643 8415
rect 33643 8381 33652 8415
rect 33600 8372 33652 8381
rect 35532 8415 35584 8424
rect 35532 8381 35541 8415
rect 35541 8381 35575 8415
rect 35575 8381 35584 8415
rect 35532 8372 35584 8381
rect 37556 8372 37608 8424
rect 32220 8236 32272 8288
rect 33968 8236 34020 8288
rect 38384 8304 38436 8356
rect 39488 8449 39497 8483
rect 39497 8449 39531 8483
rect 39531 8449 39540 8483
rect 39488 8440 39540 8449
rect 40316 8483 40368 8492
rect 40316 8449 40325 8483
rect 40325 8449 40359 8483
rect 40359 8449 40368 8483
rect 40316 8440 40368 8449
rect 41144 8483 41196 8492
rect 41144 8449 41153 8483
rect 41153 8449 41187 8483
rect 41187 8449 41196 8483
rect 41144 8440 41196 8449
rect 43352 8440 43404 8492
rect 45284 8440 45336 8492
rect 45468 8440 45520 8492
rect 40776 8372 40828 8424
rect 42524 8372 42576 8424
rect 44640 8372 44692 8424
rect 45100 8372 45152 8424
rect 48228 8508 48280 8560
rect 48412 8551 48464 8560
rect 48412 8517 48421 8551
rect 48421 8517 48455 8551
rect 48455 8517 48464 8551
rect 48412 8508 48464 8517
rect 49148 8508 49200 8560
rect 46756 8483 46808 8492
rect 46756 8449 46765 8483
rect 46765 8449 46799 8483
rect 46799 8449 46808 8483
rect 46756 8440 46808 8449
rect 46848 8483 46900 8492
rect 46848 8449 46857 8483
rect 46857 8449 46891 8483
rect 46891 8449 46900 8483
rect 46848 8440 46900 8449
rect 49332 8440 49384 8492
rect 50068 8483 50120 8492
rect 50068 8449 50077 8483
rect 50077 8449 50111 8483
rect 50111 8449 50120 8483
rect 50068 8440 50120 8449
rect 50804 8483 50856 8492
rect 50804 8449 50813 8483
rect 50813 8449 50847 8483
rect 50847 8449 50856 8483
rect 50804 8440 50856 8449
rect 51540 8440 51592 8492
rect 46940 8372 46992 8424
rect 50712 8372 50764 8424
rect 55772 8440 55824 8492
rect 40224 8236 40276 8288
rect 44180 8304 44232 8356
rect 46848 8304 46900 8356
rect 48320 8304 48372 8356
rect 41880 8279 41932 8288
rect 41880 8245 41889 8279
rect 41889 8245 41923 8279
rect 41923 8245 41932 8279
rect 41880 8236 41932 8245
rect 46940 8236 46992 8288
rect 47584 8279 47636 8288
rect 47584 8245 47593 8279
rect 47593 8245 47627 8279
rect 47627 8245 47636 8279
rect 47584 8236 47636 8245
rect 49148 8236 49200 8288
rect 49700 8304 49752 8356
rect 49884 8347 49936 8356
rect 49884 8313 49893 8347
rect 49893 8313 49927 8347
rect 49927 8313 49936 8347
rect 49884 8304 49936 8313
rect 51356 8304 51408 8356
rect 50620 8279 50672 8288
rect 50620 8245 50629 8279
rect 50629 8245 50663 8279
rect 50663 8245 50672 8279
rect 50620 8236 50672 8245
rect 52920 8304 52972 8356
rect 54392 8372 54444 8424
rect 53196 8304 53248 8356
rect 55312 8304 55364 8356
rect 8174 8134 8226 8186
rect 8238 8134 8290 8186
rect 8302 8134 8354 8186
rect 8366 8134 8418 8186
rect 8430 8134 8482 8186
rect 22622 8134 22674 8186
rect 22686 8134 22738 8186
rect 22750 8134 22802 8186
rect 22814 8134 22866 8186
rect 22878 8134 22930 8186
rect 37070 8134 37122 8186
rect 37134 8134 37186 8186
rect 37198 8134 37250 8186
rect 37262 8134 37314 8186
rect 37326 8134 37378 8186
rect 51518 8134 51570 8186
rect 51582 8134 51634 8186
rect 51646 8134 51698 8186
rect 51710 8134 51762 8186
rect 51774 8134 51826 8186
rect 1768 8032 1820 8084
rect 2044 8032 2096 8084
rect 3516 8032 3568 8084
rect 6184 8032 6236 8084
rect 10508 8032 10560 8084
rect 10968 8032 11020 8084
rect 11704 8032 11756 8084
rect 5540 7964 5592 8016
rect 9220 7964 9272 8016
rect 2964 7896 3016 7948
rect 8300 7896 8352 7948
rect 1860 7871 1912 7880
rect 1860 7837 1869 7871
rect 1869 7837 1903 7871
rect 1903 7837 1912 7871
rect 1860 7828 1912 7837
rect 3516 7828 3568 7880
rect 4344 7871 4396 7880
rect 4344 7837 4353 7871
rect 4353 7837 4387 7871
rect 4387 7837 4396 7871
rect 4344 7828 4396 7837
rect 4988 7871 5040 7880
rect 4988 7837 4997 7871
rect 4997 7837 5031 7871
rect 5031 7837 5040 7871
rect 4988 7828 5040 7837
rect 5816 7828 5868 7880
rect 5908 7871 5960 7880
rect 5908 7837 5917 7871
rect 5917 7837 5951 7871
rect 5951 7837 5960 7871
rect 7564 7871 7616 7880
rect 5908 7828 5960 7837
rect 7564 7837 7573 7871
rect 7573 7837 7607 7871
rect 7607 7837 7616 7871
rect 7564 7828 7616 7837
rect 8024 7828 8076 7880
rect 9220 7871 9272 7880
rect 9220 7837 9229 7871
rect 9229 7837 9263 7871
rect 9263 7837 9272 7871
rect 9220 7828 9272 7837
rect 9864 7828 9916 7880
rect 12440 7828 12492 7880
rect 12624 7871 12676 7880
rect 12624 7837 12633 7871
rect 12633 7837 12667 7871
rect 12667 7837 12676 7871
rect 12624 7828 12676 7837
rect 2044 7735 2096 7744
rect 2044 7701 2053 7735
rect 2053 7701 2087 7735
rect 2087 7701 2096 7735
rect 2044 7692 2096 7701
rect 2504 7735 2556 7744
rect 2504 7701 2513 7735
rect 2513 7701 2547 7735
rect 2547 7701 2556 7735
rect 2504 7692 2556 7701
rect 4712 7692 4764 7744
rect 11704 7760 11756 7812
rect 13544 7828 13596 7880
rect 14648 7964 14700 8016
rect 16212 8032 16264 8084
rect 16580 8075 16632 8084
rect 16580 8041 16589 8075
rect 16589 8041 16623 8075
rect 16623 8041 16632 8075
rect 16580 8032 16632 8041
rect 17868 8032 17920 8084
rect 17684 7964 17736 8016
rect 14832 7939 14884 7948
rect 14832 7905 14841 7939
rect 14841 7905 14875 7939
rect 14875 7905 14884 7939
rect 14832 7896 14884 7905
rect 5356 7692 5408 7744
rect 7380 7692 7432 7744
rect 8208 7692 8260 7744
rect 10048 7692 10100 7744
rect 10692 7735 10744 7744
rect 10692 7701 10701 7735
rect 10701 7701 10735 7735
rect 10735 7701 10744 7735
rect 10692 7692 10744 7701
rect 13268 7692 13320 7744
rect 14648 7760 14700 7812
rect 16396 7828 16448 7880
rect 16948 7871 17000 7880
rect 16948 7837 16957 7871
rect 16957 7837 16991 7871
rect 16991 7837 17000 7871
rect 16948 7828 17000 7837
rect 17132 7828 17184 7880
rect 18420 7828 18472 7880
rect 18788 8032 18840 8084
rect 19524 7964 19576 8016
rect 19800 8032 19852 8084
rect 21088 8032 21140 8084
rect 23020 8032 23072 8084
rect 23664 8032 23716 8084
rect 24860 8032 24912 8084
rect 25964 8032 26016 8084
rect 27620 8032 27672 8084
rect 28448 8075 28500 8084
rect 28448 8041 28457 8075
rect 28457 8041 28491 8075
rect 28491 8041 28500 8075
rect 28448 8032 28500 8041
rect 28724 8075 28776 8084
rect 28724 8041 28733 8075
rect 28733 8041 28767 8075
rect 28767 8041 28776 8075
rect 28724 8032 28776 8041
rect 30656 8032 30708 8084
rect 35072 8075 35124 8084
rect 35072 8041 35081 8075
rect 35081 8041 35115 8075
rect 35115 8041 35124 8075
rect 35072 8032 35124 8041
rect 41328 8032 41380 8084
rect 25780 7964 25832 8016
rect 26056 7964 26108 8016
rect 33232 7964 33284 8016
rect 39488 7964 39540 8016
rect 40224 8007 40276 8016
rect 40224 7973 40233 8007
rect 40233 7973 40267 8007
rect 40267 7973 40276 8007
rect 42524 8032 42576 8084
rect 43352 8032 43404 8084
rect 46296 8075 46348 8084
rect 46296 8041 46305 8075
rect 46305 8041 46339 8075
rect 46339 8041 46348 8075
rect 46296 8032 46348 8041
rect 46388 8032 46440 8084
rect 50804 8032 50856 8084
rect 51172 8075 51224 8084
rect 51172 8041 51181 8075
rect 51181 8041 51215 8075
rect 51215 8041 51224 8075
rect 51172 8032 51224 8041
rect 51356 8032 51408 8084
rect 40224 7964 40276 7973
rect 19708 7896 19760 7948
rect 19248 7871 19300 7880
rect 19248 7837 19257 7871
rect 19257 7837 19291 7871
rect 19291 7837 19300 7871
rect 19248 7828 19300 7837
rect 20168 7828 20220 7880
rect 20904 7828 20956 7880
rect 21272 7871 21324 7880
rect 21272 7837 21281 7871
rect 21281 7837 21315 7871
rect 21315 7837 21324 7871
rect 21272 7828 21324 7837
rect 23020 7896 23072 7948
rect 23296 7896 23348 7948
rect 26424 7939 26476 7948
rect 26424 7905 26433 7939
rect 26433 7905 26467 7939
rect 26467 7905 26476 7939
rect 26424 7896 26476 7905
rect 26976 7896 27028 7948
rect 24584 7871 24636 7880
rect 17960 7760 18012 7812
rect 20260 7760 20312 7812
rect 21180 7760 21232 7812
rect 22376 7760 22428 7812
rect 23480 7760 23532 7812
rect 23756 7803 23808 7812
rect 23756 7769 23765 7803
rect 23765 7769 23799 7803
rect 23799 7769 23808 7803
rect 23756 7760 23808 7769
rect 15200 7692 15252 7744
rect 19524 7692 19576 7744
rect 21640 7735 21692 7744
rect 21640 7701 21649 7735
rect 21649 7701 21683 7735
rect 21683 7701 21692 7735
rect 21640 7692 21692 7701
rect 24584 7837 24593 7871
rect 24593 7837 24627 7871
rect 24627 7837 24636 7871
rect 24584 7828 24636 7837
rect 24768 7871 24820 7880
rect 24768 7837 24777 7871
rect 24777 7837 24811 7871
rect 24811 7837 24820 7871
rect 24768 7828 24820 7837
rect 25964 7828 26016 7880
rect 27436 7828 27488 7880
rect 26792 7760 26844 7812
rect 27620 7828 27672 7880
rect 27804 7871 27856 7880
rect 27804 7837 27813 7871
rect 27813 7837 27847 7871
rect 27847 7837 27856 7871
rect 27804 7828 27856 7837
rect 27896 7871 27948 7880
rect 27896 7837 27905 7871
rect 27905 7837 27939 7871
rect 27939 7837 27948 7871
rect 28908 7871 28960 7880
rect 27896 7828 27948 7837
rect 28908 7837 28917 7871
rect 28917 7837 28951 7871
rect 28951 7837 28960 7871
rect 28908 7828 28960 7837
rect 29736 7828 29788 7880
rect 28724 7760 28776 7812
rect 30380 7760 30432 7812
rect 31300 7828 31352 7880
rect 32220 7871 32272 7880
rect 32220 7837 32229 7871
rect 32229 7837 32263 7871
rect 32263 7837 32272 7871
rect 32220 7828 32272 7837
rect 32864 7871 32916 7880
rect 32864 7837 32873 7871
rect 32873 7837 32907 7871
rect 32907 7837 32916 7871
rect 32864 7828 32916 7837
rect 33416 7828 33468 7880
rect 36176 7896 36228 7948
rect 35256 7828 35308 7880
rect 36636 7871 36688 7880
rect 36636 7837 36645 7871
rect 36645 7837 36679 7871
rect 36679 7837 36688 7871
rect 36636 7828 36688 7837
rect 36912 7828 36964 7880
rect 45284 7939 45336 7948
rect 38844 7871 38896 7880
rect 34888 7803 34940 7812
rect 34888 7769 34897 7803
rect 34897 7769 34931 7803
rect 34931 7769 34940 7803
rect 34888 7760 34940 7769
rect 38108 7760 38160 7812
rect 38844 7837 38853 7871
rect 38853 7837 38887 7871
rect 38887 7837 38896 7871
rect 38844 7828 38896 7837
rect 25228 7692 25280 7744
rect 25780 7692 25832 7744
rect 30748 7692 30800 7744
rect 31576 7692 31628 7744
rect 31852 7735 31904 7744
rect 31852 7701 31861 7735
rect 31861 7701 31895 7735
rect 31895 7701 31904 7735
rect 31852 7692 31904 7701
rect 32036 7692 32088 7744
rect 32312 7692 32364 7744
rect 37464 7692 37516 7744
rect 40408 7803 40460 7812
rect 40408 7769 40417 7803
rect 40417 7769 40451 7803
rect 40451 7769 40460 7803
rect 40408 7760 40460 7769
rect 45284 7905 45293 7939
rect 45293 7905 45327 7939
rect 45327 7905 45336 7939
rect 45284 7896 45336 7905
rect 40592 7828 40644 7880
rect 41696 7871 41748 7880
rect 41696 7837 41705 7871
rect 41705 7837 41739 7871
rect 41739 7837 41748 7871
rect 41696 7828 41748 7837
rect 43076 7871 43128 7880
rect 43076 7837 43085 7871
rect 43085 7837 43119 7871
rect 43119 7837 43128 7871
rect 43076 7828 43128 7837
rect 44180 7871 44232 7880
rect 44180 7837 44189 7871
rect 44189 7837 44223 7871
rect 44223 7837 44232 7871
rect 44180 7828 44232 7837
rect 46020 7828 46072 7880
rect 42892 7803 42944 7812
rect 42892 7769 42901 7803
rect 42901 7769 42935 7803
rect 42935 7769 42944 7803
rect 42892 7760 42944 7769
rect 40224 7692 40276 7744
rect 41420 7692 41472 7744
rect 45376 7760 45428 7812
rect 48320 7896 48372 7948
rect 49332 7964 49384 8016
rect 46940 7871 46992 7880
rect 46940 7837 46949 7871
rect 46949 7837 46983 7871
rect 46983 7837 46992 7871
rect 46940 7828 46992 7837
rect 50068 7896 50120 7948
rect 49148 7828 49200 7880
rect 49332 7828 49384 7880
rect 50344 7828 50396 7880
rect 53104 7828 53156 7880
rect 44640 7692 44692 7744
rect 47584 7692 47636 7744
rect 52460 7760 52512 7812
rect 52184 7735 52236 7744
rect 52184 7701 52193 7735
rect 52193 7701 52227 7735
rect 52227 7701 52236 7735
rect 52184 7692 52236 7701
rect 52736 7735 52788 7744
rect 52736 7701 52745 7735
rect 52745 7701 52779 7735
rect 52779 7701 52788 7735
rect 52736 7692 52788 7701
rect 54208 7692 54260 7744
rect 55312 7735 55364 7744
rect 55312 7701 55321 7735
rect 55321 7701 55355 7735
rect 55355 7701 55364 7735
rect 55312 7692 55364 7701
rect 15398 7590 15450 7642
rect 15462 7590 15514 7642
rect 15526 7590 15578 7642
rect 15590 7590 15642 7642
rect 15654 7590 15706 7642
rect 29846 7590 29898 7642
rect 29910 7590 29962 7642
rect 29974 7590 30026 7642
rect 30038 7590 30090 7642
rect 30102 7590 30154 7642
rect 44294 7590 44346 7642
rect 44358 7590 44410 7642
rect 44422 7590 44474 7642
rect 44486 7590 44538 7642
rect 44550 7590 44602 7642
rect 4252 7488 4304 7540
rect 4344 7488 4396 7540
rect 2044 7420 2096 7472
rect 1584 7395 1636 7404
rect 1584 7361 1593 7395
rect 1593 7361 1627 7395
rect 1627 7361 1636 7395
rect 1584 7352 1636 7361
rect 3424 7395 3476 7404
rect 3424 7361 3433 7395
rect 3433 7361 3467 7395
rect 3467 7361 3476 7395
rect 3424 7352 3476 7361
rect 5448 7420 5500 7472
rect 6276 7352 6328 7404
rect 6368 7352 6420 7404
rect 7748 7488 7800 7540
rect 8208 7488 8260 7540
rect 10692 7488 10744 7540
rect 15384 7488 15436 7540
rect 16948 7488 17000 7540
rect 17684 7531 17736 7540
rect 17684 7497 17693 7531
rect 17693 7497 17727 7531
rect 17727 7497 17736 7531
rect 17684 7488 17736 7497
rect 18420 7488 18472 7540
rect 24308 7488 24360 7540
rect 7564 7420 7616 7472
rect 7380 7395 7432 7404
rect 7380 7361 7389 7395
rect 7389 7361 7423 7395
rect 7423 7361 7432 7395
rect 7380 7352 7432 7361
rect 4160 7284 4212 7336
rect 5816 7284 5868 7336
rect 6000 7284 6052 7336
rect 8024 7327 8076 7336
rect 2964 7216 3016 7268
rect 5448 7216 5500 7268
rect 2228 7191 2280 7200
rect 2228 7157 2237 7191
rect 2237 7157 2271 7191
rect 2271 7157 2280 7191
rect 2228 7148 2280 7157
rect 3056 7191 3108 7200
rect 3056 7157 3065 7191
rect 3065 7157 3099 7191
rect 3099 7157 3108 7191
rect 3056 7148 3108 7157
rect 4160 7191 4212 7200
rect 4160 7157 4169 7191
rect 4169 7157 4203 7191
rect 4203 7157 4212 7191
rect 4160 7148 4212 7157
rect 5356 7148 5408 7200
rect 6736 7148 6788 7200
rect 6920 7148 6972 7200
rect 8024 7293 8033 7327
rect 8033 7293 8067 7327
rect 8067 7293 8076 7327
rect 8024 7284 8076 7293
rect 9496 7327 9548 7336
rect 9496 7293 9505 7327
rect 9505 7293 9539 7327
rect 9539 7293 9548 7327
rect 9496 7284 9548 7293
rect 14004 7420 14056 7472
rect 11796 7284 11848 7336
rect 12992 7352 13044 7404
rect 13820 7352 13872 7404
rect 14096 7395 14148 7404
rect 14096 7361 14105 7395
rect 14105 7361 14139 7395
rect 14139 7361 14148 7395
rect 14096 7352 14148 7361
rect 14188 7395 14240 7404
rect 14188 7361 14197 7395
rect 14197 7361 14231 7395
rect 14231 7361 14240 7395
rect 15384 7395 15436 7404
rect 14188 7352 14240 7361
rect 15384 7361 15393 7395
rect 15393 7361 15427 7395
rect 15427 7361 15436 7395
rect 15384 7352 15436 7361
rect 16212 7352 16264 7404
rect 17040 7352 17092 7404
rect 19248 7420 19300 7472
rect 17960 7352 18012 7404
rect 18328 7395 18380 7404
rect 18328 7361 18337 7395
rect 18337 7361 18371 7395
rect 18371 7361 18380 7395
rect 18328 7352 18380 7361
rect 18420 7352 18472 7404
rect 19432 7352 19484 7404
rect 19616 7395 19668 7404
rect 19616 7361 19625 7395
rect 19625 7361 19659 7395
rect 19659 7361 19668 7395
rect 19616 7352 19668 7361
rect 19708 7352 19760 7404
rect 21456 7352 21508 7404
rect 24584 7420 24636 7472
rect 14924 7284 14976 7336
rect 18972 7284 19024 7336
rect 21824 7284 21876 7336
rect 24308 7395 24360 7404
rect 24308 7361 24317 7395
rect 24317 7361 24351 7395
rect 24351 7361 24360 7395
rect 24308 7352 24360 7361
rect 26240 7488 26292 7540
rect 34980 7488 35032 7540
rect 25228 7352 25280 7404
rect 26056 7395 26108 7404
rect 26056 7361 26065 7395
rect 26065 7361 26099 7395
rect 26099 7361 26108 7395
rect 26056 7352 26108 7361
rect 26240 7352 26292 7404
rect 26884 7352 26936 7404
rect 25044 7327 25096 7336
rect 12072 7216 12124 7268
rect 13728 7216 13780 7268
rect 12532 7191 12584 7200
rect 12532 7157 12541 7191
rect 12541 7157 12575 7191
rect 12575 7157 12584 7191
rect 12532 7148 12584 7157
rect 12900 7148 12952 7200
rect 16304 7148 16356 7200
rect 16396 7148 16448 7200
rect 18420 7148 18472 7200
rect 19064 7148 19116 7200
rect 19156 7191 19208 7200
rect 19156 7157 19165 7191
rect 19165 7157 19199 7191
rect 19199 7157 19208 7191
rect 19156 7148 19208 7157
rect 19616 7148 19668 7200
rect 21916 7191 21968 7200
rect 21916 7157 21925 7191
rect 21925 7157 21959 7191
rect 21959 7157 21968 7191
rect 21916 7148 21968 7157
rect 22284 7216 22336 7268
rect 25044 7293 25053 7327
rect 25053 7293 25087 7327
rect 25087 7293 25096 7327
rect 25044 7284 25096 7293
rect 25136 7327 25188 7336
rect 25136 7293 25145 7327
rect 25145 7293 25179 7327
rect 25179 7293 25188 7327
rect 25136 7284 25188 7293
rect 26792 7284 26844 7336
rect 28356 7284 28408 7336
rect 29000 7395 29052 7404
rect 29000 7361 29009 7395
rect 29009 7361 29043 7395
rect 29043 7361 29052 7395
rect 29000 7352 29052 7361
rect 29644 7352 29696 7404
rect 29828 7284 29880 7336
rect 29736 7216 29788 7268
rect 31852 7352 31904 7404
rect 35992 7420 36044 7472
rect 36360 7420 36412 7472
rect 42432 7488 42484 7540
rect 46020 7531 46072 7540
rect 46020 7497 46029 7531
rect 46029 7497 46063 7531
rect 46063 7497 46072 7531
rect 46020 7488 46072 7497
rect 51172 7488 51224 7540
rect 51448 7488 51500 7540
rect 53104 7531 53156 7540
rect 53104 7497 53113 7531
rect 53113 7497 53147 7531
rect 53147 7497 53156 7531
rect 53104 7488 53156 7497
rect 38936 7420 38988 7472
rect 33968 7395 34020 7404
rect 33968 7361 33977 7395
rect 33977 7361 34011 7395
rect 34011 7361 34020 7395
rect 33968 7352 34020 7361
rect 34612 7395 34664 7404
rect 34612 7361 34621 7395
rect 34621 7361 34655 7395
rect 34655 7361 34664 7395
rect 34612 7352 34664 7361
rect 34704 7352 34756 7404
rect 37464 7395 37516 7404
rect 37464 7361 37473 7395
rect 37473 7361 37507 7395
rect 37507 7361 37516 7395
rect 37464 7352 37516 7361
rect 37556 7395 37608 7404
rect 37556 7361 37565 7395
rect 37565 7361 37599 7395
rect 37599 7361 37608 7395
rect 37556 7352 37608 7361
rect 38660 7352 38712 7404
rect 40592 7420 40644 7472
rect 40684 7395 40736 7404
rect 40684 7361 40693 7395
rect 40693 7361 40727 7395
rect 40727 7361 40736 7395
rect 40684 7352 40736 7361
rect 42892 7352 42944 7404
rect 43996 7420 44048 7472
rect 31576 7284 31628 7336
rect 35256 7327 35308 7336
rect 23296 7148 23348 7200
rect 23940 7148 23992 7200
rect 26332 7148 26384 7200
rect 27252 7148 27304 7200
rect 32312 7216 32364 7268
rect 31300 7148 31352 7200
rect 35256 7293 35265 7327
rect 35265 7293 35299 7327
rect 35299 7293 35308 7327
rect 35256 7284 35308 7293
rect 36820 7284 36872 7336
rect 37924 7284 37976 7336
rect 38936 7327 38988 7336
rect 38936 7293 38945 7327
rect 38945 7293 38979 7327
rect 38979 7293 38988 7327
rect 38936 7284 38988 7293
rect 36636 7216 36688 7268
rect 37740 7216 37792 7268
rect 38108 7259 38160 7268
rect 38108 7225 38117 7259
rect 38117 7225 38151 7259
rect 38151 7225 38160 7259
rect 38108 7216 38160 7225
rect 41420 7259 41472 7268
rect 41420 7225 41429 7259
rect 41429 7225 41463 7259
rect 41463 7225 41472 7259
rect 41420 7216 41472 7225
rect 44640 7284 44692 7336
rect 45008 7284 45060 7336
rect 45376 7395 45428 7404
rect 45376 7361 45385 7395
rect 45385 7361 45419 7395
rect 45419 7361 45428 7395
rect 45376 7352 45428 7361
rect 50344 7395 50396 7404
rect 50344 7361 50353 7395
rect 50353 7361 50387 7395
rect 50387 7361 50396 7395
rect 50344 7352 50396 7361
rect 50620 7395 50672 7404
rect 50620 7361 50629 7395
rect 50629 7361 50663 7395
rect 50663 7361 50672 7395
rect 50620 7352 50672 7361
rect 52092 7395 52144 7404
rect 52092 7361 52101 7395
rect 52101 7361 52135 7395
rect 52135 7361 52144 7395
rect 52092 7352 52144 7361
rect 55864 7420 55916 7472
rect 54208 7395 54260 7404
rect 54208 7361 54217 7395
rect 54217 7361 54251 7395
rect 54251 7361 54260 7395
rect 54208 7352 54260 7361
rect 56232 7352 56284 7404
rect 48044 7327 48096 7336
rect 48044 7293 48053 7327
rect 48053 7293 48087 7327
rect 48087 7293 48096 7327
rect 48044 7284 48096 7293
rect 49240 7284 49292 7336
rect 52368 7284 52420 7336
rect 52828 7284 52880 7336
rect 55588 7284 55640 7336
rect 57520 7284 57572 7336
rect 33600 7148 33652 7200
rect 34888 7148 34940 7200
rect 35900 7148 35952 7200
rect 36176 7148 36228 7200
rect 36912 7148 36964 7200
rect 37464 7148 37516 7200
rect 38752 7148 38804 7200
rect 42892 7148 42944 7200
rect 50068 7216 50120 7268
rect 44180 7148 44232 7200
rect 46848 7191 46900 7200
rect 46848 7157 46857 7191
rect 46857 7157 46891 7191
rect 46891 7157 46900 7191
rect 46848 7148 46900 7157
rect 50712 7148 50764 7200
rect 51264 7148 51316 7200
rect 57796 7148 57848 7200
rect 57980 7191 58032 7200
rect 57980 7157 57989 7191
rect 57989 7157 58023 7191
rect 58023 7157 58032 7191
rect 57980 7148 58032 7157
rect 8174 7046 8226 7098
rect 8238 7046 8290 7098
rect 8302 7046 8354 7098
rect 8366 7046 8418 7098
rect 8430 7046 8482 7098
rect 22622 7046 22674 7098
rect 22686 7046 22738 7098
rect 22750 7046 22802 7098
rect 22814 7046 22866 7098
rect 22878 7046 22930 7098
rect 37070 7046 37122 7098
rect 37134 7046 37186 7098
rect 37198 7046 37250 7098
rect 37262 7046 37314 7098
rect 37326 7046 37378 7098
rect 51518 7046 51570 7098
rect 51582 7046 51634 7098
rect 51646 7046 51698 7098
rect 51710 7046 51762 7098
rect 51774 7046 51826 7098
rect 5816 6944 5868 6996
rect 6184 6944 6236 6996
rect 7380 6944 7432 6996
rect 10600 6944 10652 6996
rect 4712 6876 4764 6928
rect 5356 6876 5408 6928
rect 8024 6876 8076 6928
rect 3700 6808 3752 6860
rect 10876 6808 10928 6860
rect 11796 6944 11848 6996
rect 13728 6944 13780 6996
rect 16304 6944 16356 6996
rect 18420 6944 18472 6996
rect 21824 6987 21876 6996
rect 21824 6953 21833 6987
rect 21833 6953 21867 6987
rect 21867 6953 21876 6987
rect 21824 6944 21876 6953
rect 23296 6987 23348 6996
rect 23296 6953 23305 6987
rect 23305 6953 23339 6987
rect 23339 6953 23348 6987
rect 23296 6944 23348 6953
rect 24032 6944 24084 6996
rect 24400 6944 24452 6996
rect 14372 6876 14424 6928
rect 16396 6876 16448 6928
rect 28816 6944 28868 6996
rect 29736 6987 29788 6996
rect 29736 6953 29745 6987
rect 29745 6953 29779 6987
rect 29779 6953 29788 6987
rect 29736 6944 29788 6953
rect 2136 6740 2188 6792
rect 3148 6740 3200 6792
rect 3516 6740 3568 6792
rect 3976 6740 4028 6792
rect 1860 6672 1912 6724
rect 5356 6740 5408 6792
rect 6552 6740 6604 6792
rect 6736 6783 6788 6792
rect 6736 6749 6745 6783
rect 6745 6749 6779 6783
rect 6779 6749 6788 6783
rect 6736 6740 6788 6749
rect 7288 6740 7340 6792
rect 7932 6740 7984 6792
rect 9496 6783 9548 6792
rect 9496 6749 9505 6783
rect 9505 6749 9539 6783
rect 9539 6749 9548 6783
rect 9496 6740 9548 6749
rect 9680 6740 9732 6792
rect 10324 6715 10376 6724
rect 2596 6647 2648 6656
rect 2596 6613 2605 6647
rect 2605 6613 2639 6647
rect 2639 6613 2648 6647
rect 2596 6604 2648 6613
rect 3148 6604 3200 6656
rect 4712 6604 4764 6656
rect 6000 6604 6052 6656
rect 7380 6647 7432 6656
rect 7380 6613 7389 6647
rect 7389 6613 7423 6647
rect 7423 6613 7432 6647
rect 7380 6604 7432 6613
rect 8024 6604 8076 6656
rect 8760 6604 8812 6656
rect 9128 6604 9180 6656
rect 9220 6604 9272 6656
rect 10324 6681 10333 6715
rect 10333 6681 10367 6715
rect 10367 6681 10376 6715
rect 10324 6672 10376 6681
rect 10508 6740 10560 6792
rect 14924 6808 14976 6860
rect 16948 6851 17000 6860
rect 16948 6817 16957 6851
rect 16957 6817 16991 6851
rect 16991 6817 17000 6851
rect 16948 6808 17000 6817
rect 17684 6808 17736 6860
rect 20260 6808 20312 6860
rect 22284 6851 22336 6860
rect 22284 6817 22293 6851
rect 22293 6817 22327 6851
rect 22327 6817 22336 6851
rect 22284 6808 22336 6817
rect 23388 6808 23440 6860
rect 23572 6808 23624 6860
rect 24032 6808 24084 6860
rect 24124 6808 24176 6860
rect 25136 6808 25188 6860
rect 10692 6672 10744 6724
rect 13544 6783 13596 6792
rect 13544 6749 13553 6783
rect 13553 6749 13587 6783
rect 13587 6749 13596 6783
rect 13544 6740 13596 6749
rect 14096 6783 14148 6792
rect 14096 6749 14105 6783
rect 14105 6749 14139 6783
rect 14139 6749 14148 6783
rect 14096 6740 14148 6749
rect 14648 6740 14700 6792
rect 12256 6672 12308 6724
rect 10600 6604 10652 6656
rect 11428 6604 11480 6656
rect 11520 6604 11572 6656
rect 17132 6740 17184 6792
rect 19524 6783 19576 6792
rect 16580 6672 16632 6724
rect 19524 6749 19533 6783
rect 19533 6749 19567 6783
rect 19567 6749 19576 6783
rect 19524 6740 19576 6749
rect 21640 6783 21692 6792
rect 20076 6672 20128 6724
rect 21640 6749 21649 6783
rect 21649 6749 21683 6783
rect 21683 6749 21692 6783
rect 21640 6740 21692 6749
rect 22560 6783 22612 6792
rect 22560 6749 22569 6783
rect 22569 6749 22603 6783
rect 22603 6749 22612 6783
rect 22560 6740 22612 6749
rect 24860 6740 24912 6792
rect 23572 6672 23624 6724
rect 25228 6672 25280 6724
rect 26056 6876 26108 6928
rect 26424 6876 26476 6928
rect 26976 6919 27028 6928
rect 26976 6885 26985 6919
rect 26985 6885 27019 6919
rect 27019 6885 27028 6919
rect 26976 6876 27028 6885
rect 33416 6944 33468 6996
rect 33600 6944 33652 6996
rect 36176 6944 36228 6996
rect 36360 6987 36412 6996
rect 36360 6953 36369 6987
rect 36369 6953 36403 6987
rect 36403 6953 36412 6987
rect 36360 6944 36412 6953
rect 28724 6851 28776 6860
rect 18236 6604 18288 6656
rect 18420 6604 18472 6656
rect 22100 6604 22152 6656
rect 23296 6604 23348 6656
rect 24032 6604 24084 6656
rect 28724 6817 28733 6851
rect 28733 6817 28767 6851
rect 28767 6817 28776 6851
rect 28724 6808 28776 6817
rect 29000 6783 29052 6792
rect 26424 6672 26476 6724
rect 26700 6672 26752 6724
rect 27436 6672 27488 6724
rect 29000 6749 29009 6783
rect 29009 6749 29043 6783
rect 29043 6749 29052 6783
rect 29000 6740 29052 6749
rect 32220 6876 32272 6928
rect 32036 6851 32088 6860
rect 32036 6817 32045 6851
rect 32045 6817 32079 6851
rect 32079 6817 32088 6851
rect 32036 6808 32088 6817
rect 30564 6740 30616 6792
rect 28908 6672 28960 6724
rect 30380 6672 30432 6724
rect 31852 6740 31904 6792
rect 32588 6876 32640 6928
rect 33140 6876 33192 6928
rect 37648 6944 37700 6996
rect 37740 6944 37792 6996
rect 42892 6944 42944 6996
rect 43076 6944 43128 6996
rect 48596 6987 48648 6996
rect 35808 6851 35860 6860
rect 35808 6817 35817 6851
rect 35817 6817 35851 6851
rect 35851 6817 35860 6851
rect 35808 6808 35860 6817
rect 41604 6919 41656 6928
rect 41604 6885 41613 6919
rect 41613 6885 41647 6919
rect 41647 6885 41656 6919
rect 41604 6876 41656 6885
rect 48596 6953 48605 6987
rect 48605 6953 48639 6987
rect 48639 6953 48648 6987
rect 48596 6944 48648 6953
rect 49240 6944 49292 6996
rect 51264 6987 51316 6996
rect 51264 6953 51273 6987
rect 51273 6953 51307 6987
rect 51307 6953 51316 6987
rect 51264 6944 51316 6953
rect 52368 6944 52420 6996
rect 55864 6987 55916 6996
rect 31392 6672 31444 6724
rect 32496 6740 32548 6792
rect 33876 6740 33928 6792
rect 36820 6783 36872 6792
rect 32956 6715 33008 6724
rect 29000 6604 29052 6656
rect 29460 6604 29512 6656
rect 29828 6604 29880 6656
rect 32956 6681 32965 6715
rect 32965 6681 32999 6715
rect 32999 6681 33008 6715
rect 32956 6672 33008 6681
rect 34428 6672 34480 6724
rect 36820 6749 36829 6783
rect 36829 6749 36863 6783
rect 36863 6749 36872 6783
rect 36820 6740 36872 6749
rect 37096 6783 37148 6792
rect 37096 6749 37105 6783
rect 37105 6749 37139 6783
rect 37139 6749 37148 6783
rect 37096 6740 37148 6749
rect 37280 6740 37332 6792
rect 38752 6808 38804 6860
rect 38844 6808 38896 6860
rect 40040 6808 40092 6860
rect 52276 6876 52328 6928
rect 55864 6953 55873 6987
rect 55873 6953 55907 6987
rect 55907 6953 55916 6987
rect 55864 6944 55916 6953
rect 45008 6851 45060 6860
rect 45008 6817 45017 6851
rect 45017 6817 45051 6851
rect 45051 6817 45060 6851
rect 45008 6808 45060 6817
rect 52460 6808 52512 6860
rect 54116 6808 54168 6860
rect 57796 6851 57848 6860
rect 57796 6817 57805 6851
rect 57805 6817 57839 6851
rect 57839 6817 57848 6851
rect 57796 6808 57848 6817
rect 38384 6783 38436 6792
rect 38384 6749 38393 6783
rect 38393 6749 38427 6783
rect 38427 6749 38436 6783
rect 38384 6740 38436 6749
rect 38476 6740 38528 6792
rect 41696 6740 41748 6792
rect 42432 6783 42484 6792
rect 42432 6749 42441 6783
rect 42441 6749 42475 6783
rect 42475 6749 42484 6783
rect 42432 6740 42484 6749
rect 43996 6740 44048 6792
rect 46572 6783 46624 6792
rect 32404 6604 32456 6656
rect 33232 6604 33284 6656
rect 34704 6604 34756 6656
rect 37464 6672 37516 6724
rect 35808 6604 35860 6656
rect 35992 6647 36044 6656
rect 35992 6613 36001 6647
rect 36001 6613 36035 6647
rect 36035 6613 36044 6647
rect 35992 6604 36044 6613
rect 36820 6604 36872 6656
rect 38936 6672 38988 6724
rect 40408 6715 40460 6724
rect 40408 6681 40417 6715
rect 40417 6681 40451 6715
rect 40451 6681 40460 6715
rect 40408 6672 40460 6681
rect 40868 6672 40920 6724
rect 38660 6604 38712 6656
rect 39304 6604 39356 6656
rect 41788 6672 41840 6724
rect 42616 6715 42668 6724
rect 42616 6681 42625 6715
rect 42625 6681 42659 6715
rect 42659 6681 42668 6715
rect 42616 6672 42668 6681
rect 43352 6672 43404 6724
rect 46572 6749 46581 6783
rect 46581 6749 46615 6783
rect 46615 6749 46624 6783
rect 46572 6740 46624 6749
rect 46848 6783 46900 6792
rect 46848 6749 46857 6783
rect 46857 6749 46891 6783
rect 46891 6749 46900 6783
rect 46848 6740 46900 6749
rect 41972 6604 42024 6656
rect 42708 6604 42760 6656
rect 48596 6672 48648 6724
rect 48044 6647 48096 6656
rect 48044 6613 48053 6647
rect 48053 6613 48087 6647
rect 48087 6613 48096 6647
rect 48044 6604 48096 6613
rect 49332 6783 49384 6792
rect 49332 6749 49341 6783
rect 49341 6749 49375 6783
rect 49375 6749 49384 6783
rect 49332 6740 49384 6749
rect 50528 6783 50580 6792
rect 50528 6749 50537 6783
rect 50537 6749 50571 6783
rect 50571 6749 50580 6783
rect 50528 6740 50580 6749
rect 52828 6740 52880 6792
rect 57520 6783 57572 6792
rect 52184 6672 52236 6724
rect 55680 6715 55732 6724
rect 55680 6681 55689 6715
rect 55689 6681 55723 6715
rect 55723 6681 55732 6715
rect 55680 6672 55732 6681
rect 57520 6749 57529 6783
rect 57529 6749 57563 6783
rect 57563 6749 57572 6783
rect 57520 6740 57572 6749
rect 57980 6672 58032 6724
rect 51448 6604 51500 6656
rect 52736 6604 52788 6656
rect 52920 6604 52972 6656
rect 55588 6604 55640 6656
rect 56048 6647 56100 6656
rect 56048 6613 56057 6647
rect 56057 6613 56091 6647
rect 56091 6613 56100 6647
rect 56048 6604 56100 6613
rect 15398 6502 15450 6554
rect 15462 6502 15514 6554
rect 15526 6502 15578 6554
rect 15590 6502 15642 6554
rect 15654 6502 15706 6554
rect 29846 6502 29898 6554
rect 29910 6502 29962 6554
rect 29974 6502 30026 6554
rect 30038 6502 30090 6554
rect 30102 6502 30154 6554
rect 44294 6502 44346 6554
rect 44358 6502 44410 6554
rect 44422 6502 44474 6554
rect 44486 6502 44538 6554
rect 44550 6502 44602 6554
rect 2136 6400 2188 6452
rect 5448 6400 5500 6452
rect 7840 6400 7892 6452
rect 9772 6400 9824 6452
rect 10048 6400 10100 6452
rect 11152 6400 11204 6452
rect 2136 6264 2188 6316
rect 2504 6307 2556 6316
rect 2504 6273 2513 6307
rect 2513 6273 2547 6307
rect 2547 6273 2556 6307
rect 2504 6264 2556 6273
rect 5908 6332 5960 6384
rect 6736 6332 6788 6384
rect 3884 6307 3936 6316
rect 3884 6273 3893 6307
rect 3893 6273 3927 6307
rect 3927 6273 3936 6307
rect 3884 6264 3936 6273
rect 3976 6264 4028 6316
rect 4252 6264 4304 6316
rect 4344 6196 4396 6248
rect 5172 6264 5224 6316
rect 5540 6264 5592 6316
rect 9128 6307 9180 6316
rect 9128 6273 9137 6307
rect 9137 6273 9171 6307
rect 9171 6273 9180 6307
rect 9128 6264 9180 6273
rect 4252 6128 4304 6180
rect 4804 6128 4856 6180
rect 5356 6196 5408 6248
rect 5724 6196 5776 6248
rect 9864 6264 9916 6316
rect 11428 6332 11480 6384
rect 19340 6400 19392 6452
rect 22560 6400 22612 6452
rect 23480 6443 23532 6452
rect 23480 6409 23489 6443
rect 23489 6409 23523 6443
rect 23523 6409 23532 6443
rect 23480 6400 23532 6409
rect 10600 6273 10609 6282
rect 10609 6273 10643 6282
rect 10643 6273 10652 6282
rect 10600 6230 10652 6273
rect 10968 6264 11020 6316
rect 11152 6264 11204 6316
rect 12716 6307 12768 6316
rect 12716 6273 12725 6307
rect 12725 6273 12759 6307
rect 12759 6273 12768 6307
rect 12716 6264 12768 6273
rect 5540 6128 5592 6180
rect 1952 6060 2004 6112
rect 2964 6060 3016 6112
rect 4712 6060 4764 6112
rect 5448 6060 5500 6112
rect 6736 6060 6788 6112
rect 12900 6196 12952 6248
rect 8576 6060 8628 6112
rect 9772 6060 9824 6112
rect 10968 6103 11020 6112
rect 10968 6069 10977 6103
rect 10977 6069 11011 6103
rect 11011 6069 11020 6103
rect 10968 6060 11020 6069
rect 11152 6060 11204 6112
rect 11796 6060 11848 6112
rect 14096 6264 14148 6316
rect 18328 6332 18380 6384
rect 18788 6375 18840 6384
rect 18788 6341 18797 6375
rect 18797 6341 18831 6375
rect 18831 6341 18840 6375
rect 18788 6332 18840 6341
rect 19064 6332 19116 6384
rect 14832 6264 14884 6316
rect 15108 6264 15160 6316
rect 16948 6264 17000 6316
rect 18696 6264 18748 6316
rect 19616 6307 19668 6316
rect 19616 6273 19625 6307
rect 19625 6273 19659 6307
rect 19659 6273 19668 6307
rect 19616 6264 19668 6273
rect 20260 6307 20312 6316
rect 20260 6273 20269 6307
rect 20269 6273 20303 6307
rect 20303 6273 20312 6307
rect 20260 6264 20312 6273
rect 21640 6332 21692 6384
rect 16672 6196 16724 6248
rect 17868 6239 17920 6248
rect 17868 6205 17877 6239
rect 17877 6205 17911 6239
rect 17911 6205 17920 6239
rect 17868 6196 17920 6205
rect 14188 6128 14240 6180
rect 16396 6060 16448 6112
rect 16764 6103 16816 6112
rect 16764 6069 16773 6103
rect 16773 6069 16807 6103
rect 16807 6069 16816 6103
rect 16764 6060 16816 6069
rect 17224 6103 17276 6112
rect 17224 6069 17233 6103
rect 17233 6069 17267 6103
rect 17267 6069 17276 6103
rect 17224 6060 17276 6069
rect 17408 6060 17460 6112
rect 18604 6103 18656 6112
rect 18604 6069 18613 6103
rect 18613 6069 18647 6103
rect 18647 6069 18656 6103
rect 18604 6060 18656 6069
rect 22008 6307 22060 6316
rect 22008 6273 22017 6307
rect 22017 6273 22051 6307
rect 22051 6273 22060 6307
rect 22008 6264 22060 6273
rect 22192 6307 22244 6316
rect 22192 6273 22201 6307
rect 22201 6273 22235 6307
rect 22235 6273 22244 6307
rect 23388 6307 23440 6316
rect 22192 6264 22244 6273
rect 23388 6273 23397 6307
rect 23397 6273 23431 6307
rect 23431 6273 23440 6307
rect 23388 6264 23440 6273
rect 23572 6307 23624 6316
rect 23572 6273 23581 6307
rect 23581 6273 23615 6307
rect 23615 6273 23624 6307
rect 23572 6264 23624 6273
rect 24032 6307 24084 6316
rect 24032 6273 24041 6307
rect 24041 6273 24075 6307
rect 24075 6273 24084 6307
rect 24032 6264 24084 6273
rect 24216 6307 24268 6316
rect 24216 6273 24225 6307
rect 24225 6273 24259 6307
rect 24259 6273 24268 6307
rect 24216 6264 24268 6273
rect 24676 6264 24728 6316
rect 24768 6196 24820 6248
rect 20996 6128 21048 6180
rect 24032 6128 24084 6180
rect 22100 6060 22152 6112
rect 22468 6103 22520 6112
rect 22468 6069 22477 6103
rect 22477 6069 22511 6103
rect 22511 6069 22520 6103
rect 22468 6060 22520 6069
rect 24952 6060 25004 6112
rect 25504 6307 25556 6316
rect 25504 6273 25513 6307
rect 25513 6273 25547 6307
rect 25547 6273 25556 6307
rect 25504 6264 25556 6273
rect 25872 6264 25924 6316
rect 26148 6307 26200 6316
rect 26148 6273 26157 6307
rect 26157 6273 26191 6307
rect 26191 6273 26200 6307
rect 26148 6264 26200 6273
rect 26240 6264 26292 6316
rect 28080 6307 28132 6316
rect 28080 6273 28089 6307
rect 28089 6273 28123 6307
rect 28123 6273 28132 6307
rect 28080 6264 28132 6273
rect 28816 6400 28868 6452
rect 30380 6375 30432 6384
rect 28816 6264 28868 6316
rect 29460 6307 29512 6316
rect 29460 6273 29469 6307
rect 29469 6273 29503 6307
rect 29503 6273 29512 6307
rect 29460 6264 29512 6273
rect 30380 6341 30389 6375
rect 30389 6341 30423 6375
rect 30423 6341 30432 6375
rect 30380 6332 30432 6341
rect 30472 6332 30524 6384
rect 31944 6400 31996 6452
rect 29644 6307 29696 6316
rect 29644 6273 29653 6307
rect 29653 6273 29687 6307
rect 29687 6273 29696 6307
rect 29644 6264 29696 6273
rect 27252 6128 27304 6180
rect 27436 6171 27488 6180
rect 27436 6137 27445 6171
rect 27445 6137 27479 6171
rect 27479 6137 27488 6171
rect 27436 6128 27488 6137
rect 31668 6332 31720 6384
rect 34428 6400 34480 6452
rect 34888 6400 34940 6452
rect 37004 6400 37056 6452
rect 32312 6332 32364 6384
rect 32956 6332 33008 6384
rect 33140 6332 33192 6384
rect 33876 6332 33928 6384
rect 32404 6307 32456 6316
rect 32404 6273 32413 6307
rect 32413 6273 32447 6307
rect 32447 6273 32456 6307
rect 32404 6264 32456 6273
rect 34428 6307 34480 6316
rect 34428 6273 34437 6307
rect 34437 6273 34471 6307
rect 34471 6273 34480 6307
rect 34428 6264 34480 6273
rect 34612 6307 34664 6316
rect 34612 6273 34621 6307
rect 34621 6273 34655 6307
rect 34655 6273 34664 6307
rect 34612 6264 34664 6273
rect 32588 6196 32640 6248
rect 34888 6196 34940 6248
rect 35808 6264 35860 6316
rect 35900 6264 35952 6316
rect 38476 6332 38528 6384
rect 40684 6400 40736 6452
rect 40868 6400 40920 6452
rect 46204 6400 46256 6452
rect 49976 6400 50028 6452
rect 50528 6443 50580 6452
rect 50528 6409 50537 6443
rect 50537 6409 50571 6443
rect 50571 6409 50580 6443
rect 50528 6400 50580 6409
rect 41788 6332 41840 6384
rect 37740 6307 37792 6316
rect 37740 6273 37749 6307
rect 37749 6273 37783 6307
rect 37783 6273 37792 6307
rect 37740 6264 37792 6273
rect 38292 6239 38344 6248
rect 38292 6205 38301 6239
rect 38301 6205 38335 6239
rect 38335 6205 38344 6239
rect 38292 6196 38344 6205
rect 38660 6264 38712 6316
rect 40224 6264 40276 6316
rect 41604 6264 41656 6316
rect 41696 6307 41748 6316
rect 41696 6273 41705 6307
rect 41705 6273 41739 6307
rect 41739 6273 41748 6307
rect 41696 6264 41748 6273
rect 39304 6196 39356 6248
rect 40040 6239 40092 6248
rect 40040 6205 40049 6239
rect 40049 6205 40083 6239
rect 40083 6205 40092 6239
rect 40040 6196 40092 6205
rect 41420 6196 41472 6248
rect 42616 6196 42668 6248
rect 35900 6128 35952 6180
rect 36084 6128 36136 6180
rect 36912 6128 36964 6180
rect 37004 6128 37056 6180
rect 38016 6128 38068 6180
rect 40132 6128 40184 6180
rect 44088 6332 44140 6384
rect 45100 6307 45152 6316
rect 45100 6273 45118 6307
rect 45118 6273 45152 6307
rect 45100 6264 45152 6273
rect 45376 6307 45428 6316
rect 45376 6273 45385 6307
rect 45385 6273 45419 6307
rect 45419 6273 45428 6307
rect 46848 6307 46900 6316
rect 45376 6264 45428 6273
rect 46848 6273 46857 6307
rect 46857 6273 46891 6307
rect 46891 6273 46900 6307
rect 46848 6264 46900 6273
rect 50068 6307 50120 6316
rect 50068 6273 50077 6307
rect 50077 6273 50111 6307
rect 50111 6273 50120 6307
rect 50068 6264 50120 6273
rect 50712 6307 50764 6316
rect 50712 6273 50721 6307
rect 50721 6273 50755 6307
rect 50755 6273 50764 6307
rect 50712 6264 50764 6273
rect 45836 6171 45888 6180
rect 45836 6137 45845 6171
rect 45845 6137 45879 6171
rect 45879 6137 45888 6171
rect 45836 6128 45888 6137
rect 49424 6239 49476 6248
rect 49424 6205 49433 6239
rect 49433 6205 49467 6239
rect 49467 6205 49476 6239
rect 51448 6332 51500 6384
rect 49424 6196 49476 6205
rect 28724 6060 28776 6112
rect 29920 6103 29972 6112
rect 29920 6069 29929 6103
rect 29929 6069 29963 6103
rect 29963 6069 29972 6103
rect 29920 6060 29972 6069
rect 30564 6103 30616 6112
rect 30564 6069 30573 6103
rect 30573 6069 30607 6103
rect 30607 6069 30616 6103
rect 30564 6060 30616 6069
rect 31208 6103 31260 6112
rect 31208 6069 31217 6103
rect 31217 6069 31251 6103
rect 31251 6069 31260 6103
rect 31208 6060 31260 6069
rect 33048 6060 33100 6112
rect 35164 6060 35216 6112
rect 40776 6060 40828 6112
rect 41328 6103 41380 6112
rect 41328 6069 41337 6103
rect 41337 6069 41371 6103
rect 41371 6069 41380 6103
rect 41328 6060 41380 6069
rect 42616 6060 42668 6112
rect 48044 6060 48096 6112
rect 49332 6060 49384 6112
rect 49976 6060 50028 6112
rect 52644 6264 52696 6316
rect 55404 6307 55456 6316
rect 52184 6239 52236 6248
rect 52184 6205 52193 6239
rect 52193 6205 52227 6239
rect 52227 6205 52236 6239
rect 52184 6196 52236 6205
rect 53104 6103 53156 6112
rect 53104 6069 53113 6103
rect 53113 6069 53147 6103
rect 53147 6069 53156 6103
rect 53104 6060 53156 6069
rect 54116 6239 54168 6248
rect 54116 6205 54125 6239
rect 54125 6205 54159 6239
rect 54159 6205 54168 6239
rect 55128 6239 55180 6248
rect 54116 6196 54168 6205
rect 55128 6205 55137 6239
rect 55137 6205 55171 6239
rect 55171 6205 55180 6239
rect 55128 6196 55180 6205
rect 55404 6273 55413 6307
rect 55413 6273 55447 6307
rect 55447 6273 55456 6307
rect 55404 6264 55456 6273
rect 56048 6332 56100 6384
rect 55588 6264 55640 6316
rect 56324 6264 56376 6316
rect 55956 6196 56008 6248
rect 55404 6060 55456 6112
rect 56140 6060 56192 6112
rect 56324 6103 56376 6112
rect 56324 6069 56333 6103
rect 56333 6069 56367 6103
rect 56367 6069 56376 6103
rect 56324 6060 56376 6069
rect 8174 5958 8226 6010
rect 8238 5958 8290 6010
rect 8302 5958 8354 6010
rect 8366 5958 8418 6010
rect 8430 5958 8482 6010
rect 22622 5958 22674 6010
rect 22686 5958 22738 6010
rect 22750 5958 22802 6010
rect 22814 5958 22866 6010
rect 22878 5958 22930 6010
rect 37070 5958 37122 6010
rect 37134 5958 37186 6010
rect 37198 5958 37250 6010
rect 37262 5958 37314 6010
rect 37326 5958 37378 6010
rect 51518 5958 51570 6010
rect 51582 5958 51634 6010
rect 51646 5958 51698 6010
rect 51710 5958 51762 6010
rect 51774 5958 51826 6010
rect 1860 5856 1912 5908
rect 3884 5856 3936 5908
rect 4712 5856 4764 5908
rect 7840 5856 7892 5908
rect 9772 5856 9824 5908
rect 9864 5856 9916 5908
rect 4252 5788 4304 5840
rect 6644 5831 6696 5840
rect 6644 5797 6653 5831
rect 6653 5797 6687 5831
rect 6687 5797 6696 5831
rect 6644 5788 6696 5797
rect 8576 5788 8628 5840
rect 9128 5788 9180 5840
rect 13728 5856 13780 5908
rect 3056 5720 3108 5772
rect 6368 5720 6420 5772
rect 2228 5695 2280 5704
rect 2228 5661 2237 5695
rect 2237 5661 2271 5695
rect 2271 5661 2280 5695
rect 2228 5652 2280 5661
rect 2780 5652 2832 5704
rect 3424 5652 3476 5704
rect 3700 5652 3752 5704
rect 3976 5695 4028 5704
rect 3976 5661 3980 5695
rect 3980 5661 4014 5695
rect 4014 5661 4028 5695
rect 3976 5652 4028 5661
rect 4160 5695 4212 5704
rect 4160 5661 4169 5695
rect 4169 5661 4203 5695
rect 4203 5661 4212 5695
rect 4160 5652 4212 5661
rect 5356 5652 5408 5704
rect 5540 5695 5592 5704
rect 5540 5661 5574 5695
rect 5574 5661 5592 5695
rect 5540 5652 5592 5661
rect 3056 5627 3108 5636
rect 3056 5593 3065 5627
rect 3065 5593 3099 5627
rect 3099 5593 3108 5627
rect 3056 5584 3108 5593
rect 5172 5584 5224 5636
rect 5908 5584 5960 5636
rect 10232 5720 10284 5772
rect 16764 5856 16816 5908
rect 17500 5899 17552 5908
rect 17500 5865 17509 5899
rect 17509 5865 17543 5899
rect 17543 5865 17552 5899
rect 17500 5856 17552 5865
rect 18236 5856 18288 5908
rect 18788 5856 18840 5908
rect 22008 5856 22060 5908
rect 24216 5856 24268 5908
rect 28080 5856 28132 5908
rect 29460 5856 29512 5908
rect 32312 5856 32364 5908
rect 33784 5899 33836 5908
rect 33784 5865 33793 5899
rect 33793 5865 33827 5899
rect 33827 5865 33836 5899
rect 33784 5856 33836 5865
rect 34612 5856 34664 5908
rect 36820 5856 36872 5908
rect 36912 5856 36964 5908
rect 41328 5899 41380 5908
rect 15108 5788 15160 5840
rect 20996 5788 21048 5840
rect 29736 5788 29788 5840
rect 30472 5788 30524 5840
rect 33232 5788 33284 5840
rect 36084 5788 36136 5840
rect 37648 5788 37700 5840
rect 38016 5788 38068 5840
rect 40132 5788 40184 5840
rect 7656 5695 7708 5704
rect 7656 5661 7665 5695
rect 7665 5661 7699 5695
rect 7699 5661 7708 5695
rect 7656 5652 7708 5661
rect 8668 5652 8720 5704
rect 9128 5652 9180 5704
rect 17868 5720 17920 5772
rect 9496 5584 9548 5636
rect 4068 5516 4120 5568
rect 4528 5516 4580 5568
rect 7840 5516 7892 5568
rect 10232 5516 10284 5568
rect 11704 5652 11756 5704
rect 10968 5627 11020 5636
rect 10968 5593 11002 5627
rect 11002 5593 11020 5627
rect 10968 5584 11020 5593
rect 13452 5695 13504 5704
rect 13452 5661 13461 5695
rect 13461 5661 13495 5695
rect 13495 5661 13504 5695
rect 13452 5652 13504 5661
rect 14004 5652 14056 5704
rect 14188 5652 14240 5704
rect 16396 5695 16448 5704
rect 16396 5661 16405 5695
rect 16405 5661 16439 5695
rect 16439 5661 16448 5695
rect 16396 5652 16448 5661
rect 16488 5652 16540 5704
rect 16672 5695 16724 5704
rect 16672 5661 16681 5695
rect 16681 5661 16715 5695
rect 16715 5661 16724 5695
rect 16672 5652 16724 5661
rect 17040 5652 17092 5704
rect 18236 5695 18288 5704
rect 13176 5584 13228 5636
rect 18236 5661 18245 5695
rect 18245 5661 18279 5695
rect 18279 5661 18288 5695
rect 18236 5652 18288 5661
rect 21640 5720 21692 5772
rect 23112 5763 23164 5772
rect 23112 5729 23121 5763
rect 23121 5729 23155 5763
rect 23155 5729 23164 5763
rect 23112 5720 23164 5729
rect 23296 5720 23348 5772
rect 33048 5720 33100 5772
rect 36452 5720 36504 5772
rect 18420 5695 18472 5704
rect 18420 5661 18429 5695
rect 18429 5661 18463 5695
rect 18463 5661 18472 5695
rect 18420 5652 18472 5661
rect 18696 5652 18748 5704
rect 19616 5652 19668 5704
rect 21088 5652 21140 5704
rect 21272 5695 21324 5704
rect 21272 5661 21281 5695
rect 21281 5661 21315 5695
rect 21315 5661 21324 5695
rect 21272 5652 21324 5661
rect 22468 5652 22520 5704
rect 23848 5695 23900 5704
rect 23848 5661 23857 5695
rect 23857 5661 23891 5695
rect 23891 5661 23900 5695
rect 23848 5652 23900 5661
rect 24952 5695 25004 5704
rect 24952 5661 24986 5695
rect 24986 5661 25004 5695
rect 24952 5652 25004 5661
rect 18880 5584 18932 5636
rect 19432 5627 19484 5636
rect 19432 5593 19441 5627
rect 19441 5593 19475 5627
rect 19475 5593 19484 5627
rect 19432 5584 19484 5593
rect 12716 5559 12768 5568
rect 12716 5525 12725 5559
rect 12725 5525 12759 5559
rect 12759 5525 12768 5559
rect 12716 5516 12768 5525
rect 13820 5516 13872 5568
rect 14832 5516 14884 5568
rect 17040 5559 17092 5568
rect 17040 5525 17049 5559
rect 17049 5525 17083 5559
rect 17083 5525 17092 5559
rect 17040 5516 17092 5525
rect 19524 5516 19576 5568
rect 24032 5584 24084 5636
rect 26976 5627 27028 5636
rect 26976 5593 26985 5627
rect 26985 5593 27019 5627
rect 27019 5593 27028 5627
rect 28724 5695 28776 5704
rect 28724 5661 28742 5695
rect 28742 5661 28776 5695
rect 29000 5695 29052 5704
rect 28724 5652 28776 5661
rect 29000 5661 29009 5695
rect 29009 5661 29043 5695
rect 29043 5661 29052 5695
rect 29000 5652 29052 5661
rect 29736 5695 29788 5704
rect 29736 5661 29745 5695
rect 29745 5661 29779 5695
rect 29779 5661 29788 5695
rect 29736 5652 29788 5661
rect 30380 5695 30432 5704
rect 30380 5661 30389 5695
rect 30389 5661 30423 5695
rect 30423 5661 30432 5695
rect 30380 5652 30432 5661
rect 32680 5695 32732 5704
rect 32680 5661 32689 5695
rect 32689 5661 32723 5695
rect 32723 5661 32732 5695
rect 32680 5652 32732 5661
rect 34888 5695 34940 5704
rect 34888 5661 34897 5695
rect 34897 5661 34931 5695
rect 34931 5661 34940 5695
rect 34888 5652 34940 5661
rect 26976 5584 27028 5593
rect 22192 5516 22244 5568
rect 26240 5516 26292 5568
rect 29920 5584 29972 5636
rect 32588 5584 32640 5636
rect 33324 5584 33376 5636
rect 35348 5652 35400 5704
rect 36084 5695 36136 5704
rect 36084 5661 36093 5695
rect 36093 5661 36127 5695
rect 36127 5661 36136 5695
rect 36084 5652 36136 5661
rect 38568 5695 38620 5704
rect 38568 5661 38577 5695
rect 38577 5661 38611 5695
rect 38611 5661 38620 5695
rect 38568 5652 38620 5661
rect 30748 5516 30800 5568
rect 34796 5516 34848 5568
rect 35900 5584 35952 5636
rect 40040 5720 40092 5772
rect 41328 5865 41358 5899
rect 41358 5865 41380 5899
rect 41328 5856 41380 5865
rect 42432 5856 42484 5908
rect 43996 5899 44048 5908
rect 43996 5865 44005 5899
rect 44005 5865 44039 5899
rect 44039 5865 44048 5899
rect 43996 5856 44048 5865
rect 45652 5856 45704 5908
rect 45560 5788 45612 5840
rect 49240 5788 49292 5840
rect 45376 5720 45428 5772
rect 47584 5720 47636 5772
rect 50804 5831 50856 5840
rect 50804 5797 50813 5831
rect 50813 5797 50847 5831
rect 50847 5797 50856 5831
rect 50804 5788 50856 5797
rect 53196 5788 53248 5840
rect 52552 5763 52604 5772
rect 52552 5729 52561 5763
rect 52561 5729 52595 5763
rect 52595 5729 52604 5763
rect 52552 5720 52604 5729
rect 57796 5720 57848 5772
rect 40408 5695 40460 5704
rect 40408 5661 40417 5695
rect 40417 5661 40451 5695
rect 40451 5661 40460 5695
rect 40408 5652 40460 5661
rect 42432 5652 42484 5704
rect 44180 5695 44232 5704
rect 44180 5661 44189 5695
rect 44189 5661 44223 5695
rect 44223 5661 44232 5695
rect 44180 5652 44232 5661
rect 45008 5695 45060 5704
rect 45008 5661 45017 5695
rect 45017 5661 45051 5695
rect 45051 5661 45060 5695
rect 45008 5652 45060 5661
rect 45284 5652 45336 5704
rect 47216 5695 47268 5704
rect 47216 5661 47225 5695
rect 47225 5661 47259 5695
rect 47259 5661 47268 5695
rect 47216 5652 47268 5661
rect 49240 5652 49292 5704
rect 41420 5584 41472 5636
rect 46848 5584 46900 5636
rect 52184 5652 52236 5704
rect 55220 5652 55272 5704
rect 55588 5695 55640 5704
rect 55588 5661 55597 5695
rect 55597 5661 55631 5695
rect 55631 5661 55640 5695
rect 55588 5652 55640 5661
rect 57336 5695 57388 5704
rect 57336 5661 57345 5695
rect 57345 5661 57379 5695
rect 57379 5661 57388 5695
rect 57336 5652 57388 5661
rect 37740 5516 37792 5568
rect 39120 5559 39172 5568
rect 39120 5525 39129 5559
rect 39129 5525 39163 5559
rect 39163 5525 39172 5559
rect 39120 5516 39172 5525
rect 43352 5516 43404 5568
rect 46572 5516 46624 5568
rect 48320 5516 48372 5568
rect 55956 5584 56008 5636
rect 53840 5516 53892 5568
rect 54208 5559 54260 5568
rect 54208 5525 54217 5559
rect 54217 5525 54251 5559
rect 54251 5525 54260 5559
rect 54208 5516 54260 5525
rect 55680 5516 55732 5568
rect 57980 5516 58032 5568
rect 15398 5414 15450 5466
rect 15462 5414 15514 5466
rect 15526 5414 15578 5466
rect 15590 5414 15642 5466
rect 15654 5414 15706 5466
rect 29846 5414 29898 5466
rect 29910 5414 29962 5466
rect 29974 5414 30026 5466
rect 30038 5414 30090 5466
rect 30102 5414 30154 5466
rect 44294 5414 44346 5466
rect 44358 5414 44410 5466
rect 44422 5414 44474 5466
rect 44486 5414 44538 5466
rect 44550 5414 44602 5466
rect 3976 5312 4028 5364
rect 1952 5287 2004 5296
rect 1952 5253 1961 5287
rect 1961 5253 1995 5287
rect 1995 5253 2004 5287
rect 2780 5287 2832 5296
rect 1952 5244 2004 5253
rect 2780 5253 2789 5287
rect 2789 5253 2823 5287
rect 2823 5253 2832 5287
rect 2780 5244 2832 5253
rect 3148 5287 3200 5296
rect 3148 5253 3157 5287
rect 3157 5253 3191 5287
rect 3191 5253 3200 5287
rect 3148 5244 3200 5253
rect 10048 5312 10100 5364
rect 2136 5219 2188 5228
rect 2136 5185 2145 5219
rect 2145 5185 2179 5219
rect 2179 5185 2188 5219
rect 2136 5176 2188 5185
rect 4252 5176 4304 5228
rect 5448 5244 5500 5296
rect 7380 5244 7432 5296
rect 4528 5176 4580 5228
rect 7288 5176 7340 5228
rect 5448 5108 5500 5160
rect 6828 5108 6880 5160
rect 8208 5176 8260 5228
rect 5816 5083 5868 5092
rect 5816 5049 5825 5083
rect 5825 5049 5859 5083
rect 5859 5049 5868 5083
rect 5816 5040 5868 5049
rect 4804 4972 4856 5024
rect 6000 4972 6052 5024
rect 7380 4972 7432 5024
rect 7932 4972 7984 5024
rect 10508 5244 10560 5296
rect 10600 5219 10652 5228
rect 9496 5040 9548 5092
rect 9864 5040 9916 5092
rect 10600 5185 10609 5219
rect 10609 5185 10643 5219
rect 10643 5185 10652 5219
rect 10600 5176 10652 5185
rect 10968 5040 11020 5092
rect 13728 5312 13780 5364
rect 12900 5244 12952 5296
rect 11888 5176 11940 5228
rect 14004 5176 14056 5228
rect 14924 5244 14976 5296
rect 16488 5312 16540 5364
rect 15108 5176 15160 5228
rect 16948 5312 17000 5364
rect 17408 5312 17460 5364
rect 18236 5312 18288 5364
rect 17040 5244 17092 5296
rect 17960 5244 18012 5296
rect 18880 5287 18932 5296
rect 18880 5253 18889 5287
rect 18889 5253 18923 5287
rect 18923 5253 18932 5287
rect 18880 5244 18932 5253
rect 21180 5312 21232 5364
rect 22376 5312 22428 5364
rect 19524 5244 19576 5296
rect 21456 5244 21508 5296
rect 24584 5244 24636 5296
rect 25964 5312 26016 5364
rect 27988 5312 28040 5364
rect 31300 5312 31352 5364
rect 21732 5176 21784 5228
rect 22284 5176 22336 5228
rect 23296 5219 23348 5228
rect 23296 5185 23305 5219
rect 23305 5185 23339 5219
rect 23339 5185 23348 5219
rect 23296 5176 23348 5185
rect 23388 5176 23440 5228
rect 11520 5151 11572 5160
rect 11520 5117 11529 5151
rect 11529 5117 11563 5151
rect 11563 5117 11572 5151
rect 11520 5108 11572 5117
rect 15844 5108 15896 5160
rect 16488 5108 16540 5160
rect 16948 5040 17000 5092
rect 10416 4972 10468 5024
rect 11980 4972 12032 5024
rect 15200 4972 15252 5024
rect 16764 4972 16816 5024
rect 19524 5108 19576 5160
rect 21640 5108 21692 5160
rect 23112 5108 23164 5160
rect 25504 5108 25556 5160
rect 25964 5219 26016 5228
rect 25964 5185 25973 5219
rect 25973 5185 26007 5219
rect 26007 5185 26016 5219
rect 25964 5176 26016 5185
rect 27528 5244 27580 5296
rect 26424 5176 26476 5228
rect 27712 5219 27764 5228
rect 27712 5185 27721 5219
rect 27721 5185 27755 5219
rect 27755 5185 27764 5219
rect 27712 5176 27764 5185
rect 27804 5176 27856 5228
rect 27988 5219 28040 5228
rect 27988 5185 27997 5219
rect 27997 5185 28031 5219
rect 28031 5185 28040 5219
rect 28448 5219 28500 5228
rect 27988 5176 28040 5185
rect 28448 5185 28457 5219
rect 28457 5185 28491 5219
rect 28491 5185 28500 5219
rect 28448 5176 28500 5185
rect 28724 5219 28776 5228
rect 28724 5185 28733 5219
rect 28733 5185 28767 5219
rect 28767 5185 28776 5219
rect 28724 5176 28776 5185
rect 32680 5244 32732 5296
rect 34796 5312 34848 5364
rect 38660 5312 38712 5364
rect 34520 5244 34572 5296
rect 38568 5244 38620 5296
rect 30288 5176 30340 5228
rect 19340 5015 19392 5024
rect 19340 4981 19349 5015
rect 19349 4981 19383 5015
rect 19383 4981 19392 5015
rect 19340 4972 19392 4981
rect 20904 4972 20956 5024
rect 24952 4972 25004 5024
rect 26792 4972 26844 5024
rect 26884 4972 26936 5024
rect 27712 5040 27764 5092
rect 28724 5040 28776 5092
rect 28908 5083 28960 5092
rect 28908 5049 28917 5083
rect 28917 5049 28951 5083
rect 28951 5049 28960 5083
rect 28908 5040 28960 5049
rect 27804 4972 27856 5024
rect 29460 5015 29512 5024
rect 29460 4981 29469 5015
rect 29469 4981 29503 5015
rect 29503 4981 29512 5015
rect 29460 4972 29512 4981
rect 32772 5176 32824 5228
rect 33784 5108 33836 5160
rect 36084 5176 36136 5228
rect 38752 5219 38804 5228
rect 38752 5185 38761 5219
rect 38761 5185 38795 5219
rect 38795 5185 38804 5219
rect 38752 5176 38804 5185
rect 35256 5151 35308 5160
rect 35256 5117 35265 5151
rect 35265 5117 35299 5151
rect 35299 5117 35308 5151
rect 35256 5108 35308 5117
rect 36912 5108 36964 5160
rect 31760 5040 31812 5092
rect 31668 4972 31720 5024
rect 33692 4972 33744 5024
rect 35624 4972 35676 5024
rect 37740 4972 37792 5024
rect 39028 5219 39080 5228
rect 39028 5185 39037 5219
rect 39037 5185 39071 5219
rect 39071 5185 39080 5219
rect 39028 5176 39080 5185
rect 40040 5244 40092 5296
rect 42432 5312 42484 5364
rect 46848 5355 46900 5364
rect 46848 5321 46857 5355
rect 46857 5321 46891 5355
rect 46891 5321 46900 5355
rect 46848 5312 46900 5321
rect 47584 5355 47636 5364
rect 47584 5321 47593 5355
rect 47593 5321 47627 5355
rect 47627 5321 47636 5355
rect 47584 5312 47636 5321
rect 48688 5312 48740 5364
rect 49424 5312 49476 5364
rect 49516 5312 49568 5364
rect 51448 5312 51500 5364
rect 52644 5312 52696 5364
rect 39672 5176 39724 5228
rect 44088 5244 44140 5296
rect 44456 5244 44508 5296
rect 43812 5219 43864 5228
rect 43812 5185 43846 5219
rect 43846 5185 43864 5219
rect 43812 5176 43864 5185
rect 40592 5040 40644 5092
rect 45192 5176 45244 5228
rect 48320 5244 48372 5296
rect 55680 5312 55732 5364
rect 57336 5312 57388 5364
rect 45928 5176 45980 5228
rect 47216 5176 47268 5228
rect 52092 5219 52144 5228
rect 52092 5185 52101 5219
rect 52101 5185 52135 5219
rect 52135 5185 52144 5219
rect 52092 5176 52144 5185
rect 53288 5176 53340 5228
rect 54208 5219 54260 5228
rect 54208 5185 54217 5219
rect 54217 5185 54251 5219
rect 54251 5185 54260 5219
rect 54208 5176 54260 5185
rect 54760 5176 54812 5228
rect 56324 5244 56376 5296
rect 46020 5108 46072 5160
rect 46204 5108 46256 5160
rect 49516 5108 49568 5160
rect 53196 5108 53248 5160
rect 53472 5108 53524 5160
rect 52092 5040 52144 5092
rect 55220 5108 55272 5160
rect 56140 5176 56192 5228
rect 58072 5219 58124 5228
rect 58072 5185 58081 5219
rect 58081 5185 58115 5219
rect 58115 5185 58124 5219
rect 58072 5176 58124 5185
rect 56048 5151 56100 5160
rect 56048 5117 56057 5151
rect 56057 5117 56091 5151
rect 56091 5117 56100 5151
rect 56048 5108 56100 5117
rect 55128 5040 55180 5092
rect 57704 5040 57756 5092
rect 40316 4972 40368 5024
rect 41052 4972 41104 5024
rect 42984 4972 43036 5024
rect 48136 5015 48188 5024
rect 48136 4981 48145 5015
rect 48145 4981 48179 5015
rect 48179 4981 48188 5015
rect 48136 4972 48188 4981
rect 50252 4972 50304 5024
rect 51080 5015 51132 5024
rect 51080 4981 51089 5015
rect 51089 4981 51123 5015
rect 51123 4981 51132 5015
rect 51080 4972 51132 4981
rect 51908 4972 51960 5024
rect 52000 5015 52052 5024
rect 52000 4981 52009 5015
rect 52009 4981 52043 5015
rect 52043 4981 52052 5015
rect 52000 4972 52052 4981
rect 53012 4972 53064 5024
rect 55864 4972 55916 5024
rect 8174 4870 8226 4922
rect 8238 4870 8290 4922
rect 8302 4870 8354 4922
rect 8366 4870 8418 4922
rect 8430 4870 8482 4922
rect 22622 4870 22674 4922
rect 22686 4870 22738 4922
rect 22750 4870 22802 4922
rect 22814 4870 22866 4922
rect 22878 4870 22930 4922
rect 37070 4870 37122 4922
rect 37134 4870 37186 4922
rect 37198 4870 37250 4922
rect 37262 4870 37314 4922
rect 37326 4870 37378 4922
rect 51518 4870 51570 4922
rect 51582 4870 51634 4922
rect 51646 4870 51698 4922
rect 51710 4870 51762 4922
rect 51774 4870 51826 4922
rect 2504 4607 2556 4616
rect 2504 4573 2513 4607
rect 2513 4573 2547 4607
rect 2547 4573 2556 4607
rect 2504 4564 2556 4573
rect 4068 4632 4120 4684
rect 6184 4700 6236 4752
rect 7932 4768 7984 4820
rect 8392 4768 8444 4820
rect 10416 4768 10468 4820
rect 10784 4768 10836 4820
rect 10600 4700 10652 4752
rect 6828 4675 6880 4684
rect 6828 4641 6837 4675
rect 6837 4641 6871 4675
rect 6871 4641 6880 4675
rect 6828 4632 6880 4641
rect 10048 4632 10100 4684
rect 2964 4564 3016 4616
rect 4252 4607 4304 4616
rect 4252 4573 4261 4607
rect 4261 4573 4295 4607
rect 4295 4573 4304 4607
rect 4252 4564 4304 4573
rect 5448 4564 5500 4616
rect 8392 4564 8444 4616
rect 8576 4564 8628 4616
rect 9680 4564 9732 4616
rect 1860 4539 1912 4548
rect 1860 4505 1869 4539
rect 1869 4505 1903 4539
rect 1903 4505 1912 4539
rect 1860 4496 1912 4505
rect 2136 4496 2188 4548
rect 5172 4539 5224 4548
rect 5172 4505 5206 4539
rect 5206 4505 5224 4539
rect 5172 4496 5224 4505
rect 7564 4496 7616 4548
rect 7932 4496 7984 4548
rect 8116 4496 8168 4548
rect 8668 4496 8720 4548
rect 5540 4428 5592 4480
rect 6368 4428 6420 4480
rect 9496 4496 9548 4548
rect 12992 4768 13044 4820
rect 14096 4768 14148 4820
rect 14832 4811 14884 4820
rect 14832 4777 14841 4811
rect 14841 4777 14875 4811
rect 14875 4777 14884 4811
rect 14832 4768 14884 4777
rect 17500 4768 17552 4820
rect 21456 4768 21508 4820
rect 22652 4768 22704 4820
rect 23112 4768 23164 4820
rect 23388 4768 23440 4820
rect 24492 4768 24544 4820
rect 25688 4768 25740 4820
rect 27804 4768 27856 4820
rect 29368 4768 29420 4820
rect 30288 4768 30340 4820
rect 30840 4768 30892 4820
rect 33416 4768 33468 4820
rect 36084 4768 36136 4820
rect 17868 4743 17920 4752
rect 17868 4709 17877 4743
rect 17877 4709 17911 4743
rect 17911 4709 17920 4743
rect 17868 4700 17920 4709
rect 20720 4700 20772 4752
rect 25412 4700 25464 4752
rect 34152 4743 34204 4752
rect 11704 4675 11756 4684
rect 11704 4641 11713 4675
rect 11713 4641 11747 4675
rect 11747 4641 11756 4675
rect 11704 4632 11756 4641
rect 14188 4675 14240 4684
rect 14188 4641 14197 4675
rect 14197 4641 14231 4675
rect 14231 4641 14240 4675
rect 14188 4632 14240 4641
rect 14832 4632 14884 4684
rect 16764 4675 16816 4684
rect 16764 4641 16773 4675
rect 16773 4641 16807 4675
rect 16807 4641 16816 4675
rect 16764 4632 16816 4641
rect 20628 4632 20680 4684
rect 22284 4632 22336 4684
rect 22652 4632 22704 4684
rect 14004 4564 14056 4616
rect 14924 4564 14976 4616
rect 19524 4607 19576 4616
rect 9864 4428 9916 4480
rect 12992 4428 13044 4480
rect 13728 4428 13780 4480
rect 15844 4428 15896 4480
rect 16672 4496 16724 4548
rect 18328 4496 18380 4548
rect 18420 4471 18472 4480
rect 18420 4437 18429 4471
rect 18429 4437 18463 4471
rect 18463 4437 18472 4471
rect 18420 4428 18472 4437
rect 19524 4573 19533 4607
rect 19533 4573 19567 4607
rect 19567 4573 19576 4607
rect 21364 4607 21416 4616
rect 19524 4564 19576 4573
rect 21364 4573 21373 4607
rect 21373 4573 21407 4607
rect 21407 4573 21416 4607
rect 21364 4564 21416 4573
rect 21456 4607 21508 4616
rect 21456 4573 21465 4607
rect 21465 4573 21499 4607
rect 21499 4573 21508 4607
rect 21640 4607 21692 4616
rect 21456 4564 21508 4573
rect 21640 4573 21649 4607
rect 21649 4573 21683 4607
rect 21683 4573 21692 4607
rect 21640 4564 21692 4573
rect 22560 4607 22612 4616
rect 22560 4573 22569 4607
rect 22569 4573 22603 4607
rect 22603 4573 22612 4607
rect 22560 4564 22612 4573
rect 23296 4632 23348 4684
rect 25228 4632 25280 4684
rect 19432 4496 19484 4548
rect 23112 4564 23164 4616
rect 24952 4564 25004 4616
rect 28448 4632 28500 4684
rect 34152 4709 34161 4743
rect 34161 4709 34195 4743
rect 34195 4709 34204 4743
rect 34152 4700 34204 4709
rect 35716 4700 35768 4752
rect 20168 4428 20220 4480
rect 23204 4496 23256 4548
rect 24032 4496 24084 4548
rect 25964 4564 26016 4616
rect 26608 4607 26660 4616
rect 26608 4573 26617 4607
rect 26617 4573 26651 4607
rect 26651 4573 26660 4607
rect 26608 4564 26660 4573
rect 25504 4539 25556 4548
rect 22284 4428 22336 4480
rect 22560 4428 22612 4480
rect 22652 4428 22704 4480
rect 25504 4505 25513 4539
rect 25513 4505 25547 4539
rect 25547 4505 25556 4539
rect 25504 4496 25556 4505
rect 29644 4564 29696 4616
rect 24676 4428 24728 4480
rect 27896 4471 27948 4480
rect 27896 4437 27905 4471
rect 27905 4437 27939 4471
rect 27939 4437 27948 4471
rect 27896 4428 27948 4437
rect 29920 4607 29972 4616
rect 29920 4573 29929 4607
rect 29929 4573 29963 4607
rect 29963 4573 29972 4607
rect 29920 4564 29972 4573
rect 30196 4564 30248 4616
rect 31024 4564 31076 4616
rect 36084 4632 36136 4684
rect 30288 4496 30340 4548
rect 31576 4607 31628 4616
rect 31576 4573 31585 4607
rect 31585 4573 31619 4607
rect 31619 4573 31628 4607
rect 31576 4564 31628 4573
rect 32680 4564 32732 4616
rect 31760 4496 31812 4548
rect 31668 4428 31720 4480
rect 35440 4564 35492 4616
rect 39672 4768 39724 4820
rect 41052 4768 41104 4820
rect 43812 4768 43864 4820
rect 45192 4811 45244 4820
rect 45192 4777 45201 4811
rect 45201 4777 45235 4811
rect 45235 4777 45244 4811
rect 45192 4768 45244 4777
rect 46940 4768 46992 4820
rect 51448 4768 51500 4820
rect 51908 4768 51960 4820
rect 53288 4811 53340 4820
rect 38752 4700 38804 4752
rect 36912 4632 36964 4684
rect 35532 4428 35584 4480
rect 37280 4496 37332 4548
rect 38660 4564 38712 4616
rect 41328 4700 41380 4752
rect 44456 4700 44508 4752
rect 40224 4675 40276 4684
rect 40224 4641 40233 4675
rect 40233 4641 40267 4675
rect 40267 4641 40276 4675
rect 40224 4632 40276 4641
rect 41236 4632 41288 4684
rect 42892 4632 42944 4684
rect 53288 4777 53297 4811
rect 53297 4777 53331 4811
rect 53331 4777 53340 4811
rect 53288 4768 53340 4777
rect 54760 4811 54812 4820
rect 54760 4777 54769 4811
rect 54769 4777 54803 4811
rect 54803 4777 54812 4811
rect 54760 4768 54812 4777
rect 55496 4811 55548 4820
rect 55496 4777 55505 4811
rect 55505 4777 55539 4811
rect 55539 4777 55548 4811
rect 55496 4768 55548 4777
rect 58072 4768 58124 4820
rect 55772 4700 55824 4752
rect 41052 4607 41104 4616
rect 41052 4573 41061 4607
rect 41061 4573 41095 4607
rect 41095 4573 41104 4607
rect 41052 4564 41104 4573
rect 41328 4607 41380 4616
rect 41328 4573 41337 4607
rect 41337 4573 41371 4607
rect 41371 4573 41380 4607
rect 41328 4564 41380 4573
rect 42800 4607 42852 4616
rect 42800 4573 42809 4607
rect 42809 4573 42843 4607
rect 42843 4573 42852 4607
rect 42984 4607 43036 4616
rect 42800 4564 42852 4573
rect 42984 4573 42993 4607
rect 42993 4573 43027 4607
rect 43027 4573 43036 4607
rect 42984 4564 43036 4573
rect 43168 4607 43220 4616
rect 43168 4573 43177 4607
rect 43177 4573 43211 4607
rect 43211 4573 43220 4607
rect 43168 4564 43220 4573
rect 44456 4607 44508 4616
rect 44456 4573 44465 4607
rect 44465 4573 44499 4607
rect 44499 4573 44508 4607
rect 44456 4564 44508 4573
rect 45376 4632 45428 4684
rect 48688 4675 48740 4684
rect 48688 4641 48697 4675
rect 48697 4641 48731 4675
rect 48731 4641 48740 4675
rect 48688 4632 48740 4641
rect 57796 4632 57848 4684
rect 37924 4428 37976 4480
rect 39948 4471 40000 4480
rect 39948 4437 39957 4471
rect 39957 4437 39991 4471
rect 39991 4437 40000 4471
rect 39948 4428 40000 4437
rect 45468 4539 45520 4548
rect 41236 4471 41288 4480
rect 41236 4437 41245 4471
rect 41245 4437 41279 4471
rect 41279 4437 41288 4471
rect 41236 4428 41288 4437
rect 43168 4428 43220 4480
rect 44088 4428 44140 4480
rect 45468 4505 45477 4539
rect 45477 4505 45511 4539
rect 45511 4505 45520 4539
rect 45468 4496 45520 4505
rect 45928 4607 45980 4616
rect 45928 4573 45937 4607
rect 45937 4573 45971 4607
rect 45971 4573 45980 4607
rect 45928 4564 45980 4573
rect 48412 4607 48464 4616
rect 48412 4573 48430 4607
rect 48430 4573 48464 4607
rect 48412 4564 48464 4573
rect 52460 4607 52512 4616
rect 48320 4496 48372 4548
rect 48504 4496 48556 4548
rect 48596 4496 48648 4548
rect 52460 4573 52469 4607
rect 52469 4573 52503 4607
rect 52503 4573 52512 4607
rect 52460 4564 52512 4573
rect 52552 4564 52604 4616
rect 53288 4564 53340 4616
rect 53564 4564 53616 4616
rect 55588 4564 55640 4616
rect 55956 4564 56008 4616
rect 57704 4607 57756 4616
rect 55128 4496 55180 4548
rect 46020 4471 46072 4480
rect 46020 4437 46029 4471
rect 46029 4437 46063 4471
rect 46063 4437 46072 4471
rect 46020 4428 46072 4437
rect 48136 4428 48188 4480
rect 55220 4428 55272 4480
rect 55404 4428 55456 4480
rect 57704 4573 57713 4607
rect 57713 4573 57747 4607
rect 57747 4573 57756 4607
rect 57704 4564 57756 4573
rect 57888 4471 57940 4480
rect 57888 4437 57897 4471
rect 57897 4437 57931 4471
rect 57931 4437 57940 4471
rect 57888 4428 57940 4437
rect 15398 4326 15450 4378
rect 15462 4326 15514 4378
rect 15526 4326 15578 4378
rect 15590 4326 15642 4378
rect 15654 4326 15706 4378
rect 29846 4326 29898 4378
rect 29910 4326 29962 4378
rect 29974 4326 30026 4378
rect 30038 4326 30090 4378
rect 30102 4326 30154 4378
rect 44294 4326 44346 4378
rect 44358 4326 44410 4378
rect 44422 4326 44474 4378
rect 44486 4326 44538 4378
rect 44550 4326 44602 4378
rect 2136 4224 2188 4276
rect 4436 4224 4488 4276
rect 6368 4224 6420 4276
rect 7472 4267 7524 4276
rect 7472 4233 7481 4267
rect 7481 4233 7515 4267
rect 7515 4233 7524 4267
rect 7472 4224 7524 4233
rect 7748 4224 7800 4276
rect 6276 4156 6328 4208
rect 7104 4156 7156 4208
rect 7564 4156 7616 4208
rect 1768 4088 1820 4140
rect 2688 4088 2740 4140
rect 2044 4020 2096 4072
rect 2964 4131 3016 4140
rect 2964 4097 2973 4131
rect 2973 4097 3007 4131
rect 3007 4097 3016 4131
rect 2964 4088 3016 4097
rect 3240 4088 3292 4140
rect 4344 4131 4396 4140
rect 4344 4097 4353 4131
rect 4353 4097 4387 4131
rect 4387 4097 4396 4131
rect 4344 4088 4396 4097
rect 4896 4088 4948 4140
rect 5172 4088 5224 4140
rect 6644 4088 6696 4140
rect 7288 4131 7340 4140
rect 7288 4097 7297 4131
rect 7297 4097 7331 4131
rect 7331 4097 7340 4131
rect 7288 4088 7340 4097
rect 8760 4088 8812 4140
rect 10508 4131 10560 4140
rect 10508 4097 10517 4131
rect 10517 4097 10551 4131
rect 10551 4097 10560 4131
rect 10508 4088 10560 4097
rect 17224 4224 17276 4276
rect 19432 4267 19484 4276
rect 19432 4233 19441 4267
rect 19441 4233 19475 4267
rect 19475 4233 19484 4267
rect 19432 4224 19484 4233
rect 21364 4224 21416 4276
rect 24216 4224 24268 4276
rect 24584 4224 24636 4276
rect 10968 4156 11020 4208
rect 13176 4156 13228 4208
rect 14832 4199 14884 4208
rect 14832 4165 14841 4199
rect 14841 4165 14875 4199
rect 14875 4165 14884 4199
rect 14832 4156 14884 4165
rect 14924 4156 14976 4208
rect 15108 4156 15160 4208
rect 16764 4156 16816 4208
rect 18144 4199 18196 4208
rect 13820 4088 13872 4140
rect 14093 4131 14145 4140
rect 14093 4097 14120 4131
rect 14120 4097 14145 4131
rect 14093 4088 14145 4097
rect 14188 4131 14240 4140
rect 14188 4097 14202 4131
rect 14202 4097 14236 4131
rect 14236 4097 14240 4131
rect 14188 4088 14240 4097
rect 14372 4131 14424 4140
rect 14372 4097 14381 4131
rect 14381 4097 14415 4131
rect 14415 4097 14424 4131
rect 15844 4131 15896 4140
rect 14372 4088 14424 4097
rect 15844 4097 15853 4131
rect 15853 4097 15887 4131
rect 15887 4097 15896 4131
rect 15844 4088 15896 4097
rect 5264 4020 5316 4072
rect 5816 3995 5868 4004
rect 2136 3884 2188 3936
rect 5816 3961 5825 3995
rect 5825 3961 5859 3995
rect 5859 3961 5868 3995
rect 5816 3952 5868 3961
rect 7472 3952 7524 4004
rect 8116 3952 8168 4004
rect 4804 3884 4856 3936
rect 4896 3927 4948 3936
rect 4896 3893 4905 3927
rect 4905 3893 4939 3927
rect 4939 3893 4948 3927
rect 4896 3884 4948 3893
rect 7748 3884 7800 3936
rect 11520 4063 11572 4072
rect 11520 4029 11529 4063
rect 11529 4029 11563 4063
rect 11563 4029 11572 4063
rect 11520 4020 11572 4029
rect 16304 4088 16356 4140
rect 18144 4165 18153 4199
rect 18153 4165 18187 4199
rect 18187 4165 18196 4199
rect 18144 4156 18196 4165
rect 17037 4131 17089 4140
rect 17037 4097 17064 4131
rect 17064 4097 17089 4131
rect 17037 4088 17089 4097
rect 16396 4020 16448 4072
rect 16672 4063 16724 4072
rect 16672 4029 16681 4063
rect 16681 4029 16715 4063
rect 16715 4029 16724 4063
rect 16672 4020 16724 4029
rect 13820 3884 13872 3936
rect 14924 3884 14976 3936
rect 17960 4088 18012 4140
rect 23296 4156 23348 4208
rect 17592 4020 17644 4072
rect 19156 4131 19208 4140
rect 19156 4097 19165 4131
rect 19165 4097 19199 4131
rect 19199 4097 19208 4131
rect 19156 4088 19208 4097
rect 20720 4088 20772 4140
rect 21732 4088 21784 4140
rect 16580 3884 16632 3936
rect 22284 4131 22336 4140
rect 22284 4097 22293 4131
rect 22293 4097 22327 4131
rect 22327 4097 22336 4131
rect 22284 4088 22336 4097
rect 23664 4088 23716 4140
rect 23940 4088 23992 4140
rect 24492 4088 24544 4140
rect 24768 4088 24820 4140
rect 25412 4156 25464 4208
rect 25044 4131 25096 4140
rect 25044 4097 25053 4131
rect 25053 4097 25087 4131
rect 25087 4097 25096 4131
rect 25780 4131 25832 4140
rect 25044 4088 25096 4097
rect 25780 4097 25789 4131
rect 25789 4097 25823 4131
rect 25823 4097 25832 4131
rect 25780 4088 25832 4097
rect 26056 4131 26108 4140
rect 26056 4097 26065 4131
rect 26065 4097 26099 4131
rect 26099 4097 26108 4131
rect 26056 4088 26108 4097
rect 27528 4156 27580 4208
rect 22376 4020 22428 4072
rect 23112 4020 23164 4072
rect 28724 4224 28776 4276
rect 31024 4224 31076 4276
rect 31944 4224 31996 4276
rect 27988 4156 28040 4208
rect 29368 4156 29420 4208
rect 31300 4156 31352 4208
rect 30104 4131 30156 4140
rect 30104 4097 30113 4131
rect 30113 4097 30147 4131
rect 30147 4097 30156 4131
rect 30104 4088 30156 4097
rect 30288 4131 30340 4140
rect 30288 4097 30297 4131
rect 30297 4097 30331 4131
rect 30331 4097 30340 4131
rect 30288 4088 30340 4097
rect 32772 4224 32824 4276
rect 37280 4267 37332 4276
rect 37280 4233 37289 4267
rect 37289 4233 37323 4267
rect 37323 4233 37332 4267
rect 37280 4224 37332 4233
rect 40316 4224 40368 4276
rect 41236 4224 41288 4276
rect 43996 4224 44048 4276
rect 46020 4224 46072 4276
rect 48320 4267 48372 4276
rect 48320 4233 48329 4267
rect 48329 4233 48363 4267
rect 48363 4233 48372 4267
rect 48320 4224 48372 4233
rect 52000 4224 52052 4276
rect 53564 4224 53616 4276
rect 57980 4224 58032 4276
rect 32680 4156 32732 4208
rect 32864 4156 32916 4208
rect 32220 4088 32272 4140
rect 32772 4088 32824 4140
rect 34612 4088 34664 4140
rect 35072 4088 35124 4140
rect 35808 4156 35860 4208
rect 40040 4156 40092 4208
rect 40960 4156 41012 4208
rect 31300 4063 31352 4072
rect 31300 4029 31309 4063
rect 31309 4029 31343 4063
rect 31343 4029 31352 4063
rect 31300 4020 31352 4029
rect 31576 4063 31628 4072
rect 31576 4029 31585 4063
rect 31585 4029 31619 4063
rect 31619 4029 31628 4063
rect 31576 4020 31628 4029
rect 29276 3952 29328 4004
rect 18880 3884 18932 3936
rect 19892 3927 19944 3936
rect 19892 3893 19901 3927
rect 19901 3893 19935 3927
rect 19935 3893 19944 3927
rect 19892 3884 19944 3893
rect 21640 3884 21692 3936
rect 23572 3884 23624 3936
rect 23664 3884 23716 3936
rect 25320 3884 25372 3936
rect 25688 3884 25740 3936
rect 26792 3884 26844 3936
rect 28448 3884 28500 3936
rect 33600 4020 33652 4072
rect 34428 4020 34480 4072
rect 35716 4088 35768 4140
rect 37464 4088 37516 4140
rect 36820 4020 36872 4072
rect 34060 3952 34112 4004
rect 33508 3927 33560 3936
rect 33508 3893 33517 3927
rect 33517 3893 33551 3927
rect 33551 3893 33560 3927
rect 33508 3884 33560 3893
rect 35900 3927 35952 3936
rect 35900 3893 35909 3927
rect 35909 3893 35943 3927
rect 35943 3893 35952 3927
rect 35900 3884 35952 3893
rect 35992 3884 36044 3936
rect 36176 3884 36228 3936
rect 37740 4131 37792 4140
rect 37740 4097 37749 4131
rect 37749 4097 37783 4131
rect 37783 4097 37792 4131
rect 37740 4088 37792 4097
rect 37924 4131 37976 4140
rect 37924 4097 37927 4131
rect 37927 4097 37961 4131
rect 37961 4097 37976 4131
rect 39028 4131 39080 4140
rect 37924 4088 37976 4097
rect 39028 4097 39037 4131
rect 39037 4097 39071 4131
rect 39071 4097 39080 4131
rect 39028 4088 39080 4097
rect 39304 4131 39356 4140
rect 39304 4097 39313 4131
rect 39313 4097 39347 4131
rect 39347 4097 39356 4131
rect 39304 4088 39356 4097
rect 39856 4088 39908 4140
rect 40316 4131 40368 4140
rect 40316 4097 40325 4131
rect 40325 4097 40359 4131
rect 40359 4097 40368 4131
rect 40316 4088 40368 4097
rect 40500 4088 40552 4140
rect 40684 4088 40736 4140
rect 40868 4088 40920 4140
rect 41328 4131 41380 4140
rect 41328 4097 41337 4131
rect 41337 4097 41371 4131
rect 41371 4097 41380 4131
rect 41328 4088 41380 4097
rect 42800 4088 42852 4140
rect 43168 4131 43220 4140
rect 43168 4097 43177 4131
rect 43177 4097 43211 4131
rect 43211 4097 43220 4131
rect 43168 4088 43220 4097
rect 41052 3952 41104 4004
rect 42892 4020 42944 4072
rect 43536 4088 43588 4140
rect 43996 4088 44048 4140
rect 45376 4156 45428 4208
rect 43628 4063 43680 4072
rect 43628 4029 43637 4063
rect 43637 4029 43671 4063
rect 43671 4029 43680 4063
rect 43628 4020 43680 4029
rect 44456 4131 44508 4140
rect 44456 4097 44465 4131
rect 44465 4097 44499 4131
rect 44499 4097 44508 4131
rect 44456 4088 44508 4097
rect 49608 4088 49660 4140
rect 51264 4088 51316 4140
rect 51816 4131 51868 4140
rect 51816 4097 51825 4131
rect 51825 4097 51859 4131
rect 51859 4097 51868 4131
rect 51816 4088 51868 4097
rect 52184 4131 52236 4140
rect 41512 3927 41564 3936
rect 41512 3893 41521 3927
rect 41521 3893 41555 3927
rect 41555 3893 41564 3927
rect 41512 3884 41564 3893
rect 42432 3927 42484 3936
rect 42432 3893 42441 3927
rect 42441 3893 42475 3927
rect 42475 3893 42484 3927
rect 42432 3884 42484 3893
rect 43168 3884 43220 3936
rect 52184 4097 52193 4131
rect 52193 4097 52227 4131
rect 52227 4097 52236 4131
rect 52184 4088 52236 4097
rect 54024 4131 54076 4140
rect 54024 4097 54033 4131
rect 54033 4097 54067 4131
rect 54067 4097 54076 4131
rect 54024 4088 54076 4097
rect 55496 4156 55548 4208
rect 55680 4088 55732 4140
rect 55956 4131 56008 4140
rect 55956 4097 55965 4131
rect 55965 4097 55999 4131
rect 55999 4097 56008 4131
rect 55956 4088 56008 4097
rect 57888 4131 57940 4140
rect 57888 4097 57897 4131
rect 57897 4097 57931 4131
rect 57931 4097 57940 4131
rect 57888 4088 57940 4097
rect 45008 3952 45060 4004
rect 49700 3952 49752 4004
rect 51908 3952 51960 4004
rect 53472 3952 53524 4004
rect 55128 3952 55180 4004
rect 55220 3952 55272 4004
rect 44916 3884 44968 3936
rect 45284 3884 45336 3936
rect 47768 3884 47820 3936
rect 51080 3884 51132 3936
rect 54576 3884 54628 3936
rect 56508 3927 56560 3936
rect 56508 3893 56517 3927
rect 56517 3893 56551 3927
rect 56551 3893 56560 3927
rect 56508 3884 56560 3893
rect 57796 3884 57848 3936
rect 8174 3782 8226 3834
rect 8238 3782 8290 3834
rect 8302 3782 8354 3834
rect 8366 3782 8418 3834
rect 8430 3782 8482 3834
rect 22622 3782 22674 3834
rect 22686 3782 22738 3834
rect 22750 3782 22802 3834
rect 22814 3782 22866 3834
rect 22878 3782 22930 3834
rect 37070 3782 37122 3834
rect 37134 3782 37186 3834
rect 37198 3782 37250 3834
rect 37262 3782 37314 3834
rect 37326 3782 37378 3834
rect 51518 3782 51570 3834
rect 51582 3782 51634 3834
rect 51646 3782 51698 3834
rect 51710 3782 51762 3834
rect 51774 3782 51826 3834
rect 2044 3723 2096 3732
rect 2044 3689 2053 3723
rect 2053 3689 2087 3723
rect 2087 3689 2096 3723
rect 2044 3680 2096 3689
rect 2412 3680 2464 3732
rect 4252 3680 4304 3732
rect 4804 3680 4856 3732
rect 7012 3680 7064 3732
rect 7472 3680 7524 3732
rect 7748 3680 7800 3732
rect 10048 3680 10100 3732
rect 13544 3723 13596 3732
rect 1400 3612 1452 3664
rect 2412 3544 2464 3596
rect 2780 3612 2832 3664
rect 2964 3655 3016 3664
rect 2964 3621 2973 3655
rect 2973 3621 3007 3655
rect 3007 3621 3016 3655
rect 2964 3612 3016 3621
rect 6552 3612 6604 3664
rect 7380 3612 7432 3664
rect 8484 3612 8536 3664
rect 10508 3612 10560 3664
rect 10876 3612 10928 3664
rect 4712 3544 4764 3596
rect 5264 3587 5316 3596
rect 5264 3553 5273 3587
rect 5273 3553 5307 3587
rect 5307 3553 5316 3587
rect 5264 3544 5316 3553
rect 7104 3544 7156 3596
rect 7748 3544 7800 3596
rect 2872 3476 2924 3528
rect 3792 3451 3844 3460
rect 3792 3417 3801 3451
rect 3801 3417 3835 3451
rect 3835 3417 3844 3451
rect 3792 3408 3844 3417
rect 4252 3519 4304 3528
rect 4252 3485 4261 3519
rect 4261 3485 4295 3519
rect 4295 3485 4304 3519
rect 5540 3519 5592 3528
rect 4252 3476 4304 3485
rect 5540 3485 5574 3519
rect 5574 3485 5592 3519
rect 5540 3476 5592 3485
rect 6920 3476 6972 3528
rect 7380 3476 7432 3528
rect 8116 3544 8168 3596
rect 8576 3544 8628 3596
rect 8852 3544 8904 3596
rect 9864 3544 9916 3596
rect 10784 3587 10836 3596
rect 10784 3553 10793 3587
rect 10793 3553 10827 3587
rect 10827 3553 10836 3587
rect 10784 3544 10836 3553
rect 13544 3689 13553 3723
rect 13553 3689 13587 3723
rect 13587 3689 13596 3723
rect 13544 3680 13596 3689
rect 15384 3723 15436 3732
rect 15384 3689 15393 3723
rect 15393 3689 15427 3723
rect 15427 3689 15436 3723
rect 15384 3680 15436 3689
rect 15844 3680 15896 3732
rect 14096 3612 14148 3664
rect 17040 3680 17092 3732
rect 22376 3680 22428 3732
rect 22468 3680 22520 3732
rect 23848 3680 23900 3732
rect 25136 3680 25188 3732
rect 26056 3680 26108 3732
rect 26884 3680 26936 3732
rect 27068 3680 27120 3732
rect 31208 3680 31260 3732
rect 32680 3723 32732 3732
rect 32680 3689 32689 3723
rect 32689 3689 32723 3723
rect 32723 3689 32732 3723
rect 32680 3680 32732 3689
rect 33324 3680 33376 3732
rect 34796 3723 34848 3732
rect 34796 3689 34805 3723
rect 34805 3689 34839 3723
rect 34839 3689 34848 3723
rect 34796 3680 34848 3689
rect 35256 3680 35308 3732
rect 11520 3587 11572 3596
rect 11520 3553 11529 3587
rect 11529 3553 11563 3587
rect 11563 3553 11572 3587
rect 11520 3544 11572 3553
rect 7288 3408 7340 3460
rect 5448 3340 5500 3392
rect 7472 3408 7524 3460
rect 8760 3476 8812 3528
rect 9496 3476 9548 3528
rect 10508 3476 10560 3528
rect 12532 3476 12584 3528
rect 13728 3476 13780 3528
rect 14372 3476 14424 3528
rect 17408 3612 17460 3664
rect 18420 3612 18472 3664
rect 21088 3612 21140 3664
rect 25320 3612 25372 3664
rect 14832 3519 14884 3528
rect 14832 3485 14841 3519
rect 14841 3485 14875 3519
rect 14875 3485 14884 3519
rect 14832 3476 14884 3485
rect 15292 3476 15344 3528
rect 15752 3476 15804 3528
rect 16304 3519 16356 3528
rect 8208 3340 8260 3392
rect 9680 3340 9732 3392
rect 9956 3340 10008 3392
rect 10692 3340 10744 3392
rect 10876 3340 10928 3392
rect 12716 3340 12768 3392
rect 16304 3485 16313 3519
rect 16313 3485 16347 3519
rect 16347 3485 16356 3519
rect 16304 3476 16356 3485
rect 16580 3476 16632 3528
rect 19892 3544 19944 3596
rect 17960 3519 18012 3528
rect 17960 3485 17969 3519
rect 17969 3485 18003 3519
rect 18003 3485 18012 3519
rect 17960 3476 18012 3485
rect 18328 3476 18380 3528
rect 19248 3519 19300 3528
rect 19248 3485 19257 3519
rect 19257 3485 19291 3519
rect 19291 3485 19300 3519
rect 19248 3476 19300 3485
rect 21364 3544 21416 3596
rect 17316 3408 17368 3460
rect 22100 3476 22152 3528
rect 23388 3476 23440 3528
rect 28264 3612 28316 3664
rect 30840 3612 30892 3664
rect 34612 3612 34664 3664
rect 37556 3680 37608 3732
rect 38660 3680 38712 3732
rect 39488 3612 39540 3664
rect 41972 3680 42024 3732
rect 44916 3680 44968 3732
rect 48044 3680 48096 3732
rect 52276 3723 52328 3732
rect 52276 3689 52285 3723
rect 52285 3689 52319 3723
rect 52319 3689 52328 3723
rect 52276 3680 52328 3689
rect 52552 3680 52604 3732
rect 56508 3680 56560 3732
rect 57796 3723 57848 3732
rect 57796 3689 57805 3723
rect 57805 3689 57839 3723
rect 57839 3689 57848 3723
rect 57796 3680 57848 3689
rect 27896 3544 27948 3596
rect 27620 3476 27672 3528
rect 27712 3476 27764 3528
rect 29552 3519 29604 3528
rect 29552 3485 29561 3519
rect 29561 3485 29595 3519
rect 29595 3485 29604 3519
rect 29552 3476 29604 3485
rect 37648 3544 37700 3596
rect 39948 3544 40000 3596
rect 32496 3476 32548 3528
rect 33140 3476 33192 3528
rect 34428 3476 34480 3528
rect 34888 3519 34940 3528
rect 34888 3485 34897 3519
rect 34897 3485 34931 3519
rect 34931 3485 34940 3519
rect 34888 3476 34940 3485
rect 35532 3519 35584 3528
rect 35532 3485 35541 3519
rect 35541 3485 35575 3519
rect 35575 3485 35584 3519
rect 35532 3476 35584 3485
rect 36728 3476 36780 3528
rect 16396 3340 16448 3392
rect 16948 3340 17000 3392
rect 17224 3383 17276 3392
rect 17224 3349 17233 3383
rect 17233 3349 17267 3383
rect 17267 3349 17276 3383
rect 17224 3340 17276 3349
rect 19892 3340 19944 3392
rect 21732 3340 21784 3392
rect 23572 3408 23624 3460
rect 22376 3340 22428 3392
rect 25228 3408 25280 3460
rect 27528 3408 27580 3460
rect 28172 3451 28224 3460
rect 28172 3417 28181 3451
rect 28181 3417 28215 3451
rect 28215 3417 28224 3451
rect 28172 3408 28224 3417
rect 31300 3408 31352 3460
rect 32864 3408 32916 3460
rect 35900 3408 35952 3460
rect 27344 3340 27396 3392
rect 31484 3340 31536 3392
rect 33508 3340 33560 3392
rect 38292 3519 38344 3528
rect 37464 3340 37516 3392
rect 38292 3485 38301 3519
rect 38301 3485 38335 3519
rect 38335 3485 38344 3519
rect 38292 3476 38344 3485
rect 38476 3476 38528 3528
rect 41328 3612 41380 3664
rect 40868 3476 40920 3528
rect 40960 3519 41012 3528
rect 40960 3485 40969 3519
rect 40969 3485 41003 3519
rect 41003 3485 41012 3519
rect 41512 3544 41564 3596
rect 46572 3587 46624 3596
rect 40960 3476 41012 3485
rect 41788 3476 41840 3528
rect 42616 3519 42668 3528
rect 38384 3408 38436 3460
rect 38568 3340 38620 3392
rect 40132 3408 40184 3460
rect 42616 3485 42625 3519
rect 42625 3485 42659 3519
rect 42659 3485 42668 3519
rect 42616 3476 42668 3485
rect 42708 3408 42760 3460
rect 43076 3476 43128 3528
rect 43720 3519 43772 3528
rect 43720 3485 43729 3519
rect 43729 3485 43763 3519
rect 43763 3485 43772 3519
rect 43720 3476 43772 3485
rect 43904 3519 43956 3528
rect 43904 3485 43913 3519
rect 43913 3485 43947 3519
rect 43947 3485 43956 3519
rect 43904 3476 43956 3485
rect 46572 3553 46581 3587
rect 46581 3553 46615 3587
rect 46615 3553 46624 3587
rect 46572 3544 46624 3553
rect 49608 3544 49660 3596
rect 44088 3519 44140 3528
rect 44088 3485 44097 3519
rect 44097 3485 44131 3519
rect 44131 3485 44140 3519
rect 44088 3476 44140 3485
rect 44640 3476 44692 3528
rect 46480 3408 46532 3460
rect 47216 3408 47268 3460
rect 41052 3383 41104 3392
rect 41052 3349 41061 3383
rect 41061 3349 41095 3383
rect 41095 3349 41104 3383
rect 41052 3340 41104 3349
rect 42892 3340 42944 3392
rect 45100 3340 45152 3392
rect 45652 3340 45704 3392
rect 48320 3408 48372 3460
rect 54024 3612 54076 3664
rect 55404 3612 55456 3664
rect 53288 3587 53340 3596
rect 53288 3553 53297 3587
rect 53297 3553 53331 3587
rect 53331 3553 53340 3587
rect 53288 3544 53340 3553
rect 52828 3476 52880 3528
rect 53104 3476 53156 3528
rect 51356 3408 51408 3460
rect 53932 3476 53984 3528
rect 54392 3519 54444 3528
rect 54392 3485 54401 3519
rect 54401 3485 54435 3519
rect 54435 3485 54444 3519
rect 54392 3476 54444 3485
rect 54576 3519 54628 3528
rect 54576 3485 54585 3519
rect 54585 3485 54619 3519
rect 54619 3485 54628 3519
rect 54576 3476 54628 3485
rect 52368 3340 52420 3392
rect 15398 3238 15450 3290
rect 15462 3238 15514 3290
rect 15526 3238 15578 3290
rect 15590 3238 15642 3290
rect 15654 3238 15706 3290
rect 29846 3238 29898 3290
rect 29910 3238 29962 3290
rect 29974 3238 30026 3290
rect 30038 3238 30090 3290
rect 30102 3238 30154 3290
rect 44294 3238 44346 3290
rect 44358 3238 44410 3290
rect 44422 3238 44474 3290
rect 44486 3238 44538 3290
rect 44550 3238 44602 3290
rect 1768 3136 1820 3188
rect 3792 3136 3844 3188
rect 5816 3136 5868 3188
rect 6460 3179 6512 3188
rect 6460 3145 6469 3179
rect 6469 3145 6503 3179
rect 6503 3145 6512 3179
rect 6460 3136 6512 3145
rect 7104 3179 7156 3188
rect 7104 3145 7113 3179
rect 7113 3145 7147 3179
rect 7147 3145 7156 3179
rect 7104 3136 7156 3145
rect 7472 3136 7524 3188
rect 1952 3068 2004 3120
rect 7380 3068 7432 3120
rect 1492 3000 1544 3052
rect 2964 3043 3016 3052
rect 2964 3009 2973 3043
rect 2973 3009 3007 3043
rect 3007 3009 3016 3043
rect 2964 3000 3016 3009
rect 3332 3000 3384 3052
rect 3884 3043 3936 3052
rect 3884 3009 3893 3043
rect 3893 3009 3927 3043
rect 3927 3009 3936 3043
rect 3884 3000 3936 3009
rect 4436 3000 4488 3052
rect 4620 3000 4672 3052
rect 5080 3043 5132 3052
rect 5080 3009 5089 3043
rect 5089 3009 5123 3043
rect 5123 3009 5132 3043
rect 5080 3000 5132 3009
rect 6828 3000 6880 3052
rect 9496 3136 9548 3188
rect 10692 3136 10744 3188
rect 11520 3136 11572 3188
rect 12624 3136 12676 3188
rect 2780 2864 2832 2916
rect 7380 2864 7432 2916
rect 8116 3068 8168 3120
rect 8668 3068 8720 3120
rect 8760 3043 8812 3052
rect 8760 3009 8769 3043
rect 8769 3009 8803 3043
rect 8803 3009 8812 3043
rect 8760 3000 8812 3009
rect 9220 3068 9272 3120
rect 14188 3136 14240 3188
rect 16948 3136 17000 3188
rect 17500 3136 17552 3188
rect 22192 3179 22244 3188
rect 22192 3145 22201 3179
rect 22201 3145 22235 3179
rect 22235 3145 22244 3179
rect 22192 3136 22244 3145
rect 25228 3179 25280 3188
rect 25228 3145 25237 3179
rect 25237 3145 25271 3179
rect 25271 3145 25280 3179
rect 25228 3136 25280 3145
rect 25504 3136 25556 3188
rect 25872 3136 25924 3188
rect 29000 3136 29052 3188
rect 33784 3179 33836 3188
rect 33784 3145 33793 3179
rect 33793 3145 33827 3179
rect 33827 3145 33836 3179
rect 33784 3136 33836 3145
rect 9404 3000 9456 3052
rect 9220 2932 9272 2984
rect 11704 3000 11756 3052
rect 10600 2932 10652 2984
rect 10784 2932 10836 2984
rect 8484 2864 8536 2916
rect 8760 2864 8812 2916
rect 8852 2864 8904 2916
rect 9588 2864 9640 2916
rect 11428 2864 11480 2916
rect 14372 3068 14424 3120
rect 15108 3068 15160 3120
rect 15936 3111 15988 3120
rect 15936 3077 15945 3111
rect 15945 3077 15979 3111
rect 15979 3077 15988 3111
rect 15936 3068 15988 3077
rect 18788 3068 18840 3120
rect 19064 3111 19116 3120
rect 13176 3000 13228 3052
rect 13728 3043 13780 3052
rect 13728 3009 13737 3043
rect 13737 3009 13771 3043
rect 13771 3009 13780 3043
rect 13728 3000 13780 3009
rect 14556 3000 14608 3052
rect 15292 3000 15344 3052
rect 16028 3000 16080 3052
rect 16580 3000 16632 3052
rect 17316 3043 17368 3052
rect 17316 3009 17325 3043
rect 17325 3009 17359 3043
rect 17359 3009 17368 3043
rect 17316 3000 17368 3009
rect 18052 3000 18104 3052
rect 19064 3077 19073 3111
rect 19073 3077 19107 3111
rect 19107 3077 19116 3111
rect 19064 3068 19116 3077
rect 19524 3111 19576 3120
rect 19524 3077 19533 3111
rect 19533 3077 19567 3111
rect 19567 3077 19576 3111
rect 19524 3068 19576 3077
rect 22100 3068 22152 3120
rect 23112 3068 23164 3120
rect 21824 3043 21876 3052
rect 21824 3009 21833 3043
rect 21833 3009 21867 3043
rect 21867 3009 21876 3043
rect 21824 3000 21876 3009
rect 21916 3000 21968 3052
rect 23020 3043 23072 3052
rect 23020 3009 23029 3043
rect 23029 3009 23063 3043
rect 23063 3009 23072 3043
rect 23020 3000 23072 3009
rect 24584 3000 24636 3052
rect 25504 3043 25556 3052
rect 25504 3009 25513 3043
rect 25513 3009 25547 3043
rect 25547 3009 25556 3043
rect 25504 3000 25556 3009
rect 27528 3068 27580 3120
rect 28172 3068 28224 3120
rect 30472 3068 30524 3120
rect 25688 3043 25740 3052
rect 25688 3009 25697 3043
rect 25697 3009 25731 3043
rect 25731 3009 25740 3043
rect 25688 3000 25740 3009
rect 25872 3043 25924 3052
rect 25872 3009 25881 3043
rect 25881 3009 25915 3043
rect 25915 3009 25924 3043
rect 27712 3043 27764 3052
rect 25872 3000 25924 3009
rect 27712 3009 27721 3043
rect 27721 3009 27755 3043
rect 27755 3009 27764 3043
rect 27712 3000 27764 3009
rect 29276 3043 29328 3052
rect 29276 3009 29285 3043
rect 29285 3009 29319 3043
rect 29319 3009 29328 3043
rect 29276 3000 29328 3009
rect 30840 3043 30892 3052
rect 30840 3009 30849 3043
rect 30849 3009 30883 3043
rect 30883 3009 30892 3043
rect 30840 3000 30892 3009
rect 31024 3046 31076 3055
rect 31024 3012 31033 3046
rect 31033 3012 31067 3046
rect 31067 3012 31076 3046
rect 31024 3003 31076 3012
rect 31300 3068 31352 3120
rect 32220 3068 32272 3120
rect 32496 3111 32548 3120
rect 32496 3077 32505 3111
rect 32505 3077 32539 3111
rect 32539 3077 32548 3111
rect 32496 3068 32548 3077
rect 31208 3043 31260 3052
rect 31208 3009 31217 3043
rect 31217 3009 31251 3043
rect 31251 3009 31260 3043
rect 31208 3000 31260 3009
rect 31576 3000 31628 3052
rect 34888 3136 34940 3188
rect 36728 3179 36780 3188
rect 36728 3145 36737 3179
rect 36737 3145 36771 3179
rect 36771 3145 36780 3179
rect 36728 3136 36780 3145
rect 36820 3136 36872 3188
rect 34520 3068 34572 3120
rect 35532 3068 35584 3120
rect 34796 3000 34848 3052
rect 13636 2932 13688 2984
rect 14924 2932 14976 2984
rect 3240 2839 3292 2848
rect 3240 2805 3249 2839
rect 3249 2805 3283 2839
rect 3283 2805 3292 2839
rect 3240 2796 3292 2805
rect 10416 2796 10468 2848
rect 10968 2839 11020 2848
rect 10968 2805 10977 2839
rect 10977 2805 11011 2839
rect 11011 2805 11020 2839
rect 10968 2796 11020 2805
rect 11336 2796 11388 2848
rect 19340 2932 19392 2984
rect 15936 2907 15988 2916
rect 15936 2873 15945 2907
rect 15945 2873 15979 2907
rect 15979 2873 15988 2907
rect 15936 2864 15988 2873
rect 17776 2864 17828 2916
rect 24308 2932 24360 2984
rect 28724 2932 28776 2984
rect 29092 2932 29144 2984
rect 29368 2932 29420 2984
rect 30748 2932 30800 2984
rect 31300 2932 31352 2984
rect 32312 2932 32364 2984
rect 36820 3000 36872 3052
rect 39948 3136 40000 3188
rect 41052 3136 41104 3188
rect 43904 3136 43956 3188
rect 43996 3136 44048 3188
rect 45008 3136 45060 3188
rect 45836 3136 45888 3188
rect 37464 3043 37516 3052
rect 37464 3009 37473 3043
rect 37473 3009 37507 3043
rect 37507 3009 37516 3043
rect 37648 3043 37700 3052
rect 37464 3000 37516 3009
rect 37648 3009 37657 3043
rect 37657 3009 37691 3043
rect 37691 3009 37700 3043
rect 37648 3000 37700 3009
rect 37740 3043 37792 3052
rect 37740 3009 37749 3043
rect 37749 3009 37783 3043
rect 37783 3009 37792 3043
rect 37740 3000 37792 3009
rect 35808 2932 35860 2984
rect 35900 2932 35952 2984
rect 40776 3043 40828 3052
rect 40776 3009 40785 3043
rect 40785 3009 40819 3043
rect 40819 3009 40828 3043
rect 40776 3000 40828 3009
rect 41052 3043 41104 3052
rect 41052 3009 41061 3043
rect 41061 3009 41095 3043
rect 41095 3009 41104 3043
rect 41052 3000 41104 3009
rect 42892 3068 42944 3120
rect 43812 3111 43864 3120
rect 42616 3000 42668 3052
rect 43812 3077 43821 3111
rect 43821 3077 43855 3111
rect 43855 3077 43864 3111
rect 43812 3068 43864 3077
rect 45100 3068 45152 3120
rect 49424 3068 49476 3120
rect 38292 2932 38344 2984
rect 39672 2932 39724 2984
rect 42708 2932 42760 2984
rect 43628 3000 43680 3052
rect 44180 3000 44232 3052
rect 45008 3000 45060 3052
rect 47584 2975 47636 2984
rect 47584 2941 47593 2975
rect 47593 2941 47627 2975
rect 47627 2941 47636 2975
rect 47584 2932 47636 2941
rect 49608 3000 49660 3052
rect 52828 3136 52880 3188
rect 57796 3136 57848 3188
rect 22284 2864 22336 2916
rect 25320 2864 25372 2916
rect 25504 2864 25556 2916
rect 25780 2864 25832 2916
rect 25964 2864 26016 2916
rect 31208 2864 31260 2916
rect 13452 2796 13504 2848
rect 16028 2796 16080 2848
rect 16212 2796 16264 2848
rect 17960 2839 18012 2848
rect 17960 2805 17969 2839
rect 17969 2805 18003 2839
rect 18003 2805 18012 2839
rect 17960 2796 18012 2805
rect 21548 2796 21600 2848
rect 22008 2796 22060 2848
rect 22468 2796 22520 2848
rect 26792 2796 26844 2848
rect 31760 2864 31812 2916
rect 35348 2864 35400 2916
rect 33968 2796 34020 2848
rect 34244 2796 34296 2848
rect 35532 2796 35584 2848
rect 39488 2839 39540 2848
rect 39488 2805 39497 2839
rect 39497 2805 39531 2839
rect 39531 2805 39540 2839
rect 39488 2796 39540 2805
rect 39672 2796 39724 2848
rect 43260 2864 43312 2916
rect 45284 2864 45336 2916
rect 45744 2864 45796 2916
rect 50160 2864 50212 2916
rect 52368 3000 52420 3052
rect 52828 3000 52880 3052
rect 53104 3000 53156 3052
rect 53932 3000 53984 3052
rect 54116 3043 54168 3052
rect 54116 3009 54125 3043
rect 54125 3009 54159 3043
rect 54159 3009 54168 3043
rect 54116 3000 54168 3009
rect 54760 3043 54812 3052
rect 54760 3009 54769 3043
rect 54769 3009 54803 3043
rect 54803 3009 54812 3043
rect 54760 3000 54812 3009
rect 41696 2796 41748 2848
rect 44548 2796 44600 2848
rect 44916 2839 44968 2848
rect 44916 2805 44925 2839
rect 44925 2805 44959 2839
rect 44959 2805 44968 2839
rect 44916 2796 44968 2805
rect 45652 2796 45704 2848
rect 46204 2839 46256 2848
rect 46204 2805 46213 2839
rect 46213 2805 46247 2839
rect 46247 2805 46256 2839
rect 46204 2796 46256 2805
rect 46848 2839 46900 2848
rect 46848 2805 46857 2839
rect 46857 2805 46891 2839
rect 46891 2805 46900 2839
rect 46848 2796 46900 2805
rect 48780 2796 48832 2848
rect 49332 2796 49384 2848
rect 49976 2839 50028 2848
rect 49976 2805 49985 2839
rect 49985 2805 50019 2839
rect 50019 2805 50028 2839
rect 49976 2796 50028 2805
rect 52460 2864 52512 2916
rect 53840 2864 53892 2916
rect 52184 2796 52236 2848
rect 8174 2694 8226 2746
rect 8238 2694 8290 2746
rect 8302 2694 8354 2746
rect 8366 2694 8418 2746
rect 8430 2694 8482 2746
rect 22622 2694 22674 2746
rect 22686 2694 22738 2746
rect 22750 2694 22802 2746
rect 22814 2694 22866 2746
rect 22878 2694 22930 2746
rect 37070 2694 37122 2746
rect 37134 2694 37186 2746
rect 37198 2694 37250 2746
rect 37262 2694 37314 2746
rect 37326 2694 37378 2746
rect 51518 2694 51570 2746
rect 51582 2694 51634 2746
rect 51646 2694 51698 2746
rect 51710 2694 51762 2746
rect 51774 2694 51826 2746
rect 1952 2592 2004 2644
rect 2964 2592 3016 2644
rect 4344 2592 4396 2644
rect 5816 2592 5868 2644
rect 6736 2592 6788 2644
rect 3608 2524 3660 2576
rect 6552 2524 6604 2576
rect 2228 2499 2280 2508
rect 2228 2465 2237 2499
rect 2237 2465 2271 2499
rect 2271 2465 2280 2499
rect 2228 2456 2280 2465
rect 2320 2456 2372 2508
rect 6920 2524 6972 2576
rect 3976 2431 4028 2440
rect 1676 2320 1728 2372
rect 3976 2397 3985 2431
rect 3985 2397 4019 2431
rect 4019 2397 4028 2431
rect 3976 2388 4028 2397
rect 5264 2388 5316 2440
rect 5540 2363 5592 2372
rect 5540 2329 5558 2363
rect 5558 2329 5592 2363
rect 5540 2320 5592 2329
rect 2596 2252 2648 2304
rect 7104 2456 7156 2508
rect 8116 2592 8168 2644
rect 8300 2524 8352 2576
rect 9220 2524 9272 2576
rect 10968 2592 11020 2644
rect 17776 2592 17828 2644
rect 21548 2592 21600 2644
rect 22100 2592 22152 2644
rect 27896 2592 27948 2644
rect 13820 2524 13872 2576
rect 15660 2524 15712 2576
rect 16212 2524 16264 2576
rect 9496 2456 9548 2508
rect 13268 2456 13320 2508
rect 7196 2388 7248 2440
rect 7472 2388 7524 2440
rect 8116 2388 8168 2440
rect 9036 2388 9088 2440
rect 9220 2431 9272 2440
rect 9220 2397 9229 2431
rect 9229 2397 9263 2431
rect 9263 2397 9272 2431
rect 9220 2388 9272 2397
rect 6736 2252 6788 2304
rect 10692 2431 10744 2440
rect 10692 2397 10701 2431
rect 10701 2397 10735 2431
rect 10735 2397 10744 2431
rect 10692 2388 10744 2397
rect 10968 2431 11020 2440
rect 10968 2397 10977 2431
rect 10977 2397 11011 2431
rect 11011 2397 11020 2431
rect 10968 2388 11020 2397
rect 11612 2388 11664 2440
rect 11796 2431 11848 2440
rect 11796 2397 11805 2431
rect 11805 2397 11839 2431
rect 11839 2397 11848 2431
rect 11796 2388 11848 2397
rect 13544 2431 13596 2440
rect 13544 2397 13553 2431
rect 13553 2397 13587 2431
rect 13587 2397 13596 2431
rect 13544 2388 13596 2397
rect 14372 2431 14424 2440
rect 14372 2397 14381 2431
rect 14381 2397 14415 2431
rect 14415 2397 14424 2431
rect 14372 2388 14424 2397
rect 14556 2388 14608 2440
rect 17592 2456 17644 2508
rect 17224 2431 17276 2440
rect 17224 2397 17233 2431
rect 17233 2397 17267 2431
rect 17267 2397 17276 2431
rect 17224 2388 17276 2397
rect 17684 2431 17736 2440
rect 17684 2397 17693 2431
rect 17693 2397 17727 2431
rect 17727 2397 17736 2431
rect 17684 2388 17736 2397
rect 18696 2388 18748 2440
rect 11336 2320 11388 2372
rect 21272 2524 21324 2576
rect 29552 2592 29604 2644
rect 31024 2592 31076 2644
rect 30656 2524 30708 2576
rect 20260 2431 20312 2440
rect 20260 2397 20269 2431
rect 20269 2397 20303 2431
rect 20303 2397 20312 2431
rect 20260 2388 20312 2397
rect 20536 2431 20588 2440
rect 20536 2397 20545 2431
rect 20545 2397 20579 2431
rect 20579 2397 20588 2431
rect 20536 2388 20588 2397
rect 21180 2388 21232 2440
rect 21824 2431 21876 2440
rect 21824 2397 21833 2431
rect 21833 2397 21867 2431
rect 21867 2397 21876 2431
rect 21824 2388 21876 2397
rect 22008 2431 22060 2440
rect 22008 2397 22017 2431
rect 22017 2397 22051 2431
rect 22051 2397 22060 2431
rect 22008 2388 22060 2397
rect 22100 2388 22152 2440
rect 23572 2456 23624 2508
rect 29736 2456 29788 2508
rect 30932 2456 30984 2508
rect 9220 2252 9272 2304
rect 20904 2320 20956 2372
rect 24400 2388 24452 2440
rect 24676 2431 24728 2440
rect 24676 2397 24685 2431
rect 24685 2397 24719 2431
rect 24719 2397 24728 2431
rect 24676 2388 24728 2397
rect 26976 2431 27028 2440
rect 26976 2397 26985 2431
rect 26985 2397 27019 2431
rect 27019 2397 27028 2431
rect 26976 2388 27028 2397
rect 30196 2388 30248 2440
rect 30380 2388 30432 2440
rect 33508 2592 33560 2644
rect 33968 2635 34020 2644
rect 33968 2601 33977 2635
rect 33977 2601 34011 2635
rect 34011 2601 34020 2635
rect 33968 2592 34020 2601
rect 35348 2635 35400 2644
rect 35348 2601 35357 2635
rect 35357 2601 35391 2635
rect 35391 2601 35400 2635
rect 35348 2592 35400 2601
rect 36912 2592 36964 2644
rect 37096 2592 37148 2644
rect 32036 2524 32088 2576
rect 32864 2524 32916 2576
rect 31484 2456 31536 2508
rect 36452 2524 36504 2576
rect 43720 2592 43772 2644
rect 31576 2431 31628 2440
rect 31576 2397 31585 2431
rect 31585 2397 31619 2431
rect 31619 2397 31628 2431
rect 31576 2388 31628 2397
rect 33232 2431 33284 2440
rect 33232 2397 33241 2431
rect 33241 2397 33275 2431
rect 33275 2397 33284 2431
rect 33232 2388 33284 2397
rect 33600 2388 33652 2440
rect 33692 2388 33744 2440
rect 39212 2499 39264 2508
rect 39212 2465 39221 2499
rect 39221 2465 39255 2499
rect 39255 2465 39264 2499
rect 39212 2456 39264 2465
rect 39488 2456 39540 2508
rect 46572 2592 46624 2644
rect 49516 2592 49568 2644
rect 57888 2592 57940 2644
rect 50344 2524 50396 2576
rect 50896 2524 50948 2576
rect 42708 2456 42760 2508
rect 52092 2499 52144 2508
rect 52092 2465 52101 2499
rect 52101 2465 52135 2499
rect 52135 2465 52144 2499
rect 52092 2456 52144 2465
rect 39856 2431 39908 2440
rect 14556 2295 14608 2304
rect 14556 2261 14565 2295
rect 14565 2261 14599 2295
rect 14599 2261 14608 2295
rect 14556 2252 14608 2261
rect 15292 2295 15344 2304
rect 15292 2261 15301 2295
rect 15301 2261 15335 2295
rect 15335 2261 15344 2295
rect 15292 2252 15344 2261
rect 16028 2295 16080 2304
rect 16028 2261 16037 2295
rect 16037 2261 16071 2295
rect 16071 2261 16080 2295
rect 16028 2252 16080 2261
rect 17684 2252 17736 2304
rect 19524 2295 19576 2304
rect 19524 2261 19533 2295
rect 19533 2261 19567 2295
rect 19567 2261 19576 2295
rect 29000 2320 29052 2372
rect 33324 2320 33376 2372
rect 19524 2252 19576 2261
rect 21824 2252 21876 2304
rect 22836 2252 22888 2304
rect 22928 2252 22980 2304
rect 26976 2252 27028 2304
rect 31300 2252 31352 2304
rect 32588 2252 32640 2304
rect 39856 2397 39865 2431
rect 39865 2397 39899 2431
rect 39899 2397 39908 2431
rect 39856 2388 39908 2397
rect 40500 2431 40552 2440
rect 40500 2397 40509 2431
rect 40509 2397 40543 2431
rect 40543 2397 40552 2431
rect 40500 2388 40552 2397
rect 43076 2431 43128 2440
rect 43076 2397 43085 2431
rect 43085 2397 43119 2431
rect 43119 2397 43128 2431
rect 43076 2388 43128 2397
rect 43720 2431 43772 2440
rect 43720 2397 43729 2431
rect 43729 2397 43763 2431
rect 43763 2397 43772 2431
rect 43720 2388 43772 2397
rect 43904 2388 43956 2440
rect 38016 2320 38068 2372
rect 45100 2320 45152 2372
rect 48228 2431 48280 2440
rect 48228 2397 48237 2431
rect 48237 2397 48271 2431
rect 48271 2397 48280 2431
rect 48228 2388 48280 2397
rect 48872 2431 48924 2440
rect 48872 2397 48881 2431
rect 48881 2397 48915 2431
rect 48915 2397 48924 2431
rect 48872 2388 48924 2397
rect 49516 2431 49568 2440
rect 49516 2397 49525 2431
rect 49525 2397 49559 2431
rect 49559 2397 49568 2431
rect 49516 2388 49568 2397
rect 50160 2431 50212 2440
rect 50160 2397 50169 2431
rect 50169 2397 50203 2431
rect 50203 2397 50212 2431
rect 50160 2388 50212 2397
rect 50804 2431 50856 2440
rect 50804 2397 50813 2431
rect 50813 2397 50847 2431
rect 50847 2397 50856 2431
rect 50804 2388 50856 2397
rect 51448 2431 51500 2440
rect 51448 2397 51457 2431
rect 51457 2397 51491 2431
rect 51491 2397 51500 2431
rect 51448 2388 51500 2397
rect 49424 2320 49476 2372
rect 52276 2388 52328 2440
rect 53380 2431 53432 2440
rect 53380 2397 53389 2431
rect 53389 2397 53423 2431
rect 53423 2397 53432 2431
rect 53380 2388 53432 2397
rect 54024 2431 54076 2440
rect 54024 2397 54033 2431
rect 54033 2397 54067 2431
rect 54067 2397 54076 2431
rect 54024 2388 54076 2397
rect 41788 2295 41840 2304
rect 41788 2261 41797 2295
rect 41797 2261 41831 2295
rect 41831 2261 41840 2295
rect 41788 2252 41840 2261
rect 46756 2252 46808 2304
rect 49056 2252 49108 2304
rect 49148 2252 49200 2304
rect 54668 2295 54720 2304
rect 54668 2261 54677 2295
rect 54677 2261 54711 2295
rect 54711 2261 54720 2295
rect 54668 2252 54720 2261
rect 57888 2295 57940 2304
rect 57888 2261 57897 2295
rect 57897 2261 57931 2295
rect 57931 2261 57940 2295
rect 57888 2252 57940 2261
rect 15398 2150 15450 2202
rect 15462 2150 15514 2202
rect 15526 2150 15578 2202
rect 15590 2150 15642 2202
rect 15654 2150 15706 2202
rect 29846 2150 29898 2202
rect 29910 2150 29962 2202
rect 29974 2150 30026 2202
rect 30038 2150 30090 2202
rect 30102 2150 30154 2202
rect 44294 2150 44346 2202
rect 44358 2150 44410 2202
rect 44422 2150 44474 2202
rect 44486 2150 44538 2202
rect 44550 2150 44602 2202
rect 6920 2048 6972 2100
rect 9220 2048 9272 2100
rect 20076 2048 20128 2100
rect 2136 1980 2188 2032
rect 14372 1980 14424 2032
rect 15292 1980 15344 2032
rect 20444 1980 20496 2032
rect 21088 2048 21140 2100
rect 24676 2048 24728 2100
rect 32036 2048 32088 2100
rect 33324 2048 33376 2100
rect 35072 2048 35124 2100
rect 40500 2048 40552 2100
rect 40868 2048 40920 2100
rect 42708 2048 42760 2100
rect 44732 2048 44784 2100
rect 45192 2048 45244 2100
rect 45284 2048 45336 2100
rect 53380 2048 53432 2100
rect 26240 1980 26292 2032
rect 33232 1980 33284 2032
rect 6552 1912 6604 1964
rect 8300 1912 8352 1964
rect 8760 1912 8812 1964
rect 9496 1912 9548 1964
rect 2780 1844 2832 1896
rect 8116 1844 8168 1896
rect 3516 1776 3568 1828
rect 14464 1912 14516 1964
rect 14556 1912 14608 1964
rect 19616 1912 19668 1964
rect 34796 1912 34848 1964
rect 36728 1980 36780 2032
rect 43076 1980 43128 2032
rect 44456 1980 44508 2032
rect 51448 1980 51500 2032
rect 53288 1980 53340 2032
rect 57888 1980 57940 2032
rect 13544 1844 13596 1896
rect 26148 1844 26200 1896
rect 14924 1776 14976 1828
rect 15292 1776 15344 1828
rect 5172 1708 5224 1760
rect 7104 1708 7156 1760
rect 7840 1708 7892 1760
rect 8760 1708 8812 1760
rect 10784 1708 10836 1760
rect 11612 1708 11664 1760
rect 3148 1640 3200 1692
rect 14096 1708 14148 1760
rect 14648 1708 14700 1760
rect 19524 1776 19576 1828
rect 37648 1912 37700 1964
rect 41420 1912 41472 1964
rect 48228 1912 48280 1964
rect 50344 1912 50396 1964
rect 56416 1912 56468 1964
rect 38660 1844 38712 1896
rect 45100 1844 45152 1896
rect 46112 1844 46164 1896
rect 54024 1844 54076 1896
rect 39856 1776 39908 1828
rect 43628 1776 43680 1828
rect 50804 1776 50856 1828
rect 49056 1708 49108 1760
rect 53840 1708 53892 1760
rect 54668 1708 54720 1760
rect 18144 1640 18196 1692
rect 31392 1640 31444 1692
rect 44180 1640 44232 1692
rect 44824 1640 44876 1692
rect 46664 1640 46716 1692
rect 52276 1640 52328 1692
rect 19248 1572 19300 1624
rect 27712 1572 27764 1624
rect 7472 1504 7524 1556
rect 8208 1504 8260 1556
rect 9680 1504 9732 1556
rect 10508 1504 10560 1556
rect 10600 1504 10652 1556
rect 39764 1504 39816 1556
rect 45652 1504 45704 1556
rect 7012 1368 7064 1420
rect 7472 1368 7524 1420
rect 8024 1436 8076 1488
rect 8852 1436 8904 1488
rect 9588 1436 9640 1488
rect 16028 1436 16080 1488
rect 20168 1436 20220 1488
rect 37280 1436 37332 1488
rect 38292 1436 38344 1488
rect 39212 1436 39264 1488
rect 44916 1436 44968 1488
rect 49976 1436 50028 1488
rect 54760 1436 54812 1488
rect 10968 1368 11020 1420
rect 13452 1368 13504 1420
rect 17132 1368 17184 1420
rect 24032 1368 24084 1420
rect 29460 1368 29512 1420
rect 36176 1368 36228 1420
rect 37096 1368 37148 1420
rect 41144 1368 41196 1420
rect 46848 1368 46900 1420
rect 7932 1300 7984 1352
rect 10416 1300 10468 1352
rect 10508 1300 10560 1352
rect 20536 1300 20588 1352
rect 53288 1300 53340 1352
rect 7288 1232 7340 1284
rect 7840 1232 7892 1284
rect 20260 1232 20312 1284
rect 52644 1232 52696 1284
rect 6092 1164 6144 1216
rect 8576 1164 8628 1216
rect 5908 1096 5960 1148
rect 33784 1164 33836 1216
rect 38936 1164 38988 1216
rect 43720 1164 43772 1216
rect 10416 1096 10468 1148
rect 25320 1096 25372 1148
rect 26884 1096 26936 1148
rect 40132 1096 40184 1148
rect 4896 1028 4948 1080
rect 8392 1028 8444 1080
rect 18880 1028 18932 1080
rect 35440 1028 35492 1080
rect 4528 960 4580 1012
rect 8208 960 8260 1012
rect 14832 960 14884 1012
rect 29644 960 29696 1012
rect 13176 892 13228 944
rect 26332 892 26384 944
rect 26424 892 26476 944
rect 26608 892 26660 944
rect 3240 756 3292 808
rect 7196 688 7248 740
<< metal2 >>
rect 3974 19200 4030 20000
rect 4434 19200 4490 20000
rect 4894 19200 4950 20000
rect 5354 19200 5410 20000
rect 5814 19200 5870 20000
rect 6274 19200 6330 20000
rect 6734 19200 6790 20000
rect 7194 19200 7250 20000
rect 7654 19200 7710 20000
rect 8114 19200 8170 20000
rect 8574 19200 8630 20000
rect 9034 19200 9090 20000
rect 9494 19200 9550 20000
rect 9954 19200 10010 20000
rect 10414 19200 10470 20000
rect 10874 19200 10930 20000
rect 11334 19200 11390 20000
rect 11794 19200 11850 20000
rect 12254 19200 12310 20000
rect 12714 19200 12770 20000
rect 13174 19200 13230 20000
rect 13634 19200 13690 20000
rect 14094 19200 14150 20000
rect 14554 19200 14610 20000
rect 15014 19200 15070 20000
rect 15474 19200 15530 20000
rect 15934 19200 15990 20000
rect 16394 19200 16450 20000
rect 16854 19200 16910 20000
rect 17314 19200 17370 20000
rect 17774 19200 17830 20000
rect 18234 19200 18290 20000
rect 18694 19200 18750 20000
rect 19154 19200 19210 20000
rect 19614 19200 19670 20000
rect 20074 19200 20130 20000
rect 20534 19200 20590 20000
rect 20994 19200 21050 20000
rect 21454 19200 21510 20000
rect 21914 19200 21970 20000
rect 22374 19200 22430 20000
rect 22834 19200 22890 20000
rect 23294 19200 23350 20000
rect 23754 19200 23810 20000
rect 24214 19200 24270 20000
rect 24674 19200 24730 20000
rect 25134 19200 25190 20000
rect 25594 19200 25650 20000
rect 26054 19200 26110 20000
rect 26514 19200 26570 20000
rect 26974 19200 27030 20000
rect 27434 19200 27490 20000
rect 27894 19200 27950 20000
rect 28354 19200 28410 20000
rect 28814 19200 28870 20000
rect 29274 19200 29330 20000
rect 29734 19200 29790 20000
rect 30194 19200 30250 20000
rect 30654 19200 30710 20000
rect 31114 19200 31170 20000
rect 31574 19200 31630 20000
rect 32034 19200 32090 20000
rect 32494 19200 32550 20000
rect 32954 19200 33010 20000
rect 33414 19200 33470 20000
rect 33874 19200 33930 20000
rect 34334 19200 34390 20000
rect 34794 19200 34850 20000
rect 35254 19200 35310 20000
rect 35714 19200 35770 20000
rect 36174 19200 36230 20000
rect 36634 19200 36690 20000
rect 37094 19200 37150 20000
rect 37554 19200 37610 20000
rect 38014 19200 38070 20000
rect 38474 19200 38530 20000
rect 38934 19200 38990 20000
rect 39394 19200 39450 20000
rect 39854 19200 39910 20000
rect 40314 19200 40370 20000
rect 40774 19200 40830 20000
rect 41234 19200 41290 20000
rect 41694 19200 41750 20000
rect 42154 19200 42210 20000
rect 42614 19200 42670 20000
rect 43074 19200 43130 20000
rect 43534 19200 43590 20000
rect 43994 19200 44050 20000
rect 44454 19200 44510 20000
rect 44914 19200 44970 20000
rect 45374 19200 45430 20000
rect 45834 19200 45890 20000
rect 46294 19200 46350 20000
rect 46754 19200 46810 20000
rect 47214 19200 47270 20000
rect 47674 19200 47730 20000
rect 48134 19200 48190 20000
rect 48594 19200 48650 20000
rect 49054 19200 49110 20000
rect 49514 19200 49570 20000
rect 49974 19200 50030 20000
rect 50434 19200 50490 20000
rect 50894 19200 50950 20000
rect 51354 19200 51410 20000
rect 51814 19200 51870 20000
rect 52274 19200 52330 20000
rect 52734 19200 52790 20000
rect 53194 19200 53250 20000
rect 53654 19200 53710 20000
rect 54114 19200 54170 20000
rect 54574 19200 54630 20000
rect 55034 19200 55090 20000
rect 55494 19200 55550 20000
rect 55954 19200 56010 20000
rect 4448 17202 4476 19200
rect 4908 17202 4936 19200
rect 5828 17202 5856 19200
rect 4436 17196 4488 17202
rect 4436 17138 4488 17144
rect 4896 17196 4948 17202
rect 4896 17138 4948 17144
rect 5816 17196 5868 17202
rect 5816 17138 5868 17144
rect 6288 16794 6316 19200
rect 7208 17202 7236 19200
rect 7668 17202 7696 19200
rect 8588 17202 8616 19200
rect 9048 17202 9076 19200
rect 9968 17202 9996 19200
rect 10428 17202 10456 19200
rect 7196 17196 7248 17202
rect 7196 17138 7248 17144
rect 7656 17196 7708 17202
rect 7656 17138 7708 17144
rect 8576 17196 8628 17202
rect 8576 17138 8628 17144
rect 9036 17196 9088 17202
rect 9036 17138 9088 17144
rect 9956 17196 10008 17202
rect 9956 17138 10008 17144
rect 10416 17196 10468 17202
rect 10416 17138 10468 17144
rect 8174 16892 8482 16901
rect 8174 16890 8180 16892
rect 8236 16890 8260 16892
rect 8316 16890 8340 16892
rect 8396 16890 8420 16892
rect 8476 16890 8482 16892
rect 8236 16838 8238 16890
rect 8418 16838 8420 16890
rect 8174 16836 8180 16838
rect 8236 16836 8260 16838
rect 8316 16836 8340 16838
rect 8396 16836 8420 16838
rect 8476 16836 8482 16838
rect 8174 16827 8482 16836
rect 11348 16794 11376 19200
rect 11808 17202 11836 19200
rect 12728 17202 12756 19200
rect 13188 17202 13216 19200
rect 11796 17196 11848 17202
rect 11796 17138 11848 17144
rect 12716 17196 12768 17202
rect 12716 17138 12768 17144
rect 13176 17196 13228 17202
rect 13176 17138 13228 17144
rect 14108 16794 14136 19200
rect 14568 17202 14596 19200
rect 15488 17626 15516 19200
rect 15304 17598 15516 17626
rect 15304 17202 15332 17598
rect 15398 17436 15706 17445
rect 15398 17434 15404 17436
rect 15460 17434 15484 17436
rect 15540 17434 15564 17436
rect 15620 17434 15644 17436
rect 15700 17434 15706 17436
rect 15460 17382 15462 17434
rect 15642 17382 15644 17434
rect 15398 17380 15404 17382
rect 15460 17380 15484 17382
rect 15540 17380 15564 17382
rect 15620 17380 15644 17382
rect 15700 17380 15706 17382
rect 15398 17371 15706 17380
rect 15948 17202 15976 19200
rect 14556 17196 14608 17202
rect 14556 17138 14608 17144
rect 15292 17196 15344 17202
rect 15292 17138 15344 17144
rect 15936 17196 15988 17202
rect 15936 17138 15988 17144
rect 16868 16794 16896 19200
rect 17328 17202 17356 19200
rect 18248 17202 18276 19200
rect 18708 17202 18736 19200
rect 19628 17202 19656 19200
rect 20088 17202 20116 19200
rect 17316 17196 17368 17202
rect 17316 17138 17368 17144
rect 18236 17196 18288 17202
rect 18236 17138 18288 17144
rect 18696 17196 18748 17202
rect 18696 17138 18748 17144
rect 19616 17196 19668 17202
rect 19616 17138 19668 17144
rect 20076 17196 20128 17202
rect 20076 17138 20128 17144
rect 21008 16794 21036 19200
rect 21468 17202 21496 19200
rect 22388 17202 22416 19200
rect 22848 17202 22876 19200
rect 23768 17202 23796 19200
rect 21456 17196 21508 17202
rect 21456 17138 21508 17144
rect 22376 17196 22428 17202
rect 22376 17138 22428 17144
rect 22836 17196 22888 17202
rect 22836 17138 22888 17144
rect 23756 17196 23808 17202
rect 23756 17138 23808 17144
rect 22622 16892 22930 16901
rect 22622 16890 22628 16892
rect 22684 16890 22708 16892
rect 22764 16890 22788 16892
rect 22844 16890 22868 16892
rect 22924 16890 22930 16892
rect 22684 16838 22686 16890
rect 22866 16838 22868 16890
rect 22622 16836 22628 16838
rect 22684 16836 22708 16838
rect 22764 16836 22788 16838
rect 22844 16836 22868 16838
rect 22924 16836 22930 16838
rect 22622 16827 22930 16836
rect 24228 16794 24256 19200
rect 25148 17202 25176 19200
rect 25608 17202 25636 19200
rect 26528 17202 26556 19200
rect 25136 17196 25188 17202
rect 25136 17138 25188 17144
rect 25596 17196 25648 17202
rect 25596 17138 25648 17144
rect 26516 17196 26568 17202
rect 26516 17138 26568 17144
rect 26988 16794 27016 19200
rect 27908 17202 27936 19200
rect 28368 17202 28396 19200
rect 29288 17202 29316 19200
rect 29748 17202 29776 19200
rect 29846 17436 30154 17445
rect 29846 17434 29852 17436
rect 29908 17434 29932 17436
rect 29988 17434 30012 17436
rect 30068 17434 30092 17436
rect 30148 17434 30154 17436
rect 29908 17382 29910 17434
rect 30090 17382 30092 17434
rect 29846 17380 29852 17382
rect 29908 17380 29932 17382
rect 29988 17380 30012 17382
rect 30068 17380 30092 17382
rect 30148 17380 30154 17382
rect 29846 17371 30154 17380
rect 30668 17202 30696 19200
rect 31128 17202 31156 19200
rect 32048 17202 32076 19200
rect 32508 17202 32536 19200
rect 33428 17202 33456 19200
rect 33888 17202 33916 19200
rect 34808 17202 34836 19200
rect 27896 17196 27948 17202
rect 27896 17138 27948 17144
rect 28356 17196 28408 17202
rect 28356 17138 28408 17144
rect 29276 17196 29328 17202
rect 29276 17138 29328 17144
rect 29736 17196 29788 17202
rect 29736 17138 29788 17144
rect 30656 17196 30708 17202
rect 30656 17138 30708 17144
rect 31116 17196 31168 17202
rect 31116 17138 31168 17144
rect 32036 17196 32088 17202
rect 32036 17138 32088 17144
rect 32496 17196 32548 17202
rect 32496 17138 32548 17144
rect 33416 17196 33468 17202
rect 33416 17138 33468 17144
rect 33876 17196 33928 17202
rect 33876 17138 33928 17144
rect 34796 17196 34848 17202
rect 34796 17138 34848 17144
rect 35268 17134 35296 19200
rect 35256 17128 35308 17134
rect 35256 17070 35308 17076
rect 36188 16794 36216 19200
rect 36648 17202 36676 19200
rect 37568 17202 37596 19200
rect 38028 17202 38056 19200
rect 38948 17202 38976 19200
rect 36636 17196 36688 17202
rect 36636 17138 36688 17144
rect 37556 17196 37608 17202
rect 37556 17138 37608 17144
rect 38016 17196 38068 17202
rect 38016 17138 38068 17144
rect 38936 17196 38988 17202
rect 38936 17138 38988 17144
rect 37070 16892 37378 16901
rect 37070 16890 37076 16892
rect 37132 16890 37156 16892
rect 37212 16890 37236 16892
rect 37292 16890 37316 16892
rect 37372 16890 37378 16892
rect 37132 16838 37134 16890
rect 37314 16838 37316 16890
rect 37070 16836 37076 16838
rect 37132 16836 37156 16838
rect 37212 16836 37236 16838
rect 37292 16836 37316 16838
rect 37372 16836 37378 16838
rect 37070 16827 37378 16836
rect 39408 16794 39436 19200
rect 40328 17202 40356 19200
rect 40788 17202 40816 19200
rect 41708 17202 41736 19200
rect 40316 17196 40368 17202
rect 40316 17138 40368 17144
rect 40776 17196 40828 17202
rect 40776 17138 40828 17144
rect 41696 17196 41748 17202
rect 41696 17138 41748 17144
rect 42168 17066 42196 19200
rect 43088 17202 43116 19200
rect 43076 17196 43128 17202
rect 43076 17138 43128 17144
rect 42156 17060 42208 17066
rect 42156 17002 42208 17008
rect 43548 16794 43576 19200
rect 44468 17898 44496 19200
rect 44468 17870 44680 17898
rect 44294 17436 44602 17445
rect 44294 17434 44300 17436
rect 44356 17434 44380 17436
rect 44436 17434 44460 17436
rect 44516 17434 44540 17436
rect 44596 17434 44602 17436
rect 44356 17382 44358 17434
rect 44538 17382 44540 17434
rect 44294 17380 44300 17382
rect 44356 17380 44380 17382
rect 44436 17380 44460 17382
rect 44516 17380 44540 17382
rect 44596 17380 44602 17382
rect 44294 17371 44602 17380
rect 44652 17202 44680 17870
rect 44640 17196 44692 17202
rect 44640 17138 44692 17144
rect 44928 17134 44956 19200
rect 45848 17202 45876 19200
rect 45836 17196 45888 17202
rect 45836 17138 45888 17144
rect 44916 17128 44968 17134
rect 44916 17070 44968 17076
rect 46308 16794 46336 19200
rect 47228 17202 47256 19200
rect 47688 17202 47716 19200
rect 48608 17202 48636 19200
rect 47216 17196 47268 17202
rect 47216 17138 47268 17144
rect 47676 17196 47728 17202
rect 47676 17138 47728 17144
rect 48596 17196 48648 17202
rect 48596 17138 48648 17144
rect 49068 16794 49096 19200
rect 49988 17202 50016 19200
rect 50448 17202 50476 19200
rect 51368 17202 51396 19200
rect 51828 17202 51856 19200
rect 49976 17196 50028 17202
rect 49976 17138 50028 17144
rect 50436 17196 50488 17202
rect 50436 17138 50488 17144
rect 51356 17196 51408 17202
rect 51356 17138 51408 17144
rect 51816 17196 51868 17202
rect 51816 17138 51868 17144
rect 52748 17066 52776 19200
rect 53208 17202 53236 19200
rect 53196 17196 53248 17202
rect 53196 17138 53248 17144
rect 52736 17060 52788 17066
rect 52736 17002 52788 17008
rect 51518 16892 51826 16901
rect 51518 16890 51524 16892
rect 51580 16890 51604 16892
rect 51660 16890 51684 16892
rect 51740 16890 51764 16892
rect 51820 16890 51826 16892
rect 51580 16838 51582 16890
rect 51762 16838 51764 16890
rect 51518 16836 51524 16838
rect 51580 16836 51604 16838
rect 51660 16836 51684 16838
rect 51740 16836 51764 16838
rect 51820 16836 51826 16838
rect 51518 16827 51826 16836
rect 54128 16794 54156 19200
rect 54588 17202 54616 19200
rect 55508 17202 55536 19200
rect 55968 17218 55996 19200
rect 55968 17202 56088 17218
rect 54576 17196 54628 17202
rect 54576 17138 54628 17144
rect 55496 17196 55548 17202
rect 55968 17196 56100 17202
rect 55968 17190 56048 17196
rect 55496 17138 55548 17144
rect 56048 17138 56100 17144
rect 6276 16788 6328 16794
rect 6276 16730 6328 16736
rect 11336 16788 11388 16794
rect 11336 16730 11388 16736
rect 14096 16788 14148 16794
rect 14096 16730 14148 16736
rect 16856 16788 16908 16794
rect 16856 16730 16908 16736
rect 20996 16788 21048 16794
rect 20996 16730 21048 16736
rect 24216 16788 24268 16794
rect 24216 16730 24268 16736
rect 26976 16788 27028 16794
rect 26976 16730 27028 16736
rect 36176 16788 36228 16794
rect 36176 16730 36228 16736
rect 39396 16788 39448 16794
rect 39396 16730 39448 16736
rect 43536 16788 43588 16794
rect 43536 16730 43588 16736
rect 46296 16788 46348 16794
rect 46296 16730 46348 16736
rect 49056 16788 49108 16794
rect 49056 16730 49108 16736
rect 54116 16788 54168 16794
rect 54116 16730 54168 16736
rect 15398 16348 15706 16357
rect 15398 16346 15404 16348
rect 15460 16346 15484 16348
rect 15540 16346 15564 16348
rect 15620 16346 15644 16348
rect 15700 16346 15706 16348
rect 15460 16294 15462 16346
rect 15642 16294 15644 16346
rect 15398 16292 15404 16294
rect 15460 16292 15484 16294
rect 15540 16292 15564 16294
rect 15620 16292 15644 16294
rect 15700 16292 15706 16294
rect 15398 16283 15706 16292
rect 29846 16348 30154 16357
rect 29846 16346 29852 16348
rect 29908 16346 29932 16348
rect 29988 16346 30012 16348
rect 30068 16346 30092 16348
rect 30148 16346 30154 16348
rect 29908 16294 29910 16346
rect 30090 16294 30092 16346
rect 29846 16292 29852 16294
rect 29908 16292 29932 16294
rect 29988 16292 30012 16294
rect 30068 16292 30092 16294
rect 30148 16292 30154 16294
rect 29846 16283 30154 16292
rect 44294 16348 44602 16357
rect 44294 16346 44300 16348
rect 44356 16346 44380 16348
rect 44436 16346 44460 16348
rect 44516 16346 44540 16348
rect 44596 16346 44602 16348
rect 44356 16294 44358 16346
rect 44538 16294 44540 16346
rect 44294 16292 44300 16294
rect 44356 16292 44380 16294
rect 44436 16292 44460 16294
rect 44516 16292 44540 16294
rect 44596 16292 44602 16294
rect 44294 16283 44602 16292
rect 8174 15804 8482 15813
rect 8174 15802 8180 15804
rect 8236 15802 8260 15804
rect 8316 15802 8340 15804
rect 8396 15802 8420 15804
rect 8476 15802 8482 15804
rect 8236 15750 8238 15802
rect 8418 15750 8420 15802
rect 8174 15748 8180 15750
rect 8236 15748 8260 15750
rect 8316 15748 8340 15750
rect 8396 15748 8420 15750
rect 8476 15748 8482 15750
rect 8174 15739 8482 15748
rect 22622 15804 22930 15813
rect 22622 15802 22628 15804
rect 22684 15802 22708 15804
rect 22764 15802 22788 15804
rect 22844 15802 22868 15804
rect 22924 15802 22930 15804
rect 22684 15750 22686 15802
rect 22866 15750 22868 15802
rect 22622 15748 22628 15750
rect 22684 15748 22708 15750
rect 22764 15748 22788 15750
rect 22844 15748 22868 15750
rect 22924 15748 22930 15750
rect 22622 15739 22930 15748
rect 37070 15804 37378 15813
rect 37070 15802 37076 15804
rect 37132 15802 37156 15804
rect 37212 15802 37236 15804
rect 37292 15802 37316 15804
rect 37372 15802 37378 15804
rect 37132 15750 37134 15802
rect 37314 15750 37316 15802
rect 37070 15748 37076 15750
rect 37132 15748 37156 15750
rect 37212 15748 37236 15750
rect 37292 15748 37316 15750
rect 37372 15748 37378 15750
rect 37070 15739 37378 15748
rect 51518 15804 51826 15813
rect 51518 15802 51524 15804
rect 51580 15802 51604 15804
rect 51660 15802 51684 15804
rect 51740 15802 51764 15804
rect 51820 15802 51826 15804
rect 51580 15750 51582 15802
rect 51762 15750 51764 15802
rect 51518 15748 51524 15750
rect 51580 15748 51604 15750
rect 51660 15748 51684 15750
rect 51740 15748 51764 15750
rect 51820 15748 51826 15750
rect 51518 15739 51826 15748
rect 15398 15260 15706 15269
rect 15398 15258 15404 15260
rect 15460 15258 15484 15260
rect 15540 15258 15564 15260
rect 15620 15258 15644 15260
rect 15700 15258 15706 15260
rect 15460 15206 15462 15258
rect 15642 15206 15644 15258
rect 15398 15204 15404 15206
rect 15460 15204 15484 15206
rect 15540 15204 15564 15206
rect 15620 15204 15644 15206
rect 15700 15204 15706 15206
rect 15398 15195 15706 15204
rect 29846 15260 30154 15269
rect 29846 15258 29852 15260
rect 29908 15258 29932 15260
rect 29988 15258 30012 15260
rect 30068 15258 30092 15260
rect 30148 15258 30154 15260
rect 29908 15206 29910 15258
rect 30090 15206 30092 15258
rect 29846 15204 29852 15206
rect 29908 15204 29932 15206
rect 29988 15204 30012 15206
rect 30068 15204 30092 15206
rect 30148 15204 30154 15206
rect 29846 15195 30154 15204
rect 44294 15260 44602 15269
rect 44294 15258 44300 15260
rect 44356 15258 44380 15260
rect 44436 15258 44460 15260
rect 44516 15258 44540 15260
rect 44596 15258 44602 15260
rect 44356 15206 44358 15258
rect 44538 15206 44540 15258
rect 44294 15204 44300 15206
rect 44356 15204 44380 15206
rect 44436 15204 44460 15206
rect 44516 15204 44540 15206
rect 44596 15204 44602 15206
rect 44294 15195 44602 15204
rect 8174 14716 8482 14725
rect 8174 14714 8180 14716
rect 8236 14714 8260 14716
rect 8316 14714 8340 14716
rect 8396 14714 8420 14716
rect 8476 14714 8482 14716
rect 8236 14662 8238 14714
rect 8418 14662 8420 14714
rect 8174 14660 8180 14662
rect 8236 14660 8260 14662
rect 8316 14660 8340 14662
rect 8396 14660 8420 14662
rect 8476 14660 8482 14662
rect 8174 14651 8482 14660
rect 22622 14716 22930 14725
rect 22622 14714 22628 14716
rect 22684 14714 22708 14716
rect 22764 14714 22788 14716
rect 22844 14714 22868 14716
rect 22924 14714 22930 14716
rect 22684 14662 22686 14714
rect 22866 14662 22868 14714
rect 22622 14660 22628 14662
rect 22684 14660 22708 14662
rect 22764 14660 22788 14662
rect 22844 14660 22868 14662
rect 22924 14660 22930 14662
rect 22622 14651 22930 14660
rect 37070 14716 37378 14725
rect 37070 14714 37076 14716
rect 37132 14714 37156 14716
rect 37212 14714 37236 14716
rect 37292 14714 37316 14716
rect 37372 14714 37378 14716
rect 37132 14662 37134 14714
rect 37314 14662 37316 14714
rect 37070 14660 37076 14662
rect 37132 14660 37156 14662
rect 37212 14660 37236 14662
rect 37292 14660 37316 14662
rect 37372 14660 37378 14662
rect 37070 14651 37378 14660
rect 51518 14716 51826 14725
rect 51518 14714 51524 14716
rect 51580 14714 51604 14716
rect 51660 14714 51684 14716
rect 51740 14714 51764 14716
rect 51820 14714 51826 14716
rect 51580 14662 51582 14714
rect 51762 14662 51764 14714
rect 51518 14660 51524 14662
rect 51580 14660 51604 14662
rect 51660 14660 51684 14662
rect 51740 14660 51764 14662
rect 51820 14660 51826 14662
rect 51518 14651 51826 14660
rect 15398 14172 15706 14181
rect 15398 14170 15404 14172
rect 15460 14170 15484 14172
rect 15540 14170 15564 14172
rect 15620 14170 15644 14172
rect 15700 14170 15706 14172
rect 15460 14118 15462 14170
rect 15642 14118 15644 14170
rect 15398 14116 15404 14118
rect 15460 14116 15484 14118
rect 15540 14116 15564 14118
rect 15620 14116 15644 14118
rect 15700 14116 15706 14118
rect 15398 14107 15706 14116
rect 29846 14172 30154 14181
rect 29846 14170 29852 14172
rect 29908 14170 29932 14172
rect 29988 14170 30012 14172
rect 30068 14170 30092 14172
rect 30148 14170 30154 14172
rect 29908 14118 29910 14170
rect 30090 14118 30092 14170
rect 29846 14116 29852 14118
rect 29908 14116 29932 14118
rect 29988 14116 30012 14118
rect 30068 14116 30092 14118
rect 30148 14116 30154 14118
rect 29846 14107 30154 14116
rect 44294 14172 44602 14181
rect 44294 14170 44300 14172
rect 44356 14170 44380 14172
rect 44436 14170 44460 14172
rect 44516 14170 44540 14172
rect 44596 14170 44602 14172
rect 44356 14118 44358 14170
rect 44538 14118 44540 14170
rect 44294 14116 44300 14118
rect 44356 14116 44380 14118
rect 44436 14116 44460 14118
rect 44516 14116 44540 14118
rect 44596 14116 44602 14118
rect 44294 14107 44602 14116
rect 20260 13932 20312 13938
rect 20260 13874 20312 13880
rect 3148 13864 3200 13870
rect 13360 13864 13412 13870
rect 3148 13806 3200 13812
rect 13358 13832 13360 13841
rect 13412 13832 13414 13841
rect 1492 13184 1544 13190
rect 1492 13126 1544 13132
rect 2688 13184 2740 13190
rect 2688 13126 2740 13132
rect 1400 8356 1452 8362
rect 1400 8298 1452 8304
rect 1412 3670 1440 8298
rect 1400 3664 1452 3670
rect 1400 3606 1452 3612
rect 1504 3058 1532 13126
rect 1952 12640 2004 12646
rect 1952 12582 2004 12588
rect 1964 12481 1992 12582
rect 1950 12472 2006 12481
rect 1950 12407 2006 12416
rect 1860 12232 1912 12238
rect 1860 12174 1912 12180
rect 1676 12096 1728 12102
rect 1676 12038 1728 12044
rect 1584 11552 1636 11558
rect 1584 11494 1636 11500
rect 1596 10674 1624 11494
rect 1584 10668 1636 10674
rect 1584 10610 1636 10616
rect 1596 10577 1624 10610
rect 1582 10568 1638 10577
rect 1582 10503 1638 10512
rect 1688 10062 1716 12038
rect 1766 11792 1822 11801
rect 1766 11727 1822 11736
rect 1780 10810 1808 11727
rect 1768 10804 1820 10810
rect 1768 10746 1820 10752
rect 1872 10690 1900 12174
rect 2044 11280 2096 11286
rect 2042 11248 2044 11257
rect 2096 11248 2098 11257
rect 2042 11183 2098 11192
rect 2700 11098 2728 13126
rect 3160 12714 3188 13806
rect 13358 13767 13414 13776
rect 8174 13628 8482 13637
rect 8174 13626 8180 13628
rect 8236 13626 8260 13628
rect 8316 13626 8340 13628
rect 8396 13626 8420 13628
rect 8476 13626 8482 13628
rect 8236 13574 8238 13626
rect 8418 13574 8420 13626
rect 8174 13572 8180 13574
rect 8236 13572 8260 13574
rect 8316 13572 8340 13574
rect 8396 13572 8420 13574
rect 8476 13572 8482 13574
rect 8174 13563 8482 13572
rect 11428 13320 11480 13326
rect 11428 13262 11480 13268
rect 15200 13320 15252 13326
rect 15200 13262 15252 13268
rect 5264 13252 5316 13258
rect 5264 13194 5316 13200
rect 9496 13252 9548 13258
rect 9496 13194 9548 13200
rect 3240 13184 3292 13190
rect 3240 13126 3292 13132
rect 3792 13184 3844 13190
rect 3792 13126 3844 13132
rect 4988 13184 5040 13190
rect 4988 13126 5040 13132
rect 3148 12708 3200 12714
rect 3148 12650 3200 12656
rect 3160 12238 3188 12650
rect 3148 12232 3200 12238
rect 3148 12174 3200 12180
rect 2964 12096 3016 12102
rect 2964 12038 3016 12044
rect 2976 11898 3004 12038
rect 2964 11892 3016 11898
rect 2964 11834 3016 11840
rect 2700 11070 2912 11098
rect 2596 11008 2648 11014
rect 2596 10950 2648 10956
rect 2608 10810 2636 10950
rect 2596 10804 2648 10810
rect 2596 10746 2648 10752
rect 1780 10662 1900 10690
rect 2688 10736 2740 10742
rect 2688 10678 2740 10684
rect 1676 10056 1728 10062
rect 1676 9998 1728 10004
rect 1584 8288 1636 8294
rect 1584 8230 1636 8236
rect 1596 7410 1624 8230
rect 1584 7404 1636 7410
rect 1584 7346 1636 7352
rect 1688 6914 1716 9998
rect 1780 9586 1808 10662
rect 2044 10600 2096 10606
rect 2700 10554 2728 10678
rect 2044 10542 2096 10548
rect 1860 9920 1912 9926
rect 1860 9862 1912 9868
rect 1872 9761 1900 9862
rect 1858 9752 1914 9761
rect 1858 9687 1914 9696
rect 1768 9580 1820 9586
rect 1768 9522 1820 9528
rect 1780 8401 1808 9522
rect 1952 8968 2004 8974
rect 1952 8910 2004 8916
rect 1766 8392 1822 8401
rect 1766 8327 1822 8336
rect 1860 8356 1912 8362
rect 1860 8298 1912 8304
rect 1768 8084 1820 8090
rect 1768 8026 1820 8032
rect 1596 6886 1716 6914
rect 1596 4865 1624 6886
rect 1780 6780 1808 8026
rect 1872 7886 1900 8298
rect 1860 7880 1912 7886
rect 1860 7822 1912 7828
rect 1964 6914 1992 8910
rect 2056 8498 2084 10542
rect 2608 10526 2728 10554
rect 2504 9920 2556 9926
rect 2502 9888 2504 9897
rect 2556 9888 2558 9897
rect 2502 9823 2558 9832
rect 2412 9036 2464 9042
rect 2412 8978 2464 8984
rect 2320 8560 2372 8566
rect 2320 8502 2372 8508
rect 2044 8492 2096 8498
rect 2044 8434 2096 8440
rect 2056 8090 2084 8434
rect 2044 8084 2096 8090
rect 2044 8026 2096 8032
rect 2044 7744 2096 7750
rect 2044 7686 2096 7692
rect 2056 7478 2084 7686
rect 2044 7472 2096 7478
rect 2044 7414 2096 7420
rect 2228 7200 2280 7206
rect 2228 7142 2280 7148
rect 1964 6886 2084 6914
rect 1688 6752 1808 6780
rect 1582 4856 1638 4865
rect 1582 4791 1638 4800
rect 1492 3052 1544 3058
rect 1492 2994 1544 3000
rect 1688 2378 1716 6752
rect 1860 6724 1912 6730
rect 1860 6666 1912 6672
rect 1872 5914 1900 6666
rect 1952 6112 2004 6118
rect 1952 6054 2004 6060
rect 1860 5908 1912 5914
rect 1860 5850 1912 5856
rect 1964 5302 1992 6054
rect 1952 5296 2004 5302
rect 1952 5238 2004 5244
rect 1860 4548 1912 4554
rect 1860 4490 1912 4496
rect 1766 4312 1822 4321
rect 1766 4247 1822 4256
rect 1780 4146 1808 4247
rect 1872 4185 1900 4490
rect 1858 4176 1914 4185
rect 1768 4140 1820 4146
rect 2056 4162 2084 6886
rect 2136 6792 2188 6798
rect 2136 6734 2188 6740
rect 2148 6458 2176 6734
rect 2136 6452 2188 6458
rect 2136 6394 2188 6400
rect 2136 6316 2188 6322
rect 2136 6258 2188 6264
rect 2148 5522 2176 6258
rect 2240 5710 2268 7142
rect 2228 5704 2280 5710
rect 2228 5646 2280 5652
rect 2148 5494 2268 5522
rect 2136 5228 2188 5234
rect 2136 5170 2188 5176
rect 2148 5137 2176 5170
rect 2134 5128 2190 5137
rect 2134 5063 2190 5072
rect 2136 4548 2188 4554
rect 2240 4536 2268 5494
rect 2188 4508 2268 4536
rect 2136 4490 2188 4496
rect 2148 4282 2176 4490
rect 2136 4276 2188 4282
rect 2136 4218 2188 4224
rect 1858 4111 1914 4120
rect 1964 4134 2084 4162
rect 1768 4082 1820 4088
rect 1780 3194 1808 4082
rect 1768 3188 1820 3194
rect 1768 3130 1820 3136
rect 1964 3126 1992 4134
rect 2044 4072 2096 4078
rect 2044 4014 2096 4020
rect 2056 3738 2084 4014
rect 2136 3936 2188 3942
rect 2136 3878 2188 3884
rect 2044 3732 2096 3738
rect 2044 3674 2096 3680
rect 1952 3120 2004 3126
rect 1952 3062 2004 3068
rect 1964 2650 1992 3062
rect 1952 2644 2004 2650
rect 1952 2586 2004 2592
rect 1676 2372 1728 2378
rect 1676 2314 1728 2320
rect 2148 2038 2176 3878
rect 2226 2680 2282 2689
rect 2226 2615 2282 2624
rect 2240 2514 2268 2615
rect 2332 2514 2360 8502
rect 2424 3738 2452 8978
rect 2608 8566 2636 10526
rect 2688 10464 2740 10470
rect 2688 10406 2740 10412
rect 2596 8560 2648 8566
rect 2596 8502 2648 8508
rect 2504 7744 2556 7750
rect 2504 7686 2556 7692
rect 2516 6322 2544 7686
rect 2596 6656 2648 6662
rect 2596 6598 2648 6604
rect 2608 6497 2636 6598
rect 2594 6488 2650 6497
rect 2594 6423 2650 6432
rect 2504 6316 2556 6322
rect 2504 6258 2556 6264
rect 2700 5658 2728 10406
rect 2780 9512 2832 9518
rect 2780 9454 2832 9460
rect 2792 8430 2820 9454
rect 2780 8424 2832 8430
rect 2780 8366 2832 8372
rect 2608 5630 2728 5658
rect 2780 5704 2832 5710
rect 2780 5646 2832 5652
rect 2502 4720 2558 4729
rect 2502 4655 2558 4664
rect 2516 4622 2544 4655
rect 2504 4616 2556 4622
rect 2504 4558 2556 4564
rect 2412 3732 2464 3738
rect 2412 3674 2464 3680
rect 2424 3602 2452 3674
rect 2412 3596 2464 3602
rect 2412 3538 2464 3544
rect 2228 2508 2280 2514
rect 2228 2450 2280 2456
rect 2320 2508 2372 2514
rect 2320 2450 2372 2456
rect 2608 2310 2636 5630
rect 2686 5400 2742 5409
rect 2686 5335 2742 5344
rect 2700 4146 2728 5335
rect 2792 5302 2820 5646
rect 2780 5296 2832 5302
rect 2780 5238 2832 5244
rect 2688 4140 2740 4146
rect 2688 4082 2740 4088
rect 2780 3664 2832 3670
rect 2780 3606 2832 3612
rect 2792 2922 2820 3606
rect 2884 3534 2912 11070
rect 2976 10146 3004 11834
rect 2976 10118 3188 10146
rect 2964 10056 3016 10062
rect 2964 9998 3016 10004
rect 2976 9722 3004 9998
rect 2964 9716 3016 9722
rect 2964 9658 3016 9664
rect 3160 9654 3188 10118
rect 3148 9648 3200 9654
rect 3148 9590 3200 9596
rect 3056 9580 3108 9586
rect 3056 9522 3108 9528
rect 2964 9036 3016 9042
rect 2964 8978 3016 8984
rect 2976 7954 3004 8978
rect 3068 8974 3096 9522
rect 3056 8968 3108 8974
rect 3056 8910 3108 8916
rect 2964 7948 3016 7954
rect 2964 7890 3016 7896
rect 2976 7274 3004 7890
rect 3146 7304 3202 7313
rect 2964 7268 3016 7274
rect 3146 7239 3202 7248
rect 2964 7210 3016 7216
rect 3056 7200 3108 7206
rect 3056 7142 3108 7148
rect 2964 6112 3016 6118
rect 2964 6054 3016 6060
rect 2976 4622 3004 6054
rect 3068 5778 3096 7142
rect 3160 6798 3188 7239
rect 3148 6792 3200 6798
rect 3148 6734 3200 6740
rect 3148 6656 3200 6662
rect 3148 6598 3200 6604
rect 3056 5772 3108 5778
rect 3056 5714 3108 5720
rect 3054 5672 3110 5681
rect 3054 5607 3056 5616
rect 3108 5607 3110 5616
rect 3056 5578 3108 5584
rect 3160 5302 3188 6598
rect 3148 5296 3200 5302
rect 3148 5238 3200 5244
rect 2964 4616 3016 4622
rect 2964 4558 3016 4564
rect 3252 4146 3280 13126
rect 3608 12640 3660 12646
rect 3608 12582 3660 12588
rect 3332 12232 3384 12238
rect 3332 12174 3384 12180
rect 3344 8838 3372 12174
rect 3620 11626 3648 12582
rect 3804 12481 3832 13126
rect 3976 12912 4028 12918
rect 3976 12854 4028 12860
rect 3790 12472 3846 12481
rect 3790 12407 3846 12416
rect 3884 12096 3936 12102
rect 3884 12038 3936 12044
rect 3424 11620 3476 11626
rect 3424 11562 3476 11568
rect 3608 11620 3660 11626
rect 3608 11562 3660 11568
rect 3436 9042 3464 11562
rect 3896 11354 3924 12038
rect 3884 11348 3936 11354
rect 3884 11290 3936 11296
rect 3608 11212 3660 11218
rect 3608 11154 3660 11160
rect 3516 9580 3568 9586
rect 3516 9522 3568 9528
rect 3528 9178 3556 9522
rect 3516 9172 3568 9178
rect 3516 9114 3568 9120
rect 3424 9036 3476 9042
rect 3424 8978 3476 8984
rect 3332 8832 3384 8838
rect 3332 8774 3384 8780
rect 2964 4140 3016 4146
rect 2964 4082 3016 4088
rect 3240 4140 3292 4146
rect 3240 4082 3292 4088
rect 2976 3670 3004 4082
rect 3252 4026 3280 4082
rect 3160 3998 3280 4026
rect 2964 3664 3016 3670
rect 2964 3606 3016 3612
rect 2872 3528 2924 3534
rect 2872 3470 2924 3476
rect 2780 2916 2832 2922
rect 2780 2858 2832 2864
rect 2884 2774 2912 3470
rect 2964 3052 3016 3058
rect 2964 2994 3016 3000
rect 2792 2746 2912 2774
rect 2596 2304 2648 2310
rect 2596 2246 2648 2252
rect 2136 2032 2188 2038
rect 2136 1974 2188 1980
rect 2792 1902 2820 2746
rect 2976 2650 3004 2994
rect 2964 2644 3016 2650
rect 2964 2586 3016 2592
rect 2780 1896 2832 1902
rect 2780 1838 2832 1844
rect 3160 1698 3188 3998
rect 3344 3058 3372 8774
rect 3516 8492 3568 8498
rect 3516 8434 3568 8440
rect 3424 8424 3476 8430
rect 3424 8366 3476 8372
rect 3436 7410 3464 8366
rect 3528 8090 3556 8434
rect 3516 8084 3568 8090
rect 3516 8026 3568 8032
rect 3528 7886 3556 8026
rect 3516 7880 3568 7886
rect 3516 7822 3568 7828
rect 3424 7404 3476 7410
rect 3424 7346 3476 7352
rect 3516 6792 3568 6798
rect 3516 6734 3568 6740
rect 3422 5808 3478 5817
rect 3422 5743 3478 5752
rect 3436 5710 3464 5743
rect 3424 5704 3476 5710
rect 3424 5646 3476 5652
rect 3332 3052 3384 3058
rect 3332 2994 3384 3000
rect 3240 2848 3292 2854
rect 3240 2790 3292 2796
rect 3148 1692 3200 1698
rect 3148 1634 3200 1640
rect 3252 814 3280 2790
rect 3528 1834 3556 6734
rect 3620 2582 3648 11154
rect 3792 11008 3844 11014
rect 3792 10950 3844 10956
rect 3804 10810 3832 10950
rect 3988 10810 4016 12854
rect 5000 12434 5028 13126
rect 5276 12646 5304 13194
rect 6276 13184 6328 13190
rect 6276 13126 6328 13132
rect 5908 12844 5960 12850
rect 5908 12786 5960 12792
rect 5264 12640 5316 12646
rect 5264 12582 5316 12588
rect 4632 12406 5028 12434
rect 4252 11824 4304 11830
rect 4252 11766 4304 11772
rect 4160 11076 4212 11082
rect 4160 11018 4212 11024
rect 3792 10804 3844 10810
rect 3792 10746 3844 10752
rect 3976 10804 4028 10810
rect 3976 10746 4028 10752
rect 4172 10674 4200 11018
rect 4160 10668 4212 10674
rect 4160 10610 4212 10616
rect 3792 10464 3844 10470
rect 3792 10406 3844 10412
rect 3804 8974 3832 10406
rect 4068 10260 4120 10266
rect 4068 10202 4120 10208
rect 4080 9654 4108 10202
rect 4172 10169 4200 10610
rect 4158 10160 4214 10169
rect 4158 10095 4214 10104
rect 4068 9648 4120 9654
rect 4068 9590 4120 9596
rect 3884 9580 3936 9586
rect 3884 9522 3936 9528
rect 3896 9110 3924 9522
rect 3884 9104 3936 9110
rect 3884 9046 3936 9052
rect 4080 9042 4108 9590
rect 4264 9178 4292 11766
rect 4344 11552 4396 11558
rect 4344 11494 4396 11500
rect 4252 9172 4304 9178
rect 4252 9114 4304 9120
rect 4068 9036 4120 9042
rect 4068 8978 4120 8984
rect 3792 8968 3844 8974
rect 3792 8910 3844 8916
rect 3698 7032 3754 7041
rect 3698 6967 3754 6976
rect 3712 6866 3740 6967
rect 3700 6860 3752 6866
rect 3700 6802 3752 6808
rect 3698 6352 3754 6361
rect 3698 6287 3754 6296
rect 3712 5710 3740 6287
rect 3700 5704 3752 5710
rect 3700 5646 3752 5652
rect 3804 4321 3832 8910
rect 4356 8498 4384 11494
rect 4436 11144 4488 11150
rect 4436 11086 4488 11092
rect 4448 9994 4476 11086
rect 4436 9988 4488 9994
rect 4436 9930 4488 9936
rect 4344 8492 4396 8498
rect 4344 8434 4396 8440
rect 4252 8356 4304 8362
rect 4252 8298 4304 8304
rect 4264 7546 4292 8298
rect 4344 7880 4396 7886
rect 4344 7822 4396 7828
rect 4356 7546 4384 7822
rect 4252 7540 4304 7546
rect 4252 7482 4304 7488
rect 4344 7540 4396 7546
rect 4344 7482 4396 7488
rect 4158 7440 4214 7449
rect 4158 7375 4214 7384
rect 4172 7342 4200 7375
rect 4160 7336 4212 7342
rect 4160 7278 4212 7284
rect 4160 7200 4212 7206
rect 4160 7142 4212 7148
rect 3976 6792 4028 6798
rect 3976 6734 4028 6740
rect 3988 6322 4016 6734
rect 3884 6316 3936 6322
rect 3884 6258 3936 6264
rect 3976 6316 4028 6322
rect 3976 6258 4028 6264
rect 3896 5914 3924 6258
rect 3884 5908 3936 5914
rect 3884 5850 3936 5856
rect 4172 5710 4200 7142
rect 4250 6352 4306 6361
rect 4250 6287 4252 6296
rect 4304 6287 4306 6296
rect 4252 6258 4304 6264
rect 4344 6248 4396 6254
rect 4342 6216 4344 6225
rect 4396 6216 4398 6225
rect 4252 6180 4304 6186
rect 4342 6151 4398 6160
rect 4252 6122 4304 6128
rect 4264 5846 4292 6122
rect 4252 5840 4304 5846
rect 4252 5782 4304 5788
rect 3976 5704 4028 5710
rect 3976 5646 4028 5652
rect 4160 5704 4212 5710
rect 4160 5646 4212 5652
rect 3988 5370 4016 5646
rect 4068 5568 4120 5574
rect 4068 5510 4120 5516
rect 3976 5364 4028 5370
rect 3976 5306 4028 5312
rect 4080 4690 4108 5510
rect 4252 5228 4304 5234
rect 4252 5170 4304 5176
rect 4068 4684 4120 4690
rect 4068 4626 4120 4632
rect 4264 4622 4292 5170
rect 4252 4616 4304 4622
rect 4252 4558 4304 4564
rect 3790 4312 3846 4321
rect 3790 4247 3846 4256
rect 4264 3738 4292 4558
rect 4448 4434 4476 9930
rect 4528 9512 4580 9518
rect 4528 9454 4580 9460
rect 4540 8906 4568 9454
rect 4528 8900 4580 8906
rect 4528 8842 4580 8848
rect 4540 8498 4568 8842
rect 4528 8492 4580 8498
rect 4528 8434 4580 8440
rect 4632 6882 4660 12406
rect 5172 12096 5224 12102
rect 5172 12038 5224 12044
rect 4896 11552 4948 11558
rect 4896 11494 4948 11500
rect 4908 11082 4936 11494
rect 4988 11144 5040 11150
rect 4988 11086 5040 11092
rect 4896 11076 4948 11082
rect 4896 11018 4948 11024
rect 4712 10668 4764 10674
rect 4712 10610 4764 10616
rect 4724 8634 4752 10610
rect 4896 10464 4948 10470
rect 4896 10406 4948 10412
rect 4804 9920 4856 9926
rect 4804 9862 4856 9868
rect 4816 9722 4844 9862
rect 4804 9716 4856 9722
rect 4804 9658 4856 9664
rect 4908 8974 4936 10406
rect 5000 9602 5028 11086
rect 5092 9625 5120 9685
rect 5078 9616 5134 9625
rect 5000 9574 5078 9602
rect 4896 8968 4948 8974
rect 4896 8910 4948 8916
rect 5000 8786 5028 9574
rect 5078 9551 5080 9560
rect 5132 9551 5134 9560
rect 5080 9522 5132 9528
rect 5080 9444 5132 9450
rect 5080 9386 5132 9392
rect 4816 8758 5028 8786
rect 4712 8628 4764 8634
rect 4712 8570 4764 8576
rect 4712 7744 4764 7750
rect 4712 7686 4764 7692
rect 4724 6934 4752 7686
rect 4540 6854 4660 6882
rect 4712 6928 4764 6934
rect 4712 6870 4764 6876
rect 4816 6882 4844 8758
rect 4988 8560 5040 8566
rect 4988 8502 5040 8508
rect 5000 7886 5028 8502
rect 4988 7880 5040 7886
rect 4988 7822 5040 7828
rect 4816 6854 5028 6882
rect 4540 5658 4568 6854
rect 4712 6656 4764 6662
rect 4712 6598 4764 6604
rect 4724 6118 4752 6598
rect 4804 6180 4856 6186
rect 4804 6122 4856 6128
rect 4712 6112 4764 6118
rect 4712 6054 4764 6060
rect 4724 5914 4752 6054
rect 4712 5908 4764 5914
rect 4712 5850 4764 5856
rect 4540 5630 4660 5658
rect 4528 5568 4580 5574
rect 4528 5510 4580 5516
rect 4540 5234 4568 5510
rect 4528 5228 4580 5234
rect 4528 5170 4580 5176
rect 4448 4406 4568 4434
rect 4436 4276 4488 4282
rect 4436 4218 4488 4224
rect 4344 4140 4396 4146
rect 4344 4082 4396 4088
rect 4252 3732 4304 3738
rect 4252 3674 4304 3680
rect 4252 3528 4304 3534
rect 4250 3496 4252 3505
rect 4304 3496 4306 3505
rect 3792 3460 3844 3466
rect 4250 3431 4306 3440
rect 3792 3402 3844 3408
rect 3804 3194 3832 3402
rect 3792 3188 3844 3194
rect 3792 3130 3844 3136
rect 3884 3052 3936 3058
rect 3884 2994 3936 3000
rect 3608 2576 3660 2582
rect 3608 2518 3660 2524
rect 3516 1828 3568 1834
rect 3516 1770 3568 1776
rect 3896 1737 3924 2994
rect 4356 2650 4384 4082
rect 4448 3058 4476 4218
rect 4436 3052 4488 3058
rect 4436 2994 4488 3000
rect 4344 2644 4396 2650
rect 4344 2586 4396 2592
rect 3976 2440 4028 2446
rect 3976 2382 4028 2388
rect 3988 2009 4016 2382
rect 3974 2000 4030 2009
rect 3974 1935 4030 1944
rect 3882 1728 3938 1737
rect 3882 1663 3938 1672
rect 4540 1018 4568 4406
rect 4632 3058 4660 5630
rect 4816 5030 4844 6122
rect 4804 5024 4856 5030
rect 4804 4966 4856 4972
rect 5000 4842 5028 6854
rect 4724 4814 5028 4842
rect 4724 3602 4752 4814
rect 4894 4448 4950 4457
rect 4894 4383 4950 4392
rect 4908 4146 4936 4383
rect 4896 4140 4948 4146
rect 4896 4082 4948 4088
rect 5092 4026 5120 9386
rect 5184 6322 5212 12038
rect 5172 6316 5224 6322
rect 5172 6258 5224 6264
rect 5184 5642 5212 6258
rect 5172 5636 5224 5642
rect 5172 5578 5224 5584
rect 5172 4548 5224 4554
rect 5172 4490 5224 4496
rect 5184 4146 5212 4490
rect 5172 4140 5224 4146
rect 5172 4082 5224 4088
rect 5276 4078 5304 12582
rect 5920 12170 5948 12786
rect 6288 12434 6316 13126
rect 9508 12986 9536 13194
rect 9588 13184 9640 13190
rect 9588 13126 9640 13132
rect 9680 13184 9732 13190
rect 9680 13126 9732 13132
rect 11060 13184 11112 13190
rect 11060 13126 11112 13132
rect 9496 12980 9548 12986
rect 9496 12922 9548 12928
rect 9220 12708 9272 12714
rect 9220 12650 9272 12656
rect 6552 12640 6604 12646
rect 6552 12582 6604 12588
rect 7012 12640 7064 12646
rect 7012 12582 7064 12588
rect 7932 12640 7984 12646
rect 7932 12582 7984 12588
rect 8852 12640 8904 12646
rect 8852 12582 8904 12588
rect 6564 12442 6592 12582
rect 7024 12481 7052 12582
rect 7010 12472 7066 12481
rect 6552 12436 6604 12442
rect 6288 12406 6500 12434
rect 5908 12164 5960 12170
rect 5908 12106 5960 12112
rect 5816 11552 5868 11558
rect 5814 11520 5816 11529
rect 5868 11520 5870 11529
rect 5814 11455 5870 11464
rect 5920 11286 5948 12106
rect 5908 11280 5960 11286
rect 5908 11222 5960 11228
rect 6368 11280 6420 11286
rect 6368 11222 6420 11228
rect 5816 11076 5868 11082
rect 5816 11018 5868 11024
rect 5828 10810 5856 11018
rect 5816 10804 5868 10810
rect 5816 10746 5868 10752
rect 5632 10056 5684 10062
rect 5632 9998 5684 10004
rect 5644 9722 5672 9998
rect 5632 9716 5684 9722
rect 5632 9658 5684 9664
rect 5632 9376 5684 9382
rect 5632 9318 5684 9324
rect 5448 8424 5500 8430
rect 5448 8366 5500 8372
rect 5356 7744 5408 7750
rect 5356 7686 5408 7692
rect 5368 7206 5396 7686
rect 5460 7478 5488 8366
rect 5540 8016 5592 8022
rect 5540 7958 5592 7964
rect 5448 7472 5500 7478
rect 5448 7414 5500 7420
rect 5448 7268 5500 7274
rect 5448 7210 5500 7216
rect 5356 7200 5408 7206
rect 5356 7142 5408 7148
rect 5356 6928 5408 6934
rect 5356 6870 5408 6876
rect 5368 6798 5396 6870
rect 5356 6792 5408 6798
rect 5356 6734 5408 6740
rect 5460 6458 5488 7210
rect 5448 6452 5500 6458
rect 5448 6394 5500 6400
rect 5552 6322 5580 7958
rect 5540 6316 5592 6322
rect 5540 6258 5592 6264
rect 5356 6248 5408 6254
rect 5354 6216 5356 6225
rect 5408 6216 5410 6225
rect 5354 6151 5410 6160
rect 5540 6180 5592 6186
rect 5540 6122 5592 6128
rect 5448 6112 5500 6118
rect 5448 6054 5500 6060
rect 5356 5704 5408 5710
rect 5460 5658 5488 6054
rect 5552 5710 5580 6122
rect 5408 5652 5488 5658
rect 5356 5646 5488 5652
rect 5540 5704 5592 5710
rect 5540 5646 5592 5652
rect 5368 5630 5488 5646
rect 5460 5302 5488 5630
rect 5448 5296 5500 5302
rect 5448 5238 5500 5244
rect 5460 5166 5488 5238
rect 5448 5160 5500 5166
rect 5448 5102 5500 5108
rect 5460 4622 5488 5102
rect 5448 4616 5500 4622
rect 5448 4558 5500 4564
rect 5540 4480 5592 4486
rect 5540 4422 5592 4428
rect 5264 4072 5316 4078
rect 5092 3998 5212 4026
rect 5264 4014 5316 4020
rect 4804 3936 4856 3942
rect 4804 3878 4856 3884
rect 4896 3936 4948 3942
rect 4896 3878 4948 3884
rect 4816 3738 4844 3878
rect 4804 3732 4856 3738
rect 4804 3674 4856 3680
rect 4712 3596 4764 3602
rect 4712 3538 4764 3544
rect 4620 3052 4672 3058
rect 4620 2994 4672 3000
rect 4632 2961 4660 2994
rect 4618 2952 4674 2961
rect 4618 2887 4674 2896
rect 4908 1086 4936 3878
rect 5078 3088 5134 3097
rect 5078 3023 5080 3032
rect 5132 3023 5134 3032
rect 5080 2994 5132 3000
rect 5184 1766 5212 3998
rect 5276 3602 5304 4014
rect 5264 3596 5316 3602
rect 5264 3538 5316 3544
rect 5276 2446 5304 3538
rect 5552 3534 5580 4422
rect 5540 3528 5592 3534
rect 5540 3470 5592 3476
rect 5448 3392 5500 3398
rect 5446 3360 5448 3369
rect 5500 3360 5502 3369
rect 5446 3295 5502 3304
rect 5644 2774 5672 9318
rect 6092 8968 6144 8974
rect 6092 8910 6144 8916
rect 6104 8673 6132 8910
rect 6090 8664 6146 8673
rect 6090 8599 6146 8608
rect 5816 8492 5868 8498
rect 5816 8434 5868 8440
rect 5828 8378 5856 8434
rect 6090 8392 6146 8401
rect 5828 8350 6040 8378
rect 5724 8288 5776 8294
rect 5724 8230 5776 8236
rect 5816 8288 5868 8294
rect 5816 8230 5868 8236
rect 5736 6254 5764 8230
rect 5828 7886 5856 8230
rect 5816 7880 5868 7886
rect 5816 7822 5868 7828
rect 5908 7880 5960 7886
rect 5908 7822 5960 7828
rect 5828 7342 5856 7822
rect 5816 7336 5868 7342
rect 5816 7278 5868 7284
rect 5828 7002 5856 7278
rect 5816 6996 5868 7002
rect 5816 6938 5868 6944
rect 5920 6390 5948 7822
rect 6012 7721 6040 8350
rect 6090 8327 6146 8336
rect 5998 7712 6054 7721
rect 5998 7647 6054 7656
rect 6000 7336 6052 7342
rect 6000 7278 6052 7284
rect 6012 7041 6040 7278
rect 5998 7032 6054 7041
rect 5998 6967 6054 6976
rect 6000 6656 6052 6662
rect 6000 6598 6052 6604
rect 5908 6384 5960 6390
rect 5908 6326 5960 6332
rect 5724 6248 5776 6254
rect 5724 6190 5776 6196
rect 5814 6216 5870 6225
rect 5814 6151 5870 6160
rect 5828 5137 5856 6151
rect 5908 5636 5960 5642
rect 5908 5578 5960 5584
rect 5814 5128 5870 5137
rect 5814 5063 5816 5072
rect 5868 5063 5870 5072
rect 5816 5034 5868 5040
rect 5828 5003 5856 5034
rect 5722 4992 5778 5001
rect 5722 4927 5778 4936
rect 5736 4729 5764 4927
rect 5722 4720 5778 4729
rect 5722 4655 5778 4664
rect 5814 4040 5870 4049
rect 5814 3975 5816 3984
rect 5868 3975 5870 3984
rect 5816 3946 5868 3952
rect 5816 3188 5868 3194
rect 5816 3130 5868 3136
rect 5552 2746 5672 2774
rect 5264 2440 5316 2446
rect 5264 2382 5316 2388
rect 5552 2378 5580 2746
rect 5828 2650 5856 3130
rect 5816 2644 5868 2650
rect 5816 2586 5868 2592
rect 5540 2372 5592 2378
rect 5540 2314 5592 2320
rect 5172 1760 5224 1766
rect 5172 1702 5224 1708
rect 5920 1154 5948 5578
rect 6012 5030 6040 6598
rect 6000 5024 6052 5030
rect 6000 4966 6052 4972
rect 6104 1222 6132 8327
rect 6184 8084 6236 8090
rect 6184 8026 6236 8032
rect 6196 7002 6224 8026
rect 6274 7576 6330 7585
rect 6274 7511 6330 7520
rect 6288 7410 6316 7511
rect 6380 7449 6408 11222
rect 6472 9738 6500 12406
rect 7944 12434 7972 12582
rect 8174 12540 8482 12549
rect 8174 12538 8180 12540
rect 8236 12538 8260 12540
rect 8316 12538 8340 12540
rect 8396 12538 8420 12540
rect 8476 12538 8482 12540
rect 8236 12486 8238 12538
rect 8418 12486 8420 12538
rect 8174 12484 8180 12486
rect 8236 12484 8260 12486
rect 8316 12484 8340 12486
rect 8396 12484 8420 12486
rect 8476 12484 8482 12486
rect 8174 12475 8482 12484
rect 7010 12407 7066 12416
rect 6552 12378 6604 12384
rect 7208 12406 7972 12434
rect 6920 12164 6972 12170
rect 6920 12106 6972 12112
rect 6932 11898 6960 12106
rect 6920 11892 6972 11898
rect 6920 11834 6972 11840
rect 6932 10554 6960 11834
rect 7104 11144 7156 11150
rect 7104 11086 7156 11092
rect 6840 10526 6960 10554
rect 7012 10600 7064 10606
rect 7012 10542 7064 10548
rect 6472 9710 6592 9738
rect 6460 9580 6512 9586
rect 6460 9522 6512 9528
rect 6472 8634 6500 9522
rect 6460 8628 6512 8634
rect 6460 8570 6512 8576
rect 6564 8514 6592 9710
rect 6840 9518 6868 10526
rect 6920 10464 6972 10470
rect 6920 10406 6972 10412
rect 6932 10266 6960 10406
rect 6920 10260 6972 10266
rect 6920 10202 6972 10208
rect 6828 9512 6880 9518
rect 6828 9454 6880 9460
rect 6736 9376 6788 9382
rect 6736 9318 6788 9324
rect 6748 8974 6776 9318
rect 6736 8968 6788 8974
rect 6736 8910 6788 8916
rect 6472 8486 6592 8514
rect 6366 7440 6422 7449
rect 6276 7404 6328 7410
rect 6366 7375 6368 7384
rect 6276 7346 6328 7352
rect 6420 7375 6422 7384
rect 6368 7346 6420 7352
rect 6380 7315 6408 7346
rect 6472 7154 6500 8486
rect 6550 8392 6606 8401
rect 6550 8327 6606 8336
rect 6288 7126 6500 7154
rect 6184 6996 6236 7002
rect 6184 6938 6236 6944
rect 6182 5400 6238 5409
rect 6182 5335 6238 5344
rect 6196 4758 6224 5335
rect 6184 4752 6236 4758
rect 6182 4720 6184 4729
rect 6236 4720 6238 4729
rect 6182 4655 6238 4664
rect 6288 4593 6316 7126
rect 6458 7032 6514 7041
rect 6458 6967 6514 6976
rect 6366 5808 6422 5817
rect 6366 5743 6368 5752
rect 6420 5743 6422 5752
rect 6368 5714 6420 5720
rect 6274 4584 6330 4593
rect 6274 4519 6330 4528
rect 6288 4214 6316 4519
rect 6368 4480 6420 4486
rect 6368 4422 6420 4428
rect 6380 4282 6408 4422
rect 6368 4276 6420 4282
rect 6368 4218 6420 4224
rect 6276 4208 6328 4214
rect 6276 4150 6328 4156
rect 6472 3194 6500 6967
rect 6564 6798 6592 8327
rect 6642 7848 6698 7857
rect 6642 7783 6698 7792
rect 6656 7585 6684 7783
rect 6642 7576 6698 7585
rect 6642 7511 6698 7520
rect 6734 7440 6790 7449
rect 6840 7426 6868 9454
rect 6840 7398 6960 7426
rect 6734 7375 6790 7384
rect 6748 7206 6776 7375
rect 6932 7206 6960 7398
rect 6736 7200 6788 7206
rect 6736 7142 6788 7148
rect 6920 7200 6972 7206
rect 6920 7142 6972 7148
rect 6552 6792 6604 6798
rect 6552 6734 6604 6740
rect 6736 6792 6788 6798
rect 6736 6734 6788 6740
rect 6550 6624 6606 6633
rect 6550 6559 6606 6568
rect 6564 4185 6592 6559
rect 6748 6390 6776 6734
rect 6736 6384 6788 6390
rect 6734 6352 6736 6361
rect 6788 6352 6790 6361
rect 6734 6287 6790 6296
rect 6748 6261 6776 6287
rect 6736 6112 6788 6118
rect 6736 6054 6788 6060
rect 6644 5840 6696 5846
rect 6644 5782 6696 5788
rect 6656 5681 6684 5782
rect 6642 5672 6698 5681
rect 6642 5607 6698 5616
rect 6550 4176 6606 4185
rect 6550 4111 6606 4120
rect 6644 4140 6696 4146
rect 6564 3670 6592 4111
rect 6644 4082 6696 4088
rect 6656 3913 6684 4082
rect 6642 3904 6698 3913
rect 6642 3839 6698 3848
rect 6552 3664 6604 3670
rect 6552 3606 6604 3612
rect 6460 3188 6512 3194
rect 6460 3130 6512 3136
rect 6552 2576 6604 2582
rect 6656 2553 6684 3839
rect 6748 2774 6776 6054
rect 6828 5160 6880 5166
rect 6828 5102 6880 5108
rect 6840 4690 6868 5102
rect 6918 4856 6974 4865
rect 6918 4791 6974 4800
rect 6828 4684 6880 4690
rect 6828 4626 6880 4632
rect 6826 3632 6882 3641
rect 6826 3567 6882 3576
rect 6840 3058 6868 3567
rect 6932 3534 6960 4791
rect 7024 3890 7052 10542
rect 7116 4214 7144 11086
rect 7104 4208 7156 4214
rect 7104 4150 7156 4156
rect 7024 3862 7144 3890
rect 7012 3732 7064 3738
rect 7012 3674 7064 3680
rect 6920 3528 6972 3534
rect 6920 3470 6972 3476
rect 6828 3052 6880 3058
rect 6828 2994 6880 3000
rect 6748 2746 6868 2774
rect 6736 2644 6788 2650
rect 6736 2586 6788 2592
rect 6552 2518 6604 2524
rect 6642 2544 6698 2553
rect 6564 1970 6592 2518
rect 6642 2479 6698 2488
rect 6748 2310 6776 2586
rect 6736 2304 6788 2310
rect 6736 2246 6788 2252
rect 6552 1964 6604 1970
rect 6552 1906 6604 1912
rect 6840 1873 6868 2746
rect 6920 2576 6972 2582
rect 6920 2518 6972 2524
rect 6932 2106 6960 2518
rect 6920 2100 6972 2106
rect 6920 2042 6972 2048
rect 6826 1864 6882 1873
rect 6826 1799 6882 1808
rect 7024 1426 7052 3674
rect 7116 3602 7144 3862
rect 7104 3596 7156 3602
rect 7104 3538 7156 3544
rect 7104 3188 7156 3194
rect 7104 3130 7156 3136
rect 7116 2514 7144 3130
rect 7104 2508 7156 2514
rect 7104 2450 7156 2456
rect 7116 1766 7144 2450
rect 7208 2446 7236 12406
rect 8576 12232 8628 12238
rect 8576 12174 8628 12180
rect 7840 12096 7892 12102
rect 7840 12038 7892 12044
rect 7472 11552 7524 11558
rect 7472 11494 7524 11500
rect 7656 11552 7708 11558
rect 7656 11494 7708 11500
rect 7484 11150 7512 11494
rect 7472 11144 7524 11150
rect 7472 11086 7524 11092
rect 7380 10668 7432 10674
rect 7380 10610 7432 10616
rect 7288 9648 7340 9654
rect 7288 9590 7340 9596
rect 7300 6798 7328 9590
rect 7392 9450 7420 10610
rect 7380 9444 7432 9450
rect 7380 9386 7432 9392
rect 7392 9042 7420 9386
rect 7380 9036 7432 9042
rect 7380 8978 7432 8984
rect 7380 8288 7432 8294
rect 7380 8230 7432 8236
rect 7392 7750 7420 8230
rect 7380 7744 7432 7750
rect 7380 7686 7432 7692
rect 7380 7404 7432 7410
rect 7380 7346 7432 7352
rect 7392 7002 7420 7346
rect 7380 6996 7432 7002
rect 7380 6938 7432 6944
rect 7288 6792 7340 6798
rect 7288 6734 7340 6740
rect 7380 6656 7432 6662
rect 7380 6598 7432 6604
rect 7286 5808 7342 5817
rect 7286 5743 7342 5752
rect 7300 5234 7328 5743
rect 7392 5302 7420 6598
rect 7380 5296 7432 5302
rect 7380 5238 7432 5244
rect 7288 5228 7340 5234
rect 7288 5170 7340 5176
rect 7380 5024 7432 5030
rect 7380 4966 7432 4972
rect 7288 4140 7340 4146
rect 7288 4082 7340 4088
rect 7300 3466 7328 4082
rect 7392 3670 7420 4966
rect 7484 4434 7512 11086
rect 7668 10606 7696 11494
rect 7748 11280 7800 11286
rect 7748 11222 7800 11228
rect 7760 11121 7788 11222
rect 7746 11112 7802 11121
rect 7746 11047 7802 11056
rect 7656 10600 7708 10606
rect 7656 10542 7708 10548
rect 7564 9920 7616 9926
rect 7564 9862 7616 9868
rect 7576 8974 7604 9862
rect 7564 8968 7616 8974
rect 7564 8910 7616 8916
rect 7576 8838 7604 8910
rect 7564 8832 7616 8838
rect 7564 8774 7616 8780
rect 7564 7880 7616 7886
rect 7564 7822 7616 7828
rect 7576 7478 7604 7822
rect 7564 7472 7616 7478
rect 7564 7414 7616 7420
rect 7668 7290 7696 10542
rect 7852 10010 7880 12038
rect 8588 11898 8616 12174
rect 8668 12096 8720 12102
rect 8668 12038 8720 12044
rect 8576 11892 8628 11898
rect 8576 11834 8628 11840
rect 8174 11452 8482 11461
rect 8174 11450 8180 11452
rect 8236 11450 8260 11452
rect 8316 11450 8340 11452
rect 8396 11450 8420 11452
rect 8476 11450 8482 11452
rect 8236 11398 8238 11450
rect 8418 11398 8420 11450
rect 8174 11396 8180 11398
rect 8236 11396 8260 11398
rect 8316 11396 8340 11398
rect 8396 11396 8420 11398
rect 8476 11396 8482 11398
rect 8174 11387 8482 11396
rect 8588 11082 8616 11834
rect 8576 11076 8628 11082
rect 8576 11018 8628 11024
rect 8484 11008 8536 11014
rect 8536 10956 8616 10962
rect 8484 10950 8616 10956
rect 8496 10934 8616 10950
rect 8174 10364 8482 10373
rect 8174 10362 8180 10364
rect 8236 10362 8260 10364
rect 8316 10362 8340 10364
rect 8396 10362 8420 10364
rect 8476 10362 8482 10364
rect 8236 10310 8238 10362
rect 8418 10310 8420 10362
rect 8174 10308 8180 10310
rect 8236 10308 8260 10310
rect 8316 10308 8340 10310
rect 8396 10308 8420 10310
rect 8476 10308 8482 10310
rect 8174 10299 8482 10308
rect 7760 9982 7880 10010
rect 7760 8378 7788 9982
rect 7840 9920 7892 9926
rect 7840 9862 7892 9868
rect 7852 9586 7880 9862
rect 7840 9580 7892 9586
rect 7840 9522 7892 9528
rect 7932 9512 7984 9518
rect 7932 9454 7984 9460
rect 7944 9382 7972 9454
rect 7932 9376 7984 9382
rect 7932 9318 7984 9324
rect 7944 8634 7972 9318
rect 8174 9276 8482 9285
rect 8174 9274 8180 9276
rect 8236 9274 8260 9276
rect 8316 9274 8340 9276
rect 8396 9274 8420 9276
rect 8476 9274 8482 9276
rect 8236 9222 8238 9274
rect 8418 9222 8420 9274
rect 8174 9220 8180 9222
rect 8236 9220 8260 9222
rect 8316 9220 8340 9222
rect 8396 9220 8420 9222
rect 8476 9220 8482 9222
rect 8174 9211 8482 9220
rect 8024 9104 8076 9110
rect 8024 9046 8076 9052
rect 7932 8628 7984 8634
rect 7932 8570 7984 8576
rect 7760 8350 7880 8378
rect 7748 8288 7800 8294
rect 7748 8230 7800 8236
rect 7760 7546 7788 8230
rect 7748 7540 7800 7546
rect 7748 7482 7800 7488
rect 7576 7262 7696 7290
rect 7576 4554 7604 7262
rect 7852 6610 7880 8350
rect 8036 7886 8064 9046
rect 8208 8492 8260 8498
rect 8208 8434 8260 8440
rect 8220 8401 8248 8434
rect 8206 8392 8262 8401
rect 8392 8356 8444 8362
rect 8262 8336 8392 8344
rect 8206 8327 8392 8336
rect 8220 8316 8392 8327
rect 8392 8298 8444 8304
rect 8174 8188 8482 8197
rect 8174 8186 8180 8188
rect 8236 8186 8260 8188
rect 8316 8186 8340 8188
rect 8396 8186 8420 8188
rect 8476 8186 8482 8188
rect 8236 8134 8238 8186
rect 8418 8134 8420 8186
rect 8174 8132 8180 8134
rect 8236 8132 8260 8134
rect 8316 8132 8340 8134
rect 8396 8132 8420 8134
rect 8476 8132 8482 8134
rect 8174 8123 8482 8132
rect 8300 7948 8352 7954
rect 8300 7890 8352 7896
rect 8024 7880 8076 7886
rect 8024 7822 8076 7828
rect 8208 7744 8260 7750
rect 8208 7686 8260 7692
rect 8220 7546 8248 7686
rect 8208 7540 8260 7546
rect 8208 7482 8260 7488
rect 8024 7336 8076 7342
rect 8312 7290 8340 7890
rect 8076 7284 8340 7290
rect 8024 7278 8340 7284
rect 8036 7262 8340 7278
rect 8036 6934 8064 7262
rect 8174 7100 8482 7109
rect 8174 7098 8180 7100
rect 8236 7098 8260 7100
rect 8316 7098 8340 7100
rect 8396 7098 8420 7100
rect 8476 7098 8482 7100
rect 8236 7046 8238 7098
rect 8418 7046 8420 7098
rect 8174 7044 8180 7046
rect 8236 7044 8260 7046
rect 8316 7044 8340 7046
rect 8396 7044 8420 7046
rect 8476 7044 8482 7046
rect 8174 7035 8482 7044
rect 8024 6928 8076 6934
rect 8024 6870 8076 6876
rect 7932 6792 7984 6798
rect 8588 6769 8616 10934
rect 7932 6734 7984 6740
rect 8574 6760 8630 6769
rect 7760 6582 7880 6610
rect 7760 6361 7788 6582
rect 7840 6452 7892 6458
rect 7840 6394 7892 6400
rect 7746 6352 7802 6361
rect 7746 6287 7802 6296
rect 7760 5817 7788 6287
rect 7852 5914 7880 6394
rect 7840 5908 7892 5914
rect 7840 5850 7892 5856
rect 7746 5808 7802 5817
rect 7746 5743 7802 5752
rect 7656 5704 7708 5710
rect 7654 5672 7656 5681
rect 7708 5672 7710 5681
rect 7654 5607 7710 5616
rect 7840 5568 7892 5574
rect 7840 5510 7892 5516
rect 7564 4548 7616 4554
rect 7564 4490 7616 4496
rect 7746 4448 7802 4457
rect 7484 4406 7696 4434
rect 7472 4276 7524 4282
rect 7472 4218 7524 4224
rect 7484 4185 7512 4218
rect 7564 4208 7616 4214
rect 7470 4176 7526 4185
rect 7564 4150 7616 4156
rect 7470 4111 7526 4120
rect 7472 4004 7524 4010
rect 7472 3946 7524 3952
rect 7484 3777 7512 3946
rect 7470 3768 7526 3777
rect 7470 3703 7472 3712
rect 7524 3703 7526 3712
rect 7472 3674 7524 3680
rect 7380 3664 7432 3670
rect 7484 3643 7512 3674
rect 7380 3606 7432 3612
rect 7380 3528 7432 3534
rect 7380 3470 7432 3476
rect 7288 3460 7340 3466
rect 7288 3402 7340 3408
rect 7392 3346 7420 3470
rect 7472 3460 7524 3466
rect 7472 3402 7524 3408
rect 7300 3318 7420 3346
rect 7196 2440 7248 2446
rect 7196 2382 7248 2388
rect 7104 1760 7156 1766
rect 7104 1702 7156 1708
rect 7012 1420 7064 1426
rect 7012 1362 7064 1368
rect 7300 1290 7328 3318
rect 7378 3224 7434 3233
rect 7484 3194 7512 3402
rect 7378 3159 7434 3168
rect 7472 3188 7524 3194
rect 7392 3126 7420 3159
rect 7472 3130 7524 3136
rect 7380 3120 7432 3126
rect 7380 3062 7432 3068
rect 7380 2916 7432 2922
rect 7380 2858 7432 2864
rect 7288 1284 7340 1290
rect 7288 1226 7340 1232
rect 6092 1216 6144 1222
rect 6092 1158 6144 1164
rect 5908 1148 5960 1154
rect 5908 1090 5960 1096
rect 4896 1080 4948 1086
rect 4896 1022 4948 1028
rect 4528 1012 4580 1018
rect 4528 954 4580 960
rect 7208 870 7328 898
rect 3240 808 3292 814
rect 3240 750 3292 756
rect 7208 746 7236 870
rect 7300 800 7328 870
rect 7392 800 7420 2858
rect 7472 2440 7524 2446
rect 7472 2382 7524 2388
rect 7484 1562 7512 2382
rect 7472 1556 7524 1562
rect 7472 1498 7524 1504
rect 7472 1420 7524 1426
rect 7472 1362 7524 1368
rect 7484 800 7512 1362
rect 7576 800 7604 4150
rect 7668 800 7696 4406
rect 7746 4383 7802 4392
rect 7760 4282 7788 4383
rect 7748 4276 7800 4282
rect 7748 4218 7800 4224
rect 7748 3936 7800 3942
rect 7748 3878 7800 3884
rect 7760 3738 7788 3878
rect 7748 3732 7800 3738
rect 7748 3674 7800 3680
rect 7748 3596 7800 3602
rect 7748 3538 7800 3544
rect 7760 800 7788 3538
rect 7852 1766 7880 5510
rect 7944 5030 7972 6734
rect 8574 6695 8630 6704
rect 8024 6656 8076 6662
rect 8024 6598 8076 6604
rect 7932 5024 7984 5030
rect 7932 4966 7984 4972
rect 7944 4826 7972 4966
rect 7932 4820 7984 4826
rect 7932 4762 7984 4768
rect 7932 4548 7984 4554
rect 7932 4490 7984 4496
rect 7840 1760 7892 1766
rect 7840 1702 7892 1708
rect 7944 1578 7972 4490
rect 8036 1714 8064 6598
rect 8576 6112 8628 6118
rect 8576 6054 8628 6060
rect 8174 6012 8482 6021
rect 8174 6010 8180 6012
rect 8236 6010 8260 6012
rect 8316 6010 8340 6012
rect 8396 6010 8420 6012
rect 8476 6010 8482 6012
rect 8236 5958 8238 6010
rect 8418 5958 8420 6010
rect 8174 5956 8180 5958
rect 8236 5956 8260 5958
rect 8316 5956 8340 5958
rect 8396 5956 8420 5958
rect 8476 5956 8482 5958
rect 8174 5947 8482 5956
rect 8588 5846 8616 6054
rect 8680 5953 8708 12038
rect 8760 9580 8812 9586
rect 8760 9522 8812 9528
rect 8772 9178 8800 9522
rect 8760 9172 8812 9178
rect 8760 9114 8812 9120
rect 8760 6656 8812 6662
rect 8760 6598 8812 6604
rect 8666 5944 8722 5953
rect 8666 5879 8722 5888
rect 8576 5840 8628 5846
rect 8206 5808 8262 5817
rect 8576 5782 8628 5788
rect 8206 5743 8262 5752
rect 8220 5234 8248 5743
rect 8680 5710 8708 5879
rect 8668 5704 8720 5710
rect 8668 5646 8720 5652
rect 8208 5228 8260 5234
rect 8208 5170 8260 5176
rect 8174 4924 8482 4933
rect 8174 4922 8180 4924
rect 8236 4922 8260 4924
rect 8316 4922 8340 4924
rect 8396 4922 8420 4924
rect 8476 4922 8482 4924
rect 8236 4870 8238 4922
rect 8418 4870 8420 4922
rect 8174 4868 8180 4870
rect 8236 4868 8260 4870
rect 8316 4868 8340 4870
rect 8396 4868 8420 4870
rect 8476 4868 8482 4870
rect 8174 4859 8482 4868
rect 8666 4856 8722 4865
rect 8392 4820 8444 4826
rect 8666 4791 8722 4800
rect 8392 4762 8444 4768
rect 8404 4622 8432 4762
rect 8392 4616 8444 4622
rect 8392 4558 8444 4564
rect 8576 4616 8628 4622
rect 8576 4558 8628 4564
rect 8116 4548 8168 4554
rect 8116 4490 8168 4496
rect 8128 4010 8156 4490
rect 8588 4457 8616 4558
rect 8680 4554 8708 4791
rect 8668 4548 8720 4554
rect 8668 4490 8720 4496
rect 8574 4448 8630 4457
rect 8574 4383 8630 4392
rect 8116 4004 8168 4010
rect 8116 3946 8168 3952
rect 8174 3836 8482 3845
rect 8174 3834 8180 3836
rect 8236 3834 8260 3836
rect 8316 3834 8340 3836
rect 8396 3834 8420 3836
rect 8476 3834 8482 3836
rect 8236 3782 8238 3834
rect 8418 3782 8420 3834
rect 8174 3780 8180 3782
rect 8236 3780 8260 3782
rect 8316 3780 8340 3782
rect 8396 3780 8420 3782
rect 8476 3780 8482 3782
rect 8174 3771 8482 3780
rect 8484 3664 8536 3670
rect 8484 3606 8536 3612
rect 8116 3596 8168 3602
rect 8116 3538 8168 3544
rect 8128 3126 8156 3538
rect 8208 3392 8260 3398
rect 8208 3334 8260 3340
rect 8220 3233 8248 3334
rect 8206 3224 8262 3233
rect 8206 3159 8262 3168
rect 8116 3120 8168 3126
rect 8116 3062 8168 3068
rect 8496 2922 8524 3606
rect 8588 3602 8616 4383
rect 8772 4146 8800 6598
rect 8760 4140 8812 4146
rect 8760 4082 8812 4088
rect 8666 3904 8722 3913
rect 8666 3839 8722 3848
rect 8576 3596 8628 3602
rect 8576 3538 8628 3544
rect 8680 3126 8708 3839
rect 8772 3534 8800 4082
rect 8864 3602 8892 12582
rect 9232 12442 9260 12650
rect 9220 12436 9272 12442
rect 9600 12434 9628 13126
rect 9220 12378 9272 12384
rect 9416 12406 9628 12434
rect 9692 12434 9720 13126
rect 10968 12640 11020 12646
rect 10966 12608 10968 12617
rect 11020 12608 11022 12617
rect 10966 12543 11022 12552
rect 9692 12406 9812 12434
rect 9036 11280 9088 11286
rect 9036 11222 9088 11228
rect 8944 10532 8996 10538
rect 8944 10474 8996 10480
rect 8956 3777 8984 10474
rect 8942 3768 8998 3777
rect 8942 3703 8998 3712
rect 8852 3596 8904 3602
rect 8904 3556 8984 3584
rect 8852 3538 8904 3544
rect 8760 3528 8812 3534
rect 8760 3470 8812 3476
rect 8758 3224 8814 3233
rect 8758 3159 8814 3168
rect 8668 3120 8720 3126
rect 8668 3062 8720 3068
rect 8484 2916 8536 2922
rect 8484 2858 8536 2864
rect 8574 2816 8630 2825
rect 8174 2748 8482 2757
rect 8574 2751 8630 2760
rect 8174 2746 8180 2748
rect 8236 2746 8260 2748
rect 8316 2746 8340 2748
rect 8396 2746 8420 2748
rect 8476 2746 8482 2748
rect 8236 2694 8238 2746
rect 8418 2694 8420 2746
rect 8174 2692 8180 2694
rect 8236 2692 8260 2694
rect 8316 2692 8340 2694
rect 8396 2692 8420 2694
rect 8476 2692 8482 2694
rect 8174 2683 8482 2692
rect 8116 2644 8168 2650
rect 8116 2586 8168 2592
rect 8128 2446 8156 2586
rect 8300 2576 8352 2582
rect 8300 2518 8352 2524
rect 8116 2440 8168 2446
rect 8116 2382 8168 2388
rect 8128 1902 8156 2382
rect 8312 1970 8340 2518
rect 8300 1964 8352 1970
rect 8300 1906 8352 1912
rect 8116 1896 8168 1902
rect 8116 1838 8168 1844
rect 8036 1686 8248 1714
rect 7944 1550 8156 1578
rect 8220 1562 8248 1686
rect 8024 1488 8076 1494
rect 8024 1430 8076 1436
rect 7932 1352 7984 1358
rect 7932 1294 7984 1300
rect 7840 1284 7892 1290
rect 7840 1226 7892 1232
rect 7852 800 7880 1226
rect 7944 800 7972 1294
rect 8036 800 8064 1430
rect 8128 800 8156 1550
rect 8208 1556 8260 1562
rect 8208 1498 8260 1504
rect 8588 1442 8616 2751
rect 8312 1414 8616 1442
rect 8208 1012 8260 1018
rect 8208 954 8260 960
rect 8220 800 8248 954
rect 8312 800 8340 1414
rect 8576 1216 8628 1222
rect 8576 1158 8628 1164
rect 8392 1080 8444 1086
rect 8392 1022 8444 1028
rect 8404 800 8432 1022
rect 8588 800 8616 1158
rect 8680 800 8708 3062
rect 8772 3058 8800 3159
rect 8760 3052 8812 3058
rect 8760 2994 8812 3000
rect 8760 2916 8812 2922
rect 8760 2858 8812 2864
rect 8852 2916 8904 2922
rect 8852 2858 8904 2864
rect 8772 1970 8800 2858
rect 8760 1964 8812 1970
rect 8760 1906 8812 1912
rect 8760 1760 8812 1766
rect 8760 1702 8812 1708
rect 8772 800 8800 1702
rect 8864 1494 8892 2858
rect 8852 1488 8904 1494
rect 8852 1430 8904 1436
rect 8956 800 8984 3556
rect 9048 2446 9076 11222
rect 9220 11076 9272 11082
rect 9220 11018 9272 11024
rect 9128 10056 9180 10062
rect 9128 9998 9180 10004
rect 9140 6662 9168 9998
rect 9232 8022 9260 11018
rect 9312 10668 9364 10674
rect 9312 10610 9364 10616
rect 9220 8016 9272 8022
rect 9220 7958 9272 7964
rect 9220 7880 9272 7886
rect 9220 7822 9272 7828
rect 9232 7585 9260 7822
rect 9218 7576 9274 7585
rect 9218 7511 9274 7520
rect 9128 6656 9180 6662
rect 9128 6598 9180 6604
rect 9220 6656 9272 6662
rect 9220 6598 9272 6604
rect 9126 6488 9182 6497
rect 9126 6423 9182 6432
rect 9140 6322 9168 6423
rect 9128 6316 9180 6322
rect 9128 6258 9180 6264
rect 9128 5840 9180 5846
rect 9128 5782 9180 5788
rect 9140 5710 9168 5782
rect 9128 5704 9180 5710
rect 9128 5646 9180 5652
rect 9232 4604 9260 6598
rect 9140 4576 9260 4604
rect 9036 2440 9088 2446
rect 9036 2382 9088 2388
rect 9034 2136 9090 2145
rect 9034 2071 9090 2080
rect 9048 800 9076 2071
rect 9140 800 9168 4576
rect 9218 3360 9274 3369
rect 9218 3295 9274 3304
rect 9232 3126 9260 3295
rect 9220 3120 9272 3126
rect 9220 3062 9272 3068
rect 9220 2984 9272 2990
rect 9220 2926 9272 2932
rect 9232 2582 9260 2926
rect 9220 2576 9272 2582
rect 9220 2518 9272 2524
rect 9220 2440 9272 2446
rect 9218 2408 9220 2417
rect 9272 2408 9274 2417
rect 9218 2343 9274 2352
rect 9220 2304 9272 2310
rect 9220 2246 9272 2252
rect 9232 2106 9260 2246
rect 9220 2100 9272 2106
rect 9220 2042 9272 2048
rect 9324 800 9352 10610
rect 9416 3058 9444 12406
rect 9680 11552 9732 11558
rect 9680 11494 9732 11500
rect 9588 10464 9640 10470
rect 9588 10406 9640 10412
rect 9494 8664 9550 8673
rect 9494 8599 9550 8608
rect 9508 8566 9536 8599
rect 9496 8560 9548 8566
rect 9496 8502 9548 8508
rect 9496 7336 9548 7342
rect 9494 7304 9496 7313
rect 9548 7304 9550 7313
rect 9494 7239 9550 7248
rect 9494 6896 9550 6905
rect 9494 6831 9550 6840
rect 9508 6798 9536 6831
rect 9496 6792 9548 6798
rect 9496 6734 9548 6740
rect 9600 5760 9628 10406
rect 9692 6798 9720 11494
rect 9784 9761 9812 12406
rect 10968 12368 11020 12374
rect 10968 12310 11020 12316
rect 10048 12096 10100 12102
rect 10048 12038 10100 12044
rect 10324 12096 10376 12102
rect 10324 12038 10376 12044
rect 9956 11076 10008 11082
rect 9956 11018 10008 11024
rect 9770 9752 9826 9761
rect 9770 9687 9826 9696
rect 9862 9616 9918 9625
rect 9862 9551 9864 9560
rect 9916 9551 9918 9560
rect 9864 9522 9916 9528
rect 9772 9376 9824 9382
rect 9772 9318 9824 9324
rect 9784 8838 9812 9318
rect 9772 8832 9824 8838
rect 9772 8774 9824 8780
rect 9862 7984 9918 7993
rect 9862 7919 9918 7928
rect 9876 7886 9904 7919
rect 9864 7880 9916 7886
rect 9864 7822 9916 7828
rect 9680 6792 9732 6798
rect 9680 6734 9732 6740
rect 9770 6488 9826 6497
rect 9770 6423 9772 6432
rect 9824 6423 9826 6432
rect 9772 6394 9824 6400
rect 9864 6316 9916 6322
rect 9864 6258 9916 6264
rect 9772 6112 9824 6118
rect 9770 6080 9772 6089
rect 9824 6080 9826 6089
rect 9770 6015 9826 6024
rect 9876 5914 9904 6258
rect 9772 5908 9824 5914
rect 9772 5850 9824 5856
rect 9864 5908 9916 5914
rect 9864 5850 9916 5856
rect 9784 5794 9812 5850
rect 9784 5766 9902 5794
rect 9874 5760 9902 5766
rect 9600 5732 9720 5760
rect 9874 5732 9904 5760
rect 9496 5636 9548 5642
rect 9496 5578 9548 5584
rect 9508 5409 9536 5578
rect 9692 5522 9720 5732
rect 9876 5624 9904 5732
rect 9600 5494 9720 5522
rect 9784 5596 9904 5624
rect 9494 5400 9550 5409
rect 9494 5335 9550 5344
rect 9496 5092 9548 5098
rect 9496 5034 9548 5040
rect 9508 4554 9536 5034
rect 9496 4548 9548 4554
rect 9496 4490 9548 4496
rect 9496 3528 9548 3534
rect 9496 3470 9548 3476
rect 9508 3194 9536 3470
rect 9496 3188 9548 3194
rect 9496 3130 9548 3136
rect 9404 3052 9456 3058
rect 9600 3040 9628 5494
rect 9678 5400 9734 5409
rect 9678 5335 9734 5344
rect 9692 4622 9720 5335
rect 9680 4616 9732 4622
rect 9680 4558 9732 4564
rect 9680 3392 9732 3398
rect 9680 3334 9732 3340
rect 9404 2994 9456 3000
rect 9508 3012 9628 3040
rect 9416 800 9444 2994
rect 9508 2514 9536 3012
rect 9692 2938 9720 3334
rect 9600 2922 9720 2938
rect 9588 2916 9720 2922
rect 9640 2910 9720 2916
rect 9588 2858 9640 2864
rect 9496 2508 9548 2514
rect 9496 2450 9548 2456
rect 9496 1964 9548 1970
rect 9496 1906 9548 1912
rect 9508 800 9536 1906
rect 9680 1556 9732 1562
rect 9680 1498 9732 1504
rect 9588 1488 9640 1494
rect 9588 1430 9640 1436
rect 9600 800 9628 1430
rect 9692 800 9720 1498
rect 9784 800 9812 5596
rect 9864 5092 9916 5098
rect 9864 5034 9916 5040
rect 9876 5001 9904 5034
rect 9862 4992 9918 5001
rect 9862 4927 9918 4936
rect 9864 4480 9916 4486
rect 9864 4422 9916 4428
rect 9876 3602 9904 4422
rect 9864 3596 9916 3602
rect 9864 3538 9916 3544
rect 9968 3482 9996 11018
rect 10060 10742 10088 12038
rect 10048 10736 10100 10742
rect 10048 10678 10100 10684
rect 10140 10668 10192 10674
rect 10140 10610 10192 10616
rect 10048 10056 10100 10062
rect 10048 9998 10100 10004
rect 10060 9722 10088 9998
rect 10048 9716 10100 9722
rect 10048 9658 10100 9664
rect 10046 8120 10102 8129
rect 10046 8055 10102 8064
rect 10060 7750 10088 8055
rect 10048 7744 10100 7750
rect 10048 7686 10100 7692
rect 10048 6452 10100 6458
rect 10048 6394 10100 6400
rect 10060 5370 10088 6394
rect 10048 5364 10100 5370
rect 10048 5306 10100 5312
rect 10046 5128 10102 5137
rect 10046 5063 10102 5072
rect 10060 4865 10088 5063
rect 10046 4856 10102 4865
rect 10046 4791 10102 4800
rect 10060 4690 10088 4791
rect 10048 4684 10100 4690
rect 10048 4626 10100 4632
rect 10048 3732 10100 3738
rect 10048 3674 10100 3680
rect 9876 3454 9996 3482
rect 9876 800 9904 3454
rect 9956 3392 10008 3398
rect 9956 3334 10008 3340
rect 9968 800 9996 3334
rect 10060 800 10088 3674
rect 10152 800 10180 10610
rect 10232 9920 10284 9926
rect 10232 9862 10284 9868
rect 10244 6089 10272 9862
rect 10336 9489 10364 12038
rect 10416 11552 10468 11558
rect 10416 11494 10468 11500
rect 10322 9480 10378 9489
rect 10322 9415 10378 9424
rect 10336 8498 10364 9415
rect 10428 8498 10456 11494
rect 10980 11286 11008 12310
rect 10968 11280 11020 11286
rect 10968 11222 11020 11228
rect 10784 9988 10836 9994
rect 10784 9930 10836 9936
rect 10692 9580 10744 9586
rect 10692 9522 10744 9528
rect 10600 9376 10652 9382
rect 10600 9318 10652 9324
rect 10612 9058 10640 9318
rect 10704 9178 10732 9522
rect 10692 9172 10744 9178
rect 10692 9114 10744 9120
rect 10612 9030 10732 9058
rect 10600 8968 10652 8974
rect 10598 8936 10600 8945
rect 10652 8936 10654 8945
rect 10598 8871 10654 8880
rect 10600 8832 10652 8838
rect 10600 8774 10652 8780
rect 10324 8492 10376 8498
rect 10324 8434 10376 8440
rect 10416 8492 10468 8498
rect 10416 8434 10468 8440
rect 10508 8084 10560 8090
rect 10508 8026 10560 8032
rect 10520 6798 10548 8026
rect 10612 7002 10640 8774
rect 10704 8378 10732 9030
rect 10796 8634 10824 9930
rect 10980 9518 11008 11222
rect 10968 9512 11020 9518
rect 10968 9454 11020 9460
rect 10784 8628 10836 8634
rect 10784 8570 10836 8576
rect 10796 8514 10824 8570
rect 10796 8486 10916 8514
rect 10888 8430 10916 8486
rect 10876 8424 10928 8430
rect 10704 8350 10824 8378
rect 10876 8366 10928 8372
rect 10966 8392 11022 8401
rect 10692 7744 10744 7750
rect 10692 7686 10744 7692
rect 10704 7546 10732 7686
rect 10692 7540 10744 7546
rect 10692 7482 10744 7488
rect 10600 6996 10652 7002
rect 10600 6938 10652 6944
rect 10508 6792 10560 6798
rect 10508 6734 10560 6740
rect 10324 6724 10376 6730
rect 10324 6666 10376 6672
rect 10692 6724 10744 6730
rect 10692 6666 10744 6672
rect 10230 6080 10286 6089
rect 10230 6015 10286 6024
rect 10230 5808 10286 5817
rect 10230 5743 10232 5752
rect 10284 5743 10286 5752
rect 10232 5714 10284 5720
rect 10336 5681 10364 6666
rect 10600 6656 10652 6662
rect 10600 6598 10652 6604
rect 10612 6288 10640 6598
rect 10600 6282 10652 6288
rect 10600 6224 10652 6230
rect 10322 5672 10378 5681
rect 10322 5607 10378 5616
rect 10232 5568 10284 5574
rect 10232 5510 10284 5516
rect 10244 5114 10272 5510
rect 10508 5296 10560 5302
rect 10508 5238 10560 5244
rect 10244 5086 10364 5114
rect 10336 4672 10364 5086
rect 10416 5024 10468 5030
rect 10416 4966 10468 4972
rect 10428 4826 10456 4966
rect 10416 4820 10468 4826
rect 10416 4762 10468 4768
rect 10244 4644 10364 4672
rect 10244 2802 10272 4644
rect 10322 4584 10378 4593
rect 10322 4519 10378 4528
rect 10336 3210 10364 4519
rect 10520 4146 10548 5238
rect 10600 5228 10652 5234
rect 10600 5170 10652 5176
rect 10612 4758 10640 5170
rect 10600 4752 10652 4758
rect 10600 4694 10652 4700
rect 10508 4140 10560 4146
rect 10508 4082 10560 4088
rect 10508 3664 10560 3670
rect 10508 3606 10560 3612
rect 10520 3534 10548 3606
rect 10508 3528 10560 3534
rect 10506 3496 10508 3505
rect 10560 3496 10562 3505
rect 10506 3431 10562 3440
rect 10704 3398 10732 6666
rect 10796 4826 10824 8350
rect 10966 8327 10968 8336
rect 11020 8327 11022 8336
rect 10968 8298 11020 8304
rect 10968 8084 11020 8090
rect 10968 8026 11020 8032
rect 10874 7712 10930 7721
rect 10874 7647 10930 7656
rect 10888 7313 10916 7647
rect 10874 7304 10930 7313
rect 10874 7239 10930 7248
rect 10888 6866 10916 7239
rect 10876 6860 10928 6866
rect 10876 6802 10928 6808
rect 10980 6322 11008 8026
rect 10968 6316 11020 6322
rect 10968 6258 11020 6264
rect 10968 6112 11020 6118
rect 10874 6080 10930 6089
rect 10968 6054 11020 6060
rect 10874 6015 10930 6024
rect 10784 4820 10836 4826
rect 10784 4762 10836 4768
rect 10888 3670 10916 6015
rect 10980 5642 11008 6054
rect 10968 5636 11020 5642
rect 10968 5578 11020 5584
rect 10968 5092 11020 5098
rect 10968 5034 11020 5040
rect 10980 4214 11008 5034
rect 10968 4208 11020 4214
rect 10968 4150 11020 4156
rect 10876 3664 10928 3670
rect 10876 3606 10928 3612
rect 10784 3596 10836 3602
rect 10784 3538 10836 3544
rect 10692 3392 10744 3398
rect 10692 3334 10744 3340
rect 10336 3182 10548 3210
rect 10416 2848 10468 2854
rect 10244 2774 10364 2802
rect 10416 2790 10468 2796
rect 10230 2680 10286 2689
rect 10230 2615 10286 2624
rect 10244 800 10272 2615
rect 10336 800 10364 2774
rect 10428 1442 10456 2790
rect 10520 1562 10548 3182
rect 10692 3188 10744 3194
rect 10692 3130 10744 3136
rect 10600 2984 10652 2990
rect 10704 2961 10732 3130
rect 10796 2990 10824 3538
rect 10876 3392 10928 3398
rect 10876 3334 10928 3340
rect 10784 2984 10836 2990
rect 10600 2926 10652 2932
rect 10690 2952 10746 2961
rect 10612 1562 10640 2926
rect 10784 2926 10836 2932
rect 10690 2887 10746 2896
rect 10692 2440 10744 2446
rect 10692 2382 10744 2388
rect 10508 1556 10560 1562
rect 10508 1498 10560 1504
rect 10600 1556 10652 1562
rect 10600 1498 10652 1504
rect 10428 1414 10640 1442
rect 10416 1352 10468 1358
rect 10416 1294 10468 1300
rect 10508 1352 10560 1358
rect 10508 1294 10560 1300
rect 10428 1154 10456 1294
rect 10416 1148 10468 1154
rect 10416 1090 10468 1096
rect 10520 800 10548 1294
rect 10612 800 10640 1414
rect 10704 1057 10732 2382
rect 10784 1760 10836 1766
rect 10784 1702 10836 1708
rect 10690 1048 10746 1057
rect 10690 983 10746 992
rect 10796 800 10824 1702
rect 10888 800 10916 3334
rect 10968 2848 11020 2854
rect 10968 2790 11020 2796
rect 10980 2650 11008 2790
rect 10968 2644 11020 2650
rect 10968 2586 11020 2592
rect 11072 2530 11100 13126
rect 11440 12782 11468 13262
rect 12992 13252 13044 13258
rect 12992 13194 13044 13200
rect 11612 13184 11664 13190
rect 11612 13126 11664 13132
rect 12900 13184 12952 13190
rect 12900 13126 12952 13132
rect 11428 12776 11480 12782
rect 11426 12744 11428 12753
rect 11480 12744 11482 12753
rect 11426 12679 11482 12688
rect 11152 12096 11204 12102
rect 11152 12038 11204 12044
rect 11164 9081 11192 12038
rect 11428 10600 11480 10606
rect 11428 10542 11480 10548
rect 11440 10130 11468 10542
rect 11428 10124 11480 10130
rect 11428 10066 11480 10072
rect 11244 10056 11296 10062
rect 11244 9998 11296 10004
rect 11336 10056 11388 10062
rect 11336 9998 11388 10004
rect 11256 9654 11284 9998
rect 11244 9648 11296 9654
rect 11244 9590 11296 9596
rect 11150 9072 11206 9081
rect 11150 9007 11206 9016
rect 11164 8498 11192 9007
rect 11348 8634 11376 9998
rect 11440 8974 11468 10066
rect 11428 8968 11480 8974
rect 11428 8910 11480 8916
rect 11520 8968 11572 8974
rect 11520 8910 11572 8916
rect 11336 8628 11388 8634
rect 11336 8570 11388 8576
rect 11152 8492 11204 8498
rect 11152 8434 11204 8440
rect 11244 8492 11296 8498
rect 11244 8434 11296 8440
rect 11256 8294 11284 8434
rect 11244 8288 11296 8294
rect 11244 8230 11296 8236
rect 11532 8129 11560 8910
rect 11518 8120 11574 8129
rect 11518 8055 11574 8064
rect 11428 6656 11480 6662
rect 11428 6598 11480 6604
rect 11520 6656 11572 6662
rect 11520 6598 11572 6604
rect 11152 6452 11204 6458
rect 11152 6394 11204 6400
rect 11164 6322 11192 6394
rect 11440 6390 11468 6598
rect 11532 6497 11560 6598
rect 11518 6488 11574 6497
rect 11518 6423 11574 6432
rect 11428 6384 11480 6390
rect 11428 6326 11480 6332
rect 11152 6316 11204 6322
rect 11152 6258 11204 6264
rect 11152 6112 11204 6118
rect 11152 6054 11204 6060
rect 10980 2502 11100 2530
rect 10980 2446 11008 2502
rect 10968 2440 11020 2446
rect 10968 2382 11020 2388
rect 10980 1426 11008 2382
rect 10968 1420 11020 1426
rect 10968 1362 11020 1368
rect 11164 800 11192 6054
rect 11520 5160 11572 5166
rect 11520 5102 11572 5108
rect 11532 5001 11560 5102
rect 11518 4992 11574 5001
rect 11518 4927 11574 4936
rect 11520 4072 11572 4078
rect 11520 4014 11572 4020
rect 11532 3602 11560 4014
rect 11520 3596 11572 3602
rect 11520 3538 11572 3544
rect 11532 3194 11560 3538
rect 11520 3188 11572 3194
rect 11520 3130 11572 3136
rect 11428 2916 11480 2922
rect 11428 2858 11480 2864
rect 11336 2848 11388 2854
rect 11336 2790 11388 2796
rect 11348 2378 11376 2790
rect 11336 2372 11388 2378
rect 11336 2314 11388 2320
rect 11440 800 11468 2858
rect 11624 2446 11652 13126
rect 12912 12850 12940 13126
rect 13004 12986 13032 13194
rect 14188 13184 14240 13190
rect 14188 13126 14240 13132
rect 15108 13184 15160 13190
rect 15108 13126 15160 13132
rect 12992 12980 13044 12986
rect 12992 12922 13044 12928
rect 12900 12844 12952 12850
rect 12900 12786 12952 12792
rect 11704 12640 11756 12646
rect 11704 12582 11756 12588
rect 11716 11762 11744 12582
rect 12440 12096 12492 12102
rect 12440 12038 12492 12044
rect 11704 11756 11756 11762
rect 11704 11698 11756 11704
rect 11716 8090 11744 11698
rect 12452 11558 12480 12038
rect 12440 11552 12492 11558
rect 12440 11494 12492 11500
rect 12808 11552 12860 11558
rect 12808 11494 12860 11500
rect 12348 11144 12400 11150
rect 12348 11086 12400 11092
rect 11796 10668 11848 10674
rect 11796 10610 11848 10616
rect 11808 10266 11836 10610
rect 12256 10464 12308 10470
rect 12256 10406 12308 10412
rect 11796 10260 11848 10266
rect 11796 10202 11848 10208
rect 12268 9722 12296 10406
rect 12256 9716 12308 9722
rect 12256 9658 12308 9664
rect 12268 9178 12296 9658
rect 12256 9172 12308 9178
rect 12256 9114 12308 9120
rect 11796 8832 11848 8838
rect 11796 8774 11848 8780
rect 11808 8498 11836 8774
rect 11796 8492 11848 8498
rect 11796 8434 11848 8440
rect 11808 8294 11836 8434
rect 11796 8288 11848 8294
rect 11796 8230 11848 8236
rect 11704 8084 11756 8090
rect 11704 8026 11756 8032
rect 11702 7984 11758 7993
rect 11702 7919 11758 7928
rect 11716 7818 11744 7919
rect 11704 7812 11756 7818
rect 11704 7754 11756 7760
rect 11808 7342 11836 8230
rect 11978 7440 12034 7449
rect 11978 7375 12034 7384
rect 11796 7336 11848 7342
rect 11796 7278 11848 7284
rect 11808 7002 11836 7278
rect 11796 6996 11848 7002
rect 11796 6938 11848 6944
rect 11796 6112 11848 6118
rect 11796 6054 11848 6060
rect 11886 6080 11942 6089
rect 11704 5704 11756 5710
rect 11704 5646 11756 5652
rect 11716 4690 11744 5646
rect 11704 4684 11756 4690
rect 11704 4626 11756 4632
rect 11704 3052 11756 3058
rect 11704 2994 11756 3000
rect 11716 2961 11744 2994
rect 11702 2952 11758 2961
rect 11702 2887 11758 2896
rect 11808 2774 11836 6054
rect 11886 6015 11942 6024
rect 11900 5234 11928 6015
rect 11888 5228 11940 5234
rect 11888 5170 11940 5176
rect 11992 5030 12020 7375
rect 12072 7268 12124 7274
rect 12072 7210 12124 7216
rect 11980 5024 12032 5030
rect 11980 4966 12032 4972
rect 12084 2774 12112 7210
rect 12256 6724 12308 6730
rect 12256 6666 12308 6672
rect 12162 5128 12218 5137
rect 12162 5063 12218 5072
rect 12176 3641 12204 5063
rect 12162 3632 12218 3641
rect 12162 3567 12218 3576
rect 11716 2746 11836 2774
rect 11992 2746 12112 2774
rect 11612 2440 11664 2446
rect 11612 2382 11664 2388
rect 11624 1766 11652 2382
rect 11612 1760 11664 1766
rect 11612 1702 11664 1708
rect 11716 800 11744 2746
rect 11796 2440 11848 2446
rect 11796 2382 11848 2388
rect 11808 1601 11836 2382
rect 11794 1592 11850 1601
rect 11794 1527 11850 1536
rect 11992 800 12020 2746
rect 12268 800 12296 6666
rect 12360 3482 12388 11086
rect 12452 8294 12480 11494
rect 12716 11348 12768 11354
rect 12716 11290 12768 11296
rect 12624 9920 12676 9926
rect 12624 9862 12676 9868
rect 12440 8288 12492 8294
rect 12440 8230 12492 8236
rect 12636 7886 12664 9862
rect 12728 9518 12756 11290
rect 12716 9512 12768 9518
rect 12716 9454 12768 9460
rect 12716 8968 12768 8974
rect 12716 8910 12768 8916
rect 12440 7880 12492 7886
rect 12440 7822 12492 7828
rect 12624 7880 12676 7886
rect 12624 7822 12676 7828
rect 12452 7041 12480 7822
rect 12728 7698 12756 8910
rect 12636 7670 12756 7698
rect 12532 7200 12584 7206
rect 12532 7142 12584 7148
rect 12438 7032 12494 7041
rect 12438 6967 12494 6976
rect 12544 6361 12572 7142
rect 12530 6352 12586 6361
rect 12530 6287 12586 6296
rect 12544 3534 12572 6287
rect 12532 3528 12584 3534
rect 12360 3454 12480 3482
rect 12532 3470 12584 3476
rect 12452 2774 12480 3454
rect 12636 3194 12664 7670
rect 12716 6316 12768 6322
rect 12716 6258 12768 6264
rect 12728 6225 12756 6258
rect 12714 6216 12770 6225
rect 12714 6151 12770 6160
rect 12716 5568 12768 5574
rect 12716 5510 12768 5516
rect 12728 3398 12756 5510
rect 12716 3392 12768 3398
rect 12716 3334 12768 3340
rect 12624 3188 12676 3194
rect 12624 3130 12676 3136
rect 12452 2746 12572 2774
rect 12544 800 12572 2746
rect 12820 800 12848 11494
rect 12912 7206 12940 12786
rect 13004 12730 13032 12922
rect 14200 12753 14228 13126
rect 15120 12986 15148 13126
rect 15212 12986 15240 13262
rect 16948 13252 17000 13258
rect 16948 13194 17000 13200
rect 19708 13252 19760 13258
rect 19708 13194 19760 13200
rect 15844 13184 15896 13190
rect 15844 13126 15896 13132
rect 15398 13084 15706 13093
rect 15398 13082 15404 13084
rect 15460 13082 15484 13084
rect 15540 13082 15564 13084
rect 15620 13082 15644 13084
rect 15700 13082 15706 13084
rect 15460 13030 15462 13082
rect 15642 13030 15644 13082
rect 15398 13028 15404 13030
rect 15460 13028 15484 13030
rect 15540 13028 15564 13030
rect 15620 13028 15644 13030
rect 15700 13028 15706 13030
rect 15398 13019 15706 13028
rect 15108 12980 15160 12986
rect 15108 12922 15160 12928
rect 15200 12980 15252 12986
rect 15200 12922 15252 12928
rect 14186 12744 14242 12753
rect 13004 12714 13216 12730
rect 13004 12708 13228 12714
rect 13004 12702 13176 12708
rect 14186 12679 14242 12688
rect 13176 12650 13228 12656
rect 13268 12096 13320 12102
rect 14188 12096 14240 12102
rect 13268 12038 13320 12044
rect 14186 12064 14188 12073
rect 14648 12096 14700 12102
rect 14240 12064 14242 12073
rect 13084 11144 13136 11150
rect 13084 11086 13136 11092
rect 12992 7404 13044 7410
rect 12992 7346 13044 7352
rect 12900 7200 12952 7206
rect 12900 7142 12952 7148
rect 12900 6248 12952 6254
rect 12900 6190 12952 6196
rect 12912 5302 12940 6190
rect 12900 5296 12952 5302
rect 12900 5238 12952 5244
rect 13004 4826 13032 7346
rect 12992 4820 13044 4826
rect 12992 4762 13044 4768
rect 13004 4486 13032 4762
rect 12992 4480 13044 4486
rect 12992 4422 13044 4428
rect 13096 800 13124 11086
rect 13280 11082 13308 12038
rect 14648 12038 14700 12044
rect 14186 11999 14242 12008
rect 14556 11620 14608 11626
rect 14556 11562 14608 11568
rect 13636 11552 13688 11558
rect 13636 11494 13688 11500
rect 13648 11354 13676 11494
rect 13636 11348 13688 11354
rect 13636 11290 13688 11296
rect 13636 11212 13688 11218
rect 13636 11154 13688 11160
rect 13360 11144 13412 11150
rect 13360 11086 13412 11092
rect 13268 11076 13320 11082
rect 13268 11018 13320 11024
rect 13174 10024 13230 10033
rect 13174 9959 13230 9968
rect 13188 5642 13216 9959
rect 13280 8974 13308 11018
rect 13268 8968 13320 8974
rect 13268 8910 13320 8916
rect 13268 7744 13320 7750
rect 13268 7686 13320 7692
rect 13176 5636 13228 5642
rect 13176 5578 13228 5584
rect 13188 4214 13216 5578
rect 13176 4208 13228 4214
rect 13176 4150 13228 4156
rect 13174 4040 13230 4049
rect 13174 3975 13230 3984
rect 13188 3058 13216 3975
rect 13176 3052 13228 3058
rect 13176 2994 13228 3000
rect 13188 950 13216 2994
rect 13280 2514 13308 7686
rect 13268 2508 13320 2514
rect 13268 2450 13320 2456
rect 13176 944 13228 950
rect 13176 886 13228 892
rect 13372 800 13400 11086
rect 13452 10464 13504 10470
rect 13452 10406 13504 10412
rect 13464 10033 13492 10406
rect 13450 10024 13506 10033
rect 13450 9959 13506 9968
rect 13464 9926 13492 9959
rect 13452 9920 13504 9926
rect 13452 9862 13504 9868
rect 13452 9716 13504 9722
rect 13452 9658 13504 9664
rect 13464 9625 13492 9658
rect 13450 9616 13506 9625
rect 13450 9551 13506 9560
rect 13464 8974 13492 9551
rect 13452 8968 13504 8974
rect 13452 8910 13504 8916
rect 13452 8832 13504 8838
rect 13452 8774 13504 8780
rect 13544 8832 13596 8838
rect 13544 8774 13596 8780
rect 13464 5710 13492 8774
rect 13556 8634 13584 8774
rect 13544 8628 13596 8634
rect 13544 8570 13596 8576
rect 13542 7984 13598 7993
rect 13542 7919 13598 7928
rect 13556 7886 13584 7919
rect 13544 7880 13596 7886
rect 13544 7822 13596 7828
rect 13542 7304 13598 7313
rect 13542 7239 13598 7248
rect 13556 6798 13584 7239
rect 13544 6792 13596 6798
rect 13544 6734 13596 6740
rect 13452 5704 13504 5710
rect 13452 5646 13504 5652
rect 13556 3738 13584 6734
rect 13544 3732 13596 3738
rect 13544 3674 13596 3680
rect 13648 2990 13676 11154
rect 13912 11144 13964 11150
rect 13912 11086 13964 11092
rect 13820 8900 13872 8906
rect 13820 8842 13872 8848
rect 13832 7410 13860 8842
rect 13820 7404 13872 7410
rect 13820 7346 13872 7352
rect 13728 7268 13780 7274
rect 13728 7210 13780 7216
rect 13740 7002 13768 7210
rect 13728 6996 13780 7002
rect 13728 6938 13780 6944
rect 13728 5908 13780 5914
rect 13728 5850 13780 5856
rect 13740 5370 13768 5850
rect 13820 5568 13872 5574
rect 13820 5510 13872 5516
rect 13728 5364 13780 5370
rect 13728 5306 13780 5312
rect 13832 5137 13860 5510
rect 13818 5128 13874 5137
rect 13818 5063 13874 5072
rect 13728 4480 13780 4486
rect 13728 4422 13780 4428
rect 13740 3534 13768 4422
rect 13820 4140 13872 4146
rect 13820 4082 13872 4088
rect 13832 3942 13860 4082
rect 13820 3936 13872 3942
rect 13820 3878 13872 3884
rect 13728 3528 13780 3534
rect 13728 3470 13780 3476
rect 13726 3360 13782 3369
rect 13726 3295 13782 3304
rect 13740 3058 13768 3295
rect 13728 3052 13780 3058
rect 13728 2994 13780 3000
rect 13636 2984 13688 2990
rect 13636 2926 13688 2932
rect 13452 2848 13504 2854
rect 13452 2790 13504 2796
rect 13634 2816 13690 2825
rect 13464 1426 13492 2790
rect 13634 2751 13690 2760
rect 13544 2440 13596 2446
rect 13544 2382 13596 2388
rect 13556 1902 13584 2382
rect 13544 1896 13596 1902
rect 13544 1838 13596 1844
rect 13452 1420 13504 1426
rect 13452 1362 13504 1368
rect 13648 800 13676 2751
rect 13832 2582 13860 3878
rect 13820 2576 13872 2582
rect 13820 2518 13872 2524
rect 13924 800 13952 11086
rect 14188 10736 14240 10742
rect 14188 10678 14240 10684
rect 14096 10056 14148 10062
rect 14096 9998 14148 10004
rect 14108 9654 14136 9998
rect 14200 9926 14228 10678
rect 14280 10532 14332 10538
rect 14280 10474 14332 10480
rect 14188 9920 14240 9926
rect 14188 9862 14240 9868
rect 14096 9648 14148 9654
rect 14200 9625 14228 9862
rect 14096 9590 14148 9596
rect 14186 9616 14242 9625
rect 14186 9551 14242 9560
rect 14188 9444 14240 9450
rect 14188 9386 14240 9392
rect 14200 9353 14228 9386
rect 14186 9344 14242 9353
rect 14186 9279 14242 9288
rect 14004 8424 14056 8430
rect 14004 8366 14056 8372
rect 14016 7478 14044 8366
rect 14096 8288 14148 8294
rect 14096 8230 14148 8236
rect 14004 7472 14056 7478
rect 14004 7414 14056 7420
rect 14108 7410 14136 8230
rect 14200 7410 14228 9279
rect 14096 7404 14148 7410
rect 14096 7346 14148 7352
rect 14188 7404 14240 7410
rect 14188 7346 14240 7352
rect 14096 6792 14148 6798
rect 14094 6760 14096 6769
rect 14148 6760 14150 6769
rect 14094 6695 14150 6704
rect 14096 6316 14148 6322
rect 14016 6276 14096 6304
rect 14016 5710 14044 6276
rect 14096 6258 14148 6264
rect 14188 6180 14240 6186
rect 14188 6122 14240 6128
rect 14200 5710 14228 6122
rect 14004 5704 14056 5710
rect 14004 5646 14056 5652
rect 14188 5704 14240 5710
rect 14188 5646 14240 5652
rect 14016 5234 14044 5646
rect 14004 5228 14056 5234
rect 14004 5170 14056 5176
rect 14016 4622 14044 5170
rect 14186 4856 14242 4865
rect 14096 4820 14148 4826
rect 14186 4791 14242 4800
rect 14096 4762 14148 4768
rect 14004 4616 14056 4622
rect 14004 4558 14056 4564
rect 14108 4298 14136 4762
rect 14200 4690 14228 4791
rect 14188 4684 14240 4690
rect 14188 4626 14240 4632
rect 14016 4270 14136 4298
rect 14016 2774 14044 4270
rect 14093 4140 14145 4146
rect 14093 4082 14145 4088
rect 14188 4140 14240 4146
rect 14188 4082 14240 4088
rect 14108 3670 14136 4082
rect 14096 3664 14148 3670
rect 14096 3606 14148 3612
rect 14200 3194 14228 4082
rect 14188 3188 14240 3194
rect 14188 3130 14240 3136
rect 14292 2774 14320 10474
rect 14568 9518 14596 11562
rect 14556 9512 14608 9518
rect 14556 9454 14608 9460
rect 14372 9376 14424 9382
rect 14372 9318 14424 9324
rect 14384 8378 14412 9318
rect 14556 9172 14608 9178
rect 14556 9114 14608 9120
rect 14464 8968 14516 8974
rect 14464 8910 14516 8916
rect 14476 8634 14504 8910
rect 14464 8628 14516 8634
rect 14464 8570 14516 8576
rect 14384 8350 14504 8378
rect 14370 7304 14426 7313
rect 14370 7239 14426 7248
rect 14384 6934 14412 7239
rect 14372 6928 14424 6934
rect 14372 6870 14424 6876
rect 14370 4720 14426 4729
rect 14370 4655 14426 4664
rect 14384 4146 14412 4655
rect 14372 4140 14424 4146
rect 14372 4082 14424 4088
rect 14370 4040 14426 4049
rect 14370 3975 14426 3984
rect 14384 3534 14412 3975
rect 14372 3528 14424 3534
rect 14476 3505 14504 8350
rect 14372 3470 14424 3476
rect 14462 3496 14518 3505
rect 14462 3431 14518 3440
rect 14372 3120 14424 3126
rect 14372 3062 14424 3068
rect 14384 2938 14412 3062
rect 14568 3058 14596 9114
rect 14660 8498 14688 12038
rect 15016 11552 15068 11558
rect 15016 11494 15068 11500
rect 14740 10464 14792 10470
rect 14740 10406 14792 10412
rect 14648 8492 14700 8498
rect 14648 8434 14700 8440
rect 14660 8401 14688 8434
rect 14646 8392 14702 8401
rect 14646 8327 14702 8336
rect 14648 8016 14700 8022
rect 14648 7958 14700 7964
rect 14660 7818 14688 7958
rect 14648 7812 14700 7818
rect 14648 7754 14700 7760
rect 14648 6792 14700 6798
rect 14648 6734 14700 6740
rect 14556 3052 14608 3058
rect 14556 2994 14608 3000
rect 14384 2910 14596 2938
rect 14016 2746 14136 2774
rect 14108 1766 14136 2746
rect 14200 2746 14320 2774
rect 14096 1760 14148 1766
rect 14096 1702 14148 1708
rect 14200 800 14228 2746
rect 14568 2446 14596 2910
rect 14372 2440 14424 2446
rect 14372 2382 14424 2388
rect 14556 2440 14608 2446
rect 14556 2382 14608 2388
rect 14384 2038 14412 2382
rect 14556 2304 14608 2310
rect 14556 2246 14608 2252
rect 14372 2032 14424 2038
rect 14372 1974 14424 1980
rect 14568 1970 14596 2246
rect 14464 1964 14516 1970
rect 14464 1906 14516 1912
rect 14556 1964 14608 1970
rect 14556 1906 14608 1912
rect 14476 800 14504 1906
rect 14660 1766 14688 6734
rect 14648 1760 14700 1766
rect 14648 1702 14700 1708
rect 14752 800 14780 10406
rect 14924 9920 14976 9926
rect 14924 9862 14976 9868
rect 14936 9654 14964 9862
rect 14924 9648 14976 9654
rect 14924 9590 14976 9596
rect 14832 8968 14884 8974
rect 14832 8910 14884 8916
rect 14844 7954 14872 8910
rect 14924 8900 14976 8906
rect 14924 8842 14976 8848
rect 14936 8566 14964 8842
rect 14924 8560 14976 8566
rect 14924 8502 14976 8508
rect 14832 7948 14884 7954
rect 14832 7890 14884 7896
rect 14924 7336 14976 7342
rect 14924 7278 14976 7284
rect 14936 6866 14964 7278
rect 14924 6860 14976 6866
rect 14924 6802 14976 6808
rect 14832 6316 14884 6322
rect 14832 6258 14884 6264
rect 14844 5574 14872 6258
rect 14832 5568 14884 5574
rect 14832 5510 14884 5516
rect 14922 5536 14978 5545
rect 14922 5471 14978 5480
rect 14936 5302 14964 5471
rect 14924 5296 14976 5302
rect 14924 5238 14976 5244
rect 14830 4856 14886 4865
rect 14830 4791 14832 4800
rect 14884 4791 14886 4800
rect 14832 4762 14884 4768
rect 14832 4684 14884 4690
rect 14832 4626 14884 4632
rect 14844 4214 14872 4626
rect 14924 4616 14976 4622
rect 14924 4558 14976 4564
rect 14936 4214 14964 4558
rect 14832 4208 14884 4214
rect 14830 4176 14832 4185
rect 14924 4208 14976 4214
rect 14884 4176 14886 4185
rect 14924 4150 14976 4156
rect 14830 4111 14886 4120
rect 14922 4040 14978 4049
rect 14922 3975 14978 3984
rect 14936 3942 14964 3975
rect 14924 3936 14976 3942
rect 14924 3878 14976 3884
rect 14830 3632 14886 3641
rect 14830 3567 14886 3576
rect 14844 3534 14872 3567
rect 14832 3528 14884 3534
rect 14832 3470 14884 3476
rect 14830 3224 14886 3233
rect 14830 3159 14886 3168
rect 14844 1018 14872 3159
rect 14924 2984 14976 2990
rect 14924 2926 14976 2932
rect 14936 1834 14964 2926
rect 14924 1828 14976 1834
rect 14924 1770 14976 1776
rect 14832 1012 14884 1018
rect 14832 954 14884 960
rect 15028 800 15056 11494
rect 15120 11121 15148 12922
rect 15398 11996 15706 12005
rect 15398 11994 15404 11996
rect 15460 11994 15484 11996
rect 15540 11994 15564 11996
rect 15620 11994 15644 11996
rect 15700 11994 15706 11996
rect 15460 11942 15462 11994
rect 15642 11942 15644 11994
rect 15398 11940 15404 11942
rect 15460 11940 15484 11942
rect 15540 11940 15564 11942
rect 15620 11940 15644 11942
rect 15700 11940 15706 11942
rect 15398 11931 15706 11940
rect 15752 11552 15804 11558
rect 15752 11494 15804 11500
rect 15660 11280 15712 11286
rect 15660 11222 15712 11228
rect 15672 11121 15700 11222
rect 15106 11112 15162 11121
rect 15106 11047 15162 11056
rect 15658 11112 15714 11121
rect 15658 11047 15714 11056
rect 15398 10908 15706 10917
rect 15398 10906 15404 10908
rect 15460 10906 15484 10908
rect 15540 10906 15564 10908
rect 15620 10906 15644 10908
rect 15700 10906 15706 10908
rect 15460 10854 15462 10906
rect 15642 10854 15644 10906
rect 15398 10852 15404 10854
rect 15460 10852 15484 10854
rect 15540 10852 15564 10854
rect 15620 10852 15644 10854
rect 15700 10852 15706 10854
rect 15398 10843 15706 10852
rect 15292 10464 15344 10470
rect 15292 10406 15344 10412
rect 15200 9444 15252 9450
rect 15200 9386 15252 9392
rect 15212 8498 15240 9386
rect 15108 8492 15160 8498
rect 15108 8434 15160 8440
rect 15200 8492 15252 8498
rect 15200 8434 15252 8440
rect 15120 7857 15148 8434
rect 15106 7848 15162 7857
rect 15106 7783 15162 7792
rect 15200 7744 15252 7750
rect 15200 7686 15252 7692
rect 15106 7576 15162 7585
rect 15106 7511 15162 7520
rect 15120 6769 15148 7511
rect 15212 7313 15240 7686
rect 15198 7304 15254 7313
rect 15198 7239 15254 7248
rect 15106 6760 15162 6769
rect 15106 6695 15162 6704
rect 15108 6316 15160 6322
rect 15108 6258 15160 6264
rect 15120 5846 15148 6258
rect 15108 5840 15160 5846
rect 15108 5782 15160 5788
rect 15120 5234 15148 5782
rect 15108 5228 15160 5234
rect 15108 5170 15160 5176
rect 15200 5024 15252 5030
rect 15200 4966 15252 4972
rect 15108 4208 15160 4214
rect 15108 4150 15160 4156
rect 15120 3233 15148 4150
rect 15106 3224 15162 3233
rect 15106 3159 15162 3168
rect 15108 3120 15160 3126
rect 15108 3062 15160 3068
rect 15120 2938 15148 3062
rect 15212 3040 15240 4966
rect 15304 3534 15332 10406
rect 15474 10024 15530 10033
rect 15474 9959 15530 9968
rect 15488 9926 15516 9959
rect 15476 9920 15528 9926
rect 15476 9862 15528 9868
rect 15398 9820 15706 9829
rect 15398 9818 15404 9820
rect 15460 9818 15484 9820
rect 15540 9818 15564 9820
rect 15620 9818 15644 9820
rect 15700 9818 15706 9820
rect 15460 9766 15462 9818
rect 15642 9766 15644 9818
rect 15398 9764 15404 9766
rect 15460 9764 15484 9766
rect 15540 9764 15564 9766
rect 15620 9764 15644 9766
rect 15700 9764 15706 9766
rect 15398 9755 15706 9764
rect 15382 9616 15438 9625
rect 15382 9551 15438 9560
rect 15396 9518 15424 9551
rect 15384 9512 15436 9518
rect 15384 9454 15436 9460
rect 15476 9512 15528 9518
rect 15476 9454 15528 9460
rect 15488 8838 15516 9454
rect 15568 9104 15620 9110
rect 15568 9046 15620 9052
rect 15580 8838 15608 9046
rect 15476 8832 15528 8838
rect 15476 8774 15528 8780
rect 15568 8832 15620 8838
rect 15568 8774 15620 8780
rect 15398 8732 15706 8741
rect 15398 8730 15404 8732
rect 15460 8730 15484 8732
rect 15540 8730 15564 8732
rect 15620 8730 15644 8732
rect 15700 8730 15706 8732
rect 15460 8678 15462 8730
rect 15642 8678 15644 8730
rect 15398 8676 15404 8678
rect 15460 8676 15484 8678
rect 15540 8676 15564 8678
rect 15620 8676 15644 8678
rect 15700 8676 15706 8678
rect 15398 8667 15706 8676
rect 15398 7644 15706 7653
rect 15398 7642 15404 7644
rect 15460 7642 15484 7644
rect 15540 7642 15564 7644
rect 15620 7642 15644 7644
rect 15700 7642 15706 7644
rect 15460 7590 15462 7642
rect 15642 7590 15644 7642
rect 15398 7588 15404 7590
rect 15460 7588 15484 7590
rect 15540 7588 15564 7590
rect 15620 7588 15644 7590
rect 15700 7588 15706 7590
rect 15398 7579 15706 7588
rect 15384 7540 15436 7546
rect 15384 7482 15436 7488
rect 15396 7410 15424 7482
rect 15384 7404 15436 7410
rect 15384 7346 15436 7352
rect 15398 6556 15706 6565
rect 15398 6554 15404 6556
rect 15460 6554 15484 6556
rect 15540 6554 15564 6556
rect 15620 6554 15644 6556
rect 15700 6554 15706 6556
rect 15460 6502 15462 6554
rect 15642 6502 15644 6554
rect 15398 6500 15404 6502
rect 15460 6500 15484 6502
rect 15540 6500 15564 6502
rect 15620 6500 15644 6502
rect 15700 6500 15706 6502
rect 15398 6491 15706 6500
rect 15398 5468 15706 5477
rect 15398 5466 15404 5468
rect 15460 5466 15484 5468
rect 15540 5466 15564 5468
rect 15620 5466 15644 5468
rect 15700 5466 15706 5468
rect 15460 5414 15462 5466
rect 15642 5414 15644 5466
rect 15398 5412 15404 5414
rect 15460 5412 15484 5414
rect 15540 5412 15564 5414
rect 15620 5412 15644 5414
rect 15700 5412 15706 5414
rect 15398 5403 15706 5412
rect 15398 4380 15706 4389
rect 15398 4378 15404 4380
rect 15460 4378 15484 4380
rect 15540 4378 15564 4380
rect 15620 4378 15644 4380
rect 15700 4378 15706 4380
rect 15460 4326 15462 4378
rect 15642 4326 15644 4378
rect 15398 4324 15404 4326
rect 15460 4324 15484 4326
rect 15540 4324 15564 4326
rect 15620 4324 15644 4326
rect 15700 4324 15706 4326
rect 15398 4315 15706 4324
rect 15382 3768 15438 3777
rect 15382 3703 15384 3712
rect 15436 3703 15438 3712
rect 15384 3674 15436 3680
rect 15764 3618 15792 11494
rect 15856 11218 15884 13126
rect 16960 12782 16988 13194
rect 17776 13184 17828 13190
rect 17774 13152 17776 13161
rect 18052 13184 18104 13190
rect 17828 13152 17830 13161
rect 18052 13126 18104 13132
rect 17774 13087 17830 13096
rect 17224 12844 17276 12850
rect 17224 12786 17276 12792
rect 16948 12776 17000 12782
rect 16948 12718 17000 12724
rect 17236 12646 17264 12786
rect 16120 12640 16172 12646
rect 16120 12582 16172 12588
rect 17224 12640 17276 12646
rect 17224 12582 17276 12588
rect 16132 12481 16160 12582
rect 16118 12472 16174 12481
rect 16118 12407 16174 12416
rect 17236 12434 17264 12582
rect 17236 12406 17540 12434
rect 17224 12164 17276 12170
rect 17224 12106 17276 12112
rect 16580 12096 16632 12102
rect 16580 12038 16632 12044
rect 16948 12096 17000 12102
rect 16948 12038 17000 12044
rect 16592 11626 16620 12038
rect 16580 11620 16632 11626
rect 16580 11562 16632 11568
rect 16304 11552 16356 11558
rect 16304 11494 16356 11500
rect 16028 11280 16080 11286
rect 16028 11222 16080 11228
rect 15844 11212 15896 11218
rect 15844 11154 15896 11160
rect 15844 11076 15896 11082
rect 15844 11018 15896 11024
rect 15856 10674 15884 11018
rect 15844 10668 15896 10674
rect 15844 10610 15896 10616
rect 15856 5166 15884 10610
rect 15936 10464 15988 10470
rect 15936 10406 15988 10412
rect 15844 5160 15896 5166
rect 15844 5102 15896 5108
rect 15844 4480 15896 4486
rect 15844 4422 15896 4428
rect 15856 4146 15884 4422
rect 15844 4140 15896 4146
rect 15844 4082 15896 4088
rect 15856 3738 15884 4082
rect 15844 3732 15896 3738
rect 15844 3674 15896 3680
rect 15764 3590 15884 3618
rect 15292 3528 15344 3534
rect 15292 3470 15344 3476
rect 15752 3528 15804 3534
rect 15752 3470 15804 3476
rect 15398 3292 15706 3301
rect 15398 3290 15404 3292
rect 15460 3290 15484 3292
rect 15540 3290 15564 3292
rect 15620 3290 15644 3292
rect 15700 3290 15706 3292
rect 15460 3238 15462 3290
rect 15642 3238 15644 3290
rect 15398 3236 15404 3238
rect 15460 3236 15484 3238
rect 15540 3236 15564 3238
rect 15620 3236 15644 3238
rect 15700 3236 15706 3238
rect 15398 3227 15706 3236
rect 15292 3052 15344 3058
rect 15212 3012 15292 3040
rect 15292 2994 15344 3000
rect 15120 2910 15240 2938
rect 15212 1737 15240 2910
rect 15658 2816 15714 2825
rect 15658 2751 15714 2760
rect 15672 2582 15700 2751
rect 15660 2576 15712 2582
rect 15660 2518 15712 2524
rect 15292 2304 15344 2310
rect 15292 2246 15344 2252
rect 15304 2038 15332 2246
rect 15398 2204 15706 2213
rect 15398 2202 15404 2204
rect 15460 2202 15484 2204
rect 15540 2202 15564 2204
rect 15620 2202 15644 2204
rect 15700 2202 15706 2204
rect 15460 2150 15462 2202
rect 15642 2150 15644 2202
rect 15398 2148 15404 2150
rect 15460 2148 15484 2150
rect 15540 2148 15564 2150
rect 15620 2148 15644 2150
rect 15700 2148 15706 2150
rect 15398 2139 15706 2148
rect 15764 2088 15792 3470
rect 15580 2060 15792 2088
rect 15292 2032 15344 2038
rect 15292 1974 15344 1980
rect 15292 1828 15344 1834
rect 15292 1770 15344 1776
rect 15198 1728 15254 1737
rect 15198 1663 15254 1672
rect 15304 800 15332 1770
rect 15580 800 15608 2060
rect 15856 800 15884 3590
rect 15948 3126 15976 10406
rect 15936 3120 15988 3126
rect 15936 3062 15988 3068
rect 16040 3058 16068 11222
rect 16316 11150 16344 11494
rect 16304 11144 16356 11150
rect 16304 11086 16356 11092
rect 16212 10668 16264 10674
rect 16212 10610 16264 10616
rect 16120 10532 16172 10538
rect 16120 10474 16172 10480
rect 16028 3052 16080 3058
rect 16028 2994 16080 3000
rect 15934 2952 15990 2961
rect 15934 2887 15936 2896
rect 15988 2887 15990 2896
rect 15936 2858 15988 2864
rect 16028 2848 16080 2854
rect 15948 2796 16028 2802
rect 15948 2790 16080 2796
rect 15948 2774 16068 2790
rect 15948 800 15976 2774
rect 16028 2304 16080 2310
rect 16028 2246 16080 2252
rect 16040 1494 16068 2246
rect 16028 1488 16080 1494
rect 16028 1430 16080 1436
rect 16132 800 16160 10474
rect 16224 9654 16252 10610
rect 16212 9648 16264 9654
rect 16212 9590 16264 9596
rect 16212 8832 16264 8838
rect 16212 8774 16264 8780
rect 16224 8090 16252 8774
rect 16212 8084 16264 8090
rect 16212 8026 16264 8032
rect 16224 7410 16252 8026
rect 16212 7404 16264 7410
rect 16212 7346 16264 7352
rect 16316 7290 16344 11086
rect 16592 9466 16620 11562
rect 16856 11144 16908 11150
rect 16856 11086 16908 11092
rect 16500 9450 16620 9466
rect 16488 9444 16620 9450
rect 16540 9438 16620 9444
rect 16488 9386 16540 9392
rect 16408 9166 16620 9194
rect 16408 8974 16436 9166
rect 16488 9104 16540 9110
rect 16488 9046 16540 9052
rect 16396 8968 16448 8974
rect 16396 8910 16448 8916
rect 16396 8492 16448 8498
rect 16396 8434 16448 8440
rect 16408 7886 16436 8434
rect 16396 7880 16448 7886
rect 16396 7822 16448 7828
rect 16224 7262 16344 7290
rect 16224 2854 16252 7262
rect 16408 7206 16436 7822
rect 16304 7200 16356 7206
rect 16304 7142 16356 7148
rect 16396 7200 16448 7206
rect 16396 7142 16448 7148
rect 16316 7002 16344 7142
rect 16304 6996 16356 7002
rect 16304 6938 16356 6944
rect 16396 6928 16448 6934
rect 16396 6870 16448 6876
rect 16408 6633 16436 6870
rect 16500 6746 16528 9046
rect 16592 8090 16620 9166
rect 16672 9036 16724 9042
rect 16672 8978 16724 8984
rect 16684 8566 16712 8978
rect 16672 8560 16724 8566
rect 16672 8502 16724 8508
rect 16580 8084 16632 8090
rect 16580 8026 16632 8032
rect 16500 6730 16620 6746
rect 16500 6724 16632 6730
rect 16500 6718 16580 6724
rect 16580 6666 16632 6672
rect 16394 6624 16450 6633
rect 16394 6559 16450 6568
rect 16672 6248 16724 6254
rect 16672 6190 16724 6196
rect 16396 6112 16448 6118
rect 16396 6054 16448 6060
rect 16408 5710 16436 6054
rect 16684 5710 16712 6190
rect 16764 6112 16816 6118
rect 16764 6054 16816 6060
rect 16776 5914 16804 6054
rect 16764 5908 16816 5914
rect 16764 5850 16816 5856
rect 16396 5704 16448 5710
rect 16396 5646 16448 5652
rect 16488 5704 16540 5710
rect 16488 5646 16540 5652
rect 16672 5704 16724 5710
rect 16672 5646 16724 5652
rect 16500 5370 16528 5646
rect 16488 5364 16540 5370
rect 16488 5306 16540 5312
rect 16488 5160 16540 5166
rect 16488 5102 16540 5108
rect 16304 4140 16356 4146
rect 16304 4082 16356 4088
rect 16316 3534 16344 4082
rect 16396 4072 16448 4078
rect 16396 4014 16448 4020
rect 16304 3528 16356 3534
rect 16304 3470 16356 3476
rect 16408 3398 16436 4014
rect 16396 3392 16448 3398
rect 16302 3360 16358 3369
rect 16396 3334 16448 3340
rect 16302 3295 16358 3304
rect 16212 2848 16264 2854
rect 16212 2790 16264 2796
rect 16316 2774 16344 3295
rect 16316 2746 16436 2774
rect 16212 2576 16264 2582
rect 16212 2518 16264 2524
rect 16224 800 16252 2518
rect 16408 800 16436 2746
rect 16500 800 16528 5102
rect 16776 5030 16804 5850
rect 16764 5024 16816 5030
rect 16764 4966 16816 4972
rect 16776 4690 16804 4966
rect 16764 4684 16816 4690
rect 16764 4626 16816 4632
rect 16672 4548 16724 4554
rect 16672 4490 16724 4496
rect 16684 4078 16712 4490
rect 16762 4312 16818 4321
rect 16762 4247 16818 4256
rect 16776 4214 16804 4247
rect 16764 4208 16816 4214
rect 16764 4150 16816 4156
rect 16672 4072 16724 4078
rect 16672 4014 16724 4020
rect 16580 3936 16632 3942
rect 16868 3890 16896 11086
rect 16960 9518 16988 12038
rect 17236 11558 17264 12106
rect 17224 11552 17276 11558
rect 17224 11494 17276 11500
rect 16948 9512 17000 9518
rect 16948 9454 17000 9460
rect 16960 8430 16988 9454
rect 17132 9444 17184 9450
rect 17132 9386 17184 9392
rect 17040 8968 17092 8974
rect 17040 8910 17092 8916
rect 17052 8498 17080 8910
rect 17040 8492 17092 8498
rect 17040 8434 17092 8440
rect 16948 8424 17000 8430
rect 16948 8366 17000 8372
rect 16960 7886 16988 8366
rect 17144 7886 17172 9386
rect 17236 8566 17264 11494
rect 17316 10600 17368 10606
rect 17316 10542 17368 10548
rect 17328 10062 17356 10542
rect 17408 10464 17460 10470
rect 17408 10406 17460 10412
rect 17316 10056 17368 10062
rect 17316 9998 17368 10004
rect 17328 9654 17356 9998
rect 17316 9648 17368 9654
rect 17316 9590 17368 9596
rect 17420 9586 17448 10406
rect 17408 9580 17460 9586
rect 17408 9522 17460 9528
rect 17408 8968 17460 8974
rect 17408 8910 17460 8916
rect 17420 8634 17448 8910
rect 17408 8628 17460 8634
rect 17408 8570 17460 8576
rect 17224 8560 17276 8566
rect 17224 8502 17276 8508
rect 16948 7880 17000 7886
rect 16948 7822 17000 7828
rect 17132 7880 17184 7886
rect 17132 7822 17184 7828
rect 16948 7540 17000 7546
rect 16948 7482 17000 7488
rect 16960 6866 16988 7482
rect 17040 7404 17092 7410
rect 17040 7346 17092 7352
rect 16948 6860 17000 6866
rect 16948 6802 17000 6808
rect 16960 6322 16988 6802
rect 16948 6316 17000 6322
rect 16948 6258 17000 6264
rect 17052 5710 17080 7346
rect 17314 7032 17370 7041
rect 17314 6967 17370 6976
rect 17132 6792 17184 6798
rect 17132 6734 17184 6740
rect 17040 5704 17092 5710
rect 17040 5646 17092 5652
rect 17040 5568 17092 5574
rect 17144 5545 17172 6734
rect 17224 6112 17276 6118
rect 17224 6054 17276 6060
rect 17040 5510 17092 5516
rect 17130 5536 17186 5545
rect 16948 5364 17000 5370
rect 16948 5306 17000 5312
rect 16960 5098 16988 5306
rect 17052 5302 17080 5510
rect 17130 5471 17186 5480
rect 17040 5296 17092 5302
rect 17040 5238 17092 5244
rect 16948 5092 17000 5098
rect 16948 5034 17000 5040
rect 16946 4992 17002 5001
rect 16946 4927 17002 4936
rect 16580 3878 16632 3884
rect 16592 3534 16620 3878
rect 16684 3862 16896 3890
rect 16580 3528 16632 3534
rect 16580 3470 16632 3476
rect 16592 3058 16620 3470
rect 16580 3052 16632 3058
rect 16580 2994 16632 3000
rect 16684 800 16712 3862
rect 16762 3768 16818 3777
rect 16960 3754 16988 4927
rect 17236 4282 17264 6054
rect 17224 4276 17276 4282
rect 17224 4218 17276 4224
rect 17037 4140 17089 4146
rect 17037 4082 17089 4088
rect 16762 3703 16818 3712
rect 16868 3726 16988 3754
rect 17052 3738 17080 4082
rect 17040 3732 17092 3738
rect 16776 800 16804 3703
rect 16868 2553 16896 3726
rect 17040 3674 17092 3680
rect 17328 3618 17356 6967
rect 17408 6112 17460 6118
rect 17408 6054 17460 6060
rect 17512 6066 17540 12406
rect 17684 10668 17736 10674
rect 17684 10610 17736 10616
rect 17696 10266 17724 10610
rect 17684 10260 17736 10266
rect 17684 10202 17736 10208
rect 17776 10260 17828 10266
rect 17776 10202 17828 10208
rect 17788 9722 17816 10202
rect 17776 9716 17828 9722
rect 17776 9658 17828 9664
rect 17866 9616 17922 9625
rect 17866 9551 17922 9560
rect 17880 9217 17908 9551
rect 17590 9208 17646 9217
rect 17590 9143 17646 9152
rect 17866 9208 17922 9217
rect 17866 9143 17922 9152
rect 17604 6202 17632 9143
rect 17866 8936 17922 8945
rect 17866 8871 17922 8880
rect 17774 8528 17830 8537
rect 17774 8463 17830 8472
rect 17788 8430 17816 8463
rect 17776 8424 17828 8430
rect 17776 8366 17828 8372
rect 17684 8288 17736 8294
rect 17684 8230 17736 8236
rect 17696 8022 17724 8230
rect 17880 8090 17908 8871
rect 17868 8084 17920 8090
rect 17868 8026 17920 8032
rect 17684 8016 17736 8022
rect 17684 7958 17736 7964
rect 17960 7812 18012 7818
rect 17960 7754 18012 7760
rect 17684 7540 17736 7546
rect 17684 7482 17736 7488
rect 17696 6866 17724 7482
rect 17972 7410 18000 7754
rect 17960 7404 18012 7410
rect 17960 7346 18012 7352
rect 17684 6860 17736 6866
rect 17684 6802 17736 6808
rect 17868 6248 17920 6254
rect 17604 6174 17724 6202
rect 17868 6190 17920 6196
rect 17420 5370 17448 6054
rect 17512 6038 17632 6066
rect 17498 5944 17554 5953
rect 17498 5879 17500 5888
rect 17552 5879 17554 5888
rect 17500 5850 17552 5856
rect 17408 5364 17460 5370
rect 17408 5306 17460 5312
rect 17500 4820 17552 4826
rect 17500 4762 17552 4768
rect 17052 3590 17356 3618
rect 17408 3664 17460 3670
rect 17408 3606 17460 3612
rect 16948 3392 17000 3398
rect 16948 3334 17000 3340
rect 16960 3194 16988 3334
rect 16948 3188 17000 3194
rect 16948 3130 17000 3136
rect 17052 2774 17080 3590
rect 17222 3496 17278 3505
rect 17222 3431 17278 3440
rect 17316 3460 17368 3466
rect 17236 3398 17264 3431
rect 17316 3402 17368 3408
rect 17224 3392 17276 3398
rect 17224 3334 17276 3340
rect 17328 3058 17356 3402
rect 17316 3052 17368 3058
rect 17316 2994 17368 3000
rect 16960 2746 17080 2774
rect 16854 2544 16910 2553
rect 16854 2479 16910 2488
rect 16960 800 16988 2746
rect 17222 2544 17278 2553
rect 17222 2479 17278 2488
rect 17236 2446 17264 2479
rect 17224 2440 17276 2446
rect 17224 2382 17276 2388
rect 17132 1420 17184 1426
rect 17132 1362 17184 1368
rect 17144 800 17172 1362
rect 17420 800 17448 3606
rect 17512 3194 17540 4762
rect 17604 4729 17632 6038
rect 17590 4720 17646 4729
rect 17590 4655 17646 4664
rect 17604 4078 17632 4655
rect 17592 4072 17644 4078
rect 17592 4014 17644 4020
rect 17500 3188 17552 3194
rect 17500 3130 17552 3136
rect 17696 2774 17724 6174
rect 17880 6089 17908 6190
rect 17866 6080 17922 6089
rect 17922 6038 18000 6066
rect 17866 6015 17922 6024
rect 17880 5955 17908 6015
rect 17868 5772 17920 5778
rect 17868 5714 17920 5720
rect 17880 4758 17908 5714
rect 17972 5302 18000 6038
rect 17960 5296 18012 5302
rect 17960 5238 18012 5244
rect 17958 4856 18014 4865
rect 17958 4791 18014 4800
rect 17868 4752 17920 4758
rect 17868 4694 17920 4700
rect 17972 4146 18000 4791
rect 17960 4140 18012 4146
rect 17960 4082 18012 4088
rect 17960 3528 18012 3534
rect 17960 3470 18012 3476
rect 17972 3369 18000 3470
rect 17958 3360 18014 3369
rect 17958 3295 18014 3304
rect 18064 3058 18092 13126
rect 18236 12912 18288 12918
rect 18236 12854 18288 12860
rect 18248 12646 18276 12854
rect 19064 12776 19116 12782
rect 19064 12718 19116 12724
rect 18236 12640 18288 12646
rect 18234 12608 18236 12617
rect 18288 12608 18290 12617
rect 18234 12543 18290 12552
rect 18604 12096 18656 12102
rect 18602 12064 18604 12073
rect 18788 12096 18840 12102
rect 18656 12064 18658 12073
rect 18788 12038 18840 12044
rect 18602 11999 18658 12008
rect 18236 11552 18288 11558
rect 18236 11494 18288 11500
rect 18144 10056 18196 10062
rect 18144 9998 18196 10004
rect 18156 5250 18184 9998
rect 18248 9178 18276 11494
rect 18604 11144 18656 11150
rect 18604 11086 18656 11092
rect 18420 10464 18472 10470
rect 18420 10406 18472 10412
rect 18432 9926 18460 10406
rect 18512 10056 18564 10062
rect 18512 9998 18564 10004
rect 18420 9920 18472 9926
rect 18420 9862 18472 9868
rect 18432 9722 18460 9862
rect 18420 9716 18472 9722
rect 18420 9658 18472 9664
rect 18236 9172 18288 9178
rect 18236 9114 18288 9120
rect 18248 8430 18276 9114
rect 18236 8424 18288 8430
rect 18234 8392 18236 8401
rect 18288 8392 18290 8401
rect 18234 8327 18290 8336
rect 18420 7880 18472 7886
rect 18420 7822 18472 7828
rect 18432 7546 18460 7822
rect 18420 7540 18472 7546
rect 18420 7482 18472 7488
rect 18328 7404 18380 7410
rect 18328 7346 18380 7352
rect 18420 7404 18472 7410
rect 18420 7346 18472 7352
rect 18340 6769 18368 7346
rect 18432 7206 18460 7346
rect 18420 7200 18472 7206
rect 18420 7142 18472 7148
rect 18420 6996 18472 7002
rect 18420 6938 18472 6944
rect 18326 6760 18382 6769
rect 18326 6695 18382 6704
rect 18432 6662 18460 6938
rect 18236 6656 18288 6662
rect 18420 6656 18472 6662
rect 18236 6598 18288 6604
rect 18326 6624 18382 6633
rect 18248 5914 18276 6598
rect 18420 6598 18472 6604
rect 18326 6559 18382 6568
rect 18340 6390 18368 6559
rect 18328 6384 18380 6390
rect 18328 6326 18380 6332
rect 18236 5908 18288 5914
rect 18236 5850 18288 5856
rect 18236 5704 18288 5710
rect 18236 5646 18288 5652
rect 18248 5370 18276 5646
rect 18236 5364 18288 5370
rect 18236 5306 18288 5312
rect 18156 5222 18276 5250
rect 18142 4448 18198 4457
rect 18142 4383 18198 4392
rect 18156 4214 18184 4383
rect 18144 4208 18196 4214
rect 18142 4176 18144 4185
rect 18196 4176 18198 4185
rect 18142 4111 18198 4120
rect 18052 3052 18104 3058
rect 18052 2994 18104 3000
rect 17776 2916 17828 2922
rect 17776 2858 17828 2864
rect 17604 2746 17724 2774
rect 17604 2514 17632 2746
rect 17682 2680 17738 2689
rect 17788 2650 17816 2858
rect 17960 2848 18012 2854
rect 17960 2790 18012 2796
rect 17682 2615 17738 2624
rect 17776 2644 17828 2650
rect 17592 2508 17644 2514
rect 17592 2450 17644 2456
rect 17696 2446 17724 2615
rect 17776 2586 17828 2592
rect 17684 2440 17736 2446
rect 17684 2382 17736 2388
rect 17684 2304 17736 2310
rect 17684 2246 17736 2252
rect 17696 800 17724 2246
rect 17972 800 18000 2790
rect 18064 2774 18092 2994
rect 18064 2746 18184 2774
rect 18156 1698 18184 2746
rect 18144 1692 18196 1698
rect 18144 1634 18196 1640
rect 18248 800 18276 5222
rect 18340 4554 18368 6326
rect 18432 5710 18460 6598
rect 18420 5704 18472 5710
rect 18420 5646 18472 5652
rect 18328 4548 18380 4554
rect 18328 4490 18380 4496
rect 18420 4480 18472 4486
rect 18420 4422 18472 4428
rect 18432 3670 18460 4422
rect 18420 3664 18472 3670
rect 18326 3632 18382 3641
rect 18420 3606 18472 3612
rect 18326 3567 18382 3576
rect 18340 3534 18368 3567
rect 18328 3528 18380 3534
rect 18328 3470 18380 3476
rect 18524 800 18552 9998
rect 18616 6304 18644 11086
rect 18800 11082 18828 12038
rect 18788 11076 18840 11082
rect 18788 11018 18840 11024
rect 18800 8090 18828 11018
rect 18972 9512 19024 9518
rect 18972 9454 19024 9460
rect 18984 9353 19012 9454
rect 18970 9344 19026 9353
rect 18970 9279 19026 9288
rect 18788 8084 18840 8090
rect 18788 8026 18840 8032
rect 18800 6390 18828 8026
rect 18984 7342 19012 9279
rect 18972 7336 19024 7342
rect 18972 7278 19024 7284
rect 19076 7290 19104 12718
rect 19248 12232 19300 12238
rect 19248 12174 19300 12180
rect 19260 11558 19288 12174
rect 19720 12102 19748 13194
rect 20076 12708 20128 12714
rect 20076 12650 20128 12656
rect 19984 12640 20036 12646
rect 19984 12582 20036 12588
rect 19708 12096 19760 12102
rect 19708 12038 19760 12044
rect 19248 11552 19300 11558
rect 19248 11494 19300 11500
rect 19800 11552 19852 11558
rect 19800 11494 19852 11500
rect 19260 11150 19288 11494
rect 19248 11144 19300 11150
rect 19248 11086 19300 11092
rect 19524 11076 19576 11082
rect 19524 11018 19576 11024
rect 19340 9716 19392 9722
rect 19340 9658 19392 9664
rect 19248 8288 19300 8294
rect 19248 8230 19300 8236
rect 19260 7886 19288 8230
rect 19248 7880 19300 7886
rect 19248 7822 19300 7828
rect 19248 7472 19300 7478
rect 19246 7440 19248 7449
rect 19300 7440 19302 7449
rect 19246 7375 19302 7384
rect 19076 7262 19288 7290
rect 19064 7200 19116 7206
rect 19064 7142 19116 7148
rect 19156 7200 19208 7206
rect 19156 7142 19208 7148
rect 19076 6390 19104 7142
rect 18788 6384 18840 6390
rect 18788 6326 18840 6332
rect 19064 6384 19116 6390
rect 19064 6326 19116 6332
rect 18696 6316 18748 6322
rect 18616 6276 18696 6304
rect 18616 6118 18644 6276
rect 18696 6258 18748 6264
rect 18694 6216 18750 6225
rect 18694 6151 18750 6160
rect 18604 6112 18656 6118
rect 18604 6054 18656 6060
rect 18708 5710 18736 6151
rect 18788 5908 18840 5914
rect 18788 5850 18840 5856
rect 18696 5704 18748 5710
rect 18696 5646 18748 5652
rect 18694 5128 18750 5137
rect 18694 5063 18750 5072
rect 18708 4865 18736 5063
rect 18694 4856 18750 4865
rect 18694 4791 18750 4800
rect 18708 2446 18736 4791
rect 18800 3126 18828 5850
rect 18880 5636 18932 5642
rect 18880 5578 18932 5584
rect 18892 5302 18920 5578
rect 18880 5296 18932 5302
rect 18880 5238 18932 5244
rect 19168 5137 19196 7142
rect 19154 5128 19210 5137
rect 19154 5063 19210 5072
rect 19062 4176 19118 4185
rect 19062 4111 19118 4120
rect 19156 4140 19208 4146
rect 18880 3936 18932 3942
rect 18880 3878 18932 3884
rect 18788 3120 18840 3126
rect 18788 3062 18840 3068
rect 18696 2440 18748 2446
rect 18696 2382 18748 2388
rect 18786 1864 18842 1873
rect 18786 1799 18842 1808
rect 18800 800 18828 1799
rect 18892 1086 18920 3878
rect 19076 3126 19104 4111
rect 19156 4082 19208 4088
rect 19168 4049 19196 4082
rect 19154 4040 19210 4049
rect 19154 3975 19210 3984
rect 19260 3534 19288 7262
rect 19352 6458 19380 9658
rect 19536 8809 19564 11018
rect 19708 9920 19760 9926
rect 19708 9862 19760 9868
rect 19720 9722 19748 9862
rect 19708 9716 19760 9722
rect 19708 9658 19760 9664
rect 19616 9376 19668 9382
rect 19616 9318 19668 9324
rect 19628 8974 19656 9318
rect 19616 8968 19668 8974
rect 19616 8910 19668 8916
rect 19708 8968 19760 8974
rect 19708 8910 19760 8916
rect 19522 8800 19578 8809
rect 19522 8735 19578 8744
rect 19432 8492 19484 8498
rect 19432 8434 19484 8440
rect 19444 7834 19472 8434
rect 19536 8022 19564 8735
rect 19720 8430 19748 8910
rect 19708 8424 19760 8430
rect 19708 8366 19760 8372
rect 19812 8090 19840 11494
rect 19892 9376 19944 9382
rect 19892 9318 19944 9324
rect 19904 8498 19932 9318
rect 19892 8492 19944 8498
rect 19892 8434 19944 8440
rect 19800 8084 19852 8090
rect 19800 8026 19852 8032
rect 19524 8016 19576 8022
rect 19524 7958 19576 7964
rect 19708 7948 19760 7954
rect 19708 7890 19760 7896
rect 19720 7834 19748 7890
rect 19444 7806 19748 7834
rect 19444 7410 19472 7806
rect 19524 7744 19576 7750
rect 19524 7686 19576 7692
rect 19432 7404 19484 7410
rect 19432 7346 19484 7352
rect 19430 6896 19486 6905
rect 19430 6831 19486 6840
rect 19340 6452 19392 6458
rect 19340 6394 19392 6400
rect 19444 5642 19472 6831
rect 19536 6798 19564 7686
rect 19720 7410 19748 7806
rect 19616 7404 19668 7410
rect 19616 7346 19668 7352
rect 19708 7404 19760 7410
rect 19708 7346 19760 7352
rect 19628 7290 19656 7346
rect 19812 7290 19840 8026
rect 19996 7698 20024 12582
rect 20088 12170 20116 12650
rect 20168 12368 20220 12374
rect 20168 12310 20220 12316
rect 20076 12164 20128 12170
rect 20076 12106 20128 12112
rect 20088 11898 20116 12106
rect 20076 11892 20128 11898
rect 20076 11834 20128 11840
rect 20180 11286 20208 12310
rect 20272 11558 20300 13874
rect 25412 13864 25464 13870
rect 25412 13806 25464 13812
rect 22622 13628 22930 13637
rect 22622 13626 22628 13628
rect 22684 13626 22708 13628
rect 22764 13626 22788 13628
rect 22844 13626 22868 13628
rect 22924 13626 22930 13628
rect 22684 13574 22686 13626
rect 22866 13574 22868 13626
rect 22622 13572 22628 13574
rect 22684 13572 22708 13574
rect 22764 13572 22788 13574
rect 22844 13572 22868 13574
rect 22924 13572 22930 13574
rect 22622 13563 22930 13572
rect 22284 13320 22336 13326
rect 22284 13262 22336 13268
rect 21916 12912 21968 12918
rect 21916 12854 21968 12860
rect 20720 12640 20772 12646
rect 20720 12582 20772 12588
rect 20732 12434 20760 12582
rect 20364 12406 20760 12434
rect 20260 11552 20312 11558
rect 20260 11494 20312 11500
rect 20168 11280 20220 11286
rect 20168 11222 20220 11228
rect 20180 10606 20208 11222
rect 20168 10600 20220 10606
rect 20168 10542 20220 10548
rect 20076 9580 20128 9586
rect 20076 9522 20128 9528
rect 20088 9110 20116 9522
rect 20076 9104 20128 9110
rect 20076 9046 20128 9052
rect 20076 8900 20128 8906
rect 20076 8842 20128 8848
rect 20088 8430 20116 8842
rect 20076 8424 20128 8430
rect 20076 8366 20128 8372
rect 20180 7886 20208 10542
rect 20260 10532 20312 10538
rect 20260 10474 20312 10480
rect 20272 9382 20300 10474
rect 20260 9376 20312 9382
rect 20260 9318 20312 9324
rect 20272 9042 20300 9318
rect 20260 9036 20312 9042
rect 20260 8978 20312 8984
rect 20258 8664 20314 8673
rect 20258 8599 20314 8608
rect 20272 8566 20300 8599
rect 20260 8560 20312 8566
rect 20260 8502 20312 8508
rect 20168 7880 20220 7886
rect 20168 7822 20220 7828
rect 20260 7812 20312 7818
rect 20260 7754 20312 7760
rect 20166 7712 20222 7721
rect 19996 7670 20166 7698
rect 20166 7647 20222 7656
rect 19628 7262 19840 7290
rect 19616 7200 19668 7206
rect 19616 7142 19668 7148
rect 19524 6792 19576 6798
rect 19524 6734 19576 6740
rect 19628 6322 19656 7142
rect 19616 6316 19668 6322
rect 19616 6258 19668 6264
rect 19616 5704 19668 5710
rect 19616 5646 19668 5652
rect 19432 5636 19484 5642
rect 19432 5578 19484 5584
rect 19524 5568 19576 5574
rect 19524 5510 19576 5516
rect 19338 5400 19394 5409
rect 19338 5335 19394 5344
rect 19352 5030 19380 5335
rect 19536 5302 19564 5510
rect 19524 5296 19576 5302
rect 19524 5238 19576 5244
rect 19524 5160 19576 5166
rect 19524 5102 19576 5108
rect 19340 5024 19392 5030
rect 19338 4992 19340 5001
rect 19392 4992 19394 5001
rect 19338 4927 19394 4936
rect 19536 4622 19564 5102
rect 19524 4616 19576 4622
rect 19524 4558 19576 4564
rect 19432 4548 19484 4554
rect 19432 4490 19484 4496
rect 19444 4282 19472 4490
rect 19432 4276 19484 4282
rect 19432 4218 19484 4224
rect 19248 3528 19300 3534
rect 19248 3470 19300 3476
rect 19260 3233 19288 3470
rect 19246 3224 19302 3233
rect 19246 3159 19302 3168
rect 19064 3120 19116 3126
rect 19064 3062 19116 3068
rect 19062 2952 19118 2961
rect 19062 2887 19118 2896
rect 18880 1080 18932 1086
rect 18880 1022 18932 1028
rect 19076 800 19104 2887
rect 19260 1630 19288 3159
rect 19536 3126 19564 4558
rect 19524 3120 19576 3126
rect 19524 3062 19576 3068
rect 19340 2984 19392 2990
rect 19628 2961 19656 5646
rect 19340 2926 19392 2932
rect 19614 2952 19670 2961
rect 19248 1624 19300 1630
rect 19248 1566 19300 1572
rect 19352 800 19380 2926
rect 19614 2887 19670 2896
rect 19812 2553 19840 7262
rect 20076 6724 20128 6730
rect 20076 6666 20128 6672
rect 19892 3936 19944 3942
rect 19892 3878 19944 3884
rect 19904 3602 19932 3878
rect 19892 3596 19944 3602
rect 19892 3538 19944 3544
rect 19892 3392 19944 3398
rect 19892 3334 19944 3340
rect 19798 2544 19854 2553
rect 19798 2479 19854 2488
rect 19524 2304 19576 2310
rect 19524 2246 19576 2252
rect 19536 1834 19564 2246
rect 19616 1964 19668 1970
rect 19616 1906 19668 1912
rect 19524 1828 19576 1834
rect 19524 1770 19576 1776
rect 19628 800 19656 1906
rect 19904 800 19932 3334
rect 20088 2106 20116 6666
rect 20180 4486 20208 7647
rect 20272 6866 20300 7754
rect 20260 6860 20312 6866
rect 20260 6802 20312 6808
rect 20272 6322 20300 6802
rect 20260 6316 20312 6322
rect 20260 6258 20312 6264
rect 20168 4480 20220 4486
rect 20168 4422 20220 4428
rect 20364 2774 20392 12406
rect 20536 12232 20588 12238
rect 20536 12174 20588 12180
rect 20444 10464 20496 10470
rect 20444 10406 20496 10412
rect 20456 10062 20484 10406
rect 20444 10056 20496 10062
rect 20444 9998 20496 10004
rect 20444 8968 20496 8974
rect 20444 8910 20496 8916
rect 20456 8294 20484 8910
rect 20444 8288 20496 8294
rect 20444 8230 20496 8236
rect 20272 2746 20392 2774
rect 20272 2446 20300 2746
rect 20548 2446 20576 12174
rect 20628 12096 20680 12102
rect 20628 12038 20680 12044
rect 20640 4690 20668 12038
rect 21928 11830 21956 12854
rect 22100 12844 22152 12850
rect 22100 12786 22152 12792
rect 21916 11824 21968 11830
rect 21916 11766 21968 11772
rect 20996 11688 21048 11694
rect 20996 11630 21048 11636
rect 21008 11218 21036 11630
rect 22112 11558 22140 12786
rect 22296 12102 22324 13262
rect 25044 12912 25096 12918
rect 25044 12854 25096 12860
rect 23664 12776 23716 12782
rect 23664 12718 23716 12724
rect 23480 12640 23532 12646
rect 23480 12582 23532 12588
rect 22622 12540 22930 12549
rect 22622 12538 22628 12540
rect 22684 12538 22708 12540
rect 22764 12538 22788 12540
rect 22844 12538 22868 12540
rect 22924 12538 22930 12540
rect 22684 12486 22686 12538
rect 22866 12486 22868 12538
rect 22622 12484 22628 12486
rect 22684 12484 22708 12486
rect 22764 12484 22788 12486
rect 22844 12484 22868 12486
rect 22924 12484 22930 12486
rect 22622 12475 22930 12484
rect 23492 12481 23520 12582
rect 23478 12472 23534 12481
rect 23478 12407 23534 12416
rect 22468 12232 22520 12238
rect 22468 12174 22520 12180
rect 22284 12096 22336 12102
rect 22282 12064 22284 12073
rect 22336 12064 22338 12073
rect 22282 11999 22338 12008
rect 22480 11898 22508 12174
rect 22468 11892 22520 11898
rect 22468 11834 22520 11840
rect 23112 11892 23164 11898
rect 23112 11834 23164 11840
rect 21732 11552 21784 11558
rect 22100 11552 22152 11558
rect 21732 11494 21784 11500
rect 22098 11520 22100 11529
rect 22152 11520 22154 11529
rect 21548 11280 21600 11286
rect 21548 11222 21600 11228
rect 20996 11212 21048 11218
rect 20996 11154 21048 11160
rect 20904 10124 20956 10130
rect 20904 10066 20956 10072
rect 20916 9586 20944 10066
rect 20904 9580 20956 9586
rect 20904 9522 20956 9528
rect 20720 9172 20772 9178
rect 20720 9114 20772 9120
rect 20732 8906 20760 9114
rect 20720 8900 20772 8906
rect 20720 8842 20772 8848
rect 21008 8242 21036 11154
rect 21560 11082 21588 11222
rect 21456 11076 21508 11082
rect 21456 11018 21508 11024
rect 21548 11076 21600 11082
rect 21548 11018 21600 11024
rect 21086 8936 21142 8945
rect 21086 8871 21142 8880
rect 20916 8214 21036 8242
rect 20916 7886 20944 8214
rect 21100 8090 21128 8871
rect 21180 8832 21232 8838
rect 21180 8774 21232 8780
rect 21272 8832 21324 8838
rect 21272 8774 21324 8780
rect 21088 8084 21140 8090
rect 21088 8026 21140 8032
rect 20904 7880 20956 7886
rect 20904 7822 20956 7828
rect 20916 5692 20944 7822
rect 21192 7818 21220 8774
rect 21284 8634 21312 8774
rect 21272 8628 21324 8634
rect 21272 8570 21324 8576
rect 21270 8392 21326 8401
rect 21270 8327 21326 8336
rect 21284 8294 21312 8327
rect 21272 8288 21324 8294
rect 21272 8230 21324 8236
rect 21284 7886 21312 8230
rect 21468 7993 21496 11018
rect 21640 8968 21692 8974
rect 21640 8910 21692 8916
rect 21652 8634 21680 8910
rect 21640 8628 21692 8634
rect 21640 8570 21692 8576
rect 21454 7984 21510 7993
rect 21454 7919 21510 7928
rect 21272 7880 21324 7886
rect 21272 7822 21324 7828
rect 21180 7812 21232 7818
rect 21180 7754 21232 7760
rect 21468 7410 21496 7919
rect 21640 7744 21692 7750
rect 21640 7686 21692 7692
rect 21456 7404 21508 7410
rect 21456 7346 21508 7352
rect 21652 6798 21680 7686
rect 21640 6792 21692 6798
rect 21546 6760 21602 6769
rect 21640 6734 21692 6740
rect 21546 6695 21602 6704
rect 20996 6180 21048 6186
rect 20996 6122 21048 6128
rect 21008 5846 21036 6122
rect 20996 5840 21048 5846
rect 20996 5782 21048 5788
rect 21088 5704 21140 5710
rect 20916 5664 21036 5692
rect 20904 5024 20956 5030
rect 20904 4966 20956 4972
rect 20720 4752 20772 4758
rect 20720 4694 20772 4700
rect 20628 4684 20680 4690
rect 20628 4626 20680 4632
rect 20732 4146 20760 4694
rect 20720 4140 20772 4146
rect 20720 4082 20772 4088
rect 20916 2774 20944 4966
rect 20824 2746 20944 2774
rect 21008 2774 21036 5664
rect 21088 5646 21140 5652
rect 21272 5704 21324 5710
rect 21272 5646 21324 5652
rect 21100 3670 21128 5646
rect 21180 5364 21232 5370
rect 21180 5306 21232 5312
rect 21088 3664 21140 3670
rect 21088 3606 21140 3612
rect 21008 2746 21128 2774
rect 20824 2530 20852 2746
rect 20732 2502 20852 2530
rect 20260 2440 20312 2446
rect 20260 2382 20312 2388
rect 20536 2440 20588 2446
rect 20536 2382 20588 2388
rect 20076 2100 20128 2106
rect 20076 2042 20128 2048
rect 20168 1488 20220 1494
rect 20168 1430 20220 1436
rect 20180 800 20208 1430
rect 20272 1290 20300 2382
rect 20444 2032 20496 2038
rect 20444 1974 20496 1980
rect 20260 1284 20312 1290
rect 20260 1226 20312 1232
rect 20456 800 20484 1974
rect 20548 1358 20576 2382
rect 20536 1352 20588 1358
rect 20536 1294 20588 1300
rect 20732 800 20760 2502
rect 20904 2372 20956 2378
rect 20904 2314 20956 2320
rect 20916 1170 20944 2314
rect 21100 2106 21128 2746
rect 21192 2446 21220 5306
rect 21284 4321 21312 5646
rect 21456 5296 21508 5302
rect 21456 5238 21508 5244
rect 21468 4826 21496 5238
rect 21456 4820 21508 4826
rect 21456 4762 21508 4768
rect 21468 4622 21496 4762
rect 21364 4616 21416 4622
rect 21364 4558 21416 4564
rect 21456 4616 21508 4622
rect 21456 4558 21508 4564
rect 21270 4312 21326 4321
rect 21376 4282 21404 4558
rect 21270 4247 21326 4256
rect 21364 4276 21416 4282
rect 21364 4218 21416 4224
rect 21376 3602 21404 4218
rect 21364 3596 21416 3602
rect 21364 3538 21416 3544
rect 21560 2854 21588 6695
rect 21640 6384 21692 6390
rect 21640 6326 21692 6332
rect 21652 5778 21680 6326
rect 21640 5772 21692 5778
rect 21640 5714 21692 5720
rect 21744 5234 21772 11494
rect 22098 11455 22154 11464
rect 22622 11452 22930 11461
rect 22622 11450 22628 11452
rect 22684 11450 22708 11452
rect 22764 11450 22788 11452
rect 22844 11450 22868 11452
rect 22924 11450 22930 11452
rect 22684 11398 22686 11450
rect 22866 11398 22868 11450
rect 22622 11396 22628 11398
rect 22684 11396 22708 11398
rect 22764 11396 22788 11398
rect 22844 11396 22868 11398
rect 22924 11396 22930 11398
rect 22622 11387 22930 11396
rect 22468 11348 22520 11354
rect 22468 11290 22520 11296
rect 22100 11280 22152 11286
rect 22100 11222 22152 11228
rect 22112 11150 22140 11222
rect 22100 11144 22152 11150
rect 22100 11086 22152 11092
rect 22192 11144 22244 11150
rect 22192 11086 22244 11092
rect 22100 10464 22152 10470
rect 22100 10406 22152 10412
rect 21916 9920 21968 9926
rect 21916 9862 21968 9868
rect 22008 9920 22060 9926
rect 22008 9862 22060 9868
rect 21928 9178 21956 9862
rect 22020 9722 22048 9862
rect 22008 9716 22060 9722
rect 22008 9658 22060 9664
rect 22112 9518 22140 10406
rect 22100 9512 22152 9518
rect 22020 9472 22100 9500
rect 21916 9172 21968 9178
rect 21916 9114 21968 9120
rect 21824 9104 21876 9110
rect 21824 9046 21876 9052
rect 21836 8906 21864 9046
rect 21824 8900 21876 8906
rect 21824 8842 21876 8848
rect 22020 8362 22048 9472
rect 22100 9454 22152 9460
rect 22100 8560 22152 8566
rect 22098 8528 22100 8537
rect 22152 8528 22154 8537
rect 22098 8463 22154 8472
rect 22204 8480 22232 11086
rect 22480 11082 22508 11290
rect 22468 11076 22520 11082
rect 22468 11018 22520 11024
rect 22376 10668 22428 10674
rect 22376 10610 22428 10616
rect 22284 10056 22336 10062
rect 22284 9998 22336 10004
rect 22296 9382 22324 9998
rect 22388 9722 22416 10610
rect 22376 9716 22428 9722
rect 22376 9658 22428 9664
rect 22480 9518 22508 11018
rect 23020 10464 23072 10470
rect 23020 10406 23072 10412
rect 22622 10364 22930 10373
rect 22622 10362 22628 10364
rect 22684 10362 22708 10364
rect 22764 10362 22788 10364
rect 22844 10362 22868 10364
rect 22924 10362 22930 10364
rect 22684 10310 22686 10362
rect 22866 10310 22868 10362
rect 22622 10308 22628 10310
rect 22684 10308 22708 10310
rect 22764 10308 22788 10310
rect 22844 10308 22868 10310
rect 22924 10308 22930 10310
rect 22622 10299 22930 10308
rect 22560 10124 22612 10130
rect 22560 10066 22612 10072
rect 22572 9722 22600 10066
rect 23032 10062 23060 10406
rect 23020 10056 23072 10062
rect 23020 9998 23072 10004
rect 22560 9716 22612 9722
rect 22560 9658 22612 9664
rect 22468 9512 22520 9518
rect 22468 9454 22520 9460
rect 23020 9444 23072 9450
rect 23020 9386 23072 9392
rect 22284 9376 22336 9382
rect 22284 9318 22336 9324
rect 22296 9042 22324 9318
rect 22622 9276 22930 9285
rect 22622 9274 22628 9276
rect 22684 9274 22708 9276
rect 22764 9274 22788 9276
rect 22844 9274 22868 9276
rect 22924 9274 22930 9276
rect 22684 9222 22686 9274
rect 22866 9222 22868 9274
rect 22622 9220 22628 9222
rect 22684 9220 22708 9222
rect 22764 9220 22788 9222
rect 22844 9220 22868 9222
rect 22924 9220 22930 9222
rect 22622 9211 22930 9220
rect 22284 9036 22336 9042
rect 22284 8978 22336 8984
rect 22284 8492 22336 8498
rect 22204 8452 22284 8480
rect 22284 8434 22336 8440
rect 21916 8356 21968 8362
rect 21916 8298 21968 8304
rect 22008 8356 22060 8362
rect 22008 8298 22060 8304
rect 21824 7336 21876 7342
rect 21824 7278 21876 7284
rect 21836 7002 21864 7278
rect 21928 7206 21956 8298
rect 22296 8265 22324 8434
rect 22282 8256 22338 8265
rect 22282 8191 22338 8200
rect 22622 8188 22930 8197
rect 22622 8186 22628 8188
rect 22684 8186 22708 8188
rect 22764 8186 22788 8188
rect 22844 8186 22868 8188
rect 22924 8186 22930 8188
rect 22684 8134 22686 8186
rect 22866 8134 22868 8186
rect 22622 8132 22628 8134
rect 22684 8132 22708 8134
rect 22764 8132 22788 8134
rect 22844 8132 22868 8134
rect 22924 8132 22930 8134
rect 22622 8123 22930 8132
rect 23032 8090 23060 9386
rect 23020 8084 23072 8090
rect 23020 8026 23072 8032
rect 23020 7948 23072 7954
rect 23020 7890 23072 7896
rect 22376 7812 22428 7818
rect 22376 7754 22428 7760
rect 22006 7576 22062 7585
rect 22006 7511 22062 7520
rect 21916 7200 21968 7206
rect 21916 7142 21968 7148
rect 21824 6996 21876 7002
rect 21824 6938 21876 6944
rect 22020 6440 22048 7511
rect 22284 7268 22336 7274
rect 22284 7210 22336 7216
rect 22190 6896 22246 6905
rect 22296 6866 22324 7210
rect 22190 6831 22246 6840
rect 22284 6860 22336 6866
rect 22100 6656 22152 6662
rect 22100 6598 22152 6604
rect 21928 6412 22048 6440
rect 21732 5228 21784 5234
rect 21732 5170 21784 5176
rect 21640 5160 21692 5166
rect 21640 5102 21692 5108
rect 21652 4706 21680 5102
rect 21744 4865 21772 5170
rect 21730 4856 21786 4865
rect 21730 4791 21786 4800
rect 21652 4678 21772 4706
rect 21640 4616 21692 4622
rect 21640 4558 21692 4564
rect 21652 3942 21680 4558
rect 21744 4146 21772 4678
rect 21732 4140 21784 4146
rect 21732 4082 21784 4088
rect 21640 3936 21692 3942
rect 21640 3878 21692 3884
rect 21744 3398 21772 4082
rect 21732 3392 21784 3398
rect 21732 3334 21784 3340
rect 21928 3058 21956 6412
rect 22008 6316 22060 6322
rect 22008 6258 22060 6264
rect 22020 5914 22048 6258
rect 22112 6118 22140 6598
rect 22204 6322 22232 6831
rect 22284 6802 22336 6808
rect 22192 6316 22244 6322
rect 22192 6258 22244 6264
rect 22100 6112 22152 6118
rect 22100 6054 22152 6060
rect 22008 5908 22060 5914
rect 22008 5850 22060 5856
rect 22192 5568 22244 5574
rect 22192 5510 22244 5516
rect 22100 3528 22152 3534
rect 22100 3470 22152 3476
rect 22112 3126 22140 3470
rect 22204 3194 22232 5510
rect 22388 5370 22416 7754
rect 22622 7100 22930 7109
rect 22622 7098 22628 7100
rect 22684 7098 22708 7100
rect 22764 7098 22788 7100
rect 22844 7098 22868 7100
rect 22924 7098 22930 7100
rect 22684 7046 22686 7098
rect 22866 7046 22868 7098
rect 22622 7044 22628 7046
rect 22684 7044 22708 7046
rect 22764 7044 22788 7046
rect 22844 7044 22868 7046
rect 22924 7044 22930 7046
rect 22622 7035 22930 7044
rect 22560 6792 22612 6798
rect 22560 6734 22612 6740
rect 22572 6458 22600 6734
rect 22560 6452 22612 6458
rect 22560 6394 22612 6400
rect 22468 6112 22520 6118
rect 22468 6054 22520 6060
rect 22480 5710 22508 6054
rect 22622 6012 22930 6021
rect 22622 6010 22628 6012
rect 22684 6010 22708 6012
rect 22764 6010 22788 6012
rect 22844 6010 22868 6012
rect 22924 6010 22930 6012
rect 22684 5958 22686 6010
rect 22866 5958 22868 6010
rect 22622 5956 22628 5958
rect 22684 5956 22708 5958
rect 22764 5956 22788 5958
rect 22844 5956 22868 5958
rect 22924 5956 22930 5958
rect 22622 5947 22930 5956
rect 22468 5704 22520 5710
rect 22468 5646 22520 5652
rect 22376 5364 22428 5370
rect 22376 5306 22428 5312
rect 22284 5228 22336 5234
rect 22284 5170 22336 5176
rect 22296 4690 22324 5170
rect 22622 4924 22930 4933
rect 22622 4922 22628 4924
rect 22684 4922 22708 4924
rect 22764 4922 22788 4924
rect 22844 4922 22868 4924
rect 22924 4922 22930 4924
rect 22684 4870 22686 4922
rect 22866 4870 22868 4922
rect 22622 4868 22628 4870
rect 22684 4868 22708 4870
rect 22764 4868 22788 4870
rect 22844 4868 22868 4870
rect 22924 4868 22930 4870
rect 22622 4859 22930 4868
rect 22652 4820 22704 4826
rect 22652 4762 22704 4768
rect 22558 4720 22614 4729
rect 22284 4684 22336 4690
rect 22664 4690 22692 4762
rect 22558 4655 22614 4664
rect 22652 4684 22704 4690
rect 22284 4626 22336 4632
rect 22572 4622 22600 4655
rect 22652 4626 22704 4632
rect 22560 4616 22612 4622
rect 22480 4576 22560 4604
rect 22284 4480 22336 4486
rect 22284 4422 22336 4428
rect 22296 4146 22324 4422
rect 22284 4140 22336 4146
rect 22284 4082 22336 4088
rect 22376 4072 22428 4078
rect 22376 4014 22428 4020
rect 22388 3738 22416 4014
rect 22480 3738 22508 4576
rect 22560 4558 22612 4564
rect 22560 4480 22612 4486
rect 22652 4480 22704 4486
rect 22612 4440 22652 4468
rect 22560 4422 22612 4428
rect 22652 4422 22704 4428
rect 23032 4185 23060 7890
rect 23124 5778 23152 11834
rect 23676 11642 23704 12718
rect 23940 12640 23992 12646
rect 23940 12582 23992 12588
rect 23848 12096 23900 12102
rect 23848 12038 23900 12044
rect 23676 11626 23796 11642
rect 23572 11620 23624 11626
rect 23572 11562 23624 11568
rect 23676 11620 23808 11626
rect 23676 11614 23756 11620
rect 23204 11552 23256 11558
rect 23204 11494 23256 11500
rect 23216 6905 23244 11494
rect 23388 11008 23440 11014
rect 23388 10950 23440 10956
rect 23296 10804 23348 10810
rect 23296 10746 23348 10752
rect 23308 9586 23336 10746
rect 23400 10606 23428 10950
rect 23480 10668 23532 10674
rect 23480 10610 23532 10616
rect 23388 10600 23440 10606
rect 23388 10542 23440 10548
rect 23296 9580 23348 9586
rect 23296 9522 23348 9528
rect 23296 8832 23348 8838
rect 23296 8774 23348 8780
rect 23308 8634 23336 8774
rect 23296 8628 23348 8634
rect 23296 8570 23348 8576
rect 23400 8514 23428 10542
rect 23492 9654 23520 10610
rect 23480 9648 23532 9654
rect 23480 9590 23532 9596
rect 23480 8832 23532 8838
rect 23480 8774 23532 8780
rect 23308 8486 23428 8514
rect 23308 8430 23336 8486
rect 23296 8424 23348 8430
rect 23296 8366 23348 8372
rect 23308 7954 23336 8366
rect 23296 7948 23348 7954
rect 23296 7890 23348 7896
rect 23492 7818 23520 8774
rect 23480 7812 23532 7818
rect 23480 7754 23532 7760
rect 23478 7440 23534 7449
rect 23478 7375 23534 7384
rect 23296 7200 23348 7206
rect 23296 7142 23348 7148
rect 23308 7002 23336 7142
rect 23296 6996 23348 7002
rect 23296 6938 23348 6944
rect 23202 6896 23258 6905
rect 23202 6831 23258 6840
rect 23308 6662 23336 6938
rect 23388 6860 23440 6866
rect 23388 6802 23440 6808
rect 23296 6656 23348 6662
rect 23296 6598 23348 6604
rect 23400 6322 23428 6802
rect 23492 6458 23520 7375
rect 23584 6866 23612 11562
rect 23676 11014 23704 11614
rect 23756 11562 23808 11568
rect 23664 11008 23716 11014
rect 23664 10950 23716 10956
rect 23676 8838 23704 10950
rect 23664 8832 23716 8838
rect 23664 8774 23716 8780
rect 23664 8492 23716 8498
rect 23664 8434 23716 8440
rect 23676 8090 23704 8434
rect 23664 8084 23716 8090
rect 23664 8026 23716 8032
rect 23754 7848 23810 7857
rect 23754 7783 23756 7792
rect 23808 7783 23810 7792
rect 23756 7754 23808 7760
rect 23572 6860 23624 6866
rect 23572 6802 23624 6808
rect 23860 6746 23888 12038
rect 23952 11121 23980 12582
rect 24032 12096 24084 12102
rect 24032 12038 24084 12044
rect 23938 11112 23994 11121
rect 23938 11047 23994 11056
rect 23940 8832 23992 8838
rect 23940 8774 23992 8780
rect 23952 7206 23980 8774
rect 23940 7200 23992 7206
rect 23940 7142 23992 7148
rect 24044 7002 24072 12038
rect 24492 11552 24544 11558
rect 24492 11494 24544 11500
rect 24952 11552 25004 11558
rect 25056 11540 25084 12854
rect 25136 12708 25188 12714
rect 25136 12650 25188 12656
rect 25148 12442 25176 12650
rect 25136 12436 25188 12442
rect 25424 12434 25452 13806
rect 37070 13628 37378 13637
rect 37070 13626 37076 13628
rect 37132 13626 37156 13628
rect 37212 13626 37236 13628
rect 37292 13626 37316 13628
rect 37372 13626 37378 13628
rect 37132 13574 37134 13626
rect 37314 13574 37316 13626
rect 37070 13572 37076 13574
rect 37132 13572 37156 13574
rect 37212 13572 37236 13574
rect 37292 13572 37316 13574
rect 37372 13572 37378 13574
rect 37070 13563 37378 13572
rect 51518 13628 51826 13637
rect 51518 13626 51524 13628
rect 51580 13626 51604 13628
rect 51660 13626 51684 13628
rect 51740 13626 51764 13628
rect 51820 13626 51826 13628
rect 51580 13574 51582 13626
rect 51762 13574 51764 13626
rect 51518 13572 51524 13574
rect 51580 13572 51604 13574
rect 51660 13572 51684 13574
rect 51740 13572 51764 13574
rect 51820 13572 51826 13574
rect 51518 13563 51826 13572
rect 27804 13184 27856 13190
rect 27804 13126 27856 13132
rect 27816 12434 27844 13126
rect 29846 13084 30154 13093
rect 29846 13082 29852 13084
rect 29908 13082 29932 13084
rect 29988 13082 30012 13084
rect 30068 13082 30092 13084
rect 30148 13082 30154 13084
rect 29908 13030 29910 13082
rect 30090 13030 30092 13082
rect 29846 13028 29852 13030
rect 29908 13028 29932 13030
rect 29988 13028 30012 13030
rect 30068 13028 30092 13030
rect 30148 13028 30154 13030
rect 29846 13019 30154 13028
rect 44294 13084 44602 13093
rect 44294 13082 44300 13084
rect 44356 13082 44380 13084
rect 44436 13082 44460 13084
rect 44516 13082 44540 13084
rect 44596 13082 44602 13084
rect 44356 13030 44358 13082
rect 44538 13030 44540 13082
rect 44294 13028 44300 13030
rect 44356 13028 44380 13030
rect 44436 13028 44460 13030
rect 44516 13028 44540 13030
rect 44596 13028 44602 13030
rect 44294 13019 44602 13028
rect 37070 12540 37378 12549
rect 37070 12538 37076 12540
rect 37132 12538 37156 12540
rect 37212 12538 37236 12540
rect 37292 12538 37316 12540
rect 37372 12538 37378 12540
rect 37132 12486 37134 12538
rect 37314 12486 37316 12538
rect 37070 12484 37076 12486
rect 37132 12484 37156 12486
rect 37212 12484 37236 12486
rect 37292 12484 37316 12486
rect 37372 12484 37378 12486
rect 37070 12475 37378 12484
rect 51518 12540 51826 12549
rect 51518 12538 51524 12540
rect 51580 12538 51604 12540
rect 51660 12538 51684 12540
rect 51740 12538 51764 12540
rect 51820 12538 51826 12540
rect 51580 12486 51582 12538
rect 51762 12486 51764 12538
rect 51518 12484 51524 12486
rect 51580 12484 51604 12486
rect 51660 12484 51684 12486
rect 51740 12484 51764 12486
rect 51820 12484 51826 12486
rect 51518 12475 51826 12484
rect 25424 12406 25544 12434
rect 27816 12406 27936 12434
rect 25136 12378 25188 12384
rect 25004 11512 25084 11540
rect 24952 11494 25004 11500
rect 24124 11076 24176 11082
rect 24124 11018 24176 11024
rect 24136 7449 24164 11018
rect 24216 10464 24268 10470
rect 24216 10406 24268 10412
rect 24228 9489 24256 10406
rect 24400 10056 24452 10062
rect 24400 9998 24452 10004
rect 24412 9722 24440 9998
rect 24400 9716 24452 9722
rect 24400 9658 24452 9664
rect 24214 9480 24270 9489
rect 24214 9415 24270 9424
rect 24228 8537 24256 9415
rect 24400 9036 24452 9042
rect 24400 8978 24452 8984
rect 24412 8673 24440 8978
rect 24398 8664 24454 8673
rect 24398 8599 24454 8608
rect 24214 8528 24270 8537
rect 24400 8492 24452 8498
rect 24214 8463 24216 8472
rect 24268 8463 24270 8472
rect 24216 8434 24268 8440
rect 24320 8452 24400 8480
rect 24228 8403 24256 8434
rect 24320 7546 24348 8452
rect 24400 8434 24452 8440
rect 24308 7540 24360 7546
rect 24308 7482 24360 7488
rect 24122 7440 24178 7449
rect 24320 7410 24348 7482
rect 24122 7375 24178 7384
rect 24308 7404 24360 7410
rect 24032 6996 24084 7002
rect 24032 6938 24084 6944
rect 24136 6866 24164 7375
rect 24308 7346 24360 7352
rect 24400 6996 24452 7002
rect 24400 6938 24452 6944
rect 24032 6860 24084 6866
rect 24032 6802 24084 6808
rect 24124 6860 24176 6866
rect 24124 6802 24176 6808
rect 23572 6724 23624 6730
rect 23860 6718 23980 6746
rect 23572 6666 23624 6672
rect 23480 6452 23532 6458
rect 23480 6394 23532 6400
rect 23388 6316 23440 6322
rect 23388 6258 23440 6264
rect 23112 5772 23164 5778
rect 23112 5714 23164 5720
rect 23296 5772 23348 5778
rect 23296 5714 23348 5720
rect 23124 5166 23152 5714
rect 23202 5672 23258 5681
rect 23202 5607 23258 5616
rect 23112 5160 23164 5166
rect 23112 5102 23164 5108
rect 23112 4820 23164 4826
rect 23112 4762 23164 4768
rect 23124 4622 23152 4762
rect 23112 4616 23164 4622
rect 23112 4558 23164 4564
rect 23216 4554 23244 5607
rect 23308 5234 23336 5714
rect 23296 5228 23348 5234
rect 23296 5170 23348 5176
rect 23388 5228 23440 5234
rect 23388 5170 23440 5176
rect 23400 4826 23428 5170
rect 23388 4820 23440 4826
rect 23388 4762 23440 4768
rect 23296 4684 23348 4690
rect 23296 4626 23348 4632
rect 23204 4548 23256 4554
rect 23204 4490 23256 4496
rect 23308 4214 23336 4626
rect 23296 4208 23348 4214
rect 23018 4176 23074 4185
rect 23296 4150 23348 4156
rect 23018 4111 23074 4120
rect 23112 4072 23164 4078
rect 23112 4014 23164 4020
rect 23018 3904 23074 3913
rect 22622 3836 22930 3845
rect 23018 3839 23074 3848
rect 22622 3834 22628 3836
rect 22684 3834 22708 3836
rect 22764 3834 22788 3836
rect 22844 3834 22868 3836
rect 22924 3834 22930 3836
rect 22684 3782 22686 3834
rect 22866 3782 22868 3834
rect 22622 3780 22628 3782
rect 22684 3780 22708 3782
rect 22764 3780 22788 3782
rect 22844 3780 22868 3782
rect 22924 3780 22930 3782
rect 22622 3771 22930 3780
rect 22376 3732 22428 3738
rect 22376 3674 22428 3680
rect 22468 3732 22520 3738
rect 22468 3674 22520 3680
rect 22376 3392 22428 3398
rect 22376 3334 22428 3340
rect 22192 3188 22244 3194
rect 22192 3130 22244 3136
rect 22100 3120 22152 3126
rect 22100 3062 22152 3068
rect 21824 3052 21876 3058
rect 21824 2994 21876 3000
rect 21916 3052 21968 3058
rect 21916 2994 21968 3000
rect 21548 2848 21600 2854
rect 21548 2790 21600 2796
rect 21548 2644 21600 2650
rect 21548 2586 21600 2592
rect 21272 2576 21324 2582
rect 21272 2518 21324 2524
rect 21180 2440 21232 2446
rect 21180 2382 21232 2388
rect 21088 2100 21140 2106
rect 21088 2042 21140 2048
rect 20916 1142 21036 1170
rect 21008 800 21036 1142
rect 21284 800 21312 2518
rect 21560 800 21588 2586
rect 21836 2446 21864 2994
rect 22008 2848 22060 2854
rect 22008 2790 22060 2796
rect 22020 2530 22048 2790
rect 22112 2650 22140 3062
rect 22284 2916 22336 2922
rect 22284 2858 22336 2864
rect 22100 2644 22152 2650
rect 22100 2586 22152 2592
rect 22020 2502 22140 2530
rect 22112 2446 22140 2502
rect 21824 2440 21876 2446
rect 21824 2382 21876 2388
rect 22008 2440 22060 2446
rect 22008 2382 22060 2388
rect 22100 2440 22152 2446
rect 22100 2382 22152 2388
rect 21824 2304 21876 2310
rect 22020 2281 22048 2382
rect 21824 2246 21876 2252
rect 22006 2272 22062 2281
rect 21836 800 21864 2246
rect 22006 2207 22062 2216
rect 22296 1442 22324 2858
rect 22112 1414 22324 1442
rect 22112 800 22140 1414
rect 22388 800 22416 3334
rect 23032 3058 23060 3839
rect 23124 3126 23152 4014
rect 23386 3632 23442 3641
rect 23386 3567 23442 3576
rect 23400 3534 23428 3567
rect 23388 3528 23440 3534
rect 23388 3470 23440 3476
rect 23112 3120 23164 3126
rect 23112 3062 23164 3068
rect 23020 3052 23072 3058
rect 23020 2994 23072 3000
rect 22468 2848 22520 2854
rect 22468 2790 22520 2796
rect 22480 1442 22508 2790
rect 22622 2748 22930 2757
rect 22622 2746 22628 2748
rect 22684 2746 22708 2748
rect 22764 2746 22788 2748
rect 22844 2746 22868 2748
rect 22924 2746 22930 2748
rect 22684 2694 22686 2746
rect 22866 2694 22868 2746
rect 22622 2692 22628 2694
rect 22684 2692 22708 2694
rect 22764 2692 22788 2694
rect 22844 2692 22868 2694
rect 22924 2692 22930 2694
rect 22622 2683 22930 2692
rect 22836 2304 22888 2310
rect 22836 2246 22888 2252
rect 22928 2304 22980 2310
rect 22928 2246 22980 2252
rect 22848 1465 22876 2246
rect 22834 1456 22890 1465
rect 22480 1414 22692 1442
rect 22664 800 22692 1414
rect 22834 1391 22890 1400
rect 22940 800 22968 2246
rect 23032 2145 23060 2994
rect 23018 2136 23074 2145
rect 23018 2071 23074 2080
rect 23202 2000 23258 2009
rect 23202 1935 23258 1944
rect 23216 800 23244 1935
rect 23400 1193 23428 3470
rect 23492 3346 23520 6394
rect 23584 6322 23612 6666
rect 23572 6316 23624 6322
rect 23572 6258 23624 6264
rect 23848 5704 23900 5710
rect 23848 5646 23900 5652
rect 23754 5536 23810 5545
rect 23754 5471 23810 5480
rect 23664 4140 23716 4146
rect 23664 4082 23716 4088
rect 23676 3942 23704 4082
rect 23572 3936 23624 3942
rect 23572 3878 23624 3884
rect 23664 3936 23716 3942
rect 23664 3878 23716 3884
rect 23584 3466 23612 3878
rect 23572 3460 23624 3466
rect 23572 3402 23624 3408
rect 23492 3318 23612 3346
rect 23478 3224 23534 3233
rect 23478 3159 23534 3168
rect 23386 1184 23442 1193
rect 23386 1119 23442 1128
rect 23492 800 23520 3159
rect 23584 2514 23612 3318
rect 23572 2508 23624 2514
rect 23572 2450 23624 2456
rect 23768 800 23796 5471
rect 23860 3738 23888 5646
rect 23952 4536 23980 6718
rect 24044 6662 24072 6802
rect 24032 6656 24084 6662
rect 24032 6598 24084 6604
rect 24032 6316 24084 6322
rect 24032 6258 24084 6264
rect 24216 6316 24268 6322
rect 24216 6258 24268 6264
rect 24044 6186 24072 6258
rect 24228 6225 24256 6258
rect 24214 6216 24270 6225
rect 24032 6180 24084 6186
rect 24214 6151 24270 6160
rect 24032 6122 24084 6128
rect 24044 5642 24072 6122
rect 24228 5914 24256 6151
rect 24412 6089 24440 6938
rect 24398 6080 24454 6089
rect 24398 6015 24454 6024
rect 24216 5908 24268 5914
rect 24216 5850 24268 5856
rect 24032 5636 24084 5642
rect 24032 5578 24084 5584
rect 24032 4548 24084 4554
rect 23952 4508 24032 4536
rect 23952 4457 23980 4508
rect 24032 4490 24084 4496
rect 23938 4448 23994 4457
rect 23938 4383 23994 4392
rect 24214 4448 24270 4457
rect 24214 4383 24270 4392
rect 23952 4146 23980 4383
rect 24228 4282 24256 4383
rect 24216 4276 24268 4282
rect 24216 4218 24268 4224
rect 23940 4140 23992 4146
rect 23940 4082 23992 4088
rect 23848 3732 23900 3738
rect 23848 3674 23900 3680
rect 24308 2984 24360 2990
rect 24308 2926 24360 2932
rect 24032 1420 24084 1426
rect 24032 1362 24084 1368
rect 24044 800 24072 1362
rect 24320 800 24348 2926
rect 24412 2446 24440 6015
rect 24504 4865 24532 11494
rect 24768 11280 24820 11286
rect 24768 11222 24820 11228
rect 24676 10532 24728 10538
rect 24676 10474 24728 10480
rect 24688 10062 24716 10474
rect 24676 10056 24728 10062
rect 24676 9998 24728 10004
rect 24676 8492 24728 8498
rect 24676 8434 24728 8440
rect 24582 8392 24638 8401
rect 24582 8327 24638 8336
rect 24596 8294 24624 8327
rect 24688 8294 24716 8434
rect 24584 8288 24636 8294
rect 24584 8230 24636 8236
rect 24676 8288 24728 8294
rect 24676 8230 24728 8236
rect 24780 7886 24808 11222
rect 24860 9988 24912 9994
rect 24860 9930 24912 9936
rect 24872 9722 24900 9930
rect 24860 9716 24912 9722
rect 24860 9658 24912 9664
rect 24860 8968 24912 8974
rect 24860 8910 24912 8916
rect 24872 8090 24900 8910
rect 24860 8084 24912 8090
rect 24860 8026 24912 8032
rect 24584 7880 24636 7886
rect 24584 7822 24636 7828
rect 24768 7880 24820 7886
rect 24768 7822 24820 7828
rect 24596 7478 24624 7822
rect 24584 7472 24636 7478
rect 24584 7414 24636 7420
rect 24964 6914 24992 11494
rect 25044 9376 25096 9382
rect 25044 9318 25096 9324
rect 25056 8906 25084 9318
rect 25044 8900 25096 8906
rect 25044 8842 25096 8848
rect 25148 7834 25176 12378
rect 25412 11552 25464 11558
rect 25412 11494 25464 11500
rect 25228 10668 25280 10674
rect 25228 10610 25280 10616
rect 25240 9586 25268 10610
rect 25228 9580 25280 9586
rect 25228 9522 25280 9528
rect 25240 8634 25268 9522
rect 25228 8628 25280 8634
rect 25228 8570 25280 8576
rect 25240 8362 25268 8570
rect 25228 8356 25280 8362
rect 25228 8298 25280 8304
rect 25148 7806 25360 7834
rect 25228 7744 25280 7750
rect 25228 7686 25280 7692
rect 25240 7410 25268 7686
rect 25228 7404 25280 7410
rect 25228 7346 25280 7352
rect 25044 7336 25096 7342
rect 25042 7304 25044 7313
rect 25136 7336 25188 7342
rect 25096 7304 25098 7313
rect 25136 7278 25188 7284
rect 25042 7239 25098 7248
rect 24964 6886 25084 6914
rect 24860 6792 24912 6798
rect 24674 6760 24730 6769
rect 24860 6734 24912 6740
rect 24674 6695 24730 6704
rect 24688 6322 24716 6695
rect 24676 6316 24728 6322
rect 24676 6258 24728 6264
rect 24768 6248 24820 6254
rect 24766 6216 24768 6225
rect 24820 6216 24822 6225
rect 24766 6151 24822 6160
rect 24584 5296 24636 5302
rect 24584 5238 24636 5244
rect 24766 5264 24822 5273
rect 24490 4856 24546 4865
rect 24490 4791 24492 4800
rect 24544 4791 24546 4800
rect 24492 4762 24544 4768
rect 24504 4146 24532 4762
rect 24596 4282 24624 5238
rect 24766 5199 24822 5208
rect 24676 4480 24728 4486
rect 24676 4422 24728 4428
rect 24584 4276 24636 4282
rect 24584 4218 24636 4224
rect 24492 4140 24544 4146
rect 24492 4082 24544 4088
rect 24582 3904 24638 3913
rect 24582 3839 24638 3848
rect 24596 3058 24624 3839
rect 24584 3052 24636 3058
rect 24584 2994 24636 3000
rect 24688 2774 24716 4422
rect 24780 4146 24808 5199
rect 24768 4140 24820 4146
rect 24768 4082 24820 4088
rect 24596 2746 24716 2774
rect 24400 2440 24452 2446
rect 24400 2382 24452 2388
rect 24596 800 24624 2746
rect 24676 2440 24728 2446
rect 24676 2382 24728 2388
rect 24688 2106 24716 2382
rect 24676 2100 24728 2106
rect 24676 2042 24728 2048
rect 24872 800 24900 6734
rect 24952 6112 25004 6118
rect 24952 6054 25004 6060
rect 24964 5710 24992 6054
rect 24952 5704 25004 5710
rect 24952 5646 25004 5652
rect 24952 5024 25004 5030
rect 24952 4966 25004 4972
rect 24964 4622 24992 4966
rect 24952 4616 25004 4622
rect 24952 4558 25004 4564
rect 25056 4146 25084 6886
rect 25148 6866 25176 7278
rect 25136 6860 25188 6866
rect 25136 6802 25188 6808
rect 25148 6633 25176 6802
rect 25240 6730 25268 7346
rect 25228 6724 25280 6730
rect 25228 6666 25280 6672
rect 25134 6624 25190 6633
rect 25134 6559 25190 6568
rect 25228 4684 25280 4690
rect 25228 4626 25280 4632
rect 25240 4185 25268 4626
rect 25226 4176 25282 4185
rect 25044 4140 25096 4146
rect 25226 4111 25282 4120
rect 25044 4082 25096 4088
rect 25332 3942 25360 7806
rect 25424 6769 25452 11494
rect 25516 11354 25544 12406
rect 25596 12096 25648 12102
rect 25596 12038 25648 12044
rect 25504 11348 25556 11354
rect 25504 11290 25556 11296
rect 25410 6760 25466 6769
rect 25410 6695 25466 6704
rect 25504 6316 25556 6322
rect 25504 6258 25556 6264
rect 25516 6225 25544 6258
rect 25502 6216 25558 6225
rect 25502 6151 25558 6160
rect 25608 5216 25636 12038
rect 27436 11620 27488 11626
rect 27436 11562 27488 11568
rect 26332 11348 26384 11354
rect 26332 11290 26384 11296
rect 25872 11076 25924 11082
rect 25872 11018 25924 11024
rect 25688 10056 25740 10062
rect 25688 9998 25740 10004
rect 25700 9382 25728 9998
rect 25688 9376 25740 9382
rect 25688 9318 25740 9324
rect 25700 9110 25728 9318
rect 25688 9104 25740 9110
rect 25688 9046 25740 9052
rect 25780 8016 25832 8022
rect 25780 7958 25832 7964
rect 25792 7750 25820 7958
rect 25884 7857 25912 11018
rect 26240 10804 26292 10810
rect 26240 10746 26292 10752
rect 26056 10600 26108 10606
rect 26056 10542 26108 10548
rect 26068 9586 26096 10542
rect 26252 9586 26280 10746
rect 26344 9704 26372 11290
rect 27448 11150 27476 11562
rect 27436 11144 27488 11150
rect 27436 11086 27488 11092
rect 26608 11076 26660 11082
rect 26608 11018 26660 11024
rect 26700 11076 26752 11082
rect 26700 11018 26752 11024
rect 27528 11076 27580 11082
rect 27528 11018 27580 11024
rect 26424 10464 26476 10470
rect 26424 10406 26476 10412
rect 26436 10062 26464 10406
rect 26424 10056 26476 10062
rect 26424 9998 26476 10004
rect 26344 9676 26464 9704
rect 26056 9580 26108 9586
rect 26056 9522 26108 9528
rect 26240 9580 26292 9586
rect 26240 9522 26292 9528
rect 26332 9580 26384 9586
rect 26332 9522 26384 9528
rect 26344 9178 26372 9522
rect 26332 9172 26384 9178
rect 26332 9114 26384 9120
rect 25964 8900 26016 8906
rect 26240 8900 26292 8906
rect 25964 8842 26016 8848
rect 26160 8860 26240 8888
rect 25976 8498 26004 8842
rect 26160 8634 26188 8860
rect 26240 8842 26292 8848
rect 26148 8628 26200 8634
rect 26148 8570 26200 8576
rect 26160 8498 26188 8570
rect 25964 8492 26016 8498
rect 25964 8434 26016 8440
rect 26148 8492 26200 8498
rect 26148 8434 26200 8440
rect 25976 8090 26004 8434
rect 25964 8084 26016 8090
rect 25964 8026 26016 8032
rect 25976 7886 26004 8026
rect 26056 8016 26108 8022
rect 26056 7958 26108 7964
rect 25964 7880 26016 7886
rect 25870 7848 25926 7857
rect 25964 7822 26016 7828
rect 25870 7783 25926 7792
rect 25780 7744 25832 7750
rect 25780 7686 25832 7692
rect 25884 6322 25912 7783
rect 26068 7410 26096 7958
rect 26436 7954 26464 9676
rect 26424 7948 26476 7954
rect 26424 7890 26476 7896
rect 26240 7540 26292 7546
rect 26240 7482 26292 7488
rect 26252 7410 26280 7482
rect 26056 7404 26108 7410
rect 26056 7346 26108 7352
rect 26240 7404 26292 7410
rect 26240 7346 26292 7352
rect 26056 6928 26108 6934
rect 26056 6870 26108 6876
rect 25872 6316 25924 6322
rect 25872 6258 25924 6264
rect 25964 5364 26016 5370
rect 25964 5306 26016 5312
rect 25976 5234 26004 5306
rect 25964 5228 26016 5234
rect 25608 5188 25728 5216
rect 25504 5160 25556 5166
rect 25504 5102 25556 5108
rect 25594 5128 25650 5137
rect 25412 4752 25464 4758
rect 25412 4694 25464 4700
rect 25424 4214 25452 4694
rect 25516 4554 25544 5102
rect 25594 5063 25650 5072
rect 25504 4548 25556 4554
rect 25504 4490 25556 4496
rect 25412 4208 25464 4214
rect 25412 4150 25464 4156
rect 25320 3936 25372 3942
rect 25372 3896 25544 3924
rect 25320 3878 25372 3884
rect 25136 3732 25188 3738
rect 25136 3674 25188 3680
rect 25148 800 25176 3674
rect 25320 3664 25372 3670
rect 25372 3612 25452 3618
rect 25320 3606 25452 3612
rect 25332 3590 25452 3606
rect 25228 3460 25280 3466
rect 25228 3402 25280 3408
rect 25240 3194 25268 3402
rect 25228 3188 25280 3194
rect 25228 3130 25280 3136
rect 25320 2916 25372 2922
rect 25320 2858 25372 2864
rect 25332 1154 25360 2858
rect 25320 1148 25372 1154
rect 25320 1090 25372 1096
rect 25424 800 25452 3590
rect 25516 3194 25544 3896
rect 25504 3188 25556 3194
rect 25504 3130 25556 3136
rect 25504 3052 25556 3058
rect 25504 2994 25556 3000
rect 25516 2922 25544 2994
rect 25504 2916 25556 2922
rect 25504 2858 25556 2864
rect 25608 2774 25636 5063
rect 25700 4826 25728 5188
rect 25964 5170 26016 5176
rect 25688 4820 25740 4826
rect 25688 4762 25740 4768
rect 25700 4729 25728 4762
rect 25686 4720 25742 4729
rect 25686 4655 25742 4664
rect 25700 4026 25728 4655
rect 25976 4622 26004 5170
rect 25964 4616 26016 4622
rect 25964 4558 26016 4564
rect 25778 4448 25834 4457
rect 25778 4383 25834 4392
rect 25792 4146 25820 4383
rect 26068 4264 26096 6870
rect 26252 6440 26280 7346
rect 26436 7313 26464 7890
rect 26422 7304 26478 7313
rect 26422 7239 26478 7248
rect 26332 7200 26384 7206
rect 26332 7142 26384 7148
rect 26344 6712 26372 7142
rect 26436 6934 26464 7239
rect 26424 6928 26476 6934
rect 26424 6870 26476 6876
rect 26424 6724 26476 6730
rect 26344 6684 26424 6712
rect 26424 6666 26476 6672
rect 26160 6412 26280 6440
rect 26160 6322 26188 6412
rect 26148 6316 26200 6322
rect 26148 6258 26200 6264
rect 26240 6316 26292 6322
rect 26240 6258 26292 6264
rect 26252 5574 26280 6258
rect 26240 5568 26292 5574
rect 26240 5510 26292 5516
rect 26436 5234 26464 6666
rect 26424 5228 26476 5234
rect 25976 4236 26096 4264
rect 26344 5188 26424 5216
rect 25780 4140 25832 4146
rect 25780 4082 25832 4088
rect 25700 3998 25820 4026
rect 25688 3936 25740 3942
rect 25688 3878 25740 3884
rect 25700 3058 25728 3878
rect 25688 3052 25740 3058
rect 25688 2994 25740 3000
rect 25792 2922 25820 3998
rect 25976 3618 26004 4236
rect 26056 4140 26108 4146
rect 26056 4082 26108 4088
rect 26068 3738 26096 4082
rect 26056 3732 26108 3738
rect 26056 3674 26108 3680
rect 25976 3590 26188 3618
rect 25872 3188 25924 3194
rect 25872 3130 25924 3136
rect 25884 3058 25912 3130
rect 25872 3052 25924 3058
rect 25872 2994 25924 3000
rect 25780 2916 25832 2922
rect 25780 2858 25832 2864
rect 25608 2746 25728 2774
rect 25700 800 25728 2746
rect 25884 1737 25912 2994
rect 25964 2916 26016 2922
rect 25964 2858 26016 2864
rect 25870 1728 25926 1737
rect 25870 1663 25926 1672
rect 25976 800 26004 2858
rect 26160 1902 26188 3590
rect 26240 2032 26292 2038
rect 26240 1974 26292 1980
rect 26148 1896 26200 1902
rect 26148 1838 26200 1844
rect 26252 800 26280 1974
rect 26344 950 26372 5188
rect 26424 5170 26476 5176
rect 26620 4622 26648 11018
rect 26712 7721 26740 11018
rect 27160 10668 27212 10674
rect 27160 10610 27212 10616
rect 27172 9722 27200 10610
rect 27344 9920 27396 9926
rect 27344 9862 27396 9868
rect 27160 9716 27212 9722
rect 27160 9658 27212 9664
rect 26976 9512 27028 9518
rect 26976 9454 27028 9460
rect 26790 9072 26846 9081
rect 26988 9042 27016 9454
rect 26790 9007 26846 9016
rect 26976 9036 27028 9042
rect 26804 7818 26832 9007
rect 26976 8978 27028 8984
rect 26988 8906 27016 8978
rect 27068 8968 27120 8974
rect 27068 8910 27120 8916
rect 27158 8936 27214 8945
rect 26976 8900 27028 8906
rect 26976 8842 27028 8848
rect 27080 8634 27108 8910
rect 27158 8871 27160 8880
rect 27212 8871 27214 8880
rect 27160 8842 27212 8848
rect 27068 8628 27120 8634
rect 27068 8570 27120 8576
rect 27356 8498 27384 9862
rect 27436 8832 27488 8838
rect 27436 8774 27488 8780
rect 27344 8492 27396 8498
rect 27344 8434 27396 8440
rect 27356 8265 27384 8434
rect 27342 8256 27398 8265
rect 27342 8191 27398 8200
rect 27356 7993 27384 8191
rect 27342 7984 27398 7993
rect 26976 7948 27028 7954
rect 27342 7919 27398 7928
rect 26976 7890 27028 7896
rect 26792 7812 26844 7818
rect 26792 7754 26844 7760
rect 26698 7712 26754 7721
rect 26698 7647 26754 7656
rect 26712 6730 26740 7647
rect 26790 7440 26846 7449
rect 26790 7375 26846 7384
rect 26884 7404 26936 7410
rect 26804 7342 26832 7375
rect 26988 7392 27016 7890
rect 27448 7886 27476 8774
rect 27436 7880 27488 7886
rect 27436 7822 27488 7828
rect 26936 7364 27016 7392
rect 26884 7346 26936 7352
rect 26792 7336 26844 7342
rect 26792 7278 26844 7284
rect 26988 6934 27016 7364
rect 27252 7200 27304 7206
rect 27252 7142 27304 7148
rect 26976 6928 27028 6934
rect 26976 6870 27028 6876
rect 26700 6724 26752 6730
rect 26700 6666 26752 6672
rect 27264 6186 27292 7142
rect 27434 7032 27490 7041
rect 27434 6967 27490 6976
rect 27448 6730 27476 6967
rect 27436 6724 27488 6730
rect 27436 6666 27488 6672
rect 27434 6216 27490 6225
rect 27252 6180 27304 6186
rect 27434 6151 27436 6160
rect 27252 6122 27304 6128
rect 27488 6151 27490 6160
rect 27436 6122 27488 6128
rect 26976 5636 27028 5642
rect 26976 5578 27028 5584
rect 26988 5409 27016 5578
rect 26974 5400 27030 5409
rect 26974 5335 27030 5344
rect 27540 5302 27568 11018
rect 27620 10464 27672 10470
rect 27620 10406 27672 10412
rect 27632 8090 27660 10406
rect 27804 8288 27856 8294
rect 27804 8230 27856 8236
rect 27620 8084 27672 8090
rect 27620 8026 27672 8032
rect 27632 7886 27660 8026
rect 27816 7886 27844 8230
rect 27908 7886 27936 12406
rect 36820 12096 36872 12102
rect 36820 12038 36872 12044
rect 29846 11996 30154 12005
rect 29846 11994 29852 11996
rect 29908 11994 29932 11996
rect 29988 11994 30012 11996
rect 30068 11994 30092 11996
rect 30148 11994 30154 11996
rect 29908 11942 29910 11994
rect 30090 11942 30092 11994
rect 29846 11940 29852 11942
rect 29908 11940 29932 11942
rect 29988 11940 30012 11942
rect 30068 11940 30092 11942
rect 30148 11940 30154 11942
rect 29846 11931 30154 11940
rect 36544 11688 36596 11694
rect 36544 11630 36596 11636
rect 27988 11552 28040 11558
rect 27988 11494 28040 11500
rect 35716 11552 35768 11558
rect 35716 11494 35768 11500
rect 28000 11150 28028 11494
rect 27988 11144 28040 11150
rect 35728 11121 35756 11494
rect 27988 11086 28040 11092
rect 35714 11112 35770 11121
rect 29368 11076 29420 11082
rect 29368 11018 29420 11024
rect 35164 11076 35216 11082
rect 35714 11047 35770 11056
rect 36176 11076 36228 11082
rect 35164 11018 35216 11024
rect 36176 11018 36228 11024
rect 28908 10736 28960 10742
rect 28908 10678 28960 10684
rect 28816 10668 28868 10674
rect 28816 10610 28868 10616
rect 27988 9988 28040 9994
rect 27988 9930 28040 9936
rect 28080 9988 28132 9994
rect 28080 9930 28132 9936
rect 28000 9722 28028 9930
rect 27988 9716 28040 9722
rect 27988 9658 28040 9664
rect 27988 8968 28040 8974
rect 28092 8956 28120 9930
rect 28448 9920 28500 9926
rect 28448 9862 28500 9868
rect 28460 9625 28488 9862
rect 28446 9616 28502 9625
rect 28446 9551 28448 9560
rect 28500 9551 28502 9560
rect 28448 9522 28500 9528
rect 28828 9518 28856 10610
rect 28920 9994 28948 10678
rect 29092 10532 29144 10538
rect 29092 10474 29144 10480
rect 28908 9988 28960 9994
rect 28908 9930 28960 9936
rect 29000 9580 29052 9586
rect 29000 9522 29052 9528
rect 28816 9512 28868 9518
rect 28816 9454 28868 9460
rect 28816 9376 28868 9382
rect 28816 9318 28868 9324
rect 28828 8974 28856 9318
rect 29012 9081 29040 9522
rect 28998 9072 29054 9081
rect 28998 9007 29054 9016
rect 28040 8928 28120 8956
rect 28172 8968 28224 8974
rect 27988 8910 28040 8916
rect 28172 8910 28224 8916
rect 28816 8968 28868 8974
rect 28816 8910 28868 8916
rect 28000 8809 28028 8910
rect 27986 8800 28042 8809
rect 27986 8735 28042 8744
rect 28184 8294 28212 8910
rect 29012 8634 29040 9007
rect 29000 8628 29052 8634
rect 29000 8570 29052 8576
rect 28356 8492 28408 8498
rect 28632 8492 28684 8498
rect 28408 8452 28632 8480
rect 28356 8434 28408 8440
rect 28632 8434 28684 8440
rect 28172 8288 28224 8294
rect 28172 8230 28224 8236
rect 27620 7880 27672 7886
rect 27620 7822 27672 7828
rect 27804 7880 27856 7886
rect 27896 7880 27948 7886
rect 27804 7822 27856 7828
rect 27894 7848 27896 7857
rect 27948 7848 27950 7857
rect 27950 7806 28028 7834
rect 27894 7783 27950 7792
rect 28000 5522 28028 7806
rect 28368 7342 28396 8434
rect 28448 8356 28500 8362
rect 28448 8298 28500 8304
rect 28460 8090 28488 8298
rect 28448 8084 28500 8090
rect 28448 8026 28500 8032
rect 28724 8084 28776 8090
rect 28724 8026 28776 8032
rect 28736 7818 28764 8026
rect 28908 7880 28960 7886
rect 28908 7822 28960 7828
rect 28724 7812 28776 7818
rect 28724 7754 28776 7760
rect 28356 7336 28408 7342
rect 28356 7278 28408 7284
rect 28736 6866 28764 7754
rect 28816 6996 28868 7002
rect 28816 6938 28868 6944
rect 28724 6860 28776 6866
rect 28724 6802 28776 6808
rect 28828 6458 28856 6938
rect 28920 6730 28948 7822
rect 29000 7404 29052 7410
rect 29000 7346 29052 7352
rect 29012 7313 29040 7346
rect 28998 7304 29054 7313
rect 28998 7239 29054 7248
rect 29000 6792 29052 6798
rect 29000 6734 29052 6740
rect 28908 6724 28960 6730
rect 28908 6666 28960 6672
rect 29012 6662 29040 6734
rect 29000 6656 29052 6662
rect 29000 6598 29052 6604
rect 28816 6452 28868 6458
rect 28816 6394 28868 6400
rect 28828 6322 28856 6394
rect 28080 6316 28132 6322
rect 28080 6258 28132 6264
rect 28816 6316 28868 6322
rect 28816 6258 28868 6264
rect 28092 5914 28120 6258
rect 28724 6112 28776 6118
rect 28724 6054 28776 6060
rect 28080 5908 28132 5914
rect 28080 5850 28132 5856
rect 28736 5710 28764 6054
rect 29012 5953 29040 6598
rect 28998 5944 29054 5953
rect 28998 5879 29054 5888
rect 28724 5704 28776 5710
rect 28724 5646 28776 5652
rect 29000 5704 29052 5710
rect 29000 5646 29052 5652
rect 28000 5494 28120 5522
rect 27988 5364 28040 5370
rect 27988 5306 28040 5312
rect 27528 5296 27580 5302
rect 26882 5264 26938 5273
rect 27528 5238 27580 5244
rect 26882 5199 26938 5208
rect 26896 5030 26924 5199
rect 26792 5024 26844 5030
rect 26792 4966 26844 4972
rect 26884 5024 26936 5030
rect 26884 4966 26936 4972
rect 26608 4616 26660 4622
rect 26608 4558 26660 4564
rect 26514 4312 26570 4321
rect 26514 4247 26570 4256
rect 26422 1864 26478 1873
rect 26422 1799 26478 1808
rect 26436 950 26464 1799
rect 26332 944 26384 950
rect 26332 886 26384 892
rect 26424 944 26476 950
rect 26424 886 26476 892
rect 26528 800 26556 4247
rect 26620 950 26648 4558
rect 26804 3942 26832 4966
rect 27540 4214 27568 5238
rect 28000 5234 28028 5306
rect 27712 5228 27764 5234
rect 27712 5170 27764 5176
rect 27804 5228 27856 5234
rect 27804 5170 27856 5176
rect 27988 5228 28040 5234
rect 27988 5170 28040 5176
rect 27724 5098 27752 5170
rect 27712 5092 27764 5098
rect 27712 5034 27764 5040
rect 27816 5030 27844 5170
rect 27804 5024 27856 5030
rect 27804 4966 27856 4972
rect 27816 4826 27844 4966
rect 27804 4820 27856 4826
rect 27804 4762 27856 4768
rect 27896 4480 27948 4486
rect 27896 4422 27948 4428
rect 27528 4208 27580 4214
rect 27528 4150 27580 4156
rect 26792 3936 26844 3942
rect 26792 3878 26844 3884
rect 26884 3732 26936 3738
rect 26884 3674 26936 3680
rect 27068 3732 27120 3738
rect 27068 3674 27120 3680
rect 26792 2848 26844 2854
rect 26792 2790 26844 2796
rect 26608 944 26660 950
rect 26608 886 26660 892
rect 26804 800 26832 2790
rect 26896 1154 26924 3674
rect 26976 2440 27028 2446
rect 26974 2408 26976 2417
rect 27028 2408 27030 2417
rect 26974 2343 27030 2352
rect 26988 2310 27016 2343
rect 26976 2304 27028 2310
rect 26976 2246 27028 2252
rect 26884 1148 26936 1154
rect 26884 1090 26936 1096
rect 27080 800 27108 3674
rect 27908 3602 27936 4422
rect 28000 4214 28028 5170
rect 27988 4208 28040 4214
rect 27988 4150 28040 4156
rect 27896 3596 27948 3602
rect 27896 3538 27948 3544
rect 27620 3528 27672 3534
rect 27620 3470 27672 3476
rect 27712 3528 27764 3534
rect 27712 3470 27764 3476
rect 27528 3460 27580 3466
rect 27528 3402 27580 3408
rect 27344 3392 27396 3398
rect 27344 3334 27396 3340
rect 27356 800 27384 3334
rect 27540 3126 27568 3402
rect 27528 3120 27580 3126
rect 27528 3062 27580 3068
rect 27632 800 27660 3470
rect 27724 3058 27752 3470
rect 27802 3360 27858 3369
rect 27802 3295 27858 3304
rect 27712 3052 27764 3058
rect 27712 2994 27764 3000
rect 27724 1630 27752 2994
rect 27712 1624 27764 1630
rect 27712 1566 27764 1572
rect 27816 1442 27844 3295
rect 27908 2650 27936 3538
rect 28092 2774 28120 5494
rect 28448 5228 28500 5234
rect 28448 5170 28500 5176
rect 28724 5228 28776 5234
rect 28724 5170 28776 5176
rect 28460 4690 28488 5170
rect 28736 5098 28764 5170
rect 28906 5128 28962 5137
rect 28724 5092 28776 5098
rect 28906 5063 28908 5072
rect 28724 5034 28776 5040
rect 28960 5063 28962 5072
rect 28908 5034 28960 5040
rect 28448 4684 28500 4690
rect 28448 4626 28500 4632
rect 28736 4282 28764 5034
rect 28724 4276 28776 4282
rect 28724 4218 28776 4224
rect 28448 3936 28500 3942
rect 28448 3878 28500 3884
rect 28264 3664 28316 3670
rect 28264 3606 28316 3612
rect 28172 3460 28224 3466
rect 28172 3402 28224 3408
rect 28184 3126 28212 3402
rect 28172 3120 28224 3126
rect 28172 3062 28224 3068
rect 28276 2774 28304 3606
rect 28000 2746 28120 2774
rect 28184 2746 28304 2774
rect 27896 2644 27948 2650
rect 27896 2586 27948 2592
rect 28000 2281 28028 2746
rect 27986 2272 28042 2281
rect 27986 2207 28042 2216
rect 27816 1414 27936 1442
rect 27908 800 27936 1414
rect 28184 800 28212 2746
rect 28460 800 28488 3878
rect 29012 3194 29040 5646
rect 29000 3188 29052 3194
rect 29000 3130 29052 3136
rect 29104 2990 29132 10474
rect 29184 8832 29236 8838
rect 29184 8774 29236 8780
rect 29196 8294 29224 8774
rect 29184 8288 29236 8294
rect 29184 8230 29236 8236
rect 29380 5114 29408 11018
rect 29846 10908 30154 10917
rect 29846 10906 29852 10908
rect 29908 10906 29932 10908
rect 29988 10906 30012 10908
rect 30068 10906 30092 10908
rect 30148 10906 30154 10908
rect 29908 10854 29910 10906
rect 30090 10854 30092 10906
rect 29846 10852 29852 10854
rect 29908 10852 29932 10854
rect 29988 10852 30012 10854
rect 30068 10852 30092 10854
rect 30148 10852 30154 10854
rect 29846 10843 30154 10852
rect 34612 10736 34664 10742
rect 34612 10678 34664 10684
rect 31208 10600 31260 10606
rect 31208 10542 31260 10548
rect 34520 10600 34572 10606
rect 34520 10542 34572 10548
rect 29552 10464 29604 10470
rect 29552 10406 29604 10412
rect 30196 10464 30248 10470
rect 30196 10406 30248 10412
rect 29460 9920 29512 9926
rect 29460 9862 29512 9868
rect 29472 9466 29500 9862
rect 29564 9586 29592 10406
rect 29846 9820 30154 9829
rect 29846 9818 29852 9820
rect 29908 9818 29932 9820
rect 29988 9818 30012 9820
rect 30068 9818 30092 9820
rect 30148 9818 30154 9820
rect 29908 9766 29910 9818
rect 30090 9766 30092 9818
rect 29846 9764 29852 9766
rect 29908 9764 29932 9766
rect 29988 9764 30012 9766
rect 30068 9764 30092 9766
rect 30148 9764 30154 9766
rect 29846 9755 30154 9764
rect 29552 9580 29604 9586
rect 29552 9522 29604 9528
rect 29644 9580 29696 9586
rect 29644 9522 29696 9528
rect 29656 9466 29684 9522
rect 29472 9438 29684 9466
rect 29472 8906 29500 9438
rect 30012 9376 30064 9382
rect 30012 9318 30064 9324
rect 29460 8900 29512 8906
rect 29460 8842 29512 8848
rect 30024 8838 30052 9318
rect 29552 8832 29604 8838
rect 29552 8774 29604 8780
rect 30012 8832 30064 8838
rect 30012 8774 30064 8780
rect 29458 8528 29514 8537
rect 29458 8463 29514 8472
rect 29472 6662 29500 8463
rect 29460 6656 29512 6662
rect 29460 6598 29512 6604
rect 29460 6316 29512 6322
rect 29564 6304 29592 8774
rect 29846 8732 30154 8741
rect 29846 8730 29852 8732
rect 29908 8730 29932 8732
rect 29988 8730 30012 8732
rect 30068 8730 30092 8732
rect 30148 8730 30154 8732
rect 29908 8678 29910 8730
rect 30090 8678 30092 8730
rect 29846 8676 29852 8678
rect 29908 8676 29932 8678
rect 29988 8676 30012 8678
rect 30068 8676 30092 8678
rect 30148 8676 30154 8678
rect 29846 8667 30154 8676
rect 29736 8424 29788 8430
rect 29736 8366 29788 8372
rect 29748 7886 29776 8366
rect 29736 7880 29788 7886
rect 29736 7822 29788 7828
rect 29642 7576 29698 7585
rect 29642 7511 29698 7520
rect 29656 7410 29684 7511
rect 29644 7404 29696 7410
rect 29644 7346 29696 7352
rect 29748 7274 29776 7822
rect 29846 7644 30154 7653
rect 29846 7642 29852 7644
rect 29908 7642 29932 7644
rect 29988 7642 30012 7644
rect 30068 7642 30092 7644
rect 30148 7642 30154 7644
rect 29908 7590 29910 7642
rect 30090 7590 30092 7642
rect 29846 7588 29852 7590
rect 29908 7588 29932 7590
rect 29988 7588 30012 7590
rect 30068 7588 30092 7590
rect 30148 7588 30154 7590
rect 29846 7579 30154 7588
rect 29828 7336 29880 7342
rect 29828 7278 29880 7284
rect 29736 7268 29788 7274
rect 29736 7210 29788 7216
rect 29734 7032 29790 7041
rect 29734 6967 29736 6976
rect 29788 6967 29790 6976
rect 29736 6938 29788 6944
rect 29840 6662 29868 7278
rect 29828 6656 29880 6662
rect 29828 6598 29880 6604
rect 29846 6556 30154 6565
rect 29846 6554 29852 6556
rect 29908 6554 29932 6556
rect 29988 6554 30012 6556
rect 30068 6554 30092 6556
rect 30148 6554 30154 6556
rect 29908 6502 29910 6554
rect 30090 6502 30092 6554
rect 29846 6500 29852 6502
rect 29908 6500 29932 6502
rect 29988 6500 30012 6502
rect 30068 6500 30092 6502
rect 30148 6500 30154 6502
rect 29846 6491 30154 6500
rect 29644 6316 29696 6322
rect 29564 6276 29644 6304
rect 29460 6258 29512 6264
rect 29644 6258 29696 6264
rect 29472 5914 29500 6258
rect 29920 6112 29972 6118
rect 29920 6054 29972 6060
rect 29460 5908 29512 5914
rect 29460 5850 29512 5856
rect 29748 5846 29776 5877
rect 29736 5840 29788 5846
rect 29734 5808 29736 5817
rect 29788 5808 29790 5817
rect 29734 5743 29790 5752
rect 29748 5710 29776 5743
rect 29736 5704 29788 5710
rect 29736 5646 29788 5652
rect 29932 5642 29960 6054
rect 29920 5636 29972 5642
rect 29920 5578 29972 5584
rect 29846 5468 30154 5477
rect 29846 5466 29852 5468
rect 29908 5466 29932 5468
rect 29988 5466 30012 5468
rect 30068 5466 30092 5468
rect 30148 5466 30154 5468
rect 29908 5414 29910 5466
rect 30090 5414 30092 5466
rect 29846 5412 29852 5414
rect 29908 5412 29932 5414
rect 29988 5412 30012 5414
rect 30068 5412 30092 5414
rect 30148 5412 30154 5414
rect 29846 5403 30154 5412
rect 29380 5086 29592 5114
rect 29460 5024 29512 5030
rect 29460 4966 29512 4972
rect 29368 4820 29420 4826
rect 29368 4762 29420 4768
rect 29380 4214 29408 4762
rect 29368 4208 29420 4214
rect 29182 4176 29238 4185
rect 29368 4150 29420 4156
rect 29182 4111 29238 4120
rect 28724 2984 28776 2990
rect 28724 2926 28776 2932
rect 29092 2984 29144 2990
rect 29092 2926 29144 2932
rect 28736 800 28764 2926
rect 29196 2774 29224 4111
rect 29276 4004 29328 4010
rect 29276 3946 29328 3952
rect 29288 3058 29316 3946
rect 29276 3052 29328 3058
rect 29276 2994 29328 3000
rect 29368 2984 29420 2990
rect 29368 2926 29420 2932
rect 29196 2746 29316 2774
rect 29000 2372 29052 2378
rect 29000 2314 29052 2320
rect 29012 800 29040 2314
rect 29288 800 29316 2746
rect 29380 1873 29408 2926
rect 29366 1864 29422 1873
rect 29366 1799 29422 1808
rect 29472 1426 29500 4966
rect 29564 3534 29592 5086
rect 29642 4992 29698 5001
rect 29642 4927 29698 4936
rect 29656 4622 29684 4927
rect 30208 4622 30236 10406
rect 31220 10062 31248 10542
rect 33140 10464 33192 10470
rect 33140 10406 33192 10412
rect 32312 10124 32364 10130
rect 32312 10066 32364 10072
rect 30840 10056 30892 10062
rect 30840 9998 30892 10004
rect 31208 10056 31260 10062
rect 31208 9998 31260 10004
rect 30564 9988 30616 9994
rect 30564 9930 30616 9936
rect 30288 9920 30340 9926
rect 30288 9862 30340 9868
rect 30300 9382 30328 9862
rect 30576 9654 30604 9930
rect 30852 9722 30880 9998
rect 32324 9722 32352 10066
rect 32496 9920 32548 9926
rect 32496 9862 32548 9868
rect 32588 9920 32640 9926
rect 32588 9862 32640 9868
rect 32508 9722 32536 9862
rect 30840 9716 30892 9722
rect 30840 9658 30892 9664
rect 32312 9716 32364 9722
rect 32312 9658 32364 9664
rect 32496 9716 32548 9722
rect 32496 9658 32548 9664
rect 30564 9648 30616 9654
rect 30564 9590 30616 9596
rect 31760 9648 31812 9654
rect 31760 9590 31812 9596
rect 30288 9376 30340 9382
rect 30288 9318 30340 9324
rect 30576 8974 30604 9590
rect 30748 9580 30800 9586
rect 30748 9522 30800 9528
rect 31576 9580 31628 9586
rect 31576 9522 31628 9528
rect 30760 9178 30788 9522
rect 31300 9444 31352 9450
rect 31300 9386 31352 9392
rect 31116 9376 31168 9382
rect 31116 9318 31168 9324
rect 30748 9172 30800 9178
rect 30748 9114 30800 9120
rect 30564 8968 30616 8974
rect 30564 8910 30616 8916
rect 30656 8900 30708 8906
rect 30656 8842 30708 8848
rect 30288 8492 30340 8498
rect 30340 8452 30512 8480
rect 30288 8434 30340 8440
rect 30288 8356 30340 8362
rect 30484 8344 30512 8452
rect 30564 8356 30616 8362
rect 30340 8316 30420 8344
rect 30484 8316 30564 8344
rect 30288 8298 30340 8304
rect 30392 7818 30420 8316
rect 30564 8298 30616 8304
rect 30668 8090 30696 8842
rect 31022 8528 31078 8537
rect 30840 8492 30892 8498
rect 31022 8463 31024 8472
rect 30840 8434 30892 8440
rect 31076 8463 31078 8472
rect 31024 8434 31076 8440
rect 30656 8084 30708 8090
rect 30656 8026 30708 8032
rect 30380 7812 30432 7818
rect 30380 7754 30432 7760
rect 30748 7744 30800 7750
rect 30748 7686 30800 7692
rect 30378 7576 30434 7585
rect 30378 7511 30434 7520
rect 30392 6905 30420 7511
rect 30378 6896 30434 6905
rect 30378 6831 30434 6840
rect 30564 6792 30616 6798
rect 30564 6734 30616 6740
rect 30380 6724 30432 6730
rect 30380 6666 30432 6672
rect 30392 6390 30420 6666
rect 30380 6384 30432 6390
rect 30380 6326 30432 6332
rect 30472 6384 30524 6390
rect 30472 6326 30524 6332
rect 30484 5930 30512 6326
rect 30576 6118 30604 6734
rect 30564 6112 30616 6118
rect 30564 6054 30616 6060
rect 30484 5902 30604 5930
rect 30472 5840 30524 5846
rect 30472 5782 30524 5788
rect 30380 5704 30432 5710
rect 30378 5672 30380 5681
rect 30432 5672 30434 5681
rect 30378 5607 30434 5616
rect 30288 5228 30340 5234
rect 30288 5170 30340 5176
rect 30300 4826 30328 5170
rect 30288 4820 30340 4826
rect 30288 4762 30340 4768
rect 29644 4616 29696 4622
rect 29920 4616 29972 4622
rect 29644 4558 29696 4564
rect 29748 4576 29920 4604
rect 29552 3528 29604 3534
rect 29552 3470 29604 3476
rect 29748 2774 29776 4576
rect 29920 4558 29972 4564
rect 30196 4616 30248 4622
rect 30196 4558 30248 4564
rect 30288 4548 30340 4554
rect 30288 4490 30340 4496
rect 29846 4380 30154 4389
rect 29846 4378 29852 4380
rect 29908 4378 29932 4380
rect 29988 4378 30012 4380
rect 30068 4378 30092 4380
rect 30148 4378 30154 4380
rect 29908 4326 29910 4378
rect 30090 4326 30092 4378
rect 29846 4324 29852 4326
rect 29908 4324 29932 4326
rect 29988 4324 30012 4326
rect 30068 4324 30092 4326
rect 30148 4324 30154 4326
rect 29846 4315 30154 4324
rect 30102 4176 30158 4185
rect 30300 4146 30328 4490
rect 30102 4111 30104 4120
rect 30156 4111 30158 4120
rect 30288 4140 30340 4146
rect 30104 4082 30156 4088
rect 30288 4082 30340 4088
rect 29846 3292 30154 3301
rect 29846 3290 29852 3292
rect 29908 3290 29932 3292
rect 29988 3290 30012 3292
rect 30068 3290 30092 3292
rect 30148 3290 30154 3292
rect 29908 3238 29910 3290
rect 30090 3238 30092 3290
rect 29846 3236 29852 3238
rect 29908 3236 29932 3238
rect 29988 3236 30012 3238
rect 30068 3236 30092 3238
rect 30148 3236 30154 3238
rect 29846 3227 30154 3236
rect 30484 3126 30512 5782
rect 30576 3913 30604 5902
rect 30760 5574 30788 7686
rect 30852 7041 30880 8434
rect 30838 7032 30894 7041
rect 30838 6967 30894 6976
rect 30838 6896 30894 6905
rect 30838 6831 30894 6840
rect 30748 5568 30800 5574
rect 30748 5510 30800 5516
rect 30852 4826 30880 6831
rect 31022 4856 31078 4865
rect 30840 4820 30892 4826
rect 31022 4791 31078 4800
rect 30840 4762 30892 4768
rect 31036 4622 31064 4791
rect 31024 4616 31076 4622
rect 31024 4558 31076 4564
rect 31036 4282 31064 4558
rect 31024 4276 31076 4282
rect 31024 4218 31076 4224
rect 30562 3904 30618 3913
rect 30562 3839 30618 3848
rect 30840 3664 30892 3670
rect 30840 3606 30892 3612
rect 31128 3618 31156 9318
rect 31312 8956 31340 9386
rect 31588 9178 31616 9522
rect 31576 9172 31628 9178
rect 31576 9114 31628 9120
rect 31392 8968 31444 8974
rect 31312 8928 31392 8956
rect 31392 8910 31444 8916
rect 31208 8492 31260 8498
rect 31208 8434 31260 8440
rect 31220 8362 31248 8434
rect 31404 8362 31432 8910
rect 31484 8628 31536 8634
rect 31484 8570 31536 8576
rect 31496 8537 31524 8570
rect 31482 8528 31538 8537
rect 31482 8463 31538 8472
rect 31208 8356 31260 8362
rect 31208 8298 31260 8304
rect 31392 8356 31444 8362
rect 31392 8298 31444 8304
rect 31300 7880 31352 7886
rect 31300 7822 31352 7828
rect 31312 7206 31340 7822
rect 31576 7744 31628 7750
rect 31576 7686 31628 7692
rect 31588 7342 31616 7686
rect 31576 7336 31628 7342
rect 31576 7278 31628 7284
rect 31300 7200 31352 7206
rect 31300 7142 31352 7148
rect 31392 6724 31444 6730
rect 31392 6666 31444 6672
rect 31208 6112 31260 6118
rect 31208 6054 31260 6060
rect 31220 3738 31248 6054
rect 31300 5364 31352 5370
rect 31300 5306 31352 5312
rect 31312 4214 31340 5306
rect 31300 4208 31352 4214
rect 31300 4150 31352 4156
rect 31312 4078 31340 4150
rect 31300 4072 31352 4078
rect 31300 4014 31352 4020
rect 31208 3732 31260 3738
rect 31208 3674 31260 3680
rect 30472 3120 30524 3126
rect 30472 3062 30524 3068
rect 30852 3058 30880 3606
rect 31128 3590 31248 3618
rect 31220 3369 31248 3590
rect 31300 3460 31352 3466
rect 31300 3402 31352 3408
rect 31206 3360 31262 3369
rect 31206 3295 31262 3304
rect 30840 3052 30892 3058
rect 30840 2994 30892 3000
rect 31024 3055 31076 3061
rect 31220 3058 31248 3295
rect 31312 3126 31340 3402
rect 31300 3120 31352 3126
rect 31300 3062 31352 3068
rect 31024 2997 31076 3003
rect 31208 3052 31260 3058
rect 30748 2984 30800 2990
rect 30748 2926 30800 2932
rect 29656 2746 29776 2774
rect 29552 2644 29604 2650
rect 29552 2586 29604 2592
rect 29460 1420 29512 1426
rect 29460 1362 29512 1368
rect 29564 800 29592 2586
rect 29656 1018 29684 2746
rect 30656 2576 30708 2582
rect 30656 2518 30708 2524
rect 29736 2508 29788 2514
rect 29736 2450 29788 2456
rect 29748 1306 29776 2450
rect 30196 2440 30248 2446
rect 30196 2382 30248 2388
rect 30380 2440 30432 2446
rect 30380 2382 30432 2388
rect 29846 2204 30154 2213
rect 29846 2202 29852 2204
rect 29908 2202 29932 2204
rect 29988 2202 30012 2204
rect 30068 2202 30092 2204
rect 30148 2202 30154 2204
rect 29908 2150 29910 2202
rect 30090 2150 30092 2202
rect 29846 2148 29852 2150
rect 29908 2148 29932 2150
rect 29988 2148 30012 2150
rect 30068 2148 30092 2150
rect 30148 2148 30154 2150
rect 29846 2139 30154 2148
rect 30208 1306 30236 2382
rect 29748 1278 29868 1306
rect 29644 1012 29696 1018
rect 29644 954 29696 960
rect 29840 800 29868 1278
rect 30116 1278 30236 1306
rect 30116 800 30144 1278
rect 30392 800 30420 2382
rect 30668 800 30696 2518
rect 30760 1601 30788 2926
rect 30852 2825 30880 2994
rect 30838 2816 30894 2825
rect 30838 2751 30894 2760
rect 31036 2650 31064 2997
rect 31208 2994 31260 3000
rect 31300 2984 31352 2990
rect 31300 2926 31352 2932
rect 31208 2916 31260 2922
rect 31208 2858 31260 2864
rect 31024 2644 31076 2650
rect 31024 2586 31076 2592
rect 30932 2508 30984 2514
rect 30932 2450 30984 2456
rect 30746 1592 30802 1601
rect 30746 1527 30802 1536
rect 30944 800 30972 2450
rect 31220 800 31248 2858
rect 31312 2310 31340 2926
rect 31300 2304 31352 2310
rect 31300 2246 31352 2252
rect 31404 1698 31432 6666
rect 31668 6384 31720 6390
rect 31772 6372 31800 9590
rect 32220 8288 32272 8294
rect 32218 8256 32220 8265
rect 32272 8256 32274 8265
rect 32218 8191 32274 8200
rect 32232 7886 32260 8191
rect 32220 7880 32272 7886
rect 32220 7822 32272 7828
rect 31852 7744 31904 7750
rect 31852 7686 31904 7692
rect 32036 7744 32088 7750
rect 32036 7686 32088 7692
rect 31864 7410 31892 7686
rect 31852 7404 31904 7410
rect 31852 7346 31904 7352
rect 31850 7304 31906 7313
rect 31850 7239 31906 7248
rect 31864 6798 31892 7239
rect 32048 7041 32076 7686
rect 32034 7032 32090 7041
rect 32034 6967 32090 6976
rect 32048 6866 32076 6967
rect 32232 6934 32260 7822
rect 32312 7744 32364 7750
rect 32312 7686 32364 7692
rect 32324 7274 32352 7686
rect 32312 7268 32364 7274
rect 32312 7210 32364 7216
rect 32600 6934 32628 9862
rect 32956 9580 33008 9586
rect 32956 9522 33008 9528
rect 32772 9512 32824 9518
rect 32772 9454 32824 9460
rect 32784 9110 32812 9454
rect 32968 9178 32996 9522
rect 32956 9172 33008 9178
rect 32956 9114 33008 9120
rect 33048 9172 33100 9178
rect 33048 9114 33100 9120
rect 32772 9104 32824 9110
rect 32772 9046 32824 9052
rect 33060 8498 33088 9114
rect 33152 8514 33180 10406
rect 33324 10056 33376 10062
rect 33324 9998 33376 10004
rect 33336 8974 33364 9998
rect 34152 9920 34204 9926
rect 34152 9862 34204 9868
rect 34164 9722 34192 9862
rect 34152 9716 34204 9722
rect 34152 9658 34204 9664
rect 33600 9104 33652 9110
rect 33600 9046 33652 9052
rect 33232 8968 33284 8974
rect 33232 8910 33284 8916
rect 33324 8968 33376 8974
rect 33324 8910 33376 8916
rect 33244 8634 33272 8910
rect 33336 8634 33364 8910
rect 33416 8832 33468 8838
rect 33416 8774 33468 8780
rect 33232 8628 33284 8634
rect 33232 8570 33284 8576
rect 33324 8628 33376 8634
rect 33324 8570 33376 8576
rect 33048 8492 33100 8498
rect 33152 8486 33272 8514
rect 33048 8434 33100 8440
rect 32864 8424 32916 8430
rect 32864 8366 32916 8372
rect 32876 7886 32904 8366
rect 33244 8022 33272 8486
rect 33232 8016 33284 8022
rect 33232 7958 33284 7964
rect 32864 7880 32916 7886
rect 32864 7822 32916 7828
rect 32220 6928 32272 6934
rect 32220 6870 32272 6876
rect 32588 6928 32640 6934
rect 32588 6870 32640 6876
rect 33140 6928 33192 6934
rect 33140 6870 33192 6876
rect 32036 6860 32088 6866
rect 32036 6802 32088 6808
rect 31852 6792 31904 6798
rect 32496 6792 32548 6798
rect 31852 6734 31904 6740
rect 31956 6740 32496 6746
rect 31956 6734 32548 6740
rect 31864 6497 31892 6734
rect 31956 6718 32536 6734
rect 32956 6724 33008 6730
rect 31850 6488 31906 6497
rect 31956 6458 31984 6718
rect 32956 6666 33008 6672
rect 32404 6656 32456 6662
rect 32404 6598 32456 6604
rect 31850 6423 31906 6432
rect 31944 6452 31996 6458
rect 31944 6394 31996 6400
rect 31720 6344 31800 6372
rect 32312 6384 32364 6390
rect 32310 6352 32312 6361
rect 32364 6352 32366 6361
rect 31668 6326 31720 6332
rect 32416 6322 32444 6598
rect 32968 6390 32996 6666
rect 33152 6390 33180 6870
rect 33244 6662 33272 7958
rect 33428 7886 33456 8774
rect 33612 8430 33640 9046
rect 33600 8424 33652 8430
rect 33598 8392 33600 8401
rect 33652 8392 33654 8401
rect 33598 8327 33654 8336
rect 33968 8288 34020 8294
rect 33968 8230 34020 8236
rect 33416 7880 33468 7886
rect 33416 7822 33468 7828
rect 33428 7002 33456 7822
rect 33980 7410 34008 8230
rect 33968 7404 34020 7410
rect 33968 7346 34020 7352
rect 33600 7200 33652 7206
rect 33600 7142 33652 7148
rect 33612 7002 33640 7142
rect 33416 6996 33468 7002
rect 33416 6938 33468 6944
rect 33600 6996 33652 7002
rect 33600 6938 33652 6944
rect 33232 6656 33284 6662
rect 33232 6598 33284 6604
rect 32956 6384 33008 6390
rect 32956 6326 33008 6332
rect 33140 6384 33192 6390
rect 33140 6326 33192 6332
rect 32310 6287 32366 6296
rect 32404 6316 32456 6322
rect 32324 5914 32352 6287
rect 32404 6258 32456 6264
rect 32588 6248 32640 6254
rect 32588 6190 32640 6196
rect 32600 6089 32628 6190
rect 33048 6112 33100 6118
rect 32586 6080 32642 6089
rect 33048 6054 33100 6060
rect 32586 6015 32642 6024
rect 32312 5908 32364 5914
rect 32312 5850 32364 5856
rect 32600 5642 32628 6015
rect 33060 5778 33088 6054
rect 33244 5846 33272 6598
rect 33232 5840 33284 5846
rect 33232 5782 33284 5788
rect 33048 5772 33100 5778
rect 33048 5714 33100 5720
rect 32680 5704 32732 5710
rect 32680 5646 32732 5652
rect 32588 5636 32640 5642
rect 32588 5578 32640 5584
rect 31942 5400 31998 5409
rect 31942 5335 31998 5344
rect 31760 5092 31812 5098
rect 31760 5034 31812 5040
rect 31668 5024 31720 5030
rect 31668 4966 31720 4972
rect 31574 4720 31630 4729
rect 31574 4655 31630 4664
rect 31588 4622 31616 4655
rect 31576 4616 31628 4622
rect 31576 4558 31628 4564
rect 31680 4486 31708 4966
rect 31772 4554 31800 5034
rect 31760 4548 31812 4554
rect 31760 4490 31812 4496
rect 31668 4480 31720 4486
rect 31668 4422 31720 4428
rect 31956 4282 31984 5335
rect 32692 5302 32720 5646
rect 33324 5636 33376 5642
rect 33324 5578 33376 5584
rect 32680 5296 32732 5302
rect 32680 5238 32732 5244
rect 32692 4622 32720 5238
rect 32772 5228 32824 5234
rect 32772 5170 32824 5176
rect 32680 4616 32732 4622
rect 32680 4558 32732 4564
rect 31944 4276 31996 4282
rect 31944 4218 31996 4224
rect 31576 4072 31628 4078
rect 31576 4014 31628 4020
rect 31484 3392 31536 3398
rect 31484 3334 31536 3340
rect 31496 3097 31524 3334
rect 31482 3088 31538 3097
rect 31588 3058 31616 4014
rect 31482 3023 31538 3032
rect 31576 3052 31628 3058
rect 31496 2774 31524 3023
rect 31576 2994 31628 3000
rect 31760 2916 31812 2922
rect 31760 2858 31812 2864
rect 31496 2746 31616 2774
rect 31484 2508 31536 2514
rect 31484 2450 31536 2456
rect 31392 1692 31444 1698
rect 31392 1634 31444 1640
rect 31496 800 31524 2450
rect 31588 2446 31616 2746
rect 31576 2440 31628 2446
rect 31576 2382 31628 2388
rect 31772 800 31800 2858
rect 31956 2774 31984 4218
rect 32692 4214 32720 4558
rect 32784 4282 32812 5170
rect 32772 4276 32824 4282
rect 32772 4218 32824 4224
rect 32680 4208 32732 4214
rect 32680 4150 32732 4156
rect 32220 4140 32272 4146
rect 32220 4082 32272 4088
rect 32232 3126 32260 4082
rect 32692 3738 32720 4150
rect 32784 4146 32812 4218
rect 32864 4208 32916 4214
rect 32864 4150 32916 4156
rect 32772 4140 32824 4146
rect 32772 4082 32824 4088
rect 32680 3732 32732 3738
rect 32680 3674 32732 3680
rect 32496 3528 32548 3534
rect 32496 3470 32548 3476
rect 32508 3126 32536 3470
rect 32876 3466 32904 4150
rect 33336 3738 33364 5578
rect 33612 4842 33640 6938
rect 33876 6792 33928 6798
rect 33876 6734 33928 6740
rect 33888 6390 33916 6734
rect 34428 6724 34480 6730
rect 34428 6666 34480 6672
rect 34440 6458 34468 6666
rect 34428 6452 34480 6458
rect 34428 6394 34480 6400
rect 33876 6384 33928 6390
rect 33782 6352 33838 6361
rect 33876 6326 33928 6332
rect 34440 6322 34468 6394
rect 33782 6287 33838 6296
rect 34428 6316 34480 6322
rect 33690 5944 33746 5953
rect 33796 5914 33824 6287
rect 34428 6258 34480 6264
rect 33690 5879 33746 5888
rect 33784 5908 33836 5914
rect 33704 5030 33732 5879
rect 33784 5850 33836 5856
rect 34532 5302 34560 10542
rect 34624 7410 34652 10678
rect 34796 10464 34848 10470
rect 34796 10406 34848 10412
rect 34612 7404 34664 7410
rect 34612 7346 34664 7352
rect 34704 7404 34756 7410
rect 34704 7346 34756 7352
rect 34716 6662 34744 7346
rect 34808 7018 34836 10406
rect 34980 9580 35032 9586
rect 34980 9522 35032 9528
rect 35072 9580 35124 9586
rect 35072 9522 35124 9528
rect 34888 9036 34940 9042
rect 34888 8978 34940 8984
rect 34900 7818 34928 8978
rect 34888 7812 34940 7818
rect 34888 7754 34940 7760
rect 34900 7206 34928 7754
rect 34992 7546 35020 9522
rect 35084 8634 35112 9522
rect 35072 8628 35124 8634
rect 35072 8570 35124 8576
rect 35072 8492 35124 8498
rect 35072 8434 35124 8440
rect 35084 8090 35112 8434
rect 35072 8084 35124 8090
rect 35072 8026 35124 8032
rect 34980 7540 35032 7546
rect 34980 7482 35032 7488
rect 34888 7200 34940 7206
rect 34888 7142 34940 7148
rect 34808 6990 34928 7018
rect 34704 6656 34756 6662
rect 34704 6598 34756 6604
rect 34900 6458 34928 6990
rect 34888 6452 34940 6458
rect 34888 6394 34940 6400
rect 34612 6316 34664 6322
rect 34612 6258 34664 6264
rect 34624 5914 34652 6258
rect 34900 6254 34928 6394
rect 34888 6248 34940 6254
rect 35176 6202 35204 11018
rect 35256 10736 35308 10742
rect 35256 10678 35308 10684
rect 35268 10198 35296 10678
rect 36084 10464 36136 10470
rect 36084 10406 36136 10412
rect 35256 10192 35308 10198
rect 35256 10134 35308 10140
rect 35530 9208 35586 9217
rect 35530 9143 35532 9152
rect 35584 9143 35586 9152
rect 35532 9114 35584 9120
rect 35256 8968 35308 8974
rect 35256 8910 35308 8916
rect 35268 8566 35296 8910
rect 35256 8560 35308 8566
rect 35256 8502 35308 8508
rect 35268 7886 35296 8502
rect 35544 8430 35572 9114
rect 35532 8424 35584 8430
rect 35532 8366 35584 8372
rect 35256 7880 35308 7886
rect 35256 7822 35308 7828
rect 35992 7472 36044 7478
rect 35992 7414 36044 7420
rect 35256 7336 35308 7342
rect 35308 7296 35388 7324
rect 35256 7278 35308 7284
rect 34888 6190 34940 6196
rect 34612 5908 34664 5914
rect 34612 5850 34664 5856
rect 34900 5710 34928 6190
rect 35084 6174 35204 6202
rect 34888 5704 34940 5710
rect 34888 5646 34940 5652
rect 34796 5568 34848 5574
rect 34900 5556 34928 5646
rect 34848 5528 34928 5556
rect 34796 5510 34848 5516
rect 34796 5364 34848 5370
rect 34796 5306 34848 5312
rect 34520 5296 34572 5302
rect 34150 5264 34206 5273
rect 34520 5238 34572 5244
rect 34150 5199 34206 5208
rect 33784 5160 33836 5166
rect 33784 5102 33836 5108
rect 33692 5024 33744 5030
rect 33692 4966 33744 4972
rect 33416 4820 33468 4826
rect 33612 4814 33732 4842
rect 33416 4762 33468 4768
rect 33324 3732 33376 3738
rect 33324 3674 33376 3680
rect 33140 3528 33192 3534
rect 33140 3470 33192 3476
rect 32864 3460 32916 3466
rect 32864 3402 32916 3408
rect 32220 3120 32272 3126
rect 32220 3062 32272 3068
rect 32496 3120 32548 3126
rect 32496 3062 32548 3068
rect 32312 2984 32364 2990
rect 32312 2926 32364 2932
rect 31956 2746 32076 2774
rect 32048 2582 32076 2746
rect 32036 2576 32088 2582
rect 32036 2518 32088 2524
rect 32036 2100 32088 2106
rect 32036 2042 32088 2048
rect 32048 800 32076 2042
rect 32324 800 32352 2926
rect 32864 2576 32916 2582
rect 32864 2518 32916 2524
rect 32588 2304 32640 2310
rect 32588 2246 32640 2252
rect 32600 800 32628 2246
rect 32876 800 32904 2518
rect 33152 800 33180 3470
rect 33232 2440 33284 2446
rect 33232 2382 33284 2388
rect 33244 2038 33272 2382
rect 33324 2372 33376 2378
rect 33324 2314 33376 2320
rect 33336 2106 33364 2314
rect 33324 2100 33376 2106
rect 33324 2042 33376 2048
rect 33232 2032 33284 2038
rect 33232 1974 33284 1980
rect 33428 800 33456 4762
rect 33600 4072 33652 4078
rect 33600 4014 33652 4020
rect 33508 3936 33560 3942
rect 33508 3878 33560 3884
rect 33520 3398 33548 3878
rect 33508 3392 33560 3398
rect 33508 3334 33560 3340
rect 33520 2650 33548 3334
rect 33508 2644 33560 2650
rect 33508 2586 33560 2592
rect 33612 2446 33640 4014
rect 33704 2530 33732 4814
rect 33796 3194 33824 5102
rect 34164 4758 34192 5199
rect 34532 5001 34560 5238
rect 34518 4992 34574 5001
rect 34518 4927 34574 4936
rect 34152 4752 34204 4758
rect 34152 4694 34204 4700
rect 34164 4185 34192 4694
rect 34150 4176 34206 4185
rect 34150 4111 34206 4120
rect 34612 4140 34664 4146
rect 34612 4082 34664 4088
rect 34428 4072 34480 4078
rect 34428 4014 34480 4020
rect 34060 4004 34112 4010
rect 34060 3946 34112 3952
rect 33784 3188 33836 3194
rect 33784 3130 33836 3136
rect 33968 2848 34020 2854
rect 33968 2790 34020 2796
rect 33980 2650 34008 2790
rect 33968 2644 34020 2650
rect 33968 2586 34020 2592
rect 33704 2502 33824 2530
rect 33600 2440 33652 2446
rect 33600 2382 33652 2388
rect 33692 2440 33744 2446
rect 33692 2382 33744 2388
rect 33704 800 33732 2382
rect 33796 1222 33824 2502
rect 34072 1986 34100 3946
rect 34440 3534 34468 4014
rect 34624 3670 34652 4082
rect 34808 3738 34836 5306
rect 35084 4146 35112 6174
rect 35164 6112 35216 6118
rect 35164 6054 35216 6060
rect 35176 5624 35204 6054
rect 35360 5710 35388 7296
rect 35900 7200 35952 7206
rect 35900 7142 35952 7148
rect 35806 6896 35862 6905
rect 35806 6831 35808 6840
rect 35860 6831 35862 6840
rect 35808 6802 35860 6808
rect 35808 6656 35860 6662
rect 35808 6598 35860 6604
rect 35820 6322 35848 6598
rect 35912 6322 35940 7142
rect 36004 6662 36032 7414
rect 35992 6656 36044 6662
rect 35992 6598 36044 6604
rect 35808 6316 35860 6322
rect 35808 6258 35860 6264
rect 35900 6316 35952 6322
rect 35900 6258 35952 6264
rect 35820 6202 35848 6258
rect 35820 6186 35940 6202
rect 36096 6186 36124 10406
rect 36188 9926 36216 11018
rect 36556 10810 36584 11630
rect 36636 11212 36688 11218
rect 36636 11154 36688 11160
rect 36648 11082 36676 11154
rect 36636 11076 36688 11082
rect 36636 11018 36688 11024
rect 36544 10804 36596 10810
rect 36544 10746 36596 10752
rect 36556 10062 36584 10746
rect 36544 10056 36596 10062
rect 36544 9998 36596 10004
rect 36176 9920 36228 9926
rect 36176 9862 36228 9868
rect 36360 9920 36412 9926
rect 36360 9862 36412 9868
rect 36188 9738 36216 9862
rect 36188 9710 36308 9738
rect 36280 8974 36308 9710
rect 36372 9110 36400 9862
rect 36452 9580 36504 9586
rect 36452 9522 36504 9528
rect 36464 9110 36492 9522
rect 36360 9104 36412 9110
rect 36360 9046 36412 9052
rect 36452 9104 36504 9110
rect 36452 9046 36504 9052
rect 36268 8968 36320 8974
rect 36268 8910 36320 8916
rect 36176 8900 36228 8906
rect 36176 8842 36228 8848
rect 36188 7954 36216 8842
rect 36280 8498 36308 8910
rect 36372 8498 36400 9046
rect 36268 8492 36320 8498
rect 36268 8434 36320 8440
rect 36360 8492 36412 8498
rect 36360 8434 36412 8440
rect 36176 7948 36228 7954
rect 36176 7890 36228 7896
rect 36648 7886 36676 11018
rect 36636 7880 36688 7886
rect 36636 7822 36688 7828
rect 36360 7472 36412 7478
rect 36360 7414 36412 7420
rect 36176 7200 36228 7206
rect 36176 7142 36228 7148
rect 36188 7002 36216 7142
rect 36372 7002 36400 7414
rect 36648 7274 36676 7822
rect 36832 7342 36860 12038
rect 44294 11996 44602 12005
rect 44294 11994 44300 11996
rect 44356 11994 44380 11996
rect 44436 11994 44460 11996
rect 44516 11994 44540 11996
rect 44596 11994 44602 11996
rect 44356 11942 44358 11994
rect 44538 11942 44540 11994
rect 44294 11940 44300 11942
rect 44356 11940 44380 11942
rect 44436 11940 44460 11942
rect 44516 11940 44540 11942
rect 44596 11940 44602 11942
rect 44294 11931 44602 11940
rect 45652 11756 45704 11762
rect 45652 11698 45704 11704
rect 41788 11620 41840 11626
rect 41788 11562 41840 11568
rect 37648 11552 37700 11558
rect 37648 11494 37700 11500
rect 38384 11552 38436 11558
rect 38384 11494 38436 11500
rect 37070 11452 37378 11461
rect 37070 11450 37076 11452
rect 37132 11450 37156 11452
rect 37212 11450 37236 11452
rect 37292 11450 37316 11452
rect 37372 11450 37378 11452
rect 37132 11398 37134 11450
rect 37314 11398 37316 11450
rect 37070 11396 37076 11398
rect 37132 11396 37156 11398
rect 37212 11396 37236 11398
rect 37292 11396 37316 11398
rect 37372 11396 37378 11398
rect 37070 11387 37378 11396
rect 36912 11008 36964 11014
rect 36912 10950 36964 10956
rect 36924 10606 36952 10950
rect 37464 10804 37516 10810
rect 37464 10746 37516 10752
rect 36912 10600 36964 10606
rect 36912 10542 36964 10548
rect 36924 9926 36952 10542
rect 37070 10364 37378 10373
rect 37070 10362 37076 10364
rect 37132 10362 37156 10364
rect 37212 10362 37236 10364
rect 37292 10362 37316 10364
rect 37372 10362 37378 10364
rect 37132 10310 37134 10362
rect 37314 10310 37316 10362
rect 37070 10308 37076 10310
rect 37132 10308 37156 10310
rect 37212 10308 37236 10310
rect 37292 10308 37316 10310
rect 37372 10308 37378 10310
rect 37070 10299 37378 10308
rect 36912 9920 36964 9926
rect 36912 9862 36964 9868
rect 37372 9920 37424 9926
rect 37372 9862 37424 9868
rect 37384 9722 37412 9862
rect 37372 9716 37424 9722
rect 37372 9658 37424 9664
rect 37384 9518 37412 9658
rect 37372 9512 37424 9518
rect 37372 9454 37424 9460
rect 37070 9276 37378 9285
rect 37070 9274 37076 9276
rect 37132 9274 37156 9276
rect 37212 9274 37236 9276
rect 37292 9274 37316 9276
rect 37372 9274 37378 9276
rect 37132 9222 37134 9274
rect 37314 9222 37316 9274
rect 37070 9220 37076 9222
rect 37132 9220 37156 9222
rect 37212 9220 37236 9222
rect 37292 9220 37316 9222
rect 37372 9220 37378 9222
rect 37070 9211 37378 9220
rect 37476 8974 37504 10746
rect 37556 10464 37608 10470
rect 37556 10406 37608 10412
rect 37568 9178 37596 10406
rect 37556 9172 37608 9178
rect 37556 9114 37608 9120
rect 37464 8968 37516 8974
rect 37464 8910 37516 8916
rect 36912 8832 36964 8838
rect 36912 8774 36964 8780
rect 36924 7886 36952 8774
rect 37556 8424 37608 8430
rect 37556 8366 37608 8372
rect 37070 8188 37378 8197
rect 37070 8186 37076 8188
rect 37132 8186 37156 8188
rect 37212 8186 37236 8188
rect 37292 8186 37316 8188
rect 37372 8186 37378 8188
rect 37132 8134 37134 8186
rect 37314 8134 37316 8186
rect 37070 8132 37076 8134
rect 37132 8132 37156 8134
rect 37212 8132 37236 8134
rect 37292 8132 37316 8134
rect 37372 8132 37378 8134
rect 37070 8123 37378 8132
rect 36912 7880 36964 7886
rect 36912 7822 36964 7828
rect 37464 7744 37516 7750
rect 37464 7686 37516 7692
rect 37476 7410 37504 7686
rect 37568 7410 37596 8366
rect 37464 7404 37516 7410
rect 37464 7346 37516 7352
rect 37556 7404 37608 7410
rect 37556 7346 37608 7352
rect 36820 7336 36872 7342
rect 36820 7278 36872 7284
rect 36636 7268 36688 7274
rect 36636 7210 36688 7216
rect 36912 7200 36964 7206
rect 36912 7142 36964 7148
rect 37464 7200 37516 7206
rect 37464 7142 37516 7148
rect 36924 7018 36952 7142
rect 37070 7100 37378 7109
rect 37070 7098 37076 7100
rect 37132 7098 37156 7100
rect 37212 7098 37236 7100
rect 37292 7098 37316 7100
rect 37372 7098 37378 7100
rect 37132 7046 37134 7098
rect 37314 7046 37316 7098
rect 37070 7044 37076 7046
rect 37132 7044 37156 7046
rect 37212 7044 37236 7046
rect 37292 7044 37316 7046
rect 37372 7044 37378 7046
rect 37070 7035 37378 7044
rect 36176 6996 36228 7002
rect 36176 6938 36228 6944
rect 36360 6996 36412 7002
rect 36924 6990 37044 7018
rect 36360 6938 36412 6944
rect 37016 6916 37044 6990
rect 37016 6888 37228 6916
rect 37200 6882 37228 6888
rect 37200 6854 37320 6882
rect 37292 6798 37320 6854
rect 36820 6792 36872 6798
rect 36820 6734 36872 6740
rect 37096 6792 37148 6798
rect 37096 6734 37148 6740
rect 37280 6792 37332 6798
rect 37280 6734 37332 6740
rect 36832 6662 36860 6734
rect 36820 6656 36872 6662
rect 36820 6598 36872 6604
rect 35820 6180 35952 6186
rect 35820 6174 35900 6180
rect 35900 6122 35952 6128
rect 36084 6180 36136 6186
rect 36084 6122 36136 6128
rect 35348 5704 35400 5710
rect 35348 5646 35400 5652
rect 35912 5642 35940 6122
rect 36832 5914 36860 6598
rect 37004 6452 37056 6458
rect 37004 6394 37056 6400
rect 37016 6186 37044 6394
rect 37108 6225 37136 6734
rect 37476 6730 37504 7142
rect 37660 7002 37688 11494
rect 38396 11354 38424 11494
rect 38384 11348 38436 11354
rect 38384 11290 38436 11296
rect 41144 11348 41196 11354
rect 41144 11290 41196 11296
rect 38752 11280 38804 11286
rect 38752 11222 38804 11228
rect 39488 11280 39540 11286
rect 39488 11222 39540 11228
rect 38660 11144 38712 11150
rect 38660 11086 38712 11092
rect 38200 11008 38252 11014
rect 38200 10950 38252 10956
rect 38568 11008 38620 11014
rect 38568 10950 38620 10956
rect 38212 10538 38240 10950
rect 38580 10810 38608 10950
rect 38568 10804 38620 10810
rect 38568 10746 38620 10752
rect 38672 10674 38700 11086
rect 38660 10668 38712 10674
rect 38660 10610 38712 10616
rect 38200 10532 38252 10538
rect 38200 10474 38252 10480
rect 38108 10056 38160 10062
rect 38108 9998 38160 10004
rect 38016 9988 38068 9994
rect 38016 9930 38068 9936
rect 38028 9722 38056 9930
rect 38120 9722 38148 9998
rect 38016 9716 38068 9722
rect 38016 9658 38068 9664
rect 38108 9716 38160 9722
rect 38108 9658 38160 9664
rect 38212 9602 38240 10474
rect 38672 10198 38700 10610
rect 38660 10192 38712 10198
rect 38660 10134 38712 10140
rect 38672 9654 38700 10134
rect 38120 9574 38240 9602
rect 38660 9648 38712 9654
rect 38660 9590 38712 9596
rect 38568 9580 38620 9586
rect 38120 9450 38148 9574
rect 38568 9522 38620 9528
rect 38108 9444 38160 9450
rect 38108 9386 38160 9392
rect 37832 8832 37884 8838
rect 37832 8774 37884 8780
rect 37844 8498 37872 8774
rect 38120 8498 38148 9386
rect 38580 9178 38608 9522
rect 38764 9178 38792 11222
rect 39500 10810 39528 11222
rect 40408 11076 40460 11082
rect 40408 11018 40460 11024
rect 39488 10804 39540 10810
rect 39488 10746 39540 10752
rect 39856 10464 39908 10470
rect 39856 10406 39908 10412
rect 39764 9920 39816 9926
rect 39764 9862 39816 9868
rect 38844 9376 38896 9382
rect 38844 9318 38896 9324
rect 38568 9172 38620 9178
rect 38568 9114 38620 9120
rect 38752 9172 38804 9178
rect 38752 9114 38804 9120
rect 38764 8498 38792 9114
rect 38856 9110 38884 9318
rect 39776 9110 39804 9862
rect 38844 9104 38896 9110
rect 38844 9046 38896 9052
rect 39764 9104 39816 9110
rect 39764 9046 39816 9052
rect 37832 8492 37884 8498
rect 37832 8434 37884 8440
rect 38108 8492 38160 8498
rect 38108 8434 38160 8440
rect 38752 8492 38804 8498
rect 38752 8434 38804 8440
rect 38120 7818 38148 8434
rect 38384 8356 38436 8362
rect 38384 8298 38436 8304
rect 38108 7812 38160 7818
rect 38108 7754 38160 7760
rect 37924 7336 37976 7342
rect 37924 7278 37976 7284
rect 37740 7268 37792 7274
rect 37740 7210 37792 7216
rect 37752 7002 37780 7210
rect 37648 6996 37700 7002
rect 37648 6938 37700 6944
rect 37740 6996 37792 7002
rect 37740 6938 37792 6944
rect 37464 6724 37516 6730
rect 37464 6666 37516 6672
rect 37094 6216 37150 6225
rect 36912 6180 36964 6186
rect 36912 6122 36964 6128
rect 37004 6180 37056 6186
rect 37094 6151 37150 6160
rect 37004 6122 37056 6128
rect 36924 5914 36952 6122
rect 37070 6012 37378 6021
rect 37070 6010 37076 6012
rect 37132 6010 37156 6012
rect 37212 6010 37236 6012
rect 37292 6010 37316 6012
rect 37372 6010 37378 6012
rect 37132 5958 37134 6010
rect 37314 5958 37316 6010
rect 37070 5956 37076 5958
rect 37132 5956 37156 5958
rect 37212 5956 37236 5958
rect 37292 5956 37316 5958
rect 37372 5956 37378 5958
rect 37070 5947 37378 5956
rect 36820 5908 36872 5914
rect 36820 5850 36872 5856
rect 36912 5908 36964 5914
rect 36912 5850 36964 5856
rect 37660 5846 37688 6938
rect 37740 6316 37792 6322
rect 37740 6258 37792 6264
rect 36084 5840 36136 5846
rect 37648 5840 37700 5846
rect 36136 5788 36216 5794
rect 36084 5782 36216 5788
rect 37648 5782 37700 5788
rect 36096 5766 36216 5782
rect 36188 5760 36216 5766
rect 36452 5772 36504 5778
rect 36188 5732 36452 5760
rect 36452 5714 36504 5720
rect 36084 5704 36136 5710
rect 36084 5646 36136 5652
rect 36358 5672 36414 5681
rect 35900 5636 35952 5642
rect 35176 5596 35296 5624
rect 35268 5166 35296 5596
rect 35900 5578 35952 5584
rect 36096 5234 36124 5646
rect 36358 5607 36414 5616
rect 36084 5228 36136 5234
rect 36084 5170 36136 5176
rect 35256 5160 35308 5166
rect 35256 5102 35308 5108
rect 35624 5024 35676 5030
rect 35624 4966 35676 4972
rect 35440 4616 35492 4622
rect 35440 4558 35492 4564
rect 35072 4140 35124 4146
rect 35072 4082 35124 4088
rect 34796 3732 34848 3738
rect 34796 3674 34848 3680
rect 35256 3732 35308 3738
rect 35256 3674 35308 3680
rect 34612 3664 34664 3670
rect 34612 3606 34664 3612
rect 34428 3528 34480 3534
rect 34428 3470 34480 3476
rect 34520 3120 34572 3126
rect 34520 3062 34572 3068
rect 34244 2848 34296 2854
rect 34244 2790 34296 2796
rect 33980 1958 34100 1986
rect 33784 1216 33836 1222
rect 33784 1158 33836 1164
rect 33980 800 34008 1958
rect 34256 800 34284 2790
rect 34532 800 34560 3062
rect 34624 2553 34652 3606
rect 34808 3058 34836 3674
rect 34886 3632 34942 3641
rect 34886 3567 34942 3576
rect 34900 3534 34928 3567
rect 34888 3528 34940 3534
rect 34888 3470 34940 3476
rect 34900 3194 34928 3470
rect 34888 3188 34940 3194
rect 34888 3130 34940 3136
rect 34796 3052 34848 3058
rect 34796 2994 34848 3000
rect 34610 2544 34666 2553
rect 34610 2479 34666 2488
rect 35072 2100 35124 2106
rect 35072 2042 35124 2048
rect 34796 1964 34848 1970
rect 34796 1906 34848 1912
rect 34808 800 34836 1906
rect 35084 800 35112 2042
rect 35268 1578 35296 3674
rect 35348 2916 35400 2922
rect 35348 2858 35400 2864
rect 35360 2650 35388 2858
rect 35348 2644 35400 2650
rect 35348 2586 35400 2592
rect 35268 1550 35388 1578
rect 35360 800 35388 1550
rect 35452 1086 35480 4558
rect 35532 4480 35584 4486
rect 35532 4422 35584 4428
rect 35544 3534 35572 4422
rect 35532 3528 35584 3534
rect 35532 3470 35584 3476
rect 35532 3120 35584 3126
rect 35532 3062 35584 3068
rect 35544 2854 35572 3062
rect 35532 2848 35584 2854
rect 35532 2790 35584 2796
rect 35440 1080 35492 1086
rect 35440 1022 35492 1028
rect 35636 800 35664 4966
rect 36096 4826 36124 5170
rect 36084 4820 36136 4826
rect 36084 4762 36136 4768
rect 35716 4752 35768 4758
rect 35716 4694 35768 4700
rect 35728 4146 35756 4694
rect 36084 4684 36136 4690
rect 36136 4644 36216 4672
rect 36084 4626 36136 4632
rect 35806 4448 35862 4457
rect 35806 4383 35862 4392
rect 35820 4214 35848 4383
rect 35808 4208 35860 4214
rect 35808 4150 35860 4156
rect 35716 4140 35768 4146
rect 35716 4082 35768 4088
rect 35728 3913 35756 4082
rect 36188 3942 36216 4644
rect 35900 3936 35952 3942
rect 35714 3904 35770 3913
rect 35900 3878 35952 3884
rect 35992 3936 36044 3942
rect 35992 3878 36044 3884
rect 36176 3936 36228 3942
rect 36176 3878 36228 3884
rect 35714 3839 35770 3848
rect 35728 2281 35756 3839
rect 35912 3466 35940 3878
rect 35900 3460 35952 3466
rect 35900 3402 35952 3408
rect 36004 3210 36032 3878
rect 35912 3182 36032 3210
rect 35912 3074 35940 3182
rect 35820 3046 35940 3074
rect 35820 2990 35848 3046
rect 35808 2984 35860 2990
rect 35808 2926 35860 2932
rect 35900 2984 35952 2990
rect 35900 2926 35952 2932
rect 35714 2272 35770 2281
rect 35714 2207 35770 2216
rect 35912 800 35940 2926
rect 36372 1465 36400 5607
rect 37752 5574 37780 6258
rect 37936 6225 37964 7278
rect 38108 7268 38160 7274
rect 38108 7210 38160 7216
rect 38120 6361 38148 7210
rect 38290 6896 38346 6905
rect 38290 6831 38346 6840
rect 38106 6352 38162 6361
rect 38106 6287 38162 6296
rect 38304 6254 38332 6831
rect 38396 6798 38424 8298
rect 38660 7404 38712 7410
rect 38660 7346 38712 7352
rect 38384 6792 38436 6798
rect 38384 6734 38436 6740
rect 38476 6792 38528 6798
rect 38476 6734 38528 6740
rect 38488 6390 38516 6734
rect 38672 6662 38700 7346
rect 38764 7290 38792 8434
rect 38856 7886 38884 9046
rect 39672 8968 39724 8974
rect 39672 8910 39724 8916
rect 39028 8900 39080 8906
rect 39028 8842 39080 8848
rect 39040 8634 39068 8842
rect 39684 8634 39712 8910
rect 39028 8628 39080 8634
rect 39028 8570 39080 8576
rect 39672 8628 39724 8634
rect 39672 8570 39724 8576
rect 39488 8492 39540 8498
rect 39488 8434 39540 8440
rect 39500 8022 39528 8434
rect 39488 8016 39540 8022
rect 39488 7958 39540 7964
rect 38844 7880 38896 7886
rect 38844 7822 38896 7828
rect 38936 7472 38988 7478
rect 38936 7414 38988 7420
rect 38948 7342 38976 7414
rect 38936 7336 38988 7342
rect 38764 7262 38884 7290
rect 38936 7278 38988 7284
rect 38752 7200 38804 7206
rect 38752 7142 38804 7148
rect 38764 6866 38792 7142
rect 38856 6866 38884 7262
rect 38752 6860 38804 6866
rect 38752 6802 38804 6808
rect 38844 6860 38896 6866
rect 38844 6802 38896 6808
rect 38948 6730 38976 7278
rect 38936 6724 38988 6730
rect 38936 6666 38988 6672
rect 38660 6656 38712 6662
rect 38660 6598 38712 6604
rect 39304 6656 39356 6662
rect 39304 6598 39356 6604
rect 38476 6384 38528 6390
rect 38476 6326 38528 6332
rect 38660 6316 38712 6322
rect 38660 6258 38712 6264
rect 38292 6248 38344 6254
rect 37922 6216 37978 6225
rect 38292 6190 38344 6196
rect 37922 6151 37978 6160
rect 38016 6180 38068 6186
rect 37740 5568 37792 5574
rect 37740 5510 37792 5516
rect 36912 5160 36964 5166
rect 36912 5102 36964 5108
rect 36924 4690 36952 5102
rect 37740 5024 37792 5030
rect 37740 4966 37792 4972
rect 37070 4924 37378 4933
rect 37070 4922 37076 4924
rect 37132 4922 37156 4924
rect 37212 4922 37236 4924
rect 37292 4922 37316 4924
rect 37372 4922 37378 4924
rect 37132 4870 37134 4922
rect 37314 4870 37316 4922
rect 37070 4868 37076 4870
rect 37132 4868 37156 4870
rect 37212 4868 37236 4870
rect 37292 4868 37316 4870
rect 37372 4868 37378 4870
rect 37070 4859 37378 4868
rect 36912 4684 36964 4690
rect 36912 4626 36964 4632
rect 36820 4072 36872 4078
rect 36820 4014 36872 4020
rect 36728 3528 36780 3534
rect 36728 3470 36780 3476
rect 36740 3233 36768 3470
rect 36726 3224 36782 3233
rect 36832 3194 36860 4014
rect 36726 3159 36728 3168
rect 36780 3159 36782 3168
rect 36820 3188 36872 3194
rect 36728 3130 36780 3136
rect 36820 3130 36872 3136
rect 36820 3052 36872 3058
rect 36820 2994 36872 3000
rect 36452 2576 36504 2582
rect 36452 2518 36504 2524
rect 36358 1456 36414 1465
rect 36176 1420 36228 1426
rect 36358 1391 36414 1400
rect 36176 1362 36228 1368
rect 36188 800 36216 1362
rect 36464 800 36492 2518
rect 36728 2032 36780 2038
rect 36728 1974 36780 1980
rect 36740 800 36768 1974
rect 36832 1442 36860 2994
rect 36924 2650 36952 4626
rect 37280 4548 37332 4554
rect 37280 4490 37332 4496
rect 37292 4282 37320 4490
rect 37280 4276 37332 4282
rect 37280 4218 37332 4224
rect 37752 4146 37780 4966
rect 37936 4486 37964 6151
rect 38016 6122 38068 6128
rect 38028 5846 38056 6122
rect 38016 5840 38068 5846
rect 38016 5782 38068 5788
rect 38568 5704 38620 5710
rect 38568 5646 38620 5652
rect 38580 5302 38608 5646
rect 38672 5370 38700 6258
rect 39316 6254 39344 6598
rect 39304 6248 39356 6254
rect 39304 6190 39356 6196
rect 39120 5568 39172 5574
rect 39120 5510 39172 5516
rect 38660 5364 38712 5370
rect 38660 5306 38712 5312
rect 38568 5296 38620 5302
rect 38568 5238 38620 5244
rect 38752 5228 38804 5234
rect 38752 5170 38804 5176
rect 39028 5228 39080 5234
rect 39028 5170 39080 5176
rect 38764 4758 38792 5170
rect 38752 4752 38804 4758
rect 39040 4729 39068 5170
rect 38752 4694 38804 4700
rect 39026 4720 39082 4729
rect 39026 4655 39082 4664
rect 38660 4616 38712 4622
rect 38660 4558 38712 4564
rect 37924 4480 37976 4486
rect 37924 4422 37976 4428
rect 37936 4146 37964 4422
rect 38106 4312 38162 4321
rect 38106 4247 38162 4256
rect 37464 4140 37516 4146
rect 37464 4082 37516 4088
rect 37740 4140 37792 4146
rect 37740 4082 37792 4088
rect 37924 4140 37976 4146
rect 37924 4082 37976 4088
rect 37070 3836 37378 3845
rect 37070 3834 37076 3836
rect 37132 3834 37156 3836
rect 37212 3834 37236 3836
rect 37292 3834 37316 3836
rect 37372 3834 37378 3836
rect 37132 3782 37134 3834
rect 37314 3782 37316 3834
rect 37070 3780 37076 3782
rect 37132 3780 37156 3782
rect 37212 3780 37236 3782
rect 37292 3780 37316 3782
rect 37372 3780 37378 3782
rect 37070 3771 37378 3780
rect 37476 3777 37504 4082
rect 37462 3768 37518 3777
rect 37462 3703 37518 3712
rect 37556 3732 37608 3738
rect 37476 3618 37504 3703
rect 37556 3674 37608 3680
rect 37384 3590 37504 3618
rect 37384 3369 37412 3590
rect 37464 3392 37516 3398
rect 37370 3360 37426 3369
rect 37464 3334 37516 3340
rect 37370 3295 37426 3304
rect 37476 3058 37504 3334
rect 37464 3052 37516 3058
rect 37464 2994 37516 3000
rect 37070 2748 37378 2757
rect 37070 2746 37076 2748
rect 37132 2746 37156 2748
rect 37212 2746 37236 2748
rect 37292 2746 37316 2748
rect 37372 2746 37378 2748
rect 37132 2694 37134 2746
rect 37314 2694 37316 2746
rect 37070 2692 37076 2694
rect 37132 2692 37156 2694
rect 37212 2692 37236 2694
rect 37292 2692 37316 2694
rect 37372 2692 37378 2694
rect 37070 2683 37378 2692
rect 36912 2644 36964 2650
rect 36912 2586 36964 2592
rect 37096 2644 37148 2650
rect 37096 2586 37148 2592
rect 36832 1414 37044 1442
rect 37108 1426 37136 2586
rect 37280 1488 37332 1494
rect 37280 1430 37332 1436
rect 37016 800 37044 1414
rect 37096 1420 37148 1426
rect 37096 1362 37148 1368
rect 37292 800 37320 1430
rect 37568 800 37596 3674
rect 37648 3596 37700 3602
rect 37648 3538 37700 3544
rect 37660 3058 37688 3538
rect 37738 3088 37794 3097
rect 37648 3052 37700 3058
rect 37738 3023 37740 3032
rect 37648 2994 37700 3000
rect 37792 3023 37794 3032
rect 37740 2994 37792 3000
rect 37660 1970 37688 2994
rect 37752 2825 37780 2994
rect 37738 2816 37794 2825
rect 37738 2751 37794 2760
rect 38016 2372 38068 2378
rect 38016 2314 38068 2320
rect 37648 1964 37700 1970
rect 37648 1906 37700 1912
rect 38028 1306 38056 2314
rect 37844 1278 38056 1306
rect 37844 800 37872 1278
rect 38120 800 38148 4247
rect 38672 3738 38700 4558
rect 39040 4146 39068 4655
rect 39028 4140 39080 4146
rect 39028 4082 39080 4088
rect 39132 3913 39160 5510
rect 39672 5228 39724 5234
rect 39672 5170 39724 5176
rect 39684 4826 39712 5170
rect 39672 4820 39724 4826
rect 39672 4762 39724 4768
rect 39868 4146 39896 10406
rect 40224 10056 40276 10062
rect 40224 9998 40276 10004
rect 40236 9586 40264 9998
rect 39948 9580 40000 9586
rect 39948 9522 40000 9528
rect 40224 9580 40276 9586
rect 40224 9522 40276 9528
rect 40316 9580 40368 9586
rect 40316 9522 40368 9528
rect 39960 8634 39988 9522
rect 40132 9036 40184 9042
rect 40132 8978 40184 8984
rect 40144 8838 40172 8978
rect 40328 8974 40356 9522
rect 40316 8968 40368 8974
rect 40316 8910 40368 8916
rect 40132 8832 40184 8838
rect 40132 8774 40184 8780
rect 40316 8832 40368 8838
rect 40316 8774 40368 8780
rect 39948 8628 40000 8634
rect 39948 8570 40000 8576
rect 40328 8498 40356 8774
rect 40316 8492 40368 8498
rect 40316 8434 40368 8440
rect 40224 8288 40276 8294
rect 40224 8230 40276 8236
rect 40236 8022 40264 8230
rect 40224 8016 40276 8022
rect 40420 7970 40448 11018
rect 41156 10810 41184 11290
rect 41800 10810 41828 11562
rect 43076 11552 43128 11558
rect 43076 11494 43128 11500
rect 43536 11552 43588 11558
rect 43536 11494 43588 11500
rect 41972 11076 42024 11082
rect 41972 11018 42024 11024
rect 42892 11076 42944 11082
rect 42892 11018 42944 11024
rect 41144 10804 41196 10810
rect 41144 10746 41196 10752
rect 41788 10804 41840 10810
rect 41788 10746 41840 10752
rect 41236 10532 41288 10538
rect 41236 10474 41288 10480
rect 40500 10464 40552 10470
rect 40500 10406 40552 10412
rect 40224 7958 40276 7964
rect 40328 7942 40448 7970
rect 40224 7744 40276 7750
rect 40224 7686 40276 7692
rect 39946 7440 40002 7449
rect 39946 7375 40002 7384
rect 39960 6882 39988 7375
rect 39960 6866 40080 6882
rect 39960 6860 40092 6866
rect 39960 6854 40040 6860
rect 40040 6802 40092 6808
rect 40236 6322 40264 7686
rect 40224 6316 40276 6322
rect 40224 6258 40276 6264
rect 40040 6248 40092 6254
rect 40040 6190 40092 6196
rect 40052 5778 40080 6190
rect 40132 6180 40184 6186
rect 40132 6122 40184 6128
rect 40144 5846 40172 6122
rect 40132 5840 40184 5846
rect 40132 5782 40184 5788
rect 40040 5772 40092 5778
rect 40040 5714 40092 5720
rect 40052 5302 40080 5714
rect 40040 5296 40092 5302
rect 40040 5238 40092 5244
rect 40222 5128 40278 5137
rect 40328 5114 40356 7942
rect 40408 7812 40460 7818
rect 40408 7754 40460 7760
rect 40420 6730 40448 7754
rect 40408 6724 40460 6730
rect 40408 6666 40460 6672
rect 40512 6610 40540 10406
rect 41248 9994 41276 10474
rect 41236 9988 41288 9994
rect 41236 9930 41288 9936
rect 41248 9518 41276 9930
rect 41236 9512 41288 9518
rect 41236 9454 41288 9460
rect 41328 8968 41380 8974
rect 41328 8910 41380 8916
rect 41144 8832 41196 8838
rect 41144 8774 41196 8780
rect 40776 8628 40828 8634
rect 40776 8570 40828 8576
rect 40788 8430 40816 8570
rect 41156 8498 41184 8774
rect 41144 8492 41196 8498
rect 41144 8434 41196 8440
rect 40776 8424 40828 8430
rect 40776 8366 40828 8372
rect 40592 7880 40644 7886
rect 40592 7822 40644 7828
rect 40604 7478 40632 7822
rect 40592 7472 40644 7478
rect 40592 7414 40644 7420
rect 40684 7404 40736 7410
rect 40684 7346 40736 7352
rect 40420 6582 40540 6610
rect 40420 5710 40448 6582
rect 40696 6458 40724 7346
rect 40684 6452 40736 6458
rect 40684 6394 40736 6400
rect 40788 6118 40816 8366
rect 41340 8090 41368 8910
rect 41696 8832 41748 8838
rect 41696 8774 41748 8780
rect 41328 8084 41380 8090
rect 41328 8026 41380 8032
rect 41708 7886 41736 8774
rect 41696 7880 41748 7886
rect 41696 7822 41748 7828
rect 41420 7744 41472 7750
rect 41420 7686 41472 7692
rect 41432 7274 41460 7686
rect 41420 7268 41472 7274
rect 41420 7210 41472 7216
rect 41604 6928 41656 6934
rect 41604 6870 41656 6876
rect 40868 6724 40920 6730
rect 40868 6666 40920 6672
rect 40880 6458 40908 6666
rect 40868 6452 40920 6458
rect 40868 6394 40920 6400
rect 41616 6322 41644 6870
rect 41696 6792 41748 6798
rect 41696 6734 41748 6740
rect 41708 6322 41736 6734
rect 41800 6730 41828 10746
rect 41880 8832 41932 8838
rect 41880 8774 41932 8780
rect 41892 8294 41920 8774
rect 41880 8288 41932 8294
rect 41880 8230 41932 8236
rect 41892 7585 41920 8230
rect 41878 7576 41934 7585
rect 41878 7511 41934 7520
rect 41788 6724 41840 6730
rect 41788 6666 41840 6672
rect 41800 6390 41828 6666
rect 41984 6662 42012 11018
rect 42904 10470 42932 11018
rect 42524 10464 42576 10470
rect 42524 10406 42576 10412
rect 42892 10464 42944 10470
rect 42892 10406 42944 10412
rect 42432 10056 42484 10062
rect 42432 9998 42484 10004
rect 42156 9580 42208 9586
rect 42156 9522 42208 9528
rect 42168 9178 42196 9522
rect 42444 9518 42472 9998
rect 42432 9512 42484 9518
rect 42432 9454 42484 9460
rect 42156 9172 42208 9178
rect 42156 9114 42208 9120
rect 42444 8906 42472 9454
rect 42432 8900 42484 8906
rect 42432 8842 42484 8848
rect 42536 8430 42564 10406
rect 42800 9376 42852 9382
rect 42800 9318 42852 9324
rect 42812 9178 42840 9318
rect 42800 9172 42852 9178
rect 42800 9114 42852 9120
rect 42524 8424 42576 8430
rect 42524 8366 42576 8372
rect 42536 8090 42564 8366
rect 42524 8084 42576 8090
rect 42524 8026 42576 8032
rect 42904 7857 42932 10406
rect 42984 10056 43036 10062
rect 42984 9998 43036 10004
rect 42996 9722 43024 9998
rect 42984 9716 43036 9722
rect 42984 9658 43036 9664
rect 43088 7970 43116 11494
rect 43352 11348 43404 11354
rect 43352 11290 43404 11296
rect 43364 10810 43392 11290
rect 43352 10804 43404 10810
rect 43352 10746 43404 10752
rect 43444 8968 43496 8974
rect 43444 8910 43496 8916
rect 43456 8634 43484 8910
rect 43444 8628 43496 8634
rect 43444 8570 43496 8576
rect 43352 8492 43404 8498
rect 43352 8434 43404 8440
rect 43364 8090 43392 8434
rect 43352 8084 43404 8090
rect 43352 8026 43404 8032
rect 42996 7942 43116 7970
rect 42890 7848 42946 7857
rect 42890 7783 42892 7792
rect 42944 7783 42946 7792
rect 42892 7754 42944 7760
rect 42432 7540 42484 7546
rect 42432 7482 42484 7488
rect 42444 6798 42472 7482
rect 42904 7410 42932 7754
rect 42892 7404 42944 7410
rect 42892 7346 42944 7352
rect 42892 7200 42944 7206
rect 42892 7142 42944 7148
rect 42904 7002 42932 7142
rect 42892 6996 42944 7002
rect 42892 6938 42944 6944
rect 42432 6792 42484 6798
rect 42432 6734 42484 6740
rect 42706 6760 42762 6769
rect 41972 6656 42024 6662
rect 41972 6598 42024 6604
rect 41788 6384 41840 6390
rect 41788 6326 41840 6332
rect 41604 6316 41656 6322
rect 41604 6258 41656 6264
rect 41696 6316 41748 6322
rect 41696 6258 41748 6264
rect 41420 6248 41472 6254
rect 41420 6190 41472 6196
rect 40776 6112 40828 6118
rect 40776 6054 40828 6060
rect 41328 6112 41380 6118
rect 41328 6054 41380 6060
rect 41340 5914 41368 6054
rect 41328 5908 41380 5914
rect 41328 5850 41380 5856
rect 40408 5704 40460 5710
rect 40406 5672 40408 5681
rect 40460 5672 40462 5681
rect 41432 5642 41460 6190
rect 42444 5914 42472 6734
rect 42616 6724 42668 6730
rect 42706 6695 42762 6704
rect 42616 6666 42668 6672
rect 42628 6254 42656 6666
rect 42720 6662 42748 6695
rect 42708 6656 42760 6662
rect 42708 6598 42760 6604
rect 42616 6248 42668 6254
rect 42616 6190 42668 6196
rect 42628 6118 42656 6190
rect 42616 6112 42668 6118
rect 42616 6054 42668 6060
rect 42996 5953 43024 7942
rect 43076 7880 43128 7886
rect 43076 7822 43128 7828
rect 43088 7002 43116 7822
rect 43076 6996 43128 7002
rect 43076 6938 43128 6944
rect 43352 6724 43404 6730
rect 43352 6666 43404 6672
rect 42982 5944 43038 5953
rect 42432 5908 42484 5914
rect 42432 5850 42484 5856
rect 42812 5888 42982 5896
rect 42812 5879 43038 5888
rect 42812 5868 43024 5879
rect 42432 5704 42484 5710
rect 42432 5646 42484 5652
rect 40406 5607 40462 5616
rect 41420 5636 41472 5642
rect 41420 5578 41472 5584
rect 42444 5370 42472 5646
rect 42812 5409 42840 5868
rect 42996 5819 43024 5868
rect 43364 5574 43392 6666
rect 43352 5568 43404 5574
rect 43352 5510 43404 5516
rect 42798 5400 42854 5409
rect 42432 5364 42484 5370
rect 42798 5335 42854 5344
rect 42432 5306 42484 5312
rect 40328 5086 40540 5114
rect 40222 5063 40278 5072
rect 40236 4690 40264 5063
rect 40316 5024 40368 5030
rect 40316 4966 40368 4972
rect 40224 4684 40276 4690
rect 40224 4626 40276 4632
rect 39948 4480 40000 4486
rect 39948 4422 40000 4428
rect 39960 4185 39988 4422
rect 40328 4282 40356 4966
rect 40406 4856 40462 4865
rect 40406 4791 40462 4800
rect 40316 4276 40368 4282
rect 40316 4218 40368 4224
rect 40040 4208 40092 4214
rect 39946 4176 40002 4185
rect 39304 4140 39356 4146
rect 39304 4082 39356 4088
rect 39856 4140 39908 4146
rect 40040 4150 40092 4156
rect 39946 4111 40002 4120
rect 39856 4082 39908 4088
rect 39118 3904 39174 3913
rect 39118 3839 39174 3848
rect 38660 3732 38712 3738
rect 38660 3674 38712 3680
rect 38292 3528 38344 3534
rect 38290 3496 38292 3505
rect 38476 3528 38528 3534
rect 38344 3496 38346 3505
rect 38476 3470 38528 3476
rect 38290 3431 38346 3440
rect 38384 3460 38436 3466
rect 38384 3402 38436 3408
rect 38292 2984 38344 2990
rect 38292 2926 38344 2932
rect 38304 1494 38332 2926
rect 38292 1488 38344 1494
rect 38292 1430 38344 1436
rect 38396 800 38424 3402
rect 38488 2417 38516 3470
rect 38568 3392 38620 3398
rect 38568 3334 38620 3340
rect 38474 2408 38530 2417
rect 38474 2343 38530 2352
rect 38580 2009 38608 3334
rect 39132 3233 39160 3839
rect 39118 3224 39174 3233
rect 39118 3159 39174 3168
rect 39210 2544 39266 2553
rect 39210 2479 39212 2488
rect 39264 2479 39266 2488
rect 39212 2450 39264 2456
rect 38566 2000 38622 2009
rect 38566 1935 38622 1944
rect 38580 1601 38608 1935
rect 38660 1896 38712 1902
rect 39316 1873 39344 4082
rect 39488 3664 39540 3670
rect 39488 3606 39540 3612
rect 39500 2854 39528 3606
rect 39948 3596 40000 3602
rect 39948 3538 40000 3544
rect 39960 3194 39988 3538
rect 39948 3188 40000 3194
rect 39948 3130 40000 3136
rect 39672 2984 39724 2990
rect 39672 2926 39724 2932
rect 39684 2854 39712 2926
rect 39488 2848 39540 2854
rect 39488 2790 39540 2796
rect 39672 2848 39724 2854
rect 39672 2790 39724 2796
rect 39488 2508 39540 2514
rect 39488 2450 39540 2456
rect 38660 1838 38712 1844
rect 39302 1864 39358 1873
rect 38566 1592 38622 1601
rect 38566 1527 38622 1536
rect 38672 800 38700 1838
rect 39302 1799 39358 1808
rect 39212 1488 39264 1494
rect 39212 1430 39264 1436
rect 38936 1216 38988 1222
rect 38936 1158 38988 1164
rect 38948 800 38976 1158
rect 39224 800 39252 1430
rect 39500 800 39528 2450
rect 39856 2440 39908 2446
rect 39856 2382 39908 2388
rect 39868 1834 39896 2382
rect 39856 1828 39908 1834
rect 39856 1770 39908 1776
rect 39764 1556 39816 1562
rect 39764 1498 39816 1504
rect 39776 800 39804 1498
rect 40052 800 40080 4150
rect 40328 4146 40356 4218
rect 40316 4140 40368 4146
rect 40316 4082 40368 4088
rect 40132 3460 40184 3466
rect 40132 3402 40184 3408
rect 40144 1154 40172 3402
rect 40420 2394 40448 4791
rect 40512 4146 40540 5086
rect 40592 5092 40644 5098
rect 40592 5034 40644 5040
rect 40500 4140 40552 4146
rect 40500 4082 40552 4088
rect 40328 2366 40448 2394
rect 40500 2440 40552 2446
rect 40500 2382 40552 2388
rect 40132 1148 40184 1154
rect 40132 1090 40184 1096
rect 40328 800 40356 2366
rect 40512 2106 40540 2382
rect 40500 2100 40552 2106
rect 40500 2042 40552 2048
rect 40604 800 40632 5034
rect 41052 5024 41104 5030
rect 41052 4966 41104 4972
rect 41064 4826 41092 4966
rect 41052 4820 41104 4826
rect 41052 4762 41104 4768
rect 41064 4622 41092 4762
rect 41340 4758 41368 4789
rect 41328 4752 41380 4758
rect 41326 4720 41328 4729
rect 41380 4720 41382 4729
rect 41236 4684 41288 4690
rect 41156 4644 41236 4672
rect 41052 4616 41104 4622
rect 41052 4558 41104 4564
rect 41156 4298 41184 4644
rect 41326 4655 41382 4664
rect 41236 4626 41288 4632
rect 41340 4622 41368 4655
rect 42812 4622 42840 5335
rect 43166 5128 43222 5137
rect 43166 5063 43222 5072
rect 42984 5024 43036 5030
rect 42984 4966 43036 4972
rect 42892 4684 42944 4690
rect 42892 4626 42944 4632
rect 41328 4616 41380 4622
rect 41328 4558 41380 4564
rect 42800 4616 42852 4622
rect 42800 4558 42852 4564
rect 41236 4480 41288 4486
rect 41236 4422 41288 4428
rect 42706 4448 42762 4457
rect 40972 4270 41184 4298
rect 41248 4282 41276 4422
rect 42706 4383 42762 4392
rect 41236 4276 41288 4282
rect 40972 4214 41000 4270
rect 41236 4218 41288 4224
rect 40960 4208 41012 4214
rect 40960 4150 41012 4156
rect 40684 4140 40736 4146
rect 40684 4082 40736 4088
rect 40868 4140 40920 4146
rect 40868 4082 40920 4088
rect 41328 4140 41380 4146
rect 41328 4082 41380 4088
rect 40696 3641 40724 4082
rect 40682 3632 40738 3641
rect 40880 3618 40908 4082
rect 41052 4004 41104 4010
rect 41052 3946 41104 3952
rect 40682 3567 40738 3576
rect 40788 3590 41000 3618
rect 40696 2553 40724 3567
rect 40788 3058 40816 3590
rect 40972 3534 41000 3590
rect 40868 3528 40920 3534
rect 40868 3470 40920 3476
rect 40960 3528 41012 3534
rect 40960 3470 41012 3476
rect 40880 3074 40908 3470
rect 41064 3398 41092 3946
rect 41340 3670 41368 4082
rect 41512 3936 41564 3942
rect 42432 3936 42484 3942
rect 41512 3878 41564 3884
rect 42430 3904 42432 3913
rect 42484 3904 42486 3913
rect 41328 3664 41380 3670
rect 41328 3606 41380 3612
rect 41524 3602 41552 3878
rect 42430 3839 42486 3848
rect 41972 3732 42024 3738
rect 41972 3674 42024 3680
rect 41512 3596 41564 3602
rect 41512 3538 41564 3544
rect 41788 3528 41840 3534
rect 41786 3496 41788 3505
rect 41840 3496 41842 3505
rect 41786 3431 41842 3440
rect 41052 3392 41104 3398
rect 41052 3334 41104 3340
rect 41064 3194 41092 3334
rect 41052 3188 41104 3194
rect 41052 3130 41104 3136
rect 41050 3088 41106 3097
rect 40776 3052 40828 3058
rect 40880 3046 41050 3074
rect 41050 3023 41052 3032
rect 40776 2994 40828 3000
rect 41104 3023 41106 3032
rect 41052 2994 41104 3000
rect 40788 2825 40816 2994
rect 41696 2848 41748 2854
rect 40774 2816 40830 2825
rect 41696 2790 41748 2796
rect 40774 2751 40830 2760
rect 40682 2544 40738 2553
rect 40682 2479 40738 2488
rect 40868 2100 40920 2106
rect 40868 2042 40920 2048
rect 40880 800 40908 2042
rect 41420 1964 41472 1970
rect 41420 1906 41472 1912
rect 41144 1420 41196 1426
rect 41144 1362 41196 1368
rect 41156 800 41184 1362
rect 41432 800 41460 1906
rect 41708 800 41736 2790
rect 41788 2304 41840 2310
rect 41786 2272 41788 2281
rect 41840 2272 41842 2281
rect 41786 2207 41842 2216
rect 41984 800 42012 3674
rect 42616 3528 42668 3534
rect 42616 3470 42668 3476
rect 42628 3369 42656 3470
rect 42720 3466 42748 4383
rect 42812 4146 42840 4558
rect 42800 4140 42852 4146
rect 42800 4082 42852 4088
rect 42904 4078 42932 4626
rect 42996 4622 43024 4966
rect 43180 4622 43208 5063
rect 42984 4616 43036 4622
rect 43168 4616 43220 4622
rect 42984 4558 43036 4564
rect 43088 4576 43168 4604
rect 43088 4468 43116 4576
rect 43168 4558 43220 4564
rect 42996 4440 43116 4468
rect 43168 4480 43220 4486
rect 42892 4072 42944 4078
rect 42892 4014 42944 4020
rect 42996 3516 43024 4440
rect 43168 4422 43220 4428
rect 43180 4146 43208 4422
rect 43548 4146 43576 11494
rect 43812 11076 43864 11082
rect 43812 11018 43864 11024
rect 43720 9920 43772 9926
rect 43720 9862 43772 9868
rect 43732 9382 43760 9862
rect 43720 9376 43772 9382
rect 43720 9318 43772 9324
rect 43628 8968 43680 8974
rect 43628 8910 43680 8916
rect 43640 8634 43668 8910
rect 43628 8628 43680 8634
rect 43628 8570 43680 8576
rect 43824 5352 43852 11018
rect 45008 11008 45060 11014
rect 45008 10950 45060 10956
rect 44294 10908 44602 10917
rect 44294 10906 44300 10908
rect 44356 10906 44380 10908
rect 44436 10906 44460 10908
rect 44516 10906 44540 10908
rect 44596 10906 44602 10908
rect 44356 10854 44358 10906
rect 44538 10854 44540 10906
rect 44294 10852 44300 10854
rect 44356 10852 44380 10854
rect 44436 10852 44460 10854
rect 44516 10852 44540 10854
rect 44596 10852 44602 10854
rect 44294 10843 44602 10852
rect 44088 10804 44140 10810
rect 44088 10746 44140 10752
rect 43996 10600 44048 10606
rect 43996 10542 44048 10548
rect 44008 10470 44036 10542
rect 43996 10464 44048 10470
rect 43996 10406 44048 10412
rect 44008 9382 44036 10406
rect 43996 9376 44048 9382
rect 43996 9318 44048 9324
rect 44008 7478 44036 9318
rect 43996 7472 44048 7478
rect 43996 7414 44048 7420
rect 43996 6792 44048 6798
rect 43996 6734 44048 6740
rect 44008 5914 44036 6734
rect 44100 6390 44128 10746
rect 45020 10538 45048 10950
rect 45008 10532 45060 10538
rect 45008 10474 45060 10480
rect 44180 9920 44232 9926
rect 44180 9862 44232 9868
rect 44640 9920 44692 9926
rect 44640 9862 44692 9868
rect 44192 9654 44220 9862
rect 44294 9820 44602 9829
rect 44294 9818 44300 9820
rect 44356 9818 44380 9820
rect 44436 9818 44460 9820
rect 44516 9818 44540 9820
rect 44596 9818 44602 9820
rect 44356 9766 44358 9818
rect 44538 9766 44540 9818
rect 44294 9764 44300 9766
rect 44356 9764 44380 9766
rect 44436 9764 44460 9766
rect 44516 9764 44540 9766
rect 44596 9764 44602 9766
rect 44294 9755 44602 9764
rect 44180 9648 44232 9654
rect 44180 9590 44232 9596
rect 44192 9058 44220 9590
rect 44652 9586 44680 9862
rect 45020 9586 45048 10474
rect 45468 10464 45520 10470
rect 45468 10406 45520 10412
rect 45480 9654 45508 10406
rect 45664 10062 45692 11698
rect 51518 11452 51826 11461
rect 51518 11450 51524 11452
rect 51580 11450 51604 11452
rect 51660 11450 51684 11452
rect 51740 11450 51764 11452
rect 51820 11450 51826 11452
rect 51580 11398 51582 11450
rect 51762 11398 51764 11450
rect 51518 11396 51524 11398
rect 51580 11396 51604 11398
rect 51660 11396 51684 11398
rect 51740 11396 51764 11398
rect 51820 11396 51826 11398
rect 51518 11387 51826 11396
rect 46940 10736 46992 10742
rect 46940 10678 46992 10684
rect 46756 10668 46808 10674
rect 46756 10610 46808 10616
rect 46388 10464 46440 10470
rect 46388 10406 46440 10412
rect 46400 10266 46428 10406
rect 46388 10260 46440 10266
rect 46388 10202 46440 10208
rect 46768 10062 46796 10610
rect 45652 10056 45704 10062
rect 45652 9998 45704 10004
rect 46480 10056 46532 10062
rect 46480 9998 46532 10004
rect 46756 10056 46808 10062
rect 46756 9998 46808 10004
rect 46492 9722 46520 9998
rect 46480 9716 46532 9722
rect 46480 9658 46532 9664
rect 45468 9648 45520 9654
rect 45468 9590 45520 9596
rect 44640 9580 44692 9586
rect 44640 9522 44692 9528
rect 45008 9580 45060 9586
rect 45008 9522 45060 9528
rect 44270 9072 44326 9081
rect 44192 9030 44270 9058
rect 44270 9007 44326 9016
rect 44284 8974 44312 9007
rect 44272 8968 44324 8974
rect 44652 8945 44680 9522
rect 44272 8910 44324 8916
rect 44638 8936 44694 8945
rect 44638 8871 44694 8880
rect 44294 8732 44602 8741
rect 44294 8730 44300 8732
rect 44356 8730 44380 8732
rect 44436 8730 44460 8732
rect 44516 8730 44540 8732
rect 44596 8730 44602 8732
rect 44356 8678 44358 8730
rect 44538 8678 44540 8730
rect 44294 8676 44300 8678
rect 44356 8676 44380 8678
rect 44436 8676 44460 8678
rect 44516 8676 44540 8678
rect 44596 8676 44602 8678
rect 44294 8667 44602 8676
rect 44640 8424 44692 8430
rect 44640 8366 44692 8372
rect 44180 8356 44232 8362
rect 44180 8298 44232 8304
rect 44192 7886 44220 8298
rect 44180 7880 44232 7886
rect 44180 7822 44232 7828
rect 44652 7750 44680 8366
rect 44640 7744 44692 7750
rect 44640 7686 44692 7692
rect 44294 7644 44602 7653
rect 44294 7642 44300 7644
rect 44356 7642 44380 7644
rect 44436 7642 44460 7644
rect 44516 7642 44540 7644
rect 44596 7642 44602 7644
rect 44356 7590 44358 7642
rect 44538 7590 44540 7642
rect 44294 7588 44300 7590
rect 44356 7588 44380 7590
rect 44436 7588 44460 7590
rect 44516 7588 44540 7590
rect 44596 7588 44602 7590
rect 44294 7579 44602 7588
rect 44652 7342 44680 7686
rect 45020 7342 45048 9522
rect 45480 8906 45508 9590
rect 46664 9580 46716 9586
rect 46664 9522 46716 9528
rect 46676 9178 46704 9522
rect 46768 9450 46796 9998
rect 46756 9444 46808 9450
rect 46756 9386 46808 9392
rect 46664 9172 46716 9178
rect 46664 9114 46716 9120
rect 46388 8968 46440 8974
rect 46388 8910 46440 8916
rect 46664 8968 46716 8974
rect 46664 8910 46716 8916
rect 45468 8900 45520 8906
rect 45468 8842 45520 8848
rect 45480 8498 45508 8842
rect 46296 8832 46348 8838
rect 46296 8774 46348 8780
rect 45284 8492 45336 8498
rect 45284 8434 45336 8440
rect 45468 8492 45520 8498
rect 45468 8434 45520 8440
rect 45100 8424 45152 8430
rect 45100 8366 45152 8372
rect 44640 7336 44692 7342
rect 44640 7278 44692 7284
rect 45008 7336 45060 7342
rect 45008 7278 45060 7284
rect 44180 7200 44232 7206
rect 44180 7142 44232 7148
rect 44088 6384 44140 6390
rect 44088 6326 44140 6332
rect 43996 5908 44048 5914
rect 43996 5850 44048 5856
rect 43732 5324 43852 5352
rect 43626 4720 43682 4729
rect 43626 4655 43682 4664
rect 43168 4140 43220 4146
rect 43168 4082 43220 4088
rect 43536 4140 43588 4146
rect 43536 4082 43588 4088
rect 43640 4078 43668 4655
rect 43628 4072 43680 4078
rect 43534 4040 43590 4049
rect 43628 4014 43680 4020
rect 43534 3975 43590 3984
rect 43168 3936 43220 3942
rect 43168 3878 43220 3884
rect 43076 3528 43128 3534
rect 42996 3488 43076 3516
rect 42708 3460 42760 3466
rect 42708 3402 42760 3408
rect 42614 3360 42670 3369
rect 42614 3295 42670 3304
rect 42628 3058 42656 3295
rect 42616 3052 42668 3058
rect 42616 2994 42668 3000
rect 42522 2000 42578 2009
rect 42522 1935 42578 1944
rect 42246 1864 42302 1873
rect 42246 1799 42302 1808
rect 42260 800 42288 1799
rect 42536 800 42564 1935
rect 42628 1737 42656 2994
rect 42720 2990 42748 3402
rect 42892 3392 42944 3398
rect 42892 3334 42944 3340
rect 42904 3126 42932 3334
rect 42892 3120 42944 3126
rect 42892 3062 42944 3068
rect 42708 2984 42760 2990
rect 42708 2926 42760 2932
rect 42798 2816 42854 2825
rect 42798 2751 42854 2760
rect 42708 2508 42760 2514
rect 42708 2450 42760 2456
rect 42720 2106 42748 2450
rect 42708 2100 42760 2106
rect 42708 2042 42760 2048
rect 42614 1728 42670 1737
rect 42614 1663 42670 1672
rect 42812 800 42840 2751
rect 42996 1329 43024 3488
rect 43076 3470 43128 3476
rect 43076 2440 43128 2446
rect 43076 2382 43128 2388
rect 43088 2038 43116 2382
rect 43076 2032 43128 2038
rect 43076 1974 43128 1980
rect 43180 1850 43208 3878
rect 43548 3040 43576 3975
rect 43732 3534 43760 5324
rect 44100 5302 44128 6326
rect 44192 5710 44220 7142
rect 45008 6860 45060 6866
rect 45008 6802 45060 6808
rect 44294 6556 44602 6565
rect 44294 6554 44300 6556
rect 44356 6554 44380 6556
rect 44436 6554 44460 6556
rect 44516 6554 44540 6556
rect 44596 6554 44602 6556
rect 44356 6502 44358 6554
rect 44538 6502 44540 6554
rect 44294 6500 44300 6502
rect 44356 6500 44380 6502
rect 44436 6500 44460 6502
rect 44516 6500 44540 6502
rect 44596 6500 44602 6502
rect 44294 6491 44602 6500
rect 45020 5710 45048 6802
rect 45112 6322 45140 8366
rect 45296 7954 45324 8434
rect 46308 8090 46336 8774
rect 46400 8090 46428 8910
rect 46676 8634 46704 8910
rect 46664 8628 46716 8634
rect 46952 8616 46980 10678
rect 50528 10600 50580 10606
rect 50528 10542 50580 10548
rect 48964 10464 49016 10470
rect 48964 10406 49016 10412
rect 47216 10260 47268 10266
rect 47216 10202 47268 10208
rect 46664 8570 46716 8576
rect 46768 8588 46980 8616
rect 46768 8498 46796 8588
rect 46756 8492 46808 8498
rect 46756 8434 46808 8440
rect 46848 8492 46900 8498
rect 46848 8434 46900 8440
rect 46860 8362 46888 8434
rect 46952 8430 46980 8588
rect 46940 8424 46992 8430
rect 46940 8366 46992 8372
rect 46848 8356 46900 8362
rect 46848 8298 46900 8304
rect 46940 8288 46992 8294
rect 46940 8230 46992 8236
rect 46296 8084 46348 8090
rect 46296 8026 46348 8032
rect 46388 8084 46440 8090
rect 46388 8026 46440 8032
rect 45284 7948 45336 7954
rect 45284 7890 45336 7896
rect 46952 7886 46980 8230
rect 46020 7880 46072 7886
rect 46020 7822 46072 7828
rect 46940 7880 46992 7886
rect 46940 7822 46992 7828
rect 45376 7812 45428 7818
rect 45376 7754 45428 7760
rect 45388 7410 45416 7754
rect 46032 7546 46060 7822
rect 46020 7540 46072 7546
rect 46020 7482 46072 7488
rect 45376 7404 45428 7410
rect 45376 7346 45428 7352
rect 46848 7200 46900 7206
rect 46848 7142 46900 7148
rect 46860 6798 46888 7142
rect 47228 6905 47256 10202
rect 48976 10130 49004 10406
rect 48964 10124 49016 10130
rect 48964 10066 49016 10072
rect 47676 10056 47728 10062
rect 47676 9998 47728 10004
rect 47688 9722 47716 9998
rect 48872 9920 48924 9926
rect 48872 9862 48924 9868
rect 47676 9716 47728 9722
rect 47676 9658 47728 9664
rect 48136 9580 48188 9586
rect 48136 9522 48188 9528
rect 48148 9178 48176 9522
rect 48136 9172 48188 9178
rect 48136 9114 48188 9120
rect 48228 9172 48280 9178
rect 48228 9114 48280 9120
rect 48240 8974 48268 9114
rect 48884 8974 48912 9862
rect 48976 9518 49004 10066
rect 49240 10056 49292 10062
rect 49240 9998 49292 10004
rect 48964 9512 49016 9518
rect 48964 9454 49016 9460
rect 48228 8968 48280 8974
rect 48228 8910 48280 8916
rect 48872 8968 48924 8974
rect 48872 8910 48924 8916
rect 48240 8566 48268 8910
rect 48412 8900 48464 8906
rect 48412 8842 48464 8848
rect 48424 8566 48452 8842
rect 49252 8634 49280 9998
rect 50068 9988 50120 9994
rect 50068 9930 50120 9936
rect 50080 9586 50108 9930
rect 50540 9654 50568 10542
rect 51518 10364 51826 10373
rect 51518 10362 51524 10364
rect 51580 10362 51604 10364
rect 51660 10362 51684 10364
rect 51740 10362 51764 10364
rect 51820 10362 51826 10364
rect 51580 10310 51582 10362
rect 51762 10310 51764 10362
rect 51518 10308 51524 10310
rect 51580 10308 51604 10310
rect 51660 10308 51684 10310
rect 51740 10308 51764 10310
rect 51820 10308 51826 10310
rect 51518 10299 51826 10308
rect 52276 10124 52328 10130
rect 52276 10066 52328 10072
rect 50528 9648 50580 9654
rect 50528 9590 50580 9596
rect 50068 9580 50120 9586
rect 50068 9522 50120 9528
rect 50540 9518 50568 9590
rect 51264 9580 51316 9586
rect 51264 9522 51316 9528
rect 52000 9580 52052 9586
rect 52000 9522 52052 9528
rect 49700 9512 49752 9518
rect 49700 9454 49752 9460
rect 50528 9512 50580 9518
rect 50528 9454 50580 9460
rect 49240 8628 49292 8634
rect 49240 8570 49292 8576
rect 48228 8560 48280 8566
rect 48228 8502 48280 8508
rect 48412 8560 48464 8566
rect 48412 8502 48464 8508
rect 49148 8560 49200 8566
rect 49200 8508 49280 8514
rect 49148 8502 49280 8508
rect 49160 8486 49280 8502
rect 48320 8356 48372 8362
rect 48320 8298 48372 8304
rect 47584 8288 47636 8294
rect 47584 8230 47636 8236
rect 48042 8256 48098 8265
rect 47596 7750 47624 8230
rect 48042 8191 48098 8200
rect 47584 7744 47636 7750
rect 47584 7686 47636 7692
rect 48056 7342 48084 8191
rect 48332 7954 48360 8298
rect 49148 8288 49200 8294
rect 49148 8230 49200 8236
rect 48320 7948 48372 7954
rect 48320 7890 48372 7896
rect 49160 7886 49188 8230
rect 49148 7880 49200 7886
rect 49148 7822 49200 7828
rect 49252 7342 49280 8486
rect 49332 8492 49384 8498
rect 49332 8434 49384 8440
rect 49344 8022 49372 8434
rect 49712 8362 49740 9454
rect 50528 9376 50580 9382
rect 50528 9318 50580 9324
rect 50540 9110 50568 9318
rect 51276 9178 51304 9522
rect 51448 9512 51500 9518
rect 51448 9454 51500 9460
rect 51264 9172 51316 9178
rect 51264 9114 51316 9120
rect 50528 9104 50580 9110
rect 50528 9046 50580 9052
rect 50344 8900 50396 8906
rect 50344 8842 50396 8848
rect 50712 8900 50764 8906
rect 50712 8842 50764 8848
rect 50068 8492 50120 8498
rect 50068 8434 50120 8440
rect 49700 8356 49752 8362
rect 49700 8298 49752 8304
rect 49884 8356 49936 8362
rect 49884 8298 49936 8304
rect 49896 8265 49924 8298
rect 49882 8256 49938 8265
rect 49882 8191 49938 8200
rect 49332 8016 49384 8022
rect 49332 7958 49384 7964
rect 49344 7886 49372 7958
rect 50080 7954 50108 8434
rect 50068 7948 50120 7954
rect 50068 7890 50120 7896
rect 50356 7886 50384 8842
rect 50724 8430 50752 8842
rect 51172 8832 51224 8838
rect 51172 8774 51224 8780
rect 50804 8492 50856 8498
rect 50804 8434 50856 8440
rect 50712 8424 50764 8430
rect 50712 8366 50764 8372
rect 50620 8288 50672 8294
rect 50620 8230 50672 8236
rect 49332 7880 49384 7886
rect 49332 7822 49384 7828
rect 50344 7880 50396 7886
rect 50344 7822 50396 7828
rect 50356 7410 50384 7822
rect 50632 7410 50660 8230
rect 50816 8090 50844 8434
rect 51184 8090 51212 8774
rect 51356 8356 51408 8362
rect 51356 8298 51408 8304
rect 51368 8090 51396 8298
rect 50804 8084 50856 8090
rect 50804 8026 50856 8032
rect 51172 8084 51224 8090
rect 51172 8026 51224 8032
rect 51356 8084 51408 8090
rect 51356 8026 51408 8032
rect 51184 7546 51212 8026
rect 51460 7546 51488 9454
rect 51518 9276 51826 9285
rect 51518 9274 51524 9276
rect 51580 9274 51604 9276
rect 51660 9274 51684 9276
rect 51740 9274 51764 9276
rect 51820 9274 51826 9276
rect 51580 9222 51582 9274
rect 51762 9222 51764 9274
rect 51518 9220 51524 9222
rect 51580 9220 51604 9222
rect 51660 9220 51684 9222
rect 51740 9220 51764 9222
rect 51820 9220 51826 9222
rect 51518 9211 51826 9220
rect 51540 8968 51592 8974
rect 51540 8910 51592 8916
rect 51552 8498 51580 8910
rect 52012 8634 52040 9522
rect 52288 9518 52316 10066
rect 52552 10056 52604 10062
rect 52552 9998 52604 10004
rect 53380 10056 53432 10062
rect 53380 9998 53432 10004
rect 52276 9512 52328 9518
rect 52276 9454 52328 9460
rect 52288 9042 52316 9454
rect 52564 9382 52592 9998
rect 53392 9654 53420 9998
rect 53380 9648 53432 9654
rect 53380 9590 53432 9596
rect 52552 9376 52604 9382
rect 52552 9318 52604 9324
rect 52276 9036 52328 9042
rect 52276 8978 52328 8984
rect 53392 8974 53420 9590
rect 52092 8968 52144 8974
rect 52092 8910 52144 8916
rect 53380 8968 53432 8974
rect 53380 8910 53432 8916
rect 54116 8968 54168 8974
rect 54116 8910 54168 8916
rect 52000 8628 52052 8634
rect 52000 8570 52052 8576
rect 51540 8492 51592 8498
rect 51540 8434 51592 8440
rect 51518 8188 51826 8197
rect 51518 8186 51524 8188
rect 51580 8186 51604 8188
rect 51660 8186 51684 8188
rect 51740 8186 51764 8188
rect 51820 8186 51826 8188
rect 51580 8134 51582 8186
rect 51762 8134 51764 8186
rect 51518 8132 51524 8134
rect 51580 8132 51604 8134
rect 51660 8132 51684 8134
rect 51740 8132 51764 8134
rect 51820 8132 51826 8134
rect 51518 8123 51826 8132
rect 51172 7540 51224 7546
rect 51172 7482 51224 7488
rect 51448 7540 51500 7546
rect 51448 7482 51500 7488
rect 52104 7410 52132 8910
rect 54128 8634 54156 8910
rect 54116 8628 54168 8634
rect 54116 8570 54168 8576
rect 55772 8492 55824 8498
rect 55772 8434 55824 8440
rect 54392 8424 54444 8430
rect 54392 8366 54444 8372
rect 52920 8356 52972 8362
rect 52920 8298 52972 8304
rect 53196 8356 53248 8362
rect 53196 8298 53248 8304
rect 52460 7812 52512 7818
rect 52460 7754 52512 7760
rect 52184 7744 52236 7750
rect 52184 7686 52236 7692
rect 50344 7404 50396 7410
rect 50344 7346 50396 7352
rect 50620 7404 50672 7410
rect 50620 7346 50672 7352
rect 52092 7404 52144 7410
rect 52092 7346 52144 7352
rect 48044 7336 48096 7342
rect 48044 7278 48096 7284
rect 49240 7336 49292 7342
rect 49240 7278 49292 7284
rect 48594 7032 48650 7041
rect 49252 7002 49280 7278
rect 50068 7268 50120 7274
rect 50068 7210 50120 7216
rect 48594 6967 48596 6976
rect 48648 6967 48650 6976
rect 49240 6996 49292 7002
rect 48596 6938 48648 6944
rect 49240 6938 49292 6944
rect 47214 6896 47270 6905
rect 47214 6831 47270 6840
rect 46572 6792 46624 6798
rect 46572 6734 46624 6740
rect 46848 6792 46900 6798
rect 46848 6734 46900 6740
rect 46204 6452 46256 6458
rect 46204 6394 46256 6400
rect 45100 6316 45152 6322
rect 45100 6258 45152 6264
rect 45376 6316 45428 6322
rect 45376 6258 45428 6264
rect 45388 5778 45416 6258
rect 45834 6216 45890 6225
rect 45834 6151 45836 6160
rect 45888 6151 45890 6160
rect 45836 6122 45888 6128
rect 45652 5908 45704 5914
rect 45652 5850 45704 5856
rect 45560 5840 45612 5846
rect 45664 5817 45692 5850
rect 45560 5782 45612 5788
rect 45650 5808 45706 5817
rect 45376 5772 45428 5778
rect 45376 5714 45428 5720
rect 44180 5704 44232 5710
rect 44180 5646 44232 5652
rect 45008 5704 45060 5710
rect 45008 5646 45060 5652
rect 45284 5704 45336 5710
rect 45284 5646 45336 5652
rect 44294 5468 44602 5477
rect 44294 5466 44300 5468
rect 44356 5466 44380 5468
rect 44436 5466 44460 5468
rect 44516 5466 44540 5468
rect 44596 5466 44602 5468
rect 44356 5414 44358 5466
rect 44538 5414 44540 5466
rect 44294 5412 44300 5414
rect 44356 5412 44380 5414
rect 44436 5412 44460 5414
rect 44516 5412 44540 5414
rect 44596 5412 44602 5414
rect 44294 5403 44602 5412
rect 44088 5296 44140 5302
rect 44088 5238 44140 5244
rect 44456 5296 44508 5302
rect 44456 5238 44508 5244
rect 43812 5228 43864 5234
rect 43812 5170 43864 5176
rect 43824 4826 43852 5170
rect 43812 4820 43864 4826
rect 43812 4762 43864 4768
rect 44468 4758 44496 5238
rect 45192 5228 45244 5234
rect 45192 5170 45244 5176
rect 45204 4826 45232 5170
rect 45192 4820 45244 4826
rect 45192 4762 45244 4768
rect 44456 4752 44508 4758
rect 44456 4694 44508 4700
rect 44468 4622 44496 4694
rect 44456 4616 44508 4622
rect 44456 4558 44508 4564
rect 44088 4480 44140 4486
rect 44008 4440 44088 4468
rect 44008 4282 44036 4440
rect 44088 4422 44140 4428
rect 44822 4448 44878 4457
rect 44294 4380 44602 4389
rect 44822 4383 44878 4392
rect 44294 4378 44300 4380
rect 44356 4378 44380 4380
rect 44436 4378 44460 4380
rect 44516 4378 44540 4380
rect 44596 4378 44602 4380
rect 44356 4326 44358 4378
rect 44538 4326 44540 4378
rect 44294 4324 44300 4326
rect 44356 4324 44380 4326
rect 44436 4324 44460 4326
rect 44516 4324 44540 4326
rect 44596 4324 44602 4326
rect 44086 4312 44142 4321
rect 44294 4315 44602 4324
rect 43996 4276 44048 4282
rect 44086 4247 44142 4256
rect 43996 4218 44048 4224
rect 44100 4196 44128 4247
rect 44100 4168 44220 4196
rect 43996 4140 44048 4146
rect 44048 4100 44128 4128
rect 43996 4082 44048 4088
rect 44100 3534 44128 4100
rect 43720 3528 43772 3534
rect 43720 3470 43772 3476
rect 43904 3528 43956 3534
rect 43904 3470 43956 3476
rect 44088 3528 44140 3534
rect 44088 3470 44140 3476
rect 43732 3369 43760 3470
rect 43718 3360 43774 3369
rect 43718 3295 43774 3304
rect 43628 3052 43680 3058
rect 43548 3012 43628 3040
rect 43628 2994 43680 3000
rect 43260 2916 43312 2922
rect 43260 2858 43312 2864
rect 43088 1822 43208 1850
rect 42982 1320 43038 1329
rect 42982 1255 43038 1264
rect 43088 800 43116 1822
rect 43272 1578 43300 2858
rect 43732 2650 43760 3295
rect 43916 3194 43944 3470
rect 44100 3233 44128 3470
rect 44086 3224 44142 3233
rect 43904 3188 43956 3194
rect 43904 3130 43956 3136
rect 43996 3188 44048 3194
rect 44086 3159 44142 3168
rect 43996 3130 44048 3136
rect 43812 3120 43864 3126
rect 43810 3088 43812 3097
rect 43864 3088 43866 3097
rect 43810 3023 43866 3032
rect 43720 2644 43772 2650
rect 43720 2586 43772 2592
rect 43902 2544 43958 2553
rect 43902 2479 43958 2488
rect 43916 2446 43944 2479
rect 43720 2440 43772 2446
rect 43720 2382 43772 2388
rect 43904 2440 43956 2446
rect 43904 2382 43956 2388
rect 43628 1828 43680 1834
rect 43628 1770 43680 1776
rect 43272 1550 43392 1578
rect 43364 800 43392 1550
rect 43640 800 43668 1770
rect 43732 1222 43760 2382
rect 44008 2122 44036 3130
rect 44100 2553 44128 3159
rect 44192 3058 44220 4168
rect 44456 4140 44508 4146
rect 44456 4082 44508 4088
rect 44468 4049 44496 4082
rect 44454 4040 44510 4049
rect 44454 3975 44510 3984
rect 44640 3528 44692 3534
rect 44640 3470 44692 3476
rect 44294 3292 44602 3301
rect 44294 3290 44300 3292
rect 44356 3290 44380 3292
rect 44436 3290 44460 3292
rect 44516 3290 44540 3292
rect 44596 3290 44602 3292
rect 44356 3238 44358 3290
rect 44538 3238 44540 3290
rect 44294 3236 44300 3238
rect 44356 3236 44380 3238
rect 44436 3236 44460 3238
rect 44516 3236 44540 3238
rect 44596 3236 44602 3238
rect 44294 3227 44602 3236
rect 44180 3052 44232 3058
rect 44180 2994 44232 3000
rect 44652 2972 44680 3470
rect 44560 2944 44680 2972
rect 44560 2854 44588 2944
rect 44548 2848 44600 2854
rect 44548 2790 44600 2796
rect 44086 2544 44142 2553
rect 44086 2479 44142 2488
rect 44294 2204 44602 2213
rect 44294 2202 44300 2204
rect 44356 2202 44380 2204
rect 44436 2202 44460 2204
rect 44516 2202 44540 2204
rect 44596 2202 44602 2204
rect 44356 2150 44358 2202
rect 44538 2150 44540 2202
rect 44294 2148 44300 2150
rect 44356 2148 44380 2150
rect 44436 2148 44460 2150
rect 44516 2148 44540 2150
rect 44596 2148 44602 2150
rect 44294 2139 44602 2148
rect 43916 2094 44036 2122
rect 44732 2100 44784 2106
rect 43720 1216 43772 1222
rect 43720 1158 43772 1164
rect 43916 800 43944 2094
rect 44732 2042 44784 2048
rect 44456 2032 44508 2038
rect 44456 1974 44508 1980
rect 44180 1692 44232 1698
rect 44180 1634 44232 1640
rect 44192 800 44220 1634
rect 44468 800 44496 1974
rect 44744 800 44772 2042
rect 44836 1698 44864 4383
rect 45296 4026 45324 5646
rect 45466 5264 45522 5273
rect 45466 5199 45522 5208
rect 45376 4684 45428 4690
rect 45376 4626 45428 4632
rect 45388 4214 45416 4626
rect 45480 4554 45508 5199
rect 45468 4548 45520 4554
rect 45468 4490 45520 4496
rect 45376 4208 45428 4214
rect 45376 4150 45428 4156
rect 45008 4004 45060 4010
rect 45008 3946 45060 3952
rect 45204 3998 45324 4026
rect 44916 3936 44968 3942
rect 44916 3878 44968 3884
rect 44928 3738 44956 3878
rect 44916 3732 44968 3738
rect 44916 3674 44968 3680
rect 45020 3194 45048 3946
rect 45100 3392 45152 3398
rect 45100 3334 45152 3340
rect 45008 3188 45060 3194
rect 45008 3130 45060 3136
rect 45112 3126 45140 3334
rect 45100 3120 45152 3126
rect 45100 3062 45152 3068
rect 45008 3052 45060 3058
rect 45008 2994 45060 3000
rect 44916 2848 44968 2854
rect 44916 2790 44968 2796
rect 44824 1692 44876 1698
rect 44824 1634 44876 1640
rect 44928 1494 44956 2790
rect 44916 1488 44968 1494
rect 44916 1430 44968 1436
rect 45020 800 45048 2994
rect 45100 2372 45152 2378
rect 45100 2314 45152 2320
rect 45112 1902 45140 2314
rect 45204 2106 45232 3998
rect 45284 3936 45336 3942
rect 45284 3878 45336 3884
rect 45296 2922 45324 3878
rect 45284 2916 45336 2922
rect 45284 2858 45336 2864
rect 45192 2100 45244 2106
rect 45192 2042 45244 2048
rect 45284 2100 45336 2106
rect 45284 2042 45336 2048
rect 45100 1896 45152 1902
rect 45100 1838 45152 1844
rect 45296 800 45324 2042
rect 45572 800 45600 5782
rect 45650 5743 45706 5752
rect 45928 5228 45980 5234
rect 45928 5170 45980 5176
rect 45940 4622 45968 5170
rect 46216 5166 46244 6394
rect 46584 5574 46612 6734
rect 46848 6316 46900 6322
rect 46848 6258 46900 6264
rect 46860 5642 46888 6258
rect 47228 5710 47256 6831
rect 48608 6730 48636 6938
rect 49332 6792 49384 6798
rect 49332 6734 49384 6740
rect 48596 6724 48648 6730
rect 48596 6666 48648 6672
rect 48044 6656 48096 6662
rect 48044 6598 48096 6604
rect 48056 6118 48084 6598
rect 49344 6118 49372 6734
rect 49976 6452 50028 6458
rect 49976 6394 50028 6400
rect 49424 6248 49476 6254
rect 49424 6190 49476 6196
rect 48044 6112 48096 6118
rect 48044 6054 48096 6060
rect 49332 6112 49384 6118
rect 49332 6054 49384 6060
rect 49240 5840 49292 5846
rect 49240 5782 49292 5788
rect 47584 5772 47636 5778
rect 47584 5714 47636 5720
rect 47216 5704 47268 5710
rect 47216 5646 47268 5652
rect 46848 5636 46900 5642
rect 46848 5578 46900 5584
rect 46572 5568 46624 5574
rect 46572 5510 46624 5516
rect 46860 5370 46888 5578
rect 46848 5364 46900 5370
rect 46848 5306 46900 5312
rect 47228 5234 47256 5646
rect 47596 5370 47624 5714
rect 49252 5710 49280 5782
rect 49240 5704 49292 5710
rect 49240 5646 49292 5652
rect 48320 5568 48372 5574
rect 48320 5510 48372 5516
rect 47584 5364 47636 5370
rect 47584 5306 47636 5312
rect 48332 5302 48360 5510
rect 49436 5370 49464 6190
rect 49988 6118 50016 6394
rect 50080 6322 50108 7210
rect 50712 7200 50764 7206
rect 50712 7142 50764 7148
rect 51264 7200 51316 7206
rect 51264 7142 51316 7148
rect 50528 6792 50580 6798
rect 50528 6734 50580 6740
rect 50540 6458 50568 6734
rect 50528 6452 50580 6458
rect 50528 6394 50580 6400
rect 50724 6322 50752 7142
rect 51276 7041 51304 7142
rect 51518 7100 51826 7109
rect 51518 7098 51524 7100
rect 51580 7098 51604 7100
rect 51660 7098 51684 7100
rect 51740 7098 51764 7100
rect 51820 7098 51826 7100
rect 51580 7046 51582 7098
rect 51762 7046 51764 7098
rect 51518 7044 51524 7046
rect 51580 7044 51604 7046
rect 51660 7044 51684 7046
rect 51740 7044 51764 7046
rect 51820 7044 51826 7046
rect 51262 7032 51318 7041
rect 51518 7035 51826 7044
rect 51262 6967 51264 6976
rect 51316 6967 51318 6976
rect 51264 6938 51316 6944
rect 51276 6907 51304 6938
rect 52196 6905 52224 7686
rect 52368 7336 52420 7342
rect 52368 7278 52420 7284
rect 52380 7002 52408 7278
rect 52368 6996 52420 7002
rect 52368 6938 52420 6944
rect 52276 6928 52328 6934
rect 52182 6896 52238 6905
rect 52276 6870 52328 6876
rect 52182 6831 52238 6840
rect 52184 6724 52236 6730
rect 52184 6666 52236 6672
rect 51448 6656 51500 6662
rect 51448 6598 51500 6604
rect 51460 6390 51488 6598
rect 51448 6384 51500 6390
rect 51448 6326 51500 6332
rect 50068 6316 50120 6322
rect 50068 6258 50120 6264
rect 50712 6316 50764 6322
rect 50712 6258 50764 6264
rect 52196 6254 52224 6666
rect 52184 6248 52236 6254
rect 52184 6190 52236 6196
rect 49976 6112 50028 6118
rect 49976 6054 50028 6060
rect 51518 6012 51826 6021
rect 51518 6010 51524 6012
rect 51580 6010 51604 6012
rect 51660 6010 51684 6012
rect 51740 6010 51764 6012
rect 51820 6010 51826 6012
rect 51580 5958 51582 6010
rect 51762 5958 51764 6010
rect 51518 5956 51524 5958
rect 51580 5956 51604 5958
rect 51660 5956 51684 5958
rect 51740 5956 51764 5958
rect 51820 5956 51826 5958
rect 50802 5944 50858 5953
rect 51518 5947 51826 5956
rect 50802 5879 50858 5888
rect 50816 5846 50844 5879
rect 50804 5840 50856 5846
rect 50804 5782 50856 5788
rect 52184 5704 52236 5710
rect 52184 5646 52236 5652
rect 48688 5364 48740 5370
rect 48688 5306 48740 5312
rect 49424 5364 49476 5370
rect 49424 5306 49476 5312
rect 49516 5364 49568 5370
rect 49516 5306 49568 5312
rect 51448 5364 51500 5370
rect 51448 5306 51500 5312
rect 48320 5296 48372 5302
rect 48320 5238 48372 5244
rect 47216 5228 47268 5234
rect 47216 5170 47268 5176
rect 46020 5160 46072 5166
rect 46020 5102 46072 5108
rect 46204 5160 46256 5166
rect 46204 5102 46256 5108
rect 45928 4616 45980 4622
rect 45928 4558 45980 4564
rect 46032 4486 46060 5102
rect 48136 5024 48188 5030
rect 48136 4966 48188 4972
rect 46202 4856 46258 4865
rect 46202 4791 46258 4800
rect 46940 4820 46992 4826
rect 46020 4480 46072 4486
rect 46020 4422 46072 4428
rect 46032 4282 46060 4422
rect 46020 4276 46072 4282
rect 46020 4218 46072 4224
rect 45650 3496 45706 3505
rect 45650 3431 45706 3440
rect 45664 3398 45692 3431
rect 45652 3392 45704 3398
rect 45652 3334 45704 3340
rect 45836 3188 45888 3194
rect 45836 3130 45888 3136
rect 45742 2952 45798 2961
rect 45742 2887 45744 2896
rect 45796 2887 45798 2896
rect 45744 2858 45796 2864
rect 45652 2848 45704 2854
rect 45652 2790 45704 2796
rect 45664 1562 45692 2790
rect 45652 1556 45704 1562
rect 45652 1498 45704 1504
rect 45848 800 45876 3130
rect 46216 2854 46244 4791
rect 46940 4762 46992 4768
rect 46754 4040 46810 4049
rect 46754 3975 46810 3984
rect 46570 3904 46626 3913
rect 46570 3839 46626 3848
rect 46584 3602 46612 3839
rect 46572 3596 46624 3602
rect 46572 3538 46624 3544
rect 46480 3460 46532 3466
rect 46480 3402 46532 3408
rect 46204 2848 46256 2854
rect 46204 2790 46256 2796
rect 46492 2774 46520 3402
rect 46400 2746 46520 2774
rect 46112 1896 46164 1902
rect 46112 1838 46164 1844
rect 46124 800 46152 1838
rect 46400 800 46428 2746
rect 46584 2650 46612 3538
rect 46572 2644 46624 2650
rect 46572 2586 46624 2592
rect 46768 2310 46796 3975
rect 46848 2848 46900 2854
rect 46848 2790 46900 2796
rect 46756 2304 46808 2310
rect 46756 2246 46808 2252
rect 46664 1692 46716 1698
rect 46664 1634 46716 1640
rect 46676 800 46704 1634
rect 46860 1426 46888 2790
rect 46848 1420 46900 1426
rect 46848 1362 46900 1368
rect 46952 800 46980 4762
rect 48148 4486 48176 4966
rect 48410 4720 48466 4729
rect 48700 4690 48728 5306
rect 49528 5166 49556 5306
rect 49516 5160 49568 5166
rect 49516 5102 49568 5108
rect 51078 5128 51134 5137
rect 51078 5063 51134 5072
rect 51092 5030 51120 5063
rect 50252 5024 50304 5030
rect 50252 4966 50304 4972
rect 51080 5024 51132 5030
rect 51080 4966 51132 4972
rect 48410 4655 48466 4664
rect 48688 4684 48740 4690
rect 48424 4622 48452 4655
rect 48688 4626 48740 4632
rect 48412 4616 48464 4622
rect 48412 4558 48464 4564
rect 48320 4548 48372 4554
rect 48320 4490 48372 4496
rect 48504 4548 48556 4554
rect 48504 4490 48556 4496
rect 48596 4548 48648 4554
rect 48596 4490 48648 4496
rect 48136 4480 48188 4486
rect 48136 4422 48188 4428
rect 48332 4282 48360 4490
rect 48516 4457 48544 4490
rect 48502 4448 48558 4457
rect 48502 4383 48558 4392
rect 48320 4276 48372 4282
rect 48320 4218 48372 4224
rect 47768 3936 47820 3942
rect 47768 3878 47820 3884
rect 47582 3768 47638 3777
rect 47582 3703 47638 3712
rect 47216 3460 47268 3466
rect 47216 3402 47268 3408
rect 47228 800 47256 3402
rect 47596 2990 47624 3703
rect 47584 2984 47636 2990
rect 47584 2926 47636 2932
rect 47780 1986 47808 3878
rect 48044 3732 48096 3738
rect 48044 3674 48096 3680
rect 47858 2680 47914 2689
rect 47858 2615 47914 2624
rect 47504 1958 47808 1986
rect 47504 800 47532 1958
rect 47872 1442 47900 2615
rect 47780 1414 47900 1442
rect 47780 800 47808 1414
rect 48056 800 48084 3674
rect 48320 3460 48372 3466
rect 48320 3402 48372 3408
rect 48332 3097 48360 3402
rect 48318 3088 48374 3097
rect 48318 3023 48374 3032
rect 48502 3088 48558 3097
rect 48502 3023 48558 3032
rect 48516 2774 48544 3023
rect 48424 2746 48544 2774
rect 48228 2440 48280 2446
rect 48228 2382 48280 2388
rect 48240 1970 48268 2382
rect 48228 1964 48280 1970
rect 48228 1906 48280 1912
rect 48424 1442 48452 2746
rect 48332 1414 48452 1442
rect 48332 800 48360 1414
rect 48608 800 48636 4490
rect 49608 4140 49660 4146
rect 49608 4082 49660 4088
rect 49620 3602 49648 4082
rect 49700 4004 49752 4010
rect 49700 3946 49752 3952
rect 49608 3596 49660 3602
rect 49608 3538 49660 3544
rect 49424 3120 49476 3126
rect 49424 3062 49476 3068
rect 49436 2938 49464 3062
rect 49620 3058 49648 3538
rect 49608 3052 49660 3058
rect 49608 2994 49660 3000
rect 49344 2910 49464 2938
rect 49344 2854 49372 2910
rect 48780 2848 48832 2854
rect 48780 2790 48832 2796
rect 49332 2848 49384 2854
rect 49332 2790 49384 2796
rect 48792 1442 48820 2790
rect 49620 2774 49648 2994
rect 49528 2746 49648 2774
rect 49528 2650 49556 2746
rect 49516 2644 49568 2650
rect 49516 2586 49568 2592
rect 48872 2440 48924 2446
rect 49516 2440 49568 2446
rect 48872 2382 48924 2388
rect 49514 2408 49516 2417
rect 49568 2408 49570 2417
rect 48884 1873 48912 2382
rect 49424 2372 49476 2378
rect 49514 2343 49570 2352
rect 49424 2314 49476 2320
rect 49056 2304 49108 2310
rect 49056 2246 49108 2252
rect 49148 2304 49200 2310
rect 49148 2246 49200 2252
rect 48870 1864 48926 1873
rect 48870 1799 48926 1808
rect 49068 1766 49096 2246
rect 49056 1760 49108 1766
rect 49056 1702 49108 1708
rect 48792 1414 48912 1442
rect 48884 800 48912 1414
rect 49160 800 49188 2246
rect 49436 800 49464 2314
rect 49712 800 49740 3946
rect 50160 2916 50212 2922
rect 50160 2858 50212 2864
rect 49976 2848 50028 2854
rect 49974 2816 49976 2825
rect 50028 2816 50030 2825
rect 49974 2751 50030 2760
rect 50172 2689 50200 2858
rect 50158 2680 50214 2689
rect 50158 2615 50214 2624
rect 50160 2440 50212 2446
rect 50160 2382 50212 2388
rect 50172 2009 50200 2382
rect 50158 2000 50214 2009
rect 50158 1935 50214 1944
rect 49976 1488 50028 1494
rect 49976 1430 50028 1436
rect 49988 800 50016 1430
rect 50264 800 50292 4966
rect 51460 4826 51488 5306
rect 52092 5228 52144 5234
rect 52092 5170 52144 5176
rect 52104 5098 52132 5170
rect 52092 5092 52144 5098
rect 52092 5034 52144 5040
rect 51908 5024 51960 5030
rect 51908 4966 51960 4972
rect 52000 5024 52052 5030
rect 52000 4966 52052 4972
rect 51518 4924 51826 4933
rect 51518 4922 51524 4924
rect 51580 4922 51604 4924
rect 51660 4922 51684 4924
rect 51740 4922 51764 4924
rect 51820 4922 51826 4924
rect 51580 4870 51582 4922
rect 51762 4870 51764 4922
rect 51518 4868 51524 4870
rect 51580 4868 51604 4870
rect 51660 4868 51684 4870
rect 51740 4868 51764 4870
rect 51820 4868 51826 4870
rect 51518 4859 51826 4868
rect 51920 4826 51948 4966
rect 51448 4820 51500 4826
rect 51448 4762 51500 4768
rect 51908 4820 51960 4826
rect 51908 4762 51960 4768
rect 52012 4282 52040 4966
rect 52000 4276 52052 4282
rect 52000 4218 52052 4224
rect 52104 4185 52132 5034
rect 52090 4176 52146 4185
rect 51264 4140 51316 4146
rect 51264 4082 51316 4088
rect 51816 4140 51868 4146
rect 52196 4146 52224 5646
rect 52090 4111 52146 4120
rect 52184 4140 52236 4146
rect 51816 4082 51868 4088
rect 52184 4082 52236 4088
rect 51080 3936 51132 3942
rect 51080 3878 51132 3884
rect 50526 2952 50582 2961
rect 50526 2887 50582 2896
rect 50344 2576 50396 2582
rect 50344 2518 50396 2524
rect 50356 1970 50384 2518
rect 50344 1964 50396 1970
rect 50344 1906 50396 1912
rect 50540 800 50568 2887
rect 50896 2576 50948 2582
rect 50896 2518 50948 2524
rect 50804 2440 50856 2446
rect 50804 2382 50856 2388
rect 50816 1834 50844 2382
rect 50804 1828 50856 1834
rect 50804 1770 50856 1776
rect 50908 1306 50936 2518
rect 50816 1278 50936 1306
rect 50816 800 50844 1278
rect 51092 800 51120 3878
rect 51276 1193 51304 4082
rect 51828 4049 51856 4082
rect 51814 4040 51870 4049
rect 51814 3975 51870 3984
rect 51908 4004 51960 4010
rect 51908 3946 51960 3952
rect 51518 3836 51826 3845
rect 51518 3834 51524 3836
rect 51580 3834 51604 3836
rect 51660 3834 51684 3836
rect 51740 3834 51764 3836
rect 51820 3834 51826 3836
rect 51580 3782 51582 3834
rect 51762 3782 51764 3834
rect 51518 3780 51524 3782
rect 51580 3780 51604 3782
rect 51660 3780 51684 3782
rect 51740 3780 51764 3782
rect 51820 3780 51826 3782
rect 51518 3771 51826 3780
rect 51356 3460 51408 3466
rect 51356 3402 51408 3408
rect 51262 1184 51318 1193
rect 51262 1119 51318 1128
rect 51368 800 51396 3402
rect 51518 2748 51826 2757
rect 51518 2746 51524 2748
rect 51580 2746 51604 2748
rect 51660 2746 51684 2748
rect 51740 2746 51764 2748
rect 51820 2746 51826 2748
rect 51580 2694 51582 2746
rect 51762 2694 51764 2746
rect 51518 2692 51524 2694
rect 51580 2692 51604 2694
rect 51660 2692 51684 2694
rect 51740 2692 51764 2694
rect 51820 2692 51826 2694
rect 51518 2683 51826 2692
rect 51448 2440 51500 2446
rect 51448 2382 51500 2388
rect 51460 2038 51488 2382
rect 51920 2088 51948 3946
rect 52288 3738 52316 6870
rect 52472 6866 52500 7754
rect 52736 7744 52788 7750
rect 52736 7686 52788 7692
rect 52460 6860 52512 6866
rect 52460 6802 52512 6808
rect 52472 5794 52500 6802
rect 52748 6662 52776 7686
rect 52828 7336 52880 7342
rect 52828 7278 52880 7284
rect 52840 6798 52868 7278
rect 52828 6792 52880 6798
rect 52828 6734 52880 6740
rect 52932 6662 52960 8298
rect 53104 7880 53156 7886
rect 53104 7822 53156 7828
rect 53116 7546 53144 7822
rect 53104 7540 53156 7546
rect 53104 7482 53156 7488
rect 52736 6656 52788 6662
rect 52736 6598 52788 6604
rect 52920 6656 52972 6662
rect 52920 6598 52972 6604
rect 52644 6316 52696 6322
rect 52644 6258 52696 6264
rect 52472 5778 52592 5794
rect 52472 5772 52604 5778
rect 52472 5766 52552 5772
rect 52552 5714 52604 5720
rect 52564 4622 52592 5714
rect 52656 5370 52684 6258
rect 53208 6202 53236 8298
rect 54208 7744 54260 7750
rect 54208 7686 54260 7692
rect 54220 7410 54248 7686
rect 54208 7404 54260 7410
rect 54208 7346 54260 7352
rect 54116 6860 54168 6866
rect 54116 6802 54168 6808
rect 54128 6254 54156 6802
rect 53024 6174 53236 6202
rect 54116 6248 54168 6254
rect 54116 6190 54168 6196
rect 52644 5364 52696 5370
rect 52644 5306 52696 5312
rect 53024 5030 53052 6174
rect 53104 6112 53156 6118
rect 53104 6054 53156 6060
rect 53116 5817 53144 6054
rect 53196 5840 53248 5846
rect 53102 5808 53158 5817
rect 53196 5782 53248 5788
rect 53102 5743 53158 5752
rect 53208 5166 53236 5782
rect 53840 5568 53892 5574
rect 53840 5510 53892 5516
rect 54208 5568 54260 5574
rect 54208 5510 54260 5516
rect 53288 5228 53340 5234
rect 53288 5170 53340 5176
rect 53196 5160 53248 5166
rect 53196 5102 53248 5108
rect 53012 5024 53064 5030
rect 53012 4966 53064 4972
rect 53300 4826 53328 5170
rect 53472 5160 53524 5166
rect 53472 5102 53524 5108
rect 53288 4820 53340 4826
rect 53288 4762 53340 4768
rect 52460 4616 52512 4622
rect 52460 4558 52512 4564
rect 52552 4616 52604 4622
rect 52552 4558 52604 4564
rect 53288 4616 53340 4622
rect 53288 4558 53340 4564
rect 52472 4049 52500 4558
rect 52458 4040 52514 4049
rect 52458 3975 52514 3984
rect 52276 3732 52328 3738
rect 52276 3674 52328 3680
rect 52552 3732 52604 3738
rect 52552 3674 52604 3680
rect 52368 3392 52420 3398
rect 52368 3334 52420 3340
rect 52380 3210 52408 3334
rect 51644 2060 51948 2088
rect 52012 3182 52408 3210
rect 51448 2032 51500 2038
rect 51448 1974 51500 1980
rect 51644 800 51672 2060
rect 52012 1850 52040 3182
rect 52368 3052 52420 3058
rect 52368 2994 52420 3000
rect 52184 2848 52236 2854
rect 52184 2790 52236 2796
rect 52090 2544 52146 2553
rect 52090 2479 52092 2488
rect 52144 2479 52146 2488
rect 52092 2450 52144 2456
rect 51920 1822 52040 1850
rect 51920 800 51948 1822
rect 52196 800 52224 2790
rect 52276 2440 52328 2446
rect 52276 2382 52328 2388
rect 52288 1698 52316 2382
rect 52276 1692 52328 1698
rect 52276 1634 52328 1640
rect 52380 800 52408 2994
rect 52460 2916 52512 2922
rect 52460 2858 52512 2864
rect 52472 800 52500 2858
rect 52564 800 52592 3674
rect 53300 3602 53328 4558
rect 53484 4010 53512 5102
rect 53564 4616 53616 4622
rect 53562 4584 53564 4593
rect 53616 4584 53618 4593
rect 53562 4519 53618 4528
rect 53576 4282 53604 4519
rect 53564 4276 53616 4282
rect 53564 4218 53616 4224
rect 53472 4004 53524 4010
rect 53472 3946 53524 3952
rect 53288 3596 53340 3602
rect 53288 3538 53340 3544
rect 52828 3528 52880 3534
rect 52828 3470 52880 3476
rect 53104 3528 53156 3534
rect 53104 3470 53156 3476
rect 52840 3194 52868 3470
rect 53116 3346 53144 3470
rect 52932 3318 53144 3346
rect 52828 3188 52880 3194
rect 52828 3130 52880 3136
rect 52932 3074 52960 3318
rect 52840 3058 52960 3074
rect 52828 3052 52960 3058
rect 52880 3046 52960 3052
rect 53104 3052 53156 3058
rect 52828 2994 52880 3000
rect 53104 2994 53156 3000
rect 53116 2774 53144 2994
rect 52656 2746 53144 2774
rect 52656 1290 52684 2746
rect 53300 2038 53328 3538
rect 53852 3074 53880 5510
rect 54220 5234 54248 5510
rect 54208 5228 54260 5234
rect 54208 5170 54260 5176
rect 54024 4140 54076 4146
rect 54024 4082 54076 4088
rect 54036 3670 54064 4082
rect 54024 3664 54076 3670
rect 54024 3606 54076 3612
rect 53932 3528 53984 3534
rect 53932 3470 53984 3476
rect 53760 3046 53880 3074
rect 53944 3058 53972 3470
rect 53932 3052 53984 3058
rect 53760 2802 53788 3046
rect 53932 2994 53984 3000
rect 53838 2952 53894 2961
rect 53838 2887 53840 2896
rect 53892 2887 53894 2896
rect 53840 2858 53892 2864
rect 53760 2774 53880 2802
rect 54036 2774 54064 3606
rect 54404 3534 54432 8366
rect 55312 8356 55364 8362
rect 55312 8298 55364 8304
rect 55324 7750 55352 8298
rect 55312 7744 55364 7750
rect 55312 7686 55364 7692
rect 55128 6248 55180 6254
rect 55128 6190 55180 6196
rect 54760 5228 54812 5234
rect 54760 5170 54812 5176
rect 54772 4826 54800 5170
rect 55140 5098 55168 6190
rect 55220 5704 55272 5710
rect 55220 5646 55272 5652
rect 55232 5166 55260 5646
rect 55324 5522 55352 7686
rect 55588 7336 55640 7342
rect 55588 7278 55640 7284
rect 55600 6662 55628 7278
rect 55680 6724 55732 6730
rect 55680 6666 55732 6672
rect 55588 6656 55640 6662
rect 55588 6598 55640 6604
rect 55600 6322 55628 6598
rect 55404 6316 55456 6322
rect 55404 6258 55456 6264
rect 55588 6316 55640 6322
rect 55588 6258 55640 6264
rect 55416 6118 55444 6258
rect 55404 6112 55456 6118
rect 55404 6054 55456 6060
rect 55600 5710 55628 6258
rect 55588 5704 55640 5710
rect 55588 5646 55640 5652
rect 55324 5494 55444 5522
rect 55220 5160 55272 5166
rect 55220 5102 55272 5108
rect 55128 5092 55180 5098
rect 55128 5034 55180 5040
rect 54760 4820 54812 4826
rect 54760 4762 54812 4768
rect 55140 4554 55168 5034
rect 55128 4548 55180 4554
rect 55128 4490 55180 4496
rect 55140 4010 55168 4490
rect 55232 4486 55260 5102
rect 55416 4486 55444 5494
rect 55496 4820 55548 4826
rect 55496 4762 55548 4768
rect 55220 4480 55272 4486
rect 55220 4422 55272 4428
rect 55404 4480 55456 4486
rect 55404 4422 55456 4428
rect 55218 4040 55274 4049
rect 55128 4004 55180 4010
rect 55218 3975 55220 3984
rect 55128 3946 55180 3952
rect 55272 3975 55274 3984
rect 55220 3946 55272 3952
rect 54576 3936 54628 3942
rect 54576 3878 54628 3884
rect 54588 3534 54616 3878
rect 55416 3670 55444 4422
rect 55508 4214 55536 4762
rect 55600 4622 55628 5646
rect 55692 5574 55720 6666
rect 55680 5568 55732 5574
rect 55680 5510 55732 5516
rect 55692 5370 55720 5510
rect 55680 5364 55732 5370
rect 55680 5306 55732 5312
rect 55588 4616 55640 4622
rect 55588 4558 55640 4564
rect 55496 4208 55548 4214
rect 55496 4150 55548 4156
rect 55692 4146 55720 5306
rect 55784 4758 55812 8434
rect 55864 7472 55916 7478
rect 55864 7414 55916 7420
rect 55876 7002 55904 7414
rect 56232 7404 56284 7410
rect 56284 7364 56364 7392
rect 56232 7346 56284 7352
rect 55864 6996 55916 7002
rect 55864 6938 55916 6944
rect 55876 5030 55904 6938
rect 56048 6656 56100 6662
rect 56048 6598 56100 6604
rect 56060 6390 56088 6598
rect 56048 6384 56100 6390
rect 56048 6326 56100 6332
rect 56336 6322 56364 7364
rect 57520 7336 57572 7342
rect 57520 7278 57572 7284
rect 57532 6798 57560 7278
rect 57796 7200 57848 7206
rect 57796 7142 57848 7148
rect 57980 7200 58032 7206
rect 57980 7142 58032 7148
rect 57808 6866 57836 7142
rect 57796 6860 57848 6866
rect 57796 6802 57848 6808
rect 57520 6792 57572 6798
rect 57520 6734 57572 6740
rect 56324 6316 56376 6322
rect 56324 6258 56376 6264
rect 55956 6248 56008 6254
rect 55956 6190 56008 6196
rect 55968 5642 55996 6190
rect 56336 6118 56364 6258
rect 56140 6112 56192 6118
rect 56140 6054 56192 6060
rect 56324 6112 56376 6118
rect 56324 6054 56376 6060
rect 55956 5636 56008 5642
rect 56008 5596 56088 5624
rect 55956 5578 56008 5584
rect 56060 5166 56088 5596
rect 56152 5234 56180 6054
rect 56336 5302 56364 6054
rect 57808 5778 57836 6802
rect 57992 6730 58020 7142
rect 57980 6724 58032 6730
rect 57980 6666 58032 6672
rect 57796 5772 57848 5778
rect 57796 5714 57848 5720
rect 57336 5704 57388 5710
rect 57336 5646 57388 5652
rect 57348 5370 57376 5646
rect 57336 5364 57388 5370
rect 57336 5306 57388 5312
rect 56324 5296 56376 5302
rect 56324 5238 56376 5244
rect 56140 5228 56192 5234
rect 56140 5170 56192 5176
rect 56048 5160 56100 5166
rect 56048 5102 56100 5108
rect 57704 5092 57756 5098
rect 57704 5034 57756 5040
rect 55864 5024 55916 5030
rect 55864 4966 55916 4972
rect 55772 4752 55824 4758
rect 55772 4694 55824 4700
rect 57716 4622 57744 5034
rect 57808 4690 57836 5714
rect 57980 5568 58032 5574
rect 57980 5510 58032 5516
rect 57796 4684 57848 4690
rect 57796 4626 57848 4632
rect 55956 4616 56008 4622
rect 55956 4558 56008 4564
rect 57704 4616 57756 4622
rect 57704 4558 57756 4564
rect 55968 4146 55996 4558
rect 57888 4480 57940 4486
rect 57888 4422 57940 4428
rect 57900 4146 57928 4422
rect 57992 4282 58020 5510
rect 58072 5228 58124 5234
rect 58072 5170 58124 5176
rect 58084 4826 58112 5170
rect 58072 4820 58124 4826
rect 58072 4762 58124 4768
rect 57980 4276 58032 4282
rect 57980 4218 58032 4224
rect 55680 4140 55732 4146
rect 55680 4082 55732 4088
rect 55956 4140 56008 4146
rect 55956 4082 56008 4088
rect 57888 4140 57940 4146
rect 57888 4082 57940 4088
rect 56508 3936 56560 3942
rect 56508 3878 56560 3884
rect 57796 3936 57848 3942
rect 57796 3878 57848 3884
rect 56520 3738 56548 3878
rect 57808 3738 57836 3878
rect 56508 3732 56560 3738
rect 56508 3674 56560 3680
rect 57796 3732 57848 3738
rect 57796 3674 57848 3680
rect 55404 3664 55456 3670
rect 55404 3606 55456 3612
rect 54392 3528 54444 3534
rect 54392 3470 54444 3476
rect 54576 3528 54628 3534
rect 54576 3470 54628 3476
rect 54114 3088 54170 3097
rect 54114 3023 54116 3032
rect 54168 3023 54170 3032
rect 54760 3052 54812 3058
rect 54116 2994 54168 3000
rect 54760 2994 54812 3000
rect 53380 2440 53432 2446
rect 53380 2382 53432 2388
rect 53392 2106 53420 2382
rect 53380 2100 53432 2106
rect 53380 2042 53432 2048
rect 53288 2032 53340 2038
rect 53288 1974 53340 1980
rect 53300 1358 53328 1974
rect 53852 1766 53880 2774
rect 53944 2746 54064 2774
rect 53840 1760 53892 1766
rect 53840 1702 53892 1708
rect 53944 1601 53972 2746
rect 54024 2440 54076 2446
rect 54024 2382 54076 2388
rect 54036 1902 54064 2382
rect 54668 2304 54720 2310
rect 54668 2246 54720 2252
rect 54024 1896 54076 1902
rect 54024 1838 54076 1844
rect 54680 1766 54708 2246
rect 54668 1760 54720 1766
rect 54668 1702 54720 1708
rect 53930 1592 53986 1601
rect 53930 1527 53986 1536
rect 54772 1494 54800 2994
rect 56520 2774 56548 3674
rect 57808 3194 57836 3674
rect 57796 3188 57848 3194
rect 57796 3130 57848 3136
rect 56428 2746 56548 2774
rect 57808 2774 57836 3130
rect 57808 2746 57928 2774
rect 56428 1970 56456 2746
rect 57900 2650 57928 2746
rect 57888 2644 57940 2650
rect 57888 2586 57940 2592
rect 57888 2304 57940 2310
rect 57888 2246 57940 2252
rect 57900 2038 57928 2246
rect 57888 2032 57940 2038
rect 57888 1974 57940 1980
rect 56416 1964 56468 1970
rect 56416 1906 56468 1912
rect 54760 1488 54812 1494
rect 54760 1430 54812 1436
rect 53288 1352 53340 1358
rect 53288 1294 53340 1300
rect 52644 1284 52696 1290
rect 52644 1226 52696 1232
rect 7196 740 7248 746
rect 7196 682 7248 688
rect 7286 0 7342 800
rect 7378 0 7434 800
rect 7470 0 7526 800
rect 7562 0 7618 800
rect 7654 0 7710 800
rect 7746 0 7802 800
rect 7838 0 7894 800
rect 7930 0 7986 800
rect 8022 0 8078 800
rect 8114 0 8170 800
rect 8206 0 8262 800
rect 8298 0 8354 800
rect 8390 0 8446 800
rect 8482 0 8538 800
rect 8574 0 8630 800
rect 8666 0 8722 800
rect 8758 0 8814 800
rect 8850 0 8906 800
rect 8942 0 8998 800
rect 9034 0 9090 800
rect 9126 0 9182 800
rect 9218 0 9274 800
rect 9310 0 9366 800
rect 9402 0 9458 800
rect 9494 0 9550 800
rect 9586 0 9642 800
rect 9678 0 9734 800
rect 9770 0 9826 800
rect 9862 0 9918 800
rect 9954 0 10010 800
rect 10046 0 10102 800
rect 10138 0 10194 800
rect 10230 0 10286 800
rect 10322 0 10378 800
rect 10414 0 10470 800
rect 10506 0 10562 800
rect 10598 0 10654 800
rect 10690 0 10746 800
rect 10782 0 10838 800
rect 10874 0 10930 800
rect 10966 0 11022 800
rect 11058 0 11114 800
rect 11150 0 11206 800
rect 11242 0 11298 800
rect 11334 0 11390 800
rect 11426 0 11482 800
rect 11518 0 11574 800
rect 11610 0 11666 800
rect 11702 0 11758 800
rect 11794 0 11850 800
rect 11886 0 11942 800
rect 11978 0 12034 800
rect 12070 0 12126 800
rect 12162 0 12218 800
rect 12254 0 12310 800
rect 12346 0 12402 800
rect 12438 0 12494 800
rect 12530 0 12586 800
rect 12622 0 12678 800
rect 12714 0 12770 800
rect 12806 0 12862 800
rect 12898 0 12954 800
rect 12990 0 13046 800
rect 13082 0 13138 800
rect 13174 0 13230 800
rect 13266 0 13322 800
rect 13358 0 13414 800
rect 13450 0 13506 800
rect 13542 0 13598 800
rect 13634 0 13690 800
rect 13726 0 13782 800
rect 13818 0 13874 800
rect 13910 0 13966 800
rect 14002 0 14058 800
rect 14094 0 14150 800
rect 14186 0 14242 800
rect 14278 0 14334 800
rect 14370 0 14426 800
rect 14462 0 14518 800
rect 14554 0 14610 800
rect 14646 0 14702 800
rect 14738 0 14794 800
rect 14830 0 14886 800
rect 14922 0 14978 800
rect 15014 0 15070 800
rect 15106 0 15162 800
rect 15198 0 15254 800
rect 15290 0 15346 800
rect 15382 0 15438 800
rect 15474 0 15530 800
rect 15566 0 15622 800
rect 15658 0 15714 800
rect 15750 0 15806 800
rect 15842 0 15898 800
rect 15934 0 15990 800
rect 16026 0 16082 800
rect 16118 0 16174 800
rect 16210 0 16266 800
rect 16302 0 16358 800
rect 16394 0 16450 800
rect 16486 0 16542 800
rect 16578 0 16634 800
rect 16670 0 16726 800
rect 16762 0 16818 800
rect 16854 0 16910 800
rect 16946 0 17002 800
rect 17038 0 17094 800
rect 17130 0 17186 800
rect 17222 0 17278 800
rect 17314 0 17370 800
rect 17406 0 17462 800
rect 17498 0 17554 800
rect 17590 0 17646 800
rect 17682 0 17738 800
rect 17774 0 17830 800
rect 17866 0 17922 800
rect 17958 0 18014 800
rect 18050 0 18106 800
rect 18142 0 18198 800
rect 18234 0 18290 800
rect 18326 0 18382 800
rect 18418 0 18474 800
rect 18510 0 18566 800
rect 18602 0 18658 800
rect 18694 0 18750 800
rect 18786 0 18842 800
rect 18878 0 18934 800
rect 18970 0 19026 800
rect 19062 0 19118 800
rect 19154 0 19210 800
rect 19246 0 19302 800
rect 19338 0 19394 800
rect 19430 0 19486 800
rect 19522 0 19578 800
rect 19614 0 19670 800
rect 19706 0 19762 800
rect 19798 0 19854 800
rect 19890 0 19946 800
rect 19982 0 20038 800
rect 20074 0 20130 800
rect 20166 0 20222 800
rect 20258 0 20314 800
rect 20350 0 20406 800
rect 20442 0 20498 800
rect 20534 0 20590 800
rect 20626 0 20682 800
rect 20718 0 20774 800
rect 20810 0 20866 800
rect 20902 0 20958 800
rect 20994 0 21050 800
rect 21086 0 21142 800
rect 21178 0 21234 800
rect 21270 0 21326 800
rect 21362 0 21418 800
rect 21454 0 21510 800
rect 21546 0 21602 800
rect 21638 0 21694 800
rect 21730 0 21786 800
rect 21822 0 21878 800
rect 21914 0 21970 800
rect 22006 0 22062 800
rect 22098 0 22154 800
rect 22190 0 22246 800
rect 22282 0 22338 800
rect 22374 0 22430 800
rect 22466 0 22522 800
rect 22558 0 22614 800
rect 22650 0 22706 800
rect 22742 0 22798 800
rect 22834 0 22890 800
rect 22926 0 22982 800
rect 23018 0 23074 800
rect 23110 0 23166 800
rect 23202 0 23258 800
rect 23294 0 23350 800
rect 23386 0 23442 800
rect 23478 0 23534 800
rect 23570 0 23626 800
rect 23662 0 23718 800
rect 23754 0 23810 800
rect 23846 0 23902 800
rect 23938 0 23994 800
rect 24030 0 24086 800
rect 24122 0 24178 800
rect 24214 0 24270 800
rect 24306 0 24362 800
rect 24398 0 24454 800
rect 24490 0 24546 800
rect 24582 0 24638 800
rect 24674 0 24730 800
rect 24766 0 24822 800
rect 24858 0 24914 800
rect 24950 0 25006 800
rect 25042 0 25098 800
rect 25134 0 25190 800
rect 25226 0 25282 800
rect 25318 0 25374 800
rect 25410 0 25466 800
rect 25502 0 25558 800
rect 25594 0 25650 800
rect 25686 0 25742 800
rect 25778 0 25834 800
rect 25870 0 25926 800
rect 25962 0 26018 800
rect 26054 0 26110 800
rect 26146 0 26202 800
rect 26238 0 26294 800
rect 26330 0 26386 800
rect 26422 0 26478 800
rect 26514 0 26570 800
rect 26606 0 26662 800
rect 26698 0 26754 800
rect 26790 0 26846 800
rect 26882 0 26938 800
rect 26974 0 27030 800
rect 27066 0 27122 800
rect 27158 0 27214 800
rect 27250 0 27306 800
rect 27342 0 27398 800
rect 27434 0 27490 800
rect 27526 0 27582 800
rect 27618 0 27674 800
rect 27710 0 27766 800
rect 27802 0 27858 800
rect 27894 0 27950 800
rect 27986 0 28042 800
rect 28078 0 28134 800
rect 28170 0 28226 800
rect 28262 0 28318 800
rect 28354 0 28410 800
rect 28446 0 28502 800
rect 28538 0 28594 800
rect 28630 0 28686 800
rect 28722 0 28778 800
rect 28814 0 28870 800
rect 28906 0 28962 800
rect 28998 0 29054 800
rect 29090 0 29146 800
rect 29182 0 29238 800
rect 29274 0 29330 800
rect 29366 0 29422 800
rect 29458 0 29514 800
rect 29550 0 29606 800
rect 29642 0 29698 800
rect 29734 0 29790 800
rect 29826 0 29882 800
rect 29918 0 29974 800
rect 30010 0 30066 800
rect 30102 0 30158 800
rect 30194 0 30250 800
rect 30286 0 30342 800
rect 30378 0 30434 800
rect 30470 0 30526 800
rect 30562 0 30618 800
rect 30654 0 30710 800
rect 30746 0 30802 800
rect 30838 0 30894 800
rect 30930 0 30986 800
rect 31022 0 31078 800
rect 31114 0 31170 800
rect 31206 0 31262 800
rect 31298 0 31354 800
rect 31390 0 31446 800
rect 31482 0 31538 800
rect 31574 0 31630 800
rect 31666 0 31722 800
rect 31758 0 31814 800
rect 31850 0 31906 800
rect 31942 0 31998 800
rect 32034 0 32090 800
rect 32126 0 32182 800
rect 32218 0 32274 800
rect 32310 0 32366 800
rect 32402 0 32458 800
rect 32494 0 32550 800
rect 32586 0 32642 800
rect 32678 0 32734 800
rect 32770 0 32826 800
rect 32862 0 32918 800
rect 32954 0 33010 800
rect 33046 0 33102 800
rect 33138 0 33194 800
rect 33230 0 33286 800
rect 33322 0 33378 800
rect 33414 0 33470 800
rect 33506 0 33562 800
rect 33598 0 33654 800
rect 33690 0 33746 800
rect 33782 0 33838 800
rect 33874 0 33930 800
rect 33966 0 34022 800
rect 34058 0 34114 800
rect 34150 0 34206 800
rect 34242 0 34298 800
rect 34334 0 34390 800
rect 34426 0 34482 800
rect 34518 0 34574 800
rect 34610 0 34666 800
rect 34702 0 34758 800
rect 34794 0 34850 800
rect 34886 0 34942 800
rect 34978 0 35034 800
rect 35070 0 35126 800
rect 35162 0 35218 800
rect 35254 0 35310 800
rect 35346 0 35402 800
rect 35438 0 35494 800
rect 35530 0 35586 800
rect 35622 0 35678 800
rect 35714 0 35770 800
rect 35806 0 35862 800
rect 35898 0 35954 800
rect 35990 0 36046 800
rect 36082 0 36138 800
rect 36174 0 36230 800
rect 36266 0 36322 800
rect 36358 0 36414 800
rect 36450 0 36506 800
rect 36542 0 36598 800
rect 36634 0 36690 800
rect 36726 0 36782 800
rect 36818 0 36874 800
rect 36910 0 36966 800
rect 37002 0 37058 800
rect 37094 0 37150 800
rect 37186 0 37242 800
rect 37278 0 37334 800
rect 37370 0 37426 800
rect 37462 0 37518 800
rect 37554 0 37610 800
rect 37646 0 37702 800
rect 37738 0 37794 800
rect 37830 0 37886 800
rect 37922 0 37978 800
rect 38014 0 38070 800
rect 38106 0 38162 800
rect 38198 0 38254 800
rect 38290 0 38346 800
rect 38382 0 38438 800
rect 38474 0 38530 800
rect 38566 0 38622 800
rect 38658 0 38714 800
rect 38750 0 38806 800
rect 38842 0 38898 800
rect 38934 0 38990 800
rect 39026 0 39082 800
rect 39118 0 39174 800
rect 39210 0 39266 800
rect 39302 0 39358 800
rect 39394 0 39450 800
rect 39486 0 39542 800
rect 39578 0 39634 800
rect 39670 0 39726 800
rect 39762 0 39818 800
rect 39854 0 39910 800
rect 39946 0 40002 800
rect 40038 0 40094 800
rect 40130 0 40186 800
rect 40222 0 40278 800
rect 40314 0 40370 800
rect 40406 0 40462 800
rect 40498 0 40554 800
rect 40590 0 40646 800
rect 40682 0 40738 800
rect 40774 0 40830 800
rect 40866 0 40922 800
rect 40958 0 41014 800
rect 41050 0 41106 800
rect 41142 0 41198 800
rect 41234 0 41290 800
rect 41326 0 41382 800
rect 41418 0 41474 800
rect 41510 0 41566 800
rect 41602 0 41658 800
rect 41694 0 41750 800
rect 41786 0 41842 800
rect 41878 0 41934 800
rect 41970 0 42026 800
rect 42062 0 42118 800
rect 42154 0 42210 800
rect 42246 0 42302 800
rect 42338 0 42394 800
rect 42430 0 42486 800
rect 42522 0 42578 800
rect 42614 0 42670 800
rect 42706 0 42762 800
rect 42798 0 42854 800
rect 42890 0 42946 800
rect 42982 0 43038 800
rect 43074 0 43130 800
rect 43166 0 43222 800
rect 43258 0 43314 800
rect 43350 0 43406 800
rect 43442 0 43498 800
rect 43534 0 43590 800
rect 43626 0 43682 800
rect 43718 0 43774 800
rect 43810 0 43866 800
rect 43902 0 43958 800
rect 43994 0 44050 800
rect 44086 0 44142 800
rect 44178 0 44234 800
rect 44270 0 44326 800
rect 44362 0 44418 800
rect 44454 0 44510 800
rect 44546 0 44602 800
rect 44638 0 44694 800
rect 44730 0 44786 800
rect 44822 0 44878 800
rect 44914 0 44970 800
rect 45006 0 45062 800
rect 45098 0 45154 800
rect 45190 0 45246 800
rect 45282 0 45338 800
rect 45374 0 45430 800
rect 45466 0 45522 800
rect 45558 0 45614 800
rect 45650 0 45706 800
rect 45742 0 45798 800
rect 45834 0 45890 800
rect 45926 0 45982 800
rect 46018 0 46074 800
rect 46110 0 46166 800
rect 46202 0 46258 800
rect 46294 0 46350 800
rect 46386 0 46442 800
rect 46478 0 46534 800
rect 46570 0 46626 800
rect 46662 0 46718 800
rect 46754 0 46810 800
rect 46846 0 46902 800
rect 46938 0 46994 800
rect 47030 0 47086 800
rect 47122 0 47178 800
rect 47214 0 47270 800
rect 47306 0 47362 800
rect 47398 0 47454 800
rect 47490 0 47546 800
rect 47582 0 47638 800
rect 47674 0 47730 800
rect 47766 0 47822 800
rect 47858 0 47914 800
rect 47950 0 48006 800
rect 48042 0 48098 800
rect 48134 0 48190 800
rect 48226 0 48282 800
rect 48318 0 48374 800
rect 48410 0 48466 800
rect 48502 0 48558 800
rect 48594 0 48650 800
rect 48686 0 48742 800
rect 48778 0 48834 800
rect 48870 0 48926 800
rect 48962 0 49018 800
rect 49054 0 49110 800
rect 49146 0 49202 800
rect 49238 0 49294 800
rect 49330 0 49386 800
rect 49422 0 49478 800
rect 49514 0 49570 800
rect 49606 0 49662 800
rect 49698 0 49754 800
rect 49790 0 49846 800
rect 49882 0 49938 800
rect 49974 0 50030 800
rect 50066 0 50122 800
rect 50158 0 50214 800
rect 50250 0 50306 800
rect 50342 0 50398 800
rect 50434 0 50490 800
rect 50526 0 50582 800
rect 50618 0 50674 800
rect 50710 0 50766 800
rect 50802 0 50858 800
rect 50894 0 50950 800
rect 50986 0 51042 800
rect 51078 0 51134 800
rect 51170 0 51226 800
rect 51262 0 51318 800
rect 51354 0 51410 800
rect 51446 0 51502 800
rect 51538 0 51594 800
rect 51630 0 51686 800
rect 51722 0 51778 800
rect 51814 0 51870 800
rect 51906 0 51962 800
rect 51998 0 52054 800
rect 52090 0 52146 800
rect 52182 0 52238 800
rect 52274 0 52330 800
rect 52366 0 52422 800
rect 52458 0 52514 800
rect 52550 0 52606 800
<< via2 >>
rect 8180 16890 8236 16892
rect 8260 16890 8316 16892
rect 8340 16890 8396 16892
rect 8420 16890 8476 16892
rect 8180 16838 8226 16890
rect 8226 16838 8236 16890
rect 8260 16838 8290 16890
rect 8290 16838 8302 16890
rect 8302 16838 8316 16890
rect 8340 16838 8354 16890
rect 8354 16838 8366 16890
rect 8366 16838 8396 16890
rect 8420 16838 8430 16890
rect 8430 16838 8476 16890
rect 8180 16836 8236 16838
rect 8260 16836 8316 16838
rect 8340 16836 8396 16838
rect 8420 16836 8476 16838
rect 15404 17434 15460 17436
rect 15484 17434 15540 17436
rect 15564 17434 15620 17436
rect 15644 17434 15700 17436
rect 15404 17382 15450 17434
rect 15450 17382 15460 17434
rect 15484 17382 15514 17434
rect 15514 17382 15526 17434
rect 15526 17382 15540 17434
rect 15564 17382 15578 17434
rect 15578 17382 15590 17434
rect 15590 17382 15620 17434
rect 15644 17382 15654 17434
rect 15654 17382 15700 17434
rect 15404 17380 15460 17382
rect 15484 17380 15540 17382
rect 15564 17380 15620 17382
rect 15644 17380 15700 17382
rect 22628 16890 22684 16892
rect 22708 16890 22764 16892
rect 22788 16890 22844 16892
rect 22868 16890 22924 16892
rect 22628 16838 22674 16890
rect 22674 16838 22684 16890
rect 22708 16838 22738 16890
rect 22738 16838 22750 16890
rect 22750 16838 22764 16890
rect 22788 16838 22802 16890
rect 22802 16838 22814 16890
rect 22814 16838 22844 16890
rect 22868 16838 22878 16890
rect 22878 16838 22924 16890
rect 22628 16836 22684 16838
rect 22708 16836 22764 16838
rect 22788 16836 22844 16838
rect 22868 16836 22924 16838
rect 29852 17434 29908 17436
rect 29932 17434 29988 17436
rect 30012 17434 30068 17436
rect 30092 17434 30148 17436
rect 29852 17382 29898 17434
rect 29898 17382 29908 17434
rect 29932 17382 29962 17434
rect 29962 17382 29974 17434
rect 29974 17382 29988 17434
rect 30012 17382 30026 17434
rect 30026 17382 30038 17434
rect 30038 17382 30068 17434
rect 30092 17382 30102 17434
rect 30102 17382 30148 17434
rect 29852 17380 29908 17382
rect 29932 17380 29988 17382
rect 30012 17380 30068 17382
rect 30092 17380 30148 17382
rect 37076 16890 37132 16892
rect 37156 16890 37212 16892
rect 37236 16890 37292 16892
rect 37316 16890 37372 16892
rect 37076 16838 37122 16890
rect 37122 16838 37132 16890
rect 37156 16838 37186 16890
rect 37186 16838 37198 16890
rect 37198 16838 37212 16890
rect 37236 16838 37250 16890
rect 37250 16838 37262 16890
rect 37262 16838 37292 16890
rect 37316 16838 37326 16890
rect 37326 16838 37372 16890
rect 37076 16836 37132 16838
rect 37156 16836 37212 16838
rect 37236 16836 37292 16838
rect 37316 16836 37372 16838
rect 44300 17434 44356 17436
rect 44380 17434 44436 17436
rect 44460 17434 44516 17436
rect 44540 17434 44596 17436
rect 44300 17382 44346 17434
rect 44346 17382 44356 17434
rect 44380 17382 44410 17434
rect 44410 17382 44422 17434
rect 44422 17382 44436 17434
rect 44460 17382 44474 17434
rect 44474 17382 44486 17434
rect 44486 17382 44516 17434
rect 44540 17382 44550 17434
rect 44550 17382 44596 17434
rect 44300 17380 44356 17382
rect 44380 17380 44436 17382
rect 44460 17380 44516 17382
rect 44540 17380 44596 17382
rect 51524 16890 51580 16892
rect 51604 16890 51660 16892
rect 51684 16890 51740 16892
rect 51764 16890 51820 16892
rect 51524 16838 51570 16890
rect 51570 16838 51580 16890
rect 51604 16838 51634 16890
rect 51634 16838 51646 16890
rect 51646 16838 51660 16890
rect 51684 16838 51698 16890
rect 51698 16838 51710 16890
rect 51710 16838 51740 16890
rect 51764 16838 51774 16890
rect 51774 16838 51820 16890
rect 51524 16836 51580 16838
rect 51604 16836 51660 16838
rect 51684 16836 51740 16838
rect 51764 16836 51820 16838
rect 15404 16346 15460 16348
rect 15484 16346 15540 16348
rect 15564 16346 15620 16348
rect 15644 16346 15700 16348
rect 15404 16294 15450 16346
rect 15450 16294 15460 16346
rect 15484 16294 15514 16346
rect 15514 16294 15526 16346
rect 15526 16294 15540 16346
rect 15564 16294 15578 16346
rect 15578 16294 15590 16346
rect 15590 16294 15620 16346
rect 15644 16294 15654 16346
rect 15654 16294 15700 16346
rect 15404 16292 15460 16294
rect 15484 16292 15540 16294
rect 15564 16292 15620 16294
rect 15644 16292 15700 16294
rect 29852 16346 29908 16348
rect 29932 16346 29988 16348
rect 30012 16346 30068 16348
rect 30092 16346 30148 16348
rect 29852 16294 29898 16346
rect 29898 16294 29908 16346
rect 29932 16294 29962 16346
rect 29962 16294 29974 16346
rect 29974 16294 29988 16346
rect 30012 16294 30026 16346
rect 30026 16294 30038 16346
rect 30038 16294 30068 16346
rect 30092 16294 30102 16346
rect 30102 16294 30148 16346
rect 29852 16292 29908 16294
rect 29932 16292 29988 16294
rect 30012 16292 30068 16294
rect 30092 16292 30148 16294
rect 44300 16346 44356 16348
rect 44380 16346 44436 16348
rect 44460 16346 44516 16348
rect 44540 16346 44596 16348
rect 44300 16294 44346 16346
rect 44346 16294 44356 16346
rect 44380 16294 44410 16346
rect 44410 16294 44422 16346
rect 44422 16294 44436 16346
rect 44460 16294 44474 16346
rect 44474 16294 44486 16346
rect 44486 16294 44516 16346
rect 44540 16294 44550 16346
rect 44550 16294 44596 16346
rect 44300 16292 44356 16294
rect 44380 16292 44436 16294
rect 44460 16292 44516 16294
rect 44540 16292 44596 16294
rect 8180 15802 8236 15804
rect 8260 15802 8316 15804
rect 8340 15802 8396 15804
rect 8420 15802 8476 15804
rect 8180 15750 8226 15802
rect 8226 15750 8236 15802
rect 8260 15750 8290 15802
rect 8290 15750 8302 15802
rect 8302 15750 8316 15802
rect 8340 15750 8354 15802
rect 8354 15750 8366 15802
rect 8366 15750 8396 15802
rect 8420 15750 8430 15802
rect 8430 15750 8476 15802
rect 8180 15748 8236 15750
rect 8260 15748 8316 15750
rect 8340 15748 8396 15750
rect 8420 15748 8476 15750
rect 22628 15802 22684 15804
rect 22708 15802 22764 15804
rect 22788 15802 22844 15804
rect 22868 15802 22924 15804
rect 22628 15750 22674 15802
rect 22674 15750 22684 15802
rect 22708 15750 22738 15802
rect 22738 15750 22750 15802
rect 22750 15750 22764 15802
rect 22788 15750 22802 15802
rect 22802 15750 22814 15802
rect 22814 15750 22844 15802
rect 22868 15750 22878 15802
rect 22878 15750 22924 15802
rect 22628 15748 22684 15750
rect 22708 15748 22764 15750
rect 22788 15748 22844 15750
rect 22868 15748 22924 15750
rect 37076 15802 37132 15804
rect 37156 15802 37212 15804
rect 37236 15802 37292 15804
rect 37316 15802 37372 15804
rect 37076 15750 37122 15802
rect 37122 15750 37132 15802
rect 37156 15750 37186 15802
rect 37186 15750 37198 15802
rect 37198 15750 37212 15802
rect 37236 15750 37250 15802
rect 37250 15750 37262 15802
rect 37262 15750 37292 15802
rect 37316 15750 37326 15802
rect 37326 15750 37372 15802
rect 37076 15748 37132 15750
rect 37156 15748 37212 15750
rect 37236 15748 37292 15750
rect 37316 15748 37372 15750
rect 51524 15802 51580 15804
rect 51604 15802 51660 15804
rect 51684 15802 51740 15804
rect 51764 15802 51820 15804
rect 51524 15750 51570 15802
rect 51570 15750 51580 15802
rect 51604 15750 51634 15802
rect 51634 15750 51646 15802
rect 51646 15750 51660 15802
rect 51684 15750 51698 15802
rect 51698 15750 51710 15802
rect 51710 15750 51740 15802
rect 51764 15750 51774 15802
rect 51774 15750 51820 15802
rect 51524 15748 51580 15750
rect 51604 15748 51660 15750
rect 51684 15748 51740 15750
rect 51764 15748 51820 15750
rect 15404 15258 15460 15260
rect 15484 15258 15540 15260
rect 15564 15258 15620 15260
rect 15644 15258 15700 15260
rect 15404 15206 15450 15258
rect 15450 15206 15460 15258
rect 15484 15206 15514 15258
rect 15514 15206 15526 15258
rect 15526 15206 15540 15258
rect 15564 15206 15578 15258
rect 15578 15206 15590 15258
rect 15590 15206 15620 15258
rect 15644 15206 15654 15258
rect 15654 15206 15700 15258
rect 15404 15204 15460 15206
rect 15484 15204 15540 15206
rect 15564 15204 15620 15206
rect 15644 15204 15700 15206
rect 29852 15258 29908 15260
rect 29932 15258 29988 15260
rect 30012 15258 30068 15260
rect 30092 15258 30148 15260
rect 29852 15206 29898 15258
rect 29898 15206 29908 15258
rect 29932 15206 29962 15258
rect 29962 15206 29974 15258
rect 29974 15206 29988 15258
rect 30012 15206 30026 15258
rect 30026 15206 30038 15258
rect 30038 15206 30068 15258
rect 30092 15206 30102 15258
rect 30102 15206 30148 15258
rect 29852 15204 29908 15206
rect 29932 15204 29988 15206
rect 30012 15204 30068 15206
rect 30092 15204 30148 15206
rect 44300 15258 44356 15260
rect 44380 15258 44436 15260
rect 44460 15258 44516 15260
rect 44540 15258 44596 15260
rect 44300 15206 44346 15258
rect 44346 15206 44356 15258
rect 44380 15206 44410 15258
rect 44410 15206 44422 15258
rect 44422 15206 44436 15258
rect 44460 15206 44474 15258
rect 44474 15206 44486 15258
rect 44486 15206 44516 15258
rect 44540 15206 44550 15258
rect 44550 15206 44596 15258
rect 44300 15204 44356 15206
rect 44380 15204 44436 15206
rect 44460 15204 44516 15206
rect 44540 15204 44596 15206
rect 8180 14714 8236 14716
rect 8260 14714 8316 14716
rect 8340 14714 8396 14716
rect 8420 14714 8476 14716
rect 8180 14662 8226 14714
rect 8226 14662 8236 14714
rect 8260 14662 8290 14714
rect 8290 14662 8302 14714
rect 8302 14662 8316 14714
rect 8340 14662 8354 14714
rect 8354 14662 8366 14714
rect 8366 14662 8396 14714
rect 8420 14662 8430 14714
rect 8430 14662 8476 14714
rect 8180 14660 8236 14662
rect 8260 14660 8316 14662
rect 8340 14660 8396 14662
rect 8420 14660 8476 14662
rect 22628 14714 22684 14716
rect 22708 14714 22764 14716
rect 22788 14714 22844 14716
rect 22868 14714 22924 14716
rect 22628 14662 22674 14714
rect 22674 14662 22684 14714
rect 22708 14662 22738 14714
rect 22738 14662 22750 14714
rect 22750 14662 22764 14714
rect 22788 14662 22802 14714
rect 22802 14662 22814 14714
rect 22814 14662 22844 14714
rect 22868 14662 22878 14714
rect 22878 14662 22924 14714
rect 22628 14660 22684 14662
rect 22708 14660 22764 14662
rect 22788 14660 22844 14662
rect 22868 14660 22924 14662
rect 37076 14714 37132 14716
rect 37156 14714 37212 14716
rect 37236 14714 37292 14716
rect 37316 14714 37372 14716
rect 37076 14662 37122 14714
rect 37122 14662 37132 14714
rect 37156 14662 37186 14714
rect 37186 14662 37198 14714
rect 37198 14662 37212 14714
rect 37236 14662 37250 14714
rect 37250 14662 37262 14714
rect 37262 14662 37292 14714
rect 37316 14662 37326 14714
rect 37326 14662 37372 14714
rect 37076 14660 37132 14662
rect 37156 14660 37212 14662
rect 37236 14660 37292 14662
rect 37316 14660 37372 14662
rect 51524 14714 51580 14716
rect 51604 14714 51660 14716
rect 51684 14714 51740 14716
rect 51764 14714 51820 14716
rect 51524 14662 51570 14714
rect 51570 14662 51580 14714
rect 51604 14662 51634 14714
rect 51634 14662 51646 14714
rect 51646 14662 51660 14714
rect 51684 14662 51698 14714
rect 51698 14662 51710 14714
rect 51710 14662 51740 14714
rect 51764 14662 51774 14714
rect 51774 14662 51820 14714
rect 51524 14660 51580 14662
rect 51604 14660 51660 14662
rect 51684 14660 51740 14662
rect 51764 14660 51820 14662
rect 15404 14170 15460 14172
rect 15484 14170 15540 14172
rect 15564 14170 15620 14172
rect 15644 14170 15700 14172
rect 15404 14118 15450 14170
rect 15450 14118 15460 14170
rect 15484 14118 15514 14170
rect 15514 14118 15526 14170
rect 15526 14118 15540 14170
rect 15564 14118 15578 14170
rect 15578 14118 15590 14170
rect 15590 14118 15620 14170
rect 15644 14118 15654 14170
rect 15654 14118 15700 14170
rect 15404 14116 15460 14118
rect 15484 14116 15540 14118
rect 15564 14116 15620 14118
rect 15644 14116 15700 14118
rect 29852 14170 29908 14172
rect 29932 14170 29988 14172
rect 30012 14170 30068 14172
rect 30092 14170 30148 14172
rect 29852 14118 29898 14170
rect 29898 14118 29908 14170
rect 29932 14118 29962 14170
rect 29962 14118 29974 14170
rect 29974 14118 29988 14170
rect 30012 14118 30026 14170
rect 30026 14118 30038 14170
rect 30038 14118 30068 14170
rect 30092 14118 30102 14170
rect 30102 14118 30148 14170
rect 29852 14116 29908 14118
rect 29932 14116 29988 14118
rect 30012 14116 30068 14118
rect 30092 14116 30148 14118
rect 44300 14170 44356 14172
rect 44380 14170 44436 14172
rect 44460 14170 44516 14172
rect 44540 14170 44596 14172
rect 44300 14118 44346 14170
rect 44346 14118 44356 14170
rect 44380 14118 44410 14170
rect 44410 14118 44422 14170
rect 44422 14118 44436 14170
rect 44460 14118 44474 14170
rect 44474 14118 44486 14170
rect 44486 14118 44516 14170
rect 44540 14118 44550 14170
rect 44550 14118 44596 14170
rect 44300 14116 44356 14118
rect 44380 14116 44436 14118
rect 44460 14116 44516 14118
rect 44540 14116 44596 14118
rect 13358 13812 13360 13832
rect 13360 13812 13412 13832
rect 13412 13812 13414 13832
rect 1950 12416 2006 12472
rect 1582 10512 1638 10568
rect 1766 11736 1822 11792
rect 2042 11228 2044 11248
rect 2044 11228 2096 11248
rect 2096 11228 2098 11248
rect 2042 11192 2098 11228
rect 13358 13776 13414 13812
rect 8180 13626 8236 13628
rect 8260 13626 8316 13628
rect 8340 13626 8396 13628
rect 8420 13626 8476 13628
rect 8180 13574 8226 13626
rect 8226 13574 8236 13626
rect 8260 13574 8290 13626
rect 8290 13574 8302 13626
rect 8302 13574 8316 13626
rect 8340 13574 8354 13626
rect 8354 13574 8366 13626
rect 8366 13574 8396 13626
rect 8420 13574 8430 13626
rect 8430 13574 8476 13626
rect 8180 13572 8236 13574
rect 8260 13572 8316 13574
rect 8340 13572 8396 13574
rect 8420 13572 8476 13574
rect 1858 9696 1914 9752
rect 1766 8336 1822 8392
rect 2502 9868 2504 9888
rect 2504 9868 2556 9888
rect 2556 9868 2558 9888
rect 2502 9832 2558 9868
rect 1582 4800 1638 4856
rect 1766 4256 1822 4312
rect 1858 4120 1914 4176
rect 2134 5072 2190 5128
rect 2226 2624 2282 2680
rect 2594 6432 2650 6488
rect 2502 4664 2558 4720
rect 2686 5344 2742 5400
rect 3146 7248 3202 7304
rect 3054 5636 3110 5672
rect 3054 5616 3056 5636
rect 3056 5616 3108 5636
rect 3108 5616 3110 5636
rect 3790 12416 3846 12472
rect 3422 5752 3478 5808
rect 4158 10104 4214 10160
rect 3698 6976 3754 7032
rect 3698 6296 3754 6352
rect 4158 7384 4214 7440
rect 4250 6316 4306 6352
rect 4250 6296 4252 6316
rect 4252 6296 4304 6316
rect 4304 6296 4306 6316
rect 4342 6196 4344 6216
rect 4344 6196 4396 6216
rect 4396 6196 4398 6216
rect 4342 6160 4398 6196
rect 3790 4256 3846 4312
rect 5078 9580 5134 9616
rect 5078 9560 5080 9580
rect 5080 9560 5132 9580
rect 5132 9560 5134 9580
rect 4250 3476 4252 3496
rect 4252 3476 4304 3496
rect 4304 3476 4306 3496
rect 4250 3440 4306 3476
rect 3974 1944 4030 2000
rect 3882 1672 3938 1728
rect 4894 4392 4950 4448
rect 5814 11500 5816 11520
rect 5816 11500 5868 11520
rect 5868 11500 5870 11520
rect 5814 11464 5870 11500
rect 5354 6196 5356 6216
rect 5356 6196 5408 6216
rect 5408 6196 5410 6216
rect 5354 6160 5410 6196
rect 4618 2896 4674 2952
rect 5078 3052 5134 3088
rect 5078 3032 5080 3052
rect 5080 3032 5132 3052
rect 5132 3032 5134 3052
rect 5446 3340 5448 3360
rect 5448 3340 5500 3360
rect 5500 3340 5502 3360
rect 5446 3304 5502 3340
rect 6090 8608 6146 8664
rect 6090 8336 6146 8392
rect 5998 7656 6054 7712
rect 5998 6976 6054 7032
rect 5814 6160 5870 6216
rect 5814 5092 5870 5128
rect 5814 5072 5816 5092
rect 5816 5072 5868 5092
rect 5868 5072 5870 5092
rect 5722 4936 5778 4992
rect 5722 4664 5778 4720
rect 5814 4004 5870 4040
rect 5814 3984 5816 4004
rect 5816 3984 5868 4004
rect 5868 3984 5870 4004
rect 6274 7520 6330 7576
rect 7010 12416 7066 12472
rect 8180 12538 8236 12540
rect 8260 12538 8316 12540
rect 8340 12538 8396 12540
rect 8420 12538 8476 12540
rect 8180 12486 8226 12538
rect 8226 12486 8236 12538
rect 8260 12486 8290 12538
rect 8290 12486 8302 12538
rect 8302 12486 8316 12538
rect 8340 12486 8354 12538
rect 8354 12486 8366 12538
rect 8366 12486 8396 12538
rect 8420 12486 8430 12538
rect 8430 12486 8476 12538
rect 8180 12484 8236 12486
rect 8260 12484 8316 12486
rect 8340 12484 8396 12486
rect 8420 12484 8476 12486
rect 6366 7404 6422 7440
rect 6366 7384 6368 7404
rect 6368 7384 6420 7404
rect 6420 7384 6422 7404
rect 6550 8336 6606 8392
rect 6182 5344 6238 5400
rect 6182 4700 6184 4720
rect 6184 4700 6236 4720
rect 6236 4700 6238 4720
rect 6182 4664 6238 4700
rect 6458 6976 6514 7032
rect 6366 5772 6422 5808
rect 6366 5752 6368 5772
rect 6368 5752 6420 5772
rect 6420 5752 6422 5772
rect 6274 4528 6330 4584
rect 6642 7792 6698 7848
rect 6642 7520 6698 7576
rect 6734 7384 6790 7440
rect 6550 6568 6606 6624
rect 6734 6332 6736 6352
rect 6736 6332 6788 6352
rect 6788 6332 6790 6352
rect 6734 6296 6790 6332
rect 6642 5616 6698 5672
rect 6550 4120 6606 4176
rect 6642 3848 6698 3904
rect 6918 4800 6974 4856
rect 6826 3576 6882 3632
rect 6642 2488 6698 2544
rect 6826 1808 6882 1864
rect 7286 5752 7342 5808
rect 7746 11056 7802 11112
rect 8180 11450 8236 11452
rect 8260 11450 8316 11452
rect 8340 11450 8396 11452
rect 8420 11450 8476 11452
rect 8180 11398 8226 11450
rect 8226 11398 8236 11450
rect 8260 11398 8290 11450
rect 8290 11398 8302 11450
rect 8302 11398 8316 11450
rect 8340 11398 8354 11450
rect 8354 11398 8366 11450
rect 8366 11398 8396 11450
rect 8420 11398 8430 11450
rect 8430 11398 8476 11450
rect 8180 11396 8236 11398
rect 8260 11396 8316 11398
rect 8340 11396 8396 11398
rect 8420 11396 8476 11398
rect 8180 10362 8236 10364
rect 8260 10362 8316 10364
rect 8340 10362 8396 10364
rect 8420 10362 8476 10364
rect 8180 10310 8226 10362
rect 8226 10310 8236 10362
rect 8260 10310 8290 10362
rect 8290 10310 8302 10362
rect 8302 10310 8316 10362
rect 8340 10310 8354 10362
rect 8354 10310 8366 10362
rect 8366 10310 8396 10362
rect 8420 10310 8430 10362
rect 8430 10310 8476 10362
rect 8180 10308 8236 10310
rect 8260 10308 8316 10310
rect 8340 10308 8396 10310
rect 8420 10308 8476 10310
rect 8180 9274 8236 9276
rect 8260 9274 8316 9276
rect 8340 9274 8396 9276
rect 8420 9274 8476 9276
rect 8180 9222 8226 9274
rect 8226 9222 8236 9274
rect 8260 9222 8290 9274
rect 8290 9222 8302 9274
rect 8302 9222 8316 9274
rect 8340 9222 8354 9274
rect 8354 9222 8366 9274
rect 8366 9222 8396 9274
rect 8420 9222 8430 9274
rect 8430 9222 8476 9274
rect 8180 9220 8236 9222
rect 8260 9220 8316 9222
rect 8340 9220 8396 9222
rect 8420 9220 8476 9222
rect 8206 8336 8262 8392
rect 8180 8186 8236 8188
rect 8260 8186 8316 8188
rect 8340 8186 8396 8188
rect 8420 8186 8476 8188
rect 8180 8134 8226 8186
rect 8226 8134 8236 8186
rect 8260 8134 8290 8186
rect 8290 8134 8302 8186
rect 8302 8134 8316 8186
rect 8340 8134 8354 8186
rect 8354 8134 8366 8186
rect 8366 8134 8396 8186
rect 8420 8134 8430 8186
rect 8430 8134 8476 8186
rect 8180 8132 8236 8134
rect 8260 8132 8316 8134
rect 8340 8132 8396 8134
rect 8420 8132 8476 8134
rect 8180 7098 8236 7100
rect 8260 7098 8316 7100
rect 8340 7098 8396 7100
rect 8420 7098 8476 7100
rect 8180 7046 8226 7098
rect 8226 7046 8236 7098
rect 8260 7046 8290 7098
rect 8290 7046 8302 7098
rect 8302 7046 8316 7098
rect 8340 7046 8354 7098
rect 8354 7046 8366 7098
rect 8366 7046 8396 7098
rect 8420 7046 8430 7098
rect 8430 7046 8476 7098
rect 8180 7044 8236 7046
rect 8260 7044 8316 7046
rect 8340 7044 8396 7046
rect 8420 7044 8476 7046
rect 7746 6296 7802 6352
rect 7746 5752 7802 5808
rect 7654 5652 7656 5672
rect 7656 5652 7708 5672
rect 7708 5652 7710 5672
rect 7654 5616 7710 5652
rect 7470 4120 7526 4176
rect 7470 3732 7526 3768
rect 7470 3712 7472 3732
rect 7472 3712 7524 3732
rect 7524 3712 7526 3732
rect 7378 3168 7434 3224
rect 7746 4392 7802 4448
rect 8574 6704 8630 6760
rect 8180 6010 8236 6012
rect 8260 6010 8316 6012
rect 8340 6010 8396 6012
rect 8420 6010 8476 6012
rect 8180 5958 8226 6010
rect 8226 5958 8236 6010
rect 8260 5958 8290 6010
rect 8290 5958 8302 6010
rect 8302 5958 8316 6010
rect 8340 5958 8354 6010
rect 8354 5958 8366 6010
rect 8366 5958 8396 6010
rect 8420 5958 8430 6010
rect 8430 5958 8476 6010
rect 8180 5956 8236 5958
rect 8260 5956 8316 5958
rect 8340 5956 8396 5958
rect 8420 5956 8476 5958
rect 8666 5888 8722 5944
rect 8206 5752 8262 5808
rect 8180 4922 8236 4924
rect 8260 4922 8316 4924
rect 8340 4922 8396 4924
rect 8420 4922 8476 4924
rect 8180 4870 8226 4922
rect 8226 4870 8236 4922
rect 8260 4870 8290 4922
rect 8290 4870 8302 4922
rect 8302 4870 8316 4922
rect 8340 4870 8354 4922
rect 8354 4870 8366 4922
rect 8366 4870 8396 4922
rect 8420 4870 8430 4922
rect 8430 4870 8476 4922
rect 8180 4868 8236 4870
rect 8260 4868 8316 4870
rect 8340 4868 8396 4870
rect 8420 4868 8476 4870
rect 8666 4800 8722 4856
rect 8574 4392 8630 4448
rect 8180 3834 8236 3836
rect 8260 3834 8316 3836
rect 8340 3834 8396 3836
rect 8420 3834 8476 3836
rect 8180 3782 8226 3834
rect 8226 3782 8236 3834
rect 8260 3782 8290 3834
rect 8290 3782 8302 3834
rect 8302 3782 8316 3834
rect 8340 3782 8354 3834
rect 8354 3782 8366 3834
rect 8366 3782 8396 3834
rect 8420 3782 8430 3834
rect 8430 3782 8476 3834
rect 8180 3780 8236 3782
rect 8260 3780 8316 3782
rect 8340 3780 8396 3782
rect 8420 3780 8476 3782
rect 8206 3168 8262 3224
rect 8666 3848 8722 3904
rect 10966 12588 10968 12608
rect 10968 12588 11020 12608
rect 11020 12588 11022 12608
rect 10966 12552 11022 12588
rect 8942 3712 8998 3768
rect 8758 3168 8814 3224
rect 8574 2760 8630 2816
rect 8180 2746 8236 2748
rect 8260 2746 8316 2748
rect 8340 2746 8396 2748
rect 8420 2746 8476 2748
rect 8180 2694 8226 2746
rect 8226 2694 8236 2746
rect 8260 2694 8290 2746
rect 8290 2694 8302 2746
rect 8302 2694 8316 2746
rect 8340 2694 8354 2746
rect 8354 2694 8366 2746
rect 8366 2694 8396 2746
rect 8420 2694 8430 2746
rect 8430 2694 8476 2746
rect 8180 2692 8236 2694
rect 8260 2692 8316 2694
rect 8340 2692 8396 2694
rect 8420 2692 8476 2694
rect 9218 7520 9274 7576
rect 9126 6432 9182 6488
rect 9034 2080 9090 2136
rect 9218 3304 9274 3360
rect 9218 2388 9220 2408
rect 9220 2388 9272 2408
rect 9272 2388 9274 2408
rect 9218 2352 9274 2388
rect 9494 8608 9550 8664
rect 9494 7284 9496 7304
rect 9496 7284 9548 7304
rect 9548 7284 9550 7304
rect 9494 7248 9550 7284
rect 9494 6840 9550 6896
rect 9770 9696 9826 9752
rect 9862 9580 9918 9616
rect 9862 9560 9864 9580
rect 9864 9560 9916 9580
rect 9916 9560 9918 9580
rect 9862 7928 9918 7984
rect 9770 6452 9826 6488
rect 9770 6432 9772 6452
rect 9772 6432 9824 6452
rect 9824 6432 9826 6452
rect 9770 6060 9772 6080
rect 9772 6060 9824 6080
rect 9824 6060 9826 6080
rect 9770 6024 9826 6060
rect 9494 5344 9550 5400
rect 9678 5344 9734 5400
rect 9862 4936 9918 4992
rect 10046 8064 10102 8120
rect 10046 5072 10102 5128
rect 10046 4800 10102 4856
rect 10322 9424 10378 9480
rect 10598 8916 10600 8936
rect 10600 8916 10652 8936
rect 10652 8916 10654 8936
rect 10598 8880 10654 8916
rect 10230 6024 10286 6080
rect 10230 5772 10286 5808
rect 10230 5752 10232 5772
rect 10232 5752 10284 5772
rect 10284 5752 10286 5772
rect 10322 5616 10378 5672
rect 10322 4528 10378 4584
rect 10506 3476 10508 3496
rect 10508 3476 10560 3496
rect 10560 3476 10562 3496
rect 10506 3440 10562 3476
rect 10966 8356 11022 8392
rect 10966 8336 10968 8356
rect 10968 8336 11020 8356
rect 11020 8336 11022 8356
rect 10874 7656 10930 7712
rect 10874 7248 10930 7304
rect 10874 6024 10930 6080
rect 10230 2624 10286 2680
rect 10690 2896 10746 2952
rect 10690 992 10746 1048
rect 11426 12724 11428 12744
rect 11428 12724 11480 12744
rect 11480 12724 11482 12744
rect 11426 12688 11482 12724
rect 11150 9016 11206 9072
rect 11518 8064 11574 8120
rect 11518 6432 11574 6488
rect 11518 4936 11574 4992
rect 11702 7928 11758 7984
rect 11978 7384 12034 7440
rect 11702 2896 11758 2952
rect 11886 6024 11942 6080
rect 12162 5072 12218 5128
rect 12162 3576 12218 3632
rect 11794 1536 11850 1592
rect 12438 6976 12494 7032
rect 12530 6296 12586 6352
rect 12714 6160 12770 6216
rect 15404 13082 15460 13084
rect 15484 13082 15540 13084
rect 15564 13082 15620 13084
rect 15644 13082 15700 13084
rect 15404 13030 15450 13082
rect 15450 13030 15460 13082
rect 15484 13030 15514 13082
rect 15514 13030 15526 13082
rect 15526 13030 15540 13082
rect 15564 13030 15578 13082
rect 15578 13030 15590 13082
rect 15590 13030 15620 13082
rect 15644 13030 15654 13082
rect 15654 13030 15700 13082
rect 15404 13028 15460 13030
rect 15484 13028 15540 13030
rect 15564 13028 15620 13030
rect 15644 13028 15700 13030
rect 14186 12688 14242 12744
rect 14186 12044 14188 12064
rect 14188 12044 14240 12064
rect 14240 12044 14242 12064
rect 14186 12008 14242 12044
rect 13174 9968 13230 10024
rect 13174 3984 13230 4040
rect 13450 9968 13506 10024
rect 13450 9560 13506 9616
rect 13542 7928 13598 7984
rect 13542 7248 13598 7304
rect 13818 5072 13874 5128
rect 13726 3304 13782 3360
rect 13634 2760 13690 2816
rect 14186 9560 14242 9616
rect 14186 9288 14242 9344
rect 14094 6740 14096 6760
rect 14096 6740 14148 6760
rect 14148 6740 14150 6760
rect 14094 6704 14150 6740
rect 14186 4800 14242 4856
rect 14370 7248 14426 7304
rect 14370 4664 14426 4720
rect 14370 3984 14426 4040
rect 14462 3440 14518 3496
rect 14646 8336 14702 8392
rect 14922 5480 14978 5536
rect 14830 4820 14886 4856
rect 14830 4800 14832 4820
rect 14832 4800 14884 4820
rect 14884 4800 14886 4820
rect 14830 4156 14832 4176
rect 14832 4156 14884 4176
rect 14884 4156 14886 4176
rect 14830 4120 14886 4156
rect 14922 3984 14978 4040
rect 14830 3576 14886 3632
rect 14830 3168 14886 3224
rect 15404 11994 15460 11996
rect 15484 11994 15540 11996
rect 15564 11994 15620 11996
rect 15644 11994 15700 11996
rect 15404 11942 15450 11994
rect 15450 11942 15460 11994
rect 15484 11942 15514 11994
rect 15514 11942 15526 11994
rect 15526 11942 15540 11994
rect 15564 11942 15578 11994
rect 15578 11942 15590 11994
rect 15590 11942 15620 11994
rect 15644 11942 15654 11994
rect 15654 11942 15700 11994
rect 15404 11940 15460 11942
rect 15484 11940 15540 11942
rect 15564 11940 15620 11942
rect 15644 11940 15700 11942
rect 15106 11056 15162 11112
rect 15658 11056 15714 11112
rect 15404 10906 15460 10908
rect 15484 10906 15540 10908
rect 15564 10906 15620 10908
rect 15644 10906 15700 10908
rect 15404 10854 15450 10906
rect 15450 10854 15460 10906
rect 15484 10854 15514 10906
rect 15514 10854 15526 10906
rect 15526 10854 15540 10906
rect 15564 10854 15578 10906
rect 15578 10854 15590 10906
rect 15590 10854 15620 10906
rect 15644 10854 15654 10906
rect 15654 10854 15700 10906
rect 15404 10852 15460 10854
rect 15484 10852 15540 10854
rect 15564 10852 15620 10854
rect 15644 10852 15700 10854
rect 15106 7792 15162 7848
rect 15106 7520 15162 7576
rect 15198 7248 15254 7304
rect 15106 6704 15162 6760
rect 15106 3168 15162 3224
rect 15474 9968 15530 10024
rect 15404 9818 15460 9820
rect 15484 9818 15540 9820
rect 15564 9818 15620 9820
rect 15644 9818 15700 9820
rect 15404 9766 15450 9818
rect 15450 9766 15460 9818
rect 15484 9766 15514 9818
rect 15514 9766 15526 9818
rect 15526 9766 15540 9818
rect 15564 9766 15578 9818
rect 15578 9766 15590 9818
rect 15590 9766 15620 9818
rect 15644 9766 15654 9818
rect 15654 9766 15700 9818
rect 15404 9764 15460 9766
rect 15484 9764 15540 9766
rect 15564 9764 15620 9766
rect 15644 9764 15700 9766
rect 15382 9560 15438 9616
rect 15404 8730 15460 8732
rect 15484 8730 15540 8732
rect 15564 8730 15620 8732
rect 15644 8730 15700 8732
rect 15404 8678 15450 8730
rect 15450 8678 15460 8730
rect 15484 8678 15514 8730
rect 15514 8678 15526 8730
rect 15526 8678 15540 8730
rect 15564 8678 15578 8730
rect 15578 8678 15590 8730
rect 15590 8678 15620 8730
rect 15644 8678 15654 8730
rect 15654 8678 15700 8730
rect 15404 8676 15460 8678
rect 15484 8676 15540 8678
rect 15564 8676 15620 8678
rect 15644 8676 15700 8678
rect 15404 7642 15460 7644
rect 15484 7642 15540 7644
rect 15564 7642 15620 7644
rect 15644 7642 15700 7644
rect 15404 7590 15450 7642
rect 15450 7590 15460 7642
rect 15484 7590 15514 7642
rect 15514 7590 15526 7642
rect 15526 7590 15540 7642
rect 15564 7590 15578 7642
rect 15578 7590 15590 7642
rect 15590 7590 15620 7642
rect 15644 7590 15654 7642
rect 15654 7590 15700 7642
rect 15404 7588 15460 7590
rect 15484 7588 15540 7590
rect 15564 7588 15620 7590
rect 15644 7588 15700 7590
rect 15404 6554 15460 6556
rect 15484 6554 15540 6556
rect 15564 6554 15620 6556
rect 15644 6554 15700 6556
rect 15404 6502 15450 6554
rect 15450 6502 15460 6554
rect 15484 6502 15514 6554
rect 15514 6502 15526 6554
rect 15526 6502 15540 6554
rect 15564 6502 15578 6554
rect 15578 6502 15590 6554
rect 15590 6502 15620 6554
rect 15644 6502 15654 6554
rect 15654 6502 15700 6554
rect 15404 6500 15460 6502
rect 15484 6500 15540 6502
rect 15564 6500 15620 6502
rect 15644 6500 15700 6502
rect 15404 5466 15460 5468
rect 15484 5466 15540 5468
rect 15564 5466 15620 5468
rect 15644 5466 15700 5468
rect 15404 5414 15450 5466
rect 15450 5414 15460 5466
rect 15484 5414 15514 5466
rect 15514 5414 15526 5466
rect 15526 5414 15540 5466
rect 15564 5414 15578 5466
rect 15578 5414 15590 5466
rect 15590 5414 15620 5466
rect 15644 5414 15654 5466
rect 15654 5414 15700 5466
rect 15404 5412 15460 5414
rect 15484 5412 15540 5414
rect 15564 5412 15620 5414
rect 15644 5412 15700 5414
rect 15404 4378 15460 4380
rect 15484 4378 15540 4380
rect 15564 4378 15620 4380
rect 15644 4378 15700 4380
rect 15404 4326 15450 4378
rect 15450 4326 15460 4378
rect 15484 4326 15514 4378
rect 15514 4326 15526 4378
rect 15526 4326 15540 4378
rect 15564 4326 15578 4378
rect 15578 4326 15590 4378
rect 15590 4326 15620 4378
rect 15644 4326 15654 4378
rect 15654 4326 15700 4378
rect 15404 4324 15460 4326
rect 15484 4324 15540 4326
rect 15564 4324 15620 4326
rect 15644 4324 15700 4326
rect 15382 3732 15438 3768
rect 15382 3712 15384 3732
rect 15384 3712 15436 3732
rect 15436 3712 15438 3732
rect 17774 13132 17776 13152
rect 17776 13132 17828 13152
rect 17828 13132 17830 13152
rect 17774 13096 17830 13132
rect 16118 12416 16174 12472
rect 15404 3290 15460 3292
rect 15484 3290 15540 3292
rect 15564 3290 15620 3292
rect 15644 3290 15700 3292
rect 15404 3238 15450 3290
rect 15450 3238 15460 3290
rect 15484 3238 15514 3290
rect 15514 3238 15526 3290
rect 15526 3238 15540 3290
rect 15564 3238 15578 3290
rect 15578 3238 15590 3290
rect 15590 3238 15620 3290
rect 15644 3238 15654 3290
rect 15654 3238 15700 3290
rect 15404 3236 15460 3238
rect 15484 3236 15540 3238
rect 15564 3236 15620 3238
rect 15644 3236 15700 3238
rect 15658 2760 15714 2816
rect 15404 2202 15460 2204
rect 15484 2202 15540 2204
rect 15564 2202 15620 2204
rect 15644 2202 15700 2204
rect 15404 2150 15450 2202
rect 15450 2150 15460 2202
rect 15484 2150 15514 2202
rect 15514 2150 15526 2202
rect 15526 2150 15540 2202
rect 15564 2150 15578 2202
rect 15578 2150 15590 2202
rect 15590 2150 15620 2202
rect 15644 2150 15654 2202
rect 15654 2150 15700 2202
rect 15404 2148 15460 2150
rect 15484 2148 15540 2150
rect 15564 2148 15620 2150
rect 15644 2148 15700 2150
rect 15198 1672 15254 1728
rect 15934 2916 15990 2952
rect 15934 2896 15936 2916
rect 15936 2896 15988 2916
rect 15988 2896 15990 2916
rect 16394 6568 16450 6624
rect 16302 3304 16358 3360
rect 16762 4256 16818 4312
rect 17314 6976 17370 7032
rect 17130 5480 17186 5536
rect 16946 4936 17002 4992
rect 16762 3712 16818 3768
rect 17866 9560 17922 9616
rect 17590 9152 17646 9208
rect 17866 9152 17922 9208
rect 17866 8880 17922 8936
rect 17774 8472 17830 8528
rect 17498 5908 17554 5944
rect 17498 5888 17500 5908
rect 17500 5888 17552 5908
rect 17552 5888 17554 5908
rect 17222 3440 17278 3496
rect 16854 2488 16910 2544
rect 17222 2488 17278 2544
rect 17590 4664 17646 4720
rect 17866 6024 17922 6080
rect 17958 4800 18014 4856
rect 17958 3304 18014 3360
rect 18234 12588 18236 12608
rect 18236 12588 18288 12608
rect 18288 12588 18290 12608
rect 18234 12552 18290 12588
rect 18602 12044 18604 12064
rect 18604 12044 18656 12064
rect 18656 12044 18658 12064
rect 18602 12008 18658 12044
rect 18234 8372 18236 8392
rect 18236 8372 18288 8392
rect 18288 8372 18290 8392
rect 18234 8336 18290 8372
rect 18326 6704 18382 6760
rect 18326 6568 18382 6624
rect 18142 4392 18198 4448
rect 18142 4156 18144 4176
rect 18144 4156 18196 4176
rect 18196 4156 18198 4176
rect 18142 4120 18198 4156
rect 17682 2624 17738 2680
rect 18326 3576 18382 3632
rect 18970 9288 19026 9344
rect 19246 7420 19248 7440
rect 19248 7420 19300 7440
rect 19300 7420 19302 7440
rect 19246 7384 19302 7420
rect 18694 6160 18750 6216
rect 18694 5072 18750 5128
rect 18694 4800 18750 4856
rect 19154 5072 19210 5128
rect 19062 4120 19118 4176
rect 18786 1808 18842 1864
rect 19154 3984 19210 4040
rect 19522 8744 19578 8800
rect 19430 6840 19486 6896
rect 22628 13626 22684 13628
rect 22708 13626 22764 13628
rect 22788 13626 22844 13628
rect 22868 13626 22924 13628
rect 22628 13574 22674 13626
rect 22674 13574 22684 13626
rect 22708 13574 22738 13626
rect 22738 13574 22750 13626
rect 22750 13574 22764 13626
rect 22788 13574 22802 13626
rect 22802 13574 22814 13626
rect 22814 13574 22844 13626
rect 22868 13574 22878 13626
rect 22878 13574 22924 13626
rect 22628 13572 22684 13574
rect 22708 13572 22764 13574
rect 22788 13572 22844 13574
rect 22868 13572 22924 13574
rect 20258 8608 20314 8664
rect 20166 7656 20222 7712
rect 19338 5344 19394 5400
rect 19338 4972 19340 4992
rect 19340 4972 19392 4992
rect 19392 4972 19394 4992
rect 19338 4936 19394 4972
rect 19246 3168 19302 3224
rect 19062 2896 19118 2952
rect 19614 2896 19670 2952
rect 19798 2488 19854 2544
rect 22628 12538 22684 12540
rect 22708 12538 22764 12540
rect 22788 12538 22844 12540
rect 22868 12538 22924 12540
rect 22628 12486 22674 12538
rect 22674 12486 22684 12538
rect 22708 12486 22738 12538
rect 22738 12486 22750 12538
rect 22750 12486 22764 12538
rect 22788 12486 22802 12538
rect 22802 12486 22814 12538
rect 22814 12486 22844 12538
rect 22868 12486 22878 12538
rect 22878 12486 22924 12538
rect 22628 12484 22684 12486
rect 22708 12484 22764 12486
rect 22788 12484 22844 12486
rect 22868 12484 22924 12486
rect 23478 12416 23534 12472
rect 22282 12044 22284 12064
rect 22284 12044 22336 12064
rect 22336 12044 22338 12064
rect 22282 12008 22338 12044
rect 22098 11500 22100 11520
rect 22100 11500 22152 11520
rect 22152 11500 22154 11520
rect 21086 8880 21142 8936
rect 21270 8336 21326 8392
rect 21454 7928 21510 7984
rect 21546 6704 21602 6760
rect 21270 4256 21326 4312
rect 22098 11464 22154 11500
rect 22628 11450 22684 11452
rect 22708 11450 22764 11452
rect 22788 11450 22844 11452
rect 22868 11450 22924 11452
rect 22628 11398 22674 11450
rect 22674 11398 22684 11450
rect 22708 11398 22738 11450
rect 22738 11398 22750 11450
rect 22750 11398 22764 11450
rect 22788 11398 22802 11450
rect 22802 11398 22814 11450
rect 22814 11398 22844 11450
rect 22868 11398 22878 11450
rect 22878 11398 22924 11450
rect 22628 11396 22684 11398
rect 22708 11396 22764 11398
rect 22788 11396 22844 11398
rect 22868 11396 22924 11398
rect 22098 8508 22100 8528
rect 22100 8508 22152 8528
rect 22152 8508 22154 8528
rect 22098 8472 22154 8508
rect 22628 10362 22684 10364
rect 22708 10362 22764 10364
rect 22788 10362 22844 10364
rect 22868 10362 22924 10364
rect 22628 10310 22674 10362
rect 22674 10310 22684 10362
rect 22708 10310 22738 10362
rect 22738 10310 22750 10362
rect 22750 10310 22764 10362
rect 22788 10310 22802 10362
rect 22802 10310 22814 10362
rect 22814 10310 22844 10362
rect 22868 10310 22878 10362
rect 22878 10310 22924 10362
rect 22628 10308 22684 10310
rect 22708 10308 22764 10310
rect 22788 10308 22844 10310
rect 22868 10308 22924 10310
rect 22628 9274 22684 9276
rect 22708 9274 22764 9276
rect 22788 9274 22844 9276
rect 22868 9274 22924 9276
rect 22628 9222 22674 9274
rect 22674 9222 22684 9274
rect 22708 9222 22738 9274
rect 22738 9222 22750 9274
rect 22750 9222 22764 9274
rect 22788 9222 22802 9274
rect 22802 9222 22814 9274
rect 22814 9222 22844 9274
rect 22868 9222 22878 9274
rect 22878 9222 22924 9274
rect 22628 9220 22684 9222
rect 22708 9220 22764 9222
rect 22788 9220 22844 9222
rect 22868 9220 22924 9222
rect 22282 8200 22338 8256
rect 22628 8186 22684 8188
rect 22708 8186 22764 8188
rect 22788 8186 22844 8188
rect 22868 8186 22924 8188
rect 22628 8134 22674 8186
rect 22674 8134 22684 8186
rect 22708 8134 22738 8186
rect 22738 8134 22750 8186
rect 22750 8134 22764 8186
rect 22788 8134 22802 8186
rect 22802 8134 22814 8186
rect 22814 8134 22844 8186
rect 22868 8134 22878 8186
rect 22878 8134 22924 8186
rect 22628 8132 22684 8134
rect 22708 8132 22764 8134
rect 22788 8132 22844 8134
rect 22868 8132 22924 8134
rect 22006 7520 22062 7576
rect 22190 6840 22246 6896
rect 21730 4800 21786 4856
rect 22628 7098 22684 7100
rect 22708 7098 22764 7100
rect 22788 7098 22844 7100
rect 22868 7098 22924 7100
rect 22628 7046 22674 7098
rect 22674 7046 22684 7098
rect 22708 7046 22738 7098
rect 22738 7046 22750 7098
rect 22750 7046 22764 7098
rect 22788 7046 22802 7098
rect 22802 7046 22814 7098
rect 22814 7046 22844 7098
rect 22868 7046 22878 7098
rect 22878 7046 22924 7098
rect 22628 7044 22684 7046
rect 22708 7044 22764 7046
rect 22788 7044 22844 7046
rect 22868 7044 22924 7046
rect 22628 6010 22684 6012
rect 22708 6010 22764 6012
rect 22788 6010 22844 6012
rect 22868 6010 22924 6012
rect 22628 5958 22674 6010
rect 22674 5958 22684 6010
rect 22708 5958 22738 6010
rect 22738 5958 22750 6010
rect 22750 5958 22764 6010
rect 22788 5958 22802 6010
rect 22802 5958 22814 6010
rect 22814 5958 22844 6010
rect 22868 5958 22878 6010
rect 22878 5958 22924 6010
rect 22628 5956 22684 5958
rect 22708 5956 22764 5958
rect 22788 5956 22844 5958
rect 22868 5956 22924 5958
rect 22628 4922 22684 4924
rect 22708 4922 22764 4924
rect 22788 4922 22844 4924
rect 22868 4922 22924 4924
rect 22628 4870 22674 4922
rect 22674 4870 22684 4922
rect 22708 4870 22738 4922
rect 22738 4870 22750 4922
rect 22750 4870 22764 4922
rect 22788 4870 22802 4922
rect 22802 4870 22814 4922
rect 22814 4870 22844 4922
rect 22868 4870 22878 4922
rect 22878 4870 22924 4922
rect 22628 4868 22684 4870
rect 22708 4868 22764 4870
rect 22788 4868 22844 4870
rect 22868 4868 22924 4870
rect 22558 4664 22614 4720
rect 23478 7384 23534 7440
rect 23202 6840 23258 6896
rect 23754 7812 23810 7848
rect 23754 7792 23756 7812
rect 23756 7792 23808 7812
rect 23808 7792 23810 7812
rect 23938 11056 23994 11112
rect 37076 13626 37132 13628
rect 37156 13626 37212 13628
rect 37236 13626 37292 13628
rect 37316 13626 37372 13628
rect 37076 13574 37122 13626
rect 37122 13574 37132 13626
rect 37156 13574 37186 13626
rect 37186 13574 37198 13626
rect 37198 13574 37212 13626
rect 37236 13574 37250 13626
rect 37250 13574 37262 13626
rect 37262 13574 37292 13626
rect 37316 13574 37326 13626
rect 37326 13574 37372 13626
rect 37076 13572 37132 13574
rect 37156 13572 37212 13574
rect 37236 13572 37292 13574
rect 37316 13572 37372 13574
rect 51524 13626 51580 13628
rect 51604 13626 51660 13628
rect 51684 13626 51740 13628
rect 51764 13626 51820 13628
rect 51524 13574 51570 13626
rect 51570 13574 51580 13626
rect 51604 13574 51634 13626
rect 51634 13574 51646 13626
rect 51646 13574 51660 13626
rect 51684 13574 51698 13626
rect 51698 13574 51710 13626
rect 51710 13574 51740 13626
rect 51764 13574 51774 13626
rect 51774 13574 51820 13626
rect 51524 13572 51580 13574
rect 51604 13572 51660 13574
rect 51684 13572 51740 13574
rect 51764 13572 51820 13574
rect 29852 13082 29908 13084
rect 29932 13082 29988 13084
rect 30012 13082 30068 13084
rect 30092 13082 30148 13084
rect 29852 13030 29898 13082
rect 29898 13030 29908 13082
rect 29932 13030 29962 13082
rect 29962 13030 29974 13082
rect 29974 13030 29988 13082
rect 30012 13030 30026 13082
rect 30026 13030 30038 13082
rect 30038 13030 30068 13082
rect 30092 13030 30102 13082
rect 30102 13030 30148 13082
rect 29852 13028 29908 13030
rect 29932 13028 29988 13030
rect 30012 13028 30068 13030
rect 30092 13028 30148 13030
rect 44300 13082 44356 13084
rect 44380 13082 44436 13084
rect 44460 13082 44516 13084
rect 44540 13082 44596 13084
rect 44300 13030 44346 13082
rect 44346 13030 44356 13082
rect 44380 13030 44410 13082
rect 44410 13030 44422 13082
rect 44422 13030 44436 13082
rect 44460 13030 44474 13082
rect 44474 13030 44486 13082
rect 44486 13030 44516 13082
rect 44540 13030 44550 13082
rect 44550 13030 44596 13082
rect 44300 13028 44356 13030
rect 44380 13028 44436 13030
rect 44460 13028 44516 13030
rect 44540 13028 44596 13030
rect 37076 12538 37132 12540
rect 37156 12538 37212 12540
rect 37236 12538 37292 12540
rect 37316 12538 37372 12540
rect 37076 12486 37122 12538
rect 37122 12486 37132 12538
rect 37156 12486 37186 12538
rect 37186 12486 37198 12538
rect 37198 12486 37212 12538
rect 37236 12486 37250 12538
rect 37250 12486 37262 12538
rect 37262 12486 37292 12538
rect 37316 12486 37326 12538
rect 37326 12486 37372 12538
rect 37076 12484 37132 12486
rect 37156 12484 37212 12486
rect 37236 12484 37292 12486
rect 37316 12484 37372 12486
rect 51524 12538 51580 12540
rect 51604 12538 51660 12540
rect 51684 12538 51740 12540
rect 51764 12538 51820 12540
rect 51524 12486 51570 12538
rect 51570 12486 51580 12538
rect 51604 12486 51634 12538
rect 51634 12486 51646 12538
rect 51646 12486 51660 12538
rect 51684 12486 51698 12538
rect 51698 12486 51710 12538
rect 51710 12486 51740 12538
rect 51764 12486 51774 12538
rect 51774 12486 51820 12538
rect 51524 12484 51580 12486
rect 51604 12484 51660 12486
rect 51684 12484 51740 12486
rect 51764 12484 51820 12486
rect 24214 9424 24270 9480
rect 24398 8608 24454 8664
rect 24214 8492 24270 8528
rect 24214 8472 24216 8492
rect 24216 8472 24268 8492
rect 24268 8472 24270 8492
rect 24122 7384 24178 7440
rect 23202 5616 23258 5672
rect 23018 4120 23074 4176
rect 23018 3848 23074 3904
rect 22628 3834 22684 3836
rect 22708 3834 22764 3836
rect 22788 3834 22844 3836
rect 22868 3834 22924 3836
rect 22628 3782 22674 3834
rect 22674 3782 22684 3834
rect 22708 3782 22738 3834
rect 22738 3782 22750 3834
rect 22750 3782 22764 3834
rect 22788 3782 22802 3834
rect 22802 3782 22814 3834
rect 22814 3782 22844 3834
rect 22868 3782 22878 3834
rect 22878 3782 22924 3834
rect 22628 3780 22684 3782
rect 22708 3780 22764 3782
rect 22788 3780 22844 3782
rect 22868 3780 22924 3782
rect 22006 2216 22062 2272
rect 23386 3576 23442 3632
rect 22628 2746 22684 2748
rect 22708 2746 22764 2748
rect 22788 2746 22844 2748
rect 22868 2746 22924 2748
rect 22628 2694 22674 2746
rect 22674 2694 22684 2746
rect 22708 2694 22738 2746
rect 22738 2694 22750 2746
rect 22750 2694 22764 2746
rect 22788 2694 22802 2746
rect 22802 2694 22814 2746
rect 22814 2694 22844 2746
rect 22868 2694 22878 2746
rect 22878 2694 22924 2746
rect 22628 2692 22684 2694
rect 22708 2692 22764 2694
rect 22788 2692 22844 2694
rect 22868 2692 22924 2694
rect 22834 1400 22890 1456
rect 23018 2080 23074 2136
rect 23202 1944 23258 2000
rect 23754 5480 23810 5536
rect 23478 3168 23534 3224
rect 23386 1128 23442 1184
rect 24214 6160 24270 6216
rect 24398 6024 24454 6080
rect 23938 4392 23994 4448
rect 24214 4392 24270 4448
rect 24582 8336 24638 8392
rect 25042 7284 25044 7304
rect 25044 7284 25096 7304
rect 25096 7284 25098 7304
rect 25042 7248 25098 7284
rect 24674 6704 24730 6760
rect 24766 6196 24768 6216
rect 24768 6196 24820 6216
rect 24820 6196 24822 6216
rect 24766 6160 24822 6196
rect 24490 4820 24546 4856
rect 24490 4800 24492 4820
rect 24492 4800 24544 4820
rect 24544 4800 24546 4820
rect 24766 5208 24822 5264
rect 24582 3848 24638 3904
rect 25134 6568 25190 6624
rect 25226 4120 25282 4176
rect 25410 6704 25466 6760
rect 25502 6160 25558 6216
rect 25870 7792 25926 7848
rect 25594 5072 25650 5128
rect 25686 4664 25742 4720
rect 25778 4392 25834 4448
rect 26422 7248 26478 7304
rect 25870 1672 25926 1728
rect 26790 9016 26846 9072
rect 27158 8900 27214 8936
rect 27158 8880 27160 8900
rect 27160 8880 27212 8900
rect 27212 8880 27214 8900
rect 27342 8200 27398 8256
rect 27342 7928 27398 7984
rect 26698 7656 26754 7712
rect 26790 7384 26846 7440
rect 27434 6976 27490 7032
rect 27434 6180 27490 6216
rect 27434 6160 27436 6180
rect 27436 6160 27488 6180
rect 27488 6160 27490 6180
rect 26974 5344 27030 5400
rect 29852 11994 29908 11996
rect 29932 11994 29988 11996
rect 30012 11994 30068 11996
rect 30092 11994 30148 11996
rect 29852 11942 29898 11994
rect 29898 11942 29908 11994
rect 29932 11942 29962 11994
rect 29962 11942 29974 11994
rect 29974 11942 29988 11994
rect 30012 11942 30026 11994
rect 30026 11942 30038 11994
rect 30038 11942 30068 11994
rect 30092 11942 30102 11994
rect 30102 11942 30148 11994
rect 29852 11940 29908 11942
rect 29932 11940 29988 11942
rect 30012 11940 30068 11942
rect 30092 11940 30148 11942
rect 35714 11056 35770 11112
rect 28446 9580 28502 9616
rect 28446 9560 28448 9580
rect 28448 9560 28500 9580
rect 28500 9560 28502 9580
rect 28998 9016 29054 9072
rect 27986 8744 28042 8800
rect 27894 7828 27896 7848
rect 27896 7828 27948 7848
rect 27948 7828 27950 7848
rect 27894 7792 27950 7828
rect 28998 7248 29054 7304
rect 28998 5888 29054 5944
rect 26882 5208 26938 5264
rect 26514 4256 26570 4312
rect 26422 1808 26478 1864
rect 26974 2388 26976 2408
rect 26976 2388 27028 2408
rect 27028 2388 27030 2408
rect 26974 2352 27030 2388
rect 27802 3304 27858 3360
rect 28906 5092 28962 5128
rect 28906 5072 28908 5092
rect 28908 5072 28960 5092
rect 28960 5072 28962 5092
rect 27986 2216 28042 2272
rect 29852 10906 29908 10908
rect 29932 10906 29988 10908
rect 30012 10906 30068 10908
rect 30092 10906 30148 10908
rect 29852 10854 29898 10906
rect 29898 10854 29908 10906
rect 29932 10854 29962 10906
rect 29962 10854 29974 10906
rect 29974 10854 29988 10906
rect 30012 10854 30026 10906
rect 30026 10854 30038 10906
rect 30038 10854 30068 10906
rect 30092 10854 30102 10906
rect 30102 10854 30148 10906
rect 29852 10852 29908 10854
rect 29932 10852 29988 10854
rect 30012 10852 30068 10854
rect 30092 10852 30148 10854
rect 29852 9818 29908 9820
rect 29932 9818 29988 9820
rect 30012 9818 30068 9820
rect 30092 9818 30148 9820
rect 29852 9766 29898 9818
rect 29898 9766 29908 9818
rect 29932 9766 29962 9818
rect 29962 9766 29974 9818
rect 29974 9766 29988 9818
rect 30012 9766 30026 9818
rect 30026 9766 30038 9818
rect 30038 9766 30068 9818
rect 30092 9766 30102 9818
rect 30102 9766 30148 9818
rect 29852 9764 29908 9766
rect 29932 9764 29988 9766
rect 30012 9764 30068 9766
rect 30092 9764 30148 9766
rect 29458 8472 29514 8528
rect 29852 8730 29908 8732
rect 29932 8730 29988 8732
rect 30012 8730 30068 8732
rect 30092 8730 30148 8732
rect 29852 8678 29898 8730
rect 29898 8678 29908 8730
rect 29932 8678 29962 8730
rect 29962 8678 29974 8730
rect 29974 8678 29988 8730
rect 30012 8678 30026 8730
rect 30026 8678 30038 8730
rect 30038 8678 30068 8730
rect 30092 8678 30102 8730
rect 30102 8678 30148 8730
rect 29852 8676 29908 8678
rect 29932 8676 29988 8678
rect 30012 8676 30068 8678
rect 30092 8676 30148 8678
rect 29642 7520 29698 7576
rect 29852 7642 29908 7644
rect 29932 7642 29988 7644
rect 30012 7642 30068 7644
rect 30092 7642 30148 7644
rect 29852 7590 29898 7642
rect 29898 7590 29908 7642
rect 29932 7590 29962 7642
rect 29962 7590 29974 7642
rect 29974 7590 29988 7642
rect 30012 7590 30026 7642
rect 30026 7590 30038 7642
rect 30038 7590 30068 7642
rect 30092 7590 30102 7642
rect 30102 7590 30148 7642
rect 29852 7588 29908 7590
rect 29932 7588 29988 7590
rect 30012 7588 30068 7590
rect 30092 7588 30148 7590
rect 29734 6996 29790 7032
rect 29734 6976 29736 6996
rect 29736 6976 29788 6996
rect 29788 6976 29790 6996
rect 29852 6554 29908 6556
rect 29932 6554 29988 6556
rect 30012 6554 30068 6556
rect 30092 6554 30148 6556
rect 29852 6502 29898 6554
rect 29898 6502 29908 6554
rect 29932 6502 29962 6554
rect 29962 6502 29974 6554
rect 29974 6502 29988 6554
rect 30012 6502 30026 6554
rect 30026 6502 30038 6554
rect 30038 6502 30068 6554
rect 30092 6502 30102 6554
rect 30102 6502 30148 6554
rect 29852 6500 29908 6502
rect 29932 6500 29988 6502
rect 30012 6500 30068 6502
rect 30092 6500 30148 6502
rect 29734 5788 29736 5808
rect 29736 5788 29788 5808
rect 29788 5788 29790 5808
rect 29734 5752 29790 5788
rect 29852 5466 29908 5468
rect 29932 5466 29988 5468
rect 30012 5466 30068 5468
rect 30092 5466 30148 5468
rect 29852 5414 29898 5466
rect 29898 5414 29908 5466
rect 29932 5414 29962 5466
rect 29962 5414 29974 5466
rect 29974 5414 29988 5466
rect 30012 5414 30026 5466
rect 30026 5414 30038 5466
rect 30038 5414 30068 5466
rect 30092 5414 30102 5466
rect 30102 5414 30148 5466
rect 29852 5412 29908 5414
rect 29932 5412 29988 5414
rect 30012 5412 30068 5414
rect 30092 5412 30148 5414
rect 29182 4120 29238 4176
rect 29366 1808 29422 1864
rect 29642 4936 29698 4992
rect 31022 8492 31078 8528
rect 31022 8472 31024 8492
rect 31024 8472 31076 8492
rect 31076 8472 31078 8492
rect 30378 7520 30434 7576
rect 30378 6840 30434 6896
rect 30378 5652 30380 5672
rect 30380 5652 30432 5672
rect 30432 5652 30434 5672
rect 30378 5616 30434 5652
rect 29852 4378 29908 4380
rect 29932 4378 29988 4380
rect 30012 4378 30068 4380
rect 30092 4378 30148 4380
rect 29852 4326 29898 4378
rect 29898 4326 29908 4378
rect 29932 4326 29962 4378
rect 29962 4326 29974 4378
rect 29974 4326 29988 4378
rect 30012 4326 30026 4378
rect 30026 4326 30038 4378
rect 30038 4326 30068 4378
rect 30092 4326 30102 4378
rect 30102 4326 30148 4378
rect 29852 4324 29908 4326
rect 29932 4324 29988 4326
rect 30012 4324 30068 4326
rect 30092 4324 30148 4326
rect 30102 4140 30158 4176
rect 30102 4120 30104 4140
rect 30104 4120 30156 4140
rect 30156 4120 30158 4140
rect 29852 3290 29908 3292
rect 29932 3290 29988 3292
rect 30012 3290 30068 3292
rect 30092 3290 30148 3292
rect 29852 3238 29898 3290
rect 29898 3238 29908 3290
rect 29932 3238 29962 3290
rect 29962 3238 29974 3290
rect 29974 3238 29988 3290
rect 30012 3238 30026 3290
rect 30026 3238 30038 3290
rect 30038 3238 30068 3290
rect 30092 3238 30102 3290
rect 30102 3238 30148 3290
rect 29852 3236 29908 3238
rect 29932 3236 29988 3238
rect 30012 3236 30068 3238
rect 30092 3236 30148 3238
rect 30838 6976 30894 7032
rect 30838 6840 30894 6896
rect 31022 4800 31078 4856
rect 30562 3848 30618 3904
rect 31482 8472 31538 8528
rect 31206 3304 31262 3360
rect 29852 2202 29908 2204
rect 29932 2202 29988 2204
rect 30012 2202 30068 2204
rect 30092 2202 30148 2204
rect 29852 2150 29898 2202
rect 29898 2150 29908 2202
rect 29932 2150 29962 2202
rect 29962 2150 29974 2202
rect 29974 2150 29988 2202
rect 30012 2150 30026 2202
rect 30026 2150 30038 2202
rect 30038 2150 30068 2202
rect 30092 2150 30102 2202
rect 30102 2150 30148 2202
rect 29852 2148 29908 2150
rect 29932 2148 29988 2150
rect 30012 2148 30068 2150
rect 30092 2148 30148 2150
rect 30838 2760 30894 2816
rect 30746 1536 30802 1592
rect 32218 8236 32220 8256
rect 32220 8236 32272 8256
rect 32272 8236 32274 8256
rect 32218 8200 32274 8236
rect 31850 7248 31906 7304
rect 32034 6976 32090 7032
rect 31850 6432 31906 6488
rect 32310 6332 32312 6352
rect 32312 6332 32364 6352
rect 32364 6332 32366 6352
rect 32310 6296 32366 6332
rect 33598 8372 33600 8392
rect 33600 8372 33652 8392
rect 33652 8372 33654 8392
rect 33598 8336 33654 8372
rect 32586 6024 32642 6080
rect 31942 5344 31998 5400
rect 31574 4664 31630 4720
rect 31482 3032 31538 3088
rect 33782 6296 33838 6352
rect 33690 5888 33746 5944
rect 35530 9172 35586 9208
rect 35530 9152 35532 9172
rect 35532 9152 35584 9172
rect 35584 9152 35586 9172
rect 34150 5208 34206 5264
rect 34518 4936 34574 4992
rect 34150 4120 34206 4176
rect 35806 6860 35862 6896
rect 35806 6840 35808 6860
rect 35808 6840 35860 6860
rect 35860 6840 35862 6860
rect 44300 11994 44356 11996
rect 44380 11994 44436 11996
rect 44460 11994 44516 11996
rect 44540 11994 44596 11996
rect 44300 11942 44346 11994
rect 44346 11942 44356 11994
rect 44380 11942 44410 11994
rect 44410 11942 44422 11994
rect 44422 11942 44436 11994
rect 44460 11942 44474 11994
rect 44474 11942 44486 11994
rect 44486 11942 44516 11994
rect 44540 11942 44550 11994
rect 44550 11942 44596 11994
rect 44300 11940 44356 11942
rect 44380 11940 44436 11942
rect 44460 11940 44516 11942
rect 44540 11940 44596 11942
rect 37076 11450 37132 11452
rect 37156 11450 37212 11452
rect 37236 11450 37292 11452
rect 37316 11450 37372 11452
rect 37076 11398 37122 11450
rect 37122 11398 37132 11450
rect 37156 11398 37186 11450
rect 37186 11398 37198 11450
rect 37198 11398 37212 11450
rect 37236 11398 37250 11450
rect 37250 11398 37262 11450
rect 37262 11398 37292 11450
rect 37316 11398 37326 11450
rect 37326 11398 37372 11450
rect 37076 11396 37132 11398
rect 37156 11396 37212 11398
rect 37236 11396 37292 11398
rect 37316 11396 37372 11398
rect 37076 10362 37132 10364
rect 37156 10362 37212 10364
rect 37236 10362 37292 10364
rect 37316 10362 37372 10364
rect 37076 10310 37122 10362
rect 37122 10310 37132 10362
rect 37156 10310 37186 10362
rect 37186 10310 37198 10362
rect 37198 10310 37212 10362
rect 37236 10310 37250 10362
rect 37250 10310 37262 10362
rect 37262 10310 37292 10362
rect 37316 10310 37326 10362
rect 37326 10310 37372 10362
rect 37076 10308 37132 10310
rect 37156 10308 37212 10310
rect 37236 10308 37292 10310
rect 37316 10308 37372 10310
rect 37076 9274 37132 9276
rect 37156 9274 37212 9276
rect 37236 9274 37292 9276
rect 37316 9274 37372 9276
rect 37076 9222 37122 9274
rect 37122 9222 37132 9274
rect 37156 9222 37186 9274
rect 37186 9222 37198 9274
rect 37198 9222 37212 9274
rect 37236 9222 37250 9274
rect 37250 9222 37262 9274
rect 37262 9222 37292 9274
rect 37316 9222 37326 9274
rect 37326 9222 37372 9274
rect 37076 9220 37132 9222
rect 37156 9220 37212 9222
rect 37236 9220 37292 9222
rect 37316 9220 37372 9222
rect 37076 8186 37132 8188
rect 37156 8186 37212 8188
rect 37236 8186 37292 8188
rect 37316 8186 37372 8188
rect 37076 8134 37122 8186
rect 37122 8134 37132 8186
rect 37156 8134 37186 8186
rect 37186 8134 37198 8186
rect 37198 8134 37212 8186
rect 37236 8134 37250 8186
rect 37250 8134 37262 8186
rect 37262 8134 37292 8186
rect 37316 8134 37326 8186
rect 37326 8134 37372 8186
rect 37076 8132 37132 8134
rect 37156 8132 37212 8134
rect 37236 8132 37292 8134
rect 37316 8132 37372 8134
rect 37076 7098 37132 7100
rect 37156 7098 37212 7100
rect 37236 7098 37292 7100
rect 37316 7098 37372 7100
rect 37076 7046 37122 7098
rect 37122 7046 37132 7098
rect 37156 7046 37186 7098
rect 37186 7046 37198 7098
rect 37198 7046 37212 7098
rect 37236 7046 37250 7098
rect 37250 7046 37262 7098
rect 37262 7046 37292 7098
rect 37316 7046 37326 7098
rect 37326 7046 37372 7098
rect 37076 7044 37132 7046
rect 37156 7044 37212 7046
rect 37236 7044 37292 7046
rect 37316 7044 37372 7046
rect 37094 6160 37150 6216
rect 37076 6010 37132 6012
rect 37156 6010 37212 6012
rect 37236 6010 37292 6012
rect 37316 6010 37372 6012
rect 37076 5958 37122 6010
rect 37122 5958 37132 6010
rect 37156 5958 37186 6010
rect 37186 5958 37198 6010
rect 37198 5958 37212 6010
rect 37236 5958 37250 6010
rect 37250 5958 37262 6010
rect 37262 5958 37292 6010
rect 37316 5958 37326 6010
rect 37326 5958 37372 6010
rect 37076 5956 37132 5958
rect 37156 5956 37212 5958
rect 37236 5956 37292 5958
rect 37316 5956 37372 5958
rect 36358 5616 36414 5672
rect 34886 3576 34942 3632
rect 34610 2488 34666 2544
rect 35806 4392 35862 4448
rect 35714 3848 35770 3904
rect 35714 2216 35770 2272
rect 38290 6840 38346 6896
rect 38106 6296 38162 6352
rect 37922 6160 37978 6216
rect 37076 4922 37132 4924
rect 37156 4922 37212 4924
rect 37236 4922 37292 4924
rect 37316 4922 37372 4924
rect 37076 4870 37122 4922
rect 37122 4870 37132 4922
rect 37156 4870 37186 4922
rect 37186 4870 37198 4922
rect 37198 4870 37212 4922
rect 37236 4870 37250 4922
rect 37250 4870 37262 4922
rect 37262 4870 37292 4922
rect 37316 4870 37326 4922
rect 37326 4870 37372 4922
rect 37076 4868 37132 4870
rect 37156 4868 37212 4870
rect 37236 4868 37292 4870
rect 37316 4868 37372 4870
rect 36726 3188 36782 3224
rect 36726 3168 36728 3188
rect 36728 3168 36780 3188
rect 36780 3168 36782 3188
rect 36358 1400 36414 1456
rect 39026 4664 39082 4720
rect 38106 4256 38162 4312
rect 37076 3834 37132 3836
rect 37156 3834 37212 3836
rect 37236 3834 37292 3836
rect 37316 3834 37372 3836
rect 37076 3782 37122 3834
rect 37122 3782 37132 3834
rect 37156 3782 37186 3834
rect 37186 3782 37198 3834
rect 37198 3782 37212 3834
rect 37236 3782 37250 3834
rect 37250 3782 37262 3834
rect 37262 3782 37292 3834
rect 37316 3782 37326 3834
rect 37326 3782 37372 3834
rect 37076 3780 37132 3782
rect 37156 3780 37212 3782
rect 37236 3780 37292 3782
rect 37316 3780 37372 3782
rect 37462 3712 37518 3768
rect 37370 3304 37426 3360
rect 37076 2746 37132 2748
rect 37156 2746 37212 2748
rect 37236 2746 37292 2748
rect 37316 2746 37372 2748
rect 37076 2694 37122 2746
rect 37122 2694 37132 2746
rect 37156 2694 37186 2746
rect 37186 2694 37198 2746
rect 37198 2694 37212 2746
rect 37236 2694 37250 2746
rect 37250 2694 37262 2746
rect 37262 2694 37292 2746
rect 37316 2694 37326 2746
rect 37326 2694 37372 2746
rect 37076 2692 37132 2694
rect 37156 2692 37212 2694
rect 37236 2692 37292 2694
rect 37316 2692 37372 2694
rect 37738 3052 37794 3088
rect 37738 3032 37740 3052
rect 37740 3032 37792 3052
rect 37792 3032 37794 3052
rect 37738 2760 37794 2816
rect 39946 7384 40002 7440
rect 40222 5072 40278 5128
rect 41878 7520 41934 7576
rect 42890 7812 42946 7848
rect 42890 7792 42892 7812
rect 42892 7792 42944 7812
rect 42944 7792 42946 7812
rect 40406 5652 40408 5672
rect 40408 5652 40460 5672
rect 40460 5652 40462 5672
rect 40406 5616 40462 5652
rect 42706 6704 42762 6760
rect 42982 5888 43038 5944
rect 42798 5344 42854 5400
rect 40406 4800 40462 4856
rect 39946 4120 40002 4176
rect 39118 3848 39174 3904
rect 38290 3476 38292 3496
rect 38292 3476 38344 3496
rect 38344 3476 38346 3496
rect 38290 3440 38346 3476
rect 38474 2352 38530 2408
rect 39118 3168 39174 3224
rect 39210 2508 39266 2544
rect 39210 2488 39212 2508
rect 39212 2488 39264 2508
rect 39264 2488 39266 2508
rect 38566 1944 38622 2000
rect 38566 1536 38622 1592
rect 39302 1808 39358 1864
rect 41326 4700 41328 4720
rect 41328 4700 41380 4720
rect 41380 4700 41382 4720
rect 41326 4664 41382 4700
rect 43166 5072 43222 5128
rect 42706 4392 42762 4448
rect 40682 3576 40738 3632
rect 42430 3884 42432 3904
rect 42432 3884 42484 3904
rect 42484 3884 42486 3904
rect 42430 3848 42486 3884
rect 41786 3476 41788 3496
rect 41788 3476 41840 3496
rect 41840 3476 41842 3496
rect 41786 3440 41842 3476
rect 41050 3052 41106 3088
rect 41050 3032 41052 3052
rect 41052 3032 41104 3052
rect 41104 3032 41106 3052
rect 40774 2760 40830 2816
rect 40682 2488 40738 2544
rect 41786 2252 41788 2272
rect 41788 2252 41840 2272
rect 41840 2252 41842 2272
rect 41786 2216 41842 2252
rect 44300 10906 44356 10908
rect 44380 10906 44436 10908
rect 44460 10906 44516 10908
rect 44540 10906 44596 10908
rect 44300 10854 44346 10906
rect 44346 10854 44356 10906
rect 44380 10854 44410 10906
rect 44410 10854 44422 10906
rect 44422 10854 44436 10906
rect 44460 10854 44474 10906
rect 44474 10854 44486 10906
rect 44486 10854 44516 10906
rect 44540 10854 44550 10906
rect 44550 10854 44596 10906
rect 44300 10852 44356 10854
rect 44380 10852 44436 10854
rect 44460 10852 44516 10854
rect 44540 10852 44596 10854
rect 44300 9818 44356 9820
rect 44380 9818 44436 9820
rect 44460 9818 44516 9820
rect 44540 9818 44596 9820
rect 44300 9766 44346 9818
rect 44346 9766 44356 9818
rect 44380 9766 44410 9818
rect 44410 9766 44422 9818
rect 44422 9766 44436 9818
rect 44460 9766 44474 9818
rect 44474 9766 44486 9818
rect 44486 9766 44516 9818
rect 44540 9766 44550 9818
rect 44550 9766 44596 9818
rect 44300 9764 44356 9766
rect 44380 9764 44436 9766
rect 44460 9764 44516 9766
rect 44540 9764 44596 9766
rect 51524 11450 51580 11452
rect 51604 11450 51660 11452
rect 51684 11450 51740 11452
rect 51764 11450 51820 11452
rect 51524 11398 51570 11450
rect 51570 11398 51580 11450
rect 51604 11398 51634 11450
rect 51634 11398 51646 11450
rect 51646 11398 51660 11450
rect 51684 11398 51698 11450
rect 51698 11398 51710 11450
rect 51710 11398 51740 11450
rect 51764 11398 51774 11450
rect 51774 11398 51820 11450
rect 51524 11396 51580 11398
rect 51604 11396 51660 11398
rect 51684 11396 51740 11398
rect 51764 11396 51820 11398
rect 44270 9016 44326 9072
rect 44638 8880 44694 8936
rect 44300 8730 44356 8732
rect 44380 8730 44436 8732
rect 44460 8730 44516 8732
rect 44540 8730 44596 8732
rect 44300 8678 44346 8730
rect 44346 8678 44356 8730
rect 44380 8678 44410 8730
rect 44410 8678 44422 8730
rect 44422 8678 44436 8730
rect 44460 8678 44474 8730
rect 44474 8678 44486 8730
rect 44486 8678 44516 8730
rect 44540 8678 44550 8730
rect 44550 8678 44596 8730
rect 44300 8676 44356 8678
rect 44380 8676 44436 8678
rect 44460 8676 44516 8678
rect 44540 8676 44596 8678
rect 44300 7642 44356 7644
rect 44380 7642 44436 7644
rect 44460 7642 44516 7644
rect 44540 7642 44596 7644
rect 44300 7590 44346 7642
rect 44346 7590 44356 7642
rect 44380 7590 44410 7642
rect 44410 7590 44422 7642
rect 44422 7590 44436 7642
rect 44460 7590 44474 7642
rect 44474 7590 44486 7642
rect 44486 7590 44516 7642
rect 44540 7590 44550 7642
rect 44550 7590 44596 7642
rect 44300 7588 44356 7590
rect 44380 7588 44436 7590
rect 44460 7588 44516 7590
rect 44540 7588 44596 7590
rect 43626 4664 43682 4720
rect 43534 3984 43590 4040
rect 42614 3304 42670 3360
rect 42522 1944 42578 2000
rect 42246 1808 42302 1864
rect 42798 2760 42854 2816
rect 42614 1672 42670 1728
rect 44300 6554 44356 6556
rect 44380 6554 44436 6556
rect 44460 6554 44516 6556
rect 44540 6554 44596 6556
rect 44300 6502 44346 6554
rect 44346 6502 44356 6554
rect 44380 6502 44410 6554
rect 44410 6502 44422 6554
rect 44422 6502 44436 6554
rect 44460 6502 44474 6554
rect 44474 6502 44486 6554
rect 44486 6502 44516 6554
rect 44540 6502 44550 6554
rect 44550 6502 44596 6554
rect 44300 6500 44356 6502
rect 44380 6500 44436 6502
rect 44460 6500 44516 6502
rect 44540 6500 44596 6502
rect 51524 10362 51580 10364
rect 51604 10362 51660 10364
rect 51684 10362 51740 10364
rect 51764 10362 51820 10364
rect 51524 10310 51570 10362
rect 51570 10310 51580 10362
rect 51604 10310 51634 10362
rect 51634 10310 51646 10362
rect 51646 10310 51660 10362
rect 51684 10310 51698 10362
rect 51698 10310 51710 10362
rect 51710 10310 51740 10362
rect 51764 10310 51774 10362
rect 51774 10310 51820 10362
rect 51524 10308 51580 10310
rect 51604 10308 51660 10310
rect 51684 10308 51740 10310
rect 51764 10308 51820 10310
rect 48042 8200 48098 8256
rect 49882 8200 49938 8256
rect 51524 9274 51580 9276
rect 51604 9274 51660 9276
rect 51684 9274 51740 9276
rect 51764 9274 51820 9276
rect 51524 9222 51570 9274
rect 51570 9222 51580 9274
rect 51604 9222 51634 9274
rect 51634 9222 51646 9274
rect 51646 9222 51660 9274
rect 51684 9222 51698 9274
rect 51698 9222 51710 9274
rect 51710 9222 51740 9274
rect 51764 9222 51774 9274
rect 51774 9222 51820 9274
rect 51524 9220 51580 9222
rect 51604 9220 51660 9222
rect 51684 9220 51740 9222
rect 51764 9220 51820 9222
rect 51524 8186 51580 8188
rect 51604 8186 51660 8188
rect 51684 8186 51740 8188
rect 51764 8186 51820 8188
rect 51524 8134 51570 8186
rect 51570 8134 51580 8186
rect 51604 8134 51634 8186
rect 51634 8134 51646 8186
rect 51646 8134 51660 8186
rect 51684 8134 51698 8186
rect 51698 8134 51710 8186
rect 51710 8134 51740 8186
rect 51764 8134 51774 8186
rect 51774 8134 51820 8186
rect 51524 8132 51580 8134
rect 51604 8132 51660 8134
rect 51684 8132 51740 8134
rect 51764 8132 51820 8134
rect 48594 6996 48650 7032
rect 48594 6976 48596 6996
rect 48596 6976 48648 6996
rect 48648 6976 48650 6996
rect 47214 6840 47270 6896
rect 45834 6180 45890 6216
rect 45834 6160 45836 6180
rect 45836 6160 45888 6180
rect 45888 6160 45890 6180
rect 44300 5466 44356 5468
rect 44380 5466 44436 5468
rect 44460 5466 44516 5468
rect 44540 5466 44596 5468
rect 44300 5414 44346 5466
rect 44346 5414 44356 5466
rect 44380 5414 44410 5466
rect 44410 5414 44422 5466
rect 44422 5414 44436 5466
rect 44460 5414 44474 5466
rect 44474 5414 44486 5466
rect 44486 5414 44516 5466
rect 44540 5414 44550 5466
rect 44550 5414 44596 5466
rect 44300 5412 44356 5414
rect 44380 5412 44436 5414
rect 44460 5412 44516 5414
rect 44540 5412 44596 5414
rect 44822 4392 44878 4448
rect 44300 4378 44356 4380
rect 44380 4378 44436 4380
rect 44460 4378 44516 4380
rect 44540 4378 44596 4380
rect 44300 4326 44346 4378
rect 44346 4326 44356 4378
rect 44380 4326 44410 4378
rect 44410 4326 44422 4378
rect 44422 4326 44436 4378
rect 44460 4326 44474 4378
rect 44474 4326 44486 4378
rect 44486 4326 44516 4378
rect 44540 4326 44550 4378
rect 44550 4326 44596 4378
rect 44300 4324 44356 4326
rect 44380 4324 44436 4326
rect 44460 4324 44516 4326
rect 44540 4324 44596 4326
rect 44086 4256 44142 4312
rect 43718 3304 43774 3360
rect 42982 1264 43038 1320
rect 44086 3168 44142 3224
rect 43810 3068 43812 3088
rect 43812 3068 43864 3088
rect 43864 3068 43866 3088
rect 43810 3032 43866 3068
rect 43902 2488 43958 2544
rect 44454 3984 44510 4040
rect 44300 3290 44356 3292
rect 44380 3290 44436 3292
rect 44460 3290 44516 3292
rect 44540 3290 44596 3292
rect 44300 3238 44346 3290
rect 44346 3238 44356 3290
rect 44380 3238 44410 3290
rect 44410 3238 44422 3290
rect 44422 3238 44436 3290
rect 44460 3238 44474 3290
rect 44474 3238 44486 3290
rect 44486 3238 44516 3290
rect 44540 3238 44550 3290
rect 44550 3238 44596 3290
rect 44300 3236 44356 3238
rect 44380 3236 44436 3238
rect 44460 3236 44516 3238
rect 44540 3236 44596 3238
rect 44086 2488 44142 2544
rect 44300 2202 44356 2204
rect 44380 2202 44436 2204
rect 44460 2202 44516 2204
rect 44540 2202 44596 2204
rect 44300 2150 44346 2202
rect 44346 2150 44356 2202
rect 44380 2150 44410 2202
rect 44410 2150 44422 2202
rect 44422 2150 44436 2202
rect 44460 2150 44474 2202
rect 44474 2150 44486 2202
rect 44486 2150 44516 2202
rect 44540 2150 44550 2202
rect 44550 2150 44596 2202
rect 44300 2148 44356 2150
rect 44380 2148 44436 2150
rect 44460 2148 44516 2150
rect 44540 2148 44596 2150
rect 45466 5208 45522 5264
rect 45650 5752 45706 5808
rect 51524 7098 51580 7100
rect 51604 7098 51660 7100
rect 51684 7098 51740 7100
rect 51764 7098 51820 7100
rect 51524 7046 51570 7098
rect 51570 7046 51580 7098
rect 51604 7046 51634 7098
rect 51634 7046 51646 7098
rect 51646 7046 51660 7098
rect 51684 7046 51698 7098
rect 51698 7046 51710 7098
rect 51710 7046 51740 7098
rect 51764 7046 51774 7098
rect 51774 7046 51820 7098
rect 51524 7044 51580 7046
rect 51604 7044 51660 7046
rect 51684 7044 51740 7046
rect 51764 7044 51820 7046
rect 51262 6996 51318 7032
rect 51262 6976 51264 6996
rect 51264 6976 51316 6996
rect 51316 6976 51318 6996
rect 52182 6840 52238 6896
rect 51524 6010 51580 6012
rect 51604 6010 51660 6012
rect 51684 6010 51740 6012
rect 51764 6010 51820 6012
rect 51524 5958 51570 6010
rect 51570 5958 51580 6010
rect 51604 5958 51634 6010
rect 51634 5958 51646 6010
rect 51646 5958 51660 6010
rect 51684 5958 51698 6010
rect 51698 5958 51710 6010
rect 51710 5958 51740 6010
rect 51764 5958 51774 6010
rect 51774 5958 51820 6010
rect 51524 5956 51580 5958
rect 51604 5956 51660 5958
rect 51684 5956 51740 5958
rect 51764 5956 51820 5958
rect 50802 5888 50858 5944
rect 46202 4800 46258 4856
rect 45650 3440 45706 3496
rect 45742 2916 45798 2952
rect 45742 2896 45744 2916
rect 45744 2896 45796 2916
rect 45796 2896 45798 2916
rect 46754 3984 46810 4040
rect 46570 3848 46626 3904
rect 48410 4664 48466 4720
rect 51078 5072 51134 5128
rect 48502 4392 48558 4448
rect 47582 3712 47638 3768
rect 47858 2624 47914 2680
rect 48318 3032 48374 3088
rect 48502 3032 48558 3088
rect 49514 2388 49516 2408
rect 49516 2388 49568 2408
rect 49568 2388 49570 2408
rect 49514 2352 49570 2388
rect 48870 1808 48926 1864
rect 49974 2796 49976 2816
rect 49976 2796 50028 2816
rect 50028 2796 50030 2816
rect 49974 2760 50030 2796
rect 50158 2624 50214 2680
rect 50158 1944 50214 2000
rect 51524 4922 51580 4924
rect 51604 4922 51660 4924
rect 51684 4922 51740 4924
rect 51764 4922 51820 4924
rect 51524 4870 51570 4922
rect 51570 4870 51580 4922
rect 51604 4870 51634 4922
rect 51634 4870 51646 4922
rect 51646 4870 51660 4922
rect 51684 4870 51698 4922
rect 51698 4870 51710 4922
rect 51710 4870 51740 4922
rect 51764 4870 51774 4922
rect 51774 4870 51820 4922
rect 51524 4868 51580 4870
rect 51604 4868 51660 4870
rect 51684 4868 51740 4870
rect 51764 4868 51820 4870
rect 52090 4120 52146 4176
rect 50526 2896 50582 2952
rect 51814 3984 51870 4040
rect 51524 3834 51580 3836
rect 51604 3834 51660 3836
rect 51684 3834 51740 3836
rect 51764 3834 51820 3836
rect 51524 3782 51570 3834
rect 51570 3782 51580 3834
rect 51604 3782 51634 3834
rect 51634 3782 51646 3834
rect 51646 3782 51660 3834
rect 51684 3782 51698 3834
rect 51698 3782 51710 3834
rect 51710 3782 51740 3834
rect 51764 3782 51774 3834
rect 51774 3782 51820 3834
rect 51524 3780 51580 3782
rect 51604 3780 51660 3782
rect 51684 3780 51740 3782
rect 51764 3780 51820 3782
rect 51262 1128 51318 1184
rect 51524 2746 51580 2748
rect 51604 2746 51660 2748
rect 51684 2746 51740 2748
rect 51764 2746 51820 2748
rect 51524 2694 51570 2746
rect 51570 2694 51580 2746
rect 51604 2694 51634 2746
rect 51634 2694 51646 2746
rect 51646 2694 51660 2746
rect 51684 2694 51698 2746
rect 51698 2694 51710 2746
rect 51710 2694 51740 2746
rect 51764 2694 51774 2746
rect 51774 2694 51820 2746
rect 51524 2692 51580 2694
rect 51604 2692 51660 2694
rect 51684 2692 51740 2694
rect 51764 2692 51820 2694
rect 53102 5752 53158 5808
rect 52458 3984 52514 4040
rect 52090 2508 52146 2544
rect 52090 2488 52092 2508
rect 52092 2488 52144 2508
rect 52144 2488 52146 2508
rect 53562 4564 53564 4584
rect 53564 4564 53616 4584
rect 53616 4564 53618 4584
rect 53562 4528 53618 4564
rect 53838 2916 53894 2952
rect 53838 2896 53840 2916
rect 53840 2896 53892 2916
rect 53892 2896 53894 2916
rect 55218 4004 55274 4040
rect 55218 3984 55220 4004
rect 55220 3984 55272 4004
rect 55272 3984 55274 4004
rect 54114 3052 54170 3088
rect 54114 3032 54116 3052
rect 54116 3032 54168 3052
rect 54168 3032 54170 3052
rect 53930 1536 53986 1592
<< metal3 >>
rect 15394 17440 15710 17441
rect 15394 17376 15400 17440
rect 15464 17376 15480 17440
rect 15544 17376 15560 17440
rect 15624 17376 15640 17440
rect 15704 17376 15710 17440
rect 15394 17375 15710 17376
rect 29842 17440 30158 17441
rect 29842 17376 29848 17440
rect 29912 17376 29928 17440
rect 29992 17376 30008 17440
rect 30072 17376 30088 17440
rect 30152 17376 30158 17440
rect 29842 17375 30158 17376
rect 44290 17440 44606 17441
rect 44290 17376 44296 17440
rect 44360 17376 44376 17440
rect 44440 17376 44456 17440
rect 44520 17376 44536 17440
rect 44600 17376 44606 17440
rect 44290 17375 44606 17376
rect 8170 16896 8486 16897
rect 8170 16832 8176 16896
rect 8240 16832 8256 16896
rect 8320 16832 8336 16896
rect 8400 16832 8416 16896
rect 8480 16832 8486 16896
rect 8170 16831 8486 16832
rect 22618 16896 22934 16897
rect 22618 16832 22624 16896
rect 22688 16832 22704 16896
rect 22768 16832 22784 16896
rect 22848 16832 22864 16896
rect 22928 16832 22934 16896
rect 22618 16831 22934 16832
rect 37066 16896 37382 16897
rect 37066 16832 37072 16896
rect 37136 16832 37152 16896
rect 37216 16832 37232 16896
rect 37296 16832 37312 16896
rect 37376 16832 37382 16896
rect 37066 16831 37382 16832
rect 51514 16896 51830 16897
rect 51514 16832 51520 16896
rect 51584 16832 51600 16896
rect 51664 16832 51680 16896
rect 51744 16832 51760 16896
rect 51824 16832 51830 16896
rect 51514 16831 51830 16832
rect 15394 16352 15710 16353
rect 15394 16288 15400 16352
rect 15464 16288 15480 16352
rect 15544 16288 15560 16352
rect 15624 16288 15640 16352
rect 15704 16288 15710 16352
rect 15394 16287 15710 16288
rect 29842 16352 30158 16353
rect 29842 16288 29848 16352
rect 29912 16288 29928 16352
rect 29992 16288 30008 16352
rect 30072 16288 30088 16352
rect 30152 16288 30158 16352
rect 29842 16287 30158 16288
rect 44290 16352 44606 16353
rect 44290 16288 44296 16352
rect 44360 16288 44376 16352
rect 44440 16288 44456 16352
rect 44520 16288 44536 16352
rect 44600 16288 44606 16352
rect 44290 16287 44606 16288
rect 8170 15808 8486 15809
rect 8170 15744 8176 15808
rect 8240 15744 8256 15808
rect 8320 15744 8336 15808
rect 8400 15744 8416 15808
rect 8480 15744 8486 15808
rect 8170 15743 8486 15744
rect 22618 15808 22934 15809
rect 22618 15744 22624 15808
rect 22688 15744 22704 15808
rect 22768 15744 22784 15808
rect 22848 15744 22864 15808
rect 22928 15744 22934 15808
rect 22618 15743 22934 15744
rect 37066 15808 37382 15809
rect 37066 15744 37072 15808
rect 37136 15744 37152 15808
rect 37216 15744 37232 15808
rect 37296 15744 37312 15808
rect 37376 15744 37382 15808
rect 37066 15743 37382 15744
rect 51514 15808 51830 15809
rect 51514 15744 51520 15808
rect 51584 15744 51600 15808
rect 51664 15744 51680 15808
rect 51744 15744 51760 15808
rect 51824 15744 51830 15808
rect 51514 15743 51830 15744
rect 15394 15264 15710 15265
rect 15394 15200 15400 15264
rect 15464 15200 15480 15264
rect 15544 15200 15560 15264
rect 15624 15200 15640 15264
rect 15704 15200 15710 15264
rect 15394 15199 15710 15200
rect 29842 15264 30158 15265
rect 29842 15200 29848 15264
rect 29912 15200 29928 15264
rect 29992 15200 30008 15264
rect 30072 15200 30088 15264
rect 30152 15200 30158 15264
rect 29842 15199 30158 15200
rect 44290 15264 44606 15265
rect 44290 15200 44296 15264
rect 44360 15200 44376 15264
rect 44440 15200 44456 15264
rect 44520 15200 44536 15264
rect 44600 15200 44606 15264
rect 44290 15199 44606 15200
rect 8170 14720 8486 14721
rect 8170 14656 8176 14720
rect 8240 14656 8256 14720
rect 8320 14656 8336 14720
rect 8400 14656 8416 14720
rect 8480 14656 8486 14720
rect 8170 14655 8486 14656
rect 22618 14720 22934 14721
rect 22618 14656 22624 14720
rect 22688 14656 22704 14720
rect 22768 14656 22784 14720
rect 22848 14656 22864 14720
rect 22928 14656 22934 14720
rect 22618 14655 22934 14656
rect 37066 14720 37382 14721
rect 37066 14656 37072 14720
rect 37136 14656 37152 14720
rect 37216 14656 37232 14720
rect 37296 14656 37312 14720
rect 37376 14656 37382 14720
rect 37066 14655 37382 14656
rect 51514 14720 51830 14721
rect 51514 14656 51520 14720
rect 51584 14656 51600 14720
rect 51664 14656 51680 14720
rect 51744 14656 51760 14720
rect 51824 14656 51830 14720
rect 51514 14655 51830 14656
rect 15394 14176 15710 14177
rect 15394 14112 15400 14176
rect 15464 14112 15480 14176
rect 15544 14112 15560 14176
rect 15624 14112 15640 14176
rect 15704 14112 15710 14176
rect 15394 14111 15710 14112
rect 29842 14176 30158 14177
rect 29842 14112 29848 14176
rect 29912 14112 29928 14176
rect 29992 14112 30008 14176
rect 30072 14112 30088 14176
rect 30152 14112 30158 14176
rect 29842 14111 30158 14112
rect 44290 14176 44606 14177
rect 44290 14112 44296 14176
rect 44360 14112 44376 14176
rect 44440 14112 44456 14176
rect 44520 14112 44536 14176
rect 44600 14112 44606 14176
rect 44290 14111 44606 14112
rect 13353 13836 13419 13837
rect 13302 13834 13308 13836
rect 13262 13774 13308 13834
rect 13372 13832 13419 13836
rect 13414 13776 13419 13832
rect 13302 13772 13308 13774
rect 13372 13772 13419 13776
rect 13353 13771 13419 13772
rect 8170 13632 8486 13633
rect 8170 13568 8176 13632
rect 8240 13568 8256 13632
rect 8320 13568 8336 13632
rect 8400 13568 8416 13632
rect 8480 13568 8486 13632
rect 8170 13567 8486 13568
rect 22618 13632 22934 13633
rect 22618 13568 22624 13632
rect 22688 13568 22704 13632
rect 22768 13568 22784 13632
rect 22848 13568 22864 13632
rect 22928 13568 22934 13632
rect 22618 13567 22934 13568
rect 37066 13632 37382 13633
rect 37066 13568 37072 13632
rect 37136 13568 37152 13632
rect 37216 13568 37232 13632
rect 37296 13568 37312 13632
rect 37376 13568 37382 13632
rect 37066 13567 37382 13568
rect 51514 13632 51830 13633
rect 51514 13568 51520 13632
rect 51584 13568 51600 13632
rect 51664 13568 51680 13632
rect 51744 13568 51760 13632
rect 51824 13568 51830 13632
rect 51514 13567 51830 13568
rect 17769 13156 17835 13157
rect 17718 13092 17724 13156
rect 17788 13154 17835 13156
rect 17788 13152 17880 13154
rect 17830 13096 17880 13152
rect 17788 13094 17880 13096
rect 17788 13092 17835 13094
rect 17769 13091 17835 13092
rect 15394 13088 15710 13089
rect 15394 13024 15400 13088
rect 15464 13024 15480 13088
rect 15544 13024 15560 13088
rect 15624 13024 15640 13088
rect 15704 13024 15710 13088
rect 15394 13023 15710 13024
rect 29842 13088 30158 13089
rect 29842 13024 29848 13088
rect 29912 13024 29928 13088
rect 29992 13024 30008 13088
rect 30072 13024 30088 13088
rect 30152 13024 30158 13088
rect 29842 13023 30158 13024
rect 44290 13088 44606 13089
rect 44290 13024 44296 13088
rect 44360 13024 44376 13088
rect 44440 13024 44456 13088
rect 44520 13024 44536 13088
rect 44600 13024 44606 13088
rect 44290 13023 44606 13024
rect 10726 12684 10732 12748
rect 10796 12746 10802 12748
rect 11421 12746 11487 12749
rect 10796 12744 11487 12746
rect 10796 12688 11426 12744
rect 11482 12688 11487 12744
rect 10796 12686 11487 12688
rect 10796 12684 10802 12686
rect 11421 12683 11487 12686
rect 14181 12746 14247 12749
rect 14590 12746 14596 12748
rect 14181 12744 14596 12746
rect 14181 12688 14186 12744
rect 14242 12688 14596 12744
rect 14181 12686 14596 12688
rect 14181 12683 14247 12686
rect 14590 12684 14596 12686
rect 14660 12684 14666 12748
rect 10961 12612 11027 12613
rect 10910 12548 10916 12612
rect 10980 12610 11027 12612
rect 18229 12610 18295 12613
rect 19190 12610 19196 12612
rect 10980 12608 11072 12610
rect 11022 12552 11072 12608
rect 10980 12550 11072 12552
rect 18229 12608 19196 12610
rect 18229 12552 18234 12608
rect 18290 12552 19196 12608
rect 18229 12550 19196 12552
rect 10980 12548 11027 12550
rect 10961 12547 11027 12548
rect 18229 12547 18295 12550
rect 19190 12548 19196 12550
rect 19260 12548 19266 12612
rect 8170 12544 8486 12545
rect 8170 12480 8176 12544
rect 8240 12480 8256 12544
rect 8320 12480 8336 12544
rect 8400 12480 8416 12544
rect 8480 12480 8486 12544
rect 8170 12479 8486 12480
rect 22618 12544 22934 12545
rect 22618 12480 22624 12544
rect 22688 12480 22704 12544
rect 22768 12480 22784 12544
rect 22848 12480 22864 12544
rect 22928 12480 22934 12544
rect 22618 12479 22934 12480
rect 37066 12544 37382 12545
rect 37066 12480 37072 12544
rect 37136 12480 37152 12544
rect 37216 12480 37232 12544
rect 37296 12480 37312 12544
rect 37376 12480 37382 12544
rect 37066 12479 37382 12480
rect 51514 12544 51830 12545
rect 51514 12480 51520 12544
rect 51584 12480 51600 12544
rect 51664 12480 51680 12544
rect 51744 12480 51760 12544
rect 51824 12480 51830 12544
rect 51514 12479 51830 12480
rect 1945 12476 2011 12477
rect 1894 12474 1900 12476
rect 1854 12414 1900 12474
rect 1964 12472 2011 12476
rect 2006 12416 2011 12472
rect 1894 12412 1900 12414
rect 1964 12412 2011 12416
rect 2814 12412 2820 12476
rect 2884 12474 2890 12476
rect 3785 12474 3851 12477
rect 2884 12472 3851 12474
rect 2884 12416 3790 12472
rect 3846 12416 3851 12472
rect 2884 12414 3851 12416
rect 2884 12412 2890 12414
rect 1945 12411 2011 12412
rect 3785 12411 3851 12414
rect 6678 12412 6684 12476
rect 6748 12474 6754 12476
rect 7005 12474 7071 12477
rect 6748 12472 7071 12474
rect 6748 12416 7010 12472
rect 7066 12416 7071 12472
rect 6748 12414 7071 12416
rect 6748 12412 6754 12414
rect 7005 12411 7071 12414
rect 16113 12474 16179 12477
rect 23473 12476 23539 12477
rect 16982 12474 16988 12476
rect 16113 12472 16988 12474
rect 16113 12416 16118 12472
rect 16174 12416 16988 12472
rect 16113 12414 16988 12416
rect 16113 12411 16179 12414
rect 16982 12412 16988 12414
rect 17052 12412 17058 12476
rect 23422 12474 23428 12476
rect 23382 12414 23428 12474
rect 23492 12472 23539 12476
rect 23534 12416 23539 12472
rect 23422 12412 23428 12414
rect 23492 12412 23539 12416
rect 23473 12411 23539 12412
rect 14181 12068 14247 12069
rect 18597 12068 18663 12069
rect 22277 12068 22343 12069
rect 14181 12066 14228 12068
rect 14136 12064 14228 12066
rect 14136 12008 14186 12064
rect 14136 12006 14228 12008
rect 14181 12004 14228 12006
rect 14292 12004 14298 12068
rect 18597 12066 18644 12068
rect 18552 12064 18644 12066
rect 18552 12008 18602 12064
rect 18552 12006 18644 12008
rect 18597 12004 18644 12006
rect 18708 12004 18714 12068
rect 22277 12066 22324 12068
rect 22232 12064 22324 12066
rect 22232 12008 22282 12064
rect 22232 12006 22324 12008
rect 22277 12004 22324 12006
rect 22388 12004 22394 12068
rect 14181 12003 14247 12004
rect 18597 12003 18663 12004
rect 22277 12003 22343 12004
rect 15394 12000 15710 12001
rect 15394 11936 15400 12000
rect 15464 11936 15480 12000
rect 15544 11936 15560 12000
rect 15624 11936 15640 12000
rect 15704 11936 15710 12000
rect 15394 11935 15710 11936
rect 29842 12000 30158 12001
rect 29842 11936 29848 12000
rect 29912 11936 29928 12000
rect 29992 11936 30008 12000
rect 30072 11936 30088 12000
rect 30152 11936 30158 12000
rect 29842 11935 30158 11936
rect 44290 12000 44606 12001
rect 44290 11936 44296 12000
rect 44360 11936 44376 12000
rect 44440 11936 44456 12000
rect 44520 11936 44536 12000
rect 44600 11936 44606 12000
rect 44290 11935 44606 11936
rect 1761 11794 1827 11797
rect 14590 11794 14596 11796
rect 1761 11792 14596 11794
rect 1761 11736 1766 11792
rect 1822 11736 14596 11792
rect 1761 11734 14596 11736
rect 1761 11731 1827 11734
rect 14590 11732 14596 11734
rect 14660 11732 14666 11796
rect 5809 11522 5875 11525
rect 22093 11524 22159 11525
rect 5942 11522 5948 11524
rect 5809 11520 5948 11522
rect 5809 11464 5814 11520
rect 5870 11464 5948 11520
rect 5809 11462 5948 11464
rect 5809 11459 5875 11462
rect 5942 11460 5948 11462
rect 6012 11460 6018 11524
rect 22093 11520 22140 11524
rect 22204 11522 22210 11524
rect 22093 11464 22098 11520
rect 22093 11460 22140 11464
rect 22204 11462 22250 11522
rect 22204 11460 22210 11462
rect 22093 11459 22159 11460
rect 8170 11456 8486 11457
rect 8170 11392 8176 11456
rect 8240 11392 8256 11456
rect 8320 11392 8336 11456
rect 8400 11392 8416 11456
rect 8480 11392 8486 11456
rect 8170 11391 8486 11392
rect 22618 11456 22934 11457
rect 22618 11392 22624 11456
rect 22688 11392 22704 11456
rect 22768 11392 22784 11456
rect 22848 11392 22864 11456
rect 22928 11392 22934 11456
rect 22618 11391 22934 11392
rect 37066 11456 37382 11457
rect 37066 11392 37072 11456
rect 37136 11392 37152 11456
rect 37216 11392 37232 11456
rect 37296 11392 37312 11456
rect 37376 11392 37382 11456
rect 37066 11391 37382 11392
rect 51514 11456 51830 11457
rect 51514 11392 51520 11456
rect 51584 11392 51600 11456
rect 51664 11392 51680 11456
rect 51744 11392 51760 11456
rect 51824 11392 51830 11456
rect 51514 11391 51830 11392
rect 2037 11250 2103 11253
rect 12934 11250 12940 11252
rect 2037 11248 12940 11250
rect 2037 11192 2042 11248
rect 2098 11192 12940 11248
rect 2037 11190 12940 11192
rect 2037 11187 2103 11190
rect 12934 11188 12940 11190
rect 13004 11188 13010 11252
rect 4654 11052 4660 11116
rect 4724 11114 4730 11116
rect 7741 11114 7807 11117
rect 15101 11116 15167 11117
rect 15101 11114 15148 11116
rect 4724 11112 7807 11114
rect 4724 11056 7746 11112
rect 7802 11056 7807 11112
rect 4724 11054 7807 11056
rect 15056 11112 15148 11114
rect 15056 11056 15106 11112
rect 15056 11054 15148 11056
rect 4724 11052 4730 11054
rect 7741 11051 7807 11054
rect 15101 11052 15148 11054
rect 15212 11052 15218 11116
rect 15653 11114 15719 11117
rect 18270 11114 18276 11116
rect 15653 11112 18276 11114
rect 15653 11056 15658 11112
rect 15714 11056 18276 11112
rect 15653 11054 18276 11056
rect 15101 11051 15167 11052
rect 15653 11051 15719 11054
rect 18270 11052 18276 11054
rect 18340 11052 18346 11116
rect 23054 11052 23060 11116
rect 23124 11114 23130 11116
rect 23933 11114 23999 11117
rect 23124 11112 23999 11114
rect 23124 11056 23938 11112
rect 23994 11056 23999 11112
rect 23124 11054 23999 11056
rect 23124 11052 23130 11054
rect 23933 11051 23999 11054
rect 35709 11116 35775 11117
rect 35709 11112 35756 11116
rect 35820 11114 35826 11116
rect 35709 11056 35714 11112
rect 35709 11052 35756 11056
rect 35820 11054 35866 11114
rect 35820 11052 35826 11054
rect 35709 11051 35775 11052
rect 15394 10912 15710 10913
rect 15394 10848 15400 10912
rect 15464 10848 15480 10912
rect 15544 10848 15560 10912
rect 15624 10848 15640 10912
rect 15704 10848 15710 10912
rect 15394 10847 15710 10848
rect 29842 10912 30158 10913
rect 29842 10848 29848 10912
rect 29912 10848 29928 10912
rect 29992 10848 30008 10912
rect 30072 10848 30088 10912
rect 30152 10848 30158 10912
rect 29842 10847 30158 10848
rect 44290 10912 44606 10913
rect 44290 10848 44296 10912
rect 44360 10848 44376 10912
rect 44440 10848 44456 10912
rect 44520 10848 44536 10912
rect 44600 10848 44606 10912
rect 44290 10847 44606 10848
rect 1577 10570 1643 10573
rect 9254 10570 9260 10572
rect 1577 10568 9260 10570
rect 1577 10512 1582 10568
rect 1638 10512 9260 10568
rect 1577 10510 9260 10512
rect 1577 10507 1643 10510
rect 9254 10508 9260 10510
rect 9324 10508 9330 10572
rect 8170 10368 8486 10369
rect 8170 10304 8176 10368
rect 8240 10304 8256 10368
rect 8320 10304 8336 10368
rect 8400 10304 8416 10368
rect 8480 10304 8486 10368
rect 8170 10303 8486 10304
rect 22618 10368 22934 10369
rect 22618 10304 22624 10368
rect 22688 10304 22704 10368
rect 22768 10304 22784 10368
rect 22848 10304 22864 10368
rect 22928 10304 22934 10368
rect 22618 10303 22934 10304
rect 37066 10368 37382 10369
rect 37066 10304 37072 10368
rect 37136 10304 37152 10368
rect 37216 10304 37232 10368
rect 37296 10304 37312 10368
rect 37376 10304 37382 10368
rect 37066 10303 37382 10304
rect 51514 10368 51830 10369
rect 51514 10304 51520 10368
rect 51584 10304 51600 10368
rect 51664 10304 51680 10368
rect 51744 10304 51760 10368
rect 51824 10304 51830 10368
rect 51514 10303 51830 10304
rect 4153 10162 4219 10165
rect 16614 10162 16620 10164
rect 4153 10160 16620 10162
rect 4153 10104 4158 10160
rect 4214 10104 16620 10160
rect 4153 10102 16620 10104
rect 4153 10099 4219 10102
rect 16614 10100 16620 10102
rect 16684 10100 16690 10164
rect 9070 10026 9076 10028
rect 7974 9966 9076 10026
rect 2497 9890 2563 9893
rect 7974 9890 8034 9966
rect 9070 9964 9076 9966
rect 9140 9964 9146 10028
rect 10910 9964 10916 10028
rect 10980 10026 10986 10028
rect 13169 10026 13235 10029
rect 10980 10024 13235 10026
rect 10980 9968 13174 10024
rect 13230 9968 13235 10024
rect 10980 9966 13235 9968
rect 10980 9964 10986 9966
rect 13169 9963 13235 9966
rect 13445 10026 13511 10029
rect 15469 10026 15535 10029
rect 13445 10024 15535 10026
rect 13445 9968 13450 10024
rect 13506 9968 15474 10024
rect 15530 9968 15535 10024
rect 13445 9966 15535 9968
rect 13445 9963 13511 9966
rect 15469 9963 15535 9966
rect 8886 9890 8892 9892
rect 2497 9888 8034 9890
rect 2497 9832 2502 9888
rect 2558 9832 8034 9888
rect 2497 9830 8034 9832
rect 8158 9830 8892 9890
rect 2497 9827 2563 9830
rect 1853 9754 1919 9757
rect 8158 9754 8218 9830
rect 8886 9828 8892 9830
rect 8956 9828 8962 9892
rect 15394 9824 15710 9825
rect 15394 9760 15400 9824
rect 15464 9760 15480 9824
rect 15544 9760 15560 9824
rect 15624 9760 15640 9824
rect 15704 9760 15710 9824
rect 15394 9759 15710 9760
rect 29842 9824 30158 9825
rect 29842 9760 29848 9824
rect 29912 9760 29928 9824
rect 29992 9760 30008 9824
rect 30072 9760 30088 9824
rect 30152 9760 30158 9824
rect 29842 9759 30158 9760
rect 44290 9824 44606 9825
rect 44290 9760 44296 9824
rect 44360 9760 44376 9824
rect 44440 9760 44456 9824
rect 44520 9760 44536 9824
rect 44600 9760 44606 9824
rect 44290 9759 44606 9760
rect 1853 9752 8218 9754
rect 1853 9696 1858 9752
rect 1914 9696 8218 9752
rect 1853 9694 8218 9696
rect 1853 9691 1919 9694
rect 8702 9692 8708 9756
rect 8772 9754 8778 9756
rect 9765 9754 9831 9757
rect 8772 9752 9831 9754
rect 8772 9696 9770 9752
rect 9826 9696 9831 9752
rect 8772 9694 9831 9696
rect 8772 9692 8778 9694
rect 9765 9691 9831 9694
rect 5073 9618 5139 9621
rect 9857 9618 9923 9621
rect 13445 9618 13511 9621
rect 5073 9616 13511 9618
rect 5073 9560 5078 9616
rect 5134 9560 9862 9616
rect 9918 9560 13450 9616
rect 13506 9560 13511 9616
rect 5073 9558 13511 9560
rect 5073 9555 5139 9558
rect 9857 9555 9923 9558
rect 13445 9555 13511 9558
rect 14181 9618 14247 9621
rect 15377 9618 15443 9621
rect 17861 9618 17927 9621
rect 28441 9618 28507 9621
rect 14181 9616 28507 9618
rect 14181 9560 14186 9616
rect 14242 9560 15382 9616
rect 15438 9560 17866 9616
rect 17922 9560 28446 9616
rect 28502 9560 28507 9616
rect 14181 9558 28507 9560
rect 14181 9555 14247 9558
rect 15377 9555 15443 9558
rect 17861 9555 17927 9558
rect 28441 9555 28507 9558
rect 10317 9482 10383 9485
rect 24209 9482 24275 9485
rect 10317 9480 24275 9482
rect 10317 9424 10322 9480
rect 10378 9424 24214 9480
rect 24270 9424 24275 9480
rect 10317 9422 24275 9424
rect 10317 9419 10383 9422
rect 24209 9419 24275 9422
rect 14181 9346 14247 9349
rect 18965 9346 19031 9349
rect 14181 9344 19031 9346
rect 14181 9288 14186 9344
rect 14242 9288 18970 9344
rect 19026 9288 19031 9344
rect 14181 9286 19031 9288
rect 14181 9283 14247 9286
rect 18965 9283 19031 9286
rect 8170 9280 8486 9281
rect 8170 9216 8176 9280
rect 8240 9216 8256 9280
rect 8320 9216 8336 9280
rect 8400 9216 8416 9280
rect 8480 9216 8486 9280
rect 8170 9215 8486 9216
rect 22618 9280 22934 9281
rect 22618 9216 22624 9280
rect 22688 9216 22704 9280
rect 22768 9216 22784 9280
rect 22848 9216 22864 9280
rect 22928 9216 22934 9280
rect 22618 9215 22934 9216
rect 37066 9280 37382 9281
rect 37066 9216 37072 9280
rect 37136 9216 37152 9280
rect 37216 9216 37232 9280
rect 37296 9216 37312 9280
rect 37376 9216 37382 9280
rect 37066 9215 37382 9216
rect 51514 9280 51830 9281
rect 51514 9216 51520 9280
rect 51584 9216 51600 9280
rect 51664 9216 51680 9280
rect 51744 9216 51760 9280
rect 51824 9216 51830 9280
rect 51514 9215 51830 9216
rect 17585 9210 17651 9213
rect 17861 9210 17927 9213
rect 35525 9210 35591 9213
rect 17585 9208 17927 9210
rect 17585 9152 17590 9208
rect 17646 9152 17866 9208
rect 17922 9152 17927 9208
rect 17585 9150 17927 9152
rect 17585 9147 17651 9150
rect 17861 9147 17927 9150
rect 26926 9208 35591 9210
rect 26926 9152 35530 9208
rect 35586 9152 35591 9208
rect 26926 9150 35591 9152
rect 11145 9074 11211 9077
rect 26785 9074 26851 9077
rect 11145 9072 26851 9074
rect 11145 9016 11150 9072
rect 11206 9016 26790 9072
rect 26846 9016 26851 9072
rect 11145 9014 26851 9016
rect 11145 9011 11211 9014
rect 26785 9011 26851 9014
rect 10593 8938 10659 8941
rect 17861 8938 17927 8941
rect 10593 8936 17927 8938
rect 10593 8880 10598 8936
rect 10654 8880 17866 8936
rect 17922 8880 17927 8936
rect 10593 8878 17927 8880
rect 10593 8875 10659 8878
rect 17861 8875 17927 8878
rect 21081 8938 21147 8941
rect 26926 8938 26986 9150
rect 35525 9147 35591 9150
rect 28993 9074 29059 9077
rect 44265 9074 44331 9077
rect 28993 9072 44331 9074
rect 28993 9016 28998 9072
rect 29054 9016 44270 9072
rect 44326 9016 44331 9072
rect 28993 9014 44331 9016
rect 28993 9011 29059 9014
rect 44265 9011 44331 9014
rect 21081 8936 26986 8938
rect 21081 8880 21086 8936
rect 21142 8880 26986 8936
rect 21081 8878 26986 8880
rect 27153 8938 27219 8941
rect 44633 8938 44699 8941
rect 27153 8936 44699 8938
rect 27153 8880 27158 8936
rect 27214 8880 44638 8936
rect 44694 8880 44699 8936
rect 27153 8878 44699 8880
rect 21081 8875 21147 8878
rect 27153 8875 27219 8878
rect 44633 8875 44699 8878
rect 19517 8802 19583 8805
rect 27981 8802 28047 8805
rect 19517 8800 28047 8802
rect 19517 8744 19522 8800
rect 19578 8744 27986 8800
rect 28042 8744 28047 8800
rect 19517 8742 28047 8744
rect 19517 8739 19583 8742
rect 27981 8739 28047 8742
rect 15394 8736 15710 8737
rect 15394 8672 15400 8736
rect 15464 8672 15480 8736
rect 15544 8672 15560 8736
rect 15624 8672 15640 8736
rect 15704 8672 15710 8736
rect 15394 8671 15710 8672
rect 29842 8736 30158 8737
rect 29842 8672 29848 8736
rect 29912 8672 29928 8736
rect 29992 8672 30008 8736
rect 30072 8672 30088 8736
rect 30152 8672 30158 8736
rect 29842 8671 30158 8672
rect 44290 8736 44606 8737
rect 44290 8672 44296 8736
rect 44360 8672 44376 8736
rect 44440 8672 44456 8736
rect 44520 8672 44536 8736
rect 44600 8672 44606 8736
rect 44290 8671 44606 8672
rect 6085 8666 6151 8669
rect 9489 8666 9555 8669
rect 6085 8664 9555 8666
rect 6085 8608 6090 8664
rect 6146 8608 9494 8664
rect 9550 8608 9555 8664
rect 6085 8606 9555 8608
rect 6085 8603 6151 8606
rect 9489 8603 9555 8606
rect 20253 8666 20319 8669
rect 24393 8666 24459 8669
rect 20253 8664 24459 8666
rect 20253 8608 20258 8664
rect 20314 8608 24398 8664
rect 24454 8608 24459 8664
rect 20253 8606 24459 8608
rect 20253 8603 20319 8606
rect 24393 8603 24459 8606
rect 17769 8530 17835 8533
rect 22093 8530 22159 8533
rect 17769 8528 22159 8530
rect 17769 8472 17774 8528
rect 17830 8472 22098 8528
rect 22154 8472 22159 8528
rect 17769 8470 22159 8472
rect 17769 8467 17835 8470
rect 22093 8467 22159 8470
rect 24209 8530 24275 8533
rect 29453 8530 29519 8533
rect 31017 8530 31083 8533
rect 31477 8530 31543 8533
rect 24209 8528 31543 8530
rect 24209 8472 24214 8528
rect 24270 8472 29458 8528
rect 29514 8472 31022 8528
rect 31078 8472 31482 8528
rect 31538 8472 31543 8528
rect 24209 8470 31543 8472
rect 24209 8467 24275 8470
rect 29453 8467 29519 8470
rect 31017 8467 31083 8470
rect 31477 8467 31543 8470
rect 1761 8394 1827 8397
rect 6085 8394 6151 8397
rect 1761 8392 6151 8394
rect 1761 8336 1766 8392
rect 1822 8336 6090 8392
rect 6146 8336 6151 8392
rect 1761 8334 6151 8336
rect 1761 8331 1827 8334
rect 6085 8331 6151 8334
rect 6545 8394 6611 8397
rect 8201 8394 8267 8397
rect 6545 8392 8267 8394
rect 6545 8336 6550 8392
rect 6606 8336 8206 8392
rect 8262 8336 8267 8392
rect 6545 8334 8267 8336
rect 6545 8331 6611 8334
rect 8201 8331 8267 8334
rect 10961 8394 11027 8397
rect 14641 8394 14707 8397
rect 10961 8392 14707 8394
rect 10961 8336 10966 8392
rect 11022 8336 14646 8392
rect 14702 8336 14707 8392
rect 10961 8334 14707 8336
rect 10961 8331 11027 8334
rect 14641 8331 14707 8334
rect 18229 8394 18295 8397
rect 21265 8394 21331 8397
rect 18229 8392 21331 8394
rect 18229 8336 18234 8392
rect 18290 8336 21270 8392
rect 21326 8336 21331 8392
rect 18229 8334 21331 8336
rect 18229 8331 18295 8334
rect 21265 8331 21331 8334
rect 24577 8394 24643 8397
rect 33593 8394 33659 8397
rect 24577 8392 33659 8394
rect 24577 8336 24582 8392
rect 24638 8336 33598 8392
rect 33654 8336 33659 8392
rect 24577 8334 33659 8336
rect 24577 8331 24643 8334
rect 33593 8331 33659 8334
rect 17718 8196 17724 8260
rect 17788 8258 17794 8260
rect 22277 8258 22343 8261
rect 17788 8256 22343 8258
rect 17788 8200 22282 8256
rect 22338 8200 22343 8256
rect 17788 8198 22343 8200
rect 17788 8196 17794 8198
rect 22277 8195 22343 8198
rect 27337 8258 27403 8261
rect 32213 8258 32279 8261
rect 27337 8256 32279 8258
rect 27337 8200 27342 8256
rect 27398 8200 32218 8256
rect 32274 8200 32279 8256
rect 27337 8198 32279 8200
rect 27337 8195 27403 8198
rect 32213 8195 32279 8198
rect 48037 8258 48103 8261
rect 49877 8258 49943 8261
rect 48037 8256 49943 8258
rect 48037 8200 48042 8256
rect 48098 8200 49882 8256
rect 49938 8200 49943 8256
rect 48037 8198 49943 8200
rect 48037 8195 48103 8198
rect 49877 8195 49943 8198
rect 8170 8192 8486 8193
rect 8170 8128 8176 8192
rect 8240 8128 8256 8192
rect 8320 8128 8336 8192
rect 8400 8128 8416 8192
rect 8480 8128 8486 8192
rect 8170 8127 8486 8128
rect 22618 8192 22934 8193
rect 22618 8128 22624 8192
rect 22688 8128 22704 8192
rect 22768 8128 22784 8192
rect 22848 8128 22864 8192
rect 22928 8128 22934 8192
rect 22618 8127 22934 8128
rect 37066 8192 37382 8193
rect 37066 8128 37072 8192
rect 37136 8128 37152 8192
rect 37216 8128 37232 8192
rect 37296 8128 37312 8192
rect 37376 8128 37382 8192
rect 37066 8127 37382 8128
rect 51514 8192 51830 8193
rect 51514 8128 51520 8192
rect 51584 8128 51600 8192
rect 51664 8128 51680 8192
rect 51744 8128 51760 8192
rect 51824 8128 51830 8192
rect 51514 8127 51830 8128
rect 10041 8122 10107 8125
rect 11513 8122 11579 8125
rect 10041 8120 11579 8122
rect 10041 8064 10046 8120
rect 10102 8064 11518 8120
rect 11574 8064 11579 8120
rect 10041 8062 11579 8064
rect 10041 8059 10107 8062
rect 11513 8059 11579 8062
rect 9857 7986 9923 7989
rect 11697 7986 11763 7989
rect 13537 7988 13603 7989
rect 13486 7986 13492 7988
rect 9857 7984 11763 7986
rect 9857 7928 9862 7984
rect 9918 7928 11702 7984
rect 11758 7928 11763 7984
rect 9857 7926 11763 7928
rect 13410 7926 13492 7986
rect 13556 7986 13603 7988
rect 14222 7986 14228 7988
rect 13556 7984 14228 7986
rect 13598 7928 14228 7984
rect 9857 7923 9923 7926
rect 11697 7923 11763 7926
rect 13486 7924 13492 7926
rect 13556 7926 14228 7928
rect 13556 7924 13603 7926
rect 14222 7924 14228 7926
rect 14292 7924 14298 7988
rect 21449 7986 21515 7989
rect 27337 7986 27403 7989
rect 21449 7984 27403 7986
rect 21449 7928 21454 7984
rect 21510 7928 27342 7984
rect 27398 7928 27403 7984
rect 21449 7926 27403 7928
rect 13537 7923 13603 7924
rect 21449 7923 21515 7926
rect 27337 7923 27403 7926
rect 6637 7850 6703 7853
rect 14958 7850 14964 7852
rect 6637 7848 14964 7850
rect 6637 7792 6642 7848
rect 6698 7792 14964 7848
rect 6637 7790 14964 7792
rect 6637 7787 6703 7790
rect 14958 7788 14964 7790
rect 15028 7788 15034 7852
rect 15101 7850 15167 7853
rect 23749 7850 23815 7853
rect 25865 7850 25931 7853
rect 15101 7848 25931 7850
rect 15101 7792 15106 7848
rect 15162 7792 23754 7848
rect 23810 7792 25870 7848
rect 25926 7792 25931 7848
rect 15101 7790 25931 7792
rect 15101 7787 15167 7790
rect 23749 7787 23815 7790
rect 25865 7787 25931 7790
rect 27889 7850 27955 7853
rect 42885 7850 42951 7853
rect 27889 7848 42951 7850
rect 27889 7792 27894 7848
rect 27950 7792 42890 7848
rect 42946 7792 42951 7848
rect 27889 7790 42951 7792
rect 27889 7787 27955 7790
rect 42885 7787 42951 7790
rect 5993 7714 6059 7717
rect 10869 7714 10935 7717
rect 5993 7712 10935 7714
rect 5993 7656 5998 7712
rect 6054 7656 10874 7712
rect 10930 7656 10935 7712
rect 5993 7654 10935 7656
rect 5993 7651 6059 7654
rect 10869 7651 10935 7654
rect 20161 7714 20227 7717
rect 26693 7714 26759 7717
rect 20161 7712 26759 7714
rect 20161 7656 20166 7712
rect 20222 7656 26698 7712
rect 26754 7656 26759 7712
rect 20161 7654 26759 7656
rect 20161 7651 20227 7654
rect 26693 7651 26759 7654
rect 15394 7648 15710 7649
rect 15394 7584 15400 7648
rect 15464 7584 15480 7648
rect 15544 7584 15560 7648
rect 15624 7584 15640 7648
rect 15704 7584 15710 7648
rect 15394 7583 15710 7584
rect 29842 7648 30158 7649
rect 29842 7584 29848 7648
rect 29912 7584 29928 7648
rect 29992 7584 30008 7648
rect 30072 7584 30088 7648
rect 30152 7584 30158 7648
rect 29842 7583 30158 7584
rect 44290 7648 44606 7649
rect 44290 7584 44296 7648
rect 44360 7584 44376 7648
rect 44440 7584 44456 7648
rect 44520 7584 44536 7648
rect 44600 7584 44606 7648
rect 44290 7583 44606 7584
rect 5942 7516 5948 7580
rect 6012 7578 6018 7580
rect 6269 7578 6335 7581
rect 6637 7578 6703 7581
rect 6012 7576 6703 7578
rect 6012 7520 6274 7576
rect 6330 7520 6642 7576
rect 6698 7520 6703 7576
rect 6012 7518 6703 7520
rect 6012 7516 6018 7518
rect 6269 7515 6335 7518
rect 6637 7515 6703 7518
rect 9213 7578 9279 7581
rect 15101 7578 15167 7581
rect 22001 7578 22067 7581
rect 29637 7578 29703 7581
rect 9213 7576 15167 7578
rect 9213 7520 9218 7576
rect 9274 7520 15106 7576
rect 15162 7520 15167 7576
rect 9213 7518 15167 7520
rect 9213 7515 9279 7518
rect 15101 7515 15167 7518
rect 18830 7576 29703 7578
rect 18830 7520 22006 7576
rect 22062 7520 29642 7576
rect 29698 7520 29703 7576
rect 18830 7518 29703 7520
rect 4153 7442 4219 7445
rect 6361 7442 6427 7445
rect 4153 7440 6427 7442
rect 4153 7384 4158 7440
rect 4214 7384 6366 7440
rect 6422 7384 6427 7440
rect 4153 7382 6427 7384
rect 4153 7379 4219 7382
rect 6361 7379 6427 7382
rect 6729 7442 6795 7445
rect 11973 7442 12039 7445
rect 18830 7442 18890 7518
rect 22001 7515 22067 7518
rect 29637 7515 29703 7518
rect 30373 7578 30439 7581
rect 41873 7578 41939 7581
rect 30373 7576 41939 7578
rect 30373 7520 30378 7576
rect 30434 7520 41878 7576
rect 41934 7520 41939 7576
rect 30373 7518 41939 7520
rect 30373 7515 30439 7518
rect 41873 7515 41939 7518
rect 6729 7440 12039 7442
rect 6729 7384 6734 7440
rect 6790 7384 11978 7440
rect 12034 7384 12039 7440
rect 6729 7382 12039 7384
rect 6729 7379 6795 7382
rect 11973 7379 12039 7382
rect 14966 7382 18890 7442
rect 19241 7442 19307 7445
rect 23473 7442 23539 7445
rect 19241 7440 23539 7442
rect 19241 7384 19246 7440
rect 19302 7384 23478 7440
rect 23534 7384 23539 7440
rect 19241 7382 23539 7384
rect 3141 7306 3207 7309
rect 9489 7306 9555 7309
rect 3141 7304 9555 7306
rect 3141 7248 3146 7304
rect 3202 7248 9494 7304
rect 9550 7248 9555 7304
rect 3141 7246 9555 7248
rect 3141 7243 3207 7246
rect 9489 7243 9555 7246
rect 10869 7306 10935 7309
rect 13537 7306 13603 7309
rect 10869 7304 13603 7306
rect 10869 7248 10874 7304
rect 10930 7248 13542 7304
rect 13598 7248 13603 7304
rect 10869 7246 13603 7248
rect 10869 7243 10935 7246
rect 13537 7243 13603 7246
rect 14222 7244 14228 7308
rect 14292 7306 14298 7308
rect 14365 7306 14431 7309
rect 14292 7304 14431 7306
rect 14292 7248 14370 7304
rect 14426 7248 14431 7304
rect 14292 7246 14431 7248
rect 14292 7244 14298 7246
rect 14365 7243 14431 7246
rect 14966 7170 15026 7382
rect 19241 7379 19307 7382
rect 23473 7379 23539 7382
rect 24117 7442 24183 7445
rect 26785 7442 26851 7445
rect 39941 7442 40007 7445
rect 24117 7440 40007 7442
rect 24117 7384 24122 7440
rect 24178 7384 26790 7440
rect 26846 7384 39946 7440
rect 40002 7384 40007 7440
rect 24117 7382 40007 7384
rect 24117 7379 24183 7382
rect 26785 7379 26851 7382
rect 39941 7379 40007 7382
rect 15193 7306 15259 7309
rect 25037 7306 25103 7309
rect 15193 7304 25103 7306
rect 15193 7248 15198 7304
rect 15254 7248 25042 7304
rect 25098 7248 25103 7304
rect 15193 7246 25103 7248
rect 15193 7243 15259 7246
rect 25037 7243 25103 7246
rect 26417 7306 26483 7309
rect 28993 7306 29059 7309
rect 31845 7306 31911 7309
rect 26417 7304 31911 7306
rect 26417 7248 26422 7304
rect 26478 7248 28998 7304
rect 29054 7248 31850 7304
rect 31906 7248 31911 7304
rect 26417 7246 31911 7248
rect 26417 7243 26483 7246
rect 28993 7243 29059 7246
rect 31845 7243 31911 7246
rect 8710 7110 15026 7170
rect 8170 7104 8486 7105
rect 8170 7040 8176 7104
rect 8240 7040 8256 7104
rect 8320 7040 8336 7104
rect 8400 7040 8416 7104
rect 8480 7040 8486 7104
rect 8170 7039 8486 7040
rect 3693 7034 3759 7037
rect 5993 7034 6059 7037
rect 3693 7032 6059 7034
rect 3693 6976 3698 7032
rect 3754 6976 5998 7032
rect 6054 6976 6059 7032
rect 3693 6974 6059 6976
rect 3693 6971 3759 6974
rect 5993 6971 6059 6974
rect 6453 7034 6519 7037
rect 6453 7032 8034 7034
rect 6453 6976 6458 7032
rect 6514 6976 8034 7032
rect 6453 6974 8034 6976
rect 6453 6971 6519 6974
rect 7974 6898 8034 6974
rect 8710 6898 8770 7110
rect 22618 7104 22934 7105
rect 22618 7040 22624 7104
rect 22688 7040 22704 7104
rect 22768 7040 22784 7104
rect 22848 7040 22864 7104
rect 22928 7040 22934 7104
rect 22618 7039 22934 7040
rect 37066 7104 37382 7105
rect 37066 7040 37072 7104
rect 37136 7040 37152 7104
rect 37216 7040 37232 7104
rect 37296 7040 37312 7104
rect 37376 7040 37382 7104
rect 37066 7039 37382 7040
rect 51514 7104 51830 7105
rect 51514 7040 51520 7104
rect 51584 7040 51600 7104
rect 51664 7040 51680 7104
rect 51744 7040 51760 7104
rect 51824 7040 51830 7104
rect 51514 7039 51830 7040
rect 12433 7034 12499 7037
rect 17309 7034 17375 7037
rect 12433 7032 17375 7034
rect 12433 6976 12438 7032
rect 12494 6976 17314 7032
rect 17370 6976 17375 7032
rect 12433 6974 17375 6976
rect 12433 6971 12499 6974
rect 17309 6971 17375 6974
rect 27429 7034 27495 7037
rect 29729 7034 29795 7037
rect 30833 7034 30899 7037
rect 32029 7034 32095 7037
rect 27429 7032 30666 7034
rect 27429 6976 27434 7032
rect 27490 6976 29734 7032
rect 29790 6976 30666 7032
rect 27429 6974 30666 6976
rect 27429 6971 27495 6974
rect 29729 6971 29795 6974
rect 7974 6838 8770 6898
rect 9489 6898 9555 6901
rect 19425 6898 19491 6901
rect 9489 6896 19491 6898
rect 9489 6840 9494 6896
rect 9550 6840 19430 6896
rect 19486 6840 19491 6896
rect 9489 6838 19491 6840
rect 9489 6835 9555 6838
rect 19425 6835 19491 6838
rect 22185 6898 22251 6901
rect 23197 6898 23263 6901
rect 30373 6898 30439 6901
rect 22185 6896 30439 6898
rect 22185 6840 22190 6896
rect 22246 6840 23202 6896
rect 23258 6840 30378 6896
rect 30434 6840 30439 6896
rect 22185 6838 30439 6840
rect 30606 6898 30666 6974
rect 30833 7032 32095 7034
rect 30833 6976 30838 7032
rect 30894 6976 32034 7032
rect 32090 6976 32095 7032
rect 30833 6974 32095 6976
rect 30833 6971 30899 6974
rect 32029 6971 32095 6974
rect 48589 7034 48655 7037
rect 51257 7034 51323 7037
rect 48589 7032 51323 7034
rect 48589 6976 48594 7032
rect 48650 6976 51262 7032
rect 51318 6976 51323 7032
rect 48589 6974 51323 6976
rect 48589 6971 48655 6974
rect 51257 6971 51323 6974
rect 30833 6898 30899 6901
rect 35801 6898 35867 6901
rect 38285 6898 38351 6901
rect 30606 6896 38351 6898
rect 30606 6840 30838 6896
rect 30894 6840 35806 6896
rect 35862 6840 38290 6896
rect 38346 6840 38351 6896
rect 30606 6838 38351 6840
rect 22185 6835 22251 6838
rect 23197 6835 23263 6838
rect 30373 6835 30439 6838
rect 30833 6835 30899 6838
rect 35801 6835 35867 6838
rect 38285 6835 38351 6838
rect 47209 6898 47275 6901
rect 52177 6898 52243 6901
rect 47209 6896 52243 6898
rect 47209 6840 47214 6896
rect 47270 6840 52182 6896
rect 52238 6840 52243 6896
rect 47209 6838 52243 6840
rect 47209 6835 47275 6838
rect 52177 6835 52243 6838
rect 7966 6700 7972 6764
rect 8036 6762 8042 6764
rect 8569 6762 8635 6765
rect 14089 6762 14155 6765
rect 8036 6760 8635 6762
rect 8036 6704 8574 6760
rect 8630 6704 8635 6760
rect 8036 6702 8635 6704
rect 8036 6700 8042 6702
rect 8569 6699 8635 6702
rect 12390 6760 14155 6762
rect 12390 6704 14094 6760
rect 14150 6704 14155 6760
rect 12390 6702 14155 6704
rect 6545 6626 6611 6629
rect 12390 6626 12450 6702
rect 14089 6699 14155 6702
rect 15101 6762 15167 6765
rect 17902 6762 17908 6764
rect 15101 6760 17908 6762
rect 15101 6704 15106 6760
rect 15162 6704 17908 6760
rect 15101 6702 17908 6704
rect 15101 6699 15167 6702
rect 17902 6700 17908 6702
rect 17972 6700 17978 6764
rect 18321 6762 18387 6765
rect 21541 6762 21607 6765
rect 18321 6760 21607 6762
rect 18321 6704 18326 6760
rect 18382 6704 21546 6760
rect 21602 6704 21607 6760
rect 18321 6702 21607 6704
rect 18321 6699 18387 6702
rect 21541 6699 21607 6702
rect 24669 6762 24735 6765
rect 25405 6762 25471 6765
rect 42701 6762 42767 6765
rect 24669 6760 42767 6762
rect 24669 6704 24674 6760
rect 24730 6704 25410 6760
rect 25466 6704 42706 6760
rect 42762 6704 42767 6760
rect 24669 6702 42767 6704
rect 24669 6699 24735 6702
rect 25405 6699 25471 6702
rect 42701 6699 42767 6702
rect 16389 6628 16455 6629
rect 16389 6626 16436 6628
rect 6545 6624 12450 6626
rect 6545 6568 6550 6624
rect 6606 6568 12450 6624
rect 6545 6566 12450 6568
rect 16344 6624 16436 6626
rect 16344 6568 16394 6624
rect 16344 6566 16436 6568
rect 6545 6563 6611 6566
rect 16389 6564 16436 6566
rect 16500 6564 16506 6628
rect 18321 6626 18387 6629
rect 25129 6626 25195 6629
rect 18321 6624 25195 6626
rect 18321 6568 18326 6624
rect 18382 6568 25134 6624
rect 25190 6568 25195 6624
rect 18321 6566 25195 6568
rect 16389 6563 16455 6564
rect 18321 6563 18387 6566
rect 25129 6563 25195 6566
rect 15394 6560 15710 6561
rect 15394 6496 15400 6560
rect 15464 6496 15480 6560
rect 15544 6496 15560 6560
rect 15624 6496 15640 6560
rect 15704 6496 15710 6560
rect 15394 6495 15710 6496
rect 29842 6560 30158 6561
rect 29842 6496 29848 6560
rect 29912 6496 29928 6560
rect 29992 6496 30008 6560
rect 30072 6496 30088 6560
rect 30152 6496 30158 6560
rect 29842 6495 30158 6496
rect 44290 6560 44606 6561
rect 44290 6496 44296 6560
rect 44360 6496 44376 6560
rect 44440 6496 44456 6560
rect 44520 6496 44536 6560
rect 44600 6496 44606 6560
rect 44290 6495 44606 6496
rect 2589 6490 2655 6493
rect 9121 6490 9187 6493
rect 2589 6488 9187 6490
rect 2589 6432 2594 6488
rect 2650 6432 9126 6488
rect 9182 6432 9187 6488
rect 2589 6430 9187 6432
rect 2589 6427 2655 6430
rect 9121 6427 9187 6430
rect 9765 6490 9831 6493
rect 11513 6490 11579 6493
rect 9765 6488 11579 6490
rect 9765 6432 9770 6488
rect 9826 6432 11518 6488
rect 11574 6432 11579 6488
rect 9765 6430 11579 6432
rect 9765 6427 9831 6430
rect 11513 6427 11579 6430
rect 31845 6490 31911 6493
rect 31845 6488 32506 6490
rect 31845 6432 31850 6488
rect 31906 6432 32506 6488
rect 31845 6430 32506 6432
rect 31845 6427 31911 6430
rect 3693 6354 3759 6357
rect 4245 6354 4311 6357
rect 6729 6354 6795 6357
rect 3693 6352 6795 6354
rect 3693 6296 3698 6352
rect 3754 6296 4250 6352
rect 4306 6296 6734 6352
rect 6790 6296 6795 6352
rect 3693 6294 6795 6296
rect 3693 6291 3759 6294
rect 4245 6291 4311 6294
rect 6729 6291 6795 6294
rect 7741 6354 7807 6357
rect 12198 6354 12204 6356
rect 7741 6352 12204 6354
rect 7741 6296 7746 6352
rect 7802 6296 12204 6352
rect 7741 6294 12204 6296
rect 7741 6291 7807 6294
rect 12198 6292 12204 6294
rect 12268 6292 12274 6356
rect 12525 6354 12591 6357
rect 32305 6354 32371 6357
rect 12525 6352 32371 6354
rect 12525 6296 12530 6352
rect 12586 6296 32310 6352
rect 32366 6296 32371 6352
rect 12525 6294 32371 6296
rect 32446 6354 32506 6430
rect 33777 6354 33843 6357
rect 38101 6354 38167 6357
rect 32446 6352 38167 6354
rect 32446 6296 33782 6352
rect 33838 6296 38106 6352
rect 38162 6296 38167 6352
rect 32446 6294 38167 6296
rect 12525 6291 12591 6294
rect 32305 6291 32371 6294
rect 33777 6291 33843 6294
rect 38101 6291 38167 6294
rect 4337 6218 4403 6221
rect 5349 6218 5415 6221
rect 4337 6216 5415 6218
rect 4337 6160 4342 6216
rect 4398 6160 5354 6216
rect 5410 6160 5415 6216
rect 4337 6158 5415 6160
rect 4337 6155 4403 6158
rect 5349 6155 5415 6158
rect 5809 6218 5875 6221
rect 12709 6218 12775 6221
rect 18689 6220 18755 6221
rect 5809 6216 12775 6218
rect 5809 6160 5814 6216
rect 5870 6160 12714 6216
rect 12770 6160 12775 6216
rect 5809 6158 12775 6160
rect 5809 6155 5875 6158
rect 12709 6155 12775 6158
rect 18638 6156 18644 6220
rect 18708 6218 18755 6220
rect 24209 6218 24275 6221
rect 18708 6216 18800 6218
rect 18750 6160 18800 6216
rect 18708 6158 18800 6160
rect 22050 6216 24275 6218
rect 22050 6160 24214 6216
rect 24270 6160 24275 6216
rect 22050 6158 24275 6160
rect 18708 6156 18755 6158
rect 18689 6155 18755 6156
rect 9765 6082 9831 6085
rect 9990 6082 9996 6084
rect 9765 6080 9996 6082
rect 9765 6024 9770 6080
rect 9826 6024 9996 6080
rect 9765 6022 9996 6024
rect 9765 6019 9831 6022
rect 9990 6020 9996 6022
rect 10060 6020 10066 6084
rect 10225 6082 10291 6085
rect 10869 6082 10935 6085
rect 10225 6080 10935 6082
rect 10225 6024 10230 6080
rect 10286 6024 10874 6080
rect 10930 6024 10935 6080
rect 10225 6022 10935 6024
rect 10225 6019 10291 6022
rect 10869 6019 10935 6022
rect 11881 6082 11947 6085
rect 17861 6082 17927 6085
rect 11881 6080 17927 6082
rect 11881 6024 11886 6080
rect 11942 6024 17866 6080
rect 17922 6024 17927 6080
rect 11881 6022 17927 6024
rect 11881 6019 11947 6022
rect 17861 6019 17927 6022
rect 8170 6016 8486 6017
rect 8170 5952 8176 6016
rect 8240 5952 8256 6016
rect 8320 5952 8336 6016
rect 8400 5952 8416 6016
rect 8480 5952 8486 6016
rect 8170 5951 8486 5952
rect 8661 5946 8727 5949
rect 17493 5946 17559 5949
rect 22050 5946 22110 6158
rect 24209 6155 24275 6158
rect 24761 6218 24827 6221
rect 25497 6218 25563 6221
rect 24761 6216 25563 6218
rect 24761 6160 24766 6216
rect 24822 6160 25502 6216
rect 25558 6160 25563 6216
rect 24761 6158 25563 6160
rect 24761 6155 24827 6158
rect 25497 6155 25563 6158
rect 27429 6218 27495 6221
rect 37089 6218 37155 6221
rect 27429 6216 37155 6218
rect 27429 6160 27434 6216
rect 27490 6160 37094 6216
rect 37150 6160 37155 6216
rect 27429 6158 37155 6160
rect 27429 6155 27495 6158
rect 37089 6155 37155 6158
rect 37917 6218 37983 6221
rect 45829 6218 45895 6221
rect 37917 6216 45895 6218
rect 37917 6160 37922 6216
rect 37978 6160 45834 6216
rect 45890 6160 45895 6216
rect 37917 6158 45895 6160
rect 37917 6155 37983 6158
rect 45829 6155 45895 6158
rect 24393 6082 24459 6085
rect 32581 6082 32647 6085
rect 24393 6080 32647 6082
rect 24393 6024 24398 6080
rect 24454 6024 32586 6080
rect 32642 6024 32647 6080
rect 24393 6022 32647 6024
rect 24393 6019 24459 6022
rect 32581 6019 32647 6022
rect 22618 6016 22934 6017
rect 22618 5952 22624 6016
rect 22688 5952 22704 6016
rect 22768 5952 22784 6016
rect 22848 5952 22864 6016
rect 22928 5952 22934 6016
rect 22618 5951 22934 5952
rect 37066 6016 37382 6017
rect 37066 5952 37072 6016
rect 37136 5952 37152 6016
rect 37216 5952 37232 6016
rect 37296 5952 37312 6016
rect 37376 5952 37382 6016
rect 37066 5951 37382 5952
rect 51514 6016 51830 6017
rect 51514 5952 51520 6016
rect 51584 5952 51600 6016
rect 51664 5952 51680 6016
rect 51744 5952 51760 6016
rect 51824 5952 51830 6016
rect 51514 5951 51830 5952
rect 8661 5944 22110 5946
rect 8661 5888 8666 5944
rect 8722 5888 17498 5944
rect 17554 5888 22110 5944
rect 8661 5886 22110 5888
rect 28993 5946 29059 5949
rect 33685 5946 33751 5949
rect 28993 5944 33751 5946
rect 28993 5888 28998 5944
rect 29054 5888 33690 5944
rect 33746 5888 33751 5944
rect 28993 5886 33751 5888
rect 8661 5883 8727 5886
rect 17493 5883 17559 5886
rect 28993 5883 29059 5886
rect 33685 5883 33751 5886
rect 42977 5946 43043 5949
rect 50797 5946 50863 5949
rect 42977 5944 50863 5946
rect 42977 5888 42982 5944
rect 43038 5888 50802 5944
rect 50858 5888 50863 5944
rect 42977 5886 50863 5888
rect 42977 5883 43043 5886
rect 50797 5883 50863 5886
rect 3417 5810 3483 5813
rect 6361 5810 6427 5813
rect 3417 5808 6427 5810
rect 3417 5752 3422 5808
rect 3478 5752 6366 5808
rect 6422 5752 6427 5808
rect 3417 5750 6427 5752
rect 3417 5747 3483 5750
rect 6361 5747 6427 5750
rect 7281 5810 7347 5813
rect 7741 5810 7807 5813
rect 7281 5808 7807 5810
rect 7281 5752 7286 5808
rect 7342 5752 7746 5808
rect 7802 5752 7807 5808
rect 7281 5750 7807 5752
rect 7281 5747 7347 5750
rect 7741 5747 7807 5750
rect 8201 5810 8267 5813
rect 10225 5810 10291 5813
rect 29729 5810 29795 5813
rect 8201 5808 10291 5810
rect 8201 5752 8206 5808
rect 8262 5752 10230 5808
rect 10286 5752 10291 5808
rect 8201 5750 10291 5752
rect 8201 5747 8267 5750
rect 10225 5747 10291 5750
rect 22050 5808 29795 5810
rect 22050 5752 29734 5808
rect 29790 5752 29795 5808
rect 22050 5750 29795 5752
rect 3049 5674 3115 5677
rect 6637 5674 6703 5677
rect 3049 5672 6703 5674
rect 3049 5616 3054 5672
rect 3110 5616 6642 5672
rect 6698 5616 6703 5672
rect 3049 5614 6703 5616
rect 3049 5611 3115 5614
rect 6637 5611 6703 5614
rect 7649 5674 7715 5677
rect 10317 5674 10383 5677
rect 12198 5674 12204 5676
rect 7649 5672 9690 5674
rect 7649 5616 7654 5672
rect 7710 5616 9690 5672
rect 7649 5614 9690 5616
rect 7649 5611 7715 5614
rect 9630 5538 9690 5614
rect 10317 5672 12204 5674
rect 10317 5616 10322 5672
rect 10378 5616 12204 5672
rect 10317 5614 12204 5616
rect 10317 5611 10383 5614
rect 12198 5612 12204 5614
rect 12268 5612 12274 5676
rect 12382 5612 12388 5676
rect 12452 5674 12458 5676
rect 22050 5674 22110 5750
rect 29729 5747 29795 5750
rect 45645 5810 45711 5813
rect 53097 5810 53163 5813
rect 45645 5808 53163 5810
rect 45645 5752 45650 5808
rect 45706 5752 53102 5808
rect 53158 5752 53163 5808
rect 45645 5750 53163 5752
rect 45645 5747 45711 5750
rect 53097 5747 53163 5750
rect 12452 5614 22110 5674
rect 12452 5612 12458 5614
rect 22318 5612 22324 5676
rect 22388 5674 22394 5676
rect 23197 5674 23263 5677
rect 22388 5672 23263 5674
rect 22388 5616 23202 5672
rect 23258 5616 23263 5672
rect 22388 5614 23263 5616
rect 22388 5612 22394 5614
rect 23197 5611 23263 5614
rect 23606 5612 23612 5676
rect 23676 5674 23682 5676
rect 30373 5674 30439 5677
rect 23676 5672 30439 5674
rect 23676 5616 30378 5672
rect 30434 5616 30439 5672
rect 23676 5614 30439 5616
rect 23676 5612 23682 5614
rect 30373 5611 30439 5614
rect 36353 5674 36419 5677
rect 40401 5674 40467 5677
rect 36353 5672 40467 5674
rect 36353 5616 36358 5672
rect 36414 5616 40406 5672
rect 40462 5616 40467 5672
rect 36353 5614 40467 5616
rect 36353 5611 36419 5614
rect 40401 5611 40467 5614
rect 14917 5538 14983 5541
rect 9630 5536 14983 5538
rect 9630 5480 14922 5536
rect 14978 5480 14983 5536
rect 9630 5478 14983 5480
rect 14917 5475 14983 5478
rect 17125 5538 17191 5541
rect 23749 5538 23815 5541
rect 17125 5536 23815 5538
rect 17125 5480 17130 5536
rect 17186 5480 23754 5536
rect 23810 5480 23815 5536
rect 17125 5478 23815 5480
rect 17125 5475 17191 5478
rect 23749 5475 23815 5478
rect 15394 5472 15710 5473
rect 15394 5408 15400 5472
rect 15464 5408 15480 5472
rect 15544 5408 15560 5472
rect 15624 5408 15640 5472
rect 15704 5408 15710 5472
rect 15394 5407 15710 5408
rect 29842 5472 30158 5473
rect 29842 5408 29848 5472
rect 29912 5408 29928 5472
rect 29992 5408 30008 5472
rect 30072 5408 30088 5472
rect 30152 5408 30158 5472
rect 29842 5407 30158 5408
rect 44290 5472 44606 5473
rect 44290 5408 44296 5472
rect 44360 5408 44376 5472
rect 44440 5408 44456 5472
rect 44520 5408 44536 5472
rect 44600 5408 44606 5472
rect 44290 5407 44606 5408
rect 2681 5402 2747 5405
rect 2814 5402 2820 5404
rect 2681 5400 2820 5402
rect 2681 5344 2686 5400
rect 2742 5344 2820 5400
rect 2681 5342 2820 5344
rect 2681 5339 2747 5342
rect 2814 5340 2820 5342
rect 2884 5402 2890 5404
rect 6177 5402 6243 5405
rect 2884 5400 6243 5402
rect 2884 5344 6182 5400
rect 6238 5344 6243 5400
rect 2884 5342 6243 5344
rect 2884 5340 2890 5342
rect 6177 5339 6243 5342
rect 9489 5402 9555 5405
rect 9673 5402 9739 5405
rect 9489 5400 9739 5402
rect 9489 5344 9494 5400
rect 9550 5344 9678 5400
rect 9734 5344 9739 5400
rect 9489 5342 9739 5344
rect 9489 5339 9555 5342
rect 9673 5339 9739 5342
rect 19333 5402 19399 5405
rect 26969 5402 27035 5405
rect 19333 5400 27035 5402
rect 19333 5344 19338 5400
rect 19394 5344 26974 5400
rect 27030 5344 27035 5400
rect 19333 5342 27035 5344
rect 19333 5339 19399 5342
rect 26969 5339 27035 5342
rect 31937 5402 32003 5405
rect 42793 5402 42859 5405
rect 31937 5400 42859 5402
rect 31937 5344 31942 5400
rect 31998 5344 42798 5400
rect 42854 5344 42859 5400
rect 31937 5342 42859 5344
rect 31937 5339 32003 5342
rect 42793 5339 42859 5342
rect 1894 5204 1900 5268
rect 1964 5266 1970 5268
rect 13486 5266 13492 5268
rect 1964 5206 13492 5266
rect 1964 5204 1970 5206
rect 13486 5204 13492 5206
rect 13556 5204 13562 5268
rect 24761 5266 24827 5269
rect 26877 5266 26943 5269
rect 24761 5264 26943 5266
rect 24761 5208 24766 5264
rect 24822 5208 26882 5264
rect 26938 5208 26943 5264
rect 24761 5206 26943 5208
rect 24761 5203 24827 5206
rect 26877 5203 26943 5206
rect 34145 5266 34211 5269
rect 45461 5266 45527 5269
rect 34145 5264 45527 5266
rect 34145 5208 34150 5264
rect 34206 5208 45466 5264
rect 45522 5208 45527 5264
rect 34145 5206 45527 5208
rect 34145 5203 34211 5206
rect 45461 5203 45527 5206
rect 2129 5130 2195 5133
rect 5809 5130 5875 5133
rect 10041 5130 10107 5133
rect 2129 5128 5875 5130
rect 2129 5072 2134 5128
rect 2190 5072 5814 5128
rect 5870 5072 5875 5128
rect 2129 5070 5875 5072
rect 2129 5067 2195 5070
rect 5809 5067 5875 5070
rect 7974 5128 10107 5130
rect 7974 5072 10046 5128
rect 10102 5072 10107 5128
rect 7974 5070 10107 5072
rect 5717 4994 5783 4997
rect 7974 4994 8034 5070
rect 10041 5067 10107 5070
rect 12157 5130 12223 5133
rect 13813 5130 13879 5133
rect 12157 5128 13879 5130
rect 12157 5072 12162 5128
rect 12218 5072 13818 5128
rect 13874 5072 13879 5128
rect 12157 5070 13879 5072
rect 12157 5067 12223 5070
rect 13813 5067 13879 5070
rect 16430 5068 16436 5132
rect 16500 5130 16506 5132
rect 18689 5130 18755 5133
rect 16500 5128 18755 5130
rect 16500 5072 18694 5128
rect 18750 5072 18755 5128
rect 16500 5070 18755 5072
rect 16500 5068 16506 5070
rect 18689 5067 18755 5070
rect 19149 5130 19215 5133
rect 25589 5130 25655 5133
rect 19149 5128 25655 5130
rect 19149 5072 19154 5128
rect 19210 5072 25594 5128
rect 25650 5072 25655 5128
rect 19149 5070 25655 5072
rect 19149 5067 19215 5070
rect 25589 5067 25655 5070
rect 28901 5130 28967 5133
rect 40217 5130 40283 5133
rect 28901 5128 40283 5130
rect 28901 5072 28906 5128
rect 28962 5072 40222 5128
rect 40278 5072 40283 5128
rect 28901 5070 40283 5072
rect 28901 5067 28967 5070
rect 40217 5067 40283 5070
rect 43161 5130 43227 5133
rect 51073 5130 51139 5133
rect 43161 5128 51139 5130
rect 43161 5072 43166 5128
rect 43222 5072 51078 5128
rect 51134 5072 51139 5128
rect 43161 5070 51139 5072
rect 43161 5067 43227 5070
rect 51073 5067 51139 5070
rect 5717 4992 8034 4994
rect 5717 4936 5722 4992
rect 5778 4936 8034 4992
rect 5717 4934 8034 4936
rect 9857 4994 9923 4997
rect 11513 4994 11579 4997
rect 9857 4992 11579 4994
rect 9857 4936 9862 4992
rect 9918 4936 11518 4992
rect 11574 4936 11579 4992
rect 9857 4934 11579 4936
rect 5717 4931 5783 4934
rect 9857 4931 9923 4934
rect 11513 4931 11579 4934
rect 16941 4994 17007 4997
rect 19333 4994 19399 4997
rect 29637 4994 29703 4997
rect 34513 4994 34579 4997
rect 16941 4992 19399 4994
rect 16941 4936 16946 4992
rect 17002 4936 19338 4992
rect 19394 4936 19399 4992
rect 16941 4934 19399 4936
rect 16941 4931 17007 4934
rect 19333 4931 19399 4934
rect 23016 4992 34579 4994
rect 23016 4936 29642 4992
rect 29698 4936 34518 4992
rect 34574 4936 34579 4992
rect 23016 4934 34579 4936
rect 8170 4928 8486 4929
rect 8170 4864 8176 4928
rect 8240 4864 8256 4928
rect 8320 4864 8336 4928
rect 8400 4864 8416 4928
rect 8480 4864 8486 4928
rect 8170 4863 8486 4864
rect 22618 4928 22934 4929
rect 22618 4864 22624 4928
rect 22688 4864 22704 4928
rect 22768 4864 22784 4928
rect 22848 4864 22864 4928
rect 22928 4864 22934 4928
rect 22618 4863 22934 4864
rect 1577 4858 1643 4861
rect 6913 4858 6979 4861
rect 1577 4856 6979 4858
rect 1577 4800 1582 4856
rect 1638 4800 6918 4856
rect 6974 4800 6979 4856
rect 1577 4798 6979 4800
rect 1577 4795 1643 4798
rect 6913 4795 6979 4798
rect 8661 4858 8727 4861
rect 8886 4858 8892 4860
rect 8661 4856 8892 4858
rect 8661 4800 8666 4856
rect 8722 4800 8892 4856
rect 8661 4798 8892 4800
rect 8661 4795 8727 4798
rect 8886 4796 8892 4798
rect 8956 4796 8962 4860
rect 10041 4858 10107 4861
rect 10726 4858 10732 4860
rect 10041 4856 10732 4858
rect 10041 4800 10046 4856
rect 10102 4800 10732 4856
rect 10041 4798 10732 4800
rect 10041 4795 10107 4798
rect 10726 4796 10732 4798
rect 10796 4858 10802 4860
rect 14181 4858 14247 4861
rect 10796 4856 14247 4858
rect 10796 4800 14186 4856
rect 14242 4800 14247 4856
rect 10796 4798 14247 4800
rect 10796 4796 10802 4798
rect 14181 4795 14247 4798
rect 14825 4858 14891 4861
rect 17953 4858 18019 4861
rect 14825 4856 18019 4858
rect 14825 4800 14830 4856
rect 14886 4800 17958 4856
rect 18014 4800 18019 4856
rect 14825 4798 18019 4800
rect 14825 4795 14891 4798
rect 17953 4795 18019 4798
rect 18689 4858 18755 4861
rect 21725 4858 21791 4861
rect 18689 4856 21791 4858
rect 18689 4800 18694 4856
rect 18750 4800 21730 4856
rect 21786 4800 21791 4856
rect 18689 4798 21791 4800
rect 18689 4795 18755 4798
rect 21725 4795 21791 4798
rect 2497 4722 2563 4725
rect 5717 4722 5783 4725
rect 2497 4720 5783 4722
rect 2497 4664 2502 4720
rect 2558 4664 5722 4720
rect 5778 4664 5783 4720
rect 2497 4662 5783 4664
rect 2497 4659 2563 4662
rect 5717 4659 5783 4662
rect 6177 4722 6243 4725
rect 14365 4722 14431 4725
rect 14774 4722 14780 4724
rect 6177 4720 12450 4722
rect 6177 4664 6182 4720
rect 6238 4664 12450 4720
rect 6177 4662 12450 4664
rect 6177 4659 6243 4662
rect 6269 4586 6335 4589
rect 10317 4586 10383 4589
rect 6269 4584 10383 4586
rect 6269 4528 6274 4584
rect 6330 4528 10322 4584
rect 10378 4528 10383 4584
rect 6269 4526 10383 4528
rect 12390 4586 12450 4662
rect 14365 4720 14780 4722
rect 14365 4664 14370 4720
rect 14426 4664 14780 4720
rect 14365 4662 14780 4664
rect 14365 4659 14431 4662
rect 14774 4660 14780 4662
rect 14844 4722 14850 4724
rect 17585 4722 17651 4725
rect 14844 4720 17651 4722
rect 14844 4664 17590 4720
rect 17646 4664 17651 4720
rect 14844 4662 17651 4664
rect 17956 4722 18016 4795
rect 22134 4722 22140 4724
rect 17956 4662 22140 4722
rect 14844 4660 14850 4662
rect 17585 4659 17651 4662
rect 22134 4660 22140 4662
rect 22204 4722 22210 4724
rect 22553 4722 22619 4725
rect 23016 4722 23076 4934
rect 29637 4931 29703 4934
rect 34513 4931 34579 4934
rect 37066 4928 37382 4929
rect 37066 4864 37072 4928
rect 37136 4864 37152 4928
rect 37216 4864 37232 4928
rect 37296 4864 37312 4928
rect 37376 4864 37382 4928
rect 37066 4863 37382 4864
rect 51514 4928 51830 4929
rect 51514 4864 51520 4928
rect 51584 4864 51600 4928
rect 51664 4864 51680 4928
rect 51744 4864 51760 4928
rect 51824 4864 51830 4928
rect 51514 4863 51830 4864
rect 24485 4858 24551 4861
rect 31017 4858 31083 4861
rect 24485 4856 31083 4858
rect 24485 4800 24490 4856
rect 24546 4800 31022 4856
rect 31078 4800 31083 4856
rect 24485 4798 31083 4800
rect 24485 4795 24551 4798
rect 31017 4795 31083 4798
rect 40401 4858 40467 4861
rect 46197 4858 46263 4861
rect 40401 4856 46263 4858
rect 40401 4800 40406 4856
rect 40462 4800 46202 4856
rect 46258 4800 46263 4856
rect 40401 4798 46263 4800
rect 40401 4795 40467 4798
rect 46197 4795 46263 4798
rect 22204 4720 23076 4722
rect 22204 4664 22558 4720
rect 22614 4664 23076 4720
rect 22204 4662 23076 4664
rect 25681 4722 25747 4725
rect 31569 4722 31635 4725
rect 25681 4720 31635 4722
rect 25681 4664 25686 4720
rect 25742 4664 31574 4720
rect 31630 4664 31635 4720
rect 25681 4662 31635 4664
rect 22204 4660 22210 4662
rect 22553 4659 22619 4662
rect 25681 4659 25747 4662
rect 31569 4659 31635 4662
rect 39021 4722 39087 4725
rect 41321 4722 41387 4725
rect 39021 4720 41387 4722
rect 39021 4664 39026 4720
rect 39082 4664 41326 4720
rect 41382 4664 41387 4720
rect 39021 4662 41387 4664
rect 39021 4659 39087 4662
rect 41321 4659 41387 4662
rect 43621 4722 43687 4725
rect 48405 4722 48471 4725
rect 43621 4720 48471 4722
rect 43621 4664 43626 4720
rect 43682 4664 48410 4720
rect 48466 4664 48471 4720
rect 43621 4662 48471 4664
rect 43621 4659 43687 4662
rect 48405 4659 48471 4662
rect 53557 4586 53623 4589
rect 12390 4584 53623 4586
rect 12390 4528 53562 4584
rect 53618 4528 53623 4584
rect 12390 4526 53623 4528
rect 6269 4523 6335 4526
rect 10317 4523 10383 4526
rect 53557 4523 53623 4526
rect 4889 4450 4955 4453
rect 7741 4450 7807 4453
rect 4889 4448 7807 4450
rect 4889 4392 4894 4448
rect 4950 4392 7746 4448
rect 7802 4392 7807 4448
rect 4889 4390 7807 4392
rect 4889 4387 4955 4390
rect 7741 4387 7807 4390
rect 8569 4450 8635 4453
rect 9070 4450 9076 4452
rect 8569 4448 9076 4450
rect 8569 4392 8574 4448
rect 8630 4392 9076 4448
rect 8569 4390 9076 4392
rect 8569 4387 8635 4390
rect 9070 4388 9076 4390
rect 9140 4388 9146 4452
rect 18137 4450 18203 4453
rect 23933 4450 23999 4453
rect 18137 4448 23999 4450
rect 18137 4392 18142 4448
rect 18198 4392 23938 4448
rect 23994 4392 23999 4448
rect 18137 4390 23999 4392
rect 18137 4387 18203 4390
rect 23933 4387 23999 4390
rect 24209 4450 24275 4453
rect 25773 4450 25839 4453
rect 24209 4448 25839 4450
rect 24209 4392 24214 4448
rect 24270 4392 25778 4448
rect 25834 4392 25839 4448
rect 24209 4390 25839 4392
rect 24209 4387 24275 4390
rect 25773 4387 25839 4390
rect 35801 4450 35867 4453
rect 42701 4450 42767 4453
rect 35801 4448 42767 4450
rect 35801 4392 35806 4448
rect 35862 4392 42706 4448
rect 42762 4392 42767 4448
rect 35801 4390 42767 4392
rect 35801 4387 35867 4390
rect 42701 4387 42767 4390
rect 44817 4450 44883 4453
rect 48497 4450 48563 4453
rect 44817 4448 48563 4450
rect 44817 4392 44822 4448
rect 44878 4392 48502 4448
rect 48558 4392 48563 4448
rect 44817 4390 48563 4392
rect 44817 4387 44883 4390
rect 48497 4387 48563 4390
rect 15394 4384 15710 4385
rect 15394 4320 15400 4384
rect 15464 4320 15480 4384
rect 15544 4320 15560 4384
rect 15624 4320 15640 4384
rect 15704 4320 15710 4384
rect 15394 4319 15710 4320
rect 29842 4384 30158 4385
rect 29842 4320 29848 4384
rect 29912 4320 29928 4384
rect 29992 4320 30008 4384
rect 30072 4320 30088 4384
rect 30152 4320 30158 4384
rect 29842 4319 30158 4320
rect 44290 4384 44606 4385
rect 44290 4320 44296 4384
rect 44360 4320 44376 4384
rect 44440 4320 44456 4384
rect 44520 4320 44536 4384
rect 44600 4320 44606 4384
rect 44290 4319 44606 4320
rect 1761 4314 1827 4317
rect 1894 4314 1900 4316
rect 1761 4312 1900 4314
rect 1761 4256 1766 4312
rect 1822 4256 1900 4312
rect 1761 4254 1900 4256
rect 1761 4251 1827 4254
rect 1894 4252 1900 4254
rect 1964 4252 1970 4316
rect 3785 4314 3851 4317
rect 8886 4314 8892 4316
rect 3785 4312 8892 4314
rect 3785 4256 3790 4312
rect 3846 4256 8892 4312
rect 3785 4254 8892 4256
rect 3785 4251 3851 4254
rect 8886 4252 8892 4254
rect 8956 4252 8962 4316
rect 16757 4314 16823 4317
rect 16982 4314 16988 4316
rect 16757 4312 16988 4314
rect 16757 4256 16762 4312
rect 16818 4256 16988 4312
rect 16757 4254 16988 4256
rect 16757 4251 16823 4254
rect 16982 4252 16988 4254
rect 17052 4252 17058 4316
rect 21265 4314 21331 4317
rect 26509 4314 26575 4317
rect 21265 4312 26575 4314
rect 21265 4256 21270 4312
rect 21326 4256 26514 4312
rect 26570 4256 26575 4312
rect 21265 4254 26575 4256
rect 21265 4251 21331 4254
rect 26509 4251 26575 4254
rect 38101 4314 38167 4317
rect 44081 4314 44147 4317
rect 38101 4312 44147 4314
rect 38101 4256 38106 4312
rect 38162 4256 44086 4312
rect 44142 4256 44147 4312
rect 38101 4254 44147 4256
rect 38101 4251 38167 4254
rect 44081 4251 44147 4254
rect 1853 4178 1919 4181
rect 6545 4178 6611 4181
rect 1853 4176 6611 4178
rect 1853 4120 1858 4176
rect 1914 4120 6550 4176
rect 6606 4120 6611 4176
rect 1853 4118 6611 4120
rect 1853 4115 1919 4118
rect 6545 4115 6611 4118
rect 7465 4178 7531 4181
rect 7598 4178 7604 4180
rect 7465 4176 7604 4178
rect 7465 4120 7470 4176
rect 7526 4120 7604 4176
rect 7465 4118 7604 4120
rect 7465 4115 7531 4118
rect 7598 4116 7604 4118
rect 7668 4116 7674 4180
rect 14825 4178 14891 4181
rect 18137 4178 18203 4181
rect 14825 4176 18203 4178
rect 14825 4120 14830 4176
rect 14886 4120 18142 4176
rect 18198 4120 18203 4176
rect 14825 4118 18203 4120
rect 14825 4115 14891 4118
rect 18137 4115 18203 4118
rect 19057 4178 19123 4181
rect 23013 4178 23079 4181
rect 19057 4176 23079 4178
rect 19057 4120 19062 4176
rect 19118 4120 23018 4176
rect 23074 4120 23079 4176
rect 19057 4118 23079 4120
rect 19057 4115 19123 4118
rect 23013 4115 23079 4118
rect 25221 4178 25287 4181
rect 29177 4178 29243 4181
rect 25221 4176 29243 4178
rect 25221 4120 25226 4176
rect 25282 4120 29182 4176
rect 29238 4120 29243 4176
rect 25221 4118 29243 4120
rect 25221 4115 25287 4118
rect 29177 4115 29243 4118
rect 30097 4178 30163 4181
rect 34145 4178 34211 4181
rect 30097 4176 34211 4178
rect 30097 4120 30102 4176
rect 30158 4120 34150 4176
rect 34206 4120 34211 4176
rect 30097 4118 34211 4120
rect 30097 4115 30163 4118
rect 34145 4115 34211 4118
rect 39941 4178 40007 4181
rect 52085 4178 52151 4181
rect 39941 4176 52151 4178
rect 39941 4120 39946 4176
rect 40002 4120 52090 4176
rect 52146 4120 52151 4176
rect 39941 4118 52151 4120
rect 39941 4115 40007 4118
rect 52085 4115 52151 4118
rect 5809 4042 5875 4045
rect 13169 4042 13235 4045
rect 13302 4042 13308 4044
rect 5809 4040 12450 4042
rect 5809 3984 5814 4040
rect 5870 3984 12450 4040
rect 5809 3982 12450 3984
rect 5809 3979 5875 3982
rect 6637 3908 6703 3909
rect 8661 3908 8727 3909
rect 6637 3906 6684 3908
rect 6592 3904 6684 3906
rect 6592 3848 6642 3904
rect 6592 3846 6684 3848
rect 6637 3844 6684 3846
rect 6748 3844 6754 3908
rect 8661 3906 8708 3908
rect 8616 3904 8708 3906
rect 8616 3848 8666 3904
rect 8616 3846 8708 3848
rect 8661 3844 8708 3846
rect 8772 3844 8778 3908
rect 12390 3906 12450 3982
rect 13169 4040 13308 4042
rect 13169 3984 13174 4040
rect 13230 3984 13308 4040
rect 13169 3982 13308 3984
rect 13169 3979 13235 3982
rect 13302 3980 13308 3982
rect 13372 3980 13378 4044
rect 14365 4042 14431 4045
rect 14590 4042 14596 4044
rect 14365 4040 14596 4042
rect 14365 3984 14370 4040
rect 14426 3984 14596 4040
rect 14365 3982 14596 3984
rect 14365 3979 14431 3982
rect 14590 3980 14596 3982
rect 14660 3980 14666 4044
rect 14917 4042 14983 4045
rect 19149 4044 19215 4045
rect 19149 4042 19196 4044
rect 14917 4040 19196 4042
rect 14917 3984 14922 4040
rect 14978 3984 19154 4040
rect 14917 3982 19196 3984
rect 14917 3979 14983 3982
rect 19149 3980 19196 3982
rect 19260 3980 19266 4044
rect 43529 4042 43595 4045
rect 44449 4042 44515 4045
rect 46749 4042 46815 4045
rect 22050 4040 46815 4042
rect 22050 3984 43534 4040
rect 43590 3984 44454 4040
rect 44510 3984 46754 4040
rect 46810 3984 46815 4040
rect 22050 3982 46815 3984
rect 19149 3979 19215 3980
rect 22050 3906 22110 3982
rect 43529 3979 43595 3982
rect 44449 3979 44515 3982
rect 46749 3979 46815 3982
rect 51809 4042 51875 4045
rect 52453 4042 52519 4045
rect 55213 4042 55279 4045
rect 51809 4040 55279 4042
rect 51809 3984 51814 4040
rect 51870 3984 52458 4040
rect 52514 3984 55218 4040
rect 55274 3984 55279 4040
rect 51809 3982 55279 3984
rect 51809 3979 51875 3982
rect 52453 3979 52519 3982
rect 55213 3979 55279 3982
rect 12390 3846 22110 3906
rect 23013 3908 23079 3909
rect 23013 3904 23060 3908
rect 23124 3906 23130 3908
rect 24577 3906 24643 3909
rect 30557 3906 30623 3909
rect 35709 3908 35775 3909
rect 35709 3906 35756 3908
rect 23013 3848 23018 3904
rect 23013 3844 23060 3848
rect 23124 3846 23170 3906
rect 24577 3904 30623 3906
rect 24577 3848 24582 3904
rect 24638 3848 30562 3904
rect 30618 3848 30623 3904
rect 24577 3846 30623 3848
rect 35664 3904 35756 3906
rect 35664 3848 35714 3904
rect 35664 3846 35756 3848
rect 23124 3844 23130 3846
rect 6637 3843 6703 3844
rect 8661 3843 8727 3844
rect 23013 3843 23079 3844
rect 24577 3843 24643 3846
rect 30557 3843 30623 3846
rect 35709 3844 35756 3846
rect 35820 3844 35826 3908
rect 39113 3906 39179 3909
rect 42425 3906 42491 3909
rect 46565 3906 46631 3909
rect 39113 3904 46631 3906
rect 39113 3848 39118 3904
rect 39174 3848 42430 3904
rect 42486 3848 46570 3904
rect 46626 3848 46631 3904
rect 39113 3846 46631 3848
rect 35709 3843 35775 3844
rect 39113 3843 39179 3846
rect 42425 3843 42491 3846
rect 46565 3843 46631 3846
rect 8170 3840 8486 3841
rect 8170 3776 8176 3840
rect 8240 3776 8256 3840
rect 8320 3776 8336 3840
rect 8400 3776 8416 3840
rect 8480 3776 8486 3840
rect 8170 3775 8486 3776
rect 22618 3840 22934 3841
rect 22618 3776 22624 3840
rect 22688 3776 22704 3840
rect 22768 3776 22784 3840
rect 22848 3776 22864 3840
rect 22928 3776 22934 3840
rect 22618 3775 22934 3776
rect 37066 3840 37382 3841
rect 37066 3776 37072 3840
rect 37136 3776 37152 3840
rect 37216 3776 37232 3840
rect 37296 3776 37312 3840
rect 37376 3776 37382 3840
rect 37066 3775 37382 3776
rect 51514 3840 51830 3841
rect 51514 3776 51520 3840
rect 51584 3776 51600 3840
rect 51664 3776 51680 3840
rect 51744 3776 51760 3840
rect 51824 3776 51830 3840
rect 51514 3775 51830 3776
rect 7465 3772 7531 3773
rect 7414 3770 7420 3772
rect 7374 3710 7420 3770
rect 7484 3768 7531 3772
rect 7526 3712 7531 3768
rect 7414 3708 7420 3710
rect 7484 3708 7531 3712
rect 7465 3707 7531 3708
rect 8937 3770 9003 3773
rect 9438 3770 9444 3772
rect 8937 3768 9444 3770
rect 8937 3712 8942 3768
rect 8998 3712 9444 3768
rect 8937 3710 9444 3712
rect 8937 3707 9003 3710
rect 9438 3708 9444 3710
rect 9508 3708 9514 3772
rect 15377 3770 15443 3773
rect 16430 3770 16436 3772
rect 15377 3768 16436 3770
rect 15377 3712 15382 3768
rect 15438 3712 16436 3768
rect 15377 3710 16436 3712
rect 15377 3707 15443 3710
rect 16430 3708 16436 3710
rect 16500 3708 16506 3772
rect 16614 3708 16620 3772
rect 16684 3770 16690 3772
rect 16757 3770 16823 3773
rect 16684 3768 16823 3770
rect 16684 3712 16762 3768
rect 16818 3712 16823 3768
rect 16684 3710 16823 3712
rect 16684 3708 16690 3710
rect 16757 3707 16823 3710
rect 37457 3770 37523 3773
rect 47577 3770 47643 3773
rect 37457 3768 47643 3770
rect 37457 3712 37462 3768
rect 37518 3712 47582 3768
rect 47638 3712 47643 3768
rect 37457 3710 47643 3712
rect 37457 3707 37523 3710
rect 47577 3707 47643 3710
rect 6821 3634 6887 3637
rect 12157 3634 12223 3637
rect 14825 3636 14891 3637
rect 18321 3636 18387 3637
rect 6821 3632 12223 3634
rect 6821 3576 6826 3632
rect 6882 3576 12162 3632
rect 12218 3576 12223 3632
rect 6821 3574 12223 3576
rect 6821 3571 6887 3574
rect 12157 3571 12223 3574
rect 14774 3572 14780 3636
rect 14844 3634 14891 3636
rect 14844 3632 14936 3634
rect 14886 3576 14936 3632
rect 14844 3574 14936 3576
rect 14844 3572 14891 3574
rect 18270 3572 18276 3636
rect 18340 3634 18387 3636
rect 23381 3636 23447 3637
rect 23381 3634 23428 3636
rect 18340 3632 18432 3634
rect 18382 3576 18432 3632
rect 18340 3574 18432 3576
rect 23336 3632 23428 3634
rect 23336 3576 23386 3632
rect 23336 3574 23428 3576
rect 18340 3572 18387 3574
rect 14825 3571 14891 3572
rect 18321 3571 18387 3572
rect 23381 3572 23428 3574
rect 23492 3572 23498 3636
rect 34881 3634 34947 3637
rect 40677 3634 40743 3637
rect 34881 3632 40743 3634
rect 34881 3576 34886 3632
rect 34942 3576 40682 3632
rect 40738 3576 40743 3632
rect 34881 3574 40743 3576
rect 23381 3571 23447 3572
rect 34881 3571 34947 3574
rect 40677 3571 40743 3574
rect 4245 3498 4311 3501
rect 10501 3498 10567 3501
rect 4245 3496 10567 3498
rect 4245 3440 4250 3496
rect 4306 3440 10506 3496
rect 10562 3440 10567 3496
rect 4245 3438 10567 3440
rect 4245 3435 4311 3438
rect 10501 3435 10567 3438
rect 14457 3498 14523 3501
rect 17217 3498 17283 3501
rect 38285 3498 38351 3501
rect 14457 3496 15946 3498
rect 14457 3440 14462 3496
rect 14518 3440 15946 3496
rect 14457 3438 15946 3440
rect 14457 3435 14523 3438
rect 5441 3362 5507 3365
rect 9213 3362 9279 3365
rect 5441 3360 9279 3362
rect 5441 3304 5446 3360
rect 5502 3304 9218 3360
rect 9274 3304 9279 3360
rect 5441 3302 9279 3304
rect 5441 3299 5507 3302
rect 9213 3299 9279 3302
rect 9990 3300 9996 3364
rect 10060 3362 10066 3364
rect 13721 3362 13787 3365
rect 10060 3360 13787 3362
rect 10060 3304 13726 3360
rect 13782 3304 13787 3360
rect 10060 3302 13787 3304
rect 15886 3362 15946 3438
rect 17217 3496 38351 3498
rect 17217 3440 17222 3496
rect 17278 3440 38290 3496
rect 38346 3440 38351 3496
rect 17217 3438 38351 3440
rect 17217 3435 17283 3438
rect 38285 3435 38351 3438
rect 41781 3498 41847 3501
rect 45645 3498 45711 3501
rect 41781 3496 45711 3498
rect 41781 3440 41786 3496
rect 41842 3440 45650 3496
rect 45706 3440 45711 3496
rect 41781 3438 45711 3440
rect 41781 3435 41847 3438
rect 45645 3435 45711 3438
rect 16297 3362 16363 3365
rect 15886 3360 16363 3362
rect 15886 3304 16302 3360
rect 16358 3304 16363 3360
rect 15886 3302 16363 3304
rect 10060 3300 10066 3302
rect 13721 3299 13787 3302
rect 16297 3299 16363 3302
rect 16430 3300 16436 3364
rect 16500 3362 16506 3364
rect 17953 3362 18019 3365
rect 27797 3362 27863 3365
rect 16500 3302 17234 3362
rect 16500 3300 16506 3302
rect 15394 3296 15710 3297
rect 15394 3232 15400 3296
rect 15464 3232 15480 3296
rect 15544 3232 15560 3296
rect 15624 3232 15640 3296
rect 15704 3232 15710 3296
rect 15394 3231 15710 3232
rect 7373 3228 7439 3229
rect 7373 3226 7420 3228
rect 7328 3224 7420 3226
rect 7328 3168 7378 3224
rect 7328 3166 7420 3168
rect 7373 3164 7420 3166
rect 7484 3164 7490 3228
rect 7966 3164 7972 3228
rect 8036 3226 8042 3228
rect 8201 3226 8267 3229
rect 8036 3224 8267 3226
rect 8036 3168 8206 3224
rect 8262 3168 8267 3224
rect 8036 3166 8267 3168
rect 8036 3164 8042 3166
rect 7373 3163 7439 3164
rect 8201 3163 8267 3166
rect 8753 3226 8819 3229
rect 14825 3226 14891 3229
rect 15101 3226 15167 3229
rect 8753 3224 15167 3226
rect 8753 3168 8758 3224
rect 8814 3168 14830 3224
rect 14886 3168 15106 3224
rect 15162 3168 15167 3224
rect 8753 3166 15167 3168
rect 17174 3226 17234 3302
rect 17953 3360 27863 3362
rect 17953 3304 17958 3360
rect 18014 3304 27802 3360
rect 27858 3304 27863 3360
rect 17953 3302 27863 3304
rect 17953 3299 18019 3302
rect 27797 3299 27863 3302
rect 31201 3362 31267 3365
rect 37365 3362 37431 3365
rect 31201 3360 37431 3362
rect 31201 3304 31206 3360
rect 31262 3304 37370 3360
rect 37426 3304 37431 3360
rect 31201 3302 37431 3304
rect 31201 3299 31267 3302
rect 37365 3299 37431 3302
rect 42609 3362 42675 3365
rect 43713 3362 43779 3365
rect 42609 3360 43779 3362
rect 42609 3304 42614 3360
rect 42670 3304 43718 3360
rect 43774 3304 43779 3360
rect 42609 3302 43779 3304
rect 42609 3299 42675 3302
rect 43713 3299 43779 3302
rect 29842 3296 30158 3297
rect 29842 3232 29848 3296
rect 29912 3232 29928 3296
rect 29992 3232 30008 3296
rect 30072 3232 30088 3296
rect 30152 3232 30158 3296
rect 29842 3231 30158 3232
rect 44290 3296 44606 3297
rect 44290 3232 44296 3296
rect 44360 3232 44376 3296
rect 44440 3232 44456 3296
rect 44520 3232 44536 3296
rect 44600 3232 44606 3296
rect 44290 3231 44606 3232
rect 19241 3226 19307 3229
rect 17174 3224 19307 3226
rect 17174 3168 19246 3224
rect 19302 3168 19307 3224
rect 17174 3166 19307 3168
rect 8753 3163 8819 3166
rect 14825 3163 14891 3166
rect 15101 3163 15167 3166
rect 19241 3163 19307 3166
rect 23473 3226 23539 3229
rect 23606 3226 23612 3228
rect 23473 3224 23612 3226
rect 23473 3168 23478 3224
rect 23534 3168 23612 3224
rect 23473 3166 23612 3168
rect 23473 3163 23539 3166
rect 23606 3164 23612 3166
rect 23676 3164 23682 3228
rect 36721 3226 36787 3229
rect 39113 3226 39179 3229
rect 44081 3226 44147 3229
rect 36721 3224 39179 3226
rect 36721 3168 36726 3224
rect 36782 3168 39118 3224
rect 39174 3168 39179 3224
rect 36721 3166 39179 3168
rect 36721 3163 36787 3166
rect 39113 3163 39179 3166
rect 39254 3224 44147 3226
rect 39254 3168 44086 3224
rect 44142 3168 44147 3224
rect 39254 3166 44147 3168
rect 5073 3090 5139 3093
rect 31477 3090 31543 3093
rect 37733 3090 37799 3093
rect 5073 3088 26986 3090
rect 5073 3032 5078 3088
rect 5134 3032 26986 3088
rect 5073 3030 26986 3032
rect 5073 3027 5139 3030
rect 4613 2954 4679 2957
rect 10685 2954 10751 2957
rect 11697 2954 11763 2957
rect 4613 2952 10242 2954
rect 4613 2896 4618 2952
rect 4674 2896 10242 2952
rect 4613 2894 10242 2896
rect 4613 2891 4679 2894
rect 8569 2818 8635 2821
rect 9254 2818 9260 2820
rect 8569 2816 9260 2818
rect 8569 2760 8574 2816
rect 8630 2760 9260 2816
rect 8569 2758 9260 2760
rect 8569 2755 8635 2758
rect 9254 2756 9260 2758
rect 9324 2756 9330 2820
rect 8170 2752 8486 2753
rect 8170 2688 8176 2752
rect 8240 2688 8256 2752
rect 8320 2688 8336 2752
rect 8400 2688 8416 2752
rect 8480 2688 8486 2752
rect 8170 2687 8486 2688
rect 10182 2685 10242 2894
rect 10685 2952 11763 2954
rect 10685 2896 10690 2952
rect 10746 2896 11702 2952
rect 11758 2896 11763 2952
rect 10685 2894 11763 2896
rect 10685 2891 10751 2894
rect 11697 2891 11763 2894
rect 15142 2892 15148 2956
rect 15212 2954 15218 2956
rect 15929 2954 15995 2957
rect 15212 2952 15995 2954
rect 15212 2896 15934 2952
rect 15990 2896 15995 2952
rect 15212 2894 15995 2896
rect 15212 2892 15218 2894
rect 15929 2891 15995 2894
rect 17902 2892 17908 2956
rect 17972 2954 17978 2956
rect 19057 2954 19123 2957
rect 17972 2952 19123 2954
rect 17972 2896 19062 2952
rect 19118 2896 19123 2952
rect 17972 2894 19123 2896
rect 17972 2892 17978 2894
rect 19057 2891 19123 2894
rect 19609 2954 19675 2957
rect 26926 2954 26986 3030
rect 31477 3088 37799 3090
rect 31477 3032 31482 3088
rect 31538 3032 37738 3088
rect 37794 3032 37799 3088
rect 31477 3030 37799 3032
rect 31477 3027 31543 3030
rect 37733 3027 37799 3030
rect 39254 2954 39314 3166
rect 44081 3163 44147 3166
rect 41045 3090 41111 3093
rect 43805 3090 43871 3093
rect 48313 3090 48379 3093
rect 41045 3088 41430 3090
rect 41045 3032 41050 3088
rect 41106 3032 41430 3088
rect 41045 3030 41430 3032
rect 41045 3027 41111 3030
rect 19609 2952 26802 2954
rect 19609 2896 19614 2952
rect 19670 2896 26802 2952
rect 19609 2894 26802 2896
rect 26926 2894 39314 2954
rect 41370 2954 41430 3030
rect 43805 3088 48379 3090
rect 43805 3032 43810 3088
rect 43866 3032 48318 3088
rect 48374 3032 48379 3088
rect 43805 3030 48379 3032
rect 43805 3027 43871 3030
rect 48313 3027 48379 3030
rect 48497 3090 48563 3093
rect 54109 3090 54175 3093
rect 48497 3088 54175 3090
rect 48497 3032 48502 3088
rect 48558 3032 54114 3088
rect 54170 3032 54175 3088
rect 48497 3030 54175 3032
rect 48497 3027 48563 3030
rect 54109 3027 54175 3030
rect 45737 2954 45803 2957
rect 41370 2952 45803 2954
rect 41370 2896 45742 2952
rect 45798 2896 45803 2952
rect 41370 2894 45803 2896
rect 19609 2891 19675 2894
rect 12934 2756 12940 2820
rect 13004 2818 13010 2820
rect 13629 2818 13695 2821
rect 13004 2816 13695 2818
rect 13004 2760 13634 2816
rect 13690 2760 13695 2816
rect 13004 2758 13695 2760
rect 13004 2756 13010 2758
rect 13629 2755 13695 2758
rect 14958 2756 14964 2820
rect 15028 2818 15034 2820
rect 15653 2818 15719 2821
rect 15028 2816 15719 2818
rect 15028 2760 15658 2816
rect 15714 2760 15719 2816
rect 15028 2758 15719 2760
rect 26742 2818 26802 2894
rect 45737 2891 45803 2894
rect 50521 2954 50587 2957
rect 53833 2954 53899 2957
rect 50521 2952 53899 2954
rect 50521 2896 50526 2952
rect 50582 2896 53838 2952
rect 53894 2896 53899 2952
rect 50521 2894 53899 2896
rect 50521 2891 50587 2894
rect 53833 2891 53899 2894
rect 30833 2818 30899 2821
rect 26742 2816 30899 2818
rect 26742 2760 30838 2816
rect 30894 2760 30899 2816
rect 26742 2758 30899 2760
rect 15028 2756 15034 2758
rect 15653 2755 15719 2758
rect 30833 2755 30899 2758
rect 37733 2818 37799 2821
rect 40769 2818 40835 2821
rect 37733 2816 40835 2818
rect 37733 2760 37738 2816
rect 37794 2760 40774 2816
rect 40830 2760 40835 2816
rect 37733 2758 40835 2760
rect 37733 2755 37799 2758
rect 40769 2755 40835 2758
rect 42793 2818 42859 2821
rect 49969 2818 50035 2821
rect 42793 2816 50035 2818
rect 42793 2760 42798 2816
rect 42854 2760 49974 2816
rect 50030 2760 50035 2816
rect 42793 2758 50035 2760
rect 42793 2755 42859 2758
rect 49969 2755 50035 2758
rect 22618 2752 22934 2753
rect 22618 2688 22624 2752
rect 22688 2688 22704 2752
rect 22768 2688 22784 2752
rect 22848 2688 22864 2752
rect 22928 2688 22934 2752
rect 22618 2687 22934 2688
rect 37066 2752 37382 2753
rect 37066 2688 37072 2752
rect 37136 2688 37152 2752
rect 37216 2688 37232 2752
rect 37296 2688 37312 2752
rect 37376 2688 37382 2752
rect 37066 2687 37382 2688
rect 51514 2752 51830 2753
rect 51514 2688 51520 2752
rect 51584 2688 51600 2752
rect 51664 2688 51680 2752
rect 51744 2688 51760 2752
rect 51824 2688 51830 2752
rect 51514 2687 51830 2688
rect 2221 2682 2287 2685
rect 4654 2682 4660 2684
rect 2221 2680 4660 2682
rect 2221 2624 2226 2680
rect 2282 2624 4660 2680
rect 2221 2622 4660 2624
rect 2221 2619 2287 2622
rect 4654 2620 4660 2622
rect 4724 2620 4730 2684
rect 10182 2680 10291 2685
rect 10182 2624 10230 2680
rect 10286 2624 10291 2680
rect 10182 2622 10291 2624
rect 10225 2619 10291 2622
rect 17677 2684 17743 2685
rect 17677 2680 17724 2684
rect 17788 2682 17794 2684
rect 47853 2682 47919 2685
rect 50153 2682 50219 2685
rect 17677 2624 17682 2680
rect 17677 2620 17724 2624
rect 17788 2622 17834 2682
rect 47853 2680 50219 2682
rect 47853 2624 47858 2680
rect 47914 2624 50158 2680
rect 50214 2624 50219 2680
rect 47853 2622 50219 2624
rect 17788 2620 17794 2622
rect 17677 2619 17743 2620
rect 47853 2619 47919 2622
rect 50153 2619 50219 2622
rect 6637 2546 6703 2549
rect 16849 2546 16915 2549
rect 6637 2544 16915 2546
rect 6637 2488 6642 2544
rect 6698 2488 16854 2544
rect 16910 2488 16915 2544
rect 6637 2486 16915 2488
rect 6637 2483 6703 2486
rect 16849 2483 16915 2486
rect 17217 2546 17283 2549
rect 19793 2546 19859 2549
rect 17217 2544 19859 2546
rect 17217 2488 17222 2544
rect 17278 2488 19798 2544
rect 19854 2488 19859 2544
rect 17217 2486 19859 2488
rect 17217 2483 17283 2486
rect 19793 2483 19859 2486
rect 34605 2546 34671 2549
rect 39205 2546 39271 2549
rect 34605 2544 39271 2546
rect 34605 2488 34610 2544
rect 34666 2488 39210 2544
rect 39266 2488 39271 2544
rect 34605 2486 39271 2488
rect 34605 2483 34671 2486
rect 39205 2483 39271 2486
rect 40677 2546 40743 2549
rect 43897 2546 43963 2549
rect 40677 2544 43963 2546
rect 40677 2488 40682 2544
rect 40738 2488 43902 2544
rect 43958 2488 43963 2544
rect 40677 2486 43963 2488
rect 40677 2483 40743 2486
rect 43897 2483 43963 2486
rect 44081 2546 44147 2549
rect 52085 2546 52151 2549
rect 44081 2544 52151 2546
rect 44081 2488 44086 2544
rect 44142 2488 52090 2544
rect 52146 2488 52151 2544
rect 44081 2486 52151 2488
rect 44081 2483 44147 2486
rect 52085 2483 52151 2486
rect 9213 2410 9279 2413
rect 9438 2410 9444 2412
rect 9213 2408 9444 2410
rect 9213 2352 9218 2408
rect 9274 2352 9444 2408
rect 9213 2350 9444 2352
rect 9213 2347 9279 2350
rect 9438 2348 9444 2350
rect 9508 2348 9514 2412
rect 26969 2410 27035 2413
rect 12390 2408 27035 2410
rect 12390 2352 26974 2408
rect 27030 2352 27035 2408
rect 12390 2350 27035 2352
rect 7598 2212 7604 2276
rect 7668 2274 7674 2276
rect 12390 2274 12450 2350
rect 26969 2347 27035 2350
rect 38469 2410 38535 2413
rect 49509 2410 49575 2413
rect 38469 2408 49575 2410
rect 38469 2352 38474 2408
rect 38530 2352 49514 2408
rect 49570 2352 49575 2408
rect 38469 2350 49575 2352
rect 38469 2347 38535 2350
rect 49509 2347 49575 2350
rect 7668 2214 12450 2274
rect 22001 2274 22067 2277
rect 27981 2274 28047 2277
rect 22001 2272 28047 2274
rect 22001 2216 22006 2272
rect 22062 2216 27986 2272
rect 28042 2216 28047 2272
rect 22001 2214 28047 2216
rect 7668 2212 7674 2214
rect 22001 2211 22067 2214
rect 27981 2211 28047 2214
rect 34462 2212 34468 2276
rect 34532 2274 34538 2276
rect 35709 2274 35775 2277
rect 41781 2274 41847 2277
rect 34532 2272 41847 2274
rect 34532 2216 35714 2272
rect 35770 2216 41786 2272
rect 41842 2216 41847 2272
rect 34532 2214 41847 2216
rect 34532 2212 34538 2214
rect 35709 2211 35775 2214
rect 41781 2211 41847 2214
rect 15394 2208 15710 2209
rect 15394 2144 15400 2208
rect 15464 2144 15480 2208
rect 15544 2144 15560 2208
rect 15624 2144 15640 2208
rect 15704 2144 15710 2208
rect 15394 2143 15710 2144
rect 29842 2208 30158 2209
rect 29842 2144 29848 2208
rect 29912 2144 29928 2208
rect 29992 2144 30008 2208
rect 30072 2144 30088 2208
rect 30152 2144 30158 2208
rect 29842 2143 30158 2144
rect 44290 2208 44606 2209
rect 44290 2144 44296 2208
rect 44360 2144 44376 2208
rect 44440 2144 44456 2208
rect 44520 2144 44536 2208
rect 44600 2144 44606 2208
rect 44290 2143 44606 2144
rect 8886 2076 8892 2140
rect 8956 2138 8962 2140
rect 9029 2138 9095 2141
rect 8956 2136 9095 2138
rect 8956 2080 9034 2136
rect 9090 2080 9095 2136
rect 8956 2078 9095 2080
rect 8956 2076 8962 2078
rect 9029 2075 9095 2078
rect 23013 2138 23079 2141
rect 23013 2136 23536 2138
rect 23013 2080 23018 2136
rect 23074 2080 23536 2136
rect 23013 2078 23536 2080
rect 23013 2075 23079 2078
rect 3969 2002 4035 2005
rect 23197 2002 23263 2005
rect 3969 2000 23263 2002
rect 3969 1944 3974 2000
rect 4030 1944 23202 2000
rect 23258 1944 23263 2000
rect 3969 1942 23263 1944
rect 23476 2002 23536 2078
rect 38561 2002 38627 2005
rect 23476 2000 38627 2002
rect 23476 1944 38566 2000
rect 38622 1944 38627 2000
rect 23476 1942 38627 1944
rect 3969 1939 4035 1942
rect 23197 1939 23263 1942
rect 38561 1939 38627 1942
rect 42517 2002 42583 2005
rect 50153 2002 50219 2005
rect 42517 2000 50219 2002
rect 42517 1944 42522 2000
rect 42578 1944 50158 2000
rect 50214 1944 50219 2000
rect 42517 1942 50219 1944
rect 42517 1939 42583 1942
rect 50153 1939 50219 1942
rect 6821 1866 6887 1869
rect 18781 1866 18847 1869
rect 6821 1864 18847 1866
rect 6821 1808 6826 1864
rect 6882 1808 18786 1864
rect 18842 1808 18847 1864
rect 6821 1806 18847 1808
rect 6821 1803 6887 1806
rect 18781 1803 18847 1806
rect 26417 1866 26483 1869
rect 29361 1866 29427 1869
rect 39297 1866 39363 1869
rect 26417 1864 39363 1866
rect 26417 1808 26422 1864
rect 26478 1808 29366 1864
rect 29422 1808 39302 1864
rect 39358 1808 39363 1864
rect 26417 1806 39363 1808
rect 26417 1803 26483 1806
rect 29361 1803 29427 1806
rect 39297 1803 39363 1806
rect 42241 1866 42307 1869
rect 48865 1866 48931 1869
rect 42241 1864 48931 1866
rect 42241 1808 42246 1864
rect 42302 1808 48870 1864
rect 48926 1808 48931 1864
rect 42241 1806 48931 1808
rect 42241 1803 42307 1806
rect 48865 1803 48931 1806
rect 3877 1730 3943 1733
rect 15193 1730 15259 1733
rect 3877 1728 15259 1730
rect 3877 1672 3882 1728
rect 3938 1672 15198 1728
rect 15254 1672 15259 1728
rect 3877 1670 15259 1672
rect 3877 1667 3943 1670
rect 15193 1667 15259 1670
rect 25865 1730 25931 1733
rect 42609 1730 42675 1733
rect 25865 1728 42675 1730
rect 25865 1672 25870 1728
rect 25926 1672 42614 1728
rect 42670 1672 42675 1728
rect 25865 1670 42675 1672
rect 25865 1667 25931 1670
rect 42609 1667 42675 1670
rect 11789 1594 11855 1597
rect 30741 1594 30807 1597
rect 11789 1592 30807 1594
rect 11789 1536 11794 1592
rect 11850 1536 30746 1592
rect 30802 1536 30807 1592
rect 11789 1534 30807 1536
rect 11789 1531 11855 1534
rect 30741 1531 30807 1534
rect 38561 1594 38627 1597
rect 53925 1594 53991 1597
rect 38561 1592 53991 1594
rect 38561 1536 38566 1592
rect 38622 1536 53930 1592
rect 53986 1536 53991 1592
rect 38561 1534 53991 1536
rect 38561 1531 38627 1534
rect 53925 1531 53991 1534
rect 22829 1458 22895 1461
rect 36353 1458 36419 1461
rect 22829 1456 36419 1458
rect 22829 1400 22834 1456
rect 22890 1400 36358 1456
rect 36414 1400 36419 1456
rect 22829 1398 36419 1400
rect 22829 1395 22895 1398
rect 36353 1395 36419 1398
rect 12198 1260 12204 1324
rect 12268 1322 12274 1324
rect 42977 1322 43043 1325
rect 12268 1320 43043 1322
rect 12268 1264 42982 1320
rect 43038 1264 43043 1320
rect 12268 1262 43043 1264
rect 12268 1260 12274 1262
rect 42977 1259 43043 1262
rect 23381 1186 23447 1189
rect 51257 1186 51323 1189
rect 23381 1184 51323 1186
rect 23381 1128 23386 1184
rect 23442 1128 51262 1184
rect 51318 1128 51323 1184
rect 23381 1126 51323 1128
rect 23381 1123 23447 1126
rect 51257 1123 51323 1126
rect 10685 1050 10751 1053
rect 34462 1050 34468 1052
rect 10685 1048 34468 1050
rect 10685 992 10690 1048
rect 10746 992 34468 1048
rect 10685 990 34468 992
rect 10685 987 10751 990
rect 34462 988 34468 990
rect 34532 988 34538 1052
<< via3 >>
rect 15400 17436 15464 17440
rect 15400 17380 15404 17436
rect 15404 17380 15460 17436
rect 15460 17380 15464 17436
rect 15400 17376 15464 17380
rect 15480 17436 15544 17440
rect 15480 17380 15484 17436
rect 15484 17380 15540 17436
rect 15540 17380 15544 17436
rect 15480 17376 15544 17380
rect 15560 17436 15624 17440
rect 15560 17380 15564 17436
rect 15564 17380 15620 17436
rect 15620 17380 15624 17436
rect 15560 17376 15624 17380
rect 15640 17436 15704 17440
rect 15640 17380 15644 17436
rect 15644 17380 15700 17436
rect 15700 17380 15704 17436
rect 15640 17376 15704 17380
rect 29848 17436 29912 17440
rect 29848 17380 29852 17436
rect 29852 17380 29908 17436
rect 29908 17380 29912 17436
rect 29848 17376 29912 17380
rect 29928 17436 29992 17440
rect 29928 17380 29932 17436
rect 29932 17380 29988 17436
rect 29988 17380 29992 17436
rect 29928 17376 29992 17380
rect 30008 17436 30072 17440
rect 30008 17380 30012 17436
rect 30012 17380 30068 17436
rect 30068 17380 30072 17436
rect 30008 17376 30072 17380
rect 30088 17436 30152 17440
rect 30088 17380 30092 17436
rect 30092 17380 30148 17436
rect 30148 17380 30152 17436
rect 30088 17376 30152 17380
rect 44296 17436 44360 17440
rect 44296 17380 44300 17436
rect 44300 17380 44356 17436
rect 44356 17380 44360 17436
rect 44296 17376 44360 17380
rect 44376 17436 44440 17440
rect 44376 17380 44380 17436
rect 44380 17380 44436 17436
rect 44436 17380 44440 17436
rect 44376 17376 44440 17380
rect 44456 17436 44520 17440
rect 44456 17380 44460 17436
rect 44460 17380 44516 17436
rect 44516 17380 44520 17436
rect 44456 17376 44520 17380
rect 44536 17436 44600 17440
rect 44536 17380 44540 17436
rect 44540 17380 44596 17436
rect 44596 17380 44600 17436
rect 44536 17376 44600 17380
rect 8176 16892 8240 16896
rect 8176 16836 8180 16892
rect 8180 16836 8236 16892
rect 8236 16836 8240 16892
rect 8176 16832 8240 16836
rect 8256 16892 8320 16896
rect 8256 16836 8260 16892
rect 8260 16836 8316 16892
rect 8316 16836 8320 16892
rect 8256 16832 8320 16836
rect 8336 16892 8400 16896
rect 8336 16836 8340 16892
rect 8340 16836 8396 16892
rect 8396 16836 8400 16892
rect 8336 16832 8400 16836
rect 8416 16892 8480 16896
rect 8416 16836 8420 16892
rect 8420 16836 8476 16892
rect 8476 16836 8480 16892
rect 8416 16832 8480 16836
rect 22624 16892 22688 16896
rect 22624 16836 22628 16892
rect 22628 16836 22684 16892
rect 22684 16836 22688 16892
rect 22624 16832 22688 16836
rect 22704 16892 22768 16896
rect 22704 16836 22708 16892
rect 22708 16836 22764 16892
rect 22764 16836 22768 16892
rect 22704 16832 22768 16836
rect 22784 16892 22848 16896
rect 22784 16836 22788 16892
rect 22788 16836 22844 16892
rect 22844 16836 22848 16892
rect 22784 16832 22848 16836
rect 22864 16892 22928 16896
rect 22864 16836 22868 16892
rect 22868 16836 22924 16892
rect 22924 16836 22928 16892
rect 22864 16832 22928 16836
rect 37072 16892 37136 16896
rect 37072 16836 37076 16892
rect 37076 16836 37132 16892
rect 37132 16836 37136 16892
rect 37072 16832 37136 16836
rect 37152 16892 37216 16896
rect 37152 16836 37156 16892
rect 37156 16836 37212 16892
rect 37212 16836 37216 16892
rect 37152 16832 37216 16836
rect 37232 16892 37296 16896
rect 37232 16836 37236 16892
rect 37236 16836 37292 16892
rect 37292 16836 37296 16892
rect 37232 16832 37296 16836
rect 37312 16892 37376 16896
rect 37312 16836 37316 16892
rect 37316 16836 37372 16892
rect 37372 16836 37376 16892
rect 37312 16832 37376 16836
rect 51520 16892 51584 16896
rect 51520 16836 51524 16892
rect 51524 16836 51580 16892
rect 51580 16836 51584 16892
rect 51520 16832 51584 16836
rect 51600 16892 51664 16896
rect 51600 16836 51604 16892
rect 51604 16836 51660 16892
rect 51660 16836 51664 16892
rect 51600 16832 51664 16836
rect 51680 16892 51744 16896
rect 51680 16836 51684 16892
rect 51684 16836 51740 16892
rect 51740 16836 51744 16892
rect 51680 16832 51744 16836
rect 51760 16892 51824 16896
rect 51760 16836 51764 16892
rect 51764 16836 51820 16892
rect 51820 16836 51824 16892
rect 51760 16832 51824 16836
rect 15400 16348 15464 16352
rect 15400 16292 15404 16348
rect 15404 16292 15460 16348
rect 15460 16292 15464 16348
rect 15400 16288 15464 16292
rect 15480 16348 15544 16352
rect 15480 16292 15484 16348
rect 15484 16292 15540 16348
rect 15540 16292 15544 16348
rect 15480 16288 15544 16292
rect 15560 16348 15624 16352
rect 15560 16292 15564 16348
rect 15564 16292 15620 16348
rect 15620 16292 15624 16348
rect 15560 16288 15624 16292
rect 15640 16348 15704 16352
rect 15640 16292 15644 16348
rect 15644 16292 15700 16348
rect 15700 16292 15704 16348
rect 15640 16288 15704 16292
rect 29848 16348 29912 16352
rect 29848 16292 29852 16348
rect 29852 16292 29908 16348
rect 29908 16292 29912 16348
rect 29848 16288 29912 16292
rect 29928 16348 29992 16352
rect 29928 16292 29932 16348
rect 29932 16292 29988 16348
rect 29988 16292 29992 16348
rect 29928 16288 29992 16292
rect 30008 16348 30072 16352
rect 30008 16292 30012 16348
rect 30012 16292 30068 16348
rect 30068 16292 30072 16348
rect 30008 16288 30072 16292
rect 30088 16348 30152 16352
rect 30088 16292 30092 16348
rect 30092 16292 30148 16348
rect 30148 16292 30152 16348
rect 30088 16288 30152 16292
rect 44296 16348 44360 16352
rect 44296 16292 44300 16348
rect 44300 16292 44356 16348
rect 44356 16292 44360 16348
rect 44296 16288 44360 16292
rect 44376 16348 44440 16352
rect 44376 16292 44380 16348
rect 44380 16292 44436 16348
rect 44436 16292 44440 16348
rect 44376 16288 44440 16292
rect 44456 16348 44520 16352
rect 44456 16292 44460 16348
rect 44460 16292 44516 16348
rect 44516 16292 44520 16348
rect 44456 16288 44520 16292
rect 44536 16348 44600 16352
rect 44536 16292 44540 16348
rect 44540 16292 44596 16348
rect 44596 16292 44600 16348
rect 44536 16288 44600 16292
rect 8176 15804 8240 15808
rect 8176 15748 8180 15804
rect 8180 15748 8236 15804
rect 8236 15748 8240 15804
rect 8176 15744 8240 15748
rect 8256 15804 8320 15808
rect 8256 15748 8260 15804
rect 8260 15748 8316 15804
rect 8316 15748 8320 15804
rect 8256 15744 8320 15748
rect 8336 15804 8400 15808
rect 8336 15748 8340 15804
rect 8340 15748 8396 15804
rect 8396 15748 8400 15804
rect 8336 15744 8400 15748
rect 8416 15804 8480 15808
rect 8416 15748 8420 15804
rect 8420 15748 8476 15804
rect 8476 15748 8480 15804
rect 8416 15744 8480 15748
rect 22624 15804 22688 15808
rect 22624 15748 22628 15804
rect 22628 15748 22684 15804
rect 22684 15748 22688 15804
rect 22624 15744 22688 15748
rect 22704 15804 22768 15808
rect 22704 15748 22708 15804
rect 22708 15748 22764 15804
rect 22764 15748 22768 15804
rect 22704 15744 22768 15748
rect 22784 15804 22848 15808
rect 22784 15748 22788 15804
rect 22788 15748 22844 15804
rect 22844 15748 22848 15804
rect 22784 15744 22848 15748
rect 22864 15804 22928 15808
rect 22864 15748 22868 15804
rect 22868 15748 22924 15804
rect 22924 15748 22928 15804
rect 22864 15744 22928 15748
rect 37072 15804 37136 15808
rect 37072 15748 37076 15804
rect 37076 15748 37132 15804
rect 37132 15748 37136 15804
rect 37072 15744 37136 15748
rect 37152 15804 37216 15808
rect 37152 15748 37156 15804
rect 37156 15748 37212 15804
rect 37212 15748 37216 15804
rect 37152 15744 37216 15748
rect 37232 15804 37296 15808
rect 37232 15748 37236 15804
rect 37236 15748 37292 15804
rect 37292 15748 37296 15804
rect 37232 15744 37296 15748
rect 37312 15804 37376 15808
rect 37312 15748 37316 15804
rect 37316 15748 37372 15804
rect 37372 15748 37376 15804
rect 37312 15744 37376 15748
rect 51520 15804 51584 15808
rect 51520 15748 51524 15804
rect 51524 15748 51580 15804
rect 51580 15748 51584 15804
rect 51520 15744 51584 15748
rect 51600 15804 51664 15808
rect 51600 15748 51604 15804
rect 51604 15748 51660 15804
rect 51660 15748 51664 15804
rect 51600 15744 51664 15748
rect 51680 15804 51744 15808
rect 51680 15748 51684 15804
rect 51684 15748 51740 15804
rect 51740 15748 51744 15804
rect 51680 15744 51744 15748
rect 51760 15804 51824 15808
rect 51760 15748 51764 15804
rect 51764 15748 51820 15804
rect 51820 15748 51824 15804
rect 51760 15744 51824 15748
rect 15400 15260 15464 15264
rect 15400 15204 15404 15260
rect 15404 15204 15460 15260
rect 15460 15204 15464 15260
rect 15400 15200 15464 15204
rect 15480 15260 15544 15264
rect 15480 15204 15484 15260
rect 15484 15204 15540 15260
rect 15540 15204 15544 15260
rect 15480 15200 15544 15204
rect 15560 15260 15624 15264
rect 15560 15204 15564 15260
rect 15564 15204 15620 15260
rect 15620 15204 15624 15260
rect 15560 15200 15624 15204
rect 15640 15260 15704 15264
rect 15640 15204 15644 15260
rect 15644 15204 15700 15260
rect 15700 15204 15704 15260
rect 15640 15200 15704 15204
rect 29848 15260 29912 15264
rect 29848 15204 29852 15260
rect 29852 15204 29908 15260
rect 29908 15204 29912 15260
rect 29848 15200 29912 15204
rect 29928 15260 29992 15264
rect 29928 15204 29932 15260
rect 29932 15204 29988 15260
rect 29988 15204 29992 15260
rect 29928 15200 29992 15204
rect 30008 15260 30072 15264
rect 30008 15204 30012 15260
rect 30012 15204 30068 15260
rect 30068 15204 30072 15260
rect 30008 15200 30072 15204
rect 30088 15260 30152 15264
rect 30088 15204 30092 15260
rect 30092 15204 30148 15260
rect 30148 15204 30152 15260
rect 30088 15200 30152 15204
rect 44296 15260 44360 15264
rect 44296 15204 44300 15260
rect 44300 15204 44356 15260
rect 44356 15204 44360 15260
rect 44296 15200 44360 15204
rect 44376 15260 44440 15264
rect 44376 15204 44380 15260
rect 44380 15204 44436 15260
rect 44436 15204 44440 15260
rect 44376 15200 44440 15204
rect 44456 15260 44520 15264
rect 44456 15204 44460 15260
rect 44460 15204 44516 15260
rect 44516 15204 44520 15260
rect 44456 15200 44520 15204
rect 44536 15260 44600 15264
rect 44536 15204 44540 15260
rect 44540 15204 44596 15260
rect 44596 15204 44600 15260
rect 44536 15200 44600 15204
rect 8176 14716 8240 14720
rect 8176 14660 8180 14716
rect 8180 14660 8236 14716
rect 8236 14660 8240 14716
rect 8176 14656 8240 14660
rect 8256 14716 8320 14720
rect 8256 14660 8260 14716
rect 8260 14660 8316 14716
rect 8316 14660 8320 14716
rect 8256 14656 8320 14660
rect 8336 14716 8400 14720
rect 8336 14660 8340 14716
rect 8340 14660 8396 14716
rect 8396 14660 8400 14716
rect 8336 14656 8400 14660
rect 8416 14716 8480 14720
rect 8416 14660 8420 14716
rect 8420 14660 8476 14716
rect 8476 14660 8480 14716
rect 8416 14656 8480 14660
rect 22624 14716 22688 14720
rect 22624 14660 22628 14716
rect 22628 14660 22684 14716
rect 22684 14660 22688 14716
rect 22624 14656 22688 14660
rect 22704 14716 22768 14720
rect 22704 14660 22708 14716
rect 22708 14660 22764 14716
rect 22764 14660 22768 14716
rect 22704 14656 22768 14660
rect 22784 14716 22848 14720
rect 22784 14660 22788 14716
rect 22788 14660 22844 14716
rect 22844 14660 22848 14716
rect 22784 14656 22848 14660
rect 22864 14716 22928 14720
rect 22864 14660 22868 14716
rect 22868 14660 22924 14716
rect 22924 14660 22928 14716
rect 22864 14656 22928 14660
rect 37072 14716 37136 14720
rect 37072 14660 37076 14716
rect 37076 14660 37132 14716
rect 37132 14660 37136 14716
rect 37072 14656 37136 14660
rect 37152 14716 37216 14720
rect 37152 14660 37156 14716
rect 37156 14660 37212 14716
rect 37212 14660 37216 14716
rect 37152 14656 37216 14660
rect 37232 14716 37296 14720
rect 37232 14660 37236 14716
rect 37236 14660 37292 14716
rect 37292 14660 37296 14716
rect 37232 14656 37296 14660
rect 37312 14716 37376 14720
rect 37312 14660 37316 14716
rect 37316 14660 37372 14716
rect 37372 14660 37376 14716
rect 37312 14656 37376 14660
rect 51520 14716 51584 14720
rect 51520 14660 51524 14716
rect 51524 14660 51580 14716
rect 51580 14660 51584 14716
rect 51520 14656 51584 14660
rect 51600 14716 51664 14720
rect 51600 14660 51604 14716
rect 51604 14660 51660 14716
rect 51660 14660 51664 14716
rect 51600 14656 51664 14660
rect 51680 14716 51744 14720
rect 51680 14660 51684 14716
rect 51684 14660 51740 14716
rect 51740 14660 51744 14716
rect 51680 14656 51744 14660
rect 51760 14716 51824 14720
rect 51760 14660 51764 14716
rect 51764 14660 51820 14716
rect 51820 14660 51824 14716
rect 51760 14656 51824 14660
rect 15400 14172 15464 14176
rect 15400 14116 15404 14172
rect 15404 14116 15460 14172
rect 15460 14116 15464 14172
rect 15400 14112 15464 14116
rect 15480 14172 15544 14176
rect 15480 14116 15484 14172
rect 15484 14116 15540 14172
rect 15540 14116 15544 14172
rect 15480 14112 15544 14116
rect 15560 14172 15624 14176
rect 15560 14116 15564 14172
rect 15564 14116 15620 14172
rect 15620 14116 15624 14172
rect 15560 14112 15624 14116
rect 15640 14172 15704 14176
rect 15640 14116 15644 14172
rect 15644 14116 15700 14172
rect 15700 14116 15704 14172
rect 15640 14112 15704 14116
rect 29848 14172 29912 14176
rect 29848 14116 29852 14172
rect 29852 14116 29908 14172
rect 29908 14116 29912 14172
rect 29848 14112 29912 14116
rect 29928 14172 29992 14176
rect 29928 14116 29932 14172
rect 29932 14116 29988 14172
rect 29988 14116 29992 14172
rect 29928 14112 29992 14116
rect 30008 14172 30072 14176
rect 30008 14116 30012 14172
rect 30012 14116 30068 14172
rect 30068 14116 30072 14172
rect 30008 14112 30072 14116
rect 30088 14172 30152 14176
rect 30088 14116 30092 14172
rect 30092 14116 30148 14172
rect 30148 14116 30152 14172
rect 30088 14112 30152 14116
rect 44296 14172 44360 14176
rect 44296 14116 44300 14172
rect 44300 14116 44356 14172
rect 44356 14116 44360 14172
rect 44296 14112 44360 14116
rect 44376 14172 44440 14176
rect 44376 14116 44380 14172
rect 44380 14116 44436 14172
rect 44436 14116 44440 14172
rect 44376 14112 44440 14116
rect 44456 14172 44520 14176
rect 44456 14116 44460 14172
rect 44460 14116 44516 14172
rect 44516 14116 44520 14172
rect 44456 14112 44520 14116
rect 44536 14172 44600 14176
rect 44536 14116 44540 14172
rect 44540 14116 44596 14172
rect 44596 14116 44600 14172
rect 44536 14112 44600 14116
rect 13308 13832 13372 13836
rect 13308 13776 13358 13832
rect 13358 13776 13372 13832
rect 13308 13772 13372 13776
rect 8176 13628 8240 13632
rect 8176 13572 8180 13628
rect 8180 13572 8236 13628
rect 8236 13572 8240 13628
rect 8176 13568 8240 13572
rect 8256 13628 8320 13632
rect 8256 13572 8260 13628
rect 8260 13572 8316 13628
rect 8316 13572 8320 13628
rect 8256 13568 8320 13572
rect 8336 13628 8400 13632
rect 8336 13572 8340 13628
rect 8340 13572 8396 13628
rect 8396 13572 8400 13628
rect 8336 13568 8400 13572
rect 8416 13628 8480 13632
rect 8416 13572 8420 13628
rect 8420 13572 8476 13628
rect 8476 13572 8480 13628
rect 8416 13568 8480 13572
rect 22624 13628 22688 13632
rect 22624 13572 22628 13628
rect 22628 13572 22684 13628
rect 22684 13572 22688 13628
rect 22624 13568 22688 13572
rect 22704 13628 22768 13632
rect 22704 13572 22708 13628
rect 22708 13572 22764 13628
rect 22764 13572 22768 13628
rect 22704 13568 22768 13572
rect 22784 13628 22848 13632
rect 22784 13572 22788 13628
rect 22788 13572 22844 13628
rect 22844 13572 22848 13628
rect 22784 13568 22848 13572
rect 22864 13628 22928 13632
rect 22864 13572 22868 13628
rect 22868 13572 22924 13628
rect 22924 13572 22928 13628
rect 22864 13568 22928 13572
rect 37072 13628 37136 13632
rect 37072 13572 37076 13628
rect 37076 13572 37132 13628
rect 37132 13572 37136 13628
rect 37072 13568 37136 13572
rect 37152 13628 37216 13632
rect 37152 13572 37156 13628
rect 37156 13572 37212 13628
rect 37212 13572 37216 13628
rect 37152 13568 37216 13572
rect 37232 13628 37296 13632
rect 37232 13572 37236 13628
rect 37236 13572 37292 13628
rect 37292 13572 37296 13628
rect 37232 13568 37296 13572
rect 37312 13628 37376 13632
rect 37312 13572 37316 13628
rect 37316 13572 37372 13628
rect 37372 13572 37376 13628
rect 37312 13568 37376 13572
rect 51520 13628 51584 13632
rect 51520 13572 51524 13628
rect 51524 13572 51580 13628
rect 51580 13572 51584 13628
rect 51520 13568 51584 13572
rect 51600 13628 51664 13632
rect 51600 13572 51604 13628
rect 51604 13572 51660 13628
rect 51660 13572 51664 13628
rect 51600 13568 51664 13572
rect 51680 13628 51744 13632
rect 51680 13572 51684 13628
rect 51684 13572 51740 13628
rect 51740 13572 51744 13628
rect 51680 13568 51744 13572
rect 51760 13628 51824 13632
rect 51760 13572 51764 13628
rect 51764 13572 51820 13628
rect 51820 13572 51824 13628
rect 51760 13568 51824 13572
rect 17724 13152 17788 13156
rect 17724 13096 17774 13152
rect 17774 13096 17788 13152
rect 17724 13092 17788 13096
rect 15400 13084 15464 13088
rect 15400 13028 15404 13084
rect 15404 13028 15460 13084
rect 15460 13028 15464 13084
rect 15400 13024 15464 13028
rect 15480 13084 15544 13088
rect 15480 13028 15484 13084
rect 15484 13028 15540 13084
rect 15540 13028 15544 13084
rect 15480 13024 15544 13028
rect 15560 13084 15624 13088
rect 15560 13028 15564 13084
rect 15564 13028 15620 13084
rect 15620 13028 15624 13084
rect 15560 13024 15624 13028
rect 15640 13084 15704 13088
rect 15640 13028 15644 13084
rect 15644 13028 15700 13084
rect 15700 13028 15704 13084
rect 15640 13024 15704 13028
rect 29848 13084 29912 13088
rect 29848 13028 29852 13084
rect 29852 13028 29908 13084
rect 29908 13028 29912 13084
rect 29848 13024 29912 13028
rect 29928 13084 29992 13088
rect 29928 13028 29932 13084
rect 29932 13028 29988 13084
rect 29988 13028 29992 13084
rect 29928 13024 29992 13028
rect 30008 13084 30072 13088
rect 30008 13028 30012 13084
rect 30012 13028 30068 13084
rect 30068 13028 30072 13084
rect 30008 13024 30072 13028
rect 30088 13084 30152 13088
rect 30088 13028 30092 13084
rect 30092 13028 30148 13084
rect 30148 13028 30152 13084
rect 30088 13024 30152 13028
rect 44296 13084 44360 13088
rect 44296 13028 44300 13084
rect 44300 13028 44356 13084
rect 44356 13028 44360 13084
rect 44296 13024 44360 13028
rect 44376 13084 44440 13088
rect 44376 13028 44380 13084
rect 44380 13028 44436 13084
rect 44436 13028 44440 13084
rect 44376 13024 44440 13028
rect 44456 13084 44520 13088
rect 44456 13028 44460 13084
rect 44460 13028 44516 13084
rect 44516 13028 44520 13084
rect 44456 13024 44520 13028
rect 44536 13084 44600 13088
rect 44536 13028 44540 13084
rect 44540 13028 44596 13084
rect 44596 13028 44600 13084
rect 44536 13024 44600 13028
rect 10732 12684 10796 12748
rect 14596 12684 14660 12748
rect 10916 12608 10980 12612
rect 10916 12552 10966 12608
rect 10966 12552 10980 12608
rect 10916 12548 10980 12552
rect 19196 12548 19260 12612
rect 8176 12540 8240 12544
rect 8176 12484 8180 12540
rect 8180 12484 8236 12540
rect 8236 12484 8240 12540
rect 8176 12480 8240 12484
rect 8256 12540 8320 12544
rect 8256 12484 8260 12540
rect 8260 12484 8316 12540
rect 8316 12484 8320 12540
rect 8256 12480 8320 12484
rect 8336 12540 8400 12544
rect 8336 12484 8340 12540
rect 8340 12484 8396 12540
rect 8396 12484 8400 12540
rect 8336 12480 8400 12484
rect 8416 12540 8480 12544
rect 8416 12484 8420 12540
rect 8420 12484 8476 12540
rect 8476 12484 8480 12540
rect 8416 12480 8480 12484
rect 22624 12540 22688 12544
rect 22624 12484 22628 12540
rect 22628 12484 22684 12540
rect 22684 12484 22688 12540
rect 22624 12480 22688 12484
rect 22704 12540 22768 12544
rect 22704 12484 22708 12540
rect 22708 12484 22764 12540
rect 22764 12484 22768 12540
rect 22704 12480 22768 12484
rect 22784 12540 22848 12544
rect 22784 12484 22788 12540
rect 22788 12484 22844 12540
rect 22844 12484 22848 12540
rect 22784 12480 22848 12484
rect 22864 12540 22928 12544
rect 22864 12484 22868 12540
rect 22868 12484 22924 12540
rect 22924 12484 22928 12540
rect 22864 12480 22928 12484
rect 37072 12540 37136 12544
rect 37072 12484 37076 12540
rect 37076 12484 37132 12540
rect 37132 12484 37136 12540
rect 37072 12480 37136 12484
rect 37152 12540 37216 12544
rect 37152 12484 37156 12540
rect 37156 12484 37212 12540
rect 37212 12484 37216 12540
rect 37152 12480 37216 12484
rect 37232 12540 37296 12544
rect 37232 12484 37236 12540
rect 37236 12484 37292 12540
rect 37292 12484 37296 12540
rect 37232 12480 37296 12484
rect 37312 12540 37376 12544
rect 37312 12484 37316 12540
rect 37316 12484 37372 12540
rect 37372 12484 37376 12540
rect 37312 12480 37376 12484
rect 51520 12540 51584 12544
rect 51520 12484 51524 12540
rect 51524 12484 51580 12540
rect 51580 12484 51584 12540
rect 51520 12480 51584 12484
rect 51600 12540 51664 12544
rect 51600 12484 51604 12540
rect 51604 12484 51660 12540
rect 51660 12484 51664 12540
rect 51600 12480 51664 12484
rect 51680 12540 51744 12544
rect 51680 12484 51684 12540
rect 51684 12484 51740 12540
rect 51740 12484 51744 12540
rect 51680 12480 51744 12484
rect 51760 12540 51824 12544
rect 51760 12484 51764 12540
rect 51764 12484 51820 12540
rect 51820 12484 51824 12540
rect 51760 12480 51824 12484
rect 1900 12472 1964 12476
rect 1900 12416 1950 12472
rect 1950 12416 1964 12472
rect 1900 12412 1964 12416
rect 2820 12412 2884 12476
rect 6684 12412 6748 12476
rect 16988 12412 17052 12476
rect 23428 12472 23492 12476
rect 23428 12416 23478 12472
rect 23478 12416 23492 12472
rect 23428 12412 23492 12416
rect 14228 12064 14292 12068
rect 14228 12008 14242 12064
rect 14242 12008 14292 12064
rect 14228 12004 14292 12008
rect 18644 12064 18708 12068
rect 18644 12008 18658 12064
rect 18658 12008 18708 12064
rect 18644 12004 18708 12008
rect 22324 12064 22388 12068
rect 22324 12008 22338 12064
rect 22338 12008 22388 12064
rect 22324 12004 22388 12008
rect 15400 11996 15464 12000
rect 15400 11940 15404 11996
rect 15404 11940 15460 11996
rect 15460 11940 15464 11996
rect 15400 11936 15464 11940
rect 15480 11996 15544 12000
rect 15480 11940 15484 11996
rect 15484 11940 15540 11996
rect 15540 11940 15544 11996
rect 15480 11936 15544 11940
rect 15560 11996 15624 12000
rect 15560 11940 15564 11996
rect 15564 11940 15620 11996
rect 15620 11940 15624 11996
rect 15560 11936 15624 11940
rect 15640 11996 15704 12000
rect 15640 11940 15644 11996
rect 15644 11940 15700 11996
rect 15700 11940 15704 11996
rect 15640 11936 15704 11940
rect 29848 11996 29912 12000
rect 29848 11940 29852 11996
rect 29852 11940 29908 11996
rect 29908 11940 29912 11996
rect 29848 11936 29912 11940
rect 29928 11996 29992 12000
rect 29928 11940 29932 11996
rect 29932 11940 29988 11996
rect 29988 11940 29992 11996
rect 29928 11936 29992 11940
rect 30008 11996 30072 12000
rect 30008 11940 30012 11996
rect 30012 11940 30068 11996
rect 30068 11940 30072 11996
rect 30008 11936 30072 11940
rect 30088 11996 30152 12000
rect 30088 11940 30092 11996
rect 30092 11940 30148 11996
rect 30148 11940 30152 11996
rect 30088 11936 30152 11940
rect 44296 11996 44360 12000
rect 44296 11940 44300 11996
rect 44300 11940 44356 11996
rect 44356 11940 44360 11996
rect 44296 11936 44360 11940
rect 44376 11996 44440 12000
rect 44376 11940 44380 11996
rect 44380 11940 44436 11996
rect 44436 11940 44440 11996
rect 44376 11936 44440 11940
rect 44456 11996 44520 12000
rect 44456 11940 44460 11996
rect 44460 11940 44516 11996
rect 44516 11940 44520 11996
rect 44456 11936 44520 11940
rect 44536 11996 44600 12000
rect 44536 11940 44540 11996
rect 44540 11940 44596 11996
rect 44596 11940 44600 11996
rect 44536 11936 44600 11940
rect 14596 11732 14660 11796
rect 5948 11460 6012 11524
rect 22140 11520 22204 11524
rect 22140 11464 22154 11520
rect 22154 11464 22204 11520
rect 22140 11460 22204 11464
rect 8176 11452 8240 11456
rect 8176 11396 8180 11452
rect 8180 11396 8236 11452
rect 8236 11396 8240 11452
rect 8176 11392 8240 11396
rect 8256 11452 8320 11456
rect 8256 11396 8260 11452
rect 8260 11396 8316 11452
rect 8316 11396 8320 11452
rect 8256 11392 8320 11396
rect 8336 11452 8400 11456
rect 8336 11396 8340 11452
rect 8340 11396 8396 11452
rect 8396 11396 8400 11452
rect 8336 11392 8400 11396
rect 8416 11452 8480 11456
rect 8416 11396 8420 11452
rect 8420 11396 8476 11452
rect 8476 11396 8480 11452
rect 8416 11392 8480 11396
rect 22624 11452 22688 11456
rect 22624 11396 22628 11452
rect 22628 11396 22684 11452
rect 22684 11396 22688 11452
rect 22624 11392 22688 11396
rect 22704 11452 22768 11456
rect 22704 11396 22708 11452
rect 22708 11396 22764 11452
rect 22764 11396 22768 11452
rect 22704 11392 22768 11396
rect 22784 11452 22848 11456
rect 22784 11396 22788 11452
rect 22788 11396 22844 11452
rect 22844 11396 22848 11452
rect 22784 11392 22848 11396
rect 22864 11452 22928 11456
rect 22864 11396 22868 11452
rect 22868 11396 22924 11452
rect 22924 11396 22928 11452
rect 22864 11392 22928 11396
rect 37072 11452 37136 11456
rect 37072 11396 37076 11452
rect 37076 11396 37132 11452
rect 37132 11396 37136 11452
rect 37072 11392 37136 11396
rect 37152 11452 37216 11456
rect 37152 11396 37156 11452
rect 37156 11396 37212 11452
rect 37212 11396 37216 11452
rect 37152 11392 37216 11396
rect 37232 11452 37296 11456
rect 37232 11396 37236 11452
rect 37236 11396 37292 11452
rect 37292 11396 37296 11452
rect 37232 11392 37296 11396
rect 37312 11452 37376 11456
rect 37312 11396 37316 11452
rect 37316 11396 37372 11452
rect 37372 11396 37376 11452
rect 37312 11392 37376 11396
rect 51520 11452 51584 11456
rect 51520 11396 51524 11452
rect 51524 11396 51580 11452
rect 51580 11396 51584 11452
rect 51520 11392 51584 11396
rect 51600 11452 51664 11456
rect 51600 11396 51604 11452
rect 51604 11396 51660 11452
rect 51660 11396 51664 11452
rect 51600 11392 51664 11396
rect 51680 11452 51744 11456
rect 51680 11396 51684 11452
rect 51684 11396 51740 11452
rect 51740 11396 51744 11452
rect 51680 11392 51744 11396
rect 51760 11452 51824 11456
rect 51760 11396 51764 11452
rect 51764 11396 51820 11452
rect 51820 11396 51824 11452
rect 51760 11392 51824 11396
rect 12940 11188 13004 11252
rect 4660 11052 4724 11116
rect 15148 11112 15212 11116
rect 15148 11056 15162 11112
rect 15162 11056 15212 11112
rect 15148 11052 15212 11056
rect 18276 11052 18340 11116
rect 23060 11052 23124 11116
rect 35756 11112 35820 11116
rect 35756 11056 35770 11112
rect 35770 11056 35820 11112
rect 35756 11052 35820 11056
rect 15400 10908 15464 10912
rect 15400 10852 15404 10908
rect 15404 10852 15460 10908
rect 15460 10852 15464 10908
rect 15400 10848 15464 10852
rect 15480 10908 15544 10912
rect 15480 10852 15484 10908
rect 15484 10852 15540 10908
rect 15540 10852 15544 10908
rect 15480 10848 15544 10852
rect 15560 10908 15624 10912
rect 15560 10852 15564 10908
rect 15564 10852 15620 10908
rect 15620 10852 15624 10908
rect 15560 10848 15624 10852
rect 15640 10908 15704 10912
rect 15640 10852 15644 10908
rect 15644 10852 15700 10908
rect 15700 10852 15704 10908
rect 15640 10848 15704 10852
rect 29848 10908 29912 10912
rect 29848 10852 29852 10908
rect 29852 10852 29908 10908
rect 29908 10852 29912 10908
rect 29848 10848 29912 10852
rect 29928 10908 29992 10912
rect 29928 10852 29932 10908
rect 29932 10852 29988 10908
rect 29988 10852 29992 10908
rect 29928 10848 29992 10852
rect 30008 10908 30072 10912
rect 30008 10852 30012 10908
rect 30012 10852 30068 10908
rect 30068 10852 30072 10908
rect 30008 10848 30072 10852
rect 30088 10908 30152 10912
rect 30088 10852 30092 10908
rect 30092 10852 30148 10908
rect 30148 10852 30152 10908
rect 30088 10848 30152 10852
rect 44296 10908 44360 10912
rect 44296 10852 44300 10908
rect 44300 10852 44356 10908
rect 44356 10852 44360 10908
rect 44296 10848 44360 10852
rect 44376 10908 44440 10912
rect 44376 10852 44380 10908
rect 44380 10852 44436 10908
rect 44436 10852 44440 10908
rect 44376 10848 44440 10852
rect 44456 10908 44520 10912
rect 44456 10852 44460 10908
rect 44460 10852 44516 10908
rect 44516 10852 44520 10908
rect 44456 10848 44520 10852
rect 44536 10908 44600 10912
rect 44536 10852 44540 10908
rect 44540 10852 44596 10908
rect 44596 10852 44600 10908
rect 44536 10848 44600 10852
rect 9260 10508 9324 10572
rect 8176 10364 8240 10368
rect 8176 10308 8180 10364
rect 8180 10308 8236 10364
rect 8236 10308 8240 10364
rect 8176 10304 8240 10308
rect 8256 10364 8320 10368
rect 8256 10308 8260 10364
rect 8260 10308 8316 10364
rect 8316 10308 8320 10364
rect 8256 10304 8320 10308
rect 8336 10364 8400 10368
rect 8336 10308 8340 10364
rect 8340 10308 8396 10364
rect 8396 10308 8400 10364
rect 8336 10304 8400 10308
rect 8416 10364 8480 10368
rect 8416 10308 8420 10364
rect 8420 10308 8476 10364
rect 8476 10308 8480 10364
rect 8416 10304 8480 10308
rect 22624 10364 22688 10368
rect 22624 10308 22628 10364
rect 22628 10308 22684 10364
rect 22684 10308 22688 10364
rect 22624 10304 22688 10308
rect 22704 10364 22768 10368
rect 22704 10308 22708 10364
rect 22708 10308 22764 10364
rect 22764 10308 22768 10364
rect 22704 10304 22768 10308
rect 22784 10364 22848 10368
rect 22784 10308 22788 10364
rect 22788 10308 22844 10364
rect 22844 10308 22848 10364
rect 22784 10304 22848 10308
rect 22864 10364 22928 10368
rect 22864 10308 22868 10364
rect 22868 10308 22924 10364
rect 22924 10308 22928 10364
rect 22864 10304 22928 10308
rect 37072 10364 37136 10368
rect 37072 10308 37076 10364
rect 37076 10308 37132 10364
rect 37132 10308 37136 10364
rect 37072 10304 37136 10308
rect 37152 10364 37216 10368
rect 37152 10308 37156 10364
rect 37156 10308 37212 10364
rect 37212 10308 37216 10364
rect 37152 10304 37216 10308
rect 37232 10364 37296 10368
rect 37232 10308 37236 10364
rect 37236 10308 37292 10364
rect 37292 10308 37296 10364
rect 37232 10304 37296 10308
rect 37312 10364 37376 10368
rect 37312 10308 37316 10364
rect 37316 10308 37372 10364
rect 37372 10308 37376 10364
rect 37312 10304 37376 10308
rect 51520 10364 51584 10368
rect 51520 10308 51524 10364
rect 51524 10308 51580 10364
rect 51580 10308 51584 10364
rect 51520 10304 51584 10308
rect 51600 10364 51664 10368
rect 51600 10308 51604 10364
rect 51604 10308 51660 10364
rect 51660 10308 51664 10364
rect 51600 10304 51664 10308
rect 51680 10364 51744 10368
rect 51680 10308 51684 10364
rect 51684 10308 51740 10364
rect 51740 10308 51744 10364
rect 51680 10304 51744 10308
rect 51760 10364 51824 10368
rect 51760 10308 51764 10364
rect 51764 10308 51820 10364
rect 51820 10308 51824 10364
rect 51760 10304 51824 10308
rect 16620 10100 16684 10164
rect 9076 9964 9140 10028
rect 10916 9964 10980 10028
rect 8892 9828 8956 9892
rect 15400 9820 15464 9824
rect 15400 9764 15404 9820
rect 15404 9764 15460 9820
rect 15460 9764 15464 9820
rect 15400 9760 15464 9764
rect 15480 9820 15544 9824
rect 15480 9764 15484 9820
rect 15484 9764 15540 9820
rect 15540 9764 15544 9820
rect 15480 9760 15544 9764
rect 15560 9820 15624 9824
rect 15560 9764 15564 9820
rect 15564 9764 15620 9820
rect 15620 9764 15624 9820
rect 15560 9760 15624 9764
rect 15640 9820 15704 9824
rect 15640 9764 15644 9820
rect 15644 9764 15700 9820
rect 15700 9764 15704 9820
rect 15640 9760 15704 9764
rect 29848 9820 29912 9824
rect 29848 9764 29852 9820
rect 29852 9764 29908 9820
rect 29908 9764 29912 9820
rect 29848 9760 29912 9764
rect 29928 9820 29992 9824
rect 29928 9764 29932 9820
rect 29932 9764 29988 9820
rect 29988 9764 29992 9820
rect 29928 9760 29992 9764
rect 30008 9820 30072 9824
rect 30008 9764 30012 9820
rect 30012 9764 30068 9820
rect 30068 9764 30072 9820
rect 30008 9760 30072 9764
rect 30088 9820 30152 9824
rect 30088 9764 30092 9820
rect 30092 9764 30148 9820
rect 30148 9764 30152 9820
rect 30088 9760 30152 9764
rect 44296 9820 44360 9824
rect 44296 9764 44300 9820
rect 44300 9764 44356 9820
rect 44356 9764 44360 9820
rect 44296 9760 44360 9764
rect 44376 9820 44440 9824
rect 44376 9764 44380 9820
rect 44380 9764 44436 9820
rect 44436 9764 44440 9820
rect 44376 9760 44440 9764
rect 44456 9820 44520 9824
rect 44456 9764 44460 9820
rect 44460 9764 44516 9820
rect 44516 9764 44520 9820
rect 44456 9760 44520 9764
rect 44536 9820 44600 9824
rect 44536 9764 44540 9820
rect 44540 9764 44596 9820
rect 44596 9764 44600 9820
rect 44536 9760 44600 9764
rect 8708 9692 8772 9756
rect 8176 9276 8240 9280
rect 8176 9220 8180 9276
rect 8180 9220 8236 9276
rect 8236 9220 8240 9276
rect 8176 9216 8240 9220
rect 8256 9276 8320 9280
rect 8256 9220 8260 9276
rect 8260 9220 8316 9276
rect 8316 9220 8320 9276
rect 8256 9216 8320 9220
rect 8336 9276 8400 9280
rect 8336 9220 8340 9276
rect 8340 9220 8396 9276
rect 8396 9220 8400 9276
rect 8336 9216 8400 9220
rect 8416 9276 8480 9280
rect 8416 9220 8420 9276
rect 8420 9220 8476 9276
rect 8476 9220 8480 9276
rect 8416 9216 8480 9220
rect 22624 9276 22688 9280
rect 22624 9220 22628 9276
rect 22628 9220 22684 9276
rect 22684 9220 22688 9276
rect 22624 9216 22688 9220
rect 22704 9276 22768 9280
rect 22704 9220 22708 9276
rect 22708 9220 22764 9276
rect 22764 9220 22768 9276
rect 22704 9216 22768 9220
rect 22784 9276 22848 9280
rect 22784 9220 22788 9276
rect 22788 9220 22844 9276
rect 22844 9220 22848 9276
rect 22784 9216 22848 9220
rect 22864 9276 22928 9280
rect 22864 9220 22868 9276
rect 22868 9220 22924 9276
rect 22924 9220 22928 9276
rect 22864 9216 22928 9220
rect 37072 9276 37136 9280
rect 37072 9220 37076 9276
rect 37076 9220 37132 9276
rect 37132 9220 37136 9276
rect 37072 9216 37136 9220
rect 37152 9276 37216 9280
rect 37152 9220 37156 9276
rect 37156 9220 37212 9276
rect 37212 9220 37216 9276
rect 37152 9216 37216 9220
rect 37232 9276 37296 9280
rect 37232 9220 37236 9276
rect 37236 9220 37292 9276
rect 37292 9220 37296 9276
rect 37232 9216 37296 9220
rect 37312 9276 37376 9280
rect 37312 9220 37316 9276
rect 37316 9220 37372 9276
rect 37372 9220 37376 9276
rect 37312 9216 37376 9220
rect 51520 9276 51584 9280
rect 51520 9220 51524 9276
rect 51524 9220 51580 9276
rect 51580 9220 51584 9276
rect 51520 9216 51584 9220
rect 51600 9276 51664 9280
rect 51600 9220 51604 9276
rect 51604 9220 51660 9276
rect 51660 9220 51664 9276
rect 51600 9216 51664 9220
rect 51680 9276 51744 9280
rect 51680 9220 51684 9276
rect 51684 9220 51740 9276
rect 51740 9220 51744 9276
rect 51680 9216 51744 9220
rect 51760 9276 51824 9280
rect 51760 9220 51764 9276
rect 51764 9220 51820 9276
rect 51820 9220 51824 9276
rect 51760 9216 51824 9220
rect 15400 8732 15464 8736
rect 15400 8676 15404 8732
rect 15404 8676 15460 8732
rect 15460 8676 15464 8732
rect 15400 8672 15464 8676
rect 15480 8732 15544 8736
rect 15480 8676 15484 8732
rect 15484 8676 15540 8732
rect 15540 8676 15544 8732
rect 15480 8672 15544 8676
rect 15560 8732 15624 8736
rect 15560 8676 15564 8732
rect 15564 8676 15620 8732
rect 15620 8676 15624 8732
rect 15560 8672 15624 8676
rect 15640 8732 15704 8736
rect 15640 8676 15644 8732
rect 15644 8676 15700 8732
rect 15700 8676 15704 8732
rect 15640 8672 15704 8676
rect 29848 8732 29912 8736
rect 29848 8676 29852 8732
rect 29852 8676 29908 8732
rect 29908 8676 29912 8732
rect 29848 8672 29912 8676
rect 29928 8732 29992 8736
rect 29928 8676 29932 8732
rect 29932 8676 29988 8732
rect 29988 8676 29992 8732
rect 29928 8672 29992 8676
rect 30008 8732 30072 8736
rect 30008 8676 30012 8732
rect 30012 8676 30068 8732
rect 30068 8676 30072 8732
rect 30008 8672 30072 8676
rect 30088 8732 30152 8736
rect 30088 8676 30092 8732
rect 30092 8676 30148 8732
rect 30148 8676 30152 8732
rect 30088 8672 30152 8676
rect 44296 8732 44360 8736
rect 44296 8676 44300 8732
rect 44300 8676 44356 8732
rect 44356 8676 44360 8732
rect 44296 8672 44360 8676
rect 44376 8732 44440 8736
rect 44376 8676 44380 8732
rect 44380 8676 44436 8732
rect 44436 8676 44440 8732
rect 44376 8672 44440 8676
rect 44456 8732 44520 8736
rect 44456 8676 44460 8732
rect 44460 8676 44516 8732
rect 44516 8676 44520 8732
rect 44456 8672 44520 8676
rect 44536 8732 44600 8736
rect 44536 8676 44540 8732
rect 44540 8676 44596 8732
rect 44596 8676 44600 8732
rect 44536 8672 44600 8676
rect 17724 8196 17788 8260
rect 8176 8188 8240 8192
rect 8176 8132 8180 8188
rect 8180 8132 8236 8188
rect 8236 8132 8240 8188
rect 8176 8128 8240 8132
rect 8256 8188 8320 8192
rect 8256 8132 8260 8188
rect 8260 8132 8316 8188
rect 8316 8132 8320 8188
rect 8256 8128 8320 8132
rect 8336 8188 8400 8192
rect 8336 8132 8340 8188
rect 8340 8132 8396 8188
rect 8396 8132 8400 8188
rect 8336 8128 8400 8132
rect 8416 8188 8480 8192
rect 8416 8132 8420 8188
rect 8420 8132 8476 8188
rect 8476 8132 8480 8188
rect 8416 8128 8480 8132
rect 22624 8188 22688 8192
rect 22624 8132 22628 8188
rect 22628 8132 22684 8188
rect 22684 8132 22688 8188
rect 22624 8128 22688 8132
rect 22704 8188 22768 8192
rect 22704 8132 22708 8188
rect 22708 8132 22764 8188
rect 22764 8132 22768 8188
rect 22704 8128 22768 8132
rect 22784 8188 22848 8192
rect 22784 8132 22788 8188
rect 22788 8132 22844 8188
rect 22844 8132 22848 8188
rect 22784 8128 22848 8132
rect 22864 8188 22928 8192
rect 22864 8132 22868 8188
rect 22868 8132 22924 8188
rect 22924 8132 22928 8188
rect 22864 8128 22928 8132
rect 37072 8188 37136 8192
rect 37072 8132 37076 8188
rect 37076 8132 37132 8188
rect 37132 8132 37136 8188
rect 37072 8128 37136 8132
rect 37152 8188 37216 8192
rect 37152 8132 37156 8188
rect 37156 8132 37212 8188
rect 37212 8132 37216 8188
rect 37152 8128 37216 8132
rect 37232 8188 37296 8192
rect 37232 8132 37236 8188
rect 37236 8132 37292 8188
rect 37292 8132 37296 8188
rect 37232 8128 37296 8132
rect 37312 8188 37376 8192
rect 37312 8132 37316 8188
rect 37316 8132 37372 8188
rect 37372 8132 37376 8188
rect 37312 8128 37376 8132
rect 51520 8188 51584 8192
rect 51520 8132 51524 8188
rect 51524 8132 51580 8188
rect 51580 8132 51584 8188
rect 51520 8128 51584 8132
rect 51600 8188 51664 8192
rect 51600 8132 51604 8188
rect 51604 8132 51660 8188
rect 51660 8132 51664 8188
rect 51600 8128 51664 8132
rect 51680 8188 51744 8192
rect 51680 8132 51684 8188
rect 51684 8132 51740 8188
rect 51740 8132 51744 8188
rect 51680 8128 51744 8132
rect 51760 8188 51824 8192
rect 51760 8132 51764 8188
rect 51764 8132 51820 8188
rect 51820 8132 51824 8188
rect 51760 8128 51824 8132
rect 13492 7984 13556 7988
rect 13492 7928 13542 7984
rect 13542 7928 13556 7984
rect 13492 7924 13556 7928
rect 14228 7924 14292 7988
rect 14964 7788 15028 7852
rect 15400 7644 15464 7648
rect 15400 7588 15404 7644
rect 15404 7588 15460 7644
rect 15460 7588 15464 7644
rect 15400 7584 15464 7588
rect 15480 7644 15544 7648
rect 15480 7588 15484 7644
rect 15484 7588 15540 7644
rect 15540 7588 15544 7644
rect 15480 7584 15544 7588
rect 15560 7644 15624 7648
rect 15560 7588 15564 7644
rect 15564 7588 15620 7644
rect 15620 7588 15624 7644
rect 15560 7584 15624 7588
rect 15640 7644 15704 7648
rect 15640 7588 15644 7644
rect 15644 7588 15700 7644
rect 15700 7588 15704 7644
rect 15640 7584 15704 7588
rect 29848 7644 29912 7648
rect 29848 7588 29852 7644
rect 29852 7588 29908 7644
rect 29908 7588 29912 7644
rect 29848 7584 29912 7588
rect 29928 7644 29992 7648
rect 29928 7588 29932 7644
rect 29932 7588 29988 7644
rect 29988 7588 29992 7644
rect 29928 7584 29992 7588
rect 30008 7644 30072 7648
rect 30008 7588 30012 7644
rect 30012 7588 30068 7644
rect 30068 7588 30072 7644
rect 30008 7584 30072 7588
rect 30088 7644 30152 7648
rect 30088 7588 30092 7644
rect 30092 7588 30148 7644
rect 30148 7588 30152 7644
rect 30088 7584 30152 7588
rect 44296 7644 44360 7648
rect 44296 7588 44300 7644
rect 44300 7588 44356 7644
rect 44356 7588 44360 7644
rect 44296 7584 44360 7588
rect 44376 7644 44440 7648
rect 44376 7588 44380 7644
rect 44380 7588 44436 7644
rect 44436 7588 44440 7644
rect 44376 7584 44440 7588
rect 44456 7644 44520 7648
rect 44456 7588 44460 7644
rect 44460 7588 44516 7644
rect 44516 7588 44520 7644
rect 44456 7584 44520 7588
rect 44536 7644 44600 7648
rect 44536 7588 44540 7644
rect 44540 7588 44596 7644
rect 44596 7588 44600 7644
rect 44536 7584 44600 7588
rect 5948 7516 6012 7580
rect 14228 7244 14292 7308
rect 8176 7100 8240 7104
rect 8176 7044 8180 7100
rect 8180 7044 8236 7100
rect 8236 7044 8240 7100
rect 8176 7040 8240 7044
rect 8256 7100 8320 7104
rect 8256 7044 8260 7100
rect 8260 7044 8316 7100
rect 8316 7044 8320 7100
rect 8256 7040 8320 7044
rect 8336 7100 8400 7104
rect 8336 7044 8340 7100
rect 8340 7044 8396 7100
rect 8396 7044 8400 7100
rect 8336 7040 8400 7044
rect 8416 7100 8480 7104
rect 8416 7044 8420 7100
rect 8420 7044 8476 7100
rect 8476 7044 8480 7100
rect 8416 7040 8480 7044
rect 22624 7100 22688 7104
rect 22624 7044 22628 7100
rect 22628 7044 22684 7100
rect 22684 7044 22688 7100
rect 22624 7040 22688 7044
rect 22704 7100 22768 7104
rect 22704 7044 22708 7100
rect 22708 7044 22764 7100
rect 22764 7044 22768 7100
rect 22704 7040 22768 7044
rect 22784 7100 22848 7104
rect 22784 7044 22788 7100
rect 22788 7044 22844 7100
rect 22844 7044 22848 7100
rect 22784 7040 22848 7044
rect 22864 7100 22928 7104
rect 22864 7044 22868 7100
rect 22868 7044 22924 7100
rect 22924 7044 22928 7100
rect 22864 7040 22928 7044
rect 37072 7100 37136 7104
rect 37072 7044 37076 7100
rect 37076 7044 37132 7100
rect 37132 7044 37136 7100
rect 37072 7040 37136 7044
rect 37152 7100 37216 7104
rect 37152 7044 37156 7100
rect 37156 7044 37212 7100
rect 37212 7044 37216 7100
rect 37152 7040 37216 7044
rect 37232 7100 37296 7104
rect 37232 7044 37236 7100
rect 37236 7044 37292 7100
rect 37292 7044 37296 7100
rect 37232 7040 37296 7044
rect 37312 7100 37376 7104
rect 37312 7044 37316 7100
rect 37316 7044 37372 7100
rect 37372 7044 37376 7100
rect 37312 7040 37376 7044
rect 51520 7100 51584 7104
rect 51520 7044 51524 7100
rect 51524 7044 51580 7100
rect 51580 7044 51584 7100
rect 51520 7040 51584 7044
rect 51600 7100 51664 7104
rect 51600 7044 51604 7100
rect 51604 7044 51660 7100
rect 51660 7044 51664 7100
rect 51600 7040 51664 7044
rect 51680 7100 51744 7104
rect 51680 7044 51684 7100
rect 51684 7044 51740 7100
rect 51740 7044 51744 7100
rect 51680 7040 51744 7044
rect 51760 7100 51824 7104
rect 51760 7044 51764 7100
rect 51764 7044 51820 7100
rect 51820 7044 51824 7100
rect 51760 7040 51824 7044
rect 7972 6700 8036 6764
rect 17908 6700 17972 6764
rect 16436 6624 16500 6628
rect 16436 6568 16450 6624
rect 16450 6568 16500 6624
rect 16436 6564 16500 6568
rect 15400 6556 15464 6560
rect 15400 6500 15404 6556
rect 15404 6500 15460 6556
rect 15460 6500 15464 6556
rect 15400 6496 15464 6500
rect 15480 6556 15544 6560
rect 15480 6500 15484 6556
rect 15484 6500 15540 6556
rect 15540 6500 15544 6556
rect 15480 6496 15544 6500
rect 15560 6556 15624 6560
rect 15560 6500 15564 6556
rect 15564 6500 15620 6556
rect 15620 6500 15624 6556
rect 15560 6496 15624 6500
rect 15640 6556 15704 6560
rect 15640 6500 15644 6556
rect 15644 6500 15700 6556
rect 15700 6500 15704 6556
rect 15640 6496 15704 6500
rect 29848 6556 29912 6560
rect 29848 6500 29852 6556
rect 29852 6500 29908 6556
rect 29908 6500 29912 6556
rect 29848 6496 29912 6500
rect 29928 6556 29992 6560
rect 29928 6500 29932 6556
rect 29932 6500 29988 6556
rect 29988 6500 29992 6556
rect 29928 6496 29992 6500
rect 30008 6556 30072 6560
rect 30008 6500 30012 6556
rect 30012 6500 30068 6556
rect 30068 6500 30072 6556
rect 30008 6496 30072 6500
rect 30088 6556 30152 6560
rect 30088 6500 30092 6556
rect 30092 6500 30148 6556
rect 30148 6500 30152 6556
rect 30088 6496 30152 6500
rect 44296 6556 44360 6560
rect 44296 6500 44300 6556
rect 44300 6500 44356 6556
rect 44356 6500 44360 6556
rect 44296 6496 44360 6500
rect 44376 6556 44440 6560
rect 44376 6500 44380 6556
rect 44380 6500 44436 6556
rect 44436 6500 44440 6556
rect 44376 6496 44440 6500
rect 44456 6556 44520 6560
rect 44456 6500 44460 6556
rect 44460 6500 44516 6556
rect 44516 6500 44520 6556
rect 44456 6496 44520 6500
rect 44536 6556 44600 6560
rect 44536 6500 44540 6556
rect 44540 6500 44596 6556
rect 44596 6500 44600 6556
rect 44536 6496 44600 6500
rect 12204 6292 12268 6356
rect 18644 6216 18708 6220
rect 18644 6160 18694 6216
rect 18694 6160 18708 6216
rect 18644 6156 18708 6160
rect 9996 6020 10060 6084
rect 8176 6012 8240 6016
rect 8176 5956 8180 6012
rect 8180 5956 8236 6012
rect 8236 5956 8240 6012
rect 8176 5952 8240 5956
rect 8256 6012 8320 6016
rect 8256 5956 8260 6012
rect 8260 5956 8316 6012
rect 8316 5956 8320 6012
rect 8256 5952 8320 5956
rect 8336 6012 8400 6016
rect 8336 5956 8340 6012
rect 8340 5956 8396 6012
rect 8396 5956 8400 6012
rect 8336 5952 8400 5956
rect 8416 6012 8480 6016
rect 8416 5956 8420 6012
rect 8420 5956 8476 6012
rect 8476 5956 8480 6012
rect 8416 5952 8480 5956
rect 22624 6012 22688 6016
rect 22624 5956 22628 6012
rect 22628 5956 22684 6012
rect 22684 5956 22688 6012
rect 22624 5952 22688 5956
rect 22704 6012 22768 6016
rect 22704 5956 22708 6012
rect 22708 5956 22764 6012
rect 22764 5956 22768 6012
rect 22704 5952 22768 5956
rect 22784 6012 22848 6016
rect 22784 5956 22788 6012
rect 22788 5956 22844 6012
rect 22844 5956 22848 6012
rect 22784 5952 22848 5956
rect 22864 6012 22928 6016
rect 22864 5956 22868 6012
rect 22868 5956 22924 6012
rect 22924 5956 22928 6012
rect 22864 5952 22928 5956
rect 37072 6012 37136 6016
rect 37072 5956 37076 6012
rect 37076 5956 37132 6012
rect 37132 5956 37136 6012
rect 37072 5952 37136 5956
rect 37152 6012 37216 6016
rect 37152 5956 37156 6012
rect 37156 5956 37212 6012
rect 37212 5956 37216 6012
rect 37152 5952 37216 5956
rect 37232 6012 37296 6016
rect 37232 5956 37236 6012
rect 37236 5956 37292 6012
rect 37292 5956 37296 6012
rect 37232 5952 37296 5956
rect 37312 6012 37376 6016
rect 37312 5956 37316 6012
rect 37316 5956 37372 6012
rect 37372 5956 37376 6012
rect 37312 5952 37376 5956
rect 51520 6012 51584 6016
rect 51520 5956 51524 6012
rect 51524 5956 51580 6012
rect 51580 5956 51584 6012
rect 51520 5952 51584 5956
rect 51600 6012 51664 6016
rect 51600 5956 51604 6012
rect 51604 5956 51660 6012
rect 51660 5956 51664 6012
rect 51600 5952 51664 5956
rect 51680 6012 51744 6016
rect 51680 5956 51684 6012
rect 51684 5956 51740 6012
rect 51740 5956 51744 6012
rect 51680 5952 51744 5956
rect 51760 6012 51824 6016
rect 51760 5956 51764 6012
rect 51764 5956 51820 6012
rect 51820 5956 51824 6012
rect 51760 5952 51824 5956
rect 12204 5612 12268 5676
rect 12388 5612 12452 5676
rect 22324 5612 22388 5676
rect 23612 5612 23676 5676
rect 15400 5468 15464 5472
rect 15400 5412 15404 5468
rect 15404 5412 15460 5468
rect 15460 5412 15464 5468
rect 15400 5408 15464 5412
rect 15480 5468 15544 5472
rect 15480 5412 15484 5468
rect 15484 5412 15540 5468
rect 15540 5412 15544 5468
rect 15480 5408 15544 5412
rect 15560 5468 15624 5472
rect 15560 5412 15564 5468
rect 15564 5412 15620 5468
rect 15620 5412 15624 5468
rect 15560 5408 15624 5412
rect 15640 5468 15704 5472
rect 15640 5412 15644 5468
rect 15644 5412 15700 5468
rect 15700 5412 15704 5468
rect 15640 5408 15704 5412
rect 29848 5468 29912 5472
rect 29848 5412 29852 5468
rect 29852 5412 29908 5468
rect 29908 5412 29912 5468
rect 29848 5408 29912 5412
rect 29928 5468 29992 5472
rect 29928 5412 29932 5468
rect 29932 5412 29988 5468
rect 29988 5412 29992 5468
rect 29928 5408 29992 5412
rect 30008 5468 30072 5472
rect 30008 5412 30012 5468
rect 30012 5412 30068 5468
rect 30068 5412 30072 5468
rect 30008 5408 30072 5412
rect 30088 5468 30152 5472
rect 30088 5412 30092 5468
rect 30092 5412 30148 5468
rect 30148 5412 30152 5468
rect 30088 5408 30152 5412
rect 44296 5468 44360 5472
rect 44296 5412 44300 5468
rect 44300 5412 44356 5468
rect 44356 5412 44360 5468
rect 44296 5408 44360 5412
rect 44376 5468 44440 5472
rect 44376 5412 44380 5468
rect 44380 5412 44436 5468
rect 44436 5412 44440 5468
rect 44376 5408 44440 5412
rect 44456 5468 44520 5472
rect 44456 5412 44460 5468
rect 44460 5412 44516 5468
rect 44516 5412 44520 5468
rect 44456 5408 44520 5412
rect 44536 5468 44600 5472
rect 44536 5412 44540 5468
rect 44540 5412 44596 5468
rect 44596 5412 44600 5468
rect 44536 5408 44600 5412
rect 2820 5340 2884 5404
rect 1900 5204 1964 5268
rect 13492 5204 13556 5268
rect 16436 5068 16500 5132
rect 8176 4924 8240 4928
rect 8176 4868 8180 4924
rect 8180 4868 8236 4924
rect 8236 4868 8240 4924
rect 8176 4864 8240 4868
rect 8256 4924 8320 4928
rect 8256 4868 8260 4924
rect 8260 4868 8316 4924
rect 8316 4868 8320 4924
rect 8256 4864 8320 4868
rect 8336 4924 8400 4928
rect 8336 4868 8340 4924
rect 8340 4868 8396 4924
rect 8396 4868 8400 4924
rect 8336 4864 8400 4868
rect 8416 4924 8480 4928
rect 8416 4868 8420 4924
rect 8420 4868 8476 4924
rect 8476 4868 8480 4924
rect 8416 4864 8480 4868
rect 22624 4924 22688 4928
rect 22624 4868 22628 4924
rect 22628 4868 22684 4924
rect 22684 4868 22688 4924
rect 22624 4864 22688 4868
rect 22704 4924 22768 4928
rect 22704 4868 22708 4924
rect 22708 4868 22764 4924
rect 22764 4868 22768 4924
rect 22704 4864 22768 4868
rect 22784 4924 22848 4928
rect 22784 4868 22788 4924
rect 22788 4868 22844 4924
rect 22844 4868 22848 4924
rect 22784 4864 22848 4868
rect 22864 4924 22928 4928
rect 22864 4868 22868 4924
rect 22868 4868 22924 4924
rect 22924 4868 22928 4924
rect 22864 4864 22928 4868
rect 8892 4796 8956 4860
rect 10732 4796 10796 4860
rect 14780 4660 14844 4724
rect 22140 4660 22204 4724
rect 37072 4924 37136 4928
rect 37072 4868 37076 4924
rect 37076 4868 37132 4924
rect 37132 4868 37136 4924
rect 37072 4864 37136 4868
rect 37152 4924 37216 4928
rect 37152 4868 37156 4924
rect 37156 4868 37212 4924
rect 37212 4868 37216 4924
rect 37152 4864 37216 4868
rect 37232 4924 37296 4928
rect 37232 4868 37236 4924
rect 37236 4868 37292 4924
rect 37292 4868 37296 4924
rect 37232 4864 37296 4868
rect 37312 4924 37376 4928
rect 37312 4868 37316 4924
rect 37316 4868 37372 4924
rect 37372 4868 37376 4924
rect 37312 4864 37376 4868
rect 51520 4924 51584 4928
rect 51520 4868 51524 4924
rect 51524 4868 51580 4924
rect 51580 4868 51584 4924
rect 51520 4864 51584 4868
rect 51600 4924 51664 4928
rect 51600 4868 51604 4924
rect 51604 4868 51660 4924
rect 51660 4868 51664 4924
rect 51600 4864 51664 4868
rect 51680 4924 51744 4928
rect 51680 4868 51684 4924
rect 51684 4868 51740 4924
rect 51740 4868 51744 4924
rect 51680 4864 51744 4868
rect 51760 4924 51824 4928
rect 51760 4868 51764 4924
rect 51764 4868 51820 4924
rect 51820 4868 51824 4924
rect 51760 4864 51824 4868
rect 9076 4388 9140 4452
rect 15400 4380 15464 4384
rect 15400 4324 15404 4380
rect 15404 4324 15460 4380
rect 15460 4324 15464 4380
rect 15400 4320 15464 4324
rect 15480 4380 15544 4384
rect 15480 4324 15484 4380
rect 15484 4324 15540 4380
rect 15540 4324 15544 4380
rect 15480 4320 15544 4324
rect 15560 4380 15624 4384
rect 15560 4324 15564 4380
rect 15564 4324 15620 4380
rect 15620 4324 15624 4380
rect 15560 4320 15624 4324
rect 15640 4380 15704 4384
rect 15640 4324 15644 4380
rect 15644 4324 15700 4380
rect 15700 4324 15704 4380
rect 15640 4320 15704 4324
rect 29848 4380 29912 4384
rect 29848 4324 29852 4380
rect 29852 4324 29908 4380
rect 29908 4324 29912 4380
rect 29848 4320 29912 4324
rect 29928 4380 29992 4384
rect 29928 4324 29932 4380
rect 29932 4324 29988 4380
rect 29988 4324 29992 4380
rect 29928 4320 29992 4324
rect 30008 4380 30072 4384
rect 30008 4324 30012 4380
rect 30012 4324 30068 4380
rect 30068 4324 30072 4380
rect 30008 4320 30072 4324
rect 30088 4380 30152 4384
rect 30088 4324 30092 4380
rect 30092 4324 30148 4380
rect 30148 4324 30152 4380
rect 30088 4320 30152 4324
rect 44296 4380 44360 4384
rect 44296 4324 44300 4380
rect 44300 4324 44356 4380
rect 44356 4324 44360 4380
rect 44296 4320 44360 4324
rect 44376 4380 44440 4384
rect 44376 4324 44380 4380
rect 44380 4324 44436 4380
rect 44436 4324 44440 4380
rect 44376 4320 44440 4324
rect 44456 4380 44520 4384
rect 44456 4324 44460 4380
rect 44460 4324 44516 4380
rect 44516 4324 44520 4380
rect 44456 4320 44520 4324
rect 44536 4380 44600 4384
rect 44536 4324 44540 4380
rect 44540 4324 44596 4380
rect 44596 4324 44600 4380
rect 44536 4320 44600 4324
rect 1900 4252 1964 4316
rect 8892 4252 8956 4316
rect 16988 4252 17052 4316
rect 7604 4116 7668 4180
rect 6684 3904 6748 3908
rect 6684 3848 6698 3904
rect 6698 3848 6748 3904
rect 6684 3844 6748 3848
rect 8708 3904 8772 3908
rect 8708 3848 8722 3904
rect 8722 3848 8772 3904
rect 8708 3844 8772 3848
rect 13308 3980 13372 4044
rect 14596 3980 14660 4044
rect 19196 4040 19260 4044
rect 19196 3984 19210 4040
rect 19210 3984 19260 4040
rect 19196 3980 19260 3984
rect 23060 3904 23124 3908
rect 23060 3848 23074 3904
rect 23074 3848 23124 3904
rect 23060 3844 23124 3848
rect 35756 3904 35820 3908
rect 35756 3848 35770 3904
rect 35770 3848 35820 3904
rect 35756 3844 35820 3848
rect 8176 3836 8240 3840
rect 8176 3780 8180 3836
rect 8180 3780 8236 3836
rect 8236 3780 8240 3836
rect 8176 3776 8240 3780
rect 8256 3836 8320 3840
rect 8256 3780 8260 3836
rect 8260 3780 8316 3836
rect 8316 3780 8320 3836
rect 8256 3776 8320 3780
rect 8336 3836 8400 3840
rect 8336 3780 8340 3836
rect 8340 3780 8396 3836
rect 8396 3780 8400 3836
rect 8336 3776 8400 3780
rect 8416 3836 8480 3840
rect 8416 3780 8420 3836
rect 8420 3780 8476 3836
rect 8476 3780 8480 3836
rect 8416 3776 8480 3780
rect 22624 3836 22688 3840
rect 22624 3780 22628 3836
rect 22628 3780 22684 3836
rect 22684 3780 22688 3836
rect 22624 3776 22688 3780
rect 22704 3836 22768 3840
rect 22704 3780 22708 3836
rect 22708 3780 22764 3836
rect 22764 3780 22768 3836
rect 22704 3776 22768 3780
rect 22784 3836 22848 3840
rect 22784 3780 22788 3836
rect 22788 3780 22844 3836
rect 22844 3780 22848 3836
rect 22784 3776 22848 3780
rect 22864 3836 22928 3840
rect 22864 3780 22868 3836
rect 22868 3780 22924 3836
rect 22924 3780 22928 3836
rect 22864 3776 22928 3780
rect 37072 3836 37136 3840
rect 37072 3780 37076 3836
rect 37076 3780 37132 3836
rect 37132 3780 37136 3836
rect 37072 3776 37136 3780
rect 37152 3836 37216 3840
rect 37152 3780 37156 3836
rect 37156 3780 37212 3836
rect 37212 3780 37216 3836
rect 37152 3776 37216 3780
rect 37232 3836 37296 3840
rect 37232 3780 37236 3836
rect 37236 3780 37292 3836
rect 37292 3780 37296 3836
rect 37232 3776 37296 3780
rect 37312 3836 37376 3840
rect 37312 3780 37316 3836
rect 37316 3780 37372 3836
rect 37372 3780 37376 3836
rect 37312 3776 37376 3780
rect 51520 3836 51584 3840
rect 51520 3780 51524 3836
rect 51524 3780 51580 3836
rect 51580 3780 51584 3836
rect 51520 3776 51584 3780
rect 51600 3836 51664 3840
rect 51600 3780 51604 3836
rect 51604 3780 51660 3836
rect 51660 3780 51664 3836
rect 51600 3776 51664 3780
rect 51680 3836 51744 3840
rect 51680 3780 51684 3836
rect 51684 3780 51740 3836
rect 51740 3780 51744 3836
rect 51680 3776 51744 3780
rect 51760 3836 51824 3840
rect 51760 3780 51764 3836
rect 51764 3780 51820 3836
rect 51820 3780 51824 3836
rect 51760 3776 51824 3780
rect 7420 3768 7484 3772
rect 7420 3712 7470 3768
rect 7470 3712 7484 3768
rect 7420 3708 7484 3712
rect 9444 3708 9508 3772
rect 16436 3708 16500 3772
rect 16620 3708 16684 3772
rect 14780 3632 14844 3636
rect 14780 3576 14830 3632
rect 14830 3576 14844 3632
rect 14780 3572 14844 3576
rect 18276 3632 18340 3636
rect 18276 3576 18326 3632
rect 18326 3576 18340 3632
rect 18276 3572 18340 3576
rect 23428 3632 23492 3636
rect 23428 3576 23442 3632
rect 23442 3576 23492 3632
rect 23428 3572 23492 3576
rect 9996 3300 10060 3364
rect 16436 3300 16500 3364
rect 15400 3292 15464 3296
rect 15400 3236 15404 3292
rect 15404 3236 15460 3292
rect 15460 3236 15464 3292
rect 15400 3232 15464 3236
rect 15480 3292 15544 3296
rect 15480 3236 15484 3292
rect 15484 3236 15540 3292
rect 15540 3236 15544 3292
rect 15480 3232 15544 3236
rect 15560 3292 15624 3296
rect 15560 3236 15564 3292
rect 15564 3236 15620 3292
rect 15620 3236 15624 3292
rect 15560 3232 15624 3236
rect 15640 3292 15704 3296
rect 15640 3236 15644 3292
rect 15644 3236 15700 3292
rect 15700 3236 15704 3292
rect 15640 3232 15704 3236
rect 7420 3224 7484 3228
rect 7420 3168 7434 3224
rect 7434 3168 7484 3224
rect 7420 3164 7484 3168
rect 7972 3164 8036 3228
rect 29848 3292 29912 3296
rect 29848 3236 29852 3292
rect 29852 3236 29908 3292
rect 29908 3236 29912 3292
rect 29848 3232 29912 3236
rect 29928 3292 29992 3296
rect 29928 3236 29932 3292
rect 29932 3236 29988 3292
rect 29988 3236 29992 3292
rect 29928 3232 29992 3236
rect 30008 3292 30072 3296
rect 30008 3236 30012 3292
rect 30012 3236 30068 3292
rect 30068 3236 30072 3292
rect 30008 3232 30072 3236
rect 30088 3292 30152 3296
rect 30088 3236 30092 3292
rect 30092 3236 30148 3292
rect 30148 3236 30152 3292
rect 30088 3232 30152 3236
rect 44296 3292 44360 3296
rect 44296 3236 44300 3292
rect 44300 3236 44356 3292
rect 44356 3236 44360 3292
rect 44296 3232 44360 3236
rect 44376 3292 44440 3296
rect 44376 3236 44380 3292
rect 44380 3236 44436 3292
rect 44436 3236 44440 3292
rect 44376 3232 44440 3236
rect 44456 3292 44520 3296
rect 44456 3236 44460 3292
rect 44460 3236 44516 3292
rect 44516 3236 44520 3292
rect 44456 3232 44520 3236
rect 44536 3292 44600 3296
rect 44536 3236 44540 3292
rect 44540 3236 44596 3292
rect 44596 3236 44600 3292
rect 44536 3232 44600 3236
rect 23612 3164 23676 3228
rect 9260 2756 9324 2820
rect 8176 2748 8240 2752
rect 8176 2692 8180 2748
rect 8180 2692 8236 2748
rect 8236 2692 8240 2748
rect 8176 2688 8240 2692
rect 8256 2748 8320 2752
rect 8256 2692 8260 2748
rect 8260 2692 8316 2748
rect 8316 2692 8320 2748
rect 8256 2688 8320 2692
rect 8336 2748 8400 2752
rect 8336 2692 8340 2748
rect 8340 2692 8396 2748
rect 8396 2692 8400 2748
rect 8336 2688 8400 2692
rect 8416 2748 8480 2752
rect 8416 2692 8420 2748
rect 8420 2692 8476 2748
rect 8476 2692 8480 2748
rect 8416 2688 8480 2692
rect 15148 2892 15212 2956
rect 17908 2892 17972 2956
rect 12940 2756 13004 2820
rect 14964 2756 15028 2820
rect 22624 2748 22688 2752
rect 22624 2692 22628 2748
rect 22628 2692 22684 2748
rect 22684 2692 22688 2748
rect 22624 2688 22688 2692
rect 22704 2748 22768 2752
rect 22704 2692 22708 2748
rect 22708 2692 22764 2748
rect 22764 2692 22768 2748
rect 22704 2688 22768 2692
rect 22784 2748 22848 2752
rect 22784 2692 22788 2748
rect 22788 2692 22844 2748
rect 22844 2692 22848 2748
rect 22784 2688 22848 2692
rect 22864 2748 22928 2752
rect 22864 2692 22868 2748
rect 22868 2692 22924 2748
rect 22924 2692 22928 2748
rect 22864 2688 22928 2692
rect 37072 2748 37136 2752
rect 37072 2692 37076 2748
rect 37076 2692 37132 2748
rect 37132 2692 37136 2748
rect 37072 2688 37136 2692
rect 37152 2748 37216 2752
rect 37152 2692 37156 2748
rect 37156 2692 37212 2748
rect 37212 2692 37216 2748
rect 37152 2688 37216 2692
rect 37232 2748 37296 2752
rect 37232 2692 37236 2748
rect 37236 2692 37292 2748
rect 37292 2692 37296 2748
rect 37232 2688 37296 2692
rect 37312 2748 37376 2752
rect 37312 2692 37316 2748
rect 37316 2692 37372 2748
rect 37372 2692 37376 2748
rect 37312 2688 37376 2692
rect 51520 2748 51584 2752
rect 51520 2692 51524 2748
rect 51524 2692 51580 2748
rect 51580 2692 51584 2748
rect 51520 2688 51584 2692
rect 51600 2748 51664 2752
rect 51600 2692 51604 2748
rect 51604 2692 51660 2748
rect 51660 2692 51664 2748
rect 51600 2688 51664 2692
rect 51680 2748 51744 2752
rect 51680 2692 51684 2748
rect 51684 2692 51740 2748
rect 51740 2692 51744 2748
rect 51680 2688 51744 2692
rect 51760 2748 51824 2752
rect 51760 2692 51764 2748
rect 51764 2692 51820 2748
rect 51820 2692 51824 2748
rect 51760 2688 51824 2692
rect 4660 2620 4724 2684
rect 17724 2680 17788 2684
rect 17724 2624 17738 2680
rect 17738 2624 17788 2680
rect 17724 2620 17788 2624
rect 9444 2348 9508 2412
rect 7604 2212 7668 2276
rect 34468 2212 34532 2276
rect 15400 2204 15464 2208
rect 15400 2148 15404 2204
rect 15404 2148 15460 2204
rect 15460 2148 15464 2204
rect 15400 2144 15464 2148
rect 15480 2204 15544 2208
rect 15480 2148 15484 2204
rect 15484 2148 15540 2204
rect 15540 2148 15544 2204
rect 15480 2144 15544 2148
rect 15560 2204 15624 2208
rect 15560 2148 15564 2204
rect 15564 2148 15620 2204
rect 15620 2148 15624 2204
rect 15560 2144 15624 2148
rect 15640 2204 15704 2208
rect 15640 2148 15644 2204
rect 15644 2148 15700 2204
rect 15700 2148 15704 2204
rect 15640 2144 15704 2148
rect 29848 2204 29912 2208
rect 29848 2148 29852 2204
rect 29852 2148 29908 2204
rect 29908 2148 29912 2204
rect 29848 2144 29912 2148
rect 29928 2204 29992 2208
rect 29928 2148 29932 2204
rect 29932 2148 29988 2204
rect 29988 2148 29992 2204
rect 29928 2144 29992 2148
rect 30008 2204 30072 2208
rect 30008 2148 30012 2204
rect 30012 2148 30068 2204
rect 30068 2148 30072 2204
rect 30008 2144 30072 2148
rect 30088 2204 30152 2208
rect 30088 2148 30092 2204
rect 30092 2148 30148 2204
rect 30148 2148 30152 2204
rect 30088 2144 30152 2148
rect 44296 2204 44360 2208
rect 44296 2148 44300 2204
rect 44300 2148 44356 2204
rect 44356 2148 44360 2204
rect 44296 2144 44360 2148
rect 44376 2204 44440 2208
rect 44376 2148 44380 2204
rect 44380 2148 44436 2204
rect 44436 2148 44440 2204
rect 44376 2144 44440 2148
rect 44456 2204 44520 2208
rect 44456 2148 44460 2204
rect 44460 2148 44516 2204
rect 44516 2148 44520 2204
rect 44456 2144 44520 2148
rect 44536 2204 44600 2208
rect 44536 2148 44540 2204
rect 44540 2148 44596 2204
rect 44596 2148 44600 2204
rect 44536 2144 44600 2148
rect 8892 2076 8956 2140
rect 12204 1260 12268 1324
rect 34468 988 34532 1052
<< metal4 >>
rect 8168 16896 8488 17456
rect 8168 16832 8176 16896
rect 8240 16832 8256 16896
rect 8320 16832 8336 16896
rect 8400 16832 8416 16896
rect 8480 16832 8488 16896
rect 8168 15808 8488 16832
rect 8168 15744 8176 15808
rect 8240 15744 8256 15808
rect 8320 15744 8336 15808
rect 8400 15744 8416 15808
rect 8480 15744 8488 15808
rect 8168 14720 8488 15744
rect 8168 14656 8176 14720
rect 8240 14656 8256 14720
rect 8320 14656 8336 14720
rect 8400 14656 8416 14720
rect 8480 14656 8488 14720
rect 8168 13632 8488 14656
rect 15392 17440 15712 17456
rect 15392 17376 15400 17440
rect 15464 17376 15480 17440
rect 15544 17376 15560 17440
rect 15624 17376 15640 17440
rect 15704 17376 15712 17440
rect 15392 16352 15712 17376
rect 15392 16288 15400 16352
rect 15464 16288 15480 16352
rect 15544 16288 15560 16352
rect 15624 16288 15640 16352
rect 15704 16288 15712 16352
rect 15392 15264 15712 16288
rect 15392 15200 15400 15264
rect 15464 15200 15480 15264
rect 15544 15200 15560 15264
rect 15624 15200 15640 15264
rect 15704 15200 15712 15264
rect 15392 14176 15712 15200
rect 15392 14112 15400 14176
rect 15464 14112 15480 14176
rect 15544 14112 15560 14176
rect 15624 14112 15640 14176
rect 15704 14112 15712 14176
rect 13307 13836 13373 13837
rect 13307 13772 13308 13836
rect 13372 13772 13373 13836
rect 13307 13771 13373 13772
rect 8168 13568 8176 13632
rect 8240 13568 8256 13632
rect 8320 13568 8336 13632
rect 8400 13568 8416 13632
rect 8480 13568 8488 13632
rect 8168 12544 8488 13568
rect 10731 12748 10797 12749
rect 10731 12684 10732 12748
rect 10796 12684 10797 12748
rect 10731 12683 10797 12684
rect 8168 12480 8176 12544
rect 8240 12480 8256 12544
rect 8320 12480 8336 12544
rect 8400 12480 8416 12544
rect 8480 12480 8488 12544
rect 1899 12476 1965 12477
rect 1899 12412 1900 12476
rect 1964 12412 1965 12476
rect 1899 12411 1965 12412
rect 2819 12476 2885 12477
rect 2819 12412 2820 12476
rect 2884 12412 2885 12476
rect 2819 12411 2885 12412
rect 6683 12476 6749 12477
rect 6683 12412 6684 12476
rect 6748 12412 6749 12476
rect 6683 12411 6749 12412
rect 1902 5269 1962 12411
rect 2822 5405 2882 12411
rect 5947 11524 6013 11525
rect 5947 11460 5948 11524
rect 6012 11460 6013 11524
rect 5947 11459 6013 11460
rect 4659 11116 4725 11117
rect 4659 11052 4660 11116
rect 4724 11052 4725 11116
rect 4659 11051 4725 11052
rect 2819 5404 2885 5405
rect 2819 5340 2820 5404
rect 2884 5340 2885 5404
rect 2819 5339 2885 5340
rect 1899 5268 1965 5269
rect 1899 5204 1900 5268
rect 1964 5204 1965 5268
rect 1899 5203 1965 5204
rect 1902 4317 1962 5203
rect 1899 4316 1965 4317
rect 1899 4252 1900 4316
rect 1964 4252 1965 4316
rect 1899 4251 1965 4252
rect 4662 2685 4722 11051
rect 5950 7581 6010 11459
rect 5947 7580 6013 7581
rect 5947 7516 5948 7580
rect 6012 7516 6013 7580
rect 5947 7515 6013 7516
rect 6686 3909 6746 12411
rect 8168 11456 8488 12480
rect 8168 11392 8176 11456
rect 8240 11392 8256 11456
rect 8320 11392 8336 11456
rect 8400 11392 8416 11456
rect 8480 11392 8488 11456
rect 8168 10368 8488 11392
rect 9259 10572 9325 10573
rect 9259 10508 9260 10572
rect 9324 10508 9325 10572
rect 9259 10507 9325 10508
rect 8168 10304 8176 10368
rect 8240 10304 8256 10368
rect 8320 10304 8336 10368
rect 8400 10304 8416 10368
rect 8480 10304 8488 10368
rect 8168 9280 8488 10304
rect 9075 10028 9141 10029
rect 9075 9964 9076 10028
rect 9140 9964 9141 10028
rect 9075 9963 9141 9964
rect 8891 9892 8957 9893
rect 8891 9828 8892 9892
rect 8956 9828 8957 9892
rect 8891 9827 8957 9828
rect 8707 9756 8773 9757
rect 8707 9692 8708 9756
rect 8772 9692 8773 9756
rect 8707 9691 8773 9692
rect 8168 9216 8176 9280
rect 8240 9216 8256 9280
rect 8320 9216 8336 9280
rect 8400 9216 8416 9280
rect 8480 9216 8488 9280
rect 8168 8192 8488 9216
rect 8168 8128 8176 8192
rect 8240 8128 8256 8192
rect 8320 8128 8336 8192
rect 8400 8128 8416 8192
rect 8480 8128 8488 8192
rect 8168 7104 8488 8128
rect 8168 7040 8176 7104
rect 8240 7040 8256 7104
rect 8320 7040 8336 7104
rect 8400 7040 8416 7104
rect 8480 7040 8488 7104
rect 7971 6764 8037 6765
rect 7971 6700 7972 6764
rect 8036 6700 8037 6764
rect 7971 6699 8037 6700
rect 7603 4180 7669 4181
rect 7603 4116 7604 4180
rect 7668 4116 7669 4180
rect 7603 4115 7669 4116
rect 6683 3908 6749 3909
rect 6683 3844 6684 3908
rect 6748 3844 6749 3908
rect 6683 3843 6749 3844
rect 7419 3772 7485 3773
rect 7419 3708 7420 3772
rect 7484 3708 7485 3772
rect 7419 3707 7485 3708
rect 7422 3229 7482 3707
rect 7419 3228 7485 3229
rect 7419 3164 7420 3228
rect 7484 3164 7485 3228
rect 7419 3163 7485 3164
rect 4659 2684 4725 2685
rect 4659 2620 4660 2684
rect 4724 2620 4725 2684
rect 4659 2619 4725 2620
rect 7606 2277 7666 4115
rect 7974 3229 8034 6699
rect 8168 6016 8488 7040
rect 8168 5952 8176 6016
rect 8240 5952 8256 6016
rect 8320 5952 8336 6016
rect 8400 5952 8416 6016
rect 8480 5952 8488 6016
rect 8168 4928 8488 5952
rect 8168 4864 8176 4928
rect 8240 4864 8256 4928
rect 8320 4864 8336 4928
rect 8400 4864 8416 4928
rect 8480 4864 8488 4928
rect 8168 3840 8488 4864
rect 8710 3909 8770 9691
rect 8894 4861 8954 9827
rect 8891 4860 8957 4861
rect 8891 4796 8892 4860
rect 8956 4796 8957 4860
rect 8891 4795 8957 4796
rect 9078 4453 9138 9963
rect 9075 4452 9141 4453
rect 9075 4388 9076 4452
rect 9140 4388 9141 4452
rect 9075 4387 9141 4388
rect 8891 4316 8957 4317
rect 8891 4252 8892 4316
rect 8956 4252 8957 4316
rect 8891 4251 8957 4252
rect 8707 3908 8773 3909
rect 8707 3844 8708 3908
rect 8772 3844 8773 3908
rect 8707 3843 8773 3844
rect 8168 3776 8176 3840
rect 8240 3776 8256 3840
rect 8320 3776 8336 3840
rect 8400 3776 8416 3840
rect 8480 3776 8488 3840
rect 7971 3228 8037 3229
rect 7971 3164 7972 3228
rect 8036 3164 8037 3228
rect 7971 3163 8037 3164
rect 8168 2752 8488 3776
rect 8168 2688 8176 2752
rect 8240 2688 8256 2752
rect 8320 2688 8336 2752
rect 8400 2688 8416 2752
rect 8480 2688 8488 2752
rect 7603 2276 7669 2277
rect 7603 2212 7604 2276
rect 7668 2212 7669 2276
rect 7603 2211 7669 2212
rect 8168 2128 8488 2688
rect 8894 2141 8954 4251
rect 9262 2821 9322 10507
rect 9995 6084 10061 6085
rect 9995 6020 9996 6084
rect 10060 6020 10061 6084
rect 9995 6019 10061 6020
rect 9443 3772 9509 3773
rect 9443 3708 9444 3772
rect 9508 3708 9509 3772
rect 9443 3707 9509 3708
rect 9259 2820 9325 2821
rect 9259 2756 9260 2820
rect 9324 2756 9325 2820
rect 9259 2755 9325 2756
rect 9446 2413 9506 3707
rect 9998 3365 10058 6019
rect 10734 4861 10794 12683
rect 10915 12612 10981 12613
rect 10915 12548 10916 12612
rect 10980 12548 10981 12612
rect 10915 12547 10981 12548
rect 10918 10029 10978 12547
rect 12939 11252 13005 11253
rect 12939 11188 12940 11252
rect 13004 11188 13005 11252
rect 12939 11187 13005 11188
rect 10915 10028 10981 10029
rect 10915 9964 10916 10028
rect 10980 9964 10981 10028
rect 10915 9963 10981 9964
rect 12203 6356 12269 6357
rect 12203 6292 12204 6356
rect 12268 6292 12269 6356
rect 12203 6291 12269 6292
rect 12206 5810 12266 6291
rect 12206 5750 12450 5810
rect 12390 5677 12450 5750
rect 12203 5676 12269 5677
rect 12203 5612 12204 5676
rect 12268 5612 12269 5676
rect 12203 5611 12269 5612
rect 12387 5676 12453 5677
rect 12387 5612 12388 5676
rect 12452 5612 12453 5676
rect 12387 5611 12453 5612
rect 10731 4860 10797 4861
rect 10731 4796 10732 4860
rect 10796 4796 10797 4860
rect 10731 4795 10797 4796
rect 9995 3364 10061 3365
rect 9995 3300 9996 3364
rect 10060 3300 10061 3364
rect 9995 3299 10061 3300
rect 9443 2412 9509 2413
rect 9443 2348 9444 2412
rect 9508 2348 9509 2412
rect 9443 2347 9509 2348
rect 8891 2140 8957 2141
rect 8891 2076 8892 2140
rect 8956 2076 8957 2140
rect 8891 2075 8957 2076
rect 12206 1325 12266 5611
rect 12942 2821 13002 11187
rect 13310 4045 13370 13771
rect 15392 13088 15712 14112
rect 22616 16896 22936 17456
rect 22616 16832 22624 16896
rect 22688 16832 22704 16896
rect 22768 16832 22784 16896
rect 22848 16832 22864 16896
rect 22928 16832 22936 16896
rect 22616 15808 22936 16832
rect 22616 15744 22624 15808
rect 22688 15744 22704 15808
rect 22768 15744 22784 15808
rect 22848 15744 22864 15808
rect 22928 15744 22936 15808
rect 22616 14720 22936 15744
rect 22616 14656 22624 14720
rect 22688 14656 22704 14720
rect 22768 14656 22784 14720
rect 22848 14656 22864 14720
rect 22928 14656 22936 14720
rect 22616 13632 22936 14656
rect 22616 13568 22624 13632
rect 22688 13568 22704 13632
rect 22768 13568 22784 13632
rect 22848 13568 22864 13632
rect 22928 13568 22936 13632
rect 17723 13156 17789 13157
rect 17723 13092 17724 13156
rect 17788 13092 17789 13156
rect 17723 13091 17789 13092
rect 15392 13024 15400 13088
rect 15464 13024 15480 13088
rect 15544 13024 15560 13088
rect 15624 13024 15640 13088
rect 15704 13024 15712 13088
rect 14595 12748 14661 12749
rect 14595 12684 14596 12748
rect 14660 12684 14661 12748
rect 14595 12683 14661 12684
rect 14227 12068 14293 12069
rect 14227 12004 14228 12068
rect 14292 12004 14293 12068
rect 14227 12003 14293 12004
rect 14230 7989 14290 12003
rect 14598 11797 14658 12683
rect 15392 12000 15712 13024
rect 16987 12476 17053 12477
rect 16987 12412 16988 12476
rect 17052 12412 17053 12476
rect 16987 12411 17053 12412
rect 15392 11936 15400 12000
rect 15464 11936 15480 12000
rect 15544 11936 15560 12000
rect 15624 11936 15640 12000
rect 15704 11936 15712 12000
rect 14595 11796 14661 11797
rect 14595 11732 14596 11796
rect 14660 11732 14661 11796
rect 14595 11731 14661 11732
rect 13491 7988 13557 7989
rect 13491 7924 13492 7988
rect 13556 7924 13557 7988
rect 13491 7923 13557 7924
rect 14227 7988 14293 7989
rect 14227 7924 14228 7988
rect 14292 7924 14293 7988
rect 14227 7923 14293 7924
rect 13494 5269 13554 7923
rect 14230 7309 14290 7923
rect 14227 7308 14293 7309
rect 14227 7244 14228 7308
rect 14292 7244 14293 7308
rect 14227 7243 14293 7244
rect 13491 5268 13557 5269
rect 13491 5204 13492 5268
rect 13556 5204 13557 5268
rect 13491 5203 13557 5204
rect 14598 4045 14658 11731
rect 15147 11116 15213 11117
rect 15147 11052 15148 11116
rect 15212 11052 15213 11116
rect 15147 11051 15213 11052
rect 14963 7852 15029 7853
rect 14963 7788 14964 7852
rect 15028 7788 15029 7852
rect 14963 7787 15029 7788
rect 14779 4724 14845 4725
rect 14779 4660 14780 4724
rect 14844 4660 14845 4724
rect 14779 4659 14845 4660
rect 13307 4044 13373 4045
rect 13307 3980 13308 4044
rect 13372 3980 13373 4044
rect 13307 3979 13373 3980
rect 14595 4044 14661 4045
rect 14595 3980 14596 4044
rect 14660 3980 14661 4044
rect 14595 3979 14661 3980
rect 14782 3637 14842 4659
rect 14779 3636 14845 3637
rect 14779 3572 14780 3636
rect 14844 3572 14845 3636
rect 14779 3571 14845 3572
rect 14966 2821 15026 7787
rect 15150 2957 15210 11051
rect 15392 10912 15712 11936
rect 15392 10848 15400 10912
rect 15464 10848 15480 10912
rect 15544 10848 15560 10912
rect 15624 10848 15640 10912
rect 15704 10848 15712 10912
rect 15392 9824 15712 10848
rect 16619 10164 16685 10165
rect 16619 10100 16620 10164
rect 16684 10100 16685 10164
rect 16619 10099 16685 10100
rect 15392 9760 15400 9824
rect 15464 9760 15480 9824
rect 15544 9760 15560 9824
rect 15624 9760 15640 9824
rect 15704 9760 15712 9824
rect 15392 8736 15712 9760
rect 15392 8672 15400 8736
rect 15464 8672 15480 8736
rect 15544 8672 15560 8736
rect 15624 8672 15640 8736
rect 15704 8672 15712 8736
rect 15392 7648 15712 8672
rect 15392 7584 15400 7648
rect 15464 7584 15480 7648
rect 15544 7584 15560 7648
rect 15624 7584 15640 7648
rect 15704 7584 15712 7648
rect 15392 6560 15712 7584
rect 16435 6628 16501 6629
rect 16435 6564 16436 6628
rect 16500 6564 16501 6628
rect 16435 6563 16501 6564
rect 15392 6496 15400 6560
rect 15464 6496 15480 6560
rect 15544 6496 15560 6560
rect 15624 6496 15640 6560
rect 15704 6496 15712 6560
rect 15392 5472 15712 6496
rect 15392 5408 15400 5472
rect 15464 5408 15480 5472
rect 15544 5408 15560 5472
rect 15624 5408 15640 5472
rect 15704 5408 15712 5472
rect 15392 4384 15712 5408
rect 16438 5133 16498 6563
rect 16435 5132 16501 5133
rect 16435 5068 16436 5132
rect 16500 5068 16501 5132
rect 16435 5067 16501 5068
rect 15392 4320 15400 4384
rect 15464 4320 15480 4384
rect 15544 4320 15560 4384
rect 15624 4320 15640 4384
rect 15704 4320 15712 4384
rect 15392 3296 15712 4320
rect 16622 3773 16682 10099
rect 16990 4317 17050 12411
rect 17726 8261 17786 13091
rect 19195 12612 19261 12613
rect 19195 12548 19196 12612
rect 19260 12548 19261 12612
rect 19195 12547 19261 12548
rect 18643 12068 18709 12069
rect 18643 12004 18644 12068
rect 18708 12004 18709 12068
rect 18643 12003 18709 12004
rect 18275 11116 18341 11117
rect 18275 11052 18276 11116
rect 18340 11052 18341 11116
rect 18275 11051 18341 11052
rect 17723 8260 17789 8261
rect 17723 8196 17724 8260
rect 17788 8196 17789 8260
rect 17723 8195 17789 8196
rect 16987 4316 17053 4317
rect 16987 4252 16988 4316
rect 17052 4252 17053 4316
rect 16987 4251 17053 4252
rect 16435 3772 16501 3773
rect 16435 3708 16436 3772
rect 16500 3708 16501 3772
rect 16435 3707 16501 3708
rect 16619 3772 16685 3773
rect 16619 3708 16620 3772
rect 16684 3708 16685 3772
rect 16619 3707 16685 3708
rect 16438 3365 16498 3707
rect 16435 3364 16501 3365
rect 16435 3300 16436 3364
rect 16500 3300 16501 3364
rect 16435 3299 16501 3300
rect 15392 3232 15400 3296
rect 15464 3232 15480 3296
rect 15544 3232 15560 3296
rect 15624 3232 15640 3296
rect 15704 3232 15712 3296
rect 15147 2956 15213 2957
rect 15147 2892 15148 2956
rect 15212 2892 15213 2956
rect 15147 2891 15213 2892
rect 12939 2820 13005 2821
rect 12939 2756 12940 2820
rect 13004 2756 13005 2820
rect 12939 2755 13005 2756
rect 14963 2820 15029 2821
rect 14963 2756 14964 2820
rect 15028 2756 15029 2820
rect 14963 2755 15029 2756
rect 15392 2208 15712 3232
rect 17726 2685 17786 8195
rect 17907 6764 17973 6765
rect 17907 6700 17908 6764
rect 17972 6700 17973 6764
rect 17907 6699 17973 6700
rect 17910 2957 17970 6699
rect 18278 3637 18338 11051
rect 18646 6221 18706 12003
rect 18643 6220 18709 6221
rect 18643 6156 18644 6220
rect 18708 6156 18709 6220
rect 18643 6155 18709 6156
rect 19198 4045 19258 12547
rect 22616 12544 22936 13568
rect 22616 12480 22624 12544
rect 22688 12480 22704 12544
rect 22768 12480 22784 12544
rect 22848 12480 22864 12544
rect 22928 12480 22936 12544
rect 22323 12068 22389 12069
rect 22323 12004 22324 12068
rect 22388 12004 22389 12068
rect 22323 12003 22389 12004
rect 22139 11524 22205 11525
rect 22139 11460 22140 11524
rect 22204 11460 22205 11524
rect 22139 11459 22205 11460
rect 22142 4725 22202 11459
rect 22326 5677 22386 12003
rect 22616 11456 22936 12480
rect 29840 17440 30160 17456
rect 29840 17376 29848 17440
rect 29912 17376 29928 17440
rect 29992 17376 30008 17440
rect 30072 17376 30088 17440
rect 30152 17376 30160 17440
rect 29840 16352 30160 17376
rect 29840 16288 29848 16352
rect 29912 16288 29928 16352
rect 29992 16288 30008 16352
rect 30072 16288 30088 16352
rect 30152 16288 30160 16352
rect 29840 15264 30160 16288
rect 29840 15200 29848 15264
rect 29912 15200 29928 15264
rect 29992 15200 30008 15264
rect 30072 15200 30088 15264
rect 30152 15200 30160 15264
rect 29840 14176 30160 15200
rect 29840 14112 29848 14176
rect 29912 14112 29928 14176
rect 29992 14112 30008 14176
rect 30072 14112 30088 14176
rect 30152 14112 30160 14176
rect 29840 13088 30160 14112
rect 29840 13024 29848 13088
rect 29912 13024 29928 13088
rect 29992 13024 30008 13088
rect 30072 13024 30088 13088
rect 30152 13024 30160 13088
rect 23427 12476 23493 12477
rect 23427 12412 23428 12476
rect 23492 12412 23493 12476
rect 23427 12411 23493 12412
rect 22616 11392 22624 11456
rect 22688 11392 22704 11456
rect 22768 11392 22784 11456
rect 22848 11392 22864 11456
rect 22928 11392 22936 11456
rect 22616 10368 22936 11392
rect 23059 11116 23125 11117
rect 23059 11052 23060 11116
rect 23124 11052 23125 11116
rect 23059 11051 23125 11052
rect 22616 10304 22624 10368
rect 22688 10304 22704 10368
rect 22768 10304 22784 10368
rect 22848 10304 22864 10368
rect 22928 10304 22936 10368
rect 22616 9280 22936 10304
rect 22616 9216 22624 9280
rect 22688 9216 22704 9280
rect 22768 9216 22784 9280
rect 22848 9216 22864 9280
rect 22928 9216 22936 9280
rect 22616 8192 22936 9216
rect 22616 8128 22624 8192
rect 22688 8128 22704 8192
rect 22768 8128 22784 8192
rect 22848 8128 22864 8192
rect 22928 8128 22936 8192
rect 22616 7104 22936 8128
rect 22616 7040 22624 7104
rect 22688 7040 22704 7104
rect 22768 7040 22784 7104
rect 22848 7040 22864 7104
rect 22928 7040 22936 7104
rect 22616 6016 22936 7040
rect 22616 5952 22624 6016
rect 22688 5952 22704 6016
rect 22768 5952 22784 6016
rect 22848 5952 22864 6016
rect 22928 5952 22936 6016
rect 22323 5676 22389 5677
rect 22323 5612 22324 5676
rect 22388 5612 22389 5676
rect 22323 5611 22389 5612
rect 22616 4928 22936 5952
rect 22616 4864 22624 4928
rect 22688 4864 22704 4928
rect 22768 4864 22784 4928
rect 22848 4864 22864 4928
rect 22928 4864 22936 4928
rect 22139 4724 22205 4725
rect 22139 4660 22140 4724
rect 22204 4660 22205 4724
rect 22139 4659 22205 4660
rect 19195 4044 19261 4045
rect 19195 3980 19196 4044
rect 19260 3980 19261 4044
rect 19195 3979 19261 3980
rect 22616 3840 22936 4864
rect 23062 3909 23122 11051
rect 23059 3908 23125 3909
rect 23059 3844 23060 3908
rect 23124 3844 23125 3908
rect 23059 3843 23125 3844
rect 22616 3776 22624 3840
rect 22688 3776 22704 3840
rect 22768 3776 22784 3840
rect 22848 3776 22864 3840
rect 22928 3776 22936 3840
rect 18275 3636 18341 3637
rect 18275 3572 18276 3636
rect 18340 3572 18341 3636
rect 18275 3571 18341 3572
rect 17907 2956 17973 2957
rect 17907 2892 17908 2956
rect 17972 2892 17973 2956
rect 17907 2891 17973 2892
rect 22616 2752 22936 3776
rect 23430 3637 23490 12411
rect 29840 12000 30160 13024
rect 29840 11936 29848 12000
rect 29912 11936 29928 12000
rect 29992 11936 30008 12000
rect 30072 11936 30088 12000
rect 30152 11936 30160 12000
rect 29840 10912 30160 11936
rect 37064 16896 37384 17456
rect 37064 16832 37072 16896
rect 37136 16832 37152 16896
rect 37216 16832 37232 16896
rect 37296 16832 37312 16896
rect 37376 16832 37384 16896
rect 37064 15808 37384 16832
rect 37064 15744 37072 15808
rect 37136 15744 37152 15808
rect 37216 15744 37232 15808
rect 37296 15744 37312 15808
rect 37376 15744 37384 15808
rect 37064 14720 37384 15744
rect 37064 14656 37072 14720
rect 37136 14656 37152 14720
rect 37216 14656 37232 14720
rect 37296 14656 37312 14720
rect 37376 14656 37384 14720
rect 37064 13632 37384 14656
rect 37064 13568 37072 13632
rect 37136 13568 37152 13632
rect 37216 13568 37232 13632
rect 37296 13568 37312 13632
rect 37376 13568 37384 13632
rect 37064 12544 37384 13568
rect 37064 12480 37072 12544
rect 37136 12480 37152 12544
rect 37216 12480 37232 12544
rect 37296 12480 37312 12544
rect 37376 12480 37384 12544
rect 37064 11456 37384 12480
rect 37064 11392 37072 11456
rect 37136 11392 37152 11456
rect 37216 11392 37232 11456
rect 37296 11392 37312 11456
rect 37376 11392 37384 11456
rect 35755 11116 35821 11117
rect 35755 11052 35756 11116
rect 35820 11052 35821 11116
rect 35755 11051 35821 11052
rect 29840 10848 29848 10912
rect 29912 10848 29928 10912
rect 29992 10848 30008 10912
rect 30072 10848 30088 10912
rect 30152 10848 30160 10912
rect 29840 9824 30160 10848
rect 29840 9760 29848 9824
rect 29912 9760 29928 9824
rect 29992 9760 30008 9824
rect 30072 9760 30088 9824
rect 30152 9760 30160 9824
rect 29840 8736 30160 9760
rect 29840 8672 29848 8736
rect 29912 8672 29928 8736
rect 29992 8672 30008 8736
rect 30072 8672 30088 8736
rect 30152 8672 30160 8736
rect 29840 7648 30160 8672
rect 29840 7584 29848 7648
rect 29912 7584 29928 7648
rect 29992 7584 30008 7648
rect 30072 7584 30088 7648
rect 30152 7584 30160 7648
rect 29840 6560 30160 7584
rect 29840 6496 29848 6560
rect 29912 6496 29928 6560
rect 29992 6496 30008 6560
rect 30072 6496 30088 6560
rect 30152 6496 30160 6560
rect 23611 5676 23677 5677
rect 23611 5612 23612 5676
rect 23676 5612 23677 5676
rect 23611 5611 23677 5612
rect 23427 3636 23493 3637
rect 23427 3572 23428 3636
rect 23492 3572 23493 3636
rect 23427 3571 23493 3572
rect 23614 3229 23674 5611
rect 29840 5472 30160 6496
rect 29840 5408 29848 5472
rect 29912 5408 29928 5472
rect 29992 5408 30008 5472
rect 30072 5408 30088 5472
rect 30152 5408 30160 5472
rect 29840 4384 30160 5408
rect 29840 4320 29848 4384
rect 29912 4320 29928 4384
rect 29992 4320 30008 4384
rect 30072 4320 30088 4384
rect 30152 4320 30160 4384
rect 29840 3296 30160 4320
rect 35758 3909 35818 11051
rect 37064 10368 37384 11392
rect 37064 10304 37072 10368
rect 37136 10304 37152 10368
rect 37216 10304 37232 10368
rect 37296 10304 37312 10368
rect 37376 10304 37384 10368
rect 37064 9280 37384 10304
rect 37064 9216 37072 9280
rect 37136 9216 37152 9280
rect 37216 9216 37232 9280
rect 37296 9216 37312 9280
rect 37376 9216 37384 9280
rect 37064 8192 37384 9216
rect 37064 8128 37072 8192
rect 37136 8128 37152 8192
rect 37216 8128 37232 8192
rect 37296 8128 37312 8192
rect 37376 8128 37384 8192
rect 37064 7104 37384 8128
rect 37064 7040 37072 7104
rect 37136 7040 37152 7104
rect 37216 7040 37232 7104
rect 37296 7040 37312 7104
rect 37376 7040 37384 7104
rect 37064 6016 37384 7040
rect 37064 5952 37072 6016
rect 37136 5952 37152 6016
rect 37216 5952 37232 6016
rect 37296 5952 37312 6016
rect 37376 5952 37384 6016
rect 37064 4928 37384 5952
rect 37064 4864 37072 4928
rect 37136 4864 37152 4928
rect 37216 4864 37232 4928
rect 37296 4864 37312 4928
rect 37376 4864 37384 4928
rect 35755 3908 35821 3909
rect 35755 3844 35756 3908
rect 35820 3844 35821 3908
rect 35755 3843 35821 3844
rect 29840 3232 29848 3296
rect 29912 3232 29928 3296
rect 29992 3232 30008 3296
rect 30072 3232 30088 3296
rect 30152 3232 30160 3296
rect 23611 3228 23677 3229
rect 23611 3164 23612 3228
rect 23676 3164 23677 3228
rect 23611 3163 23677 3164
rect 22616 2688 22624 2752
rect 22688 2688 22704 2752
rect 22768 2688 22784 2752
rect 22848 2688 22864 2752
rect 22928 2688 22936 2752
rect 17723 2684 17789 2685
rect 17723 2620 17724 2684
rect 17788 2620 17789 2684
rect 17723 2619 17789 2620
rect 15392 2144 15400 2208
rect 15464 2144 15480 2208
rect 15544 2144 15560 2208
rect 15624 2144 15640 2208
rect 15704 2144 15712 2208
rect 15392 2128 15712 2144
rect 22616 2128 22936 2688
rect 29840 2208 30160 3232
rect 37064 3840 37384 4864
rect 37064 3776 37072 3840
rect 37136 3776 37152 3840
rect 37216 3776 37232 3840
rect 37296 3776 37312 3840
rect 37376 3776 37384 3840
rect 37064 2752 37384 3776
rect 37064 2688 37072 2752
rect 37136 2688 37152 2752
rect 37216 2688 37232 2752
rect 37296 2688 37312 2752
rect 37376 2688 37384 2752
rect 34467 2276 34533 2277
rect 34467 2212 34468 2276
rect 34532 2212 34533 2276
rect 34467 2211 34533 2212
rect 29840 2144 29848 2208
rect 29912 2144 29928 2208
rect 29992 2144 30008 2208
rect 30072 2144 30088 2208
rect 30152 2144 30160 2208
rect 29840 2128 30160 2144
rect 12203 1324 12269 1325
rect 12203 1260 12204 1324
rect 12268 1260 12269 1324
rect 12203 1259 12269 1260
rect 34470 1053 34530 2211
rect 37064 2128 37384 2688
rect 44288 17440 44608 17456
rect 44288 17376 44296 17440
rect 44360 17376 44376 17440
rect 44440 17376 44456 17440
rect 44520 17376 44536 17440
rect 44600 17376 44608 17440
rect 44288 16352 44608 17376
rect 44288 16288 44296 16352
rect 44360 16288 44376 16352
rect 44440 16288 44456 16352
rect 44520 16288 44536 16352
rect 44600 16288 44608 16352
rect 44288 15264 44608 16288
rect 44288 15200 44296 15264
rect 44360 15200 44376 15264
rect 44440 15200 44456 15264
rect 44520 15200 44536 15264
rect 44600 15200 44608 15264
rect 44288 14176 44608 15200
rect 44288 14112 44296 14176
rect 44360 14112 44376 14176
rect 44440 14112 44456 14176
rect 44520 14112 44536 14176
rect 44600 14112 44608 14176
rect 44288 13088 44608 14112
rect 44288 13024 44296 13088
rect 44360 13024 44376 13088
rect 44440 13024 44456 13088
rect 44520 13024 44536 13088
rect 44600 13024 44608 13088
rect 44288 12000 44608 13024
rect 44288 11936 44296 12000
rect 44360 11936 44376 12000
rect 44440 11936 44456 12000
rect 44520 11936 44536 12000
rect 44600 11936 44608 12000
rect 44288 10912 44608 11936
rect 44288 10848 44296 10912
rect 44360 10848 44376 10912
rect 44440 10848 44456 10912
rect 44520 10848 44536 10912
rect 44600 10848 44608 10912
rect 44288 9824 44608 10848
rect 44288 9760 44296 9824
rect 44360 9760 44376 9824
rect 44440 9760 44456 9824
rect 44520 9760 44536 9824
rect 44600 9760 44608 9824
rect 44288 8736 44608 9760
rect 44288 8672 44296 8736
rect 44360 8672 44376 8736
rect 44440 8672 44456 8736
rect 44520 8672 44536 8736
rect 44600 8672 44608 8736
rect 44288 7648 44608 8672
rect 44288 7584 44296 7648
rect 44360 7584 44376 7648
rect 44440 7584 44456 7648
rect 44520 7584 44536 7648
rect 44600 7584 44608 7648
rect 44288 6560 44608 7584
rect 44288 6496 44296 6560
rect 44360 6496 44376 6560
rect 44440 6496 44456 6560
rect 44520 6496 44536 6560
rect 44600 6496 44608 6560
rect 44288 5472 44608 6496
rect 44288 5408 44296 5472
rect 44360 5408 44376 5472
rect 44440 5408 44456 5472
rect 44520 5408 44536 5472
rect 44600 5408 44608 5472
rect 44288 4384 44608 5408
rect 44288 4320 44296 4384
rect 44360 4320 44376 4384
rect 44440 4320 44456 4384
rect 44520 4320 44536 4384
rect 44600 4320 44608 4384
rect 44288 3296 44608 4320
rect 44288 3232 44296 3296
rect 44360 3232 44376 3296
rect 44440 3232 44456 3296
rect 44520 3232 44536 3296
rect 44600 3232 44608 3296
rect 44288 2208 44608 3232
rect 44288 2144 44296 2208
rect 44360 2144 44376 2208
rect 44440 2144 44456 2208
rect 44520 2144 44536 2208
rect 44600 2144 44608 2208
rect 44288 2128 44608 2144
rect 51512 16896 51832 17456
rect 51512 16832 51520 16896
rect 51584 16832 51600 16896
rect 51664 16832 51680 16896
rect 51744 16832 51760 16896
rect 51824 16832 51832 16896
rect 51512 15808 51832 16832
rect 51512 15744 51520 15808
rect 51584 15744 51600 15808
rect 51664 15744 51680 15808
rect 51744 15744 51760 15808
rect 51824 15744 51832 15808
rect 51512 14720 51832 15744
rect 51512 14656 51520 14720
rect 51584 14656 51600 14720
rect 51664 14656 51680 14720
rect 51744 14656 51760 14720
rect 51824 14656 51832 14720
rect 51512 13632 51832 14656
rect 51512 13568 51520 13632
rect 51584 13568 51600 13632
rect 51664 13568 51680 13632
rect 51744 13568 51760 13632
rect 51824 13568 51832 13632
rect 51512 12544 51832 13568
rect 51512 12480 51520 12544
rect 51584 12480 51600 12544
rect 51664 12480 51680 12544
rect 51744 12480 51760 12544
rect 51824 12480 51832 12544
rect 51512 11456 51832 12480
rect 51512 11392 51520 11456
rect 51584 11392 51600 11456
rect 51664 11392 51680 11456
rect 51744 11392 51760 11456
rect 51824 11392 51832 11456
rect 51512 10368 51832 11392
rect 51512 10304 51520 10368
rect 51584 10304 51600 10368
rect 51664 10304 51680 10368
rect 51744 10304 51760 10368
rect 51824 10304 51832 10368
rect 51512 9280 51832 10304
rect 51512 9216 51520 9280
rect 51584 9216 51600 9280
rect 51664 9216 51680 9280
rect 51744 9216 51760 9280
rect 51824 9216 51832 9280
rect 51512 8192 51832 9216
rect 51512 8128 51520 8192
rect 51584 8128 51600 8192
rect 51664 8128 51680 8192
rect 51744 8128 51760 8192
rect 51824 8128 51832 8192
rect 51512 7104 51832 8128
rect 51512 7040 51520 7104
rect 51584 7040 51600 7104
rect 51664 7040 51680 7104
rect 51744 7040 51760 7104
rect 51824 7040 51832 7104
rect 51512 6016 51832 7040
rect 51512 5952 51520 6016
rect 51584 5952 51600 6016
rect 51664 5952 51680 6016
rect 51744 5952 51760 6016
rect 51824 5952 51832 6016
rect 51512 4928 51832 5952
rect 51512 4864 51520 4928
rect 51584 4864 51600 4928
rect 51664 4864 51680 4928
rect 51744 4864 51760 4928
rect 51824 4864 51832 4928
rect 51512 3840 51832 4864
rect 51512 3776 51520 3840
rect 51584 3776 51600 3840
rect 51664 3776 51680 3840
rect 51744 3776 51760 3840
rect 51824 3776 51832 3840
rect 51512 2752 51832 3776
rect 51512 2688 51520 2752
rect 51584 2688 51600 2752
rect 51664 2688 51680 2752
rect 51744 2688 51760 2752
rect 51824 2688 51832 2752
rect 51512 2128 51832 2688
rect 34467 1052 34533 1053
rect 34467 988 34468 1052
rect 34532 988 34533 1052
rect 34467 987 34533 988
use sky130_fd_sc_hd__diode_2  ANTENNA__0398__A dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 32568 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0400__B
timestamp 1649977179
transform -1 0 21252 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0401__A
timestamp 1649977179
transform 1 0 27784 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0402__A
timestamp 1649977179
transform 1 0 26956 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0404__A
timestamp 1649977179
transform -1 0 15180 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0404__B
timestamp 1649977179
transform -1 0 15732 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0407__A1
timestamp 1649977179
transform 1 0 33304 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0408__A2
timestamp 1649977179
transform -1 0 33304 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0408__C1
timestamp 1649977179
transform 1 0 33396 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0409__A1
timestamp 1649977179
transform -1 0 48208 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0409__B1
timestamp 1649977179
transform 1 0 41768 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0410__A1
timestamp 1649977179
transform -1 0 42044 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0412__A1
timestamp 1649977179
transform -1 0 42596 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0412__A2
timestamp 1649977179
transform -1 0 36156 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0413__A
timestamp 1649977179
transform 1 0 37812 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0414__A1
timestamp 1649977179
transform 1 0 34500 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0414__A2
timestamp 1649977179
transform 1 0 43240 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0414__B1
timestamp 1649977179
transform 1 0 42964 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0415__A1
timestamp 1649977179
transform 1 0 39836 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0416__A
timestamp 1649977179
transform 1 0 37260 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0416__C_N
timestamp 1649977179
transform 1 0 36432 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0417__A
timestamp 1649977179
transform 1 0 18584 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0417__B
timestamp 1649977179
transform -1 0 19412 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0418__A
timestamp 1649977179
transform 1 0 35236 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0419__A_N
timestamp 1649977179
transform 1 0 33764 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0419__B
timestamp 1649977179
transform 1 0 33672 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0420__A
timestamp 1649977179
transform 1 0 30636 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0421__B
timestamp 1649977179
transform -1 0 31648 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0422__A
timestamp 1649977179
transform 1 0 27232 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0422__B
timestamp 1649977179
transform 1 0 23736 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0427__A
timestamp 1649977179
transform 1 0 27968 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0428__B
timestamp 1649977179
transform -1 0 43148 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0430__A_N
timestamp 1649977179
transform 1 0 26312 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0431__A
timestamp 1649977179
transform 1 0 28704 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0432__A
timestamp 1649977179
transform -1 0 47288 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0433__B
timestamp 1649977179
transform 1 0 25392 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0435__A
timestamp 1649977179
transform -1 0 13340 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0436__A2
timestamp 1649977179
transform 1 0 22080 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0438__A
timestamp 1649977179
transform 1 0 28796 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0443__A
timestamp 1649977179
transform -1 0 9936 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0443__B
timestamp 1649977179
transform -1 0 10764 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0446__A
timestamp 1649977179
transform 1 0 24564 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0448__A
timestamp 1649977179
transform -1 0 45172 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0449__A
timestamp 1649977179
transform -1 0 23828 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0459__A
timestamp 1649977179
transform -1 0 54832 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0470__C
timestamp 1649977179
transform -1 0 49680 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0475__A
timestamp 1649977179
transform -1 0 58236 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0479__A2
timestamp 1649977179
transform 1 0 54096 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0482__A2
timestamp 1649977179
transform -1 0 53728 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0483__C
timestamp 1649977179
transform 1 0 55292 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0485__A
timestamp 1649977179
transform 1 0 22080 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0486__A
timestamp 1649977179
transform 1 0 10304 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0486__B
timestamp 1649977179
transform -1 0 11408 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0488__A
timestamp 1649977179
transform 1 0 3404 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0490__A
timestamp 1649977179
transform -1 0 3680 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0490__B
timestamp 1649977179
transform 1 0 2392 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0493__A
timestamp 1649977179
transform -1 0 3128 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0495__A
timestamp 1649977179
transform 1 0 18676 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0497__A
timestamp 1649977179
transform 1 0 14536 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0500__A
timestamp 1649977179
transform 1 0 22080 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0502__A
timestamp 1649977179
transform 1 0 36708 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0503__A
timestamp 1649977179
transform -1 0 34224 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0505__A
timestamp 1649977179
transform 1 0 37812 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0508__A
timestamp 1649977179
transform 1 0 32016 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0510__A
timestamp 1649977179
transform 1 0 23644 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0512__A
timestamp 1649977179
transform -1 0 19320 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0514__A
timestamp 1649977179
transform 1 0 25944 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0516__A
timestamp 1649977179
transform -1 0 38732 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0516__B
timestamp 1649977179
transform -1 0 38180 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0519__A
timestamp 1649977179
transform 1 0 21160 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0524__A
timestamp 1649977179
transform 1 0 42596 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0525__A
timestamp 1649977179
transform -1 0 51796 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0529__A
timestamp 1649977179
transform 1 0 23736 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0530__A
timestamp 1649977179
transform 1 0 2852 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0532__A
timestamp 1649977179
transform -1 0 3956 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0532__B
timestamp 1649977179
transform 1 0 4324 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0534__A
timestamp 1649977179
transform -1 0 3220 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0536__A
timestamp 1649977179
transform 1 0 13524 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0538__A
timestamp 1649977179
transform 1 0 22632 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0540__A
timestamp 1649977179
transform 1 0 38824 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0541__A
timestamp 1649977179
transform -1 0 40572 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0543__A
timestamp 1649977179
transform 1 0 29532 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0545__A
timestamp 1649977179
transform -1 0 16376 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0547__A
timestamp 1649977179
transform 1 0 39836 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0547__B
timestamp 1649977179
transform -1 0 39284 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0549__A
timestamp 1649977179
transform 1 0 17204 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0551__A
timestamp 1649977179
transform 1 0 50508 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0557__A
timestamp 1649977179
transform 1 0 20884 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0558__A
timestamp 1649977179
transform -1 0 4968 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0560__A
timestamp 1649977179
transform 1 0 5704 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0560__B
timestamp 1649977179
transform 1 0 5796 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0562__A
timestamp 1649977179
transform -1 0 4140 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0564__A
timestamp 1649977179
transform 1 0 10948 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0566__A
timestamp 1649977179
transform 1 0 20148 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0568__A
timestamp 1649977179
transform 1 0 36524 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0569__A
timestamp 1649977179
transform -1 0 39100 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0571__A
timestamp 1649977179
transform 1 0 34684 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0573__A
timestamp 1649977179
transform 1 0 18584 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0575__A
timestamp 1649977179
transform 1 0 37444 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0575__B
timestamp 1649977179
transform 1 0 38364 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0577__A
timestamp 1649977179
transform -1 0 18308 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0579__A
timestamp 1649977179
transform 1 0 46920 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0585__A
timestamp 1649977179
transform 1 0 20516 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0596__A
timestamp 1649977179
transform 1 0 37260 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0597__A
timestamp 1649977179
transform -1 0 37444 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0599__A
timestamp 1649977179
transform 1 0 34684 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0601__A
timestamp 1649977179
transform -1 0 17204 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0603__A
timestamp 1649977179
transform 1 0 36156 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0603__B
timestamp 1649977179
transform -1 0 40848 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0605__A
timestamp 1649977179
transform -1 0 13432 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0609__A
timestamp 1649977179
transform 1 0 43884 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0613__A
timestamp 1649977179
transform -1 0 1564 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0614__A
timestamp 1649977179
transform 1 0 6808 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0616__A
timestamp 1649977179
transform -1 0 10120 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0618__A
timestamp 1649977179
transform -1 0 7820 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0620__A
timestamp 1649977179
transform 1 0 13432 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0622__A
timestamp 1649977179
transform 1 0 28244 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0625__A
timestamp 1649977179
transform -1 0 23368 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0627__A
timestamp 1649977179
transform -1 0 45172 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0629__A
timestamp 1649977179
transform 1 0 45264 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0629__B
timestamp 1649977179
transform -1 0 46000 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0631__A
timestamp 1649977179
transform 1 0 24380 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0632__A
timestamp 1649977179
transform 1 0 11776 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0634__A
timestamp 1649977179
transform -1 0 12144 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0636__A
timestamp 1649977179
transform 1 0 12328 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0638__A
timestamp 1649977179
transform 1 0 10856 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0640__A
timestamp 1649977179
transform -1 0 30820 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0643__A
timestamp 1649977179
transform -1 0 21620 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0645__A
timestamp 1649977179
transform -1 0 47748 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0647__A
timestamp 1649977179
transform 1 0 26220 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0649__A
timestamp 1649977179
transform 1 0 41032 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0653__B
timestamp 1649977179
transform -1 0 6532 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0655__B
timestamp 1649977179
transform -1 0 22448 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0656__A
timestamp 1649977179
transform -1 0 40756 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0657__A
timestamp 1649977179
transform 1 0 27600 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0659__A
timestamp 1649977179
transform 1 0 42412 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0661__A
timestamp 1649977179
transform -1 0 31556 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0664__A
timestamp 1649977179
transform 1 0 24840 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0666__A
timestamp 1649977179
transform 1 0 39468 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0668__A
timestamp 1649977179
transform -1 0 45172 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0668__B
timestamp 1649977179
transform 1 0 44160 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0671__A_N
timestamp 1649977179
transform -1 0 15180 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0672__B
timestamp 1649977179
transform -1 0 1564 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0678__A
timestamp 1649977179
transform -1 0 2760 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0679__A
timestamp 1649977179
transform 1 0 9936 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0681__A1
timestamp 1649977179
transform -1 0 3956 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0681__C1
timestamp 1649977179
transform -1 0 3312 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0686__B
timestamp 1649977179
transform -1 0 3496 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0687__A
timestamp 1649977179
transform -1 0 30728 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0688__A
timestamp 1649977179
transform -1 0 44528 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0690__A
timestamp 1649977179
transform -1 0 27140 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0693__A1
timestamp 1649977179
transform 1 0 18124 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0693__C1
timestamp 1649977179
transform 1 0 19228 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0695__A1
timestamp 1649977179
transform 1 0 22172 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0695__C1
timestamp 1649977179
transform 1 0 21988 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0697__A1
timestamp 1649977179
transform -1 0 30176 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0697__C1
timestamp 1649977179
transform -1 0 23920 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0700__A
timestamp 1649977179
transform 1 0 14076 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0701__A1
timestamp 1649977179
transform -1 0 25208 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0701__C1
timestamp 1649977179
transform -1 0 24656 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0703__A1
timestamp 1649977179
transform 1 0 26036 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0703__C1
timestamp 1649977179
transform -1 0 32292 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0705__A
timestamp 1649977179
transform -1 0 40572 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0706__A
timestamp 1649977179
transform -1 0 40204 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0708__A1
timestamp 1649977179
transform -1 0 53176 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0708__C1
timestamp 1649977179
transform -1 0 53728 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0710__A1
timestamp 1649977179
transform 1 0 50968 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0710__C1
timestamp 1649977179
transform 1 0 50784 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0712__A1
timestamp 1649977179
transform -1 0 52256 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0712__C1
timestamp 1649977179
transform -1 0 42964 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0714__A
timestamp 1649977179
transform 1 0 17572 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0715__A1
timestamp 1649977179
transform -1 0 35788 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0715__C1
timestamp 1649977179
transform -1 0 46000 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0717__A1
timestamp 1649977179
transform -1 0 47748 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0717__C1
timestamp 1649977179
transform 1 0 37076 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0720__B
timestamp 1649977179
transform 1 0 15272 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0723__A
timestamp 1649977179
transform -1 0 19964 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0725__A1
timestamp 1649977179
transform 1 0 13524 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0725__C1
timestamp 1649977179
transform -1 0 14628 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0727__A1
timestamp 1649977179
transform -1 0 14260 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0727__C1
timestamp 1649977179
transform -1 0 15180 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0729__A1
timestamp 1649977179
transform -1 0 16192 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0729__C1
timestamp 1649977179
transform -1 0 17204 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0731__A
timestamp 1649977179
transform 1 0 23644 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0732__A1
timestamp 1649977179
transform -1 0 21988 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0732__C1
timestamp 1649977179
transform -1 0 22724 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0734__A1
timestamp 1649977179
transform -1 0 25760 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0734__C1
timestamp 1649977179
transform 1 0 25024 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0737__A
timestamp 1649977179
transform -1 0 29716 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0739__A1
timestamp 1649977179
transform -1 0 54832 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0739__C1
timestamp 1649977179
transform 1 0 56396 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0741__A1
timestamp 1649977179
transform -1 0 54096 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0741__C1
timestamp 1649977179
transform 1 0 43884 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0743__A1
timestamp 1649977179
transform -1 0 43516 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0743__C1
timestamp 1649977179
transform -1 0 57408 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0746__A1
timestamp 1649977179
transform -1 0 41952 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0746__C1
timestamp 1649977179
transform 1 0 35052 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0748__A1
timestamp 1649977179
transform -1 0 31556 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0748__C1
timestamp 1649977179
transform -1 0 39376 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0749__A
timestamp 1649977179
transform 1 0 46368 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0753__A
timestamp 1649977179
transform -1 0 4968 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0756__A
timestamp 1649977179
transform -1 0 19412 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0756__B
timestamp 1649977179
transform 1 0 19228 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0758__B
timestamp 1649977179
transform 1 0 4600 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0761__C1
timestamp 1649977179
transform -1 0 11040 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0762__A1
timestamp 1649977179
transform -1 0 18124 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0763__C1
timestamp 1649977179
transform -1 0 10488 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0766__C1
timestamp 1649977179
transform 1 0 18492 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0769__A1
timestamp 1649977179
transform -1 0 22724 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0771__A
timestamp 1649977179
transform -1 0 30452 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0773__A
timestamp 1649977179
transform 1 0 17480 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0774__A1
timestamp 1649977179
transform -1 0 25760 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0775__A
timestamp 1649977179
transform 1 0 19320 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0776__A1
timestamp 1649977179
transform -1 0 23920 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0785__A1
timestamp 1649977179
transform -1 0 11684 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0789__A1
timestamp 1649977179
transform -1 0 5336 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0793__C1
timestamp 1649977179
transform -1 0 11500 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0795__C1
timestamp 1649977179
transform 1 0 4048 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0798__A
timestamp 1649977179
transform -1 0 52348 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0799__CLK
timestamp 1649977179
transform 1 0 6440 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0800__CLK
timestamp 1649977179
transform 1 0 20792 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0801__CLK
timestamp 1649977179
transform 1 0 23092 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0802__CLK
timestamp 1649977179
transform 1 0 34684 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0803__CLK
timestamp 1649977179
transform -1 0 28796 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0804__CLK
timestamp 1649977179
transform 1 0 36616 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0805__CLK
timestamp 1649977179
transform 1 0 56948 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0806__CLK
timestamp 1649977179
transform 1 0 43332 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0807__CLK
timestamp 1649977179
transform -1 0 54464 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0808__CLK
timestamp 1649977179
transform 1 0 39836 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0809__CLK
timestamp 1649977179
transform 1 0 47564 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0810__CLK
timestamp 1649977179
transform 1 0 12972 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0811__CLK
timestamp 1649977179
transform -1 0 12788 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0812__CLK
timestamp 1649977179
transform -1 0 17020 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0813__CLK
timestamp 1649977179
transform 1 0 19964 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0814__CLK
timestamp 1649977179
transform 1 0 12420 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0815__CLK
timestamp 1649977179
transform -1 0 58052 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0816__CLK
timestamp 1649977179
transform 1 0 57776 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0817__CLK
timestamp 1649977179
transform -1 0 57408 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0818__CLK
timestamp 1649977179
transform -1 0 47104 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0819__CLK
timestamp 1649977179
transform 1 0 42412 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0820__CLK
timestamp 1649977179
transform -1 0 36800 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0820__SET_B
timestamp 1649977179
transform 1 0 33856 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0821__CLK
timestamp 1649977179
transform -1 0 38548 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0822__CLK
timestamp 1649977179
transform 1 0 41124 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0823__CLK
timestamp 1649977179
transform 1 0 35604 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0824__CLK
timestamp 1649977179
transform 1 0 5152 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0825__CLK
timestamp 1649977179
transform 1 0 8280 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0826__CLK
timestamp 1649977179
transform 1 0 9476 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0827__CLK
timestamp 1649977179
transform 1 0 21344 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0828__CLK
timestamp 1649977179
transform 1 0 23092 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0829__CLK
timestamp 1649977179
transform 1 0 39008 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0830__CLK
timestamp 1649977179
transform 1 0 16652 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0831__CLK
timestamp 1649977179
transform -1 0 26496 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0832__CLK
timestamp 1649977179
transform 1 0 6348 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0833__CLK
timestamp 1649977179
transform 1 0 5704 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0834__CLK
timestamp 1649977179
transform 1 0 12144 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0835__CLK
timestamp 1649977179
transform 1 0 9108 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0836__CLK
timestamp 1649977179
transform 1 0 6532 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0837__CLK
timestamp 1649977179
transform 1 0 5704 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0838__CLK
timestamp 1649977179
transform -1 0 1564 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0839__CLK
timestamp 1649977179
transform -1 0 6900 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0885__GATE_N
timestamp 1649977179
transform -1 0 3956 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0893__GATE_N
timestamp 1649977179
transform 1 0 8648 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0899__GATE_N
timestamp 1649977179
transform 1 0 11500 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0918__CLK
timestamp 1649977179
transform 1 0 44436 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0919__CLK
timestamp 1649977179
transform 1 0 48208 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0920__CLK
timestamp 1649977179
transform 1 0 52716 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0921__CLK
timestamp 1649977179
transform 1 0 48760 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0923__GATE_N
timestamp 1649977179
transform 1 0 53268 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0926__GATE_N
timestamp 1649977179
transform -1 0 58052 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0927__GATE_N
timestamp 1649977179
transform 1 0 54556 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0929__D
timestamp 1649977179
transform -1 0 20792 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0929__GATE_N
timestamp 1649977179
transform -1 0 20424 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1138__A
timestamp 1649977179
transform 1 0 12972 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1139__A
timestamp 1649977179
transform -1 0 2024 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1140__A
timestamp 1649977179
transform 1 0 17388 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1141__A
timestamp 1649977179
transform 1 0 14076 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_wb_clk_i_A
timestamp 1649977179
transform -1 0 26680 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input1_A
timestamp 1649977179
transform -1 0 2208 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input2_A
timestamp 1649977179
transform -1 0 2116 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input3_A
timestamp 1649977179
transform -1 0 3220 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input4_A
timestamp 1649977179
transform -1 0 16836 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input5_A
timestamp 1649977179
transform -1 0 5888 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input6_A
timestamp 1649977179
transform -1 0 2668 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input7_A
timestamp 1649977179
transform -1 0 18124 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input8_A
timestamp 1649977179
transform -1 0 4232 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input9_A
timestamp 1649977179
transform -1 0 9016 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input10_A
timestamp 1649977179
transform -1 0 9016 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input11_A
timestamp 1649977179
transform -1 0 2668 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input12_A
timestamp 1649977179
transform -1 0 10212 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input13_A
timestamp 1649977179
transform -1 0 11040 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input14_A
timestamp 1649977179
transform -1 0 6532 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input15_A
timestamp 1649977179
transform -1 0 7912 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input16_A
timestamp 1649977179
transform -1 0 2024 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input17_A
timestamp 1649977179
transform -1 0 10028 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input18_A
timestamp 1649977179
transform -1 0 3404 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input19_A
timestamp 1649977179
transform -1 0 9476 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input20_A
timestamp 1649977179
transform -1 0 6072 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input21_A
timestamp 1649977179
transform -1 0 9384 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input22_A
timestamp 1649977179
transform -1 0 5336 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input23_A
timestamp 1649977179
transform -1 0 10948 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input24_A
timestamp 1649977179
transform -1 0 12052 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input25_A
timestamp 1649977179
transform -1 0 8280 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input26_A
timestamp 1649977179
transform -1 0 7728 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input27_A
timestamp 1649977179
transform -1 0 6532 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output28_A
timestamp 1649977179
transform -1 0 13524 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output31_A
timestamp 1649977179
transform -1 0 15732 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output32_A
timestamp 1649977179
transform 1 0 21160 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output33_A
timestamp 1649977179
transform -1 0 17480 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output34_A
timestamp 1649977179
transform -1 0 26312 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output35_A
timestamp 1649977179
transform -1 0 17848 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output36_A
timestamp 1649977179
transform -1 0 21344 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output38_A
timestamp 1649977179
transform -1 0 23552 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output39_A
timestamp 1649977179
transform -1 0 18860 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output40_A
timestamp 1649977179
transform -1 0 24104 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output41_A
timestamp 1649977179
transform -1 0 24564 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output42_A
timestamp 1649977179
transform -1 0 14076 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output43_A
timestamp 1649977179
transform -1 0 18400 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output56_A
timestamp 1649977179
transform -1 0 7268 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output57_A
timestamp 1649977179
transform -1 0 8464 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output58_A
timestamp 1649977179
transform -1 0 7176 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_repeater72_A
timestamp 1649977179
transform -1 0 5888 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_repeater80_A
timestamp 1649977179
transform -1 0 35604 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 1380 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 1748 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13
timestamp 1649977179
transform 1 0 2300 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 3128 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32
timestamp 1649977179
transform 1 0 4048 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_52
timestamp 1649977179
transform 1 0 5888 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_57 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 6348 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_66
timestamp 1649977179
transform 1 0 7176 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_80
timestamp 1649977179
transform 1 0 8464 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_92
timestamp 1649977179
transform 1 0 9568 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_108
timestamp 1649977179
transform 1 0 11040 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_123 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 12420 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_131
timestamp 1649977179
transform 1 0 13156 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_136
timestamp 1649977179
transform 1 0 13616 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_141
timestamp 1649977179
transform 1 0 14076 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_148
timestamp 1649977179
transform 1 0 14720 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_156
timestamp 1649977179
transform 1 0 15456 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_164
timestamp 1649977179
transform 1 0 16192 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_169
timestamp 1649977179
transform 1 0 16652 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_176
timestamp 1649977179
transform 1 0 17296 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_184
timestamp 1649977179
transform 1 0 18032 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_192
timestamp 1649977179
transform 1 0 18768 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_197
timestamp 1649977179
transform 1 0 19228 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_212
timestamp 1649977179
transform 1 0 20608 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_220
timestamp 1649977179
transform 1 0 21344 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_230
timestamp 1649977179
transform 1 0 22264 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_239
timestamp 1649977179
transform 1 0 23092 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_247
timestamp 1649977179
transform 1 0 23828 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_251
timestamp 1649977179
transform 1 0 24196 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_257
timestamp 1649977179
transform 1 0 24748 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_265
timestamp 1649977179
transform 1 0 25484 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_269
timestamp 1649977179
transform 1 0 25852 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_276
timestamp 1649977179
transform 1 0 26496 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_283
timestamp 1649977179
transform 1 0 27140 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_290
timestamp 1649977179
transform 1 0 27784 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_297
timestamp 1649977179
transform 1 0 28428 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_304
timestamp 1649977179
transform 1 0 29072 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_309
timestamp 1649977179
transform 1 0 29532 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_315
timestamp 1649977179
transform 1 0 30084 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_322
timestamp 1649977179
transform 1 0 30728 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_332
timestamp 1649977179
transform 1 0 31648 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_339
timestamp 1649977179
transform 1 0 32292 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_353
timestamp 1649977179
transform 1 0 33580 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_360
timestamp 1649977179
transform 1 0 34224 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_368
timestamp 1649977179
transform 1 0 34960 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_375
timestamp 1649977179
transform 1 0 35604 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_382
timestamp 1649977179
transform 1 0 36248 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_388
timestamp 1649977179
transform 1 0 36800 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_396
timestamp 1649977179
transform 1 0 37536 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_403
timestamp 1649977179
transform 1 0 38180 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_410
timestamp 1649977179
transform 1 0 38824 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_416
timestamp 1649977179
transform 1 0 39376 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_424
timestamp 1649977179
transform 1 0 40112 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_431
timestamp 1649977179
transform 1 0 40756 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_438
timestamp 1649977179
transform 1 0 41400 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_444
timestamp 1649977179
transform 1 0 41952 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_452
timestamp 1649977179
transform 1 0 42688 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_459
timestamp 1649977179
transform 1 0 43332 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_466
timestamp 1649977179
transform 1 0 43976 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_472
timestamp 1649977179
transform 1 0 44528 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_480
timestamp 1649977179
transform 1 0 45264 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_487
timestamp 1649977179
transform 1 0 45908 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_494
timestamp 1649977179
transform 1 0 46552 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_500
timestamp 1649977179
transform 1 0 47104 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_508
timestamp 1649977179
transform 1 0 47840 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_515
timestamp 1649977179
transform 1 0 48484 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_522
timestamp 1649977179
transform 1 0 49128 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_528
timestamp 1649977179
transform 1 0 49680 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_536
timestamp 1649977179
transform 1 0 50416 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_543
timestamp 1649977179
transform 1 0 51060 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_550
timestamp 1649977179
transform 1 0 51704 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_556
timestamp 1649977179
transform 1 0 52256 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_564
timestamp 1649977179
transform 1 0 52992 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_571
timestamp 1649977179
transform 1 0 53636 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_578
timestamp 1649977179
transform 1 0 54280 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_584
timestamp 1649977179
transform 1 0 54832 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_592
timestamp 1649977179
transform 1 0 55568 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_599
timestamp 1649977179
transform 1 0 56212 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_606
timestamp 1649977179
transform 1 0 56856 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_612
timestamp 1649977179
transform 1 0 57408 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_619
timestamp 1649977179
transform 1 0 58052 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_5
timestamp 1649977179
transform 1 0 1564 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_13
timestamp 1649977179
transform 1 0 2300 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_24
timestamp 1649977179
transform 1 0 3312 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_35
timestamp 1649977179
transform 1 0 4324 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_39
timestamp 1649977179
transform 1 0 4692 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_44
timestamp 1649977179
transform 1 0 5152 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_52
timestamp 1649977179
transform 1 0 5888 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_59
timestamp 1649977179
transform 1 0 6532 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_73
timestamp 1649977179
transform 1 0 7820 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_87
timestamp 1649977179
transform 1 0 9108 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_101
timestamp 1649977179
transform 1 0 10396 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_108
timestamp 1649977179
transform 1 0 11040 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_119
timestamp 1649977179
transform 1 0 12052 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_125
timestamp 1649977179
transform 1 0 12604 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_133
timestamp 1649977179
transform 1 0 13340 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_141
timestamp 1649977179
transform 1 0 14076 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_149
timestamp 1649977179
transform 1 0 14812 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_163
timestamp 1649977179
transform 1 0 16100 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_167
timestamp 1649977179
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_169 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 16652 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_177
timestamp 1649977179
transform 1 0 17388 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_181
timestamp 1649977179
transform 1 0 17756 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_1_186
timestamp 1649977179
transform 1 0 18216 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_196
timestamp 1649977179
transform 1 0 19136 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_220
timestamp 1649977179
transform 1 0 21344 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_230
timestamp 1649977179
transform 1 0 22264 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_234
timestamp 1649977179
transform 1 0 22632 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_239
timestamp 1649977179
transform 1 0 23092 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_247
timestamp 1649977179
transform 1 0 23828 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_1_258
timestamp 1649977179
transform 1 0 24840 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_270
timestamp 1649977179
transform 1 0 25944 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_276
timestamp 1649977179
transform 1 0 26496 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_284
timestamp 1649977179
transform 1 0 27232 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_288
timestamp 1649977179
transform 1 0 27600 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_292
timestamp 1649977179
transform 1 0 27968 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_299
timestamp 1649977179
transform 1 0 28612 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_313
timestamp 1649977179
transform 1 0 29900 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_319
timestamp 1649977179
transform 1 0 30452 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_331
timestamp 1649977179
transform 1 0 31556 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_335
timestamp 1649977179
transform 1 0 31924 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_337
timestamp 1649977179
transform 1 0 32108 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_361
timestamp 1649977179
transform 1 0 34316 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_375
timestamp 1649977179
transform 1 0 35604 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_382
timestamp 1649977179
transform 1 0 36248 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_388
timestamp 1649977179
transform 1 0 36800 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_399
timestamp 1649977179
transform 1 0 37812 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_406
timestamp 1649977179
transform 1 0 38456 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_413
timestamp 1649977179
transform 1 0 39100 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_420
timestamp 1649977179
transform 1 0 39744 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_427
timestamp 1649977179
transform 1 0 40388 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_437
timestamp 1649977179
transform 1 0 41308 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_444
timestamp 1649977179
transform 1 0 41952 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_452
timestamp 1649977179
transform 1 0 42688 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_456
timestamp 1649977179
transform 1 0 43056 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_465
timestamp 1649977179
transform 1 0 43884 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_472
timestamp 1649977179
transform 1 0 44528 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_479
timestamp 1649977179
transform 1 0 45172 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_486
timestamp 1649977179
transform 1 0 45816 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_493
timestamp 1649977179
transform 1 0 46460 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_500
timestamp 1649977179
transform 1 0 47104 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_507
timestamp 1649977179
transform 1 0 47748 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_527
timestamp 1649977179
transform 1 0 49588 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_534
timestamp 1649977179
transform 1 0 50232 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_541
timestamp 1649977179
transform 1 0 50876 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_548
timestamp 1649977179
transform 1 0 51520 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_555
timestamp 1649977179
transform 1 0 52164 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_559
timestamp 1649977179
transform 1 0 52532 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_565
timestamp 1649977179
transform 1 0 53084 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_572
timestamp 1649977179
transform 1 0 53728 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_579
timestamp 1649977179
transform 1 0 54372 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_586
timestamp 1649977179
transform 1 0 55016 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_593
timestamp 1649977179
transform 1 0 55660 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_600
timestamp 1649977179
transform 1 0 56304 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_607
timestamp 1649977179
transform 1 0 56948 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_615
timestamp 1649977179
transform 1 0 57684 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_1_619
timestamp 1649977179
transform 1 0 58052 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_2_3
timestamp 1649977179
transform 1 0 1380 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_11
timestamp 1649977179
transform 1 0 2116 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_21
timestamp 1649977179
transform 1 0 3036 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp 1649977179
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_37
timestamp 1649977179
transform 1 0 4508 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_2_61
timestamp 1649977179
transform 1 0 6716 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_67
timestamp 1649977179
transform 1 0 7268 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_75
timestamp 1649977179
transform 1 0 8004 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_83
timestamp 1649977179
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_85
timestamp 1649977179
transform 1 0 8924 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_96
timestamp 1649977179
transform 1 0 9936 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_108
timestamp 1649977179
transform 1 0 11040 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_112
timestamp 1649977179
transform 1 0 11408 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_129
timestamp 1649977179
transform 1 0 12972 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_136
timestamp 1649977179
transform 1 0 13616 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_141
timestamp 1649977179
transform 1 0 14076 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_150
timestamp 1649977179
transform 1 0 14904 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_156
timestamp 1649977179
transform 1 0 15456 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_166
timestamp 1649977179
transform 1 0 16376 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_177
timestamp 1649977179
transform 1 0 17388 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_184
timestamp 1649977179
transform 1 0 18032 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_192
timestamp 1649977179
transform 1 0 18768 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_207
timestamp 1649977179
transform 1 0 20148 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_213
timestamp 1649977179
transform 1 0 20700 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_234
timestamp 1649977179
transform 1 0 22632 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_242
timestamp 1649977179
transform 1 0 23368 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_248
timestamp 1649977179
transform 1 0 23920 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_253
timestamp 1649977179
transform 1 0 24380 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_260
timestamp 1649977179
transform 1 0 25024 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_280
timestamp 1649977179
transform 1 0 26864 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_287
timestamp 1649977179
transform 1 0 27508 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_291
timestamp 1649977179
transform 1 0 27876 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_296
timestamp 1649977179
transform 1 0 28336 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_304
timestamp 1649977179
transform 1 0 29072 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_319
timestamp 1649977179
transform 1 0 30452 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_2_347
timestamp 1649977179
transform 1 0 33028 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_353
timestamp 1649977179
transform 1 0 33580 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_360
timestamp 1649977179
transform 1 0 34224 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_368
timestamp 1649977179
transform 1 0 34960 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_2_390
timestamp 1649977179
transform 1 0 36984 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_394
timestamp 1649977179
transform 1 0 37352 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_412
timestamp 1649977179
transform 1 0 39008 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_421
timestamp 1649977179
transform 1 0 39836 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_429
timestamp 1649977179
transform 1 0 40572 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_439
timestamp 1649977179
transform 1 0 41492 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_446
timestamp 1649977179
transform 1 0 42136 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_450
timestamp 1649977179
transform 1 0 42504 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_459
timestamp 1649977179
transform 1 0 43332 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_471
timestamp 1649977179
transform 1 0 44436 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_475
timestamp 1649977179
transform 1 0 44804 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_477
timestamp 1649977179
transform 1 0 44988 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_495
timestamp 1649977179
transform 1 0 46644 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_502
timestamp 1649977179
transform 1 0 47288 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_2_526
timestamp 1649977179
transform 1 0 49496 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_2_536
timestamp 1649977179
transform 1 0 50416 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_543
timestamp 1649977179
transform 1 0 51060 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_550
timestamp 1649977179
transform 1 0 51704 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_2_568
timestamp 1649977179
transform 1 0 53360 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_575
timestamp 1649977179
transform 1 0 54004 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_583
timestamp 1649977179
transform 1 0 54740 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_587
timestamp 1649977179
transform 1 0 55108 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_592
timestamp 1649977179
transform 1 0 55568 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_599
timestamp 1649977179
transform 1 0 56212 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_606
timestamp 1649977179
transform 1 0 56856 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_612
timestamp 1649977179
transform 1 0 57408 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_618
timestamp 1649977179
transform 1 0 57960 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_624
timestamp 1649977179
transform 1 0 58512 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_3
timestamp 1649977179
transform 1 0 1380 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_7
timestamp 1649977179
transform 1 0 1748 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_11
timestamp 1649977179
transform 1 0 2116 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_23
timestamp 1649977179
transform 1 0 3220 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_31
timestamp 1649977179
transform 1 0 3956 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_36
timestamp 1649977179
transform 1 0 4416 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_44
timestamp 1649977179
transform 1 0 5152 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_52
timestamp 1649977179
transform 1 0 5888 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_57
timestamp 1649977179
transform 1 0 6348 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_62
timestamp 1649977179
transform 1 0 6808 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_71
timestamp 1649977179
transform 1 0 7636 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_91
timestamp 1649977179
transform 1 0 9476 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_97
timestamp 1649977179
transform 1 0 10028 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_3_106
timestamp 1649977179
transform 1 0 10856 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_3_129
timestamp 1649977179
transform 1 0 12972 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_3_145
timestamp 1649977179
transform 1 0 14444 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_153
timestamp 1649977179
transform 1 0 15180 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_157
timestamp 1649977179
transform 1 0 15548 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_164
timestamp 1649977179
transform 1 0 16192 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_177
timestamp 1649977179
transform 1 0 17388 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_183
timestamp 1649977179
transform 1 0 17940 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_188
timestamp 1649977179
transform 1 0 18400 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_200
timestamp 1649977179
transform 1 0 19504 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_220
timestamp 1649977179
transform 1 0 21344 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_233
timestamp 1649977179
transform 1 0 22540 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_3_242
timestamp 1649977179
transform 1 0 23368 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_250
timestamp 1649977179
transform 1 0 24104 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_3_264
timestamp 1649977179
transform 1 0 25392 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_274
timestamp 1649977179
transform 1 0 26312 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_3_281
timestamp 1649977179
transform 1 0 26956 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_299
timestamp 1649977179
transform 1 0 28612 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_307
timestamp 1649977179
transform 1 0 29348 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_311
timestamp 1649977179
transform 1 0 29716 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_318
timestamp 1649977179
transform 1 0 30360 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_332
timestamp 1649977179
transform 1 0 31648 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_353
timestamp 1649977179
transform 1 0 33580 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_367
timestamp 1649977179
transform 1 0 34868 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_379
timestamp 1649977179
transform 1 0 35972 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_386
timestamp 1649977179
transform 1 0 36616 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_3_401
timestamp 1649977179
transform 1 0 37996 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_405
timestamp 1649977179
transform 1 0 38364 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_416
timestamp 1649977179
transform 1 0 39376 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_430
timestamp 1649977179
transform 1 0 40664 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_440
timestamp 1649977179
transform 1 0 41584 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_3_451
timestamp 1649977179
transform 1 0 42596 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_463
timestamp 1649977179
transform 1 0 43700 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_475
timestamp 1649977179
transform 1 0 44804 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_482
timestamp 1649977179
transform 1 0 45448 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_489
timestamp 1649977179
transform 1 0 46092 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_496
timestamp 1649977179
transform 1 0 46736 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_3_508
timestamp 1649977179
transform 1 0 47840 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_512
timestamp 1649977179
transform 1 0 48208 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_529
timestamp 1649977179
transform 1 0 49772 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_536
timestamp 1649977179
transform 1 0 50416 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_543
timestamp 1649977179
transform 1 0 51060 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_549
timestamp 1649977179
transform 1 0 51612 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_556
timestamp 1649977179
transform 1 0 52256 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_564
timestamp 1649977179
transform 1 0 52992 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_571
timestamp 1649977179
transform 1 0 53636 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_581
timestamp 1649977179
transform 1 0 54556 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_590
timestamp 1649977179
transform 1 0 55384 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_597
timestamp 1649977179
transform 1 0 56028 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_603
timestamp 1649977179
transform 1 0 56580 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_609
timestamp 1649977179
transform 1 0 57132 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_615
timestamp 1649977179
transform 1 0 57684 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_620
timestamp 1649977179
transform 1 0 58144 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_624
timestamp 1649977179
transform 1 0 58512 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_4_3
timestamp 1649977179
transform 1 0 1380 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_11
timestamp 1649977179
transform 1 0 2116 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_23
timestamp 1649977179
transform 1 0 3220 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 1649977179
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_29
timestamp 1649977179
transform 1 0 3772 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_37
timestamp 1649977179
transform 1 0 4508 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_58
timestamp 1649977179
transform 1 0 6440 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_4_78
timestamp 1649977179
transform 1 0 8280 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_4_90
timestamp 1649977179
transform 1 0 9384 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_99
timestamp 1649977179
transform 1 0 10212 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_111
timestamp 1649977179
transform 1 0 11316 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_131
timestamp 1649977179
transform 1 0 13156 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_139
timestamp 1649977179
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_143
timestamp 1649977179
transform 1 0 14260 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_151
timestamp 1649977179
transform 1 0 14996 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_171
timestamp 1649977179
transform 1 0 16836 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_4_183
timestamp 1649977179
transform 1 0 17940 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_191
timestamp 1649977179
transform 1 0 18676 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_195
timestamp 1649977179
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_4_197
timestamp 1649977179
transform 1 0 19228 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_216
timestamp 1649977179
transform 1 0 20976 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_4_226
timestamp 1649977179
transform 1 0 21896 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_232
timestamp 1649977179
transform 1 0 22448 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_241
timestamp 1649977179
transform 1 0 23276 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_248
timestamp 1649977179
transform 1 0 23920 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_257
timestamp 1649977179
transform 1 0 24748 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_267
timestamp 1649977179
transform 1 0 25668 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_273
timestamp 1649977179
transform 1 0 26220 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_297
timestamp 1649977179
transform 1 0 28428 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_304
timestamp 1649977179
transform 1 0 29072 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_317
timestamp 1649977179
transform 1 0 30268 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_323
timestamp 1649977179
transform 1 0 30820 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_335
timestamp 1649977179
transform 1 0 31924 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_343
timestamp 1649977179
transform 1 0 32660 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_360
timestamp 1649977179
transform 1 0 34224 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_367
timestamp 1649977179
transform 1 0 34868 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_374
timestamp 1649977179
transform 1 0 35512 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_378
timestamp 1649977179
transform 1 0 35880 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_4_387
timestamp 1649977179
transform 1 0 36708 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_4_409
timestamp 1649977179
transform 1 0 38732 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_416
timestamp 1649977179
transform 1 0 39376 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_428
timestamp 1649977179
transform 1 0 40480 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_438
timestamp 1649977179
transform 1 0 41400 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_445
timestamp 1649977179
transform 1 0 42044 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_4_461
timestamp 1649977179
transform 1 0 43516 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_465
timestamp 1649977179
transform 1 0 43884 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_472
timestamp 1649977179
transform 1 0 44528 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_483
timestamp 1649977179
transform 1 0 45540 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_493
timestamp 1649977179
transform 1 0 46460 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_501
timestamp 1649977179
transform 1 0 47196 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_518
timestamp 1649977179
transform 1 0 48760 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_4_525
timestamp 1649977179
transform 1 0 49404 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_531
timestamp 1649977179
transform 1 0 49956 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_536
timestamp 1649977179
transform 1 0 50416 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_4_543
timestamp 1649977179
transform 1 0 51060 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_549
timestamp 1649977179
transform 1 0 51612 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_562
timestamp 1649977179
transform 1 0 52808 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_570
timestamp 1649977179
transform 1 0 53544 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_576
timestamp 1649977179
transform 1 0 54096 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_580
timestamp 1649977179
transform 1 0 54464 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_584
timestamp 1649977179
transform 1 0 54832 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_594
timestamp 1649977179
transform 1 0 55752 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_598
timestamp 1649977179
transform 1 0 56120 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_611
timestamp 1649977179
transform 1 0 57316 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_4_618
timestamp 1649977179
transform 1 0 57960 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_624
timestamp 1649977179
transform 1 0 58512 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_5
timestamp 1649977179
transform 1 0 1564 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_14
timestamp 1649977179
transform 1 0 2392 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_23
timestamp 1649977179
transform 1 0 3220 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_27
timestamp 1649977179
transform 1 0 3588 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_32
timestamp 1649977179
transform 1 0 4048 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_52
timestamp 1649977179
transform 1 0 5888 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_59
timestamp 1649977179
transform 1 0 6532 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_67
timestamp 1649977179
transform 1 0 7268 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_87
timestamp 1649977179
transform 1 0 9108 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_96
timestamp 1649977179
transform 1 0 9936 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_108
timestamp 1649977179
transform 1 0 11040 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_123
timestamp 1649977179
transform 1 0 12420 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_137
timestamp 1649977179
transform 1 0 13708 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_151
timestamp 1649977179
transform 1 0 14996 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_5_164
timestamp 1649977179
transform 1 0 16192 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_185
timestamp 1649977179
transform 1 0 18124 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_194
timestamp 1649977179
transform 1 0 18952 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_200
timestamp 1649977179
transform 1 0 19504 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_220
timestamp 1649977179
transform 1 0 21344 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_229
timestamp 1649977179
transform 1 0 22172 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_233
timestamp 1649977179
transform 1 0 22540 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_237
timestamp 1649977179
transform 1 0 22908 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_257
timestamp 1649977179
transform 1 0 24748 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_5_271
timestamp 1649977179
transform 1 0 26036 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_279
timestamp 1649977179
transform 1 0 26772 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_283
timestamp 1649977179
transform 1 0 27140 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_293
timestamp 1649977179
transform 1 0 28060 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_303
timestamp 1649977179
transform 1 0 28980 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_307
timestamp 1649977179
transform 1 0 29348 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_311
timestamp 1649977179
transform 1 0 29716 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_315
timestamp 1649977179
transform 1 0 30084 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_332
timestamp 1649977179
transform 1 0 31648 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_343
timestamp 1649977179
transform 1 0 32660 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_351
timestamp 1649977179
transform 1 0 33396 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_376
timestamp 1649977179
transform 1 0 35696 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_384
timestamp 1649977179
transform 1 0 36432 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_388
timestamp 1649977179
transform 1 0 36800 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_393
timestamp 1649977179
transform 1 0 37260 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_5_398
timestamp 1649977179
transform 1 0 37720 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_406
timestamp 1649977179
transform 1 0 38456 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_413
timestamp 1649977179
transform 1 0 39100 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_417
timestamp 1649977179
transform 1 0 39468 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_434
timestamp 1649977179
transform 1 0 41032 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_5_441
timestamp 1649977179
transform 1 0 41676 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_447
timestamp 1649977179
transform 1 0 42228 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_452
timestamp 1649977179
transform 1 0 42688 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_460
timestamp 1649977179
transform 1 0 43424 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_477
timestamp 1649977179
transform 1 0 44988 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_487
timestamp 1649977179
transform 1 0 45908 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_495
timestamp 1649977179
transform 1 0 46644 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_500
timestamp 1649977179
transform 1 0 47104 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_507
timestamp 1649977179
transform 1 0 47748 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_531
timestamp 1649977179
transform 1 0 49956 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_538
timestamp 1649977179
transform 1 0 50600 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_544
timestamp 1649977179
transform 1 0 51152 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_5_555
timestamp 1649977179
transform 1 0 52164 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_559
timestamp 1649977179
transform 1 0 52532 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_569
timestamp 1649977179
transform 1 0 53452 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_580
timestamp 1649977179
transform 1 0 54464 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_5_590
timestamp 1649977179
transform 1 0 55384 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_5_601
timestamp 1649977179
transform 1 0 56396 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_608
timestamp 1649977179
transform 1 0 57040 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_5_620
timestamp 1649977179
transform 1 0 58144 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_624
timestamp 1649977179
transform 1 0 58512 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_3
timestamp 1649977179
transform 1 0 1380 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_8
timestamp 1649977179
transform 1 0 1840 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_15
timestamp 1649977179
transform 1 0 2484 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_24
timestamp 1649977179
transform 1 0 3312 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_6_37
timestamp 1649977179
transform 1 0 4508 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_6_61
timestamp 1649977179
transform 1 0 6716 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_67
timestamp 1649977179
transform 1 0 7268 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_72
timestamp 1649977179
transform 1 0 7728 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_80
timestamp 1649977179
transform 1 0 8464 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_89
timestamp 1649977179
transform 1 0 9292 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_6_98
timestamp 1649977179
transform 1 0 10120 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_6_120
timestamp 1649977179
transform 1 0 12144 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_128
timestamp 1649977179
transform 1 0 12880 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_136
timestamp 1649977179
transform 1 0 13616 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_6_157
timestamp 1649977179
transform 1 0 15548 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_165
timestamp 1649977179
transform 1 0 16284 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_174
timestamp 1649977179
transform 1 0 17112 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_180
timestamp 1649977179
transform 1 0 17664 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_192
timestamp 1649977179
transform 1 0 18768 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_6_202
timestamp 1649977179
transform 1 0 19688 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_6_213
timestamp 1649977179
transform 1 0 20700 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_220
timestamp 1649977179
transform 1 0 21344 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_240
timestamp 1649977179
transform 1 0 23184 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_244
timestamp 1649977179
transform 1 0 23552 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_248
timestamp 1649977179
transform 1 0 23920 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_6_253
timestamp 1649977179
transform 1 0 24380 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_6_272
timestamp 1649977179
transform 1 0 26128 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_278
timestamp 1649977179
transform 1 0 26680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_284
timestamp 1649977179
transform 1 0 27232 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_304
timestamp 1649977179
transform 1 0 29072 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_314
timestamp 1649977179
transform 1 0 29992 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_6_321
timestamp 1649977179
transform 1 0 30636 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_327
timestamp 1649977179
transform 1 0 31188 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_344
timestamp 1649977179
transform 1 0 32752 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_350
timestamp 1649977179
transform 1 0 33304 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_6_356
timestamp 1649977179
transform 1 0 33856 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_6_369
timestamp 1649977179
transform 1 0 35052 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_376
timestamp 1649977179
transform 1 0 35696 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_401
timestamp 1649977179
transform 1 0 37996 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_408
timestamp 1649977179
transform 1 0 38640 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_6_414
timestamp 1649977179
transform 1 0 39192 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_6_423
timestamp 1649977179
transform 1 0 40020 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_430
timestamp 1649977179
transform 1 0 40664 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_454
timestamp 1649977179
transform 1 0 42872 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_6_460
timestamp 1649977179
transform 1 0 43424 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_6_469
timestamp 1649977179
transform 1 0 44252 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_475
timestamp 1649977179
transform 1 0 44804 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_480
timestamp 1649977179
transform 1 0 45264 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_487
timestamp 1649977179
transform 1 0 45908 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_6_494
timestamp 1649977179
transform 1 0 46552 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_500
timestamp 1649977179
transform 1 0 47104 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_504
timestamp 1649977179
transform 1 0 47472 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_528
timestamp 1649977179
transform 1 0 49680 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_536
timestamp 1649977179
transform 1 0 50416 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_6_542
timestamp 1649977179
transform 1 0 50968 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_6_560
timestamp 1649977179
transform 1 0 52624 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_566
timestamp 1649977179
transform 1 0 53176 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_572
timestamp 1649977179
transform 1 0 53728 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_6_579
timestamp 1649977179
transform 1 0 54372 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_587
timestamp 1649977179
transform 1 0 55108 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_599
timestamp 1649977179
transform 1 0 56212 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_615
timestamp 1649977179
transform 1 0 57684 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_621
timestamp 1649977179
transform 1 0 58236 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_3
timestamp 1649977179
transform 1 0 1380 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_7
timestamp 1649977179
transform 1 0 1748 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_11
timestamp 1649977179
transform 1 0 2116 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_18
timestamp 1649977179
transform 1 0 2760 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_34
timestamp 1649977179
transform 1 0 4232 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_46
timestamp 1649977179
transform 1 0 5336 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_52
timestamp 1649977179
transform 1 0 5888 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_7_57
timestamp 1649977179
transform 1 0 6348 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_7_63
timestamp 1649977179
transform 1 0 6900 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_79
timestamp 1649977179
transform 1 0 8372 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_83
timestamp 1649977179
transform 1 0 8740 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_96
timestamp 1649977179
transform 1 0 9936 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_108
timestamp 1649977179
transform 1 0 11040 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_7_117
timestamp 1649977179
transform 1 0 11868 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_125
timestamp 1649977179
transform 1 0 12604 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_130
timestamp 1649977179
transform 1 0 13064 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_142
timestamp 1649977179
transform 1 0 14168 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_7_151
timestamp 1649977179
transform 1 0 14996 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_159
timestamp 1649977179
transform 1 0 15732 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_164
timestamp 1649977179
transform 1 0 16192 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_171
timestamp 1649977179
transform 1 0 16836 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_183
timestamp 1649977179
transform 1 0 17940 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_187
timestamp 1649977179
transform 1 0 18308 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_193
timestamp 1649977179
transform 1 0 18860 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_7_204
timestamp 1649977179
transform 1 0 19872 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_220
timestamp 1649977179
transform 1 0 21344 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_7_233
timestamp 1649977179
transform 1 0 22540 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_241
timestamp 1649977179
transform 1 0 23276 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_245
timestamp 1649977179
transform 1 0 23644 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_254
timestamp 1649977179
transform 1 0 24472 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_266
timestamp 1649977179
transform 1 0 25576 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_7_273
timestamp 1649977179
transform 1 0 26220 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_279
timestamp 1649977179
transform 1 0 26772 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_7_281
timestamp 1649977179
transform 1 0 26956 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_7_287
timestamp 1649977179
transform 1 0 27508 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_7_299
timestamp 1649977179
transform 1 0 28612 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_305
timestamp 1649977179
transform 1 0 29164 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_314
timestamp 1649977179
transform 1 0 29992 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_323
timestamp 1649977179
transform 1 0 30820 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_7_330
timestamp 1649977179
transform 1 0 31464 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_7_343
timestamp 1649977179
transform 1 0 32660 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_351
timestamp 1649977179
transform 1 0 33396 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_357
timestamp 1649977179
transform 1 0 33948 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_367
timestamp 1649977179
transform 1 0 34868 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_7_375
timestamp 1649977179
transform 1 0 35604 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_7_386
timestamp 1649977179
transform 1 0 36616 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_7_393
timestamp 1649977179
transform 1 0 37260 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_399
timestamp 1649977179
transform 1 0 37812 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_424
timestamp 1649977179
transform 1 0 40112 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_428
timestamp 1649977179
transform 1 0 40480 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_432
timestamp 1649977179
transform 1 0 40848 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_436
timestamp 1649977179
transform 1 0 41216 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_443
timestamp 1649977179
transform 1 0 41860 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_447
timestamp 1649977179
transform 1 0 42228 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_451
timestamp 1649977179
transform 1 0 42596 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_7_457
timestamp 1649977179
transform 1 0 43148 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_7_482
timestamp 1649977179
transform 1 0 45448 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_7_488
timestamp 1649977179
transform 1 0 46000 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_496
timestamp 1649977179
transform 1 0 46736 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_500
timestamp 1649977179
transform 1 0 47104 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_505
timestamp 1649977179
transform 1 0 47564 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_526
timestamp 1649977179
transform 1 0 49496 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_533
timestamp 1649977179
transform 1 0 50140 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_540
timestamp 1649977179
transform 1 0 50784 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_556
timestamp 1649977179
transform 1 0 52256 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_561
timestamp 1649977179
transform 1 0 52716 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_577
timestamp 1649977179
transform 1 0 54188 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_591
timestamp 1649977179
transform 1 0 55476 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_601
timestamp 1649977179
transform 1 0 56396 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_7_608
timestamp 1649977179
transform 1 0 57040 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_7_620
timestamp 1649977179
transform 1 0 58144 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_624
timestamp 1649977179
transform 1 0 58512 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_3
timestamp 1649977179
transform 1 0 1380 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_10
timestamp 1649977179
transform 1 0 2024 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_17
timestamp 1649977179
transform 1 0 2668 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_24
timestamp 1649977179
transform 1 0 3312 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_8_41
timestamp 1649977179
transform 1 0 4876 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_8_50
timestamp 1649977179
transform 1 0 5704 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_57
timestamp 1649977179
transform 1 0 6348 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_8_69
timestamp 1649977179
transform 1 0 7452 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_75
timestamp 1649977179
transform 1 0 8004 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_80
timestamp 1649977179
transform 1 0 8464 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_8_85
timestamp 1649977179
transform 1 0 8924 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_8_92
timestamp 1649977179
transform 1 0 9568 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_96
timestamp 1649977179
transform 1 0 9936 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_8_101
timestamp 1649977179
transform 1 0 10396 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_107
timestamp 1649977179
transform 1 0 10948 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_120
timestamp 1649977179
transform 1 0 12144 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_136
timestamp 1649977179
transform 1 0 13616 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_8_145
timestamp 1649977179
transform 1 0 14444 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_8_154
timestamp 1649977179
transform 1 0 15272 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_161
timestamp 1649977179
transform 1 0 15916 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_168
timestamp 1649977179
transform 1 0 16560 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_184
timestamp 1649977179
transform 1 0 18032 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_188
timestamp 1649977179
transform 1 0 18400 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_192
timestamp 1649977179
transform 1 0 18768 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_8_209
timestamp 1649977179
transform 1 0 20332 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_215
timestamp 1649977179
transform 1 0 20884 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_219
timestamp 1649977179
transform 1 0 21252 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_226
timestamp 1649977179
transform 1 0 21896 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_242
timestamp 1649977179
transform 1 0 23368 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_248
timestamp 1649977179
transform 1 0 23920 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_255
timestamp 1649977179
transform 1 0 24564 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_264
timestamp 1649977179
transform 1 0 25392 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_273
timestamp 1649977179
transform 1 0 26220 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_282
timestamp 1649977179
transform 1 0 27048 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_290
timestamp 1649977179
transform 1 0 27784 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_304
timestamp 1649977179
transform 1 0 29072 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_315
timestamp 1649977179
transform 1 0 30084 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_324
timestamp 1649977179
transform 1 0 30912 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_328
timestamp 1649977179
transform 1 0 31280 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_331
timestamp 1649977179
transform 1 0 31556 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_342
timestamp 1649977179
transform 1 0 32568 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_8_350
timestamp 1649977179
transform 1 0 33304 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_356
timestamp 1649977179
transform 1 0 33856 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_360
timestamp 1649977179
transform 1 0 34224 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_365
timestamp 1649977179
transform 1 0 34684 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_373
timestamp 1649977179
transform 1 0 35420 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_384
timestamp 1649977179
transform 1 0 36432 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_400
timestamp 1649977179
transform 1 0 37904 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_404
timestamp 1649977179
transform 1 0 38272 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_408
timestamp 1649977179
transform 1 0 38640 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_416
timestamp 1649977179
transform 1 0 39376 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_421
timestamp 1649977179
transform 1 0 39836 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_8_429
timestamp 1649977179
transform 1 0 40572 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_8_441
timestamp 1649977179
transform 1 0 41676 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_447
timestamp 1649977179
transform 1 0 42228 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_452
timestamp 1649977179
transform 1 0 42688 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_8_472
timestamp 1649977179
transform 1 0 44528 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_489
timestamp 1649977179
transform 1 0 46092 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_493
timestamp 1649977179
transform 1 0 46460 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_506
timestamp 1649977179
transform 1 0 47656 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_512
timestamp 1649977179
transform 1 0 48208 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_528
timestamp 1649977179
transform 1 0 49680 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_533
timestamp 1649977179
transform 1 0 50140 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_546
timestamp 1649977179
transform 1 0 51336 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_8_554
timestamp 1649977179
transform 1 0 52072 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_8_574
timestamp 1649977179
transform 1 0 53912 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_8_580
timestamp 1649977179
transform 1 0 54464 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_8_589
timestamp 1649977179
transform 1 0 55292 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_8_598
timestamp 1649977179
transform 1 0 56120 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_604
timestamp 1649977179
transform 1 0 56672 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_617
timestamp 1649977179
transform 1 0 57868 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_3
timestamp 1649977179
transform 1 0 1380 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_8
timestamp 1649977179
transform 1 0 1840 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_17
timestamp 1649977179
transform 1 0 2668 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_9_26
timestamp 1649977179
transform 1 0 3496 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_32
timestamp 1649977179
transform 1 0 4048 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_45
timestamp 1649977179
transform 1 0 5244 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_52
timestamp 1649977179
transform 1 0 5888 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_62
timestamp 1649977179
transform 1 0 6808 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_71
timestamp 1649977179
transform 1 0 7636 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_87
timestamp 1649977179
transform 1 0 9108 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_9_96
timestamp 1649977179
transform 1 0 9936 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_104
timestamp 1649977179
transform 1 0 10672 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_108
timestamp 1649977179
transform 1 0 11040 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_118
timestamp 1649977179
transform 1 0 11960 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_126
timestamp 1649977179
transform 1 0 12696 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_134
timestamp 1649977179
transform 1 0 13432 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_138
timestamp 1649977179
transform 1 0 13800 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_144
timestamp 1649977179
transform 1 0 14352 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_9_164
timestamp 1649977179
transform 1 0 16192 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_169
timestamp 1649977179
transform 1 0 16652 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_176
timestamp 1649977179
transform 1 0 17296 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_183
timestamp 1649977179
transform 1 0 17940 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_190
timestamp 1649977179
transform 1 0 18584 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_197
timestamp 1649977179
transform 1 0 19228 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_211
timestamp 1649977179
transform 1 0 20516 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_220
timestamp 1649977179
transform 1 0 21344 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_225
timestamp 1649977179
transform 1 0 21804 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_229
timestamp 1649977179
transform 1 0 22172 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_9_245
timestamp 1649977179
transform 1 0 23644 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_251
timestamp 1649977179
transform 1 0 24196 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_255
timestamp 1649977179
transform 1 0 24564 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_276
timestamp 1649977179
transform 1 0 26496 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_9_291
timestamp 1649977179
transform 1 0 27876 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_297
timestamp 1649977179
transform 1 0 28428 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_305
timestamp 1649977179
transform 1 0 29164 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_9_323
timestamp 1649977179
transform 1 0 30820 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_9_332
timestamp 1649977179
transform 1 0 31648 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_9_337
timestamp 1649977179
transform 1 0 32108 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_9_352
timestamp 1649977179
transform 1 0 33488 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_356
timestamp 1649977179
transform 1 0 33856 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_360
timestamp 1649977179
transform 1 0 34224 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_367
timestamp 1649977179
transform 1 0 34868 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_9_383
timestamp 1649977179
transform 1 0 36340 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_391
timestamp 1649977179
transform 1 0 37076 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_398
timestamp 1649977179
transform 1 0 37720 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_406
timestamp 1649977179
transform 1 0 38456 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_410
timestamp 1649977179
transform 1 0 38824 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_423
timestamp 1649977179
transform 1 0 40020 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_9_439
timestamp 1649977179
transform 1 0 41492 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_447
timestamp 1649977179
transform 1 0 42228 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_449
timestamp 1649977179
transform 1 0 42412 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_456
timestamp 1649977179
transform 1 0 43056 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_465
timestamp 1649977179
transform 1 0 43884 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_474
timestamp 1649977179
transform 1 0 44712 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_478
timestamp 1649977179
transform 1 0 45080 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_484
timestamp 1649977179
transform 1 0 45632 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_491
timestamp 1649977179
transform 1 0 46276 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_9_498
timestamp 1649977179
transform 1 0 46920 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_9_505
timestamp 1649977179
transform 1 0 47564 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_509
timestamp 1649977179
transform 1 0 47932 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_9_515
timestamp 1649977179
transform 1 0 48484 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_521
timestamp 1649977179
transform 1 0 49036 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_527
timestamp 1649977179
transform 1 0 49588 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_9_547
timestamp 1649977179
transform 1 0 51428 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_551
timestamp 1649977179
transform 1 0 51796 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_556
timestamp 1649977179
transform 1 0 52256 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_9_566
timestamp 1649977179
transform 1 0 53176 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_9_586
timestamp 1649977179
transform 1 0 55016 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_592
timestamp 1649977179
transform 1 0 55568 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_596
timestamp 1649977179
transform 1 0 55936 0 -1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_9_603 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 56580 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_9_615
timestamp 1649977179
transform 1 0 57684 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_620
timestamp 1649977179
transform 1 0 58144 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_624
timestamp 1649977179
transform 1 0 58512 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_3
timestamp 1649977179
transform 1 0 1380 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_7
timestamp 1649977179
transform 1 0 1748 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_11
timestamp 1649977179
transform 1 0 2116 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_10_20
timestamp 1649977179
transform 1 0 2944 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_10_31
timestamp 1649977179
transform 1 0 3956 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_38
timestamp 1649977179
transform 1 0 4600 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_45
timestamp 1649977179
transform 1 0 5244 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_10_61
timestamp 1649977179
transform 1 0 6716 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_69
timestamp 1649977179
transform 1 0 7452 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_73
timestamp 1649977179
transform 1 0 7820 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_80
timestamp 1649977179
transform 1 0 8464 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_85
timestamp 1649977179
transform 1 0 8924 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_89
timestamp 1649977179
transform 1 0 9292 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_105
timestamp 1649977179
transform 1 0 10764 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_109
timestamp 1649977179
transform 1 0 11132 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_113
timestamp 1649977179
transform 1 0 11500 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_129
timestamp 1649977179
transform 1 0 12972 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_136
timestamp 1649977179
transform 1 0 13616 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_141
timestamp 1649977179
transform 1 0 14076 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_145
timestamp 1649977179
transform 1 0 14444 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_10_161
timestamp 1649977179
transform 1 0 15916 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_167
timestamp 1649977179
transform 1 0 16468 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_173
timestamp 1649977179
transform 1 0 17020 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_181
timestamp 1649977179
transform 1 0 17756 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_185
timestamp 1649977179
transform 1 0 18124 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_192
timestamp 1649977179
transform 1 0 18768 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_200
timestamp 1649977179
transform 1 0 19504 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_204
timestamp 1649977179
transform 1 0 19872 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_215
timestamp 1649977179
transform 1 0 20884 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_224
timestamp 1649977179
transform 1 0 21712 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_230
timestamp 1649977179
transform 1 0 22264 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_10_238
timestamp 1649977179
transform 1 0 23000 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_244
timestamp 1649977179
transform 1 0 23552 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_248
timestamp 1649977179
transform 1 0 23920 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_10_258
timestamp 1649977179
transform 1 0 24840 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_264
timestamp 1649977179
transform 1 0 25392 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_270
timestamp 1649977179
transform 1 0 25944 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_276
timestamp 1649977179
transform 1 0 26496 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_283
timestamp 1649977179
transform 1 0 27140 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_292
timestamp 1649977179
transform 1 0 27968 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_303
timestamp 1649977179
transform 1 0 28980 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_307
timestamp 1649977179
transform 1 0 29348 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_309
timestamp 1649977179
transform 1 0 29532 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_317
timestamp 1649977179
transform 1 0 30268 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_323
timestamp 1649977179
transform 1 0 30820 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_330
timestamp 1649977179
transform 1 0 31464 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_339
timestamp 1649977179
transform 1 0 32292 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_346
timestamp 1649977179
transform 1 0 32936 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_353
timestamp 1649977179
transform 1 0 33580 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_360
timestamp 1649977179
transform 1 0 34224 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_10_370
timestamp 1649977179
transform 1 0 35144 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_376
timestamp 1649977179
transform 1 0 35696 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_387
timestamp 1649977179
transform 1 0 36708 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_10_395
timestamp 1649977179
transform 1 0 37444 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_10_406
timestamp 1649977179
transform 1 0 38456 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_415
timestamp 1649977179
transform 1 0 39284 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_419
timestamp 1649977179
transform 1 0 39652 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_421
timestamp 1649977179
transform 1 0 39836 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_10_429
timestamp 1649977179
transform 1 0 40572 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_437
timestamp 1649977179
transform 1 0 41308 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_450
timestamp 1649977179
transform 1 0 42504 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_10_459
timestamp 1649977179
transform 1 0 43332 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_467
timestamp 1649977179
transform 1 0 44068 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_471
timestamp 1649977179
transform 1 0 44436 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_475
timestamp 1649977179
transform 1 0 44804 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_10_477
timestamp 1649977179
transform 1 0 44988 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_10_492
timestamp 1649977179
transform 1 0 46368 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_10_499
timestamp 1649977179
transform 1 0 47012 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_10_510
timestamp 1649977179
transform 1 0 48024 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_519
timestamp 1649977179
transform 1 0 48852 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_528
timestamp 1649977179
transform 1 0 49680 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_545
timestamp 1649977179
transform 1 0 51244 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_551
timestamp 1649977179
transform 1 0 51796 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_557
timestamp 1649977179
transform 1 0 52348 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_563
timestamp 1649977179
transform 1 0 52900 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_569
timestamp 1649977179
transform 1 0 53452 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_573
timestamp 1649977179
transform 1 0 53820 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_577
timestamp 1649977179
transform 1 0 54188 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_583
timestamp 1649977179
transform 1 0 54740 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_587
timestamp 1649977179
transform 1 0 55108 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_591
timestamp 1649977179
transform 1 0 55476 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_603
timestamp 1649977179
transform 1 0 56580 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_615
timestamp 1649977179
transform 1 0 57684 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_623
timestamp 1649977179
transform 1 0 58420 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_3
timestamp 1649977179
transform 1 0 1380 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_8
timestamp 1649977179
transform 1 0 1840 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_11_17
timestamp 1649977179
transform 1 0 2668 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_23
timestamp 1649977179
transform 1 0 3220 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_11_29
timestamp 1649977179
transform 1 0 3772 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_11_40
timestamp 1649977179
transform 1 0 4784 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_48
timestamp 1649977179
transform 1 0 5520 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_52
timestamp 1649977179
transform 1 0 5888 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_69
timestamp 1649977179
transform 1 0 7452 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_11_78
timestamp 1649977179
transform 1 0 8280 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_11_91
timestamp 1649977179
transform 1 0 9476 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_97
timestamp 1649977179
transform 1 0 10028 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_101
timestamp 1649977179
transform 1 0 10396 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_108
timestamp 1649977179
transform 1 0 11040 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_118
timestamp 1649977179
transform 1 0 11960 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_122
timestamp 1649977179
transform 1 0 12328 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_128
timestamp 1649977179
transform 1 0 12880 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_134
timestamp 1649977179
transform 1 0 13432 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_141
timestamp 1649977179
transform 1 0 14076 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_148
timestamp 1649977179
transform 1 0 14720 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_155
timestamp 1649977179
transform 1 0 15364 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_164
timestamp 1649977179
transform 1 0 16192 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_169
timestamp 1649977179
transform 1 0 16652 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_176
timestamp 1649977179
transform 1 0 17296 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_185
timestamp 1649977179
transform 1 0 18124 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_189
timestamp 1649977179
transform 1 0 18492 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_193
timestamp 1649977179
transform 1 0 18860 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_202
timestamp 1649977179
transform 1 0 19688 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_11_218
timestamp 1649977179
transform 1 0 21160 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_11_225
timestamp 1649977179
transform 1 0 21804 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_232
timestamp 1649977179
transform 1 0 22448 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_241
timestamp 1649977179
transform 1 0 23276 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_248
timestamp 1649977179
transform 1 0 23920 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_255
timestamp 1649977179
transform 1 0 24564 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_11_271
timestamp 1649977179
transform 1 0 26036 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_279
timestamp 1649977179
transform 1 0 26772 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_281
timestamp 1649977179
transform 1 0 26956 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_287
timestamp 1649977179
transform 1 0 27508 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_11_300
timestamp 1649977179
transform 1 0 28704 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_310
timestamp 1649977179
transform 1 0 29624 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_319
timestamp 1649977179
transform 1 0 30452 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_326
timestamp 1649977179
transform 1 0 31096 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_332
timestamp 1649977179
transform 1 0 31648 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_11_340
timestamp 1649977179
transform 1 0 32384 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_348
timestamp 1649977179
transform 1 0 33120 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_354
timestamp 1649977179
transform 1 0 33672 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_363
timestamp 1649977179
transform 1 0 34500 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_370
timestamp 1649977179
transform 1 0 35144 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_11_384
timestamp 1649977179
transform 1 0 36432 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_11_395
timestamp 1649977179
transform 1 0 37444 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_404
timestamp 1649977179
transform 1 0 38272 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_413
timestamp 1649977179
transform 1 0 39100 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_420
timestamp 1649977179
transform 1 0 39744 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_427
timestamp 1649977179
transform 1 0 40388 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_431
timestamp 1649977179
transform 1 0 40756 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_444
timestamp 1649977179
transform 1 0 41952 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_454
timestamp 1649977179
transform 1 0 42872 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_461
timestamp 1649977179
transform 1 0 43516 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_11_468
timestamp 1649977179
transform 1 0 44160 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_11_477
timestamp 1649977179
transform 1 0 44988 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_491
timestamp 1649977179
transform 1 0 46276 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_500
timestamp 1649977179
transform 1 0 47104 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_507
timestamp 1649977179
transform 1 0 47748 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_511
timestamp 1649977179
transform 1 0 48116 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_516
timestamp 1649977179
transform 1 0 48576 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_520
timestamp 1649977179
transform 1 0 48944 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_526
timestamp 1649977179
transform 1 0 49496 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_534
timestamp 1649977179
transform 1 0 50232 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_11_541
timestamp 1649977179
transform 1 0 50876 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_11_552
timestamp 1649977179
transform 1 0 51888 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_11_566
timestamp 1649977179
transform 1 0 53176 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_572
timestamp 1649977179
transform 1 0 53728 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_578
timestamp 1649977179
transform 1 0 54280 0 -1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_11_584
timestamp 1649977179
transform 1 0 54832 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_596
timestamp 1649977179
transform 1 0 55936 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_608
timestamp 1649977179
transform 1 0 57040 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_11_617
timestamp 1649977179
transform 1 0 57868 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_3
timestamp 1649977179
transform 1 0 1380 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_8
timestamp 1649977179
transform 1 0 1840 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_15
timestamp 1649977179
transform 1 0 2484 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_24
timestamp 1649977179
transform 1 0 3312 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_29
timestamp 1649977179
transform 1 0 3772 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_34
timestamp 1649977179
transform 1 0 4232 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_50
timestamp 1649977179
transform 1 0 5704 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_57
timestamp 1649977179
transform 1 0 6348 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_64
timestamp 1649977179
transform 1 0 6992 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_80
timestamp 1649977179
transform 1 0 8464 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_85
timestamp 1649977179
transform 1 0 8924 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_90
timestamp 1649977179
transform 1 0 9384 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_97
timestamp 1649977179
transform 1 0 10028 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_106
timestamp 1649977179
transform 1 0 10856 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_122
timestamp 1649977179
transform 1 0 12328 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_129
timestamp 1649977179
transform 1 0 12972 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_136
timestamp 1649977179
transform 1 0 13616 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_141
timestamp 1649977179
transform 1 0 14076 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_154
timestamp 1649977179
transform 1 0 15272 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_161
timestamp 1649977179
transform 1 0 15916 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_170
timestamp 1649977179
transform 1 0 16744 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_186
timestamp 1649977179
transform 1 0 18216 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_192
timestamp 1649977179
transform 1 0 18768 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_197
timestamp 1649977179
transform 1 0 19228 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_204
timestamp 1649977179
transform 1 0 19872 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_213
timestamp 1649977179
transform 1 0 20700 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_219
timestamp 1649977179
transform 1 0 21252 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_226
timestamp 1649977179
transform 1 0 21896 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_242
timestamp 1649977179
transform 1 0 23368 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_248
timestamp 1649977179
transform 1 0 23920 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_253
timestamp 1649977179
transform 1 0 24380 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_257
timestamp 1649977179
transform 1 0 24748 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_261
timestamp 1649977179
transform 1 0 25116 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_268
timestamp 1649977179
transform 1 0 25760 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_275
timestamp 1649977179
transform 1 0 26404 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_12_284
timestamp 1649977179
transform 1 0 27232 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_12_295
timestamp 1649977179
transform 1 0 28244 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_304
timestamp 1649977179
transform 1 0 29072 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_309
timestamp 1649977179
transform 1 0 29532 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_323
timestamp 1649977179
transform 1 0 30820 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_332
timestamp 1649977179
transform 1 0 31648 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_12_338
timestamp 1649977179
transform 1 0 32200 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_12_347
timestamp 1649977179
transform 1 0 33028 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_354
timestamp 1649977179
transform 1 0 33672 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_360
timestamp 1649977179
transform 1 0 34224 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_367
timestamp 1649977179
transform 1 0 34868 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_12_376
timestamp 1649977179
transform 1 0 35696 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_12_389
timestamp 1649977179
transform 1 0 36892 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_393
timestamp 1649977179
transform 1 0 37260 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_399
timestamp 1649977179
transform 1 0 37812 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_406
timestamp 1649977179
transform 1 0 38456 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_410
timestamp 1649977179
transform 1 0 38824 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_416
timestamp 1649977179
transform 1 0 39376 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_426
timestamp 1649977179
transform 1 0 40296 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_433
timestamp 1649977179
transform 1 0 40940 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_440
timestamp 1649977179
transform 1 0 41584 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_447
timestamp 1649977179
transform 1 0 42228 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_463
timestamp 1649977179
transform 1 0 43700 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_472
timestamp 1649977179
transform 1 0 44528 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_479
timestamp 1649977179
transform 1 0 45172 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_483
timestamp 1649977179
transform 1 0 45540 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_496
timestamp 1649977179
transform 1 0 46736 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_502
timestamp 1649977179
transform 1 0 47288 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_506
timestamp 1649977179
transform 1 0 47656 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_512
timestamp 1649977179
transform 1 0 48208 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_528
timestamp 1649977179
transform 1 0 49680 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_533
timestamp 1649977179
transform 1 0 50140 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_541
timestamp 1649977179
transform 1 0 50876 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_12_550
timestamp 1649977179
transform 1 0 51704 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_556
timestamp 1649977179
transform 1 0 52256 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_570
timestamp 1649977179
transform 1 0 53544 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_12_577
timestamp 1649977179
transform 1 0 54188 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_12_585
timestamp 1649977179
transform 1 0 54924 0 1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_12_589
timestamp 1649977179
transform 1 0 55292 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_601
timestamp 1649977179
transform 1 0 56396 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_613
timestamp 1649977179
transform 1 0 57500 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_3
timestamp 1649977179
transform 1 0 1380 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_10
timestamp 1649977179
transform 1 0 2024 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_19
timestamp 1649977179
transform 1 0 2852 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_13_35
timestamp 1649977179
transform 1 0 4324 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_41
timestamp 1649977179
transform 1 0 4876 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_45
timestamp 1649977179
transform 1 0 5244 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_52
timestamp 1649977179
transform 1 0 5888 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_13_62
timestamp 1649977179
transform 1 0 6808 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_70
timestamp 1649977179
transform 1 0 7544 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_76
timestamp 1649977179
transform 1 0 8096 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_92
timestamp 1649977179
transform 1 0 9568 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_98
timestamp 1649977179
transform 1 0 10120 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_107
timestamp 1649977179
transform 1 0 10948 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_111
timestamp 1649977179
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_118
timestamp 1649977179
transform 1 0 11960 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_13_131
timestamp 1649977179
transform 1 0 13156 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_13_142
timestamp 1649977179
transform 1 0 14168 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_151
timestamp 1649977179
transform 1 0 14996 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_13_160
timestamp 1649977179
transform 1 0 15824 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_13_169
timestamp 1649977179
transform 1 0 16652 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_173
timestamp 1649977179
transform 1 0 17020 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_186
timestamp 1649977179
transform 1 0 18216 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_194
timestamp 1649977179
transform 1 0 18952 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_200
timestamp 1649977179
transform 1 0 19504 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_13_216
timestamp 1649977179
transform 1 0 20976 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_225
timestamp 1649977179
transform 1 0 21804 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_232
timestamp 1649977179
transform 1 0 22448 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_241
timestamp 1649977179
transform 1 0 23276 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_247
timestamp 1649977179
transform 1 0 23828 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_254
timestamp 1649977179
transform 1 0 24472 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_13_263
timestamp 1649977179
transform 1 0 25300 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_13_276
timestamp 1649977179
transform 1 0 26496 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_293
timestamp 1649977179
transform 1 0 28060 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_302
timestamp 1649977179
transform 1 0 28888 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_318
timestamp 1649977179
transform 1 0 30360 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_325
timestamp 1649977179
transform 1 0 31004 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_331
timestamp 1649977179
transform 1 0 31556 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_335
timestamp 1649977179
transform 1 0 31924 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_340
timestamp 1649977179
transform 1 0 32384 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_356
timestamp 1649977179
transform 1 0 33856 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_372
timestamp 1649977179
transform 1 0 35328 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_388
timestamp 1649977179
transform 1 0 36800 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_393
timestamp 1649977179
transform 1 0 37260 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_401
timestamp 1649977179
transform 1 0 37996 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_13_408
timestamp 1649977179
transform 1 0 38640 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_13_426
timestamp 1649977179
transform 1 0 40296 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_432
timestamp 1649977179
transform 1 0 40848 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_13_441
timestamp 1649977179
transform 1 0 41676 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_447
timestamp 1649977179
transform 1 0 42228 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_461
timestamp 1649977179
transform 1 0 43516 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_468
timestamp 1649977179
transform 1 0 44160 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_472
timestamp 1649977179
transform 1 0 44528 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_476
timestamp 1649977179
transform 1 0 44896 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_13_489
timestamp 1649977179
transform 1 0 46092 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_13_496
timestamp 1649977179
transform 1 0 46736 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_13_508
timestamp 1649977179
transform 1 0 47840 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_512
timestamp 1649977179
transform 1 0 48208 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_516
timestamp 1649977179
transform 1 0 48576 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_533
timestamp 1649977179
transform 1 0 50140 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_13_539
timestamp 1649977179
transform 1 0 50692 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_545
timestamp 1649977179
transform 1 0 51244 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_549
timestamp 1649977179
transform 1 0 51612 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_556
timestamp 1649977179
transform 1 0 52256 0 -1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_13_574
timestamp 1649977179
transform 1 0 53912 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_586
timestamp 1649977179
transform 1 0 55016 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_598
timestamp 1649977179
transform 1 0 56120 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_610
timestamp 1649977179
transform 1 0 57224 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_13_617
timestamp 1649977179
transform 1 0 57868 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_14_3
timestamp 1649977179
transform 1 0 1380 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_14_9
timestamp 1649977179
transform 1 0 1932 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_16
timestamp 1649977179
transform 1 0 2576 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_23
timestamp 1649977179
transform 1 0 3220 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_27
timestamp 1649977179
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_14_41
timestamp 1649977179
transform 1 0 4876 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_14_52
timestamp 1649977179
transform 1 0 5888 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_14_68
timestamp 1649977179
transform 1 0 7360 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_76
timestamp 1649977179
transform 1 0 8096 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_80
timestamp 1649977179
transform 1 0 8464 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_85
timestamp 1649977179
transform 1 0 8924 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_89
timestamp 1649977179
transform 1 0 9292 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_93
timestamp 1649977179
transform 1 0 9660 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_100
timestamp 1649977179
transform 1 0 10304 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_107
timestamp 1649977179
transform 1 0 10948 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_114
timestamp 1649977179
transform 1 0 11592 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_130
timestamp 1649977179
transform 1 0 13064 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_136
timestamp 1649977179
transform 1 0 13616 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_14_144
timestamp 1649977179
transform 1 0 14352 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_14_162
timestamp 1649977179
transform 1 0 16008 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_166
timestamp 1649977179
transform 1 0 16376 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_170
timestamp 1649977179
transform 1 0 16744 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_177
timestamp 1649977179
transform 1 0 17388 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_181
timestamp 1649977179
transform 1 0 17756 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_185
timestamp 1649977179
transform 1 0 18124 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_192
timestamp 1649977179
transform 1 0 18768 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_197
timestamp 1649977179
transform 1 0 19228 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_201
timestamp 1649977179
transform 1 0 19596 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_214
timestamp 1649977179
transform 1 0 20792 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_221
timestamp 1649977179
transform 1 0 21436 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_225
timestamp 1649977179
transform 1 0 21804 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_229
timestamp 1649977179
transform 1 0 22172 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_14_245
timestamp 1649977179
transform 1 0 23644 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_251
timestamp 1649977179
transform 1 0 24196 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_14_265
timestamp 1649977179
transform 1 0 25484 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_271
timestamp 1649977179
transform 1 0 26036 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_284
timestamp 1649977179
transform 1 0 27232 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_290
timestamp 1649977179
transform 1 0 27784 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_294
timestamp 1649977179
transform 1 0 28152 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_297
timestamp 1649977179
transform 1 0 28428 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_303
timestamp 1649977179
transform 1 0 28980 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_307
timestamp 1649977179
transform 1 0 29348 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_311
timestamp 1649977179
transform 1 0 29716 0 1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_14_327
timestamp 1649977179
transform 1 0 31188 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_14_339
timestamp 1649977179
transform 1 0 32292 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_14_344
timestamp 1649977179
transform 1 0 32752 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_360
timestamp 1649977179
transform 1 0 34224 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_367
timestamp 1649977179
transform 1 0 34868 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_14_373
timestamp 1649977179
transform 1 0 35420 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_14_385
timestamp 1649977179
transform 1 0 36524 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_393
timestamp 1649977179
transform 1 0 37260 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_406
timestamp 1649977179
transform 1 0 38456 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_14_412
timestamp 1649977179
transform 1 0 39008 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_14_423
timestamp 1649977179
transform 1 0 40020 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_429
timestamp 1649977179
transform 1 0 40572 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_433
timestamp 1649977179
transform 1 0 40940 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_14_436
timestamp 1649977179
transform 1 0 41216 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_444
timestamp 1649977179
transform 1 0 41952 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_448
timestamp 1649977179
transform 1 0 42320 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_464
timestamp 1649977179
transform 1 0 43792 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_14_470
timestamp 1649977179
transform 1 0 44344 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_14_479
timestamp 1649977179
transform 1 0 45172 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_483
timestamp 1649977179
transform 1 0 45540 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_14_497
timestamp 1649977179
transform 1 0 46828 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_14_516
timestamp 1649977179
transform 1 0 48576 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_520
timestamp 1649977179
transform 1 0 48944 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_14_524
timestamp 1649977179
transform 1 0 49312 0 1 9792
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_14_533
timestamp 1649977179
transform 1 0 50140 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_545
timestamp 1649977179
transform 1 0 51244 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_14_553
timestamp 1649977179
transform 1 0 51980 0 1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_14_569
timestamp 1649977179
transform 1 0 53452 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_581
timestamp 1649977179
transform 1 0 54556 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_587
timestamp 1649977179
transform 1 0 55108 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_589
timestamp 1649977179
transform 1 0 55292 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_601
timestamp 1649977179
transform 1 0 56396 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_613
timestamp 1649977179
transform 1 0 57500 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_15_3
timestamp 1649977179
transform 1 0 1380 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_8
timestamp 1649977179
transform 1 0 1840 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_15_15
timestamp 1649977179
transform 1 0 2484 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_15_25
timestamp 1649977179
transform 1 0 3404 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_15_32
timestamp 1649977179
transform 1 0 4048 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_38
timestamp 1649977179
transform 1 0 4600 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_42
timestamp 1649977179
transform 1 0 4968 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_15_52
timestamp 1649977179
transform 1 0 5888 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_59
timestamp 1649977179
transform 1 0 6532 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_66
timestamp 1649977179
transform 1 0 7176 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_73
timestamp 1649977179
transform 1 0 7820 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_80
timestamp 1649977179
transform 1 0 8464 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_86
timestamp 1649977179
transform 1 0 9016 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_15_93
timestamp 1649977179
transform 1 0 9660 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_15_102
timestamp 1649977179
transform 1 0 10488 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_108
timestamp 1649977179
transform 1 0 11040 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_15_125
timestamp 1649977179
transform 1 0 12604 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_15_136
timestamp 1649977179
transform 1 0 13616 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_143
timestamp 1649977179
transform 1 0 14260 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_150
timestamp 1649977179
transform 1 0 14904 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_157
timestamp 1649977179
transform 1 0 15548 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_164
timestamp 1649977179
transform 1 0 16192 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_172
timestamp 1649977179
transform 1 0 16928 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_176
timestamp 1649977179
transform 1 0 17296 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_15_189
timestamp 1649977179
transform 1 0 18492 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_195
timestamp 1649977179
transform 1 0 19044 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_198
timestamp 1649977179
transform 1 0 19320 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_207
timestamp 1649977179
transform 1 0 20148 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_214
timestamp 1649977179
transform 1 0 20792 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_220
timestamp 1649977179
transform 1 0 21344 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_15_225
timestamp 1649977179
transform 1 0 21804 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_15_230
timestamp 1649977179
transform 1 0 22264 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_15_237
timestamp 1649977179
transform 1 0 22908 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_15_246
timestamp 1649977179
transform 1 0 23736 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_254
timestamp 1649977179
transform 1 0 24472 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_257
timestamp 1649977179
transform 1 0 24748 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_265
timestamp 1649977179
transform 1 0 25484 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_269
timestamp 1649977179
transform 1 0 25852 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_275
timestamp 1649977179
transform 1 0 26404 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_279
timestamp 1649977179
transform 1 0 26772 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_284
timestamp 1649977179
transform 1 0 27232 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_15_294
timestamp 1649977179
transform 1 0 28152 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_15_302
timestamp 1649977179
transform 1 0 28888 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_306
timestamp 1649977179
transform 1 0 29256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_310
timestamp 1649977179
transform 1 0 29624 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_316
timestamp 1649977179
transform 1 0 30176 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_15_322
timestamp 1649977179
transform 1 0 30728 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_15_334
timestamp 1649977179
transform 1 0 31832 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_15_337
timestamp 1649977179
transform 1 0 32108 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_15_349
timestamp 1649977179
transform 1 0 33212 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_352
timestamp 1649977179
transform 1 0 33488 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_358
timestamp 1649977179
transform 1 0 34040 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_362
timestamp 1649977179
transform 1 0 34408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_365
timestamp 1649977179
transform 1 0 34684 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_15_375
timestamp 1649977179
transform 1 0 35604 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_381
timestamp 1649977179
transform 1 0 36156 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_387
timestamp 1649977179
transform 1 0 36708 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_391
timestamp 1649977179
transform 1 0 37076 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_395
timestamp 1649977179
transform 1 0 37444 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_401
timestamp 1649977179
transform 1 0 37996 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_407
timestamp 1649977179
transform 1 0 38548 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_413
timestamp 1649977179
transform 1 0 39100 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_419
timestamp 1649977179
transform 1 0 39652 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_425
timestamp 1649977179
transform 1 0 40204 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_431
timestamp 1649977179
transform 1 0 40756 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_437
timestamp 1649977179
transform 1 0 41308 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_441
timestamp 1649977179
transform 1 0 41676 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_444
timestamp 1649977179
transform 1 0 41952 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_451
timestamp 1649977179
transform 1 0 42596 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_15_457
timestamp 1649977179
transform 1 0 43148 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_15_467
timestamp 1649977179
transform 1 0 44068 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_15_473
timestamp 1649977179
transform 1 0 44620 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_479
timestamp 1649977179
transform 1 0 45172 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_482
timestamp 1649977179
transform 1 0 45448 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_488
timestamp 1649977179
transform 1 0 46000 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_494
timestamp 1649977179
transform 1 0 46552 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_500
timestamp 1649977179
transform 1 0 47104 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_508
timestamp 1649977179
transform 1 0 47840 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_514
timestamp 1649977179
transform 1 0 48392 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_15_520
timestamp 1649977179
transform 1 0 48944 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_532
timestamp 1649977179
transform 1 0 50048 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_544
timestamp 1649977179
transform 1 0 51152 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_556
timestamp 1649977179
transform 1 0 52256 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_15_561
timestamp 1649977179
transform 1 0 52716 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_573
timestamp 1649977179
transform 1 0 53820 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_585
timestamp 1649977179
transform 1 0 54924 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_597
timestamp 1649977179
transform 1 0 56028 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_609
timestamp 1649977179
transform 1 0 57132 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_615
timestamp 1649977179
transform 1 0 57684 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_617
timestamp 1649977179
transform 1 0 57868 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_16_3
timestamp 1649977179
transform 1 0 1380 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_7
timestamp 1649977179
transform 1 0 1748 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_11
timestamp 1649977179
transform 1 0 2116 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_17
timestamp 1649977179
transform 1 0 2668 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_23
timestamp 1649977179
transform 1 0 3220 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_27
timestamp 1649977179
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_16_29
timestamp 1649977179
transform 1 0 3772 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_16_34
timestamp 1649977179
transform 1 0 4232 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_16_42
timestamp 1649977179
transform 1 0 4968 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_50
timestamp 1649977179
transform 1 0 5704 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_53
timestamp 1649977179
transform 1 0 5980 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_59
timestamp 1649977179
transform 1 0 6532 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_16_66
timestamp 1649977179
transform 1 0 7176 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_16_75
timestamp 1649977179
transform 1 0 8004 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_83
timestamp 1649977179
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_85
timestamp 1649977179
transform 1 0 8924 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_89
timestamp 1649977179
transform 1 0 9292 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_93
timestamp 1649977179
transform 1 0 9660 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_16_99
timestamp 1649977179
transform 1 0 10212 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_16_109
timestamp 1649977179
transform 1 0 11132 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_115
timestamp 1649977179
transform 1 0 11684 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_122
timestamp 1649977179
transform 1 0 12328 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_129
timestamp 1649977179
transform 1 0 12972 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_136
timestamp 1649977179
transform 1 0 13616 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_144
timestamp 1649977179
transform 1 0 14352 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_148
timestamp 1649977179
transform 1 0 14720 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_152
timestamp 1649977179
transform 1 0 15088 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_159
timestamp 1649977179
transform 1 0 15732 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_166
timestamp 1649977179
transform 1 0 16376 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_173
timestamp 1649977179
transform 1 0 17020 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_179
timestamp 1649977179
transform 1 0 17572 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_185
timestamp 1649977179
transform 1 0 18124 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_189
timestamp 1649977179
transform 1 0 18492 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_192
timestamp 1649977179
transform 1 0 18768 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_16_199
timestamp 1649977179
transform 1 0 19412 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_16_209
timestamp 1649977179
transform 1 0 20332 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_16_217
timestamp 1649977179
transform 1 0 21068 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_223
timestamp 1649977179
transform 1 0 21620 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_227
timestamp 1649977179
transform 1 0 21988 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_230
timestamp 1649977179
transform 1 0 22264 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_236
timestamp 1649977179
transform 1 0 22816 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_242
timestamp 1649977179
transform 1 0 23368 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_248
timestamp 1649977179
transform 1 0 23920 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_253
timestamp 1649977179
transform 1 0 24380 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_257
timestamp 1649977179
transform 1 0 24748 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_260
timestamp 1649977179
transform 1 0 25024 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_266
timestamp 1649977179
transform 1 0 25576 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_272
timestamp 1649977179
transform 1 0 26128 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_16_278
timestamp 1649977179
transform 1 0 26680 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_16_286
timestamp 1649977179
transform 1 0 27416 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_16_292
timestamp 1649977179
transform 1 0 27968 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_298
timestamp 1649977179
transform 1 0 28520 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_16_301
timestamp 1649977179
transform 1 0 28796 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_307
timestamp 1649977179
transform 1 0 29348 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_311
timestamp 1649977179
transform 1 0 29716 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_323
timestamp 1649977179
transform 1 0 30820 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_335
timestamp 1649977179
transform 1 0 31924 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_347
timestamp 1649977179
transform 1 0 33028 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_359
timestamp 1649977179
transform 1 0 34132 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_363
timestamp 1649977179
transform 1 0 34500 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_365
timestamp 1649977179
transform 1 0 34684 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_371
timestamp 1649977179
transform 1 0 35236 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_377
timestamp 1649977179
transform 1 0 35788 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_383
timestamp 1649977179
transform 1 0 36340 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_16_389
timestamp 1649977179
transform 1 0 36892 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_16_397
timestamp 1649977179
transform 1 0 37628 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_403
timestamp 1649977179
transform 1 0 38180 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_409
timestamp 1649977179
transform 1 0 38732 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_415
timestamp 1649977179
transform 1 0 39284 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_419
timestamp 1649977179
transform 1 0 39652 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_423
timestamp 1649977179
transform 1 0 40020 0 1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_16_429
timestamp 1649977179
transform 1 0 40572 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_16_441
timestamp 1649977179
transform 1 0 41676 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_16_445
timestamp 1649977179
transform 1 0 42044 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_16_453
timestamp 1649977179
transform 1 0 42780 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_16_461
timestamp 1649977179
transform 1 0 43516 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_16_467
timestamp 1649977179
transform 1 0 44068 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_475
timestamp 1649977179
transform 1 0 44804 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_479
timestamp 1649977179
transform 1 0 45172 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_491
timestamp 1649977179
transform 1 0 46276 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_503
timestamp 1649977179
transform 1 0 47380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_515
timestamp 1649977179
transform 1 0 48484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_527
timestamp 1649977179
transform 1 0 49588 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_531
timestamp 1649977179
transform 1 0 49956 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_533
timestamp 1649977179
transform 1 0 50140 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_545
timestamp 1649977179
transform 1 0 51244 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_557
timestamp 1649977179
transform 1 0 52348 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_569
timestamp 1649977179
transform 1 0 53452 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_581
timestamp 1649977179
transform 1 0 54556 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_587
timestamp 1649977179
transform 1 0 55108 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_589
timestamp 1649977179
transform 1 0 55292 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_601
timestamp 1649977179
transform 1 0 56396 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_613
timestamp 1649977179
transform 1 0 57500 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_3
timestamp 1649977179
transform 1 0 1380 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_7
timestamp 1649977179
transform 1 0 1748 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_10
timestamp 1649977179
transform 1 0 2024 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_18
timestamp 1649977179
transform 1 0 2760 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_21
timestamp 1649977179
transform 1 0 3036 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_27
timestamp 1649977179
transform 1 0 3588 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_17_33
timestamp 1649977179
transform 1 0 4140 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_39
timestamp 1649977179
transform 1 0 4692 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_42
timestamp 1649977179
transform 1 0 4968 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_17_52
timestamp 1649977179
transform 1 0 5888 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_57
timestamp 1649977179
transform 1 0 6348 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_61
timestamp 1649977179
transform 1 0 6716 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_17_64
timestamp 1649977179
transform 1 0 6992 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_17_72
timestamp 1649977179
transform 1 0 7728 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_78
timestamp 1649977179
transform 1 0 8280 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_84
timestamp 1649977179
transform 1 0 8832 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_90
timestamp 1649977179
transform 1 0 9384 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_96
timestamp 1649977179
transform 1 0 9936 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_102
timestamp 1649977179
transform 1 0 10488 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_108
timestamp 1649977179
transform 1 0 11040 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_17_113
timestamp 1649977179
transform 1 0 11500 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_17_118
timestamp 1649977179
transform 1 0 11960 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_124
timestamp 1649977179
transform 1 0 12512 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_131
timestamp 1649977179
transform 1 0 13156 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_17_137
timestamp 1649977179
transform 1 0 13708 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_145
timestamp 1649977179
transform 1 0 14444 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_148
timestamp 1649977179
transform 1 0 14720 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_17_155
timestamp 1649977179
transform 1 0 15364 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_17_164
timestamp 1649977179
transform 1 0 16192 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_171
timestamp 1649977179
transform 1 0 16836 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_17_177
timestamp 1649977179
transform 1 0 17388 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_17_187
timestamp 1649977179
transform 1 0 18308 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_193
timestamp 1649977179
transform 1 0 18860 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_17_199
timestamp 1649977179
transform 1 0 19412 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_17_207
timestamp 1649977179
transform 1 0 20148 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_213
timestamp 1649977179
transform 1 0 20700 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_217
timestamp 1649977179
transform 1 0 21068 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_220
timestamp 1649977179
transform 1 0 21344 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_225
timestamp 1649977179
transform 1 0 21804 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_229
timestamp 1649977179
transform 1 0 22172 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_235
timestamp 1649977179
transform 1 0 22724 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_241
timestamp 1649977179
transform 1 0 23276 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_17_247
timestamp 1649977179
transform 1 0 23828 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_253
timestamp 1649977179
transform 1 0 24380 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_256
timestamp 1649977179
transform 1 0 24656 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_262
timestamp 1649977179
transform 1 0 25208 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_268
timestamp 1649977179
transform 1 0 25760 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_17_274
timestamp 1649977179
transform 1 0 26312 0 -1 11968
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_17_281
timestamp 1649977179
transform 1 0 26956 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_293
timestamp 1649977179
transform 1 0 28060 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_305
timestamp 1649977179
transform 1 0 29164 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_317
timestamp 1649977179
transform 1 0 30268 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_329
timestamp 1649977179
transform 1 0 31372 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_335
timestamp 1649977179
transform 1 0 31924 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_337
timestamp 1649977179
transform 1 0 32108 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_349
timestamp 1649977179
transform 1 0 33212 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_361
timestamp 1649977179
transform 1 0 34316 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_17_373
timestamp 1649977179
transform 1 0 35420 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_17_377
timestamp 1649977179
transform 1 0 35788 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_383
timestamp 1649977179
transform 1 0 36340 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_17_386
timestamp 1649977179
transform 1 0 36616 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_17_395
timestamp 1649977179
transform 1 0 37444 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_401
timestamp 1649977179
transform 1 0 37996 0 -1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_17_407
timestamp 1649977179
transform 1 0 38548 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_419
timestamp 1649977179
transform 1 0 39652 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_431
timestamp 1649977179
transform 1 0 40756 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_443
timestamp 1649977179
transform 1 0 41860 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_447
timestamp 1649977179
transform 1 0 42228 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_449
timestamp 1649977179
transform 1 0 42412 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_455
timestamp 1649977179
transform 1 0 42964 0 -1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_17_461
timestamp 1649977179
transform 1 0 43516 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_473
timestamp 1649977179
transform 1 0 44620 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_485
timestamp 1649977179
transform 1 0 45724 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_497
timestamp 1649977179
transform 1 0 46828 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_503
timestamp 1649977179
transform 1 0 47380 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_505
timestamp 1649977179
transform 1 0 47564 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_517
timestamp 1649977179
transform 1 0 48668 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_529
timestamp 1649977179
transform 1 0 49772 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_541
timestamp 1649977179
transform 1 0 50876 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_553
timestamp 1649977179
transform 1 0 51980 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_559
timestamp 1649977179
transform 1 0 52532 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_561
timestamp 1649977179
transform 1 0 52716 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_573
timestamp 1649977179
transform 1 0 53820 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_585
timestamp 1649977179
transform 1 0 54924 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_597
timestamp 1649977179
transform 1 0 56028 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_609
timestamp 1649977179
transform 1 0 57132 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_615
timestamp 1649977179
transform 1 0 57684 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_617
timestamp 1649977179
transform 1 0 57868 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_18_5
timestamp 1649977179
transform 1 0 1564 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_11
timestamp 1649977179
transform 1 0 2116 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_17
timestamp 1649977179
transform 1 0 2668 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_23
timestamp 1649977179
transform 1 0 3220 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp 1649977179
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_31
timestamp 1649977179
transform 1 0 3956 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_18_37
timestamp 1649977179
transform 1 0 4508 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_43
timestamp 1649977179
transform 1 0 5060 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_46
timestamp 1649977179
transform 1 0 5336 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_18_52
timestamp 1649977179
transform 1 0 5888 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_58
timestamp 1649977179
transform 1 0 6440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_61
timestamp 1649977179
transform 1 0 6716 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_67
timestamp 1649977179
transform 1 0 7268 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_73
timestamp 1649977179
transform 1 0 7820 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_77
timestamp 1649977179
transform 1 0 8188 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_80
timestamp 1649977179
transform 1 0 8464 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_85
timestamp 1649977179
transform 1 0 8924 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_18_89
timestamp 1649977179
transform 1 0 9292 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_95
timestamp 1649977179
transform 1 0 9844 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_98
timestamp 1649977179
transform 1 0 10120 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_102
timestamp 1649977179
transform 1 0 10488 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_105
timestamp 1649977179
transform 1 0 10764 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_109
timestamp 1649977179
transform 1 0 11132 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_18_112
timestamp 1649977179
transform 1 0 11408 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_18_120
timestamp 1649977179
transform 1 0 12144 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_128
timestamp 1649977179
transform 1 0 12880 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_131
timestamp 1649977179
transform 1 0 13156 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_139
timestamp 1649977179
transform 1 0 13892 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_143
timestamp 1649977179
transform 1 0 14260 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_18_153
timestamp 1649977179
transform 1 0 15180 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_159
timestamp 1649977179
transform 1 0 15732 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_163
timestamp 1649977179
transform 1 0 16100 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_18_166
timestamp 1649977179
transform 1 0 16376 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_172
timestamp 1649977179
transform 1 0 16928 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_175
timestamp 1649977179
transform 1 0 17204 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_18_185
timestamp 1649977179
transform 1 0 18124 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_191
timestamp 1649977179
transform 1 0 18676 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_195
timestamp 1649977179
transform 1 0 19044 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_199
timestamp 1649977179
transform 1 0 19412 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_207
timestamp 1649977179
transform 1 0 20148 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_210
timestamp 1649977179
transform 1 0 20424 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_216
timestamp 1649977179
transform 1 0 20976 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_18_222
timestamp 1649977179
transform 1 0 21528 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_228
timestamp 1649977179
transform 1 0 22080 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_231
timestamp 1649977179
transform 1 0 22356 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_18_241
timestamp 1649977179
transform 1 0 23276 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_247
timestamp 1649977179
transform 1 0 23828 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_251
timestamp 1649977179
transform 1 0 24196 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_255
timestamp 1649977179
transform 1 0 24564 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_259
timestamp 1649977179
transform 1 0 24932 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_262
timestamp 1649977179
transform 1 0 25208 0 1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_18_268
timestamp 1649977179
transform 1 0 25760 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_280
timestamp 1649977179
transform 1 0 26864 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_292
timestamp 1649977179
transform 1 0 27968 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_304
timestamp 1649977179
transform 1 0 29072 0 1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_18_309
timestamp 1649977179
transform 1 0 29532 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_321
timestamp 1649977179
transform 1 0 30636 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_333
timestamp 1649977179
transform 1 0 31740 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_345
timestamp 1649977179
transform 1 0 32844 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_357
timestamp 1649977179
transform 1 0 33948 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_363
timestamp 1649977179
transform 1 0 34500 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_365
timestamp 1649977179
transform 1 0 34684 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_377
timestamp 1649977179
transform 1 0 35788 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_18_389
timestamp 1649977179
transform 1 0 36892 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_18_393
timestamp 1649977179
transform 1 0 37260 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_405
timestamp 1649977179
transform 1 0 38364 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_18_417
timestamp 1649977179
transform 1 0 39468 0 1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_18_421
timestamp 1649977179
transform 1 0 39836 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_433
timestamp 1649977179
transform 1 0 40940 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_445
timestamp 1649977179
transform 1 0 42044 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_457
timestamp 1649977179
transform 1 0 43148 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_469
timestamp 1649977179
transform 1 0 44252 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_475
timestamp 1649977179
transform 1 0 44804 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_477
timestamp 1649977179
transform 1 0 44988 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_489
timestamp 1649977179
transform 1 0 46092 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_501
timestamp 1649977179
transform 1 0 47196 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_513
timestamp 1649977179
transform 1 0 48300 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_525
timestamp 1649977179
transform 1 0 49404 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_531
timestamp 1649977179
transform 1 0 49956 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_533
timestamp 1649977179
transform 1 0 50140 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_545
timestamp 1649977179
transform 1 0 51244 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_557
timestamp 1649977179
transform 1 0 52348 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_569
timestamp 1649977179
transform 1 0 53452 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_581
timestamp 1649977179
transform 1 0 54556 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_587
timestamp 1649977179
transform 1 0 55108 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_589
timestamp 1649977179
transform 1 0 55292 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_601
timestamp 1649977179
transform 1 0 56396 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_613
timestamp 1649977179
transform 1 0 57500 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_3
timestamp 1649977179
transform 1 0 1380 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_7
timestamp 1649977179
transform 1 0 1748 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_10
timestamp 1649977179
transform 1 0 2024 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_16
timestamp 1649977179
transform 1 0 2576 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_22
timestamp 1649977179
transform 1 0 3128 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_28
timestamp 1649977179
transform 1 0 3680 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_34
timestamp 1649977179
transform 1 0 4232 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_40
timestamp 1649977179
transform 1 0 4784 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_46
timestamp 1649977179
transform 1 0 5336 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_52
timestamp 1649977179
transform 1 0 5888 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_57
timestamp 1649977179
transform 1 0 6348 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_60
timestamp 1649977179
transform 1 0 6624 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_19_66
timestamp 1649977179
transform 1 0 7176 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_19_74
timestamp 1649977179
transform 1 0 7912 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_80
timestamp 1649977179
transform 1 0 8464 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_86
timestamp 1649977179
transform 1 0 9016 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_90
timestamp 1649977179
transform 1 0 9384 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_19_93
timestamp 1649977179
transform 1 0 9660 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_99
timestamp 1649977179
transform 1 0 10212 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_102
timestamp 1649977179
transform 1 0 10488 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_108
timestamp 1649977179
transform 1 0 11040 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_115
timestamp 1649977179
transform 1 0 11684 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_119
timestamp 1649977179
transform 1 0 12052 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_19_122
timestamp 1649977179
transform 1 0 12328 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_128
timestamp 1649977179
transform 1 0 12880 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_131
timestamp 1649977179
transform 1 0 13156 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_19_137
timestamp 1649977179
transform 1 0 13708 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_19_147
timestamp 1649977179
transform 1 0 14628 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_19_153
timestamp 1649977179
transform 1 0 15180 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_161
timestamp 1649977179
transform 1 0 15916 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_164
timestamp 1649977179
transform 1 0 16192 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_169
timestamp 1649977179
transform 1 0 16652 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_175
timestamp 1649977179
transform 1 0 17204 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_181
timestamp 1649977179
transform 1 0 17756 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_187
timestamp 1649977179
transform 1 0 18308 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_193
timestamp 1649977179
transform 1 0 18860 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_199
timestamp 1649977179
transform 1 0 19412 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_19_205
timestamp 1649977179
transform 1 0 19964 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_211
timestamp 1649977179
transform 1 0 20516 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_214
timestamp 1649977179
transform 1 0 20792 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_220
timestamp 1649977179
transform 1 0 21344 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_19_227
timestamp 1649977179
transform 1 0 21988 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_19_235
timestamp 1649977179
transform 1 0 22724 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_241
timestamp 1649977179
transform 1 0 23276 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_244
timestamp 1649977179
transform 1 0 23552 0 -1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_19_250
timestamp 1649977179
transform 1 0 24104 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_262
timestamp 1649977179
transform 1 0 25208 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_274
timestamp 1649977179
transform 1 0 26312 0 -1 13056
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_19_281
timestamp 1649977179
transform 1 0 26956 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_293
timestamp 1649977179
transform 1 0 28060 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_305
timestamp 1649977179
transform 1 0 29164 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_317
timestamp 1649977179
transform 1 0 30268 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_329
timestamp 1649977179
transform 1 0 31372 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_335
timestamp 1649977179
transform 1 0 31924 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_337
timestamp 1649977179
transform 1 0 32108 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_349
timestamp 1649977179
transform 1 0 33212 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_361
timestamp 1649977179
transform 1 0 34316 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_373
timestamp 1649977179
transform 1 0 35420 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_385
timestamp 1649977179
transform 1 0 36524 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_391
timestamp 1649977179
transform 1 0 37076 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_393
timestamp 1649977179
transform 1 0 37260 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_405
timestamp 1649977179
transform 1 0 38364 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_417
timestamp 1649977179
transform 1 0 39468 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_429
timestamp 1649977179
transform 1 0 40572 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_441
timestamp 1649977179
transform 1 0 41676 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_447
timestamp 1649977179
transform 1 0 42228 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_449
timestamp 1649977179
transform 1 0 42412 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_461
timestamp 1649977179
transform 1 0 43516 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_473
timestamp 1649977179
transform 1 0 44620 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_485
timestamp 1649977179
transform 1 0 45724 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_497
timestamp 1649977179
transform 1 0 46828 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_503
timestamp 1649977179
transform 1 0 47380 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_505
timestamp 1649977179
transform 1 0 47564 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_517
timestamp 1649977179
transform 1 0 48668 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_529
timestamp 1649977179
transform 1 0 49772 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_541
timestamp 1649977179
transform 1 0 50876 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_553
timestamp 1649977179
transform 1 0 51980 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_559
timestamp 1649977179
transform 1 0 52532 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_561
timestamp 1649977179
transform 1 0 52716 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_573
timestamp 1649977179
transform 1 0 53820 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_585
timestamp 1649977179
transform 1 0 54924 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_597
timestamp 1649977179
transform 1 0 56028 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_609
timestamp 1649977179
transform 1 0 57132 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_615
timestamp 1649977179
transform 1 0 57684 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_617
timestamp 1649977179
transform 1 0 57868 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_20_3
timestamp 1649977179
transform 1 0 1380 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_9
timestamp 1649977179
transform 1 0 1932 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_12
timestamp 1649977179
transform 1 0 2208 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_18
timestamp 1649977179
transform 1 0 2760 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_24
timestamp 1649977179
transform 1 0 3312 0 1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_20_31
timestamp 1649977179
transform 1 0 3956 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_43
timestamp 1649977179
transform 1 0 5060 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_20_46
timestamp 1649977179
transform 1 0 5336 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_20_54
timestamp 1649977179
transform 1 0 6072 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_60
timestamp 1649977179
transform 1 0 6624 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_63
timestamp 1649977179
transform 1 0 6900 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_75
timestamp 1649977179
transform 1 0 8004 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_83
timestamp 1649977179
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_85
timestamp 1649977179
transform 1 0 8924 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_91
timestamp 1649977179
transform 1 0 9476 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_97
timestamp 1649977179
transform 1 0 10028 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_20_107
timestamp 1649977179
transform 1 0 10948 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_113
timestamp 1649977179
transform 1 0 11500 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_20_119
timestamp 1649977179
transform 1 0 12052 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_20_127
timestamp 1649977179
transform 1 0 12788 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_20_133
timestamp 1649977179
transform 1 0 13340 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_139
timestamp 1649977179
transform 1 0 13892 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_143
timestamp 1649977179
transform 1 0 14260 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_20_153
timestamp 1649977179
transform 1 0 15180 0 1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_20_159
timestamp 1649977179
transform 1 0 15732 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_173
timestamp 1649977179
transform 1 0 17020 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_179
timestamp 1649977179
transform 1 0 17572 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_182
timestamp 1649977179
transform 1 0 17848 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_188
timestamp 1649977179
transform 1 0 18400 0 1 13056
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_20_197
timestamp 1649977179
transform 1 0 19228 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_209
timestamp 1649977179
transform 1 0 20332 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_221
timestamp 1649977179
transform 1 0 21436 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_229
timestamp 1649977179
transform 1 0 22172 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_232
timestamp 1649977179
transform 1 0 22448 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_244
timestamp 1649977179
transform 1 0 23552 0 1 13056
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_20_253
timestamp 1649977179
transform 1 0 24380 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_265
timestamp 1649977179
transform 1 0 25484 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_277
timestamp 1649977179
transform 1 0 26588 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_289
timestamp 1649977179
transform 1 0 27692 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_301
timestamp 1649977179
transform 1 0 28796 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_307
timestamp 1649977179
transform 1 0 29348 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_309
timestamp 1649977179
transform 1 0 29532 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_321
timestamp 1649977179
transform 1 0 30636 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_333
timestamp 1649977179
transform 1 0 31740 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_345
timestamp 1649977179
transform 1 0 32844 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_357
timestamp 1649977179
transform 1 0 33948 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_363
timestamp 1649977179
transform 1 0 34500 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_365
timestamp 1649977179
transform 1 0 34684 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_377
timestamp 1649977179
transform 1 0 35788 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_389
timestamp 1649977179
transform 1 0 36892 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_401
timestamp 1649977179
transform 1 0 37996 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_413
timestamp 1649977179
transform 1 0 39100 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_419
timestamp 1649977179
transform 1 0 39652 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_421
timestamp 1649977179
transform 1 0 39836 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_433
timestamp 1649977179
transform 1 0 40940 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_445
timestamp 1649977179
transform 1 0 42044 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_457
timestamp 1649977179
transform 1 0 43148 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_469
timestamp 1649977179
transform 1 0 44252 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_475
timestamp 1649977179
transform 1 0 44804 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_477
timestamp 1649977179
transform 1 0 44988 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_489
timestamp 1649977179
transform 1 0 46092 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_501
timestamp 1649977179
transform 1 0 47196 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_513
timestamp 1649977179
transform 1 0 48300 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_525
timestamp 1649977179
transform 1 0 49404 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_531
timestamp 1649977179
transform 1 0 49956 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_533
timestamp 1649977179
transform 1 0 50140 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_545
timestamp 1649977179
transform 1 0 51244 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_557
timestamp 1649977179
transform 1 0 52348 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_569
timestamp 1649977179
transform 1 0 53452 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_581
timestamp 1649977179
transform 1 0 54556 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_587
timestamp 1649977179
transform 1 0 55108 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_589
timestamp 1649977179
transform 1 0 55292 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_601
timestamp 1649977179
transform 1 0 56396 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_613
timestamp 1649977179
transform 1 0 57500 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_3
timestamp 1649977179
transform 1 0 1380 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_15
timestamp 1649977179
transform 1 0 2484 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_23
timestamp 1649977179
transform 1 0 3220 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_26
timestamp 1649977179
transform 1 0 3496 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_38
timestamp 1649977179
transform 1 0 4600 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_50
timestamp 1649977179
transform 1 0 5704 0 -1 14144
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_21_57
timestamp 1649977179
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_69
timestamp 1649977179
transform 1 0 7452 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_81
timestamp 1649977179
transform 1 0 8556 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_93
timestamp 1649977179
transform 1 0 9660 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_105
timestamp 1649977179
transform 1 0 10764 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_111
timestamp 1649977179
transform 1 0 11316 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_113
timestamp 1649977179
transform 1 0 11500 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_125
timestamp 1649977179
transform 1 0 12604 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_21_135
timestamp 1649977179
transform 1 0 13524 0 -1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_21_141
timestamp 1649977179
transform 1 0 14076 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_153
timestamp 1649977179
transform 1 0 15180 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_21_165
timestamp 1649977179
transform 1 0 16284 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_21_169
timestamp 1649977179
transform 1 0 16652 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_175
timestamp 1649977179
transform 1 0 17204 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_178
timestamp 1649977179
transform 1 0 17480 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_190
timestamp 1649977179
transform 1 0 18584 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_202
timestamp 1649977179
transform 1 0 19688 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_214
timestamp 1649977179
transform 1 0 20792 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_222
timestamp 1649977179
transform 1 0 21528 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_21_225
timestamp 1649977179
transform 1 0 21804 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_237
timestamp 1649977179
transform 1 0 22908 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_249
timestamp 1649977179
transform 1 0 24012 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_261
timestamp 1649977179
transform 1 0 25116 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_273
timestamp 1649977179
transform 1 0 26220 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_279
timestamp 1649977179
transform 1 0 26772 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_281
timestamp 1649977179
transform 1 0 26956 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_293
timestamp 1649977179
transform 1 0 28060 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_305
timestamp 1649977179
transform 1 0 29164 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_317
timestamp 1649977179
transform 1 0 30268 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_329
timestamp 1649977179
transform 1 0 31372 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_335
timestamp 1649977179
transform 1 0 31924 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_337
timestamp 1649977179
transform 1 0 32108 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_349
timestamp 1649977179
transform 1 0 33212 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_361
timestamp 1649977179
transform 1 0 34316 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_373
timestamp 1649977179
transform 1 0 35420 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_385
timestamp 1649977179
transform 1 0 36524 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_391
timestamp 1649977179
transform 1 0 37076 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_393
timestamp 1649977179
transform 1 0 37260 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_405
timestamp 1649977179
transform 1 0 38364 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_417
timestamp 1649977179
transform 1 0 39468 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_429
timestamp 1649977179
transform 1 0 40572 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_441
timestamp 1649977179
transform 1 0 41676 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_447
timestamp 1649977179
transform 1 0 42228 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_449
timestamp 1649977179
transform 1 0 42412 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_461
timestamp 1649977179
transform 1 0 43516 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_473
timestamp 1649977179
transform 1 0 44620 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_485
timestamp 1649977179
transform 1 0 45724 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_497
timestamp 1649977179
transform 1 0 46828 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_503
timestamp 1649977179
transform 1 0 47380 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_505
timestamp 1649977179
transform 1 0 47564 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_517
timestamp 1649977179
transform 1 0 48668 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_529
timestamp 1649977179
transform 1 0 49772 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_541
timestamp 1649977179
transform 1 0 50876 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_553
timestamp 1649977179
transform 1 0 51980 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_559
timestamp 1649977179
transform 1 0 52532 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_561
timestamp 1649977179
transform 1 0 52716 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_573
timestamp 1649977179
transform 1 0 53820 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_585
timestamp 1649977179
transform 1 0 54924 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_597
timestamp 1649977179
transform 1 0 56028 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_609
timestamp 1649977179
transform 1 0 57132 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_615
timestamp 1649977179
transform 1 0 57684 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_617
timestamp 1649977179
transform 1 0 57868 0 -1 14144
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_22_3
timestamp 1649977179
transform 1 0 1380 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_15
timestamp 1649977179
transform 1 0 2484 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_27
timestamp 1649977179
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_29
timestamp 1649977179
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_41
timestamp 1649977179
transform 1 0 4876 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_53
timestamp 1649977179
transform 1 0 5980 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_65
timestamp 1649977179
transform 1 0 7084 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_77
timestamp 1649977179
transform 1 0 8188 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_83
timestamp 1649977179
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_85
timestamp 1649977179
transform 1 0 8924 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_97
timestamp 1649977179
transform 1 0 10028 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_109
timestamp 1649977179
transform 1 0 11132 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_121
timestamp 1649977179
transform 1 0 12236 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_133
timestamp 1649977179
transform 1 0 13340 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_139
timestamp 1649977179
transform 1 0 13892 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_141
timestamp 1649977179
transform 1 0 14076 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_153
timestamp 1649977179
transform 1 0 15180 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_165
timestamp 1649977179
transform 1 0 16284 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_177
timestamp 1649977179
transform 1 0 17388 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_189
timestamp 1649977179
transform 1 0 18492 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_195
timestamp 1649977179
transform 1 0 19044 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_197
timestamp 1649977179
transform 1 0 19228 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_209
timestamp 1649977179
transform 1 0 20332 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_221
timestamp 1649977179
transform 1 0 21436 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_233
timestamp 1649977179
transform 1 0 22540 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_245
timestamp 1649977179
transform 1 0 23644 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_251
timestamp 1649977179
transform 1 0 24196 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_253
timestamp 1649977179
transform 1 0 24380 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_265
timestamp 1649977179
transform 1 0 25484 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_277
timestamp 1649977179
transform 1 0 26588 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_289
timestamp 1649977179
transform 1 0 27692 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_301
timestamp 1649977179
transform 1 0 28796 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_307
timestamp 1649977179
transform 1 0 29348 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_309
timestamp 1649977179
transform 1 0 29532 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_321
timestamp 1649977179
transform 1 0 30636 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_333
timestamp 1649977179
transform 1 0 31740 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_345
timestamp 1649977179
transform 1 0 32844 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_357
timestamp 1649977179
transform 1 0 33948 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_363
timestamp 1649977179
transform 1 0 34500 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_365
timestamp 1649977179
transform 1 0 34684 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_377
timestamp 1649977179
transform 1 0 35788 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_389
timestamp 1649977179
transform 1 0 36892 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_401
timestamp 1649977179
transform 1 0 37996 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_413
timestamp 1649977179
transform 1 0 39100 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_419
timestamp 1649977179
transform 1 0 39652 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_421
timestamp 1649977179
transform 1 0 39836 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_433
timestamp 1649977179
transform 1 0 40940 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_445
timestamp 1649977179
transform 1 0 42044 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_457
timestamp 1649977179
transform 1 0 43148 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_469
timestamp 1649977179
transform 1 0 44252 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_475
timestamp 1649977179
transform 1 0 44804 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_477
timestamp 1649977179
transform 1 0 44988 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_489
timestamp 1649977179
transform 1 0 46092 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_501
timestamp 1649977179
transform 1 0 47196 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_513
timestamp 1649977179
transform 1 0 48300 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_525
timestamp 1649977179
transform 1 0 49404 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_531
timestamp 1649977179
transform 1 0 49956 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_533
timestamp 1649977179
transform 1 0 50140 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_545
timestamp 1649977179
transform 1 0 51244 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_557
timestamp 1649977179
transform 1 0 52348 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_569
timestamp 1649977179
transform 1 0 53452 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_581
timestamp 1649977179
transform 1 0 54556 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_587
timestamp 1649977179
transform 1 0 55108 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_589
timestamp 1649977179
transform 1 0 55292 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_601
timestamp 1649977179
transform 1 0 56396 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_613
timestamp 1649977179
transform 1 0 57500 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_3
timestamp 1649977179
transform 1 0 1380 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_15
timestamp 1649977179
transform 1 0 2484 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_27
timestamp 1649977179
transform 1 0 3588 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_39
timestamp 1649977179
transform 1 0 4692 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_51
timestamp 1649977179
transform 1 0 5796 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_55
timestamp 1649977179
transform 1 0 6164 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_57
timestamp 1649977179
transform 1 0 6348 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_69
timestamp 1649977179
transform 1 0 7452 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_81
timestamp 1649977179
transform 1 0 8556 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_93
timestamp 1649977179
transform 1 0 9660 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_105
timestamp 1649977179
transform 1 0 10764 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_111
timestamp 1649977179
transform 1 0 11316 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_113
timestamp 1649977179
transform 1 0 11500 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_125
timestamp 1649977179
transform 1 0 12604 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_137
timestamp 1649977179
transform 1 0 13708 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_149
timestamp 1649977179
transform 1 0 14812 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_161
timestamp 1649977179
transform 1 0 15916 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_167
timestamp 1649977179
transform 1 0 16468 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_169
timestamp 1649977179
transform 1 0 16652 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_181
timestamp 1649977179
transform 1 0 17756 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_193
timestamp 1649977179
transform 1 0 18860 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_205
timestamp 1649977179
transform 1 0 19964 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_217
timestamp 1649977179
transform 1 0 21068 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_223
timestamp 1649977179
transform 1 0 21620 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_225
timestamp 1649977179
transform 1 0 21804 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_237
timestamp 1649977179
transform 1 0 22908 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_249
timestamp 1649977179
transform 1 0 24012 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_261
timestamp 1649977179
transform 1 0 25116 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_273
timestamp 1649977179
transform 1 0 26220 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_279
timestamp 1649977179
transform 1 0 26772 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_281
timestamp 1649977179
transform 1 0 26956 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_293
timestamp 1649977179
transform 1 0 28060 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_305
timestamp 1649977179
transform 1 0 29164 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_317
timestamp 1649977179
transform 1 0 30268 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_329
timestamp 1649977179
transform 1 0 31372 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_335
timestamp 1649977179
transform 1 0 31924 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_337
timestamp 1649977179
transform 1 0 32108 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_349
timestamp 1649977179
transform 1 0 33212 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_361
timestamp 1649977179
transform 1 0 34316 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_373
timestamp 1649977179
transform 1 0 35420 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_385
timestamp 1649977179
transform 1 0 36524 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_391
timestamp 1649977179
transform 1 0 37076 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_393
timestamp 1649977179
transform 1 0 37260 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_405
timestamp 1649977179
transform 1 0 38364 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_417
timestamp 1649977179
transform 1 0 39468 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_429
timestamp 1649977179
transform 1 0 40572 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_441
timestamp 1649977179
transform 1 0 41676 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_447
timestamp 1649977179
transform 1 0 42228 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_449
timestamp 1649977179
transform 1 0 42412 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_461
timestamp 1649977179
transform 1 0 43516 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_473
timestamp 1649977179
transform 1 0 44620 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_485
timestamp 1649977179
transform 1 0 45724 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_497
timestamp 1649977179
transform 1 0 46828 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_503
timestamp 1649977179
transform 1 0 47380 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_505
timestamp 1649977179
transform 1 0 47564 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_517
timestamp 1649977179
transform 1 0 48668 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_529
timestamp 1649977179
transform 1 0 49772 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_541
timestamp 1649977179
transform 1 0 50876 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_553
timestamp 1649977179
transform 1 0 51980 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_559
timestamp 1649977179
transform 1 0 52532 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_561
timestamp 1649977179
transform 1 0 52716 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_573
timestamp 1649977179
transform 1 0 53820 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_585
timestamp 1649977179
transform 1 0 54924 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_597
timestamp 1649977179
transform 1 0 56028 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_609
timestamp 1649977179
transform 1 0 57132 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_615
timestamp 1649977179
transform 1 0 57684 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_617
timestamp 1649977179
transform 1 0 57868 0 -1 15232
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_24_3
timestamp 1649977179
transform 1 0 1380 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_15
timestamp 1649977179
transform 1 0 2484 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_27
timestamp 1649977179
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_29
timestamp 1649977179
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_41
timestamp 1649977179
transform 1 0 4876 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_53
timestamp 1649977179
transform 1 0 5980 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_65
timestamp 1649977179
transform 1 0 7084 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_77
timestamp 1649977179
transform 1 0 8188 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_83
timestamp 1649977179
transform 1 0 8740 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_85
timestamp 1649977179
transform 1 0 8924 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_97
timestamp 1649977179
transform 1 0 10028 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_109
timestamp 1649977179
transform 1 0 11132 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_121
timestamp 1649977179
transform 1 0 12236 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_133
timestamp 1649977179
transform 1 0 13340 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_139
timestamp 1649977179
transform 1 0 13892 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_141
timestamp 1649977179
transform 1 0 14076 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_153
timestamp 1649977179
transform 1 0 15180 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_165
timestamp 1649977179
transform 1 0 16284 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_177
timestamp 1649977179
transform 1 0 17388 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_189
timestamp 1649977179
transform 1 0 18492 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_195
timestamp 1649977179
transform 1 0 19044 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_197
timestamp 1649977179
transform 1 0 19228 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_209
timestamp 1649977179
transform 1 0 20332 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_221
timestamp 1649977179
transform 1 0 21436 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_233
timestamp 1649977179
transform 1 0 22540 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_245
timestamp 1649977179
transform 1 0 23644 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_251
timestamp 1649977179
transform 1 0 24196 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_253
timestamp 1649977179
transform 1 0 24380 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_265
timestamp 1649977179
transform 1 0 25484 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_277
timestamp 1649977179
transform 1 0 26588 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_289
timestamp 1649977179
transform 1 0 27692 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_301
timestamp 1649977179
transform 1 0 28796 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_307
timestamp 1649977179
transform 1 0 29348 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_309
timestamp 1649977179
transform 1 0 29532 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_321
timestamp 1649977179
transform 1 0 30636 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_333
timestamp 1649977179
transform 1 0 31740 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_345
timestamp 1649977179
transform 1 0 32844 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_357
timestamp 1649977179
transform 1 0 33948 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_363
timestamp 1649977179
transform 1 0 34500 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_365
timestamp 1649977179
transform 1 0 34684 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_377
timestamp 1649977179
transform 1 0 35788 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_389
timestamp 1649977179
transform 1 0 36892 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_401
timestamp 1649977179
transform 1 0 37996 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_413
timestamp 1649977179
transform 1 0 39100 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_419
timestamp 1649977179
transform 1 0 39652 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_421
timestamp 1649977179
transform 1 0 39836 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_433
timestamp 1649977179
transform 1 0 40940 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_445
timestamp 1649977179
transform 1 0 42044 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_457
timestamp 1649977179
transform 1 0 43148 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_469
timestamp 1649977179
transform 1 0 44252 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_475
timestamp 1649977179
transform 1 0 44804 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_477
timestamp 1649977179
transform 1 0 44988 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_489
timestamp 1649977179
transform 1 0 46092 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_501
timestamp 1649977179
transform 1 0 47196 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_513
timestamp 1649977179
transform 1 0 48300 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_525
timestamp 1649977179
transform 1 0 49404 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_531
timestamp 1649977179
transform 1 0 49956 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_533
timestamp 1649977179
transform 1 0 50140 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_545
timestamp 1649977179
transform 1 0 51244 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_557
timestamp 1649977179
transform 1 0 52348 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_569
timestamp 1649977179
transform 1 0 53452 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_581
timestamp 1649977179
transform 1 0 54556 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_587
timestamp 1649977179
transform 1 0 55108 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_589
timestamp 1649977179
transform 1 0 55292 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_601
timestamp 1649977179
transform 1 0 56396 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_613
timestamp 1649977179
transform 1 0 57500 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_3
timestamp 1649977179
transform 1 0 1380 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_15
timestamp 1649977179
transform 1 0 2484 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_27
timestamp 1649977179
transform 1 0 3588 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_39
timestamp 1649977179
transform 1 0 4692 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_51
timestamp 1649977179
transform 1 0 5796 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_55
timestamp 1649977179
transform 1 0 6164 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_57
timestamp 1649977179
transform 1 0 6348 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_69
timestamp 1649977179
transform 1 0 7452 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_81
timestamp 1649977179
transform 1 0 8556 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_93
timestamp 1649977179
transform 1 0 9660 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_105
timestamp 1649977179
transform 1 0 10764 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_111
timestamp 1649977179
transform 1 0 11316 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_113
timestamp 1649977179
transform 1 0 11500 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_125
timestamp 1649977179
transform 1 0 12604 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_137
timestamp 1649977179
transform 1 0 13708 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_149
timestamp 1649977179
transform 1 0 14812 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_161
timestamp 1649977179
transform 1 0 15916 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_167
timestamp 1649977179
transform 1 0 16468 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_169
timestamp 1649977179
transform 1 0 16652 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_181
timestamp 1649977179
transform 1 0 17756 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_193
timestamp 1649977179
transform 1 0 18860 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_205
timestamp 1649977179
transform 1 0 19964 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_217
timestamp 1649977179
transform 1 0 21068 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_223
timestamp 1649977179
transform 1 0 21620 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_225
timestamp 1649977179
transform 1 0 21804 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_237
timestamp 1649977179
transform 1 0 22908 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_249
timestamp 1649977179
transform 1 0 24012 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_261
timestamp 1649977179
transform 1 0 25116 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_273
timestamp 1649977179
transform 1 0 26220 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_279
timestamp 1649977179
transform 1 0 26772 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_281
timestamp 1649977179
transform 1 0 26956 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_293
timestamp 1649977179
transform 1 0 28060 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_305
timestamp 1649977179
transform 1 0 29164 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_317
timestamp 1649977179
transform 1 0 30268 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_329
timestamp 1649977179
transform 1 0 31372 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_335
timestamp 1649977179
transform 1 0 31924 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_337
timestamp 1649977179
transform 1 0 32108 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_349
timestamp 1649977179
transform 1 0 33212 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_361
timestamp 1649977179
transform 1 0 34316 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_373
timestamp 1649977179
transform 1 0 35420 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_385
timestamp 1649977179
transform 1 0 36524 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_391
timestamp 1649977179
transform 1 0 37076 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_393
timestamp 1649977179
transform 1 0 37260 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_405
timestamp 1649977179
transform 1 0 38364 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_417
timestamp 1649977179
transform 1 0 39468 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_429
timestamp 1649977179
transform 1 0 40572 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_441
timestamp 1649977179
transform 1 0 41676 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_447
timestamp 1649977179
transform 1 0 42228 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_449
timestamp 1649977179
transform 1 0 42412 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_461
timestamp 1649977179
transform 1 0 43516 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_473
timestamp 1649977179
transform 1 0 44620 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_485
timestamp 1649977179
transform 1 0 45724 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_497
timestamp 1649977179
transform 1 0 46828 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_503
timestamp 1649977179
transform 1 0 47380 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_505
timestamp 1649977179
transform 1 0 47564 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_517
timestamp 1649977179
transform 1 0 48668 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_529
timestamp 1649977179
transform 1 0 49772 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_541
timestamp 1649977179
transform 1 0 50876 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_553
timestamp 1649977179
transform 1 0 51980 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_559
timestamp 1649977179
transform 1 0 52532 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_561
timestamp 1649977179
transform 1 0 52716 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_573
timestamp 1649977179
transform 1 0 53820 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_585
timestamp 1649977179
transform 1 0 54924 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_597
timestamp 1649977179
transform 1 0 56028 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_609
timestamp 1649977179
transform 1 0 57132 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_615
timestamp 1649977179
transform 1 0 57684 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_617
timestamp 1649977179
transform 1 0 57868 0 -1 16320
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_26_3
timestamp 1649977179
transform 1 0 1380 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_15
timestamp 1649977179
transform 1 0 2484 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_27
timestamp 1649977179
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_29
timestamp 1649977179
transform 1 0 3772 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_41
timestamp 1649977179
transform 1 0 4876 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_53
timestamp 1649977179
transform 1 0 5980 0 1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_26_60
timestamp 1649977179
transform 1 0 6624 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_72
timestamp 1649977179
transform 1 0 7728 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_85
timestamp 1649977179
transform 1 0 8924 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_97
timestamp 1649977179
transform 1 0 10028 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_26_109
timestamp 1649977179
transform 1 0 11132 0 1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_26_115
timestamp 1649977179
transform 1 0 11684 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_127
timestamp 1649977179
transform 1 0 12788 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_139
timestamp 1649977179
transform 1 0 13892 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_26_141
timestamp 1649977179
transform 1 0 14076 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_145
timestamp 1649977179
transform 1 0 14444 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_157
timestamp 1649977179
transform 1 0 15548 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_26_169
timestamp 1649977179
transform 1 0 16652 0 1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_26_175
timestamp 1649977179
transform 1 0 17204 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_187
timestamp 1649977179
transform 1 0 18308 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_195
timestamp 1649977179
transform 1 0 19044 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_197
timestamp 1649977179
transform 1 0 19228 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_209
timestamp 1649977179
transform 1 0 20332 0 1 16320
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_26_220
timestamp 1649977179
transform 1 0 21344 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_232
timestamp 1649977179
transform 1 0 22448 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_244
timestamp 1649977179
transform 1 0 23552 0 1 16320
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_26_256
timestamp 1649977179
transform 1 0 24656 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_268
timestamp 1649977179
transform 1 0 25760 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_26_280
timestamp 1649977179
transform 1 0 26864 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_26_285
timestamp 1649977179
transform 1 0 27324 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_297
timestamp 1649977179
transform 1 0 28428 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_26_305
timestamp 1649977179
transform 1 0 29164 0 1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_26_309
timestamp 1649977179
transform 1 0 29532 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_321
timestamp 1649977179
transform 1 0 30636 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_333
timestamp 1649977179
transform 1 0 31740 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_345
timestamp 1649977179
transform 1 0 32844 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_357
timestamp 1649977179
transform 1 0 33948 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_363
timestamp 1649977179
transform 1 0 34500 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_365
timestamp 1649977179
transform 1 0 34684 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_377
timestamp 1649977179
transform 1 0 35788 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_381
timestamp 1649977179
transform 1 0 36156 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_385
timestamp 1649977179
transform 1 0 36524 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_397
timestamp 1649977179
transform 1 0 37628 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_409
timestamp 1649977179
transform 1 0 38732 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_26_417
timestamp 1649977179
transform 1 0 39468 0 1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_26_424
timestamp 1649977179
transform 1 0 40112 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_436
timestamp 1649977179
transform 1 0 41216 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_448
timestamp 1649977179
transform 1 0 42320 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_26_460
timestamp 1649977179
transform 1 0 43424 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_26_465
timestamp 1649977179
transform 1 0 43884 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_26_473
timestamp 1649977179
transform 1 0 44620 0 1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_26_477
timestamp 1649977179
transform 1 0 44988 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_26_489
timestamp 1649977179
transform 1 0 46092 0 1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_26_495
timestamp 1649977179
transform 1 0 46644 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_507
timestamp 1649977179
transform 1 0 47748 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_26_519
timestamp 1649977179
transform 1 0 48852 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_26_525
timestamp 1649977179
transform 1 0 49404 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_531
timestamp 1649977179
transform 1 0 49956 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_533
timestamp 1649977179
transform 1 0 50140 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_545
timestamp 1649977179
transform 1 0 51244 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_557
timestamp 1649977179
transform 1 0 52348 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_569
timestamp 1649977179
transform 1 0 53452 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_26_580
timestamp 1649977179
transform 1 0 54464 0 1 16320
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_26_589
timestamp 1649977179
transform 1 0 55292 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_601
timestamp 1649977179
transform 1 0 56396 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_613
timestamp 1649977179
transform 1 0 57500 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_3
timestamp 1649977179
transform 1 0 1380 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_15
timestamp 1649977179
transform 1 0 2484 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_27_27
timestamp 1649977179
transform 1 0 3588 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_27_29
timestamp 1649977179
transform 1 0 3772 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_27_38
timestamp 1649977179
transform 1 0 4600 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_45
timestamp 1649977179
transform 1 0 5244 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_52
timestamp 1649977179
transform 1 0 5888 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_27_57
timestamp 1649977179
transform 1 0 6348 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_27_66
timestamp 1649977179
transform 1 0 7176 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_73
timestamp 1649977179
transform 1 0 7820 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_80
timestamp 1649977179
transform 1 0 8464 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_85
timestamp 1649977179
transform 1 0 8924 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_90
timestamp 1649977179
transform 1 0 9384 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_94
timestamp 1649977179
transform 1 0 9752 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_98
timestamp 1649977179
transform 1 0 10120 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_27_105
timestamp 1649977179
transform 1 0 10764 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_111
timestamp 1649977179
transform 1 0 11316 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_113
timestamp 1649977179
transform 1 0 11500 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_120
timestamp 1649977179
transform 1 0 12144 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_124
timestamp 1649977179
transform 1 0 12512 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_128
timestamp 1649977179
transform 1 0 12880 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_135
timestamp 1649977179
transform 1 0 13524 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_139
timestamp 1649977179
transform 1 0 13892 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_27_141
timestamp 1649977179
transform 1 0 14076 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_27_150
timestamp 1649977179
transform 1 0 14904 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_157
timestamp 1649977179
transform 1 0 15548 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_164
timestamp 1649977179
transform 1 0 16192 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_27_169
timestamp 1649977179
transform 1 0 16652 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_27_178
timestamp 1649977179
transform 1 0 17480 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_185
timestamp 1649977179
transform 1 0 18124 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_192
timestamp 1649977179
transform 1 0 18768 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_27_197
timestamp 1649977179
transform 1 0 19228 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_27_203
timestamp 1649977179
transform 1 0 19780 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_27_210
timestamp 1649977179
transform 1 0 20424 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_216
timestamp 1649977179
transform 1 0 20976 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_220
timestamp 1649977179
transform 1 0 21344 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_225
timestamp 1649977179
transform 1 0 21804 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_229
timestamp 1649977179
transform 1 0 22172 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_233
timestamp 1649977179
transform 1 0 22540 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_240
timestamp 1649977179
transform 1 0 23184 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_244
timestamp 1649977179
transform 1 0 23552 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_248
timestamp 1649977179
transform 1 0 23920 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_27_253
timestamp 1649977179
transform 1 0 24380 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_27_262
timestamp 1649977179
transform 1 0 25208 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_269
timestamp 1649977179
transform 1 0 25852 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_276
timestamp 1649977179
transform 1 0 26496 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_27_281
timestamp 1649977179
transform 1 0 26956 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_27_290
timestamp 1649977179
transform 1 0 27784 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_297
timestamp 1649977179
transform 1 0 28428 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_304
timestamp 1649977179
transform 1 0 29072 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_27_309
timestamp 1649977179
transform 1 0 29532 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_27_315
timestamp 1649977179
transform 1 0 30084 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_319
timestamp 1649977179
transform 1 0 30452 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_323
timestamp 1649977179
transform 1 0 30820 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_27_330
timestamp 1649977179
transform 1 0 31464 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_27_340
timestamp 1649977179
transform 1 0 32384 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_347
timestamp 1649977179
transform 1 0 33028 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_351
timestamp 1649977179
transform 1 0 33396 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_355
timestamp 1649977179
transform 1 0 33764 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_363
timestamp 1649977179
transform 1 0 34500 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_368
timestamp 1649977179
transform 1 0 34960 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_375
timestamp 1649977179
transform 1 0 35604 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_27_382
timestamp 1649977179
transform 1 0 36248 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_390
timestamp 1649977179
transform 1 0 36984 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_396
timestamp 1649977179
transform 1 0 37536 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_403
timestamp 1649977179
transform 1 0 38180 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_27_410
timestamp 1649977179
transform 1 0 38824 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_418
timestamp 1649977179
transform 1 0 39560 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_424
timestamp 1649977179
transform 1 0 40112 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_431
timestamp 1649977179
transform 1 0 40756 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_27_438
timestamp 1649977179
transform 1 0 41400 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_446
timestamp 1649977179
transform 1 0 42136 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_452
timestamp 1649977179
transform 1 0 42688 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_459
timestamp 1649977179
transform 1 0 43332 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_27_466
timestamp 1649977179
transform 1 0 43976 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_474
timestamp 1649977179
transform 1 0 44712 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_480
timestamp 1649977179
transform 1 0 45264 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_487
timestamp 1649977179
transform 1 0 45908 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_27_494
timestamp 1649977179
transform 1 0 46552 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_502
timestamp 1649977179
transform 1 0 47288 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_508
timestamp 1649977179
transform 1 0 47840 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_515
timestamp 1649977179
transform 1 0 48484 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_27_522
timestamp 1649977179
transform 1 0 49128 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_530
timestamp 1649977179
transform 1 0 49864 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_536
timestamp 1649977179
transform 1 0 50416 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_543
timestamp 1649977179
transform 1 0 51060 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_27_550
timestamp 1649977179
transform 1 0 51704 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_558
timestamp 1649977179
transform 1 0 52440 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_564
timestamp 1649977179
transform 1 0 52992 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_571
timestamp 1649977179
transform 1 0 53636 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_27_578
timestamp 1649977179
transform 1 0 54280 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_586
timestamp 1649977179
transform 1 0 55016 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_592
timestamp 1649977179
transform 1 0 55568 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_599
timestamp 1649977179
transform 1 0 56212 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_27_606
timestamp 1649977179
transform 1 0 56856 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_614
timestamp 1649977179
transform 1 0 57592 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_27_617
timestamp 1649977179
transform 1 0 57868 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1649977179
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1649977179
transform -1 0 58880 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1649977179
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1649977179
transform -1 0 58880 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1649977179
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1649977179
transform -1 0 58880 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1649977179
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1649977179
transform -1 0 58880 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1649977179
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1649977179
transform -1 0 58880 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1649977179
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1649977179
transform -1 0 58880 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1649977179
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1649977179
transform -1 0 58880 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1649977179
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1649977179
transform -1 0 58880 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1649977179
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1649977179
transform -1 0 58880 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1649977179
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1649977179
transform -1 0 58880 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1649977179
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1649977179
transform -1 0 58880 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1649977179
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1649977179
transform -1 0 58880 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1649977179
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1649977179
transform -1 0 58880 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1649977179
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1649977179
transform -1 0 58880 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1649977179
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1649977179
transform -1 0 58880 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1649977179
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1649977179
transform -1 0 58880 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1649977179
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1649977179
transform -1 0 58880 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1649977179
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1649977179
transform -1 0 58880 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1649977179
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1649977179
transform -1 0 58880 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1649977179
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1649977179
transform -1 0 58880 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1649977179
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1649977179
transform -1 0 58880 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1649977179
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1649977179
transform -1 0 58880 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1649977179
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1649977179
transform -1 0 58880 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1649977179
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1649977179
transform -1 0 58880 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1649977179
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1649977179
transform -1 0 58880 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1649977179
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1649977179
transform -1 0 58880 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1649977179
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1649977179
transform -1 0 58880 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1649977179
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1649977179
transform -1 0 58880 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_56 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_57
timestamp 1649977179
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_58
timestamp 1649977179
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_59
timestamp 1649977179
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_60
timestamp 1649977179
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_61
timestamp 1649977179
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_62
timestamp 1649977179
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_63
timestamp 1649977179
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_64
timestamp 1649977179
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_65
timestamp 1649977179
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_66
timestamp 1649977179
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_67
timestamp 1649977179
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_68
timestamp 1649977179
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_69
timestamp 1649977179
transform 1 0 37168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_70
timestamp 1649977179
transform 1 0 39744 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_71
timestamp 1649977179
transform 1 0 42320 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_72
timestamp 1649977179
transform 1 0 44896 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_73
timestamp 1649977179
transform 1 0 47472 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_74
timestamp 1649977179
transform 1 0 50048 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_75
timestamp 1649977179
transform 1 0 52624 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_76
timestamp 1649977179
transform 1 0 55200 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_77
timestamp 1649977179
transform 1 0 57776 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_78
timestamp 1649977179
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_79
timestamp 1649977179
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_80
timestamp 1649977179
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_81
timestamp 1649977179
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_82
timestamp 1649977179
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_83
timestamp 1649977179
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_84
timestamp 1649977179
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_85
timestamp 1649977179
transform 1 0 42320 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_86
timestamp 1649977179
transform 1 0 47472 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_87
timestamp 1649977179
transform 1 0 52624 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_88
timestamp 1649977179
transform 1 0 57776 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_89
timestamp 1649977179
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_90
timestamp 1649977179
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_91
timestamp 1649977179
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_92
timestamp 1649977179
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_93
timestamp 1649977179
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_94
timestamp 1649977179
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_95
timestamp 1649977179
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_96
timestamp 1649977179
transform 1 0 39744 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_97
timestamp 1649977179
transform 1 0 44896 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_98
timestamp 1649977179
transform 1 0 50048 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_99
timestamp 1649977179
transform 1 0 55200 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_100
timestamp 1649977179
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_101
timestamp 1649977179
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_102
timestamp 1649977179
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_103
timestamp 1649977179
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_104
timestamp 1649977179
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_105
timestamp 1649977179
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_106
timestamp 1649977179
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_107
timestamp 1649977179
transform 1 0 42320 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_108
timestamp 1649977179
transform 1 0 47472 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_109
timestamp 1649977179
transform 1 0 52624 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_110
timestamp 1649977179
transform 1 0 57776 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_111
timestamp 1649977179
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_112
timestamp 1649977179
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_113
timestamp 1649977179
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_114
timestamp 1649977179
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_115
timestamp 1649977179
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_116
timestamp 1649977179
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_117
timestamp 1649977179
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_118
timestamp 1649977179
transform 1 0 39744 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_119
timestamp 1649977179
transform 1 0 44896 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_120
timestamp 1649977179
transform 1 0 50048 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_121
timestamp 1649977179
transform 1 0 55200 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_122
timestamp 1649977179
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_123
timestamp 1649977179
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_124
timestamp 1649977179
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_125
timestamp 1649977179
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_126
timestamp 1649977179
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_127
timestamp 1649977179
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_128
timestamp 1649977179
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_129
timestamp 1649977179
transform 1 0 42320 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130
timestamp 1649977179
transform 1 0 47472 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 1649977179
transform 1 0 52624 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 1649977179
transform 1 0 57776 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 1649977179
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 1649977179
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1649977179
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1649977179
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1649977179
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1649977179
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1649977179
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1649977179
transform 1 0 39744 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1649977179
transform 1 0 44896 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1649977179
transform 1 0 50048 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1649977179
transform 1 0 55200 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1649977179
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1649977179
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1649977179
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1649977179
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1649977179
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1649977179
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1649977179
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1649977179
transform 1 0 42320 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1649977179
transform 1 0 47472 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1649977179
transform 1 0 52624 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1649977179
transform 1 0 57776 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1649977179
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1649977179
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1649977179
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1649977179
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1649977179
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1649977179
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1649977179
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1649977179
transform 1 0 39744 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1649977179
transform 1 0 44896 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1649977179
transform 1 0 50048 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1649977179
transform 1 0 55200 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1649977179
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1649977179
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1649977179
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1649977179
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1649977179
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1649977179
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1649977179
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1649977179
transform 1 0 42320 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1649977179
transform 1 0 47472 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1649977179
transform 1 0 52624 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1649977179
transform 1 0 57776 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1649977179
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1649977179
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1649977179
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1649977179
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1649977179
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1649977179
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1649977179
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1649977179
transform 1 0 39744 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1649977179
transform 1 0 44896 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1649977179
transform 1 0 50048 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1649977179
transform 1 0 55200 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1649977179
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1649977179
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1649977179
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1649977179
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1649977179
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1649977179
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1649977179
transform 1 0 37168 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1649977179
transform 1 0 42320 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1649977179
transform 1 0 47472 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1649977179
transform 1 0 52624 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1649977179
transform 1 0 57776 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1649977179
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1649977179
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1649977179
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1649977179
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1649977179
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1649977179
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1649977179
transform 1 0 34592 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1649977179
transform 1 0 39744 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1649977179
transform 1 0 44896 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1649977179
transform 1 0 50048 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1649977179
transform 1 0 55200 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1649977179
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1649977179
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1649977179
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1649977179
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1649977179
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1649977179
transform 1 0 32016 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1649977179
transform 1 0 37168 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1649977179
transform 1 0 42320 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1649977179
transform 1 0 47472 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1649977179
transform 1 0 52624 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1649977179
transform 1 0 57776 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1649977179
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1649977179
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1649977179
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1649977179
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1649977179
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1649977179
transform 1 0 29440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1649977179
transform 1 0 34592 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1649977179
transform 1 0 39744 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1649977179
transform 1 0 44896 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1649977179
transform 1 0 50048 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1649977179
transform 1 0 55200 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1649977179
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1649977179
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1649977179
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1649977179
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1649977179
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1649977179
transform 1 0 32016 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1649977179
transform 1 0 37168 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1649977179
transform 1 0 42320 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1649977179
transform 1 0 47472 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1649977179
transform 1 0 52624 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1649977179
transform 1 0 57776 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1649977179
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1649977179
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1649977179
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1649977179
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1649977179
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1649977179
transform 1 0 29440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1649977179
transform 1 0 34592 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1649977179
transform 1 0 39744 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1649977179
transform 1 0 44896 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1649977179
transform 1 0 50048 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1649977179
transform 1 0 55200 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1649977179
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1649977179
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1649977179
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1649977179
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1649977179
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1649977179
transform 1 0 32016 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1649977179
transform 1 0 37168 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1649977179
transform 1 0 42320 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1649977179
transform 1 0 47472 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1649977179
transform 1 0 52624 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1649977179
transform 1 0 57776 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1649977179
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1649977179
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1649977179
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1649977179
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1649977179
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1649977179
transform 1 0 29440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1649977179
transform 1 0 34592 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1649977179
transform 1 0 39744 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1649977179
transform 1 0 44896 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1649977179
transform 1 0 50048 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1649977179
transform 1 0 55200 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1649977179
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1649977179
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1649977179
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1649977179
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1649977179
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1649977179
transform 1 0 32016 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1649977179
transform 1 0 37168 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1649977179
transform 1 0 42320 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1649977179
transform 1 0 47472 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1649977179
transform 1 0 52624 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1649977179
transform 1 0 57776 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1649977179
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1649977179
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1649977179
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1649977179
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1649977179
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1649977179
transform 1 0 29440 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1649977179
transform 1 0 34592 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1649977179
transform 1 0 39744 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1649977179
transform 1 0 44896 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1649977179
transform 1 0 50048 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1649977179
transform 1 0 55200 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1649977179
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1649977179
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1649977179
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1649977179
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1649977179
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1649977179
transform 1 0 32016 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1649977179
transform 1 0 37168 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1649977179
transform 1 0 42320 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1649977179
transform 1 0 47472 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1649977179
transform 1 0 52624 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1649977179
transform 1 0 57776 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1649977179
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1649977179
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1649977179
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1649977179
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1649977179
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1649977179
transform 1 0 29440 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1649977179
transform 1 0 34592 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1649977179
transform 1 0 39744 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1649977179
transform 1 0 44896 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1649977179
transform 1 0 50048 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1649977179
transform 1 0 55200 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1649977179
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1649977179
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1649977179
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1649977179
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1649977179
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1649977179
transform 1 0 32016 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1649977179
transform 1 0 37168 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1649977179
transform 1 0 42320 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1649977179
transform 1 0 47472 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1649977179
transform 1 0 52624 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1649977179
transform 1 0 57776 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1649977179
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1649977179
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1649977179
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1649977179
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1649977179
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1649977179
transform 1 0 29440 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1649977179
transform 1 0 34592 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1649977179
transform 1 0 39744 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1649977179
transform 1 0 44896 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1649977179
transform 1 0 50048 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1649977179
transform 1 0 55200 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1649977179
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1649977179
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1649977179
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1649977179
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1649977179
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1649977179
transform 1 0 32016 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1649977179
transform 1 0 37168 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1649977179
transform 1 0 42320 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1649977179
transform 1 0 47472 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1649977179
transform 1 0 52624 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1649977179
transform 1 0 57776 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1649977179
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1649977179
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1649977179
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1649977179
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1649977179
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1649977179
transform 1 0 29440 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1649977179
transform 1 0 34592 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1649977179
transform 1 0 39744 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1649977179
transform 1 0 44896 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1649977179
transform 1 0 50048 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1649977179
transform 1 0 55200 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1649977179
transform 1 0 3680 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1649977179
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1649977179
transform 1 0 8832 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1649977179
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1649977179
transform 1 0 13984 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1649977179
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1649977179
transform 1 0 19136 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1649977179
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1649977179
transform 1 0 24288 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1649977179
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1649977179
transform 1 0 29440 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1649977179
transform 1 0 32016 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1649977179
transform 1 0 34592 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1649977179
transform 1 0 37168 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1649977179
transform 1 0 39744 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1649977179
transform 1 0 42320 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1649977179
transform 1 0 44896 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1649977179
transform 1 0 47472 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1649977179
transform 1 0 50048 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1649977179
transform 1 0 52624 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1649977179
transform 1 0 55200 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1649977179
transform 1 0 57776 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  _0398_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 33396 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0399_
timestamp 1649977179
transform 1 0 42320 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _0400_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 23644 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0401_
timestamp 1649977179
transform 1 0 27416 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0402_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 29072 0 1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__nand2_2  _0403_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 30452 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0404_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 15364 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0405_
timestamp 1649977179
transform 1 0 12328 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _0406_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 30360 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _0407_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 32936 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__a211oi_1  _0408_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 32108 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _0409_
timestamp 1649977179
transform -1 0 41676 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _0410_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 41308 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _0411_
timestamp 1649977179
transform 1 0 29900 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _0412_
timestamp 1649977179
transform 1 0 35236 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__nor3_1  _0413_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 37444 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _0414_
timestamp 1649977179
transform 1 0 34684 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _0415_
timestamp 1649977179
transform -1 0 34868 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__or3b_2  _0416_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 35788 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0417_
timestamp 1649977179
transform -1 0 18768 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0418_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 34592 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__nand2b_2  _0419_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 32568 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__or2b_1  _0420_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 30084 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _0421_
timestamp 1649977179
transform -1 0 31096 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _0422_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 26588 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0423_
timestamp 1649977179
transform -1 0 34224 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _0424_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 35236 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _0425_
timestamp 1649977179
transform 1 0 37076 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__or2b_2  _0426_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 28980 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_2  _0427_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 27508 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0428_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 42872 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0429_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 43884 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__nand2b_2  _0430_
timestamp 1649977179
transform -1 0 29164 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_2  _0431_
timestamp 1649977179
transform -1 0 28704 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0432_
timestamp 1649977179
transform -1 0 46276 0 -1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__or2_1  _0433_
timestamp 1649977179
transform -1 0 25392 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _0434_
timestamp 1649977179
transform -1 0 26220 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0435_
timestamp 1649977179
transform -1 0 13616 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__a31oi_4  _0436_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 26496 0 -1 7616
box -38 -48 1602 592
use sky130_fd_sc_hd__nor2_1  _0437_
timestamp 1649977179
transform 1 0 24288 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0438_
timestamp 1649977179
transform -1 0 28244 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0439_
timestamp 1649977179
transform -1 0 25944 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0440_
timestamp 1649977179
transform -1 0 25116 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _0441_
timestamp 1649977179
transform 1 0 29072 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0442_
timestamp 1649977179
transform -1 0 31464 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0443_
timestamp 1649977179
transform -1 0 10396 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0444_
timestamp 1649977179
transform -1 0 8280 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0445_
timestamp 1649977179
transform -1 0 5888 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0446_
timestamp 1649977179
transform -1 0 24564 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0447_
timestamp 1649977179
transform 1 0 26772 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0448_
timestamp 1649977179
transform -1 0 44896 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _0449_
timestamp 1649977179
transform -1 0 25300 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0450_
timestamp 1649977179
transform 1 0 21160 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0451_
timestamp 1649977179
transform 1 0 34684 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0452_
timestamp 1649977179
transform 1 0 34868 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0453_
timestamp 1649977179
transform -1 0 55476 0 -1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__inv_2  _0454_
timestamp 1649977179
transform 1 0 54096 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0455_
timestamp 1649977179
transform 1 0 55292 0 1 5440
box -38 -48 958 592
use sky130_fd_sc_hd__nor2_1  _0456_
timestamp 1649977179
transform -1 0 56028 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0457_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 55384 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _0458_
timestamp 1649977179
transform -1 0 54740 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _0459_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 52716 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0460_
timestamp 1649977179
transform 1 0 56764 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _0461_
timestamp 1649977179
transform 1 0 55936 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0462_
timestamp 1649977179
transform -1 0 57960 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0463_
timestamp 1649977179
transform 1 0 57868 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0464_
timestamp 1649977179
transform 1 0 56304 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0465_
timestamp 1649977179
transform 1 0 57868 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0466_
timestamp 1649977179
transform 1 0 55660 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0467_
timestamp 1649977179
transform 1 0 57868 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__or4_2  _0468_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 16744 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _0469_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 40572 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__nor4_4  _0470_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 37444 0 1 3264
box -38 -48 1602 592
use sky130_fd_sc_hd__or4_1  _0471_
timestamp 1649977179
transform 1 0 28428 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0472_
timestamp 1649977179
transform -1 0 45540 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__or4_2  _0473_
timestamp 1649977179
transform -1 0 40480 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0474_
timestamp 1649977179
transform -1 0 52164 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _0475_
timestamp 1649977179
transform -1 0 53544 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0476_
timestamp 1649977179
transform -1 0 54832 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _0477_
timestamp 1649977179
transform -1 0 56396 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0478_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 55384 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__a21boi_1  _0479_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 54556 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _0480_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 53820 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__o2bb2a_1  _0481_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 52716 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _0482_
timestamp 1649977179
transform -1 0 52256 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _0483_
timestamp 1649977179
transform 1 0 55292 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0484_
timestamp 1649977179
transform 1 0 57868 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0485_
timestamp 1649977179
transform -1 0 22448 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0486_
timestamp 1649977179
transform -1 0 11040 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0487_
timestamp 1649977179
transform 1 0 8188 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0488_
timestamp 1649977179
transform -1 0 3312 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0489_
timestamp 1649977179
transform -1 0 2484 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0490_
timestamp 1649977179
transform -1 0 2668 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0491_
timestamp 1649977179
transform -1 0 2484 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0492_
timestamp 1649977179
transform 1 0 6072 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0493_
timestamp 1649977179
transform -1 0 2944 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0494_
timestamp 1649977179
transform -1 0 2760 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0495_
timestamp 1649977179
transform -1 0 18124 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0496_
timestamp 1649977179
transform -1 0 9384 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0497_
timestamp 1649977179
transform 1 0 14536 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0498_
timestamp 1649977179
transform -1 0 16744 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0499_
timestamp 1649977179
transform -1 0 25852 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0500_
timestamp 1649977179
transform 1 0 21988 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0501_
timestamp 1649977179
transform -1 0 22908 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0502_
timestamp 1649977179
transform -1 0 36708 0 1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__nor2_1  _0503_
timestamp 1649977179
transform -1 0 33580 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0504_
timestamp 1649977179
transform -1 0 39744 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0505_
timestamp 1649977179
transform 1 0 37352 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0506_
timestamp 1649977179
transform 1 0 38364 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0507_
timestamp 1649977179
transform -1 0 32384 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0508_
timestamp 1649977179
transform 1 0 31188 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0509_
timestamp 1649977179
transform -1 0 32384 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0510_
timestamp 1649977179
transform -1 0 23644 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0511_
timestamp 1649977179
transform 1 0 17020 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0512_
timestamp 1649977179
transform -1 0 19688 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0513_
timestamp 1649977179
transform -1 0 19504 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0514_
timestamp 1649977179
transform -1 0 26220 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0515_
timestamp 1649977179
transform 1 0 29900 0 -1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _0516_
timestamp 1649977179
transform 1 0 37996 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0517_
timestamp 1649977179
transform -1 0 41584 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0518_
timestamp 1649977179
transform 1 0 21896 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0519_
timestamp 1649977179
transform -1 0 20700 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0520_
timestamp 1649977179
transform -1 0 18860 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0521_
timestamp 1649977179
transform -1 0 44436 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0522_
timestamp 1649977179
transform -1 0 48852 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0523_
timestamp 1649977179
transform -1 0 48024 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0524_
timestamp 1649977179
transform -1 0 43056 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0525_
timestamp 1649977179
transform 1 0 48024 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0526_
timestamp 1649977179
transform 1 0 49864 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0527_
timestamp 1649977179
transform 1 0 52716 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0528_
timestamp 1649977179
transform 1 0 53912 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0529_
timestamp 1649977179
transform -1 0 23000 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _0530_
timestamp 1649977179
transform 1 0 2392 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0531_
timestamp 1649977179
transform -1 0 3220 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0532_
timestamp 1649977179
transform -1 0 3496 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0533_
timestamp 1649977179
transform -1 0 1840 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0534_
timestamp 1649977179
transform -1 0 2668 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0535_
timestamp 1649977179
transform -1 0 1840 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0536_
timestamp 1649977179
transform 1 0 12696 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0537_
timestamp 1649977179
transform -1 0 14352 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0538_
timestamp 1649977179
transform 1 0 22816 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0539_
timestamp 1649977179
transform -1 0 23736 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0540_
timestamp 1649977179
transform 1 0 37628 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _0541_
timestamp 1649977179
transform 1 0 39836 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0542_
timestamp 1649977179
transform 1 0 40112 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0543_
timestamp 1649977179
transform 1 0 28612 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0544_
timestamp 1649977179
transform -1 0 31004 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0545_
timestamp 1649977179
transform -1 0 16192 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0546_
timestamp 1649977179
transform -1 0 11040 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0547_
timestamp 1649977179
transform 1 0 38824 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0548_
timestamp 1649977179
transform -1 0 40848 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0549_
timestamp 1649977179
transform -1 0 16744 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0550_
timestamp 1649977179
transform -1 0 14720 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0551_
timestamp 1649977179
transform 1 0 49220 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0552_
timestamp 1649977179
transform 1 0 50600 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0553_
timestamp 1649977179
transform 1 0 52716 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0554_
timestamp 1649977179
transform -1 0 54188 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0555_
timestamp 1649977179
transform -1 0 51704 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0556_
timestamp 1649977179
transform -1 0 51612 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0557_
timestamp 1649977179
transform -1 0 20884 0 1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _0558_
timestamp 1649977179
transform 1 0 4324 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0559_
timestamp 1649977179
transform -1 0 4968 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0560_
timestamp 1649977179
transform -1 0 6808 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0561_
timestamp 1649977179
transform -1 0 4600 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0562_
timestamp 1649977179
transform -1 0 3772 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0563_
timestamp 1649977179
transform -1 0 2116 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0564_
timestamp 1649977179
transform -1 0 10948 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0565_
timestamp 1649977179
transform -1 0 10304 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0566_
timestamp 1649977179
transform 1 0 19688 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0567_
timestamp 1649977179
transform 1 0 20516 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0568_
timestamp 1649977179
transform 1 0 36156 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _0569_
timestamp 1649977179
transform 1 0 38916 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0570_
timestamp 1649977179
transform -1 0 42228 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0571_
timestamp 1649977179
transform -1 0 33672 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0572_
timestamp 1649977179
transform -1 0 33028 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0573_
timestamp 1649977179
transform 1 0 21252 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0574_
timestamp 1649977179
transform -1 0 21896 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0575_
timestamp 1649977179
transform 1 0 37812 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0576_
timestamp 1649977179
transform -1 0 38640 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0577_
timestamp 1649977179
transform -1 0 18124 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0578_
timestamp 1649977179
transform -1 0 14444 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0579_
timestamp 1649977179
transform 1 0 46644 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0580_
timestamp 1649977179
transform 1 0 46736 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0581_
timestamp 1649977179
transform 1 0 49128 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0582_
timestamp 1649977179
transform 1 0 50508 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0583_
timestamp 1649977179
transform 1 0 47748 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0584_
timestamp 1649977179
transform -1 0 48576 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0585_
timestamp 1649977179
transform 1 0 19596 0 -1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _0586_
timestamp 1649977179
transform -1 0 8096 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0587_
timestamp 1649977179
transform -1 0 6992 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0588_
timestamp 1649977179
transform -1 0 14352 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0589_
timestamp 1649977179
transform -1 0 10028 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0590_
timestamp 1649977179
transform -1 0 9476 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0591_
timestamp 1649977179
transform -1 0 5244 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0592_
timestamp 1649977179
transform -1 0 11960 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0593_
timestamp 1649977179
transform -1 0 10948 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0594_
timestamp 1649977179
transform 1 0 19044 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0595_
timestamp 1649977179
transform -1 0 19872 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0596_
timestamp 1649977179
transform 1 0 35512 0 -1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _0597_
timestamp 1649977179
transform 1 0 36432 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0598_
timestamp 1649977179
transform 1 0 38180 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0599_
timestamp 1649977179
transform -1 0 34500 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0600_
timestamp 1649977179
transform -1 0 34224 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0601_
timestamp 1649977179
transform -1 0 17020 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0602_
timestamp 1649977179
transform -1 0 15916 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0603_
timestamp 1649977179
transform -1 0 37720 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0604_
timestamp 1649977179
transform -1 0 34224 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0605_
timestamp 1649977179
transform -1 0 17296 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0606_
timestamp 1649977179
transform -1 0 14076 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0607_
timestamp 1649977179
transform -1 0 49496 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0608_
timestamp 1649977179
transform 1 0 49036 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0609_
timestamp 1649977179
transform 1 0 43424 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0610_
timestamp 1649977179
transform 1 0 43976 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0611_
timestamp 1649977179
transform 1 0 51428 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0612_
timestamp 1649977179
transform -1 0 52256 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0613_
timestamp 1649977179
transform -1 0 18768 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _0614_
timestamp 1649977179
transform -1 0 6808 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0615_
timestamp 1649977179
transform -1 0 5888 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0616_
timestamp 1649977179
transform -1 0 9936 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0617_
timestamp 1649977179
transform -1 0 2668 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0618_
timestamp 1649977179
transform -1 0 7636 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0619_
timestamp 1649977179
transform -1 0 2024 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0620_
timestamp 1649977179
transform 1 0 15364 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0621_
timestamp 1649977179
transform -1 0 16928 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0622_
timestamp 1649977179
transform 1 0 28428 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0623_
timestamp 1649977179
transform -1 0 29624 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0624_
timestamp 1649977179
transform 1 0 18768 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _0625_
timestamp 1649977179
transform -1 0 23276 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0626_
timestamp 1649977179
transform -1 0 21896 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0627_
timestamp 1649977179
transform 1 0 45172 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0628_
timestamp 1649977179
transform 1 0 46000 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0629_
timestamp 1649977179
transform 1 0 45632 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0630_
timestamp 1649977179
transform -1 0 47840 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0631_
timestamp 1649977179
transform 1 0 26956 0 -1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _0632_
timestamp 1649977179
transform -1 0 11960 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0633_
timestamp 1649977179
transform -1 0 6348 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0634_
timestamp 1649977179
transform -1 0 11960 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0635_
timestamp 1649977179
transform -1 0 7820 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0636_
timestamp 1649977179
transform -1 0 12880 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0637_
timestamp 1649977179
transform -1 0 11592 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0638_
timestamp 1649977179
transform -1 0 10856 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0639_
timestamp 1649977179
transform -1 0 8464 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0640_
timestamp 1649977179
transform 1 0 29992 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0641_
timestamp 1649977179
transform 1 0 32660 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0642_
timestamp 1649977179
transform -1 0 40572 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _0643_
timestamp 1649977179
transform -1 0 21344 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0644_
timestamp 1649977179
transform -1 0 19872 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0645_
timestamp 1649977179
transform 1 0 44252 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0646_
timestamp 1649977179
transform -1 0 46920 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0647_
timestamp 1649977179
transform 1 0 26036 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0648_
timestamp 1649977179
transform 1 0 26956 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0649_
timestamp 1649977179
transform 1 0 41216 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0650_
timestamp 1649977179
transform 1 0 43884 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0651_
timestamp 1649977179
transform -1 0 23092 0 1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0652_
timestamp 1649977179
transform -1 0 18584 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0653_
timestamp 1649977179
transform 1 0 21804 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0654_
timestamp 1649977179
transform -1 0 27508 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0655_
timestamp 1649977179
transform 1 0 21804 0 1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0656_
timestamp 1649977179
transform -1 0 40664 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0657_
timestamp 1649977179
transform -1 0 27508 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0658_
timestamp 1649977179
transform -1 0 26404 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0659_
timestamp 1649977179
transform 1 0 42412 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0660_
timestamp 1649977179
transform -1 0 43516 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0661_
timestamp 1649977179
transform -1 0 32292 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0662_
timestamp 1649977179
transform -1 0 31648 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0663_
timestamp 1649977179
transform -1 0 39376 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _0664_
timestamp 1649977179
transform -1 0 24840 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0665_
timestamp 1649977179
transform -1 0 23920 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0666_
timestamp 1649977179
transform 1 0 38640 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0667_
timestamp 1649977179
transform -1 0 40940 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0668_
timestamp 1649977179
transform 1 0 44068 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0669_
timestamp 1649977179
transform 1 0 46460 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0670_
timestamp 1649977179
transform -1 0 2300 0 1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and4bb_1  _0671_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 16100 0 -1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__nand2_1  _0672_
timestamp 1649977179
transform 1 0 1564 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0673_
timestamp 1649977179
transform 1 0 1564 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0674_
timestamp 1649977179
transform 1 0 8924 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _0675_
timestamp 1649977179
transform -1 0 7176 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0676_
timestamp 1649977179
transform 1 0 11500 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__nor3_1  _0677_
timestamp 1649977179
transform -1 0 2116 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__or4_1  _0678_
timestamp 1649977179
transform 1 0 2484 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0679_
timestamp 1649977179
transform 1 0 13340 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0680_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 14628 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _0681_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 2484 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__or3b_1  _0682_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 8004 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_2  _0683_
timestamp 1649977179
transform -1 0 7636 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0684_
timestamp 1649977179
transform 1 0 2668 0 1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__nor4b_1  _0685_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 8924 0 1 2176
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _0686_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 2668 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0687_
timestamp 1649977179
transform 1 0 28980 0 -1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__nand2_1  _0688_
timestamp 1649977179
transform 1 0 34684 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0689_
timestamp 1649977179
transform -1 0 33396 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0690_
timestamp 1649977179
transform -1 0 31648 0 -1 4352
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0691_
timestamp 1649977179
transform 1 0 33948 0 -1 4352
box -38 -48 958 592
use sky130_fd_sc_hd__a21o_1  _0692_
timestamp 1649977179
transform 1 0 25116 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _0693_
timestamp 1649977179
transform -1 0 19504 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _0694_
timestamp 1649977179
transform 1 0 25484 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _0695_
timestamp 1649977179
transform -1 0 23276 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _0696_
timestamp 1649977179
transform 1 0 32108 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _0697_
timestamp 1649977179
transform -1 0 30268 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _0698_
timestamp 1649977179
transform 1 0 27508 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _0699_
timestamp 1649977179
transform -1 0 15180 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0700_
timestamp 1649977179
transform 1 0 24380 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _0701_
timestamp 1649977179
transform -1 0 25392 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _0702_
timestamp 1649977179
transform -1 0 30360 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _0703_
timestamp 1649977179
transform -1 0 31924 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0704_
timestamp 1649977179
transform 1 0 34684 0 -1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0705_
timestamp 1649977179
transform -1 0 40664 0 -1 4352
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0706_
timestamp 1649977179
transform -1 0 39376 0 -1 4352
box -38 -48 958 592
use sky130_fd_sc_hd__a21o_1  _0707_
timestamp 1649977179
transform -1 0 46460 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _0708_
timestamp 1649977179
transform -1 0 44804 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _0709_
timestamp 1649977179
transform 1 0 45356 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _0710_
timestamp 1649977179
transform -1 0 43516 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _0711_
timestamp 1649977179
transform 1 0 43976 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _0712_
timestamp 1649977179
transform -1 0 43700 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _0713_
timestamp 1649977179
transform 1 0 40848 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _0714_
timestamp 1649977179
transform 1 0 18032 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _0715_
timestamp 1649977179
transform -1 0 36708 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _0716_
timestamp 1649977179
transform 1 0 38548 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _0717_
timestamp 1649977179
transform 1 0 37260 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _0718_
timestamp 1649977179
transform -1 0 9660 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_2  _0719_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 10304 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _0720_
timestamp 1649977179
transform 1 0 27692 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0721_
timestamp 1649977179
transform -1 0 28336 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0722_
timestamp 1649977179
transform -1 0 29348 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0723_
timestamp 1649977179
transform 1 0 19228 0 1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__a21o_1  _0724_
timestamp 1649977179
transform 1 0 16836 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _0725_
timestamp 1649977179
transform 1 0 13708 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _0726_
timestamp 1649977179
transform 1 0 15824 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _0727_
timestamp 1649977179
transform 1 0 14168 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _0728_
timestamp 1649977179
transform 1 0 15640 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _0729_
timestamp 1649977179
transform 1 0 16652 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _0730_
timestamp 1649977179
transform -1 0 21896 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _0731_
timestamp 1649977179
transform 1 0 23736 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _0732_
timestamp 1649977179
transform 1 0 21804 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _0733_
timestamp 1649977179
transform -1 0 26312 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _0734_
timestamp 1649977179
transform 1 0 25208 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _0735_
timestamp 1649977179
transform 1 0 28704 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0736_
timestamp 1649977179
transform -1 0 33580 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0737_
timestamp 1649977179
transform 1 0 29532 0 1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__a21o_1  _0738_
timestamp 1649977179
transform -1 0 41492 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _0739_
timestamp 1649977179
transform -1 0 43884 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _0740_
timestamp 1649977179
transform -1 0 41584 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _0741_
timestamp 1649977179
transform -1 0 43332 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _0742_
timestamp 1649977179
transform -1 0 41308 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _0743_
timestamp 1649977179
transform -1 0 44436 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _0744_
timestamp 1649977179
transform 1 0 37260 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _0745_
timestamp 1649977179
transform -1 0 13616 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _0746_
timestamp 1649977179
transform -1 0 35972 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _0747_
timestamp 1649977179
transform 1 0 31096 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _0748_
timestamp 1649977179
transform -1 0 31556 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _0749_
timestamp 1649977179
transform -1 0 47104 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0750_
timestamp 1649977179
transform -1 0 37720 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0751_
timestamp 1649977179
transform -1 0 42688 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0752_
timestamp 1649977179
transform -1 0 38640 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0753_
timestamp 1649977179
transform 1 0 4968 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__or4b_1  _0754_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 3772 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _0755_
timestamp 1649977179
transform 1 0 4140 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _0756_
timestamp 1649977179
transform -1 0 18860 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__and4bb_1  _0757_
timestamp 1649977179
transform -1 0 7820 0 -1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__and4_1  _0758_
timestamp 1649977179
transform 1 0 3680 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0759_
timestamp 1649977179
transform 1 0 11500 0 -1 5440
box -38 -48 958 592
use sky130_fd_sc_hd__or2_1  _0760_
timestamp 1649977179
transform -1 0 9936 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0761_
timestamp 1649977179
transform 1 0 10304 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__a21bo_1  _0762_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 17940 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _0763_
timestamp 1649977179
transform 1 0 10120 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _0764_
timestamp 1649977179
transform 1 0 17572 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _0765_
timestamp 1649977179
transform -1 0 18952 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0766_
timestamp 1649977179
transform -1 0 18768 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0767_
timestamp 1649977179
transform 1 0 19228 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _0768_
timestamp 1649977179
transform 1 0 15824 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _0769_
timestamp 1649977179
transform -1 0 22540 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0770_
timestamp 1649977179
transform 1 0 12788 0 -1 5440
box -38 -48 958 592
use sky130_fd_sc_hd__or2_1  _0771_
timestamp 1649977179
transform 1 0 29532 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0772_
timestamp 1649977179
transform -1 0 29992 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0773_
timestamp 1649977179
transform 1 0 24012 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0774_
timestamp 1649977179
transform 1 0 24840 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0775_
timestamp 1649977179
transform 1 0 26772 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0776_
timestamp 1649977179
transform -1 0 28612 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _0777_
timestamp 1649977179
transform 1 0 3680 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _0778_
timestamp 1649977179
transform 1 0 15732 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0779_
timestamp 1649977179
transform -1 0 17112 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0780_
timestamp 1649977179
transform -1 0 14996 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0781_
timestamp 1649977179
transform 1 0 14076 0 -1 5440
box -38 -48 958 592
use sky130_fd_sc_hd__o211a_1  _0782_
timestamp 1649977179
transform -1 0 14168 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  _0783_
timestamp 1649977179
transform 1 0 1840 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0784_
timestamp 1649977179
transform 1 0 9660 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0785_
timestamp 1649977179
transform -1 0 11040 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0786_
timestamp 1649977179
transform 1 0 2760 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0787_
timestamp 1649977179
transform -1 0 7452 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0788_
timestamp 1649977179
transform 1 0 2852 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0789_
timestamp 1649977179
transform -1 0 5336 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0790_
timestamp 1649977179
transform 1 0 1932 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0791_
timestamp 1649977179
transform -1 0 4508 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0792_
timestamp 1649977179
transform 1 0 9752 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0793_
timestamp 1649977179
transform -1 0 11316 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0794_
timestamp 1649977179
transform -1 0 2116 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0795_
timestamp 1649977179
transform -1 0 3220 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _0796_
timestamp 1649977179
transform 1 0 46828 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0797_
timestamp 1649977179
transform 1 0 50140 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0798_
timestamp 1649977179
transform 1 0 47196 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_2  _0799_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 4876 0 1 4352
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _0800_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 19504 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0801_
timestamp 1649977179
transform 1 0 23276 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0802_
timestamp 1649977179
transform 1 0 30176 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0803_
timestamp 1649977179
transform 1 0 27140 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0804_
timestamp 1649977179
transform 1 0 32752 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0805_
timestamp 1649977179
transform -1 0 49772 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0806_
timestamp 1649977179
transform 1 0 43516 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0807_
timestamp 1649977179
transform -1 0 48760 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0808_
timestamp 1649977179
transform 1 0 39560 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0809_
timestamp 1649977179
transform 1 0 37260 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0810_
timestamp 1649977179
transform 1 0 11500 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0811_
timestamp 1649977179
transform 1 0 11500 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0812_
timestamp 1649977179
transform -1 0 16836 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0813_
timestamp 1649977179
transform -1 0 21344 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0814_
timestamp 1649977179
transform 1 0 25392 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0815_
timestamp 1649977179
transform -1 0 49496 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0816_
timestamp 1649977179
transform -1 0 46644 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0817_
timestamp 1649977179
transform -1 0 49588 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0818_
timestamp 1649977179
transform 1 0 35512 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0819_
timestamp 1649977179
transform 1 0 32108 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfstp_1  _0820_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 35696 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _0821_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 40112 0 -1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _0822_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 41032 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _0823_
timestamp 1649977179
transform 1 0 36064 0 1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__dfxtp_1  _0824_
timestamp 1649977179
transform -1 0 5888 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0825_
timestamp 1649977179
transform 1 0 6808 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0826_
timestamp 1649977179
transform -1 0 9476 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0827_
timestamp 1649977179
transform -1 0 21344 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0828_
timestamp 1649977179
transform -1 0 23184 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0829_
timestamp 1649977179
transform -1 0 32752 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0830_
timestamp 1649977179
transform 1 0 24656 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0831_
timestamp 1649977179
transform -1 0 29072 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0832_
timestamp 1649977179
transform -1 0 18124 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0833_
timestamp 1649977179
transform 1 0 14076 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0834_
timestamp 1649977179
transform 1 0 10672 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0835_
timestamp 1649977179
transform 1 0 7636 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0836_
timestamp 1649977179
transform 1 0 5244 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0837_
timestamp 1649977179
transform 1 0 4416 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0838_
timestamp 1649977179
transform 1 0 11684 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0839_
timestamp 1649977179
transform 1 0 5244 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dlxtn_1  _0840_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 19228 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _0841_
timestamp 1649977179
transform 1 0 17388 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _0842_
timestamp 1649977179
transform -1 0 38456 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _0843_
timestamp 1649977179
transform 1 0 50140 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _0844_
timestamp 1649977179
transform -1 0 4232 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _0845_
timestamp 1649977179
transform 1 0 41400 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _0846_
timestamp 1649977179
transform 1 0 5612 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _0847_
timestamp 1649977179
transform 1 0 33120 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _0848_
timestamp 1649977179
transform 1 0 22540 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _0849_
timestamp 1649977179
transform -1 0 49680 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _0850_
timestamp 1649977179
transform 1 0 20056 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _0851_
timestamp 1649977179
transform 1 0 3220 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_2  _0852_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 52348 0 1 8704
box -38 -48 1234 592
use sky130_fd_sc_hd__dlxtn_1  _0853_
timestamp 1649977179
transform 1 0 15088 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _0854_
timestamp 1649977179
transform 1 0 14904 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _0855_
timestamp 1649977179
transform -1 0 40296 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _0856_
timestamp 1649977179
transform 1 0 50324 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _0857_
timestamp 1649977179
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _0858_
timestamp 1649977179
transform 1 0 40388 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _0859_
timestamp 1649977179
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _0860_
timestamp 1649977179
transform -1 0 31188 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _0861_
timestamp 1649977179
transform 1 0 24380 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _0862_
timestamp 1649977179
transform 1 0 53912 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _0863_
timestamp 1649977179
transform 1 0 17112 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _0864_
timestamp 1649977179
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_2  _0865_
timestamp 1649977179
transform 1 0 52256 0 1 9792
box -38 -48 1234 592
use sky130_fd_sc_hd__dlxtn_1  _0866_
timestamp 1649977179
transform 1 0 22540 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _0867_
timestamp 1649977179
transform 1 0 11500 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _0868_
timestamp 1649977179
transform 1 0 42412 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _0869_
timestamp 1649977179
transform -1 0 46736 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _0870_
timestamp 1649977179
transform 1 0 7268 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _0871_
timestamp 1649977179
transform 1 0 38916 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _0872_
timestamp 1649977179
transform -1 0 5244 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _0873_
timestamp 1649977179
transform 1 0 32752 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _0874_
timestamp 1649977179
transform -1 0 20792 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _0875_
timestamp 1649977179
transform 1 0 50232 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _0876_
timestamp 1649977179
transform 1 0 14812 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _0877_
timestamp 1649977179
transform 1 0 4600 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_2  _0878_
timestamp 1649977179
transform 1 0 48944 0 -1 9792
box -38 -48 1234 592
use sky130_fd_sc_hd__dlxtn_1  _0879_
timestamp 1649977179
transform 1 0 16928 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _0880_
timestamp 1649977179
transform 1 0 11960 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _0881_
timestamp 1649977179
transform -1 0 36800 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _0882_
timestamp 1649977179
transform 1 0 48576 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _0883_
timestamp 1649977179
transform -1 0 13616 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _0884_
timestamp 1649977179
transform 1 0 35236 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _0885_
timestamp 1649977179
transform 1 0 9660 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _0886_
timestamp 1649977179
transform -1 0 35328 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _0887_
timestamp 1649977179
transform -1 0 20976 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _0888_
timestamp 1649977179
transform -1 0 44528 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _0889_
timestamp 1649977179
transform 1 0 14168 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _0890_
timestamp 1649977179
transform 1 0 8464 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_2  _0891_
timestamp 1649977179
transform 1 0 52716 0 -1 9792
box -38 -48 1234 592
use sky130_fd_sc_hd__dlxtn_1  _0892_
timestamp 1649977179
transform 1 0 8832 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _0893_
timestamp 1649977179
transform 1 0 8004 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _0894_
timestamp 1649977179
transform 1 0 6256 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _0895_
timestamp 1649977179
transform 1 0 11224 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _0896_
timestamp 1649977179
transform -1 0 43700 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _0897_
timestamp 1649977179
transform 1 0 11040 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _0898_
timestamp 1649977179
transform 1 0 32384 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _0899_
timestamp 1649977179
transform -1 0 12972 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _0900_
timestamp 1649977179
transform -1 0 30820 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _0901_
timestamp 1649977179
transform 1 0 26956 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _0902_
timestamp 1649977179
transform 1 0 46552 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _0903_
timestamp 1649977179
transform -1 0 26036 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _0904_
timestamp 1649977179
transform 1 0 7360 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_2  _0905_
timestamp 1649977179
transform -1 0 46828 0 1 9792
box -38 -48 1234 592
use sky130_fd_sc_hd__dlxtn_1  _0906_
timestamp 1649977179
transform 1 0 20240 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _0907_
timestamp 1649977179
transform 1 0 17112 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _0908_
timestamp 1649977179
transform 1 0 42688 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _0909_
timestamp 1649977179
transform 1 0 45264 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _0910_
timestamp 1649977179
transform 1 0 36800 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _0911_
timestamp 1649977179
transform 1 0 29256 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _0912_
timestamp 1649977179
transform 1 0 26128 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _0913_
timestamp 1649977179
transform 1 0 44988 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _0914_
timestamp 1649977179
transform 1 0 22264 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_2  _0915_
timestamp 1649977179
transform 1 0 47380 0 1 9792
box -38 -48 1234 592
use sky130_fd_sc_hd__dlxtn_1  _0916_
timestamp 1649977179
transform 1 0 22264 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _0917_
timestamp 1649977179
transform 1 0 40848 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_2  _0918_
timestamp 1649977179
transform -1 0 45448 0 -1 6528
box -38 -48 1602 592
use sky130_fd_sc_hd__dfrtp_1  _0919_
timestamp 1649977179
transform -1 0 49496 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0920_
timestamp 1649977179
transform 1 0 47840 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0921_
timestamp 1649977179
transform -1 0 49956 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dlxtn_1  _0922_
timestamp 1649977179
transform -1 0 52256 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _0923_
timestamp 1649977179
transform -1 0 52624 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _0924_
timestamp 1649977179
transform -1 0 57684 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _0925_
timestamp 1649977179
transform -1 0 54188 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _0926_
timestamp 1649977179
transform -1 0 53360 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _0927_
timestamp 1649977179
transform -1 0 52808 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _0928_
timestamp 1649977179
transform -1 0 57316 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _0929_
timestamp 1649977179
transform -1 0 20608 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _0930_
timestamp 1649977179
transform -1 0 53912 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _0931_
timestamp 1649977179
transform -1 0 57868 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  _1138_
timestamp 1649977179
transform -1 0 12972 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1139_
timestamp 1649977179
transform -1 0 2116 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1140_
timestamp 1649977179
transform -1 0 15732 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1141_
timestamp 1649977179
transform -1 0 13616 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_wb_clk_i dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 26588 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_0__f_wb_clk_i
timestamp 1649977179
transform 1 0 20792 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_1__f_wb_clk_i
timestamp 1649977179
transform -1 0 21344 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_2__f_wb_clk_i
timestamp 1649977179
transform 1 0 31188 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_3__f_wb_clk_i
timestamp 1649977179
transform 1 0 32476 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__buf_2  input1
timestamp 1649977179
transform -1 0 2300 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1649977179
transform -1 0 1932 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1649977179
transform -1 0 2576 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1649977179
transform 1 0 16100 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1649977179
transform -1 0 5888 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1649977179
transform -1 0 2024 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1649977179
transform 1 0 15916 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp 1649977179
transform -1 0 4048 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input9
timestamp 1649977179
transform 1 0 9016 0 1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input10
timestamp 1649977179
transform -1 0 9660 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input11
timestamp 1649977179
transform -1 0 2484 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input12
timestamp 1649977179
transform 1 0 9384 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input13
timestamp 1649977179
transform 1 0 10212 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input14
timestamp 1649977179
transform 1 0 6900 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input15
timestamp 1649977179
transform 1 0 7544 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input16
timestamp 1649977179
transform -1 0 1840 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input17
timestamp 1649977179
transform -1 0 9108 0 -1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input18
timestamp 1649977179
transform -1 0 4232 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input19
timestamp 1649977179
transform 1 0 9476 0 -1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input20
timestamp 1649977179
transform 1 0 5520 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input21
timestamp 1649977179
transform 1 0 10028 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input22
timestamp 1649977179
transform 1 0 4784 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input23
timestamp 1649977179
transform -1 0 11040 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input24
timestamp 1649977179
transform 1 0 11500 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input25
timestamp 1649977179
transform 1 0 8188 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input26
timestamp 1649977179
transform 1 0 7728 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input27
timestamp 1649977179
transform 1 0 7544 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output28
timestamp 1649977179
transform -1 0 13340 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output29
timestamp 1649977179
transform 1 0 18400 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output30
timestamp 1649977179
transform 1 0 15824 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output31
timestamp 1649977179
transform 1 0 15088 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output32
timestamp 1649977179
transform 1 0 21804 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output33
timestamp 1649977179
transform -1 0 17296 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output34
timestamp 1649977179
transform -1 0 24748 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output35
timestamp 1649977179
transform 1 0 17664 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output36
timestamp 1649977179
transform -1 0 21344 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output37
timestamp 1649977179
transform -1 0 23828 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output38
timestamp 1649977179
transform -1 0 23368 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output39
timestamp 1649977179
transform -1 0 18676 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output40
timestamp 1649977179
transform -1 0 23092 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output41
timestamp 1649977179
transform -1 0 23828 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output42
timestamp 1649977179
transform -1 0 13616 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output43
timestamp 1649977179
transform -1 0 18216 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output44
timestamp 1649977179
transform 1 0 14444 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output45
timestamp 1649977179
transform 1 0 14352 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output46
timestamp 1649977179
transform -1 0 4416 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output47
timestamp 1649977179
transform -1 0 8464 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output48
timestamp 1649977179
transform 1 0 11500 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output49
timestamp 1649977179
transform 1 0 13708 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output50
timestamp 1649977179
transform 1 0 12696 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output51
timestamp 1649977179
transform 1 0 13064 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output52
timestamp 1649977179
transform 1 0 14076 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output53
timestamp 1649977179
transform -1 0 5152 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output54
timestamp 1649977179
transform -1 0 7728 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output55
timestamp 1649977179
transform -1 0 9568 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output56
timestamp 1649977179
transform -1 0 7268 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output57
timestamp 1649977179
transform -1 0 8464 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output58
timestamp 1649977179
transform -1 0 6808 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output59
timestamp 1649977179
transform -1 0 9292 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output60
timestamp 1649977179
transform -1 0 5888 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output61
timestamp 1649977179
transform 1 0 12512 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  pixel_macro_90 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 4600 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_91
timestamp 1649977179
transform 1 0 5612 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_92
timestamp 1649977179
transform 1 0 6900 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_93
timestamp 1649977179
transform 1 0 8188 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_94
timestamp 1649977179
transform -1 0 10120 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_95
timestamp 1649977179
transform -1 0 11684 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_96
timestamp 1649977179
transform -1 0 12880 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_97
timestamp 1649977179
transform -1 0 14444 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_98
timestamp 1649977179
transform 1 0 15272 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_99
timestamp 1649977179
transform -1 0 17204 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_100
timestamp 1649977179
transform 1 0 17848 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_101
timestamp 1649977179
transform -1 0 19780 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_102
timestamp 1649977179
transform -1 0 21344 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_103
timestamp 1649977179
transform -1 0 22540 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_104
timestamp 1649977179
transform -1 0 23920 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_105
timestamp 1649977179
transform 1 0 24932 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_106
timestamp 1649977179
transform 1 0 26220 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_107
timestamp 1649977179
transform 1 0 27508 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_108
timestamp 1649977179
transform 1 0 28796 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_109
timestamp 1649977179
transform -1 0 30820 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_110
timestamp 1649977179
transform -1 0 32384 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_111
timestamp 1649977179
transform -1 0 33764 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_112
timestamp 1649977179
transform -1 0 35604 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_113
timestamp 1649977179
transform -1 0 36524 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_114
timestamp 1649977179
transform -1 0 38180 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_115
timestamp 1649977179
transform -1 0 40112 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_116
timestamp 1649977179
transform -1 0 40756 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_117
timestamp 1649977179
transform -1 0 42688 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_118
timestamp 1649977179
transform -1 0 43976 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_119
timestamp 1649977179
transform -1 0 45264 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_120
timestamp 1649977179
transform -1 0 46552 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_121
timestamp 1649977179
transform -1 0 47840 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_122
timestamp 1649977179
transform -1 0 49128 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_123
timestamp 1649977179
transform -1 0 50416 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_124
timestamp 1649977179
transform -1 0 51704 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_125
timestamp 1649977179
transform -1 0 53636 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_126
timestamp 1649977179
transform -1 0 54464 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_127
timestamp 1649977179
transform -1 0 56212 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_128
timestamp 1649977179
transform -1 0 5244 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_129
timestamp 1649977179
transform -1 0 6624 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_130
timestamp 1649977179
transform -1 0 7820 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_131
timestamp 1649977179
transform -1 0 9384 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_132
timestamp 1649977179
transform -1 0 10764 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_133
timestamp 1649977179
transform -1 0 12144 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_134
timestamp 1649977179
transform -1 0 13524 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_135
timestamp 1649977179
transform -1 0 14904 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_136
timestamp 1649977179
transform -1 0 16192 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_137
timestamp 1649977179
transform -1 0 17480 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_138
timestamp 1649977179
transform 1 0 18492 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_139
timestamp 1649977179
transform -1 0 20424 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_140
timestamp 1649977179
transform 1 0 21068 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_141
timestamp 1649977179
transform -1 0 23184 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_142
timestamp 1649977179
transform -1 0 24656 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_143
timestamp 1649977179
transform -1 0 25852 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_144
timestamp 1649977179
transform -1 0 27324 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_145
timestamp 1649977179
transform 1 0 28152 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_146
timestamp 1649977179
transform -1 0 30084 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_147
timestamp 1649977179
transform -1 0 31464 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_148
timestamp 1649977179
transform -1 0 33028 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_149
timestamp 1649977179
transform -1 0 34960 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_150
timestamp 1649977179
transform -1 0 36248 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_151
timestamp 1649977179
transform -1 0 37536 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_152
timestamp 1649977179
transform -1 0 38824 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_153
timestamp 1649977179
transform -1 0 40112 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_154
timestamp 1649977179
transform -1 0 41400 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_155
timestamp 1649977179
transform -1 0 43332 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_156
timestamp 1649977179
transform -1 0 43884 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_157
timestamp 1649977179
transform -1 0 45908 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_158
timestamp 1649977179
transform -1 0 46644 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_159
timestamp 1649977179
transform -1 0 48484 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_160
timestamp 1649977179
transform -1 0 49404 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_161
timestamp 1649977179
transform -1 0 51060 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_162
timestamp 1649977179
transform -1 0 52992 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_163
timestamp 1649977179
transform -1 0 54280 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_164
timestamp 1649977179
transform -1 0 55568 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_165
timestamp 1649977179
transform -1 0 56856 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_166
timestamp 1649977179
transform -1 0 56856 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_167
timestamp 1649977179
transform -1 0 56948 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_168
timestamp 1649977179
transform -1 0 56212 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_169
timestamp 1649977179
transform 1 0 17848 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_170
timestamp 1649977179
transform -1 0 18768 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_171
timestamp 1649977179
transform 1 0 6624 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_172
timestamp 1649977179
transform 1 0 9016 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_173
timestamp 1649977179
transform 1 0 3772 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_174
timestamp 1649977179
transform -1 0 30636 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_175
timestamp 1649977179
transform 1 0 16284 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_176
timestamp 1649977179
transform -1 0 29716 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_177
timestamp 1649977179
transform 1 0 10764 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_178
timestamp 1649977179
transform -1 0 29072 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_179
timestamp 1649977179
transform 1 0 20976 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_180
timestamp 1649977179
transform 1 0 23644 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_181
timestamp 1649977179
transform 1 0 20424 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_182
timestamp 1649977179
transform 1 0 18952 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_183
timestamp 1649977179
transform -1 0 28612 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_184
timestamp 1649977179
transform 1 0 18492 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_185
timestamp 1649977179
transform 1 0 21068 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_186
timestamp 1649977179
transform -1 0 27232 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_187
timestamp 1649977179
transform -1 0 31464 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_188
timestamp 1649977179
transform 1 0 23092 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_189
timestamp 1649977179
transform 1 0 27232 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_190
timestamp 1649977179
transform 1 0 17756 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_191
timestamp 1649977179
transform 1 0 24748 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_192
timestamp 1649977179
transform 1 0 22632 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_193
timestamp 1649977179
transform 1 0 24564 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_194
timestamp 1649977179
transform 1 0 26220 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_195
timestamp 1649977179
transform 1 0 23644 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_196
timestamp 1649977179
transform 1 0 25576 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_197
timestamp 1649977179
transform 1 0 27508 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_198
timestamp 1649977179
transform 1 0 28152 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_199
timestamp 1649977179
transform -1 0 30728 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_200
timestamp 1649977179
transform 1 0 28796 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_201
timestamp 1649977179
transform 1 0 29808 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_202
timestamp 1649977179
transform -1 0 34224 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_203
timestamp 1649977179
transform -1 0 34960 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_204
timestamp 1649977179
transform -1 0 35604 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_205
timestamp 1649977179
transform -1 0 37536 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_206
timestamp 1649977179
transform -1 0 36248 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_207
timestamp 1649977179
transform -1 0 38180 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_208
timestamp 1649977179
transform -1 0 36248 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_209
timestamp 1649977179
transform -1 0 34224 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_210
timestamp 1649977179
transform -1 0 35512 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_211
timestamp 1649977179
transform -1 0 38824 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_212
timestamp 1649977179
transform -1 0 36616 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_213
timestamp 1649977179
transform -1 0 38456 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_214
timestamp 1649977179
transform -1 0 39100 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_215
timestamp 1649977179
transform -1 0 40112 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_216
timestamp 1649977179
transform -1 0 40756 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_217
timestamp 1649977179
transform -1 0 39744 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_218
timestamp 1649977179
transform -1 0 36800 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_219
timestamp 1649977179
transform -1 0 40388 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_220
timestamp 1649977179
transform -1 0 42688 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_221
timestamp 1649977179
transform -1 0 41400 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_222
timestamp 1649977179
transform -1 0 43332 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_223
timestamp 1649977179
transform -1 0 41952 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_224
timestamp 1649977179
transform -1 0 42688 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_225
timestamp 1649977179
transform -1 0 39376 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_226
timestamp 1649977179
transform -1 0 45264 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_227
timestamp 1649977179
transform -1 0 44528 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_228
timestamp 1649977179
transform -1 0 42136 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_229
timestamp 1649977179
transform -1 0 45908 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_230
timestamp 1649977179
transform -1 0 43976 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_231
timestamp 1649977179
transform -1 0 45172 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_232
timestamp 1649977179
transform -1 0 46552 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_233
timestamp 1649977179
transform -1 0 45816 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_234
timestamp 1649977179
transform -1 0 42044 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_235
timestamp 1649977179
transform -1 0 46460 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_236
timestamp 1649977179
transform -1 0 41676 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_237
timestamp 1649977179
transform -1 0 47840 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_238
timestamp 1649977179
transform -1 0 47104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_239
timestamp 1649977179
transform -1 0 48484 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_240
timestamp 1649977179
transform -1 0 47288 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_241
timestamp 1649977179
transform -1 0 45448 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_242
timestamp 1649977179
transform -1 0 49128 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_243
timestamp 1649977179
transform -1 0 50416 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_244
timestamp 1649977179
transform -1 0 50232 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_245
timestamp 1649977179
transform -1 0 46092 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_246
timestamp 1649977179
transform -1 0 47840 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_247
timestamp 1649977179
transform -1 0 51060 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_248
timestamp 1649977179
transform -1 0 46736 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_249
timestamp 1649977179
transform -1 0 49404 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_250
timestamp 1649977179
transform -1 0 51704 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_251
timestamp 1649977179
transform -1 0 45908 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_252
timestamp 1649977179
transform -1 0 50876 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_253
timestamp 1649977179
transform -1 0 53636 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_254
timestamp 1649977179
transform -1 0 46552 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_255
timestamp 1649977179
transform -1 0 51520 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_256
timestamp 1649977179
transform -1 0 54280 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_257
timestamp 1649977179
transform -1 0 50416 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_258
timestamp 1649977179
transform -1 0 52992 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_259
timestamp 1649977179
transform -1 0 50416 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_260
timestamp 1649977179
transform -1 0 51704 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_261
timestamp 1649977179
transform -1 0 50416 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_262
timestamp 1649977179
transform -1 0 53728 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_263
timestamp 1649977179
transform -1 0 51060 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_264
timestamp 1649977179
transform -1 0 54372 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_265
timestamp 1649977179
transform -1 0 51060 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_266
timestamp 1649977179
transform -1 0 52164 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_267
timestamp 1649977179
transform -1 0 55568 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_268
timestamp 1649977179
transform -1 0 56212 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_269
timestamp 1649977179
transform -1 0 51060 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_270
timestamp 1649977179
transform -1 0 55016 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_271
timestamp 1649977179
transform -1 0 50600 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_272
timestamp 1649977179
transform -1 0 55660 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_273
timestamp 1649977179
transform -1 0 56856 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_274
timestamp 1649977179
transform -1 0 52992 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_275
timestamp 1649977179
transform -1 0 54004 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_276
timestamp 1649977179
transform -1 0 53636 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_277
timestamp 1649977179
transform -1 0 55568 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_278
timestamp 1649977179
transform -1 0 56304 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_279
timestamp 1649977179
transform 1 0 12052 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_280
timestamp 1649977179
transform -1 0 13156 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_281
timestamp 1649977179
transform 1 0 12696 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_282
timestamp 1649977179
transform -1 0 13616 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_283
timestamp 1649977179
transform 1 0 1840 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_284
timestamp 1649977179
transform -1 0 14352 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_285
timestamp 1649977179
transform 1 0 13340 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_286
timestamp 1649977179
transform 1 0 3036 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_287
timestamp 1649977179
transform 1 0 13984 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_288
timestamp 1649977179
transform -1 0 15364 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_289
timestamp 1649977179
transform 1 0 14812 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_290
timestamp 1649977179
transform 1 0 14628 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_291
timestamp 1649977179
transform -1 0 16192 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_292
timestamp 1649977179
transform 1 0 15272 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_293
timestamp 1649977179
transform 1 0 13892 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_294
timestamp 1649977179
transform -1 0 17020 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  pixel_macro_295
timestamp 1649977179
transform 1 0 11224 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  repeater62
timestamp 1649977179
transform 1 0 17112 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  repeater63
timestamp 1649977179
transform -1 0 47840 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  repeater64
timestamp 1649977179
transform 1 0 42044 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  repeater65
timestamp 1649977179
transform 1 0 6900 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  repeater66
timestamp 1649977179
transform 1 0 24196 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  repeater67
timestamp 1649977179
transform -1 0 25760 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  repeater68
timestamp 1649977179
transform 1 0 5612 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  repeater69
timestamp 1649977179
transform -1 0 45264 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  repeater70
timestamp 1649977179
transform 1 0 33396 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  repeater71
timestamp 1649977179
transform -1 0 35696 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  repeater72
timestamp 1649977179
transform -1 0 5704 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  repeater73
timestamp 1649977179
transform -1 0 52256 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  repeater74
timestamp 1649977179
transform -1 0 50232 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  repeater75
timestamp 1649977179
transform 1 0 15640 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  repeater76
timestamp 1649977179
transform -1 0 15272 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  repeater77
timestamp 1649977179
transform -1 0 50876 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  repeater78
timestamp 1649977179
transform -1 0 40572 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  repeater79
timestamp 1649977179
transform -1 0 48576 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  repeater80
timestamp 1649977179
transform -1 0 35420 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  repeater81
timestamp 1649977179
transform 1 0 17664 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  repeater82
timestamp 1649977179
transform 1 0 51704 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  repeater83
timestamp 1649977179
transform 1 0 56764 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  repeater84
timestamp 1649977179
transform -1 0 55936 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  repeater85
timestamp 1649977179
transform 1 0 21896 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  repeater86
timestamp 1649977179
transform 1 0 26864 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  repeater87
timestamp 1649977179
transform -1 0 44988 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  repeater88
timestamp 1649977179
transform -1 0 36616 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  repeater89
timestamp 1649977179
transform -1 0 38456 0 -1 7616
box -38 -48 406 592
<< labels >>
flabel metal2 s 3974 19200 4030 20000 0 FreeSans 224 90 0 0 io_in[0]
port 0 nsew signal input
flabel metal2 s 17774 19200 17830 20000 0 FreeSans 224 90 0 0 io_in[10]
port 1 nsew signal input
flabel metal2 s 19154 19200 19210 20000 0 FreeSans 224 90 0 0 io_in[11]
port 2 nsew signal input
flabel metal2 s 20534 19200 20590 20000 0 FreeSans 224 90 0 0 io_in[12]
port 3 nsew signal input
flabel metal2 s 21914 19200 21970 20000 0 FreeSans 224 90 0 0 io_in[13]
port 4 nsew signal input
flabel metal2 s 23294 19200 23350 20000 0 FreeSans 224 90 0 0 io_in[14]
port 5 nsew signal input
flabel metal2 s 24674 19200 24730 20000 0 FreeSans 224 90 0 0 io_in[15]
port 6 nsew signal input
flabel metal2 s 26054 19200 26110 20000 0 FreeSans 224 90 0 0 io_in[16]
port 7 nsew signal input
flabel metal2 s 27434 19200 27490 20000 0 FreeSans 224 90 0 0 io_in[17]
port 8 nsew signal input
flabel metal2 s 28814 19200 28870 20000 0 FreeSans 224 90 0 0 io_in[18]
port 9 nsew signal input
flabel metal2 s 30194 19200 30250 20000 0 FreeSans 224 90 0 0 io_in[19]
port 10 nsew signal input
flabel metal2 s 5354 19200 5410 20000 0 FreeSans 224 90 0 0 io_in[1]
port 11 nsew signal input
flabel metal2 s 31574 19200 31630 20000 0 FreeSans 224 90 0 0 io_in[20]
port 12 nsew signal input
flabel metal2 s 32954 19200 33010 20000 0 FreeSans 224 90 0 0 io_in[21]
port 13 nsew signal input
flabel metal2 s 34334 19200 34390 20000 0 FreeSans 224 90 0 0 io_in[22]
port 14 nsew signal input
flabel metal2 s 35714 19200 35770 20000 0 FreeSans 224 90 0 0 io_in[23]
port 15 nsew signal input
flabel metal2 s 37094 19200 37150 20000 0 FreeSans 224 90 0 0 io_in[24]
port 16 nsew signal input
flabel metal2 s 38474 19200 38530 20000 0 FreeSans 224 90 0 0 io_in[25]
port 17 nsew signal input
flabel metal2 s 39854 19200 39910 20000 0 FreeSans 224 90 0 0 io_in[26]
port 18 nsew signal input
flabel metal2 s 41234 19200 41290 20000 0 FreeSans 224 90 0 0 io_in[27]
port 19 nsew signal input
flabel metal2 s 42614 19200 42670 20000 0 FreeSans 224 90 0 0 io_in[28]
port 20 nsew signal input
flabel metal2 s 43994 19200 44050 20000 0 FreeSans 224 90 0 0 io_in[29]
port 21 nsew signal input
flabel metal2 s 6734 19200 6790 20000 0 FreeSans 224 90 0 0 io_in[2]
port 22 nsew signal input
flabel metal2 s 45374 19200 45430 20000 0 FreeSans 224 90 0 0 io_in[30]
port 23 nsew signal input
flabel metal2 s 46754 19200 46810 20000 0 FreeSans 224 90 0 0 io_in[31]
port 24 nsew signal input
flabel metal2 s 48134 19200 48190 20000 0 FreeSans 224 90 0 0 io_in[32]
port 25 nsew signal input
flabel metal2 s 49514 19200 49570 20000 0 FreeSans 224 90 0 0 io_in[33]
port 26 nsew signal input
flabel metal2 s 50894 19200 50950 20000 0 FreeSans 224 90 0 0 io_in[34]
port 27 nsew signal input
flabel metal2 s 52274 19200 52330 20000 0 FreeSans 224 90 0 0 io_in[35]
port 28 nsew signal input
flabel metal2 s 53654 19200 53710 20000 0 FreeSans 224 90 0 0 io_in[36]
port 29 nsew signal input
flabel metal2 s 55034 19200 55090 20000 0 FreeSans 224 90 0 0 io_in[37]
port 30 nsew signal input
flabel metal2 s 8114 19200 8170 20000 0 FreeSans 224 90 0 0 io_in[3]
port 31 nsew signal input
flabel metal2 s 9494 19200 9550 20000 0 FreeSans 224 90 0 0 io_in[4]
port 32 nsew signal input
flabel metal2 s 10874 19200 10930 20000 0 FreeSans 224 90 0 0 io_in[5]
port 33 nsew signal input
flabel metal2 s 12254 19200 12310 20000 0 FreeSans 224 90 0 0 io_in[6]
port 34 nsew signal input
flabel metal2 s 13634 19200 13690 20000 0 FreeSans 224 90 0 0 io_in[7]
port 35 nsew signal input
flabel metal2 s 15014 19200 15070 20000 0 FreeSans 224 90 0 0 io_in[8]
port 36 nsew signal input
flabel metal2 s 16394 19200 16450 20000 0 FreeSans 224 90 0 0 io_in[9]
port 37 nsew signal input
flabel metal2 s 4434 19200 4490 20000 0 FreeSans 224 90 0 0 io_oeb[0]
port 38 nsew signal tristate
flabel metal2 s 18234 19200 18290 20000 0 FreeSans 224 90 0 0 io_oeb[10]
port 39 nsew signal tristate
flabel metal2 s 19614 19200 19670 20000 0 FreeSans 224 90 0 0 io_oeb[11]
port 40 nsew signal tristate
flabel metal2 s 20994 19200 21050 20000 0 FreeSans 224 90 0 0 io_oeb[12]
port 41 nsew signal tristate
flabel metal2 s 22374 19200 22430 20000 0 FreeSans 224 90 0 0 io_oeb[13]
port 42 nsew signal tristate
flabel metal2 s 23754 19200 23810 20000 0 FreeSans 224 90 0 0 io_oeb[14]
port 43 nsew signal tristate
flabel metal2 s 25134 19200 25190 20000 0 FreeSans 224 90 0 0 io_oeb[15]
port 44 nsew signal tristate
flabel metal2 s 26514 19200 26570 20000 0 FreeSans 224 90 0 0 io_oeb[16]
port 45 nsew signal tristate
flabel metal2 s 27894 19200 27950 20000 0 FreeSans 224 90 0 0 io_oeb[17]
port 46 nsew signal tristate
flabel metal2 s 29274 19200 29330 20000 0 FreeSans 224 90 0 0 io_oeb[18]
port 47 nsew signal tristate
flabel metal2 s 30654 19200 30710 20000 0 FreeSans 224 90 0 0 io_oeb[19]
port 48 nsew signal tristate
flabel metal2 s 5814 19200 5870 20000 0 FreeSans 224 90 0 0 io_oeb[1]
port 49 nsew signal tristate
flabel metal2 s 32034 19200 32090 20000 0 FreeSans 224 90 0 0 io_oeb[20]
port 50 nsew signal tristate
flabel metal2 s 33414 19200 33470 20000 0 FreeSans 224 90 0 0 io_oeb[21]
port 51 nsew signal tristate
flabel metal2 s 34794 19200 34850 20000 0 FreeSans 224 90 0 0 io_oeb[22]
port 52 nsew signal tristate
flabel metal2 s 36174 19200 36230 20000 0 FreeSans 224 90 0 0 io_oeb[23]
port 53 nsew signal tristate
flabel metal2 s 37554 19200 37610 20000 0 FreeSans 224 90 0 0 io_oeb[24]
port 54 nsew signal tristate
flabel metal2 s 38934 19200 38990 20000 0 FreeSans 224 90 0 0 io_oeb[25]
port 55 nsew signal tristate
flabel metal2 s 40314 19200 40370 20000 0 FreeSans 224 90 0 0 io_oeb[26]
port 56 nsew signal tristate
flabel metal2 s 41694 19200 41750 20000 0 FreeSans 224 90 0 0 io_oeb[27]
port 57 nsew signal tristate
flabel metal2 s 43074 19200 43130 20000 0 FreeSans 224 90 0 0 io_oeb[28]
port 58 nsew signal tristate
flabel metal2 s 44454 19200 44510 20000 0 FreeSans 224 90 0 0 io_oeb[29]
port 59 nsew signal tristate
flabel metal2 s 7194 19200 7250 20000 0 FreeSans 224 90 0 0 io_oeb[2]
port 60 nsew signal tristate
flabel metal2 s 45834 19200 45890 20000 0 FreeSans 224 90 0 0 io_oeb[30]
port 61 nsew signal tristate
flabel metal2 s 47214 19200 47270 20000 0 FreeSans 224 90 0 0 io_oeb[31]
port 62 nsew signal tristate
flabel metal2 s 48594 19200 48650 20000 0 FreeSans 224 90 0 0 io_oeb[32]
port 63 nsew signal tristate
flabel metal2 s 49974 19200 50030 20000 0 FreeSans 224 90 0 0 io_oeb[33]
port 64 nsew signal tristate
flabel metal2 s 51354 19200 51410 20000 0 FreeSans 224 90 0 0 io_oeb[34]
port 65 nsew signal tristate
flabel metal2 s 52734 19200 52790 20000 0 FreeSans 224 90 0 0 io_oeb[35]
port 66 nsew signal tristate
flabel metal2 s 54114 19200 54170 20000 0 FreeSans 224 90 0 0 io_oeb[36]
port 67 nsew signal tristate
flabel metal2 s 55494 19200 55550 20000 0 FreeSans 224 90 0 0 io_oeb[37]
port 68 nsew signal tristate
flabel metal2 s 8574 19200 8630 20000 0 FreeSans 224 90 0 0 io_oeb[3]
port 69 nsew signal tristate
flabel metal2 s 9954 19200 10010 20000 0 FreeSans 224 90 0 0 io_oeb[4]
port 70 nsew signal tristate
flabel metal2 s 11334 19200 11390 20000 0 FreeSans 224 90 0 0 io_oeb[5]
port 71 nsew signal tristate
flabel metal2 s 12714 19200 12770 20000 0 FreeSans 224 90 0 0 io_oeb[6]
port 72 nsew signal tristate
flabel metal2 s 14094 19200 14150 20000 0 FreeSans 224 90 0 0 io_oeb[7]
port 73 nsew signal tristate
flabel metal2 s 15474 19200 15530 20000 0 FreeSans 224 90 0 0 io_oeb[8]
port 74 nsew signal tristate
flabel metal2 s 16854 19200 16910 20000 0 FreeSans 224 90 0 0 io_oeb[9]
port 75 nsew signal tristate
flabel metal2 s 4894 19200 4950 20000 0 FreeSans 224 90 0 0 io_out[0]
port 76 nsew signal tristate
flabel metal2 s 18694 19200 18750 20000 0 FreeSans 224 90 0 0 io_out[10]
port 77 nsew signal tristate
flabel metal2 s 20074 19200 20130 20000 0 FreeSans 224 90 0 0 io_out[11]
port 78 nsew signal tristate
flabel metal2 s 21454 19200 21510 20000 0 FreeSans 224 90 0 0 io_out[12]
port 79 nsew signal tristate
flabel metal2 s 22834 19200 22890 20000 0 FreeSans 224 90 0 0 io_out[13]
port 80 nsew signal tristate
flabel metal2 s 24214 19200 24270 20000 0 FreeSans 224 90 0 0 io_out[14]
port 81 nsew signal tristate
flabel metal2 s 25594 19200 25650 20000 0 FreeSans 224 90 0 0 io_out[15]
port 82 nsew signal tristate
flabel metal2 s 26974 19200 27030 20000 0 FreeSans 224 90 0 0 io_out[16]
port 83 nsew signal tristate
flabel metal2 s 28354 19200 28410 20000 0 FreeSans 224 90 0 0 io_out[17]
port 84 nsew signal tristate
flabel metal2 s 29734 19200 29790 20000 0 FreeSans 224 90 0 0 io_out[18]
port 85 nsew signal tristate
flabel metal2 s 31114 19200 31170 20000 0 FreeSans 224 90 0 0 io_out[19]
port 86 nsew signal tristate
flabel metal2 s 6274 19200 6330 20000 0 FreeSans 224 90 0 0 io_out[1]
port 87 nsew signal tristate
flabel metal2 s 32494 19200 32550 20000 0 FreeSans 224 90 0 0 io_out[20]
port 88 nsew signal tristate
flabel metal2 s 33874 19200 33930 20000 0 FreeSans 224 90 0 0 io_out[21]
port 89 nsew signal tristate
flabel metal2 s 35254 19200 35310 20000 0 FreeSans 224 90 0 0 io_out[22]
port 90 nsew signal tristate
flabel metal2 s 36634 19200 36690 20000 0 FreeSans 224 90 0 0 io_out[23]
port 91 nsew signal tristate
flabel metal2 s 38014 19200 38070 20000 0 FreeSans 224 90 0 0 io_out[24]
port 92 nsew signal tristate
flabel metal2 s 39394 19200 39450 20000 0 FreeSans 224 90 0 0 io_out[25]
port 93 nsew signal tristate
flabel metal2 s 40774 19200 40830 20000 0 FreeSans 224 90 0 0 io_out[26]
port 94 nsew signal tristate
flabel metal2 s 42154 19200 42210 20000 0 FreeSans 224 90 0 0 io_out[27]
port 95 nsew signal tristate
flabel metal2 s 43534 19200 43590 20000 0 FreeSans 224 90 0 0 io_out[28]
port 96 nsew signal tristate
flabel metal2 s 44914 19200 44970 20000 0 FreeSans 224 90 0 0 io_out[29]
port 97 nsew signal tristate
flabel metal2 s 7654 19200 7710 20000 0 FreeSans 224 90 0 0 io_out[2]
port 98 nsew signal tristate
flabel metal2 s 46294 19200 46350 20000 0 FreeSans 224 90 0 0 io_out[30]
port 99 nsew signal tristate
flabel metal2 s 47674 19200 47730 20000 0 FreeSans 224 90 0 0 io_out[31]
port 100 nsew signal tristate
flabel metal2 s 49054 19200 49110 20000 0 FreeSans 224 90 0 0 io_out[32]
port 101 nsew signal tristate
flabel metal2 s 50434 19200 50490 20000 0 FreeSans 224 90 0 0 io_out[33]
port 102 nsew signal tristate
flabel metal2 s 51814 19200 51870 20000 0 FreeSans 224 90 0 0 io_out[34]
port 103 nsew signal tristate
flabel metal2 s 53194 19200 53250 20000 0 FreeSans 224 90 0 0 io_out[35]
port 104 nsew signal tristate
flabel metal2 s 54574 19200 54630 20000 0 FreeSans 224 90 0 0 io_out[36]
port 105 nsew signal tristate
flabel metal2 s 55954 19200 56010 20000 0 FreeSans 224 90 0 0 io_out[37]
port 106 nsew signal tristate
flabel metal2 s 9034 19200 9090 20000 0 FreeSans 224 90 0 0 io_out[3]
port 107 nsew signal tristate
flabel metal2 s 10414 19200 10470 20000 0 FreeSans 224 90 0 0 io_out[4]
port 108 nsew signal tristate
flabel metal2 s 11794 19200 11850 20000 0 FreeSans 224 90 0 0 io_out[5]
port 109 nsew signal tristate
flabel metal2 s 13174 19200 13230 20000 0 FreeSans 224 90 0 0 io_out[6]
port 110 nsew signal tristate
flabel metal2 s 14554 19200 14610 20000 0 FreeSans 224 90 0 0 io_out[7]
port 111 nsew signal tristate
flabel metal2 s 15934 19200 15990 20000 0 FreeSans 224 90 0 0 io_out[8]
port 112 nsew signal tristate
flabel metal2 s 17314 19200 17370 20000 0 FreeSans 224 90 0 0 io_out[9]
port 113 nsew signal tristate
flabel metal2 s 52366 0 52422 800 0 FreeSans 224 90 0 0 irq[0]
port 114 nsew signal tristate
flabel metal2 s 52458 0 52514 800 0 FreeSans 224 90 0 0 irq[1]
port 115 nsew signal tristate
flabel metal2 s 52550 0 52606 800 0 FreeSans 224 90 0 0 irq[2]
port 116 nsew signal tristate
flabel metal2 s 17038 0 17094 800 0 FreeSans 224 90 0 0 la_data_in[0]
port 117 nsew signal input
flabel metal2 s 44638 0 44694 800 0 FreeSans 224 90 0 0 la_data_in[100]
port 118 nsew signal input
flabel metal2 s 44914 0 44970 800 0 FreeSans 224 90 0 0 la_data_in[101]
port 119 nsew signal input
flabel metal2 s 45190 0 45246 800 0 FreeSans 224 90 0 0 la_data_in[102]
port 120 nsew signal input
flabel metal2 s 45466 0 45522 800 0 FreeSans 224 90 0 0 la_data_in[103]
port 121 nsew signal input
flabel metal2 s 45742 0 45798 800 0 FreeSans 224 90 0 0 la_data_in[104]
port 122 nsew signal input
flabel metal2 s 46018 0 46074 800 0 FreeSans 224 90 0 0 la_data_in[105]
port 123 nsew signal input
flabel metal2 s 46294 0 46350 800 0 FreeSans 224 90 0 0 la_data_in[106]
port 124 nsew signal input
flabel metal2 s 46570 0 46626 800 0 FreeSans 224 90 0 0 la_data_in[107]
port 125 nsew signal input
flabel metal2 s 46846 0 46902 800 0 FreeSans 224 90 0 0 la_data_in[108]
port 126 nsew signal input
flabel metal2 s 47122 0 47178 800 0 FreeSans 224 90 0 0 la_data_in[109]
port 127 nsew signal input
flabel metal2 s 19798 0 19854 800 0 FreeSans 224 90 0 0 la_data_in[10]
port 128 nsew signal input
flabel metal2 s 47398 0 47454 800 0 FreeSans 224 90 0 0 la_data_in[110]
port 129 nsew signal input
flabel metal2 s 47674 0 47730 800 0 FreeSans 224 90 0 0 la_data_in[111]
port 130 nsew signal input
flabel metal2 s 47950 0 48006 800 0 FreeSans 224 90 0 0 la_data_in[112]
port 131 nsew signal input
flabel metal2 s 48226 0 48282 800 0 FreeSans 224 90 0 0 la_data_in[113]
port 132 nsew signal input
flabel metal2 s 48502 0 48558 800 0 FreeSans 224 90 0 0 la_data_in[114]
port 133 nsew signal input
flabel metal2 s 48778 0 48834 800 0 FreeSans 224 90 0 0 la_data_in[115]
port 134 nsew signal input
flabel metal2 s 49054 0 49110 800 0 FreeSans 224 90 0 0 la_data_in[116]
port 135 nsew signal input
flabel metal2 s 49330 0 49386 800 0 FreeSans 224 90 0 0 la_data_in[117]
port 136 nsew signal input
flabel metal2 s 49606 0 49662 800 0 FreeSans 224 90 0 0 la_data_in[118]
port 137 nsew signal input
flabel metal2 s 49882 0 49938 800 0 FreeSans 224 90 0 0 la_data_in[119]
port 138 nsew signal input
flabel metal2 s 20074 0 20130 800 0 FreeSans 224 90 0 0 la_data_in[11]
port 139 nsew signal input
flabel metal2 s 50158 0 50214 800 0 FreeSans 224 90 0 0 la_data_in[120]
port 140 nsew signal input
flabel metal2 s 50434 0 50490 800 0 FreeSans 224 90 0 0 la_data_in[121]
port 141 nsew signal input
flabel metal2 s 50710 0 50766 800 0 FreeSans 224 90 0 0 la_data_in[122]
port 142 nsew signal input
flabel metal2 s 50986 0 51042 800 0 FreeSans 224 90 0 0 la_data_in[123]
port 143 nsew signal input
flabel metal2 s 51262 0 51318 800 0 FreeSans 224 90 0 0 la_data_in[124]
port 144 nsew signal input
flabel metal2 s 51538 0 51594 800 0 FreeSans 224 90 0 0 la_data_in[125]
port 145 nsew signal input
flabel metal2 s 51814 0 51870 800 0 FreeSans 224 90 0 0 la_data_in[126]
port 146 nsew signal input
flabel metal2 s 52090 0 52146 800 0 FreeSans 224 90 0 0 la_data_in[127]
port 147 nsew signal input
flabel metal2 s 20350 0 20406 800 0 FreeSans 224 90 0 0 la_data_in[12]
port 148 nsew signal input
flabel metal2 s 20626 0 20682 800 0 FreeSans 224 90 0 0 la_data_in[13]
port 149 nsew signal input
flabel metal2 s 20902 0 20958 800 0 FreeSans 224 90 0 0 la_data_in[14]
port 150 nsew signal input
flabel metal2 s 21178 0 21234 800 0 FreeSans 224 90 0 0 la_data_in[15]
port 151 nsew signal input
flabel metal2 s 21454 0 21510 800 0 FreeSans 224 90 0 0 la_data_in[16]
port 152 nsew signal input
flabel metal2 s 21730 0 21786 800 0 FreeSans 224 90 0 0 la_data_in[17]
port 153 nsew signal input
flabel metal2 s 22006 0 22062 800 0 FreeSans 224 90 0 0 la_data_in[18]
port 154 nsew signal input
flabel metal2 s 22282 0 22338 800 0 FreeSans 224 90 0 0 la_data_in[19]
port 155 nsew signal input
flabel metal2 s 17314 0 17370 800 0 FreeSans 224 90 0 0 la_data_in[1]
port 156 nsew signal input
flabel metal2 s 22558 0 22614 800 0 FreeSans 224 90 0 0 la_data_in[20]
port 157 nsew signal input
flabel metal2 s 22834 0 22890 800 0 FreeSans 224 90 0 0 la_data_in[21]
port 158 nsew signal input
flabel metal2 s 23110 0 23166 800 0 FreeSans 224 90 0 0 la_data_in[22]
port 159 nsew signal input
flabel metal2 s 23386 0 23442 800 0 FreeSans 224 90 0 0 la_data_in[23]
port 160 nsew signal input
flabel metal2 s 23662 0 23718 800 0 FreeSans 224 90 0 0 la_data_in[24]
port 161 nsew signal input
flabel metal2 s 23938 0 23994 800 0 FreeSans 224 90 0 0 la_data_in[25]
port 162 nsew signal input
flabel metal2 s 24214 0 24270 800 0 FreeSans 224 90 0 0 la_data_in[26]
port 163 nsew signal input
flabel metal2 s 24490 0 24546 800 0 FreeSans 224 90 0 0 la_data_in[27]
port 164 nsew signal input
flabel metal2 s 24766 0 24822 800 0 FreeSans 224 90 0 0 la_data_in[28]
port 165 nsew signal input
flabel metal2 s 25042 0 25098 800 0 FreeSans 224 90 0 0 la_data_in[29]
port 166 nsew signal input
flabel metal2 s 17590 0 17646 800 0 FreeSans 224 90 0 0 la_data_in[2]
port 167 nsew signal input
flabel metal2 s 25318 0 25374 800 0 FreeSans 224 90 0 0 la_data_in[30]
port 168 nsew signal input
flabel metal2 s 25594 0 25650 800 0 FreeSans 224 90 0 0 la_data_in[31]
port 169 nsew signal input
flabel metal2 s 25870 0 25926 800 0 FreeSans 224 90 0 0 la_data_in[32]
port 170 nsew signal input
flabel metal2 s 26146 0 26202 800 0 FreeSans 224 90 0 0 la_data_in[33]
port 171 nsew signal input
flabel metal2 s 26422 0 26478 800 0 FreeSans 224 90 0 0 la_data_in[34]
port 172 nsew signal input
flabel metal2 s 26698 0 26754 800 0 FreeSans 224 90 0 0 la_data_in[35]
port 173 nsew signal input
flabel metal2 s 26974 0 27030 800 0 FreeSans 224 90 0 0 la_data_in[36]
port 174 nsew signal input
flabel metal2 s 27250 0 27306 800 0 FreeSans 224 90 0 0 la_data_in[37]
port 175 nsew signal input
flabel metal2 s 27526 0 27582 800 0 FreeSans 224 90 0 0 la_data_in[38]
port 176 nsew signal input
flabel metal2 s 27802 0 27858 800 0 FreeSans 224 90 0 0 la_data_in[39]
port 177 nsew signal input
flabel metal2 s 17866 0 17922 800 0 FreeSans 224 90 0 0 la_data_in[3]
port 178 nsew signal input
flabel metal2 s 28078 0 28134 800 0 FreeSans 224 90 0 0 la_data_in[40]
port 179 nsew signal input
flabel metal2 s 28354 0 28410 800 0 FreeSans 224 90 0 0 la_data_in[41]
port 180 nsew signal input
flabel metal2 s 28630 0 28686 800 0 FreeSans 224 90 0 0 la_data_in[42]
port 181 nsew signal input
flabel metal2 s 28906 0 28962 800 0 FreeSans 224 90 0 0 la_data_in[43]
port 182 nsew signal input
flabel metal2 s 29182 0 29238 800 0 FreeSans 224 90 0 0 la_data_in[44]
port 183 nsew signal input
flabel metal2 s 29458 0 29514 800 0 FreeSans 224 90 0 0 la_data_in[45]
port 184 nsew signal input
flabel metal2 s 29734 0 29790 800 0 FreeSans 224 90 0 0 la_data_in[46]
port 185 nsew signal input
flabel metal2 s 30010 0 30066 800 0 FreeSans 224 90 0 0 la_data_in[47]
port 186 nsew signal input
flabel metal2 s 30286 0 30342 800 0 FreeSans 224 90 0 0 la_data_in[48]
port 187 nsew signal input
flabel metal2 s 30562 0 30618 800 0 FreeSans 224 90 0 0 la_data_in[49]
port 188 nsew signal input
flabel metal2 s 18142 0 18198 800 0 FreeSans 224 90 0 0 la_data_in[4]
port 189 nsew signal input
flabel metal2 s 30838 0 30894 800 0 FreeSans 224 90 0 0 la_data_in[50]
port 190 nsew signal input
flabel metal2 s 31114 0 31170 800 0 FreeSans 224 90 0 0 la_data_in[51]
port 191 nsew signal input
flabel metal2 s 31390 0 31446 800 0 FreeSans 224 90 0 0 la_data_in[52]
port 192 nsew signal input
flabel metal2 s 31666 0 31722 800 0 FreeSans 224 90 0 0 la_data_in[53]
port 193 nsew signal input
flabel metal2 s 31942 0 31998 800 0 FreeSans 224 90 0 0 la_data_in[54]
port 194 nsew signal input
flabel metal2 s 32218 0 32274 800 0 FreeSans 224 90 0 0 la_data_in[55]
port 195 nsew signal input
flabel metal2 s 32494 0 32550 800 0 FreeSans 224 90 0 0 la_data_in[56]
port 196 nsew signal input
flabel metal2 s 32770 0 32826 800 0 FreeSans 224 90 0 0 la_data_in[57]
port 197 nsew signal input
flabel metal2 s 33046 0 33102 800 0 FreeSans 224 90 0 0 la_data_in[58]
port 198 nsew signal input
flabel metal2 s 33322 0 33378 800 0 FreeSans 224 90 0 0 la_data_in[59]
port 199 nsew signal input
flabel metal2 s 18418 0 18474 800 0 FreeSans 224 90 0 0 la_data_in[5]
port 200 nsew signal input
flabel metal2 s 33598 0 33654 800 0 FreeSans 224 90 0 0 la_data_in[60]
port 201 nsew signal input
flabel metal2 s 33874 0 33930 800 0 FreeSans 224 90 0 0 la_data_in[61]
port 202 nsew signal input
flabel metal2 s 34150 0 34206 800 0 FreeSans 224 90 0 0 la_data_in[62]
port 203 nsew signal input
flabel metal2 s 34426 0 34482 800 0 FreeSans 224 90 0 0 la_data_in[63]
port 204 nsew signal input
flabel metal2 s 34702 0 34758 800 0 FreeSans 224 90 0 0 la_data_in[64]
port 205 nsew signal input
flabel metal2 s 34978 0 35034 800 0 FreeSans 224 90 0 0 la_data_in[65]
port 206 nsew signal input
flabel metal2 s 35254 0 35310 800 0 FreeSans 224 90 0 0 la_data_in[66]
port 207 nsew signal input
flabel metal2 s 35530 0 35586 800 0 FreeSans 224 90 0 0 la_data_in[67]
port 208 nsew signal input
flabel metal2 s 35806 0 35862 800 0 FreeSans 224 90 0 0 la_data_in[68]
port 209 nsew signal input
flabel metal2 s 36082 0 36138 800 0 FreeSans 224 90 0 0 la_data_in[69]
port 210 nsew signal input
flabel metal2 s 18694 0 18750 800 0 FreeSans 224 90 0 0 la_data_in[6]
port 211 nsew signal input
flabel metal2 s 36358 0 36414 800 0 FreeSans 224 90 0 0 la_data_in[70]
port 212 nsew signal input
flabel metal2 s 36634 0 36690 800 0 FreeSans 224 90 0 0 la_data_in[71]
port 213 nsew signal input
flabel metal2 s 36910 0 36966 800 0 FreeSans 224 90 0 0 la_data_in[72]
port 214 nsew signal input
flabel metal2 s 37186 0 37242 800 0 FreeSans 224 90 0 0 la_data_in[73]
port 215 nsew signal input
flabel metal2 s 37462 0 37518 800 0 FreeSans 224 90 0 0 la_data_in[74]
port 216 nsew signal input
flabel metal2 s 37738 0 37794 800 0 FreeSans 224 90 0 0 la_data_in[75]
port 217 nsew signal input
flabel metal2 s 38014 0 38070 800 0 FreeSans 224 90 0 0 la_data_in[76]
port 218 nsew signal input
flabel metal2 s 38290 0 38346 800 0 FreeSans 224 90 0 0 la_data_in[77]
port 219 nsew signal input
flabel metal2 s 38566 0 38622 800 0 FreeSans 224 90 0 0 la_data_in[78]
port 220 nsew signal input
flabel metal2 s 38842 0 38898 800 0 FreeSans 224 90 0 0 la_data_in[79]
port 221 nsew signal input
flabel metal2 s 18970 0 19026 800 0 FreeSans 224 90 0 0 la_data_in[7]
port 222 nsew signal input
flabel metal2 s 39118 0 39174 800 0 FreeSans 224 90 0 0 la_data_in[80]
port 223 nsew signal input
flabel metal2 s 39394 0 39450 800 0 FreeSans 224 90 0 0 la_data_in[81]
port 224 nsew signal input
flabel metal2 s 39670 0 39726 800 0 FreeSans 224 90 0 0 la_data_in[82]
port 225 nsew signal input
flabel metal2 s 39946 0 40002 800 0 FreeSans 224 90 0 0 la_data_in[83]
port 226 nsew signal input
flabel metal2 s 40222 0 40278 800 0 FreeSans 224 90 0 0 la_data_in[84]
port 227 nsew signal input
flabel metal2 s 40498 0 40554 800 0 FreeSans 224 90 0 0 la_data_in[85]
port 228 nsew signal input
flabel metal2 s 40774 0 40830 800 0 FreeSans 224 90 0 0 la_data_in[86]
port 229 nsew signal input
flabel metal2 s 41050 0 41106 800 0 FreeSans 224 90 0 0 la_data_in[87]
port 230 nsew signal input
flabel metal2 s 41326 0 41382 800 0 FreeSans 224 90 0 0 la_data_in[88]
port 231 nsew signal input
flabel metal2 s 41602 0 41658 800 0 FreeSans 224 90 0 0 la_data_in[89]
port 232 nsew signal input
flabel metal2 s 19246 0 19302 800 0 FreeSans 224 90 0 0 la_data_in[8]
port 233 nsew signal input
flabel metal2 s 41878 0 41934 800 0 FreeSans 224 90 0 0 la_data_in[90]
port 234 nsew signal input
flabel metal2 s 42154 0 42210 800 0 FreeSans 224 90 0 0 la_data_in[91]
port 235 nsew signal input
flabel metal2 s 42430 0 42486 800 0 FreeSans 224 90 0 0 la_data_in[92]
port 236 nsew signal input
flabel metal2 s 42706 0 42762 800 0 FreeSans 224 90 0 0 la_data_in[93]
port 237 nsew signal input
flabel metal2 s 42982 0 43038 800 0 FreeSans 224 90 0 0 la_data_in[94]
port 238 nsew signal input
flabel metal2 s 43258 0 43314 800 0 FreeSans 224 90 0 0 la_data_in[95]
port 239 nsew signal input
flabel metal2 s 43534 0 43590 800 0 FreeSans 224 90 0 0 la_data_in[96]
port 240 nsew signal input
flabel metal2 s 43810 0 43866 800 0 FreeSans 224 90 0 0 la_data_in[97]
port 241 nsew signal input
flabel metal2 s 44086 0 44142 800 0 FreeSans 224 90 0 0 la_data_in[98]
port 242 nsew signal input
flabel metal2 s 44362 0 44418 800 0 FreeSans 224 90 0 0 la_data_in[99]
port 243 nsew signal input
flabel metal2 s 19522 0 19578 800 0 FreeSans 224 90 0 0 la_data_in[9]
port 244 nsew signal input
flabel metal2 s 17130 0 17186 800 0 FreeSans 224 90 0 0 la_data_out[0]
port 245 nsew signal tristate
flabel metal2 s 44730 0 44786 800 0 FreeSans 224 90 0 0 la_data_out[100]
port 246 nsew signal tristate
flabel metal2 s 45006 0 45062 800 0 FreeSans 224 90 0 0 la_data_out[101]
port 247 nsew signal tristate
flabel metal2 s 45282 0 45338 800 0 FreeSans 224 90 0 0 la_data_out[102]
port 248 nsew signal tristate
flabel metal2 s 45558 0 45614 800 0 FreeSans 224 90 0 0 la_data_out[103]
port 249 nsew signal tristate
flabel metal2 s 45834 0 45890 800 0 FreeSans 224 90 0 0 la_data_out[104]
port 250 nsew signal tristate
flabel metal2 s 46110 0 46166 800 0 FreeSans 224 90 0 0 la_data_out[105]
port 251 nsew signal tristate
flabel metal2 s 46386 0 46442 800 0 FreeSans 224 90 0 0 la_data_out[106]
port 252 nsew signal tristate
flabel metal2 s 46662 0 46718 800 0 FreeSans 224 90 0 0 la_data_out[107]
port 253 nsew signal tristate
flabel metal2 s 46938 0 46994 800 0 FreeSans 224 90 0 0 la_data_out[108]
port 254 nsew signal tristate
flabel metal2 s 47214 0 47270 800 0 FreeSans 224 90 0 0 la_data_out[109]
port 255 nsew signal tristate
flabel metal2 s 19890 0 19946 800 0 FreeSans 224 90 0 0 la_data_out[10]
port 256 nsew signal tristate
flabel metal2 s 47490 0 47546 800 0 FreeSans 224 90 0 0 la_data_out[110]
port 257 nsew signal tristate
flabel metal2 s 47766 0 47822 800 0 FreeSans 224 90 0 0 la_data_out[111]
port 258 nsew signal tristate
flabel metal2 s 48042 0 48098 800 0 FreeSans 224 90 0 0 la_data_out[112]
port 259 nsew signal tristate
flabel metal2 s 48318 0 48374 800 0 FreeSans 224 90 0 0 la_data_out[113]
port 260 nsew signal tristate
flabel metal2 s 48594 0 48650 800 0 FreeSans 224 90 0 0 la_data_out[114]
port 261 nsew signal tristate
flabel metal2 s 48870 0 48926 800 0 FreeSans 224 90 0 0 la_data_out[115]
port 262 nsew signal tristate
flabel metal2 s 49146 0 49202 800 0 FreeSans 224 90 0 0 la_data_out[116]
port 263 nsew signal tristate
flabel metal2 s 49422 0 49478 800 0 FreeSans 224 90 0 0 la_data_out[117]
port 264 nsew signal tristate
flabel metal2 s 49698 0 49754 800 0 FreeSans 224 90 0 0 la_data_out[118]
port 265 nsew signal tristate
flabel metal2 s 49974 0 50030 800 0 FreeSans 224 90 0 0 la_data_out[119]
port 266 nsew signal tristate
flabel metal2 s 20166 0 20222 800 0 FreeSans 224 90 0 0 la_data_out[11]
port 267 nsew signal tristate
flabel metal2 s 50250 0 50306 800 0 FreeSans 224 90 0 0 la_data_out[120]
port 268 nsew signal tristate
flabel metal2 s 50526 0 50582 800 0 FreeSans 224 90 0 0 la_data_out[121]
port 269 nsew signal tristate
flabel metal2 s 50802 0 50858 800 0 FreeSans 224 90 0 0 la_data_out[122]
port 270 nsew signal tristate
flabel metal2 s 51078 0 51134 800 0 FreeSans 224 90 0 0 la_data_out[123]
port 271 nsew signal tristate
flabel metal2 s 51354 0 51410 800 0 FreeSans 224 90 0 0 la_data_out[124]
port 272 nsew signal tristate
flabel metal2 s 51630 0 51686 800 0 FreeSans 224 90 0 0 la_data_out[125]
port 273 nsew signal tristate
flabel metal2 s 51906 0 51962 800 0 FreeSans 224 90 0 0 la_data_out[126]
port 274 nsew signal tristate
flabel metal2 s 52182 0 52238 800 0 FreeSans 224 90 0 0 la_data_out[127]
port 275 nsew signal tristate
flabel metal2 s 20442 0 20498 800 0 FreeSans 224 90 0 0 la_data_out[12]
port 276 nsew signal tristate
flabel metal2 s 20718 0 20774 800 0 FreeSans 224 90 0 0 la_data_out[13]
port 277 nsew signal tristate
flabel metal2 s 20994 0 21050 800 0 FreeSans 224 90 0 0 la_data_out[14]
port 278 nsew signal tristate
flabel metal2 s 21270 0 21326 800 0 FreeSans 224 90 0 0 la_data_out[15]
port 279 nsew signal tristate
flabel metal2 s 21546 0 21602 800 0 FreeSans 224 90 0 0 la_data_out[16]
port 280 nsew signal tristate
flabel metal2 s 21822 0 21878 800 0 FreeSans 224 90 0 0 la_data_out[17]
port 281 nsew signal tristate
flabel metal2 s 22098 0 22154 800 0 FreeSans 224 90 0 0 la_data_out[18]
port 282 nsew signal tristate
flabel metal2 s 22374 0 22430 800 0 FreeSans 224 90 0 0 la_data_out[19]
port 283 nsew signal tristate
flabel metal2 s 17406 0 17462 800 0 FreeSans 224 90 0 0 la_data_out[1]
port 284 nsew signal tristate
flabel metal2 s 22650 0 22706 800 0 FreeSans 224 90 0 0 la_data_out[20]
port 285 nsew signal tristate
flabel metal2 s 22926 0 22982 800 0 FreeSans 224 90 0 0 la_data_out[21]
port 286 nsew signal tristate
flabel metal2 s 23202 0 23258 800 0 FreeSans 224 90 0 0 la_data_out[22]
port 287 nsew signal tristate
flabel metal2 s 23478 0 23534 800 0 FreeSans 224 90 0 0 la_data_out[23]
port 288 nsew signal tristate
flabel metal2 s 23754 0 23810 800 0 FreeSans 224 90 0 0 la_data_out[24]
port 289 nsew signal tristate
flabel metal2 s 24030 0 24086 800 0 FreeSans 224 90 0 0 la_data_out[25]
port 290 nsew signal tristate
flabel metal2 s 24306 0 24362 800 0 FreeSans 224 90 0 0 la_data_out[26]
port 291 nsew signal tristate
flabel metal2 s 24582 0 24638 800 0 FreeSans 224 90 0 0 la_data_out[27]
port 292 nsew signal tristate
flabel metal2 s 24858 0 24914 800 0 FreeSans 224 90 0 0 la_data_out[28]
port 293 nsew signal tristate
flabel metal2 s 25134 0 25190 800 0 FreeSans 224 90 0 0 la_data_out[29]
port 294 nsew signal tristate
flabel metal2 s 17682 0 17738 800 0 FreeSans 224 90 0 0 la_data_out[2]
port 295 nsew signal tristate
flabel metal2 s 25410 0 25466 800 0 FreeSans 224 90 0 0 la_data_out[30]
port 296 nsew signal tristate
flabel metal2 s 25686 0 25742 800 0 FreeSans 224 90 0 0 la_data_out[31]
port 297 nsew signal tristate
flabel metal2 s 25962 0 26018 800 0 FreeSans 224 90 0 0 la_data_out[32]
port 298 nsew signal tristate
flabel metal2 s 26238 0 26294 800 0 FreeSans 224 90 0 0 la_data_out[33]
port 299 nsew signal tristate
flabel metal2 s 26514 0 26570 800 0 FreeSans 224 90 0 0 la_data_out[34]
port 300 nsew signal tristate
flabel metal2 s 26790 0 26846 800 0 FreeSans 224 90 0 0 la_data_out[35]
port 301 nsew signal tristate
flabel metal2 s 27066 0 27122 800 0 FreeSans 224 90 0 0 la_data_out[36]
port 302 nsew signal tristate
flabel metal2 s 27342 0 27398 800 0 FreeSans 224 90 0 0 la_data_out[37]
port 303 nsew signal tristate
flabel metal2 s 27618 0 27674 800 0 FreeSans 224 90 0 0 la_data_out[38]
port 304 nsew signal tristate
flabel metal2 s 27894 0 27950 800 0 FreeSans 224 90 0 0 la_data_out[39]
port 305 nsew signal tristate
flabel metal2 s 17958 0 18014 800 0 FreeSans 224 90 0 0 la_data_out[3]
port 306 nsew signal tristate
flabel metal2 s 28170 0 28226 800 0 FreeSans 224 90 0 0 la_data_out[40]
port 307 nsew signal tristate
flabel metal2 s 28446 0 28502 800 0 FreeSans 224 90 0 0 la_data_out[41]
port 308 nsew signal tristate
flabel metal2 s 28722 0 28778 800 0 FreeSans 224 90 0 0 la_data_out[42]
port 309 nsew signal tristate
flabel metal2 s 28998 0 29054 800 0 FreeSans 224 90 0 0 la_data_out[43]
port 310 nsew signal tristate
flabel metal2 s 29274 0 29330 800 0 FreeSans 224 90 0 0 la_data_out[44]
port 311 nsew signal tristate
flabel metal2 s 29550 0 29606 800 0 FreeSans 224 90 0 0 la_data_out[45]
port 312 nsew signal tristate
flabel metal2 s 29826 0 29882 800 0 FreeSans 224 90 0 0 la_data_out[46]
port 313 nsew signal tristate
flabel metal2 s 30102 0 30158 800 0 FreeSans 224 90 0 0 la_data_out[47]
port 314 nsew signal tristate
flabel metal2 s 30378 0 30434 800 0 FreeSans 224 90 0 0 la_data_out[48]
port 315 nsew signal tristate
flabel metal2 s 30654 0 30710 800 0 FreeSans 224 90 0 0 la_data_out[49]
port 316 nsew signal tristate
flabel metal2 s 18234 0 18290 800 0 FreeSans 224 90 0 0 la_data_out[4]
port 317 nsew signal tristate
flabel metal2 s 30930 0 30986 800 0 FreeSans 224 90 0 0 la_data_out[50]
port 318 nsew signal tristate
flabel metal2 s 31206 0 31262 800 0 FreeSans 224 90 0 0 la_data_out[51]
port 319 nsew signal tristate
flabel metal2 s 31482 0 31538 800 0 FreeSans 224 90 0 0 la_data_out[52]
port 320 nsew signal tristate
flabel metal2 s 31758 0 31814 800 0 FreeSans 224 90 0 0 la_data_out[53]
port 321 nsew signal tristate
flabel metal2 s 32034 0 32090 800 0 FreeSans 224 90 0 0 la_data_out[54]
port 322 nsew signal tristate
flabel metal2 s 32310 0 32366 800 0 FreeSans 224 90 0 0 la_data_out[55]
port 323 nsew signal tristate
flabel metal2 s 32586 0 32642 800 0 FreeSans 224 90 0 0 la_data_out[56]
port 324 nsew signal tristate
flabel metal2 s 32862 0 32918 800 0 FreeSans 224 90 0 0 la_data_out[57]
port 325 nsew signal tristate
flabel metal2 s 33138 0 33194 800 0 FreeSans 224 90 0 0 la_data_out[58]
port 326 nsew signal tristate
flabel metal2 s 33414 0 33470 800 0 FreeSans 224 90 0 0 la_data_out[59]
port 327 nsew signal tristate
flabel metal2 s 18510 0 18566 800 0 FreeSans 224 90 0 0 la_data_out[5]
port 328 nsew signal tristate
flabel metal2 s 33690 0 33746 800 0 FreeSans 224 90 0 0 la_data_out[60]
port 329 nsew signal tristate
flabel metal2 s 33966 0 34022 800 0 FreeSans 224 90 0 0 la_data_out[61]
port 330 nsew signal tristate
flabel metal2 s 34242 0 34298 800 0 FreeSans 224 90 0 0 la_data_out[62]
port 331 nsew signal tristate
flabel metal2 s 34518 0 34574 800 0 FreeSans 224 90 0 0 la_data_out[63]
port 332 nsew signal tristate
flabel metal2 s 34794 0 34850 800 0 FreeSans 224 90 0 0 la_data_out[64]
port 333 nsew signal tristate
flabel metal2 s 35070 0 35126 800 0 FreeSans 224 90 0 0 la_data_out[65]
port 334 nsew signal tristate
flabel metal2 s 35346 0 35402 800 0 FreeSans 224 90 0 0 la_data_out[66]
port 335 nsew signal tristate
flabel metal2 s 35622 0 35678 800 0 FreeSans 224 90 0 0 la_data_out[67]
port 336 nsew signal tristate
flabel metal2 s 35898 0 35954 800 0 FreeSans 224 90 0 0 la_data_out[68]
port 337 nsew signal tristate
flabel metal2 s 36174 0 36230 800 0 FreeSans 224 90 0 0 la_data_out[69]
port 338 nsew signal tristate
flabel metal2 s 18786 0 18842 800 0 FreeSans 224 90 0 0 la_data_out[6]
port 339 nsew signal tristate
flabel metal2 s 36450 0 36506 800 0 FreeSans 224 90 0 0 la_data_out[70]
port 340 nsew signal tristate
flabel metal2 s 36726 0 36782 800 0 FreeSans 224 90 0 0 la_data_out[71]
port 341 nsew signal tristate
flabel metal2 s 37002 0 37058 800 0 FreeSans 224 90 0 0 la_data_out[72]
port 342 nsew signal tristate
flabel metal2 s 37278 0 37334 800 0 FreeSans 224 90 0 0 la_data_out[73]
port 343 nsew signal tristate
flabel metal2 s 37554 0 37610 800 0 FreeSans 224 90 0 0 la_data_out[74]
port 344 nsew signal tristate
flabel metal2 s 37830 0 37886 800 0 FreeSans 224 90 0 0 la_data_out[75]
port 345 nsew signal tristate
flabel metal2 s 38106 0 38162 800 0 FreeSans 224 90 0 0 la_data_out[76]
port 346 nsew signal tristate
flabel metal2 s 38382 0 38438 800 0 FreeSans 224 90 0 0 la_data_out[77]
port 347 nsew signal tristate
flabel metal2 s 38658 0 38714 800 0 FreeSans 224 90 0 0 la_data_out[78]
port 348 nsew signal tristate
flabel metal2 s 38934 0 38990 800 0 FreeSans 224 90 0 0 la_data_out[79]
port 349 nsew signal tristate
flabel metal2 s 19062 0 19118 800 0 FreeSans 224 90 0 0 la_data_out[7]
port 350 nsew signal tristate
flabel metal2 s 39210 0 39266 800 0 FreeSans 224 90 0 0 la_data_out[80]
port 351 nsew signal tristate
flabel metal2 s 39486 0 39542 800 0 FreeSans 224 90 0 0 la_data_out[81]
port 352 nsew signal tristate
flabel metal2 s 39762 0 39818 800 0 FreeSans 224 90 0 0 la_data_out[82]
port 353 nsew signal tristate
flabel metal2 s 40038 0 40094 800 0 FreeSans 224 90 0 0 la_data_out[83]
port 354 nsew signal tristate
flabel metal2 s 40314 0 40370 800 0 FreeSans 224 90 0 0 la_data_out[84]
port 355 nsew signal tristate
flabel metal2 s 40590 0 40646 800 0 FreeSans 224 90 0 0 la_data_out[85]
port 356 nsew signal tristate
flabel metal2 s 40866 0 40922 800 0 FreeSans 224 90 0 0 la_data_out[86]
port 357 nsew signal tristate
flabel metal2 s 41142 0 41198 800 0 FreeSans 224 90 0 0 la_data_out[87]
port 358 nsew signal tristate
flabel metal2 s 41418 0 41474 800 0 FreeSans 224 90 0 0 la_data_out[88]
port 359 nsew signal tristate
flabel metal2 s 41694 0 41750 800 0 FreeSans 224 90 0 0 la_data_out[89]
port 360 nsew signal tristate
flabel metal2 s 19338 0 19394 800 0 FreeSans 224 90 0 0 la_data_out[8]
port 361 nsew signal tristate
flabel metal2 s 41970 0 42026 800 0 FreeSans 224 90 0 0 la_data_out[90]
port 362 nsew signal tristate
flabel metal2 s 42246 0 42302 800 0 FreeSans 224 90 0 0 la_data_out[91]
port 363 nsew signal tristate
flabel metal2 s 42522 0 42578 800 0 FreeSans 224 90 0 0 la_data_out[92]
port 364 nsew signal tristate
flabel metal2 s 42798 0 42854 800 0 FreeSans 224 90 0 0 la_data_out[93]
port 365 nsew signal tristate
flabel metal2 s 43074 0 43130 800 0 FreeSans 224 90 0 0 la_data_out[94]
port 366 nsew signal tristate
flabel metal2 s 43350 0 43406 800 0 FreeSans 224 90 0 0 la_data_out[95]
port 367 nsew signal tristate
flabel metal2 s 43626 0 43682 800 0 FreeSans 224 90 0 0 la_data_out[96]
port 368 nsew signal tristate
flabel metal2 s 43902 0 43958 800 0 FreeSans 224 90 0 0 la_data_out[97]
port 369 nsew signal tristate
flabel metal2 s 44178 0 44234 800 0 FreeSans 224 90 0 0 la_data_out[98]
port 370 nsew signal tristate
flabel metal2 s 44454 0 44510 800 0 FreeSans 224 90 0 0 la_data_out[99]
port 371 nsew signal tristate
flabel metal2 s 19614 0 19670 800 0 FreeSans 224 90 0 0 la_data_out[9]
port 372 nsew signal tristate
flabel metal2 s 17222 0 17278 800 0 FreeSans 224 90 0 0 la_oenb[0]
port 373 nsew signal input
flabel metal2 s 44822 0 44878 800 0 FreeSans 224 90 0 0 la_oenb[100]
port 374 nsew signal input
flabel metal2 s 45098 0 45154 800 0 FreeSans 224 90 0 0 la_oenb[101]
port 375 nsew signal input
flabel metal2 s 45374 0 45430 800 0 FreeSans 224 90 0 0 la_oenb[102]
port 376 nsew signal input
flabel metal2 s 45650 0 45706 800 0 FreeSans 224 90 0 0 la_oenb[103]
port 377 nsew signal input
flabel metal2 s 45926 0 45982 800 0 FreeSans 224 90 0 0 la_oenb[104]
port 378 nsew signal input
flabel metal2 s 46202 0 46258 800 0 FreeSans 224 90 0 0 la_oenb[105]
port 379 nsew signal input
flabel metal2 s 46478 0 46534 800 0 FreeSans 224 90 0 0 la_oenb[106]
port 380 nsew signal input
flabel metal2 s 46754 0 46810 800 0 FreeSans 224 90 0 0 la_oenb[107]
port 381 nsew signal input
flabel metal2 s 47030 0 47086 800 0 FreeSans 224 90 0 0 la_oenb[108]
port 382 nsew signal input
flabel metal2 s 47306 0 47362 800 0 FreeSans 224 90 0 0 la_oenb[109]
port 383 nsew signal input
flabel metal2 s 19982 0 20038 800 0 FreeSans 224 90 0 0 la_oenb[10]
port 384 nsew signal input
flabel metal2 s 47582 0 47638 800 0 FreeSans 224 90 0 0 la_oenb[110]
port 385 nsew signal input
flabel metal2 s 47858 0 47914 800 0 FreeSans 224 90 0 0 la_oenb[111]
port 386 nsew signal input
flabel metal2 s 48134 0 48190 800 0 FreeSans 224 90 0 0 la_oenb[112]
port 387 nsew signal input
flabel metal2 s 48410 0 48466 800 0 FreeSans 224 90 0 0 la_oenb[113]
port 388 nsew signal input
flabel metal2 s 48686 0 48742 800 0 FreeSans 224 90 0 0 la_oenb[114]
port 389 nsew signal input
flabel metal2 s 48962 0 49018 800 0 FreeSans 224 90 0 0 la_oenb[115]
port 390 nsew signal input
flabel metal2 s 49238 0 49294 800 0 FreeSans 224 90 0 0 la_oenb[116]
port 391 nsew signal input
flabel metal2 s 49514 0 49570 800 0 FreeSans 224 90 0 0 la_oenb[117]
port 392 nsew signal input
flabel metal2 s 49790 0 49846 800 0 FreeSans 224 90 0 0 la_oenb[118]
port 393 nsew signal input
flabel metal2 s 50066 0 50122 800 0 FreeSans 224 90 0 0 la_oenb[119]
port 394 nsew signal input
flabel metal2 s 20258 0 20314 800 0 FreeSans 224 90 0 0 la_oenb[11]
port 395 nsew signal input
flabel metal2 s 50342 0 50398 800 0 FreeSans 224 90 0 0 la_oenb[120]
port 396 nsew signal input
flabel metal2 s 50618 0 50674 800 0 FreeSans 224 90 0 0 la_oenb[121]
port 397 nsew signal input
flabel metal2 s 50894 0 50950 800 0 FreeSans 224 90 0 0 la_oenb[122]
port 398 nsew signal input
flabel metal2 s 51170 0 51226 800 0 FreeSans 224 90 0 0 la_oenb[123]
port 399 nsew signal input
flabel metal2 s 51446 0 51502 800 0 FreeSans 224 90 0 0 la_oenb[124]
port 400 nsew signal input
flabel metal2 s 51722 0 51778 800 0 FreeSans 224 90 0 0 la_oenb[125]
port 401 nsew signal input
flabel metal2 s 51998 0 52054 800 0 FreeSans 224 90 0 0 la_oenb[126]
port 402 nsew signal input
flabel metal2 s 52274 0 52330 800 0 FreeSans 224 90 0 0 la_oenb[127]
port 403 nsew signal input
flabel metal2 s 20534 0 20590 800 0 FreeSans 224 90 0 0 la_oenb[12]
port 404 nsew signal input
flabel metal2 s 20810 0 20866 800 0 FreeSans 224 90 0 0 la_oenb[13]
port 405 nsew signal input
flabel metal2 s 21086 0 21142 800 0 FreeSans 224 90 0 0 la_oenb[14]
port 406 nsew signal input
flabel metal2 s 21362 0 21418 800 0 FreeSans 224 90 0 0 la_oenb[15]
port 407 nsew signal input
flabel metal2 s 21638 0 21694 800 0 FreeSans 224 90 0 0 la_oenb[16]
port 408 nsew signal input
flabel metal2 s 21914 0 21970 800 0 FreeSans 224 90 0 0 la_oenb[17]
port 409 nsew signal input
flabel metal2 s 22190 0 22246 800 0 FreeSans 224 90 0 0 la_oenb[18]
port 410 nsew signal input
flabel metal2 s 22466 0 22522 800 0 FreeSans 224 90 0 0 la_oenb[19]
port 411 nsew signal input
flabel metal2 s 17498 0 17554 800 0 FreeSans 224 90 0 0 la_oenb[1]
port 412 nsew signal input
flabel metal2 s 22742 0 22798 800 0 FreeSans 224 90 0 0 la_oenb[20]
port 413 nsew signal input
flabel metal2 s 23018 0 23074 800 0 FreeSans 224 90 0 0 la_oenb[21]
port 414 nsew signal input
flabel metal2 s 23294 0 23350 800 0 FreeSans 224 90 0 0 la_oenb[22]
port 415 nsew signal input
flabel metal2 s 23570 0 23626 800 0 FreeSans 224 90 0 0 la_oenb[23]
port 416 nsew signal input
flabel metal2 s 23846 0 23902 800 0 FreeSans 224 90 0 0 la_oenb[24]
port 417 nsew signal input
flabel metal2 s 24122 0 24178 800 0 FreeSans 224 90 0 0 la_oenb[25]
port 418 nsew signal input
flabel metal2 s 24398 0 24454 800 0 FreeSans 224 90 0 0 la_oenb[26]
port 419 nsew signal input
flabel metal2 s 24674 0 24730 800 0 FreeSans 224 90 0 0 la_oenb[27]
port 420 nsew signal input
flabel metal2 s 24950 0 25006 800 0 FreeSans 224 90 0 0 la_oenb[28]
port 421 nsew signal input
flabel metal2 s 25226 0 25282 800 0 FreeSans 224 90 0 0 la_oenb[29]
port 422 nsew signal input
flabel metal2 s 17774 0 17830 800 0 FreeSans 224 90 0 0 la_oenb[2]
port 423 nsew signal input
flabel metal2 s 25502 0 25558 800 0 FreeSans 224 90 0 0 la_oenb[30]
port 424 nsew signal input
flabel metal2 s 25778 0 25834 800 0 FreeSans 224 90 0 0 la_oenb[31]
port 425 nsew signal input
flabel metal2 s 26054 0 26110 800 0 FreeSans 224 90 0 0 la_oenb[32]
port 426 nsew signal input
flabel metal2 s 26330 0 26386 800 0 FreeSans 224 90 0 0 la_oenb[33]
port 427 nsew signal input
flabel metal2 s 26606 0 26662 800 0 FreeSans 224 90 0 0 la_oenb[34]
port 428 nsew signal input
flabel metal2 s 26882 0 26938 800 0 FreeSans 224 90 0 0 la_oenb[35]
port 429 nsew signal input
flabel metal2 s 27158 0 27214 800 0 FreeSans 224 90 0 0 la_oenb[36]
port 430 nsew signal input
flabel metal2 s 27434 0 27490 800 0 FreeSans 224 90 0 0 la_oenb[37]
port 431 nsew signal input
flabel metal2 s 27710 0 27766 800 0 FreeSans 224 90 0 0 la_oenb[38]
port 432 nsew signal input
flabel metal2 s 27986 0 28042 800 0 FreeSans 224 90 0 0 la_oenb[39]
port 433 nsew signal input
flabel metal2 s 18050 0 18106 800 0 FreeSans 224 90 0 0 la_oenb[3]
port 434 nsew signal input
flabel metal2 s 28262 0 28318 800 0 FreeSans 224 90 0 0 la_oenb[40]
port 435 nsew signal input
flabel metal2 s 28538 0 28594 800 0 FreeSans 224 90 0 0 la_oenb[41]
port 436 nsew signal input
flabel metal2 s 28814 0 28870 800 0 FreeSans 224 90 0 0 la_oenb[42]
port 437 nsew signal input
flabel metal2 s 29090 0 29146 800 0 FreeSans 224 90 0 0 la_oenb[43]
port 438 nsew signal input
flabel metal2 s 29366 0 29422 800 0 FreeSans 224 90 0 0 la_oenb[44]
port 439 nsew signal input
flabel metal2 s 29642 0 29698 800 0 FreeSans 224 90 0 0 la_oenb[45]
port 440 nsew signal input
flabel metal2 s 29918 0 29974 800 0 FreeSans 224 90 0 0 la_oenb[46]
port 441 nsew signal input
flabel metal2 s 30194 0 30250 800 0 FreeSans 224 90 0 0 la_oenb[47]
port 442 nsew signal input
flabel metal2 s 30470 0 30526 800 0 FreeSans 224 90 0 0 la_oenb[48]
port 443 nsew signal input
flabel metal2 s 30746 0 30802 800 0 FreeSans 224 90 0 0 la_oenb[49]
port 444 nsew signal input
flabel metal2 s 18326 0 18382 800 0 FreeSans 224 90 0 0 la_oenb[4]
port 445 nsew signal input
flabel metal2 s 31022 0 31078 800 0 FreeSans 224 90 0 0 la_oenb[50]
port 446 nsew signal input
flabel metal2 s 31298 0 31354 800 0 FreeSans 224 90 0 0 la_oenb[51]
port 447 nsew signal input
flabel metal2 s 31574 0 31630 800 0 FreeSans 224 90 0 0 la_oenb[52]
port 448 nsew signal input
flabel metal2 s 31850 0 31906 800 0 FreeSans 224 90 0 0 la_oenb[53]
port 449 nsew signal input
flabel metal2 s 32126 0 32182 800 0 FreeSans 224 90 0 0 la_oenb[54]
port 450 nsew signal input
flabel metal2 s 32402 0 32458 800 0 FreeSans 224 90 0 0 la_oenb[55]
port 451 nsew signal input
flabel metal2 s 32678 0 32734 800 0 FreeSans 224 90 0 0 la_oenb[56]
port 452 nsew signal input
flabel metal2 s 32954 0 33010 800 0 FreeSans 224 90 0 0 la_oenb[57]
port 453 nsew signal input
flabel metal2 s 33230 0 33286 800 0 FreeSans 224 90 0 0 la_oenb[58]
port 454 nsew signal input
flabel metal2 s 33506 0 33562 800 0 FreeSans 224 90 0 0 la_oenb[59]
port 455 nsew signal input
flabel metal2 s 18602 0 18658 800 0 FreeSans 224 90 0 0 la_oenb[5]
port 456 nsew signal input
flabel metal2 s 33782 0 33838 800 0 FreeSans 224 90 0 0 la_oenb[60]
port 457 nsew signal input
flabel metal2 s 34058 0 34114 800 0 FreeSans 224 90 0 0 la_oenb[61]
port 458 nsew signal input
flabel metal2 s 34334 0 34390 800 0 FreeSans 224 90 0 0 la_oenb[62]
port 459 nsew signal input
flabel metal2 s 34610 0 34666 800 0 FreeSans 224 90 0 0 la_oenb[63]
port 460 nsew signal input
flabel metal2 s 34886 0 34942 800 0 FreeSans 224 90 0 0 la_oenb[64]
port 461 nsew signal input
flabel metal2 s 35162 0 35218 800 0 FreeSans 224 90 0 0 la_oenb[65]
port 462 nsew signal input
flabel metal2 s 35438 0 35494 800 0 FreeSans 224 90 0 0 la_oenb[66]
port 463 nsew signal input
flabel metal2 s 35714 0 35770 800 0 FreeSans 224 90 0 0 la_oenb[67]
port 464 nsew signal input
flabel metal2 s 35990 0 36046 800 0 FreeSans 224 90 0 0 la_oenb[68]
port 465 nsew signal input
flabel metal2 s 36266 0 36322 800 0 FreeSans 224 90 0 0 la_oenb[69]
port 466 nsew signal input
flabel metal2 s 18878 0 18934 800 0 FreeSans 224 90 0 0 la_oenb[6]
port 467 nsew signal input
flabel metal2 s 36542 0 36598 800 0 FreeSans 224 90 0 0 la_oenb[70]
port 468 nsew signal input
flabel metal2 s 36818 0 36874 800 0 FreeSans 224 90 0 0 la_oenb[71]
port 469 nsew signal input
flabel metal2 s 37094 0 37150 800 0 FreeSans 224 90 0 0 la_oenb[72]
port 470 nsew signal input
flabel metal2 s 37370 0 37426 800 0 FreeSans 224 90 0 0 la_oenb[73]
port 471 nsew signal input
flabel metal2 s 37646 0 37702 800 0 FreeSans 224 90 0 0 la_oenb[74]
port 472 nsew signal input
flabel metal2 s 37922 0 37978 800 0 FreeSans 224 90 0 0 la_oenb[75]
port 473 nsew signal input
flabel metal2 s 38198 0 38254 800 0 FreeSans 224 90 0 0 la_oenb[76]
port 474 nsew signal input
flabel metal2 s 38474 0 38530 800 0 FreeSans 224 90 0 0 la_oenb[77]
port 475 nsew signal input
flabel metal2 s 38750 0 38806 800 0 FreeSans 224 90 0 0 la_oenb[78]
port 476 nsew signal input
flabel metal2 s 39026 0 39082 800 0 FreeSans 224 90 0 0 la_oenb[79]
port 477 nsew signal input
flabel metal2 s 19154 0 19210 800 0 FreeSans 224 90 0 0 la_oenb[7]
port 478 nsew signal input
flabel metal2 s 39302 0 39358 800 0 FreeSans 224 90 0 0 la_oenb[80]
port 479 nsew signal input
flabel metal2 s 39578 0 39634 800 0 FreeSans 224 90 0 0 la_oenb[81]
port 480 nsew signal input
flabel metal2 s 39854 0 39910 800 0 FreeSans 224 90 0 0 la_oenb[82]
port 481 nsew signal input
flabel metal2 s 40130 0 40186 800 0 FreeSans 224 90 0 0 la_oenb[83]
port 482 nsew signal input
flabel metal2 s 40406 0 40462 800 0 FreeSans 224 90 0 0 la_oenb[84]
port 483 nsew signal input
flabel metal2 s 40682 0 40738 800 0 FreeSans 224 90 0 0 la_oenb[85]
port 484 nsew signal input
flabel metal2 s 40958 0 41014 800 0 FreeSans 224 90 0 0 la_oenb[86]
port 485 nsew signal input
flabel metal2 s 41234 0 41290 800 0 FreeSans 224 90 0 0 la_oenb[87]
port 486 nsew signal input
flabel metal2 s 41510 0 41566 800 0 FreeSans 224 90 0 0 la_oenb[88]
port 487 nsew signal input
flabel metal2 s 41786 0 41842 800 0 FreeSans 224 90 0 0 la_oenb[89]
port 488 nsew signal input
flabel metal2 s 19430 0 19486 800 0 FreeSans 224 90 0 0 la_oenb[8]
port 489 nsew signal input
flabel metal2 s 42062 0 42118 800 0 FreeSans 224 90 0 0 la_oenb[90]
port 490 nsew signal input
flabel metal2 s 42338 0 42394 800 0 FreeSans 224 90 0 0 la_oenb[91]
port 491 nsew signal input
flabel metal2 s 42614 0 42670 800 0 FreeSans 224 90 0 0 la_oenb[92]
port 492 nsew signal input
flabel metal2 s 42890 0 42946 800 0 FreeSans 224 90 0 0 la_oenb[93]
port 493 nsew signal input
flabel metal2 s 43166 0 43222 800 0 FreeSans 224 90 0 0 la_oenb[94]
port 494 nsew signal input
flabel metal2 s 43442 0 43498 800 0 FreeSans 224 90 0 0 la_oenb[95]
port 495 nsew signal input
flabel metal2 s 43718 0 43774 800 0 FreeSans 224 90 0 0 la_oenb[96]
port 496 nsew signal input
flabel metal2 s 43994 0 44050 800 0 FreeSans 224 90 0 0 la_oenb[97]
port 497 nsew signal input
flabel metal2 s 44270 0 44326 800 0 FreeSans 224 90 0 0 la_oenb[98]
port 498 nsew signal input
flabel metal2 s 44546 0 44602 800 0 FreeSans 224 90 0 0 la_oenb[99]
port 499 nsew signal input
flabel metal2 s 19706 0 19762 800 0 FreeSans 224 90 0 0 la_oenb[9]
port 500 nsew signal input
flabel metal4 s 8168 2128 8488 17456 0 FreeSans 1920 90 0 0 vccd1
port 501 nsew power bidirectional
flabel metal4 s 22616 2128 22936 17456 0 FreeSans 1920 90 0 0 vccd1
port 501 nsew power bidirectional
flabel metal4 s 37064 2128 37384 17456 0 FreeSans 1920 90 0 0 vccd1
port 501 nsew power bidirectional
flabel metal4 s 51512 2128 51832 17456 0 FreeSans 1920 90 0 0 vccd1
port 501 nsew power bidirectional
flabel metal4 s 15392 2128 15712 17456 0 FreeSans 1920 90 0 0 vssd1
port 502 nsew ground bidirectional
flabel metal4 s 29840 2128 30160 17456 0 FreeSans 1920 90 0 0 vssd1
port 502 nsew ground bidirectional
flabel metal4 s 44288 2128 44608 17456 0 FreeSans 1920 90 0 0 vssd1
port 502 nsew ground bidirectional
flabel metal2 s 7286 0 7342 800 0 FreeSans 224 90 0 0 wb_clk_i
port 503 nsew signal input
flabel metal2 s 7378 0 7434 800 0 FreeSans 224 90 0 0 wb_rst_i
port 504 nsew signal input
flabel metal2 s 7470 0 7526 800 0 FreeSans 224 90 0 0 wbs_ack_o
port 505 nsew signal tristate
flabel metal2 s 7838 0 7894 800 0 FreeSans 224 90 0 0 wbs_adr_i[0]
port 506 nsew signal input
flabel metal2 s 10966 0 11022 800 0 FreeSans 224 90 0 0 wbs_adr_i[10]
port 507 nsew signal input
flabel metal2 s 11242 0 11298 800 0 FreeSans 224 90 0 0 wbs_adr_i[11]
port 508 nsew signal input
flabel metal2 s 11518 0 11574 800 0 FreeSans 224 90 0 0 wbs_adr_i[12]
port 509 nsew signal input
flabel metal2 s 11794 0 11850 800 0 FreeSans 224 90 0 0 wbs_adr_i[13]
port 510 nsew signal input
flabel metal2 s 12070 0 12126 800 0 FreeSans 224 90 0 0 wbs_adr_i[14]
port 511 nsew signal input
flabel metal2 s 12346 0 12402 800 0 FreeSans 224 90 0 0 wbs_adr_i[15]
port 512 nsew signal input
flabel metal2 s 12622 0 12678 800 0 FreeSans 224 90 0 0 wbs_adr_i[16]
port 513 nsew signal input
flabel metal2 s 12898 0 12954 800 0 FreeSans 224 90 0 0 wbs_adr_i[17]
port 514 nsew signal input
flabel metal2 s 13174 0 13230 800 0 FreeSans 224 90 0 0 wbs_adr_i[18]
port 515 nsew signal input
flabel metal2 s 13450 0 13506 800 0 FreeSans 224 90 0 0 wbs_adr_i[19]
port 516 nsew signal input
flabel metal2 s 8206 0 8262 800 0 FreeSans 224 90 0 0 wbs_adr_i[1]
port 517 nsew signal input
flabel metal2 s 13726 0 13782 800 0 FreeSans 224 90 0 0 wbs_adr_i[20]
port 518 nsew signal input
flabel metal2 s 14002 0 14058 800 0 FreeSans 224 90 0 0 wbs_adr_i[21]
port 519 nsew signal input
flabel metal2 s 14278 0 14334 800 0 FreeSans 224 90 0 0 wbs_adr_i[22]
port 520 nsew signal input
flabel metal2 s 14554 0 14610 800 0 FreeSans 224 90 0 0 wbs_adr_i[23]
port 521 nsew signal input
flabel metal2 s 14830 0 14886 800 0 FreeSans 224 90 0 0 wbs_adr_i[24]
port 522 nsew signal input
flabel metal2 s 15106 0 15162 800 0 FreeSans 224 90 0 0 wbs_adr_i[25]
port 523 nsew signal input
flabel metal2 s 15382 0 15438 800 0 FreeSans 224 90 0 0 wbs_adr_i[26]
port 524 nsew signal input
flabel metal2 s 15658 0 15714 800 0 FreeSans 224 90 0 0 wbs_adr_i[27]
port 525 nsew signal input
flabel metal2 s 15934 0 15990 800 0 FreeSans 224 90 0 0 wbs_adr_i[28]
port 526 nsew signal input
flabel metal2 s 16210 0 16266 800 0 FreeSans 224 90 0 0 wbs_adr_i[29]
port 527 nsew signal input
flabel metal2 s 8574 0 8630 800 0 FreeSans 224 90 0 0 wbs_adr_i[2]
port 528 nsew signal input
flabel metal2 s 16486 0 16542 800 0 FreeSans 224 90 0 0 wbs_adr_i[30]
port 529 nsew signal input
flabel metal2 s 16762 0 16818 800 0 FreeSans 224 90 0 0 wbs_adr_i[31]
port 530 nsew signal input
flabel metal2 s 8942 0 8998 800 0 FreeSans 224 90 0 0 wbs_adr_i[3]
port 531 nsew signal input
flabel metal2 s 9310 0 9366 800 0 FreeSans 224 90 0 0 wbs_adr_i[4]
port 532 nsew signal input
flabel metal2 s 9586 0 9642 800 0 FreeSans 224 90 0 0 wbs_adr_i[5]
port 533 nsew signal input
flabel metal2 s 9862 0 9918 800 0 FreeSans 224 90 0 0 wbs_adr_i[6]
port 534 nsew signal input
flabel metal2 s 10138 0 10194 800 0 FreeSans 224 90 0 0 wbs_adr_i[7]
port 535 nsew signal input
flabel metal2 s 10414 0 10470 800 0 FreeSans 224 90 0 0 wbs_adr_i[8]
port 536 nsew signal input
flabel metal2 s 10690 0 10746 800 0 FreeSans 224 90 0 0 wbs_adr_i[9]
port 537 nsew signal input
flabel metal2 s 7562 0 7618 800 0 FreeSans 224 90 0 0 wbs_cyc_i
port 538 nsew signal input
flabel metal2 s 7930 0 7986 800 0 FreeSans 224 90 0 0 wbs_dat_i[0]
port 539 nsew signal input
flabel metal2 s 11058 0 11114 800 0 FreeSans 224 90 0 0 wbs_dat_i[10]
port 540 nsew signal input
flabel metal2 s 11334 0 11390 800 0 FreeSans 224 90 0 0 wbs_dat_i[11]
port 541 nsew signal input
flabel metal2 s 11610 0 11666 800 0 FreeSans 224 90 0 0 wbs_dat_i[12]
port 542 nsew signal input
flabel metal2 s 11886 0 11942 800 0 FreeSans 224 90 0 0 wbs_dat_i[13]
port 543 nsew signal input
flabel metal2 s 12162 0 12218 800 0 FreeSans 224 90 0 0 wbs_dat_i[14]
port 544 nsew signal input
flabel metal2 s 12438 0 12494 800 0 FreeSans 224 90 0 0 wbs_dat_i[15]
port 545 nsew signal input
flabel metal2 s 12714 0 12770 800 0 FreeSans 224 90 0 0 wbs_dat_i[16]
port 546 nsew signal input
flabel metal2 s 12990 0 13046 800 0 FreeSans 224 90 0 0 wbs_dat_i[17]
port 547 nsew signal input
flabel metal2 s 13266 0 13322 800 0 FreeSans 224 90 0 0 wbs_dat_i[18]
port 548 nsew signal input
flabel metal2 s 13542 0 13598 800 0 FreeSans 224 90 0 0 wbs_dat_i[19]
port 549 nsew signal input
flabel metal2 s 8298 0 8354 800 0 FreeSans 224 90 0 0 wbs_dat_i[1]
port 550 nsew signal input
flabel metal2 s 13818 0 13874 800 0 FreeSans 224 90 0 0 wbs_dat_i[20]
port 551 nsew signal input
flabel metal2 s 14094 0 14150 800 0 FreeSans 224 90 0 0 wbs_dat_i[21]
port 552 nsew signal input
flabel metal2 s 14370 0 14426 800 0 FreeSans 224 90 0 0 wbs_dat_i[22]
port 553 nsew signal input
flabel metal2 s 14646 0 14702 800 0 FreeSans 224 90 0 0 wbs_dat_i[23]
port 554 nsew signal input
flabel metal2 s 14922 0 14978 800 0 FreeSans 224 90 0 0 wbs_dat_i[24]
port 555 nsew signal input
flabel metal2 s 15198 0 15254 800 0 FreeSans 224 90 0 0 wbs_dat_i[25]
port 556 nsew signal input
flabel metal2 s 15474 0 15530 800 0 FreeSans 224 90 0 0 wbs_dat_i[26]
port 557 nsew signal input
flabel metal2 s 15750 0 15806 800 0 FreeSans 224 90 0 0 wbs_dat_i[27]
port 558 nsew signal input
flabel metal2 s 16026 0 16082 800 0 FreeSans 224 90 0 0 wbs_dat_i[28]
port 559 nsew signal input
flabel metal2 s 16302 0 16358 800 0 FreeSans 224 90 0 0 wbs_dat_i[29]
port 560 nsew signal input
flabel metal2 s 8666 0 8722 800 0 FreeSans 224 90 0 0 wbs_dat_i[2]
port 561 nsew signal input
flabel metal2 s 16578 0 16634 800 0 FreeSans 224 90 0 0 wbs_dat_i[30]
port 562 nsew signal input
flabel metal2 s 16854 0 16910 800 0 FreeSans 224 90 0 0 wbs_dat_i[31]
port 563 nsew signal input
flabel metal2 s 9034 0 9090 800 0 FreeSans 224 90 0 0 wbs_dat_i[3]
port 564 nsew signal input
flabel metal2 s 9402 0 9458 800 0 FreeSans 224 90 0 0 wbs_dat_i[4]
port 565 nsew signal input
flabel metal2 s 9678 0 9734 800 0 FreeSans 224 90 0 0 wbs_dat_i[5]
port 566 nsew signal input
flabel metal2 s 9954 0 10010 800 0 FreeSans 224 90 0 0 wbs_dat_i[6]
port 567 nsew signal input
flabel metal2 s 10230 0 10286 800 0 FreeSans 224 90 0 0 wbs_dat_i[7]
port 568 nsew signal input
flabel metal2 s 10506 0 10562 800 0 FreeSans 224 90 0 0 wbs_dat_i[8]
port 569 nsew signal input
flabel metal2 s 10782 0 10838 800 0 FreeSans 224 90 0 0 wbs_dat_i[9]
port 570 nsew signal input
flabel metal2 s 8022 0 8078 800 0 FreeSans 224 90 0 0 wbs_dat_o[0]
port 571 nsew signal tristate
flabel metal2 s 11150 0 11206 800 0 FreeSans 224 90 0 0 wbs_dat_o[10]
port 572 nsew signal tristate
flabel metal2 s 11426 0 11482 800 0 FreeSans 224 90 0 0 wbs_dat_o[11]
port 573 nsew signal tristate
flabel metal2 s 11702 0 11758 800 0 FreeSans 224 90 0 0 wbs_dat_o[12]
port 574 nsew signal tristate
flabel metal2 s 11978 0 12034 800 0 FreeSans 224 90 0 0 wbs_dat_o[13]
port 575 nsew signal tristate
flabel metal2 s 12254 0 12310 800 0 FreeSans 224 90 0 0 wbs_dat_o[14]
port 576 nsew signal tristate
flabel metal2 s 12530 0 12586 800 0 FreeSans 224 90 0 0 wbs_dat_o[15]
port 577 nsew signal tristate
flabel metal2 s 12806 0 12862 800 0 FreeSans 224 90 0 0 wbs_dat_o[16]
port 578 nsew signal tristate
flabel metal2 s 13082 0 13138 800 0 FreeSans 224 90 0 0 wbs_dat_o[17]
port 579 nsew signal tristate
flabel metal2 s 13358 0 13414 800 0 FreeSans 224 90 0 0 wbs_dat_o[18]
port 580 nsew signal tristate
flabel metal2 s 13634 0 13690 800 0 FreeSans 224 90 0 0 wbs_dat_o[19]
port 581 nsew signal tristate
flabel metal2 s 8390 0 8446 800 0 FreeSans 224 90 0 0 wbs_dat_o[1]
port 582 nsew signal tristate
flabel metal2 s 13910 0 13966 800 0 FreeSans 224 90 0 0 wbs_dat_o[20]
port 583 nsew signal tristate
flabel metal2 s 14186 0 14242 800 0 FreeSans 224 90 0 0 wbs_dat_o[21]
port 584 nsew signal tristate
flabel metal2 s 14462 0 14518 800 0 FreeSans 224 90 0 0 wbs_dat_o[22]
port 585 nsew signal tristate
flabel metal2 s 14738 0 14794 800 0 FreeSans 224 90 0 0 wbs_dat_o[23]
port 586 nsew signal tristate
flabel metal2 s 15014 0 15070 800 0 FreeSans 224 90 0 0 wbs_dat_o[24]
port 587 nsew signal tristate
flabel metal2 s 15290 0 15346 800 0 FreeSans 224 90 0 0 wbs_dat_o[25]
port 588 nsew signal tristate
flabel metal2 s 15566 0 15622 800 0 FreeSans 224 90 0 0 wbs_dat_o[26]
port 589 nsew signal tristate
flabel metal2 s 15842 0 15898 800 0 FreeSans 224 90 0 0 wbs_dat_o[27]
port 590 nsew signal tristate
flabel metal2 s 16118 0 16174 800 0 FreeSans 224 90 0 0 wbs_dat_o[28]
port 591 nsew signal tristate
flabel metal2 s 16394 0 16450 800 0 FreeSans 224 90 0 0 wbs_dat_o[29]
port 592 nsew signal tristate
flabel metal2 s 8758 0 8814 800 0 FreeSans 224 90 0 0 wbs_dat_o[2]
port 593 nsew signal tristate
flabel metal2 s 16670 0 16726 800 0 FreeSans 224 90 0 0 wbs_dat_o[30]
port 594 nsew signal tristate
flabel metal2 s 16946 0 17002 800 0 FreeSans 224 90 0 0 wbs_dat_o[31]
port 595 nsew signal tristate
flabel metal2 s 9126 0 9182 800 0 FreeSans 224 90 0 0 wbs_dat_o[3]
port 596 nsew signal tristate
flabel metal2 s 9494 0 9550 800 0 FreeSans 224 90 0 0 wbs_dat_o[4]
port 597 nsew signal tristate
flabel metal2 s 9770 0 9826 800 0 FreeSans 224 90 0 0 wbs_dat_o[5]
port 598 nsew signal tristate
flabel metal2 s 10046 0 10102 800 0 FreeSans 224 90 0 0 wbs_dat_o[6]
port 599 nsew signal tristate
flabel metal2 s 10322 0 10378 800 0 FreeSans 224 90 0 0 wbs_dat_o[7]
port 600 nsew signal tristate
flabel metal2 s 10598 0 10654 800 0 FreeSans 224 90 0 0 wbs_dat_o[8]
port 601 nsew signal tristate
flabel metal2 s 10874 0 10930 800 0 FreeSans 224 90 0 0 wbs_dat_o[9]
port 602 nsew signal tristate
flabel metal2 s 8114 0 8170 800 0 FreeSans 224 90 0 0 wbs_sel_i[0]
port 603 nsew signal input
flabel metal2 s 8482 0 8538 800 0 FreeSans 224 90 0 0 wbs_sel_i[1]
port 604 nsew signal input
flabel metal2 s 8850 0 8906 800 0 FreeSans 224 90 0 0 wbs_sel_i[2]
port 605 nsew signal input
flabel metal2 s 9218 0 9274 800 0 FreeSans 224 90 0 0 wbs_sel_i[3]
port 606 nsew signal input
flabel metal2 s 7654 0 7710 800 0 FreeSans 224 90 0 0 wbs_stb_i
port 607 nsew signal input
flabel metal2 s 7746 0 7802 800 0 FreeSans 224 90 0 0 wbs_we_i
port 608 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 60000 20000
<< end >>
