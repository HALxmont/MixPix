magic
tech sky130B
magscale 1 2
timestamp 1667845509
<< metal1 >>
rect 71774 702992 71780 703044
rect 71832 703032 71838 703044
rect 72970 703032 72976 703044
rect 71832 703004 72976 703032
rect 71832 702992 71838 703004
rect 72970 702992 72976 703004
rect 73028 702992 73034 703044
rect 137830 700816 137836 700868
rect 137888 700856 137894 700868
rect 157334 700856 157340 700868
rect 137888 700828 157340 700856
rect 137888 700816 137894 700828
rect 157334 700816 157340 700828
rect 157392 700816 157398 700868
rect 155954 700748 155960 700800
rect 156012 700788 156018 700800
rect 202782 700788 202788 700800
rect 156012 700760 202788 700788
rect 156012 700748 156018 700760
rect 202782 700748 202788 700760
rect 202840 700748 202846 700800
rect 89162 700680 89168 700732
rect 89220 700720 89226 700732
rect 160738 700720 160744 700732
rect 89220 700692 160744 700720
rect 89220 700680 89226 700692
rect 160738 700680 160744 700692
rect 160796 700680 160802 700732
rect 154574 700612 154580 700664
rect 154632 700652 154638 700664
rect 267642 700652 267648 700664
rect 154632 700624 267648 700652
rect 154632 700612 154638 700624
rect 267642 700612 267648 700624
rect 267700 700612 267706 700664
rect 24302 700544 24308 700596
rect 24360 700584 24366 700596
rect 162210 700584 162216 700596
rect 24360 700556 162216 700584
rect 24360 700544 24366 700556
rect 162210 700544 162216 700556
rect 162268 700544 162274 700596
rect 8110 700476 8116 700528
rect 8168 700516 8174 700528
rect 162118 700516 162124 700528
rect 8168 700488 162124 700516
rect 8168 700476 8174 700488
rect 162118 700476 162124 700488
rect 162176 700476 162182 700528
rect 153286 700408 153292 700460
rect 153344 700448 153350 700460
rect 332502 700448 332508 700460
rect 153344 700420 332508 700448
rect 153344 700408 153350 700420
rect 332502 700408 332508 700420
rect 332560 700408 332566 700460
rect 153102 700340 153108 700392
rect 153160 700380 153166 700392
rect 413646 700380 413652 700392
rect 153160 700352 413652 700380
rect 153160 700340 153166 700352
rect 413646 700340 413652 700352
rect 413704 700340 413710 700392
rect 148318 700272 148324 700324
rect 148376 700312 148382 700324
rect 543458 700312 543464 700324
rect 148376 700284 543464 700312
rect 148376 700272 148382 700284
rect 543458 700272 543464 700284
rect 543516 700272 543522 700324
rect 559650 700312 559656 700324
rect 547846 700284 559656 700312
rect 542998 700204 543004 700256
rect 543056 700244 543062 700256
rect 547846 700244 547874 700284
rect 559650 700272 559656 700284
rect 559708 700272 559714 700324
rect 543056 700216 547874 700244
rect 543056 700204 543062 700216
rect 105446 699660 105452 699712
rect 105504 699700 105510 699712
rect 106918 699700 106924 699712
rect 105504 699672 106924 699700
rect 105504 699660 105510 699672
rect 106918 699660 106924 699672
rect 106976 699660 106982 699712
rect 396718 699660 396724 699712
rect 396776 699700 396782 699712
rect 397454 699700 397460 699712
rect 396776 699672 397460 699700
rect 396776 699660 396782 699672
rect 397454 699660 397460 699672
rect 397512 699660 397518 699712
rect 428458 699660 428464 699712
rect 428516 699700 428522 699712
rect 429838 699700 429844 699712
rect 428516 699672 429844 699700
rect 428516 699660 428522 699672
rect 429838 699660 429844 699672
rect 429896 699660 429902 699712
rect 146294 696940 146300 696992
rect 146352 696980 146358 696992
rect 580166 696980 580172 696992
rect 146352 696952 580172 696980
rect 146352 696940 146358 696952
rect 580166 696940 580172 696952
rect 580224 696940 580230 696992
rect 3418 683204 3424 683256
rect 3476 683244 3482 683256
rect 162302 683244 162308 683256
rect 3476 683216 162308 683244
rect 3476 683204 3482 683216
rect 162302 683204 162308 683216
rect 162360 683204 162366 683256
rect 146938 683136 146944 683188
rect 146996 683176 147002 683188
rect 580166 683176 580172 683188
rect 146996 683148 580172 683176
rect 146996 683136 147002 683148
rect 580166 683136 580172 683148
rect 580224 683136 580230 683188
rect 3510 670692 3516 670744
rect 3568 670732 3574 670744
rect 163498 670732 163504 670744
rect 3568 670704 163504 670732
rect 3568 670692 3574 670704
rect 163498 670692 163504 670704
rect 163556 670692 163562 670744
rect 185578 670692 185584 670744
rect 185636 670732 185642 670744
rect 580166 670732 580172 670744
rect 185636 670704 580172 670732
rect 185636 670692 185642 670704
rect 580166 670692 580172 670704
rect 580224 670692 580230 670744
rect 149054 660288 149060 660340
rect 149112 660328 149118 660340
rect 462314 660328 462320 660340
rect 149112 660300 462320 660328
rect 149112 660288 149118 660300
rect 462314 660288 462320 660300
rect 462372 660288 462378 660340
rect 3418 656888 3424 656940
rect 3476 656928 3482 656940
rect 163590 656928 163596 656940
rect 3476 656900 163596 656928
rect 3476 656888 3482 656900
rect 163590 656888 163596 656900
rect 163648 656888 163654 656940
rect 184198 643084 184204 643136
rect 184256 643124 184262 643136
rect 580166 643124 580172 643136
rect 184256 643096 580172 643124
rect 184256 643084 184262 643096
rect 580166 643084 580172 643096
rect 580224 643084 580230 643136
rect 3418 632068 3424 632120
rect 3476 632108 3482 632120
rect 164234 632108 164240 632120
rect 3476 632080 164240 632108
rect 3476 632068 3482 632080
rect 164234 632068 164240 632080
rect 164292 632068 164298 632120
rect 203518 630640 203524 630692
rect 203576 630680 203582 630692
rect 580166 630680 580172 630692
rect 203576 630652 580172 630680
rect 203576 630640 203582 630652
rect 580166 630640 580172 630652
rect 580224 630640 580230 630692
rect 3142 618264 3148 618316
rect 3200 618304 3206 618316
rect 164878 618304 164884 618316
rect 3200 618276 164884 618304
rect 3200 618264 3206 618276
rect 164878 618264 164884 618276
rect 164936 618264 164942 618316
rect 143626 616836 143632 616888
rect 143684 616876 143690 616888
rect 580166 616876 580172 616888
rect 143684 616848 580172 616876
rect 143684 616836 143690 616848
rect 580166 616836 580172 616848
rect 580224 616836 580230 616888
rect 3234 605820 3240 605872
rect 3292 605860 3298 605872
rect 164970 605860 164976 605872
rect 3292 605832 164976 605860
rect 3292 605820 3298 605832
rect 164970 605820 164976 605832
rect 165028 605820 165034 605872
rect 142154 590656 142160 590708
rect 142212 590696 142218 590708
rect 579798 590696 579804 590708
rect 142212 590668 579804 590696
rect 142212 590656 142218 590668
rect 579798 590656 579804 590668
rect 579856 590656 579862 590708
rect 3326 579640 3332 579692
rect 3384 579680 3390 579692
rect 165614 579680 165620 579692
rect 3384 579652 165620 579680
rect 3384 579640 3390 579652
rect 165614 579640 165620 579652
rect 165672 579640 165678 579692
rect 144178 576852 144184 576904
rect 144236 576892 144242 576904
rect 580166 576892 580172 576904
rect 144236 576864 580172 576892
rect 144236 576852 144242 576864
rect 580166 576852 580172 576864
rect 580224 576852 580230 576904
rect 3418 565836 3424 565888
rect 3476 565876 3482 565888
rect 167638 565876 167644 565888
rect 3476 565848 167644 565876
rect 3476 565836 3482 565848
rect 167638 565836 167644 565848
rect 167696 565836 167702 565888
rect 142798 563048 142804 563100
rect 142856 563088 142862 563100
rect 579798 563088 579804 563100
rect 142856 563060 579804 563088
rect 142856 563048 142862 563060
rect 579798 563048 579804 563060
rect 579856 563048 579862 563100
rect 3418 553392 3424 553444
rect 3476 553432 3482 553444
rect 166258 553432 166264 553444
rect 3476 553404 166264 553432
rect 3476 553392 3482 553404
rect 166258 553392 166264 553404
rect 166316 553392 166322 553444
rect 178678 536800 178684 536852
rect 178736 536840 178742 536852
rect 580166 536840 580172 536852
rect 178736 536812 580172 536840
rect 178736 536800 178742 536812
rect 580166 536800 580172 536812
rect 580224 536800 580230 536852
rect 3418 527144 3424 527196
rect 3476 527184 3482 527196
rect 166994 527184 167000 527196
rect 3476 527156 167000 527184
rect 3476 527144 3482 527156
rect 166994 527144 167000 527156
rect 167052 527144 167058 527196
rect 142890 524424 142896 524476
rect 142948 524464 142954 524476
rect 580166 524464 580172 524476
rect 142948 524436 580172 524464
rect 142948 524424 142954 524436
rect 580166 524424 580172 524436
rect 580224 524424 580230 524476
rect 3418 514768 3424 514820
rect 3476 514808 3482 514820
rect 8938 514808 8944 514820
rect 3476 514780 8944 514808
rect 3476 514768 3482 514780
rect 8938 514768 8944 514780
rect 8996 514768 9002 514820
rect 181438 510620 181444 510672
rect 181496 510660 181502 510672
rect 580166 510660 580172 510672
rect 181496 510632 580172 510660
rect 181496 510620 181502 510632
rect 580166 510620 580172 510632
rect 580224 510620 580230 510672
rect 3050 500964 3056 501016
rect 3108 501004 3114 501016
rect 167730 501004 167736 501016
rect 3108 500976 167736 501004
rect 3108 500964 3114 500976
rect 167730 500964 167736 500976
rect 167788 500964 167794 501016
rect 139394 484372 139400 484424
rect 139452 484412 139458 484424
rect 580166 484412 580172 484424
rect 139452 484384 580172 484412
rect 139452 484372 139458 484384
rect 580166 484372 580172 484384
rect 580224 484372 580230 484424
rect 140038 470568 140044 470620
rect 140096 470608 140102 470620
rect 579982 470608 579988 470620
rect 140096 470580 579988 470608
rect 140096 470568 140102 470580
rect 579982 470568 579988 470580
rect 580040 470568 580046 470620
rect 3510 462340 3516 462392
rect 3568 462380 3574 462392
rect 170398 462380 170404 462392
rect 3568 462352 170404 462380
rect 3568 462340 3574 462352
rect 170398 462340 170404 462352
rect 170456 462340 170462 462392
rect 180058 456764 180064 456816
rect 180116 456804 180122 456816
rect 580166 456804 580172 456816
rect 180116 456776 580172 456804
rect 180116 456764 180122 456776
rect 580166 456764 580172 456776
rect 580224 456764 580230 456816
rect 3142 448536 3148 448588
rect 3200 448576 3206 448588
rect 170490 448576 170496 448588
rect 3200 448548 170496 448576
rect 3200 448536 3206 448548
rect 170490 448536 170496 448548
rect 170548 448536 170554 448588
rect 157426 447788 157432 447840
rect 157484 447828 157490 447840
rect 169754 447828 169760 447840
rect 157484 447800 169760 447828
rect 157484 447788 157490 447800
rect 169754 447788 169760 447800
rect 169812 447788 169818 447840
rect 138658 430584 138664 430636
rect 138716 430624 138722 430636
rect 580166 430624 580172 430636
rect 138716 430596 580172 430624
rect 138716 430584 138722 430596
rect 580166 430584 580172 430596
rect 580224 430584 580230 430636
rect 3510 422288 3516 422340
rect 3568 422328 3574 422340
rect 169754 422328 169760 422340
rect 3568 422300 169760 422328
rect 3568 422288 3574 422300
rect 169754 422288 169760 422300
rect 169812 422288 169818 422340
rect 138750 418140 138756 418192
rect 138808 418180 138814 418192
rect 580166 418180 580172 418192
rect 138808 418152 580172 418180
rect 138808 418140 138814 418152
rect 580166 418140 580172 418152
rect 580224 418140 580230 418192
rect 2866 409844 2872 409896
rect 2924 409884 2930 409896
rect 171778 409884 171784 409896
rect 2924 409856 171784 409884
rect 2924 409844 2930 409856
rect 171778 409844 171784 409856
rect 171836 409844 171842 409896
rect 199378 404336 199384 404388
rect 199436 404376 199442 404388
rect 580166 404376 580172 404388
rect 199436 404348 580172 404376
rect 199436 404336 199442 404348
rect 580166 404336 580172 404348
rect 580224 404336 580230 404388
rect 3510 397468 3516 397520
rect 3568 397508 3574 397520
rect 171134 397508 171140 397520
rect 3568 397480 171140 397508
rect 3568 397468 3574 397480
rect 171134 397468 171140 397480
rect 171192 397468 171198 397520
rect 182818 378156 182824 378208
rect 182876 378196 182882 378208
rect 580166 378196 580172 378208
rect 182876 378168 580172 378196
rect 182876 378156 182882 378168
rect 580166 378156 580172 378168
rect 580224 378156 580230 378208
rect 2774 371288 2780 371340
rect 2832 371328 2838 371340
rect 4798 371328 4804 371340
rect 2832 371300 4804 371328
rect 2832 371288 2838 371300
rect 4798 371288 4804 371300
rect 4856 371288 4862 371340
rect 3142 357416 3148 357468
rect 3200 357456 3206 357468
rect 10318 357456 10324 357468
rect 3200 357428 10324 357456
rect 3200 357416 3206 357428
rect 10318 357416 10324 357428
rect 10376 357416 10382 357468
rect 135254 351908 135260 351960
rect 135312 351948 135318 351960
rect 580166 351948 580172 351960
rect 135312 351920 580172 351948
rect 135312 351908 135318 351920
rect 580166 351908 580172 351920
rect 580224 351908 580230 351960
rect 3510 345176 3516 345228
rect 3568 345216 3574 345228
rect 7558 345216 7564 345228
rect 3568 345188 7564 345216
rect 3568 345176 3574 345188
rect 7558 345176 7564 345188
rect 7616 345176 7622 345228
rect 134518 324300 134524 324352
rect 134576 324340 134582 324352
rect 580166 324340 580172 324352
rect 134576 324312 580172 324340
rect 134576 324300 134582 324312
rect 580166 324300 580172 324312
rect 580224 324300 580230 324352
rect 3326 318792 3332 318844
rect 3384 318832 3390 318844
rect 173894 318832 173900 318844
rect 3384 318804 173900 318832
rect 3384 318792 3390 318804
rect 173894 318792 173900 318804
rect 173952 318792 173958 318844
rect 135898 311856 135904 311908
rect 135956 311896 135962 311908
rect 579982 311896 579988 311908
rect 135956 311868 579988 311896
rect 135956 311856 135962 311868
rect 579982 311856 579988 311868
rect 580040 311856 580046 311908
rect 3510 304988 3516 305040
rect 3568 305028 3574 305040
rect 175918 305028 175924 305040
rect 3568 305000 175924 305028
rect 3568 304988 3574 305000
rect 175918 304988 175924 305000
rect 175976 304988 175982 305040
rect 134610 298120 134616 298172
rect 134668 298160 134674 298172
rect 580166 298160 580172 298172
rect 134668 298132 580172 298160
rect 134668 298120 134674 298132
rect 580166 298120 580172 298132
rect 580224 298120 580230 298172
rect 3510 292544 3516 292596
rect 3568 292584 3574 292596
rect 174538 292584 174544 292596
rect 3568 292556 174544 292584
rect 3568 292544 3574 292556
rect 174538 292544 174544 292556
rect 174596 292544 174602 292596
rect 10318 289076 10324 289128
rect 10376 289116 10382 289128
rect 173158 289116 173164 289128
rect 10376 289088 173164 289116
rect 10376 289076 10382 289088
rect 173158 289076 173164 289088
rect 173216 289076 173222 289128
rect 145558 287648 145564 287700
rect 145616 287688 145622 287700
rect 203518 287688 203524 287700
rect 145616 287660 203524 287688
rect 145616 287648 145622 287660
rect 203518 287648 203524 287660
rect 203576 287648 203582 287700
rect 137278 286288 137284 286340
rect 137336 286328 137342 286340
rect 182818 286328 182824 286340
rect 137336 286300 182824 286328
rect 137336 286288 137342 286300
rect 182818 286288 182824 286300
rect 182876 286288 182882 286340
rect 186314 284928 186320 284980
rect 186372 284968 186378 284980
rect 187142 284968 187148 284980
rect 186372 284940 187148 284968
rect 186372 284928 186378 284940
rect 187142 284928 187148 284940
rect 187200 284968 187206 284980
rect 396718 284968 396724 284980
rect 187200 284940 396724 284968
rect 187200 284928 187206 284940
rect 396718 284928 396724 284940
rect 396776 284928 396782 284980
rect 150434 284316 150440 284368
rect 150492 284356 150498 284368
rect 186314 284356 186320 284368
rect 150492 284328 186320 284356
rect 150492 284316 150498 284328
rect 186314 284316 186320 284328
rect 186372 284316 186378 284368
rect 147950 283568 147956 283620
rect 148008 283608 148014 283620
rect 527174 283608 527180 283620
rect 148008 283580 527180 283608
rect 148008 283568 148014 283580
rect 527174 283568 527180 283580
rect 527232 283568 527238 283620
rect 145098 282140 145104 282192
rect 145156 282180 145162 282192
rect 184198 282180 184204 282192
rect 145156 282152 184204 282180
rect 145156 282140 145162 282152
rect 184198 282140 184204 282152
rect 184256 282140 184262 282192
rect 140774 280780 140780 280832
rect 140832 280820 140838 280832
rect 178678 280820 178684 280832
rect 140832 280792 178684 280820
rect 140832 280780 140838 280792
rect 178678 280780 178684 280792
rect 178736 280780 178742 280832
rect 40034 279420 40040 279472
rect 40092 279460 40098 279472
rect 160094 279460 160100 279472
rect 40092 279432 160100 279460
rect 40092 279420 40098 279432
rect 160094 279420 160100 279432
rect 160152 279420 160158 279472
rect 204162 276632 204168 276684
rect 204220 276672 204226 276684
rect 299474 276672 299480 276684
rect 204220 276644 299480 276672
rect 204220 276632 204226 276644
rect 299474 276632 299480 276644
rect 299532 276632 299538 276684
rect 153378 276020 153384 276072
rect 153436 276060 153442 276072
rect 203058 276060 203064 276072
rect 153436 276032 203064 276060
rect 153436 276020 153442 276032
rect 203058 276020 203064 276032
rect 203116 276060 203122 276072
rect 204162 276060 204168 276072
rect 203116 276032 204168 276060
rect 203116 276020 203122 276032
rect 204162 276020 204168 276032
rect 204220 276020 204226 276072
rect 204806 275272 204812 275324
rect 204864 275312 204870 275324
rect 364334 275312 364340 275324
rect 204864 275284 364340 275312
rect 204864 275272 204870 275284
rect 364334 275272 364340 275284
rect 364392 275272 364398 275324
rect 151814 274660 151820 274712
rect 151872 274700 151878 274712
rect 204530 274700 204536 274712
rect 151872 274672 204536 274700
rect 151872 274660 151878 274672
rect 204530 274660 204536 274672
rect 204588 274700 204594 274712
rect 204806 274700 204812 274712
rect 204588 274672 204812 274700
rect 204588 274660 204594 274672
rect 204806 274660 204812 274672
rect 204864 274660 204870 274712
rect 8938 273980 8944 274032
rect 8996 274020 9002 274032
rect 169018 274020 169024 274032
rect 8996 273992 169024 274020
rect 8996 273980 9002 273992
rect 169018 273980 169024 273992
rect 169076 273980 169082 274032
rect 151078 273912 151084 273964
rect 151136 273952 151142 273964
rect 428458 273952 428464 273964
rect 151136 273924 428464 273952
rect 151136 273912 151142 273924
rect 428458 273912 428464 273924
rect 428516 273912 428522 273964
rect 133138 271872 133144 271924
rect 133196 271912 133202 271924
rect 580166 271912 580172 271924
rect 133196 271884 580172 271912
rect 133196 271872 133202 271884
rect 580166 271872 580172 271884
rect 580224 271872 580230 271924
rect 7558 271192 7564 271244
rect 7616 271232 7622 271244
rect 173250 271232 173256 271244
rect 7616 271204 173256 271232
rect 7616 271192 7622 271204
rect 173250 271192 173256 271204
rect 173308 271192 173314 271244
rect 149146 271124 149152 271176
rect 149204 271164 149210 271176
rect 494054 271164 494060 271176
rect 149204 271136 494060 271164
rect 149204 271124 149210 271136
rect 494054 271124 494060 271136
rect 494112 271124 494118 271176
rect 71774 269764 71780 269816
rect 71832 269804 71838 269816
rect 121454 269804 121460 269816
rect 71832 269776 121460 269804
rect 71832 269764 71838 269776
rect 121454 269764 121460 269776
rect 121512 269764 121518 269816
rect 147766 269764 147772 269816
rect 147824 269804 147830 269816
rect 542998 269804 543004 269816
rect 147824 269776 543004 269804
rect 147824 269764 147830 269776
rect 542998 269764 543004 269776
rect 543056 269764 543062 269816
rect 121454 269084 121460 269136
rect 121512 269124 121518 269136
rect 122374 269124 122380 269136
rect 121512 269096 122380 269124
rect 121512 269084 121518 269096
rect 122374 269084 122380 269096
rect 122432 269124 122438 269136
rect 158714 269124 158720 269136
rect 122432 269096 158720 269124
rect 122432 269084 122438 269096
rect 158714 269084 158720 269096
rect 158772 269084 158778 269136
rect 146202 268404 146208 268456
rect 146260 268444 146266 268456
rect 185578 268444 185584 268456
rect 146260 268416 185584 268444
rect 146260 268404 146266 268416
rect 185578 268404 185584 268416
rect 185636 268404 185642 268456
rect 4798 268336 4804 268388
rect 4856 268376 4862 268388
rect 172698 268376 172704 268388
rect 4856 268348 172704 268376
rect 4856 268336 4862 268348
rect 172698 268336 172704 268348
rect 172756 268336 172762 268388
rect 137830 266976 137836 267028
rect 137888 267016 137894 267028
rect 199378 267016 199384 267028
rect 137888 266988 199384 267016
rect 137888 266976 137894 266988
rect 199378 266976 199384 266988
rect 199436 266976 199442 267028
rect 3050 266364 3056 266416
rect 3108 266404 3114 266416
rect 175918 266404 175924 266416
rect 3108 266376 175924 266404
rect 3108 266364 3114 266376
rect 175918 266364 175924 266376
rect 175976 266364 175982 266416
rect 174538 265752 174544 265804
rect 174596 265792 174602 265804
rect 174596 265764 190454 265792
rect 174596 265752 174602 265764
rect 141694 265684 141700 265736
rect 141752 265724 141758 265736
rect 181438 265724 181444 265736
rect 141752 265696 181444 265724
rect 141752 265684 141758 265696
rect 181438 265684 181444 265696
rect 181496 265684 181502 265736
rect 3418 265616 3424 265668
rect 3476 265656 3482 265668
rect 169202 265656 169208 265668
rect 3476 265628 169208 265656
rect 3476 265616 3482 265628
rect 169202 265616 169208 265628
rect 169260 265616 169266 265668
rect 190426 265656 190454 265764
rect 192018 265656 192024 265668
rect 190426 265628 192024 265656
rect 192018 265616 192024 265628
rect 192076 265616 192082 265668
rect 173250 265548 173256 265600
rect 173308 265588 173314 265600
rect 192110 265588 192116 265600
rect 173308 265560 192116 265588
rect 173308 265548 173314 265560
rect 192110 265548 192116 265560
rect 192168 265548 192174 265600
rect 175826 265480 175832 265532
rect 175884 265520 175890 265532
rect 199194 265520 199200 265532
rect 175884 265492 199200 265520
rect 175884 265480 175890 265492
rect 199194 265480 199200 265492
rect 199252 265480 199258 265532
rect 170398 265412 170404 265464
rect 170456 265452 170462 265464
rect 170674 265452 170680 265464
rect 170456 265424 170680 265452
rect 170456 265412 170462 265424
rect 170674 265412 170680 265424
rect 170732 265452 170738 265464
rect 195054 265452 195060 265464
rect 170732 265424 195060 265452
rect 170732 265412 170738 265424
rect 195054 265412 195060 265424
rect 195112 265412 195118 265464
rect 171778 265344 171784 265396
rect 171836 265384 171842 265396
rect 196618 265384 196624 265396
rect 171836 265356 196624 265384
rect 171836 265344 171842 265356
rect 196618 265344 196624 265356
rect 196676 265344 196682 265396
rect 167822 265276 167828 265328
rect 167880 265316 167886 265328
rect 193582 265316 193588 265328
rect 167880 265288 193588 265316
rect 167880 265276 167886 265288
rect 193582 265276 193588 265288
rect 193640 265276 193646 265328
rect 162302 265208 162308 265260
rect 162360 265248 162366 265260
rect 188246 265248 188252 265260
rect 162360 265220 188252 265248
rect 162360 265208 162366 265220
rect 188246 265208 188252 265220
rect 188304 265208 188310 265260
rect 169110 265140 169116 265192
rect 169168 265180 169174 265192
rect 196250 265180 196256 265192
rect 169168 265152 196256 265180
rect 169168 265140 169174 265152
rect 196250 265140 196256 265152
rect 196308 265140 196314 265192
rect 167454 265072 167460 265124
rect 167512 265112 167518 265124
rect 194962 265112 194968 265124
rect 167512 265084 194968 265112
rect 167512 265072 167518 265084
rect 194962 265072 194968 265084
rect 195020 265072 195026 265124
rect 164878 265004 164884 265056
rect 164936 265044 164942 265056
rect 165338 265044 165344 265056
rect 164936 265016 165344 265044
rect 164936 265004 164942 265016
rect 165338 265004 165344 265016
rect 165396 265044 165402 265056
rect 196434 265044 196440 265056
rect 165396 265016 196440 265044
rect 165396 265004 165402 265016
rect 196434 265004 196440 265016
rect 196492 265004 196498 265056
rect 152182 264936 152188 264988
rect 152240 264976 152246 264988
rect 153102 264976 153108 264988
rect 152240 264948 153108 264976
rect 152240 264936 152246 264948
rect 153102 264936 153108 264948
rect 153160 264976 153166 264988
rect 187510 264976 187516 264988
rect 153160 264948 187516 264976
rect 153160 264936 153166 264948
rect 187510 264936 187516 264948
rect 187568 264936 187574 264988
rect 120810 264256 120816 264308
rect 120868 264296 120874 264308
rect 139486 264296 139492 264308
rect 120868 264268 139492 264296
rect 120868 264256 120874 264268
rect 139486 264256 139492 264268
rect 139544 264296 139550 264308
rect 139544 264268 142154 264296
rect 139544 264256 139550 264268
rect 106918 264188 106924 264240
rect 106976 264228 106982 264240
rect 121454 264228 121460 264240
rect 106976 264200 121460 264228
rect 106976 264188 106982 264200
rect 121454 264188 121460 264200
rect 121512 264188 121518 264240
rect 142126 264228 142154 264268
rect 180058 264228 180064 264240
rect 142126 264200 180064 264228
rect 180058 264188 180064 264200
rect 180116 264188 180122 264240
rect 118234 264120 118240 264172
rect 118292 264160 118298 264172
rect 134242 264160 134248 264172
rect 118292 264132 134248 264160
rect 118292 264120 118298 264132
rect 134242 264120 134248 264132
rect 134300 264160 134306 264172
rect 134610 264160 134616 264172
rect 134300 264132 134616 264160
rect 134300 264120 134306 264132
rect 134610 264120 134616 264132
rect 134668 264120 134674 264172
rect 115566 264052 115572 264104
rect 115624 264092 115630 264104
rect 133138 264092 133144 264104
rect 115624 264064 133144 264092
rect 115624 264052 115630 264064
rect 133138 264052 133144 264064
rect 133196 264052 133202 264104
rect 120902 263984 120908 264036
rect 120960 264024 120966 264036
rect 141142 264024 141148 264036
rect 120960 263996 141148 264024
rect 120960 263984 120966 263996
rect 141142 263984 141148 263996
rect 141200 264024 141206 264036
rect 141694 264024 141700 264036
rect 141200 263996 141700 264024
rect 141200 263984 141206 263996
rect 141694 263984 141700 263996
rect 141752 263984 141758 264036
rect 115382 263916 115388 263968
rect 115440 263956 115446 263968
rect 137186 263956 137192 263968
rect 115440 263928 137192 263956
rect 115440 263916 115446 263928
rect 137186 263916 137192 263928
rect 137244 263916 137250 263968
rect 119798 263848 119804 263900
rect 119856 263888 119862 263900
rect 142614 263888 142620 263900
rect 119856 263860 142620 263888
rect 119856 263848 119862 263860
rect 142614 263848 142620 263860
rect 142672 263848 142678 263900
rect 122558 263780 122564 263832
rect 122616 263820 122622 263832
rect 148502 263820 148508 263832
rect 122616 263792 148508 263820
rect 122616 263780 122622 263792
rect 148502 263780 148508 263792
rect 148560 263780 148566 263832
rect 119706 263712 119712 263764
rect 119764 263752 119770 263764
rect 146202 263752 146208 263764
rect 119764 263724 146208 263752
rect 119764 263712 119770 263724
rect 146202 263712 146208 263724
rect 146260 263712 146266 263764
rect 120718 263644 120724 263696
rect 120776 263684 120782 263696
rect 151078 263684 151084 263696
rect 120776 263656 151084 263684
rect 120776 263644 120782 263656
rect 151078 263644 151084 263656
rect 151136 263644 151142 263696
rect 172698 263644 172704 263696
rect 172756 263684 172762 263696
rect 189350 263684 189356 263696
rect 172756 263656 189356 263684
rect 172756 263644 172762 263656
rect 189350 263644 189356 263656
rect 189408 263644 189414 263696
rect 121454 263576 121460 263628
rect 121512 263616 121518 263628
rect 122006 263616 122012 263628
rect 121512 263588 122012 263616
rect 121512 263576 121518 263588
rect 122006 263576 122012 263588
rect 122064 263616 122070 263628
rect 159082 263616 159088 263628
rect 122064 263588 159088 263616
rect 122064 263576 122070 263588
rect 159082 263576 159088 263588
rect 159140 263576 159146 263628
rect 173158 263576 173164 263628
rect 173216 263616 173222 263628
rect 173710 263616 173716 263628
rect 173216 263588 173716 263616
rect 173216 263576 173222 263588
rect 173710 263576 173716 263588
rect 173768 263616 173774 263628
rect 197906 263616 197912 263628
rect 173768 263588 197912 263616
rect 173768 263576 173774 263588
rect 197906 263576 197912 263588
rect 197964 263576 197970 263628
rect 137462 263508 137468 263560
rect 137520 263548 137526 263560
rect 580258 263548 580264 263560
rect 137520 263520 580264 263548
rect 137520 263508 137526 263520
rect 580258 263508 580264 263520
rect 580316 263508 580322 263560
rect 150434 263440 150440 263492
rect 150492 263480 150498 263492
rect 151354 263480 151360 263492
rect 150492 263452 151360 263480
rect 150492 263440 150498 263452
rect 151354 263440 151360 263452
rect 151412 263440 151418 263492
rect 193122 263440 193128 263492
rect 193180 263480 193186 263492
rect 218054 263480 218060 263492
rect 193180 263452 218060 263480
rect 193180 263440 193186 263452
rect 218054 263440 218060 263452
rect 218112 263440 218118 263492
rect 163406 263236 163412 263288
rect 163464 263276 163470 263288
rect 163590 263276 163596 263288
rect 163464 263248 163596 263276
rect 163464 263236 163470 263248
rect 163590 263236 163596 263248
rect 163648 263236 163654 263288
rect 170214 263032 170220 263084
rect 170272 263072 170278 263084
rect 170490 263072 170496 263084
rect 170272 263044 170496 263072
rect 170272 263032 170278 263044
rect 170490 263032 170496 263044
rect 170548 263072 170554 263084
rect 192294 263072 192300 263084
rect 170548 263044 192300 263072
rect 170548 263032 170554 263044
rect 192294 263032 192300 263044
rect 192352 263032 192358 263084
rect 116762 262964 116768 263016
rect 116820 263004 116826 263016
rect 131114 263004 131120 263016
rect 116820 262976 131120 263004
rect 116820 262964 116826 262976
rect 131114 262964 131120 262976
rect 131172 262964 131178 263016
rect 132034 262964 132040 263016
rect 132092 263004 132098 263016
rect 580350 263004 580356 263016
rect 132092 262976 580356 263004
rect 132092 262964 132098 262976
rect 580350 262964 580356 262976
rect 580408 262964 580414 263016
rect 3418 262896 3424 262948
rect 3476 262936 3482 262948
rect 178494 262936 178500 262948
rect 3476 262908 178500 262936
rect 3476 262896 3482 262908
rect 178494 262896 178500 262908
rect 178552 262896 178558 262948
rect 179230 262896 179236 262948
rect 179288 262936 179294 262948
rect 189534 262936 189540 262948
rect 179288 262908 189540 262936
rect 179288 262896 179294 262908
rect 189534 262896 189540 262908
rect 189592 262896 189598 262948
rect 113818 262828 113824 262880
rect 113876 262868 113882 262880
rect 131758 262868 131764 262880
rect 113876 262840 131764 262868
rect 113876 262828 113882 262840
rect 131758 262828 131764 262840
rect 131816 262868 131822 262880
rect 580442 262868 580448 262880
rect 131816 262840 580448 262868
rect 131816 262828 131822 262840
rect 580442 262828 580448 262840
rect 580500 262828 580506 262880
rect 113910 262760 113916 262812
rect 113968 262800 113974 262812
rect 134518 262800 134524 262812
rect 113968 262772 134524 262800
rect 113968 262760 113974 262772
rect 134518 262760 134524 262772
rect 134576 262800 134582 262812
rect 134794 262800 134800 262812
rect 134576 262772 134800 262800
rect 134576 262760 134582 262772
rect 134794 262760 134800 262772
rect 134852 262760 134858 262812
rect 163406 262760 163412 262812
rect 163464 262800 163470 262812
rect 192386 262800 192392 262812
rect 163464 262772 192392 262800
rect 163464 262760 163470 262772
rect 192386 262760 192392 262772
rect 192444 262760 192450 262812
rect 116670 262692 116676 262744
rect 116728 262732 116734 262744
rect 127710 262732 127716 262744
rect 116728 262704 127716 262732
rect 116728 262692 116734 262704
rect 127710 262692 127716 262704
rect 127768 262692 127774 262744
rect 162026 262692 162032 262744
rect 162084 262732 162090 262744
rect 193766 262732 193772 262744
rect 162084 262704 193772 262732
rect 162084 262692 162090 262704
rect 193766 262692 193772 262704
rect 193824 262692 193830 262744
rect 115290 262624 115296 262676
rect 115348 262664 115354 262676
rect 129826 262664 129832 262676
rect 115348 262636 129832 262664
rect 115348 262624 115354 262636
rect 129826 262624 129832 262636
rect 129884 262624 129890 262676
rect 153194 262624 153200 262676
rect 153252 262664 153258 262676
rect 158714 262664 158720 262676
rect 153252 262636 158720 262664
rect 153252 262624 153258 262636
rect 158714 262624 158720 262636
rect 158772 262624 158778 262676
rect 162210 262624 162216 262676
rect 162268 262664 162274 262676
rect 195146 262664 195152 262676
rect 162268 262636 195152 262664
rect 162268 262624 162274 262636
rect 195146 262624 195152 262636
rect 195204 262624 195210 262676
rect 112898 262556 112904 262608
rect 112956 262596 112962 262608
rect 128722 262596 128728 262608
rect 112956 262568 128728 262596
rect 112956 262556 112962 262568
rect 128722 262556 128728 262568
rect 128780 262556 128786 262608
rect 157150 262556 157156 262608
rect 157208 262596 157214 262608
rect 192478 262596 192484 262608
rect 157208 262568 192484 262596
rect 157208 262556 157214 262568
rect 192478 262556 192484 262568
rect 192536 262596 192542 262608
rect 193122 262596 193128 262608
rect 192536 262568 193128 262596
rect 192536 262556 192542 262568
rect 193122 262556 193128 262568
rect 193180 262556 193186 262608
rect 121914 262488 121920 262540
rect 121972 262528 121978 262540
rect 144178 262528 144184 262540
rect 121972 262500 144184 262528
rect 121972 262488 121978 262500
rect 144178 262488 144184 262500
rect 144236 262488 144242 262540
rect 160738 262488 160744 262540
rect 160796 262528 160802 262540
rect 200574 262528 200580 262540
rect 160796 262500 200580 262528
rect 160796 262488 160802 262500
rect 200574 262488 200580 262500
rect 200632 262488 200638 262540
rect 3510 262420 3516 262472
rect 3568 262460 3574 262472
rect 176746 262460 176752 262472
rect 3568 262432 176752 262460
rect 3568 262420 3574 262432
rect 176746 262420 176752 262432
rect 176804 262420 176810 262472
rect 180150 262420 180156 262472
rect 180208 262460 180214 262472
rect 193490 262460 193496 262472
rect 180208 262432 193496 262460
rect 180208 262420 180214 262432
rect 193490 262420 193496 262432
rect 193548 262420 193554 262472
rect 118142 262352 118148 262404
rect 118200 262392 118206 262404
rect 129274 262392 129280 262404
rect 118200 262364 129280 262392
rect 118200 262352 118206 262364
rect 129274 262352 129280 262364
rect 129332 262352 129338 262404
rect 182910 262352 182916 262404
rect 182968 262392 182974 262404
rect 182968 262364 190454 262392
rect 182968 262352 182974 262364
rect 190426 262336 190454 262364
rect 184566 262284 184572 262336
rect 184624 262324 184630 262336
rect 189166 262324 189172 262336
rect 184624 262296 189172 262324
rect 184624 262284 184630 262296
rect 189166 262284 189172 262296
rect 189224 262284 189230 262336
rect 190426 262296 190460 262336
rect 190454 262284 190460 262296
rect 190512 262284 190518 262336
rect 122466 262216 122472 262268
rect 122524 262256 122530 262268
rect 125962 262256 125968 262268
rect 122524 262228 125968 262256
rect 122524 262216 122530 262228
rect 125962 262216 125968 262228
rect 126020 262216 126026 262268
rect 181254 262216 181260 262268
rect 181312 262256 181318 262268
rect 187786 262256 187792 262268
rect 181312 262228 187792 262256
rect 181312 262216 181318 262228
rect 187786 262216 187792 262228
rect 187844 262216 187850 262268
rect 129826 261400 129832 261452
rect 129884 261440 129890 261452
rect 188338 261440 188344 261452
rect 129884 261412 188344 261440
rect 129884 261400 129890 261412
rect 188338 261400 188344 261412
rect 188396 261400 188402 261452
rect 176746 261332 176752 261384
rect 176804 261372 176810 261384
rect 197998 261372 198004 261384
rect 176804 261344 198004 261372
rect 176804 261332 176810 261344
rect 197998 261332 198004 261344
rect 198056 261332 198062 261384
rect 131114 261264 131120 261316
rect 131172 261304 131178 261316
rect 471238 261304 471244 261316
rect 131172 261276 471244 261304
rect 131172 261264 131178 261276
rect 471238 261264 471244 261276
rect 471296 261264 471302 261316
rect 184014 261196 184020 261248
rect 184072 261236 184078 261248
rect 199010 261236 199016 261248
rect 184072 261208 199016 261236
rect 184072 261196 184078 261208
rect 199010 261196 199016 261208
rect 199068 261196 199074 261248
rect 118050 261128 118056 261180
rect 118108 261168 118114 261180
rect 132862 261168 132868 261180
rect 118108 261140 132868 261168
rect 118108 261128 118114 261140
rect 132862 261128 132868 261140
rect 132920 261128 132926 261180
rect 180518 261128 180524 261180
rect 180576 261168 180582 261180
rect 198090 261168 198096 261180
rect 180576 261140 198096 261168
rect 180576 261128 180582 261140
rect 198090 261128 198096 261140
rect 198148 261128 198154 261180
rect 111242 261060 111248 261112
rect 111300 261100 111306 261112
rect 132034 261100 132040 261112
rect 111300 261072 132040 261100
rect 111300 261060 111306 261072
rect 132034 261060 132040 261072
rect 132092 261060 132098 261112
rect 178494 261060 178500 261112
rect 178552 261100 178558 261112
rect 199102 261100 199108 261112
rect 178552 261072 199108 261100
rect 178552 261060 178558 261072
rect 199102 261060 199108 261072
rect 199160 261060 199166 261112
rect 111426 260992 111432 261044
rect 111484 261032 111490 261044
rect 130378 261032 130384 261044
rect 111484 261004 130384 261032
rect 111484 260992 111490 261004
rect 130378 260992 130384 261004
rect 130436 260992 130442 261044
rect 181990 260992 181996 261044
rect 182048 261032 182054 261044
rect 197814 261032 197820 261044
rect 182048 261004 197820 261032
rect 182048 260992 182054 261004
rect 197814 260992 197820 261004
rect 197872 260992 197878 261044
rect 4798 260924 4804 260976
rect 4856 260964 4862 260976
rect 176194 260964 176200 260976
rect 4856 260936 176200 260964
rect 4856 260924 4862 260936
rect 176194 260924 176200 260936
rect 176252 260964 176258 260976
rect 190914 260964 190920 260976
rect 176252 260936 190920 260964
rect 176252 260924 176258 260936
rect 190914 260924 190920 260936
rect 190972 260924 190978 260976
rect 112622 260856 112628 260908
rect 112680 260896 112686 260908
rect 133966 260896 133972 260908
rect 112680 260868 133972 260896
rect 112680 260856 112686 260868
rect 133966 260856 133972 260868
rect 134024 260856 134030 260908
rect 177574 260856 177580 260908
rect 177632 260896 177638 260908
rect 191006 260896 191012 260908
rect 177632 260868 191012 260896
rect 177632 260856 177638 260868
rect 191006 260856 191012 260868
rect 191064 260856 191070 260908
rect 119338 260788 119344 260840
rect 119396 260828 119402 260840
rect 124306 260828 124312 260840
rect 119396 260800 124312 260828
rect 119396 260788 119402 260800
rect 124306 260788 124312 260800
rect 124364 260788 124370 260840
rect 173894 260380 173900 260432
rect 173952 260420 173958 260432
rect 173952 260392 180794 260420
rect 173952 260380 173958 260392
rect 180766 260352 180794 260392
rect 185578 260380 185584 260432
rect 185636 260420 185642 260432
rect 190730 260420 190736 260432
rect 185636 260392 190736 260420
rect 185636 260380 185642 260392
rect 190730 260380 190736 260392
rect 190788 260380 190794 260432
rect 187878 260352 187884 260364
rect 180766 260324 187884 260352
rect 187878 260312 187884 260324
rect 187936 260312 187942 260364
rect 167702 260256 171134 260284
rect 167702 260228 167730 260256
rect 116578 260176 116584 260228
rect 116636 260216 116642 260228
rect 135254 260216 135260 260228
rect 116636 260188 135260 260216
rect 116636 260176 116642 260188
rect 135254 260176 135260 260188
rect 135312 260216 135318 260228
rect 136220 260216 136226 260228
rect 135312 260188 136226 260216
rect 135312 260176 135318 260188
rect 136220 260176 136226 260188
rect 136278 260176 136284 260228
rect 157334 260176 157340 260228
rect 157392 260216 157398 260228
rect 158300 260216 158306 260228
rect 157392 260188 158306 260216
rect 157392 260176 157398 260188
rect 158300 260176 158306 260188
rect 158358 260176 158364 260228
rect 166994 260176 167000 260228
rect 167052 260216 167058 260228
rect 167684 260216 167690 260228
rect 167052 260188 167690 260216
rect 167052 260176 167058 260188
rect 167684 260176 167690 260188
rect 167742 260176 167748 260228
rect 169754 260176 169760 260228
rect 169812 260216 169818 260228
rect 170996 260216 171002 260228
rect 169812 260188 171002 260216
rect 169812 260176 169818 260188
rect 170996 260176 171002 260188
rect 171054 260176 171060 260228
rect 171106 260216 171134 260256
rect 175918 260244 175924 260296
rect 175976 260284 175982 260296
rect 175976 260256 176240 260284
rect 175976 260244 175982 260256
rect 176102 260216 176108 260228
rect 171106 260188 176108 260216
rect 176102 260176 176108 260188
rect 176160 260176 176166 260228
rect 176212 260216 176240 260256
rect 178402 260244 178408 260296
rect 178460 260284 178466 260296
rect 189626 260284 189632 260296
rect 178460 260256 189632 260284
rect 178460 260244 178466 260256
rect 189626 260244 189632 260256
rect 189684 260244 189690 260296
rect 187326 260216 187332 260228
rect 176212 260188 187332 260216
rect 187326 260176 187332 260188
rect 187384 260176 187390 260228
rect 132908 260108 132914 260160
rect 132966 260148 132972 260160
rect 485038 260148 485044 260160
rect 132966 260120 485044 260148
rect 132966 260108 132972 260120
rect 485038 260108 485044 260120
rect 485096 260108 485102 260160
rect 114002 260040 114008 260092
rect 114060 260080 114066 260092
rect 126836 260080 126842 260092
rect 114060 260052 126842 260080
rect 114060 260040 114066 260052
rect 126836 260040 126842 260052
rect 126894 260040 126900 260092
rect 170996 260040 171002 260092
rect 171054 260080 171060 260092
rect 185578 260080 185584 260092
rect 171054 260052 185584 260080
rect 171054 260040 171060 260052
rect 185578 260040 185584 260052
rect 185636 260040 185642 260092
rect 185670 260040 185676 260092
rect 185728 260080 185734 260092
rect 190822 260080 190828 260092
rect 185728 260052 190828 260080
rect 185728 260040 185734 260052
rect 190822 260040 190828 260052
rect 190880 260040 190886 260092
rect 113634 259972 113640 260024
rect 113692 260012 113698 260024
rect 128354 260012 128360 260024
rect 113692 259984 128360 260012
rect 113692 259972 113698 259984
rect 128354 259972 128360 259984
rect 128412 259972 128418 260024
rect 189442 260012 189448 260024
rect 171612 259984 189448 260012
rect 117866 259904 117872 259956
rect 117924 259944 117930 259956
rect 142154 259944 142160 259956
rect 117924 259916 142160 259944
rect 117924 259904 117930 259916
rect 142154 259904 142160 259916
rect 142212 259944 142218 259956
rect 143074 259944 143080 259956
rect 142212 259916 143080 259944
rect 142212 259904 142218 259916
rect 143074 259904 143080 259916
rect 143132 259904 143138 259956
rect 119430 259836 119436 259888
rect 119488 259876 119494 259888
rect 146294 259876 146300 259888
rect 119488 259848 146300 259876
rect 119488 259836 119494 259848
rect 146294 259836 146300 259848
rect 146352 259836 146358 259888
rect 169478 259836 169484 259888
rect 169536 259876 169542 259888
rect 171612 259876 171640 259984
rect 189442 259972 189448 259984
rect 189500 259972 189506 260024
rect 171686 259904 171692 259956
rect 171744 259944 171750 259956
rect 193674 259944 193680 259956
rect 171744 259916 188108 259944
rect 171744 259904 171750 259916
rect 169536 259848 171640 259876
rect 169536 259836 169542 259848
rect 176102 259836 176108 259888
rect 176160 259876 176166 259888
rect 185670 259876 185676 259888
rect 176160 259848 185676 259876
rect 176160 259836 176166 259848
rect 185670 259836 185676 259848
rect 185728 259836 185734 259888
rect 119522 259768 119528 259820
rect 119580 259808 119586 259820
rect 149146 259808 149152 259820
rect 119580 259780 149152 259808
rect 119580 259768 119586 259780
rect 149146 259768 149152 259780
rect 149204 259768 149210 259820
rect 158070 259768 158076 259820
rect 158128 259808 158134 259820
rect 187970 259808 187976 259820
rect 158128 259780 187976 259808
rect 158128 259768 158134 259780
rect 187970 259768 187976 259780
rect 188028 259768 188034 259820
rect 188080 259808 188108 259916
rect 190426 259916 193680 259944
rect 190426 259808 190454 259916
rect 193674 259904 193680 259916
rect 193732 259904 193738 259956
rect 188080 259780 190454 259808
rect 119614 259700 119620 259752
rect 119672 259740 119678 259752
rect 153194 259740 153200 259752
rect 119672 259712 153200 259740
rect 119672 259700 119678 259712
rect 153194 259700 153200 259712
rect 153252 259700 153258 259752
rect 158622 259700 158628 259752
rect 158680 259740 158686 259752
rect 188154 259740 188160 259752
rect 158680 259712 188160 259740
rect 158680 259700 158686 259712
rect 188154 259700 188160 259712
rect 188212 259700 188218 259752
rect 134334 259632 134340 259684
rect 134392 259672 134398 259684
rect 187694 259672 187700 259684
rect 134392 259644 187700 259672
rect 134392 259632 134398 259644
rect 187694 259632 187700 259644
rect 187752 259632 187758 259684
rect 120534 259564 120540 259616
rect 120592 259604 120598 259616
rect 178034 259604 178040 259616
rect 120592 259576 178040 259604
rect 120592 259564 120598 259576
rect 178034 259564 178040 259576
rect 178092 259564 178098 259616
rect 181806 259564 181812 259616
rect 181864 259604 181870 259616
rect 203426 259604 203432 259616
rect 181864 259576 203432 259604
rect 181864 259564 181870 259576
rect 203426 259564 203432 259576
rect 203484 259564 203490 259616
rect 7558 259496 7564 259548
rect 7616 259536 7622 259548
rect 177298 259536 177304 259548
rect 7616 259508 177304 259536
rect 7616 259496 7622 259508
rect 177298 259496 177304 259508
rect 177356 259496 177362 259548
rect 183462 259496 183468 259548
rect 183520 259536 183526 259548
rect 206094 259536 206100 259548
rect 183520 259508 206100 259536
rect 183520 259496 183526 259508
rect 206094 259496 206100 259508
rect 206152 259496 206158 259548
rect 117958 259428 117964 259480
rect 118016 259468 118022 259480
rect 139394 259468 139400 259480
rect 118016 259440 139400 259468
rect 118016 259428 118022 259440
rect 139394 259428 139400 259440
rect 139452 259468 139458 259480
rect 139762 259468 139768 259480
rect 139452 259440 139768 259468
rect 139452 259428 139458 259440
rect 139762 259428 139768 259440
rect 139820 259428 139826 259480
rect 184934 259428 184940 259480
rect 184992 259468 184998 259480
rect 196526 259468 196532 259480
rect 184992 259440 196532 259468
rect 184992 259428 184998 259440
rect 196526 259428 196532 259440
rect 196584 259428 196590 259480
rect 187694 259360 187700 259412
rect 187752 259400 187758 259412
rect 580166 259400 580172 259412
rect 187752 259372 580172 259400
rect 187752 259360 187758 259372
rect 580166 259360 580172 259372
rect 580224 259360 580230 259412
rect 187786 258476 187792 258528
rect 187844 258516 187850 258528
rect 188062 258516 188068 258528
rect 187844 258488 188068 258516
rect 187844 258476 187850 258488
rect 188062 258476 188068 258488
rect 188120 258476 188126 258528
rect 485038 245556 485044 245608
rect 485096 245596 485102 245608
rect 580166 245596 580172 245608
rect 485096 245568 580172 245596
rect 485096 245556 485102 245568
rect 580166 245556 580172 245568
rect 580224 245556 580230 245608
rect 2774 241204 2780 241256
rect 2832 241244 2838 241256
rect 4798 241244 4804 241256
rect 2832 241216 4804 241244
rect 2832 241204 2838 241216
rect 4798 241204 4804 241216
rect 4856 241204 4862 241256
rect 3510 215092 3516 215144
rect 3568 215132 3574 215144
rect 7558 215132 7564 215144
rect 3568 215104 7564 215132
rect 3568 215092 3574 215104
rect 7558 215092 7564 215104
rect 7616 215092 7622 215144
rect 471238 206932 471244 206984
rect 471296 206972 471302 206984
rect 579798 206972 579804 206984
rect 471296 206944 579804 206972
rect 471296 206932 471302 206944
rect 579798 206932 579804 206944
rect 579856 206932 579862 206984
rect 142126 201096 147168 201124
rect 124186 200960 128354 200988
rect 124186 200716 124214 200960
rect 122806 200688 124214 200716
rect 128326 200716 128354 200960
rect 142126 200920 142154 201096
rect 132328 200892 142154 200920
rect 132328 200852 132356 200892
rect 132144 200824 132356 200852
rect 142126 200824 147076 200852
rect 132144 200728 132172 200824
rect 142126 200784 142154 200824
rect 132236 200756 142154 200784
rect 132236 200728 132264 200756
rect 130838 200716 130844 200728
rect 128326 200688 130844 200716
rect 104434 200540 104440 200592
rect 104492 200580 104498 200592
rect 122806 200580 122834 200688
rect 130838 200676 130844 200688
rect 130896 200676 130902 200728
rect 132034 200716 132040 200728
rect 131040 200688 132040 200716
rect 104492 200552 122834 200580
rect 104492 200540 104498 200552
rect 119062 200472 119068 200524
rect 119120 200512 119126 200524
rect 131040 200512 131068 200688
rect 132034 200676 132040 200688
rect 132092 200676 132098 200728
rect 132126 200676 132132 200728
rect 132184 200676 132190 200728
rect 132218 200676 132224 200728
rect 132276 200676 132282 200728
rect 132328 200688 139394 200716
rect 131114 200608 131120 200660
rect 131172 200648 131178 200660
rect 132328 200648 132356 200688
rect 131172 200620 132356 200648
rect 131172 200608 131178 200620
rect 132034 200540 132040 200592
rect 132092 200580 132098 200592
rect 132218 200580 132224 200592
rect 132092 200552 132224 200580
rect 132092 200540 132098 200552
rect 132218 200540 132224 200552
rect 132276 200540 132282 200592
rect 119120 200484 131068 200512
rect 139366 200512 139394 200688
rect 139366 200484 145236 200512
rect 119120 200472 119126 200484
rect 113082 200404 113088 200456
rect 113140 200444 113146 200456
rect 113140 200416 143074 200444
rect 113140 200404 113146 200416
rect 112990 200336 112996 200388
rect 113048 200376 113054 200388
rect 113048 200348 141188 200376
rect 113048 200336 113054 200348
rect 119890 200268 119896 200320
rect 119948 200308 119954 200320
rect 132126 200308 132132 200320
rect 119948 200280 132132 200308
rect 119948 200268 119954 200280
rect 132126 200268 132132 200280
rect 132184 200268 132190 200320
rect 118602 200200 118608 200252
rect 118660 200240 118666 200252
rect 141160 200240 141188 200348
rect 118660 200212 139394 200240
rect 141160 200212 142982 200240
rect 118660 200200 118666 200212
rect 130838 200064 130844 200116
rect 130896 200104 130902 200116
rect 130896 200076 138290 200104
rect 130896 200064 130902 200076
rect 124186 200008 135806 200036
rect 102870 199656 102876 199708
rect 102928 199696 102934 199708
rect 124186 199696 124214 200008
rect 102928 199668 124214 199696
rect 125980 199940 135668 199968
rect 102928 199656 102934 199668
rect 105998 199588 106004 199640
rect 106056 199628 106062 199640
rect 125980 199628 126008 199940
rect 132908 199860 132914 199912
rect 132966 199860 132972 199912
rect 133000 199860 133006 199912
rect 133058 199860 133064 199912
rect 133276 199900 133282 199912
rect 133110 199872 133282 199900
rect 126054 199724 126060 199776
rect 126112 199764 126118 199776
rect 132926 199764 132954 199860
rect 126112 199736 132954 199764
rect 126112 199724 126118 199736
rect 130746 199656 130752 199708
rect 130804 199696 130810 199708
rect 133018 199696 133046 199860
rect 130804 199668 133046 199696
rect 130804 199656 130810 199668
rect 106056 199600 126008 199628
rect 106056 199588 106062 199600
rect 130654 199588 130660 199640
rect 130712 199628 130718 199640
rect 133110 199628 133138 199872
rect 133276 199860 133282 199872
rect 133334 199860 133340 199912
rect 133460 199860 133466 199912
rect 133518 199860 133524 199912
rect 133644 199860 133650 199912
rect 133702 199860 133708 199912
rect 133736 199860 133742 199912
rect 133794 199860 133800 199912
rect 133920 199860 133926 199912
rect 133978 199860 133984 199912
rect 134196 199860 134202 199912
rect 134254 199860 134260 199912
rect 134472 199860 134478 199912
rect 134530 199860 134536 199912
rect 134748 199860 134754 199912
rect 134806 199860 134812 199912
rect 135024 199860 135030 199912
rect 135082 199860 135088 199912
rect 135116 199860 135122 199912
rect 135174 199860 135180 199912
rect 135208 199860 135214 199912
rect 135266 199860 135272 199912
rect 135300 199860 135306 199912
rect 135358 199860 135364 199912
rect 135392 199860 135398 199912
rect 135450 199860 135456 199912
rect 133478 199640 133506 199860
rect 133662 199776 133690 199860
rect 133644 199724 133650 199776
rect 133702 199724 133708 199776
rect 133754 199708 133782 199860
rect 133938 199776 133966 199860
rect 134012 199792 134018 199844
rect 134070 199792 134076 199844
rect 133874 199724 133880 199776
rect 133932 199736 133966 199776
rect 133932 199724 133938 199736
rect 133754 199668 133788 199708
rect 133782 199656 133788 199668
rect 133840 199656 133846 199708
rect 130712 199600 133138 199628
rect 130712 199588 130718 199600
rect 133414 199588 133420 199640
rect 133472 199600 133506 199640
rect 133472 199588 133478 199600
rect 133598 199588 133604 199640
rect 133656 199628 133662 199640
rect 134030 199628 134058 199792
rect 134214 199708 134242 199860
rect 134490 199708 134518 199860
rect 134150 199656 134156 199708
rect 134208 199668 134242 199708
rect 134208 199656 134214 199668
rect 134426 199656 134432 199708
rect 134484 199668 134518 199708
rect 134766 199708 134794 199860
rect 135042 199832 135070 199860
rect 134996 199804 135070 199832
rect 134766 199668 134800 199708
rect 134484 199656 134490 199668
rect 134794 199656 134800 199668
rect 134852 199656 134858 199708
rect 134996 199640 135024 199804
rect 135134 199776 135162 199860
rect 135070 199724 135076 199776
rect 135128 199736 135162 199776
rect 135128 199724 135134 199736
rect 135226 199640 135254 199860
rect 135318 199640 135346 199860
rect 135410 199640 135438 199860
rect 135640 199832 135668 199940
rect 135778 199912 135806 200008
rect 135870 199940 137462 199968
rect 135760 199860 135766 199912
rect 135818 199860 135824 199912
rect 135870 199832 135898 199940
rect 136036 199860 136042 199912
rect 136094 199860 136100 199912
rect 136128 199860 136134 199912
rect 136186 199900 136192 199912
rect 136588 199900 136594 199912
rect 136186 199872 136450 199900
rect 136186 199860 136192 199872
rect 135640 199804 135898 199832
rect 136054 199832 136082 199860
rect 136054 199804 136128 199832
rect 136100 199776 136128 199804
rect 136312 199792 136318 199844
rect 136370 199792 136376 199844
rect 135484 199724 135490 199776
rect 135542 199724 135548 199776
rect 136082 199724 136088 199776
rect 136140 199724 136146 199776
rect 135502 199696 135530 199724
rect 136330 199696 136358 199792
rect 135502 199668 136358 199696
rect 133656 199600 134058 199628
rect 133656 199588 133662 199600
rect 134978 199588 134984 199640
rect 135036 199588 135042 199640
rect 135162 199588 135168 199640
rect 135220 199600 135254 199640
rect 135220 199588 135226 199600
rect 135300 199588 135306 199640
rect 135358 199588 135364 199640
rect 135410 199600 135444 199640
rect 135438 199588 135444 199600
rect 135496 199588 135502 199640
rect 136174 199588 136180 199640
rect 136232 199628 136238 199640
rect 136422 199628 136450 199872
rect 136560 199860 136594 199900
rect 136646 199860 136652 199912
rect 136680 199860 136686 199912
rect 136738 199860 136744 199912
rect 136772 199860 136778 199912
rect 136830 199860 136836 199912
rect 137232 199860 137238 199912
rect 137290 199860 137296 199912
rect 137324 199860 137330 199912
rect 137382 199860 137388 199912
rect 136560 199640 136588 199860
rect 136698 199832 136726 199860
rect 136652 199804 136726 199832
rect 136652 199708 136680 199804
rect 136790 199776 136818 199860
rect 136726 199724 136732 199776
rect 136784 199736 136818 199776
rect 136784 199724 136790 199736
rect 136634 199656 136640 199708
rect 136692 199656 136698 199708
rect 137250 199640 137278 199860
rect 136232 199600 136450 199628
rect 136232 199588 136238 199600
rect 136542 199588 136548 199640
rect 136600 199588 136606 199640
rect 137186 199588 137192 199640
rect 137244 199600 137278 199640
rect 137244 199588 137250 199600
rect 137342 199572 137370 199860
rect 114922 199520 114928 199572
rect 114980 199560 114986 199572
rect 132954 199560 132960 199572
rect 114980 199532 132960 199560
rect 114980 199520 114986 199532
rect 132954 199520 132960 199532
rect 133012 199520 133018 199572
rect 133690 199520 133696 199572
rect 133748 199560 133754 199572
rect 136818 199560 136824 199572
rect 133748 199532 136824 199560
rect 133748 199520 133754 199532
rect 136818 199520 136824 199532
rect 136876 199520 136882 199572
rect 137278 199520 137284 199572
rect 137336 199532 137370 199572
rect 137434 199560 137462 199940
rect 138262 199912 138290 200076
rect 139366 200036 139394 200212
rect 139366 200008 141970 200036
rect 141942 199968 141970 200008
rect 139044 199940 139394 199968
rect 137784 199860 137790 199912
rect 137842 199860 137848 199912
rect 137876 199860 137882 199912
rect 137934 199860 137940 199912
rect 137968 199860 137974 199912
rect 138026 199860 138032 199912
rect 138060 199860 138066 199912
rect 138118 199900 138124 199912
rect 138118 199860 138152 199900
rect 138244 199860 138250 199912
rect 138302 199860 138308 199912
rect 138520 199860 138526 199912
rect 138578 199860 138584 199912
rect 138704 199900 138710 199912
rect 138630 199872 138710 199900
rect 137508 199792 137514 199844
rect 137566 199792 137572 199844
rect 137600 199792 137606 199844
rect 137658 199792 137664 199844
rect 137526 199640 137554 199792
rect 137618 199696 137646 199792
rect 137618 199668 137692 199696
rect 137664 199640 137692 199668
rect 137802 199640 137830 199860
rect 137894 199776 137922 199860
rect 137986 199832 138014 199860
rect 137986 199804 138060 199832
rect 138032 199776 138060 199804
rect 137894 199736 137928 199776
rect 137922 199724 137928 199736
rect 137980 199724 137986 199776
rect 138014 199724 138020 199776
rect 138072 199724 138078 199776
rect 138124 199640 138152 199860
rect 138428 199792 138434 199844
rect 138486 199792 138492 199844
rect 138446 199696 138474 199792
rect 138400 199668 138474 199696
rect 137526 199600 137560 199640
rect 137554 199588 137560 199600
rect 137612 199588 137618 199640
rect 137646 199588 137652 199640
rect 137704 199588 137710 199640
rect 137738 199588 137744 199640
rect 137796 199600 137830 199640
rect 137796 199588 137802 199600
rect 138106 199588 138112 199640
rect 138164 199588 138170 199640
rect 138400 199572 138428 199668
rect 138538 199640 138566 199860
rect 138474 199588 138480 199640
rect 138532 199600 138566 199640
rect 138532 199588 138538 199600
rect 138630 199572 138658 199872
rect 138704 199860 138710 199872
rect 138762 199860 138768 199912
rect 138796 199860 138802 199912
rect 138854 199860 138860 199912
rect 138888 199860 138894 199912
rect 138946 199860 138952 199912
rect 138814 199776 138842 199860
rect 138750 199724 138756 199776
rect 138808 199736 138842 199776
rect 138808 199724 138814 199736
rect 138906 199708 138934 199860
rect 138842 199656 138848 199708
rect 138900 199668 138934 199708
rect 138900 199656 138906 199668
rect 139044 199640 139072 199940
rect 139366 199912 139394 199940
rect 139458 199940 139946 199968
rect 139164 199860 139170 199912
rect 139222 199860 139228 199912
rect 139348 199860 139354 199912
rect 139406 199860 139412 199912
rect 139026 199588 139032 199640
rect 139084 199588 139090 199640
rect 139182 199628 139210 199860
rect 139302 199628 139308 199640
rect 139182 199600 139308 199628
rect 139302 199588 139308 199600
rect 139360 199588 139366 199640
rect 137830 199560 137836 199572
rect 137434 199532 137836 199560
rect 137336 199520 137342 199532
rect 137830 199520 137836 199532
rect 137888 199520 137894 199572
rect 138382 199520 138388 199572
rect 138440 199520 138446 199572
rect 138630 199532 138664 199572
rect 138658 199520 138664 199532
rect 138716 199520 138722 199572
rect 138750 199520 138756 199572
rect 138808 199560 138814 199572
rect 139458 199560 139486 199940
rect 139918 199912 139946 199940
rect 140654 199940 141326 199968
rect 139532 199860 139538 199912
rect 139590 199860 139596 199912
rect 139716 199860 139722 199912
rect 139774 199860 139780 199912
rect 139808 199860 139814 199912
rect 139866 199860 139872 199912
rect 139900 199860 139906 199912
rect 139958 199860 139964 199912
rect 139992 199860 139998 199912
rect 140050 199860 140056 199912
rect 140176 199860 140182 199912
rect 140234 199860 140240 199912
rect 140360 199860 140366 199912
rect 140418 199860 140424 199912
rect 140452 199860 140458 199912
rect 140510 199860 140516 199912
rect 139550 199708 139578 199860
rect 139734 199776 139762 199860
rect 139670 199724 139676 199776
rect 139728 199736 139762 199776
rect 139826 199776 139854 199860
rect 140010 199776 140038 199860
rect 139826 199736 139860 199776
rect 139728 199724 139734 199736
rect 139854 199724 139860 199736
rect 139912 199724 139918 199776
rect 139946 199724 139952 199776
rect 140004 199736 140038 199776
rect 140004 199724 140010 199736
rect 139550 199668 139584 199708
rect 139578 199656 139584 199668
rect 139636 199656 139642 199708
rect 140038 199588 140044 199640
rect 140096 199628 140102 199640
rect 140194 199628 140222 199860
rect 140378 199832 140406 199860
rect 140096 199600 140222 199628
rect 140332 199804 140406 199832
rect 140096 199588 140102 199600
rect 138808 199532 139486 199560
rect 138808 199520 138814 199532
rect 140222 199520 140228 199572
rect 140280 199560 140286 199572
rect 140332 199560 140360 199804
rect 140470 199776 140498 199860
rect 140406 199724 140412 199776
rect 140464 199736 140498 199776
rect 140464 199724 140470 199736
rect 140654 199628 140682 199940
rect 141298 199912 141326 199940
rect 141390 199940 141878 199968
rect 141942 199940 142154 199968
rect 140728 199860 140734 199912
rect 140786 199860 140792 199912
rect 140820 199860 140826 199912
rect 140878 199900 140884 199912
rect 140878 199860 140912 199900
rect 141004 199860 141010 199912
rect 141062 199860 141068 199912
rect 141280 199860 141286 199912
rect 141338 199860 141344 199912
rect 140746 199776 140774 199860
rect 140728 199724 140734 199776
rect 140786 199724 140792 199776
rect 140884 199708 140912 199860
rect 141022 199832 141050 199860
rect 141390 199832 141418 199940
rect 141464 199860 141470 199912
rect 141522 199860 141528 199912
rect 141740 199860 141746 199912
rect 141798 199860 141804 199912
rect 141022 199804 141418 199832
rect 141482 199708 141510 199860
rect 140866 199656 140872 199708
rect 140924 199656 140930 199708
rect 141418 199656 141424 199708
rect 141476 199668 141510 199708
rect 141476 199656 141482 199668
rect 141602 199628 141608 199640
rect 140654 199600 141608 199628
rect 141602 199588 141608 199600
rect 141660 199588 141666 199640
rect 141758 199572 141786 199860
rect 141850 199640 141878 199940
rect 142016 199860 142022 199912
rect 142074 199860 142080 199912
rect 141924 199792 141930 199844
rect 141982 199792 141988 199844
rect 141942 199696 141970 199792
rect 142034 199764 142062 199860
rect 142126 199832 142154 199940
rect 142678 199940 142890 199968
rect 142678 199912 142706 199940
rect 142200 199860 142206 199912
rect 142258 199900 142264 199912
rect 142258 199872 142522 199900
rect 142258 199860 142264 199872
rect 142126 199804 142384 199832
rect 142034 199736 142292 199764
rect 142154 199696 142160 199708
rect 141942 199668 142160 199696
rect 142154 199656 142160 199668
rect 142212 199656 142218 199708
rect 141850 199600 141884 199640
rect 141878 199588 141884 199600
rect 141936 199588 141942 199640
rect 141970 199588 141976 199640
rect 142028 199628 142034 199640
rect 142028 199600 142154 199628
rect 142028 199588 142034 199600
rect 140280 199532 140360 199560
rect 140280 199520 140286 199532
rect 141142 199520 141148 199572
rect 141200 199560 141206 199572
rect 141510 199560 141516 199572
rect 141200 199532 141516 199560
rect 141200 199520 141206 199532
rect 141510 199520 141516 199532
rect 141568 199520 141574 199572
rect 141758 199532 141792 199572
rect 141786 199520 141792 199532
rect 141844 199520 141850 199572
rect 142126 199560 142154 199600
rect 142264 199560 142292 199736
rect 142356 199628 142384 199804
rect 142494 199776 142522 199872
rect 142568 199860 142574 199912
rect 142626 199860 142632 199912
rect 142660 199860 142666 199912
rect 142718 199860 142724 199912
rect 142752 199860 142758 199912
rect 142810 199860 142816 199912
rect 142476 199724 142482 199776
rect 142534 199724 142540 199776
rect 142586 199696 142614 199860
rect 142586 199668 142660 199696
rect 142522 199628 142528 199640
rect 142356 199600 142528 199628
rect 142522 199588 142528 199600
rect 142580 199588 142586 199640
rect 142632 199572 142660 199668
rect 142770 199640 142798 199860
rect 142862 199832 142890 199940
rect 142954 199912 142982 200212
rect 142936 199860 142942 199912
rect 142994 199860 143000 199912
rect 143046 199832 143074 200416
rect 145208 199968 145236 200484
rect 147048 200036 147076 200824
rect 147140 200172 147168 201096
rect 154546 201096 184244 201124
rect 154546 200784 154574 201096
rect 153902 200756 154574 200784
rect 158686 200756 167684 200784
rect 147140 200144 151814 200172
rect 147048 200008 148778 200036
rect 143552 199940 144454 199968
rect 145208 199940 145282 199968
rect 143120 199860 143126 199912
rect 143178 199860 143184 199912
rect 142862 199804 143074 199832
rect 143138 199764 143166 199860
rect 143212 199792 143218 199844
rect 143270 199792 143276 199844
rect 143304 199792 143310 199844
rect 143362 199792 143368 199844
rect 143396 199792 143402 199844
rect 143454 199832 143460 199844
rect 143454 199792 143488 199832
rect 143092 199736 143166 199764
rect 143092 199708 143120 199736
rect 143230 199708 143258 199792
rect 143074 199656 143080 199708
rect 143132 199656 143138 199708
rect 143166 199656 143172 199708
rect 143224 199668 143258 199708
rect 143224 199656 143230 199668
rect 143322 199640 143350 199792
rect 143460 199640 143488 199792
rect 143552 199640 143580 199940
rect 144426 199912 144454 199940
rect 143672 199860 143678 199912
rect 143730 199860 143736 199912
rect 143764 199860 143770 199912
rect 143822 199860 143828 199912
rect 144040 199860 144046 199912
rect 144098 199860 144104 199912
rect 144132 199860 144138 199912
rect 144190 199860 144196 199912
rect 144408 199860 144414 199912
rect 144466 199860 144472 199912
rect 144500 199860 144506 199912
rect 144558 199860 144564 199912
rect 144592 199860 144598 199912
rect 144650 199860 144656 199912
rect 145052 199860 145058 199912
rect 145110 199860 145116 199912
rect 145144 199860 145150 199912
rect 145202 199860 145208 199912
rect 143690 199640 143718 199860
rect 143782 199776 143810 199860
rect 143782 199736 143816 199776
rect 143810 199724 143816 199736
rect 143868 199724 143874 199776
rect 142706 199588 142712 199640
rect 142764 199600 142798 199640
rect 142764 199588 142770 199600
rect 143258 199588 143264 199640
rect 143316 199600 143350 199640
rect 143316 199588 143322 199600
rect 143442 199588 143448 199640
rect 143500 199588 143506 199640
rect 143534 199588 143540 199640
rect 143592 199588 143598 199640
rect 143690 199600 143724 199640
rect 143718 199588 143724 199600
rect 143776 199588 143782 199640
rect 142126 199532 142292 199560
rect 142614 199520 142620 199572
rect 142672 199520 142678 199572
rect 143350 199520 143356 199572
rect 143408 199560 143414 199572
rect 143408 199532 143488 199560
rect 143408 199520 143414 199532
rect 118326 199452 118332 199504
rect 118384 199492 118390 199504
rect 142430 199492 142436 199504
rect 118384 199464 142436 199492
rect 118384 199452 118390 199464
rect 142430 199452 142436 199464
rect 142488 199452 142494 199504
rect 122466 199384 122472 199436
rect 122524 199424 122530 199436
rect 126606 199424 126612 199436
rect 122524 199396 126612 199424
rect 122524 199384 122530 199396
rect 126606 199384 126612 199396
rect 126664 199384 126670 199436
rect 127894 199384 127900 199436
rect 127952 199424 127958 199436
rect 135162 199424 135168 199436
rect 127952 199396 135168 199424
rect 127952 199384 127958 199396
rect 135162 199384 135168 199396
rect 135220 199384 135226 199436
rect 143350 199424 143356 199436
rect 135824 199396 143356 199424
rect 135824 199368 135852 199396
rect 143350 199384 143356 199396
rect 143408 199384 143414 199436
rect 143460 199424 143488 199532
rect 143902 199520 143908 199572
rect 143960 199560 143966 199572
rect 144058 199560 144086 199860
rect 143960 199532 144086 199560
rect 144150 199572 144178 199860
rect 144518 199708 144546 199860
rect 144454 199656 144460 199708
rect 144512 199668 144546 199708
rect 144512 199656 144518 199668
rect 144610 199640 144638 199860
rect 144776 199792 144782 199844
rect 144834 199792 144840 199844
rect 144546 199588 144552 199640
rect 144604 199600 144638 199640
rect 144604 199588 144610 199600
rect 144150 199532 144184 199572
rect 143960 199520 143966 199532
rect 144178 199520 144184 199532
rect 144236 199520 144242 199572
rect 144638 199520 144644 199572
rect 144696 199560 144702 199572
rect 144794 199560 144822 199792
rect 145070 199764 145098 199860
rect 145024 199736 145098 199764
rect 145024 199640 145052 199736
rect 145162 199708 145190 199860
rect 145098 199656 145104 199708
rect 145156 199668 145190 199708
rect 145156 199656 145162 199668
rect 145006 199588 145012 199640
rect 145064 199588 145070 199640
rect 145254 199628 145282 199940
rect 146542 199940 146754 199968
rect 146542 199912 146570 199940
rect 145328 199860 145334 199912
rect 145386 199860 145392 199912
rect 145604 199860 145610 199912
rect 145662 199860 145668 199912
rect 145788 199860 145794 199912
rect 145846 199860 145852 199912
rect 145880 199860 145886 199912
rect 145938 199860 145944 199912
rect 146064 199900 146070 199912
rect 146036 199860 146070 199900
rect 146122 199860 146128 199912
rect 146156 199860 146162 199912
rect 146214 199860 146220 199912
rect 146524 199860 146530 199912
rect 146582 199860 146588 199912
rect 146616 199860 146622 199912
rect 146674 199860 146680 199912
rect 145116 199600 145282 199628
rect 144696 199532 144822 199560
rect 144696 199520 144702 199532
rect 145116 199424 145144 199600
rect 145346 199572 145374 199860
rect 145466 199588 145472 199640
rect 145524 199628 145530 199640
rect 145622 199628 145650 199860
rect 145806 199764 145834 199860
rect 145524 199600 145650 199628
rect 145760 199736 145834 199764
rect 145524 199588 145530 199600
rect 145760 199572 145788 199736
rect 145898 199708 145926 199860
rect 145834 199656 145840 199708
rect 145892 199668 145926 199708
rect 145892 199656 145898 199668
rect 146036 199572 146064 199860
rect 146174 199832 146202 199860
rect 146128 199804 146202 199832
rect 146128 199708 146156 199804
rect 146202 199724 146208 199776
rect 146260 199764 146266 199776
rect 146634 199764 146662 199860
rect 146260 199736 146662 199764
rect 146260 199724 146266 199736
rect 146110 199656 146116 199708
rect 146168 199656 146174 199708
rect 146726 199640 146754 199940
rect 146818 199940 147352 199968
rect 146818 199912 146846 199940
rect 146800 199860 146806 199912
rect 146858 199860 146864 199912
rect 146892 199860 146898 199912
rect 146950 199860 146956 199912
rect 146984 199860 146990 199912
rect 147042 199860 147048 199912
rect 146910 199776 146938 199860
rect 146846 199724 146852 199776
rect 146904 199736 146938 199776
rect 146904 199724 146910 199736
rect 147002 199708 147030 199860
rect 146938 199656 146944 199708
rect 146996 199668 147030 199708
rect 146996 199656 147002 199668
rect 146726 199600 146760 199640
rect 146754 199588 146760 199600
rect 146812 199588 146818 199640
rect 145282 199520 145288 199572
rect 145340 199532 145374 199572
rect 145340 199520 145346 199532
rect 145742 199520 145748 199572
rect 145800 199520 145806 199572
rect 146018 199520 146024 199572
rect 146076 199520 146082 199572
rect 147324 199436 147352 199940
rect 148750 199912 148778 200008
rect 148842 200008 151262 200036
rect 147812 199860 147818 199912
rect 147870 199860 147876 199912
rect 148364 199860 148370 199912
rect 148422 199860 148428 199912
rect 148456 199860 148462 199912
rect 148514 199860 148520 199912
rect 148640 199860 148646 199912
rect 148698 199860 148704 199912
rect 148732 199860 148738 199912
rect 148790 199860 148796 199912
rect 147674 199588 147680 199640
rect 147732 199628 147738 199640
rect 147830 199628 147858 199860
rect 148382 199776 148410 199860
rect 148474 199832 148502 199860
rect 148474 199804 148548 199832
rect 148520 199776 148548 199804
rect 148658 199776 148686 199860
rect 148382 199736 148416 199776
rect 148410 199724 148416 199736
rect 148468 199724 148474 199776
rect 148502 199724 148508 199776
rect 148560 199724 148566 199776
rect 148594 199724 148600 199776
rect 148652 199736 148686 199776
rect 148652 199724 148658 199736
rect 147732 199600 147858 199628
rect 147732 199588 147738 199600
rect 147398 199452 147404 199504
rect 147456 199492 147462 199504
rect 147582 199492 147588 199504
rect 147456 199464 147588 199492
rect 147456 199452 147462 199464
rect 147582 199452 147588 199464
rect 147640 199452 147646 199504
rect 143460 199396 145144 199424
rect 147306 199384 147312 199436
rect 147364 199384 147370 199436
rect 121362 199316 121368 199368
rect 121420 199356 121426 199368
rect 121420 199328 135760 199356
rect 121420 199316 121426 199328
rect 132126 199248 132132 199300
rect 132184 199288 132190 199300
rect 132770 199288 132776 199300
rect 132184 199260 132776 199288
rect 132184 199248 132190 199260
rect 132770 199248 132776 199260
rect 132828 199248 132834 199300
rect 132954 199248 132960 199300
rect 133012 199288 133018 199300
rect 133690 199288 133696 199300
rect 133012 199260 133696 199288
rect 133012 199248 133018 199260
rect 133690 199248 133696 199260
rect 133748 199248 133754 199300
rect 135732 199288 135760 199328
rect 135806 199316 135812 199368
rect 135864 199316 135870 199368
rect 142154 199356 142160 199368
rect 135916 199328 142160 199356
rect 135916 199288 135944 199328
rect 142154 199316 142160 199328
rect 142212 199316 142218 199368
rect 142522 199316 142528 199368
rect 142580 199356 142586 199368
rect 142580 199328 145236 199356
rect 142580 199316 142586 199328
rect 135732 199260 135944 199288
rect 139486 199248 139492 199300
rect 139544 199288 139550 199300
rect 145098 199288 145104 199300
rect 139544 199260 145104 199288
rect 139544 199248 139550 199260
rect 145098 199248 145104 199260
rect 145156 199248 145162 199300
rect 145208 199288 145236 199328
rect 146386 199316 146392 199368
rect 146444 199356 146450 199368
rect 147398 199356 147404 199368
rect 146444 199328 147404 199356
rect 146444 199316 146450 199328
rect 147398 199316 147404 199328
rect 147456 199316 147462 199368
rect 148842 199288 148870 200008
rect 149578 199940 149790 199968
rect 149578 199912 149606 199940
rect 149008 199860 149014 199912
rect 149066 199860 149072 199912
rect 149284 199860 149290 199912
rect 149342 199860 149348 199912
rect 149468 199860 149474 199912
rect 149526 199860 149532 199912
rect 149560 199860 149566 199912
rect 149618 199860 149624 199912
rect 149652 199860 149658 199912
rect 149710 199860 149716 199912
rect 149026 199572 149054 199860
rect 149302 199640 149330 199860
rect 149486 199640 149514 199860
rect 149302 199600 149336 199640
rect 149330 199588 149336 199600
rect 149388 199588 149394 199640
rect 149486 199600 149520 199640
rect 149514 199588 149520 199600
rect 149572 199588 149578 199640
rect 148962 199520 148968 199572
rect 149020 199532 149054 199572
rect 149020 199520 149026 199532
rect 149146 199520 149152 199572
rect 149204 199560 149210 199572
rect 149670 199560 149698 199860
rect 149204 199532 149698 199560
rect 149204 199520 149210 199532
rect 149606 199452 149612 199504
rect 149664 199492 149670 199504
rect 149762 199492 149790 199940
rect 149664 199464 149790 199492
rect 149900 199940 150986 199968
rect 149664 199452 149670 199464
rect 145208 199260 148870 199288
rect 118418 199180 118424 199232
rect 118476 199220 118482 199232
rect 145650 199220 145656 199232
rect 118476 199192 145656 199220
rect 118476 199180 118482 199192
rect 145650 199180 145656 199192
rect 145708 199180 145714 199232
rect 117130 199112 117136 199164
rect 117188 199152 117194 199164
rect 145374 199152 145380 199164
rect 117188 199124 145380 199152
rect 117188 199112 117194 199124
rect 145374 199112 145380 199124
rect 145432 199112 145438 199164
rect 114370 199044 114376 199096
rect 114428 199084 114434 199096
rect 142338 199084 142344 199096
rect 114428 199056 142344 199084
rect 114428 199044 114434 199056
rect 142338 199044 142344 199056
rect 142396 199044 142402 199096
rect 143350 199044 143356 199096
rect 143408 199084 143414 199096
rect 149900 199084 149928 199940
rect 150958 199912 150986 199940
rect 151234 199912 151262 200008
rect 151786 199912 151814 200144
rect 152798 199940 153010 199968
rect 152798 199912 152826 199940
rect 150112 199860 150118 199912
rect 150170 199860 150176 199912
rect 150940 199860 150946 199912
rect 150998 199860 151004 199912
rect 151216 199860 151222 199912
rect 151274 199860 151280 199912
rect 151768 199860 151774 199912
rect 151826 199860 151832 199912
rect 151952 199860 151958 199912
rect 152010 199860 152016 199912
rect 152228 199900 152234 199912
rect 152200 199860 152234 199900
rect 152286 199860 152292 199912
rect 152320 199860 152326 199912
rect 152378 199860 152384 199912
rect 152412 199860 152418 199912
rect 152470 199860 152476 199912
rect 152688 199860 152694 199912
rect 152746 199860 152752 199912
rect 152780 199860 152786 199912
rect 152838 199860 152844 199912
rect 152872 199860 152878 199912
rect 152930 199860 152936 199912
rect 150130 199764 150158 199860
rect 151970 199832 151998 199860
rect 151970 199804 152136 199832
rect 151998 199764 152004 199776
rect 150130 199736 152004 199764
rect 151998 199724 152004 199736
rect 152056 199724 152062 199776
rect 151906 199656 151912 199708
rect 151964 199696 151970 199708
rect 152108 199696 152136 199804
rect 151964 199668 152136 199696
rect 151964 199656 151970 199668
rect 152200 199640 152228 199860
rect 152338 199832 152366 199860
rect 152292 199804 152366 199832
rect 152292 199776 152320 199804
rect 152430 199776 152458 199860
rect 152274 199724 152280 199776
rect 152332 199724 152338 199776
rect 152366 199724 152372 199776
rect 152424 199736 152458 199776
rect 152706 199776 152734 199860
rect 152890 199776 152918 199860
rect 152706 199736 152740 199776
rect 152424 199724 152430 199736
rect 152734 199724 152740 199736
rect 152792 199724 152798 199776
rect 152826 199724 152832 199776
rect 152884 199736 152918 199776
rect 152884 199724 152890 199736
rect 152182 199588 152188 199640
rect 152240 199588 152246 199640
rect 152982 199628 153010 199940
rect 153258 199940 153838 199968
rect 153056 199860 153062 199912
rect 153114 199860 153120 199912
rect 152798 199600 153010 199628
rect 152798 199504 152826 199600
rect 152734 199452 152740 199504
rect 152792 199464 152826 199504
rect 153074 199492 153102 199860
rect 153258 199560 153286 199940
rect 153810 199912 153838 199940
rect 153902 199912 153930 200756
rect 158686 200648 158714 200756
rect 167656 200716 167684 200756
rect 184216 200728 184244 201096
rect 158594 200620 158714 200648
rect 164206 200688 165614 200716
rect 167656 200688 177896 200716
rect 158594 200512 158622 200620
rect 164206 200580 164234 200688
rect 165586 200648 165614 200688
rect 177758 200648 177764 200660
rect 165586 200620 177764 200648
rect 177758 200608 177764 200620
rect 177816 200608 177822 200660
rect 177868 200648 177896 200688
rect 184198 200676 184204 200728
rect 184256 200676 184262 200728
rect 180058 200648 180064 200660
rect 177868 200620 180064 200648
rect 180058 200608 180064 200620
rect 180116 200608 180122 200660
rect 178034 200580 178040 200592
rect 157628 200484 158622 200512
rect 158686 200552 164234 200580
rect 169726 200552 178040 200580
rect 157628 200036 157656 200484
rect 158686 200444 158714 200552
rect 155282 200008 156782 200036
rect 153332 199860 153338 199912
rect 153390 199860 153396 199912
rect 153424 199860 153430 199912
rect 153482 199900 153488 199912
rect 153482 199872 153562 199900
rect 153482 199860 153488 199872
rect 153350 199776 153378 199860
rect 153350 199736 153384 199776
rect 153378 199724 153384 199736
rect 153436 199724 153442 199776
rect 153534 199640 153562 199872
rect 153608 199860 153614 199912
rect 153666 199860 153672 199912
rect 153700 199860 153706 199912
rect 153758 199860 153764 199912
rect 153792 199860 153798 199912
rect 153850 199860 153856 199912
rect 153884 199860 153890 199912
rect 153942 199860 153948 199912
rect 153976 199860 153982 199912
rect 154034 199860 154040 199912
rect 154252 199860 154258 199912
rect 154310 199900 154316 199912
rect 154436 199900 154442 199912
rect 154310 199860 154344 199900
rect 153626 199776 153654 199860
rect 153718 199832 153746 199860
rect 153718 199804 153792 199832
rect 153626 199736 153660 199776
rect 153654 199724 153660 199736
rect 153712 199724 153718 199776
rect 153764 199708 153792 199804
rect 153994 199776 154022 199860
rect 153930 199724 153936 199776
rect 153988 199736 154022 199776
rect 153988 199724 153994 199736
rect 153746 199656 153752 199708
rect 153804 199656 153810 199708
rect 154316 199640 154344 199860
rect 154408 199860 154442 199900
rect 154494 199860 154500 199912
rect 155172 199860 155178 199912
rect 155230 199860 155236 199912
rect 153534 199600 153568 199640
rect 153562 199588 153568 199600
rect 153620 199588 153626 199640
rect 154298 199588 154304 199640
rect 154356 199588 154362 199640
rect 153838 199560 153844 199572
rect 153258 199532 153844 199560
rect 153838 199520 153844 199532
rect 153896 199520 153902 199572
rect 154114 199520 154120 199572
rect 154172 199560 154178 199572
rect 154408 199560 154436 199860
rect 155190 199708 155218 199860
rect 155282 199832 155310 200008
rect 155356 199860 155362 199912
rect 155414 199860 155420 199912
rect 155448 199860 155454 199912
rect 155506 199860 155512 199912
rect 155724 199900 155730 199912
rect 155696 199860 155730 199900
rect 155782 199860 155788 199912
rect 155816 199860 155822 199912
rect 155874 199860 155880 199912
rect 155908 199860 155914 199912
rect 155966 199860 155972 199912
rect 156368 199860 156374 199912
rect 156426 199860 156432 199912
rect 156460 199860 156466 199912
rect 156518 199860 156524 199912
rect 156552 199860 156558 199912
rect 156610 199860 156616 199912
rect 155374 199832 155402 199860
rect 155282 199804 155402 199832
rect 155466 199776 155494 199860
rect 155402 199724 155408 199776
rect 155460 199736 155494 199776
rect 155460 199724 155466 199736
rect 155190 199668 155224 199708
rect 155218 199656 155224 199668
rect 155276 199656 155282 199708
rect 155696 199640 155724 199860
rect 155834 199832 155862 199860
rect 155788 199804 155862 199832
rect 155788 199776 155816 199804
rect 155926 199776 155954 199860
rect 155770 199724 155776 199776
rect 155828 199724 155834 199776
rect 155862 199724 155868 199776
rect 155920 199736 155954 199776
rect 155920 199724 155926 199736
rect 155678 199588 155684 199640
rect 155736 199588 155742 199640
rect 154172 199532 154436 199560
rect 154172 199520 154178 199532
rect 153194 199492 153200 199504
rect 153074 199464 153200 199492
rect 152792 199452 152798 199464
rect 153194 199452 153200 199464
rect 153252 199452 153258 199504
rect 156230 199452 156236 199504
rect 156288 199492 156294 199504
rect 156386 199492 156414 199860
rect 156288 199464 156414 199492
rect 156288 199452 156294 199464
rect 156478 199436 156506 199860
rect 156570 199640 156598 199860
rect 156570 199600 156604 199640
rect 156598 199588 156604 199600
rect 156656 199588 156662 199640
rect 156754 199560 156782 200008
rect 157214 200008 157656 200036
rect 157720 200416 158714 200444
rect 161722 200484 168098 200512
rect 156846 199940 157150 199968
rect 156846 199696 156874 199940
rect 157122 199912 157150 199940
rect 156920 199860 156926 199912
rect 156978 199860 156984 199912
rect 157012 199860 157018 199912
rect 157070 199860 157076 199912
rect 157104 199860 157110 199912
rect 157162 199860 157168 199912
rect 156938 199764 156966 199860
rect 157030 199832 157058 199860
rect 157214 199832 157242 200008
rect 157472 199860 157478 199912
rect 157530 199860 157536 199912
rect 157030 199804 157242 199832
rect 157490 199776 157518 199860
rect 156938 199736 157196 199764
rect 157490 199736 157524 199776
rect 157058 199696 157064 199708
rect 156846 199668 157064 199696
rect 157058 199656 157064 199668
rect 157116 199656 157122 199708
rect 156966 199588 156972 199640
rect 157024 199628 157030 199640
rect 157168 199628 157196 199736
rect 157518 199724 157524 199736
rect 157576 199724 157582 199776
rect 157024 199600 157196 199628
rect 157024 199588 157030 199600
rect 157720 199560 157748 200416
rect 158318 199940 158898 199968
rect 158318 199912 158346 199940
rect 157840 199860 157846 199912
rect 157898 199860 157904 199912
rect 158024 199860 158030 199912
rect 158082 199860 158088 199912
rect 158300 199860 158306 199912
rect 158358 199860 158364 199912
rect 158392 199860 158398 199912
rect 158450 199860 158456 199912
rect 158576 199900 158582 199912
rect 158548 199860 158582 199900
rect 158634 199860 158640 199912
rect 158668 199860 158674 199912
rect 158726 199860 158732 199912
rect 158760 199860 158766 199912
rect 158818 199860 158824 199912
rect 156754 199532 157748 199560
rect 157858 199560 157886 199860
rect 158042 199640 158070 199860
rect 158410 199708 158438 199860
rect 158548 199708 158576 199860
rect 158686 199832 158714 199860
rect 158640 199804 158714 199832
rect 158640 199776 158668 199804
rect 158778 199776 158806 199860
rect 158622 199724 158628 199776
rect 158680 199724 158686 199776
rect 158714 199724 158720 199776
rect 158772 199736 158806 199776
rect 158772 199724 158778 199736
rect 158346 199656 158352 199708
rect 158404 199668 158438 199708
rect 158404 199656 158410 199668
rect 158530 199656 158536 199708
rect 158588 199656 158594 199708
rect 157978 199588 157984 199640
rect 158036 199600 158070 199640
rect 158870 199628 158898 199940
rect 161722 199912 161750 200484
rect 168070 200376 168098 200484
rect 169726 200376 169754 200552
rect 178034 200540 178040 200552
rect 178092 200540 178098 200592
rect 178126 200540 178132 200592
rect 178184 200580 178190 200592
rect 191926 200580 191932 200592
rect 178184 200552 191932 200580
rect 178184 200540 178190 200552
rect 191926 200540 191932 200552
rect 191984 200540 191990 200592
rect 177942 200472 177948 200524
rect 178000 200512 178006 200524
rect 193214 200512 193220 200524
rect 178000 200484 193220 200512
rect 178000 200472 178006 200484
rect 193214 200472 193220 200484
rect 193272 200472 193278 200524
rect 180334 200444 180340 200456
rect 168070 200348 169754 200376
rect 170186 200416 180340 200444
rect 170186 200308 170214 200416
rect 180334 200404 180340 200416
rect 180392 200404 180398 200456
rect 178402 200376 178408 200388
rect 168070 200280 170214 200308
rect 170370 200348 178408 200376
rect 165586 200008 168006 200036
rect 162274 199940 162762 199968
rect 158944 199860 158950 199912
rect 159002 199860 159008 199912
rect 159036 199860 159042 199912
rect 159094 199860 159100 199912
rect 159128 199860 159134 199912
rect 159186 199900 159192 199912
rect 159186 199872 159496 199900
rect 159186 199860 159192 199872
rect 158962 199708 158990 199860
rect 159054 199832 159082 199860
rect 159054 199804 159128 199832
rect 159100 199708 159128 199804
rect 158962 199668 158996 199708
rect 158990 199656 158996 199668
rect 159048 199656 159054 199708
rect 159082 199656 159088 199708
rect 159140 199656 159146 199708
rect 159468 199640 159496 199872
rect 159588 199860 159594 199912
rect 159646 199860 159652 199912
rect 159772 199860 159778 199912
rect 159830 199860 159836 199912
rect 159864 199860 159870 199912
rect 159922 199860 159928 199912
rect 160048 199860 160054 199912
rect 160106 199860 160112 199912
rect 160140 199860 160146 199912
rect 160198 199860 160204 199912
rect 160232 199860 160238 199912
rect 160290 199860 160296 199912
rect 160324 199860 160330 199912
rect 160382 199900 160388 199912
rect 160692 199900 160698 199912
rect 160382 199872 160600 199900
rect 160382 199860 160388 199872
rect 159606 199776 159634 199860
rect 159606 199736 159640 199776
rect 159634 199724 159640 199736
rect 159692 199724 159698 199776
rect 159790 199640 159818 199860
rect 159266 199628 159272 199640
rect 158870 199600 159272 199628
rect 158036 199588 158042 199600
rect 159266 199588 159272 199600
rect 159324 199588 159330 199640
rect 159450 199588 159456 199640
rect 159508 199588 159514 199640
rect 159726 199588 159732 199640
rect 159784 199600 159818 199640
rect 159784 199588 159790 199600
rect 158622 199560 158628 199572
rect 157858 199532 158628 199560
rect 158622 199520 158628 199532
rect 158680 199520 158686 199572
rect 158806 199520 158812 199572
rect 158864 199560 158870 199572
rect 159882 199560 159910 199860
rect 158864 199532 159910 199560
rect 158864 199520 158870 199532
rect 160066 199492 160094 199860
rect 160158 199776 160186 199860
rect 160250 199832 160278 199860
rect 160250 199804 160324 199832
rect 160296 199776 160324 199804
rect 160158 199736 160192 199776
rect 160186 199724 160192 199736
rect 160244 199724 160250 199776
rect 160278 199724 160284 199776
rect 160336 199724 160342 199776
rect 160572 199560 160600 199872
rect 160664 199860 160698 199900
rect 160750 199860 160756 199912
rect 160876 199860 160882 199912
rect 160934 199860 160940 199912
rect 161060 199860 161066 199912
rect 161118 199860 161124 199912
rect 161152 199860 161158 199912
rect 161210 199860 161216 199912
rect 161612 199900 161618 199912
rect 161584 199860 161618 199900
rect 161670 199860 161676 199912
rect 161704 199860 161710 199912
rect 161762 199860 161768 199912
rect 161796 199860 161802 199912
rect 161854 199860 161860 199912
rect 161888 199860 161894 199912
rect 161946 199860 161952 199912
rect 160664 199776 160692 199860
rect 160646 199724 160652 199776
rect 160704 199724 160710 199776
rect 160894 199764 160922 199860
rect 161078 199764 161106 199860
rect 160848 199736 160922 199764
rect 161032 199736 161106 199764
rect 160848 199640 160876 199736
rect 161032 199640 161060 199736
rect 161170 199708 161198 199860
rect 161106 199656 161112 199708
rect 161164 199668 161198 199708
rect 161164 199656 161170 199668
rect 160830 199588 160836 199640
rect 160888 199588 160894 199640
rect 161014 199588 161020 199640
rect 161072 199588 161078 199640
rect 161474 199560 161480 199572
rect 160572 199532 161480 199560
rect 161474 199520 161480 199532
rect 161532 199520 161538 199572
rect 160462 199492 160468 199504
rect 160066 199464 160468 199492
rect 160462 199452 160468 199464
rect 160520 199452 160526 199504
rect 161584 199492 161612 199860
rect 161658 199724 161664 199776
rect 161716 199764 161722 199776
rect 161814 199764 161842 199860
rect 161716 199736 161842 199764
rect 161716 199724 161722 199736
rect 161906 199708 161934 199860
rect 162072 199792 162078 199844
rect 162130 199792 162136 199844
rect 161842 199656 161848 199708
rect 161900 199668 161934 199708
rect 161900 199656 161906 199668
rect 162090 199572 162118 199792
rect 162274 199696 162302 199940
rect 162734 199912 162762 199940
rect 162826 199940 163222 199968
rect 162624 199900 162630 199912
rect 162026 199520 162032 199572
rect 162084 199532 162118 199572
rect 162228 199668 162302 199696
rect 162366 199872 162630 199900
rect 162228 199560 162256 199668
rect 162366 199640 162394 199872
rect 162624 199860 162630 199872
rect 162682 199860 162688 199912
rect 162716 199860 162722 199912
rect 162774 199860 162780 199912
rect 162532 199792 162538 199844
rect 162590 199792 162596 199844
rect 162302 199588 162308 199640
rect 162360 199600 162394 199640
rect 162360 199588 162366 199600
rect 162550 199572 162578 199792
rect 162826 199640 162854 199940
rect 163194 199912 163222 199940
rect 162900 199860 162906 199912
rect 162958 199860 162964 199912
rect 163084 199860 163090 199912
rect 163142 199860 163148 199912
rect 163176 199860 163182 199912
rect 163234 199860 163240 199912
rect 163268 199860 163274 199912
rect 163326 199860 163332 199912
rect 163360 199860 163366 199912
rect 163418 199900 163424 199912
rect 163820 199900 163826 199912
rect 163418 199872 163590 199900
rect 163418 199860 163424 199872
rect 162762 199588 162768 199640
rect 162820 199600 162854 199640
rect 162918 199628 162946 199860
rect 163102 199776 163130 199860
rect 163286 199776 163314 199860
rect 163452 199832 163458 199844
rect 163102 199736 163136 199776
rect 163130 199724 163136 199736
rect 163188 199724 163194 199776
rect 163222 199724 163228 199776
rect 163280 199736 163314 199776
rect 163424 199792 163458 199832
rect 163510 199792 163516 199844
rect 163280 199724 163286 199736
rect 163424 199708 163452 199792
rect 163562 199764 163590 199872
rect 163792 199860 163826 199900
rect 163878 199860 163884 199912
rect 163912 199860 163918 199912
rect 163970 199860 163976 199912
rect 164372 199860 164378 199912
rect 164430 199900 164436 199912
rect 164430 199872 164694 199900
rect 164430 199860 164436 199872
rect 163636 199792 163642 199844
rect 163694 199792 163700 199844
rect 163516 199736 163590 199764
rect 163406 199656 163412 199708
rect 163464 199656 163470 199708
rect 163038 199628 163044 199640
rect 162918 199600 163044 199628
rect 162820 199588 162826 199600
rect 163038 199588 163044 199600
rect 163096 199588 163102 199640
rect 162394 199560 162400 199572
rect 162228 199532 162400 199560
rect 162084 199520 162090 199532
rect 162394 199520 162400 199532
rect 162452 199520 162458 199572
rect 162486 199520 162492 199572
rect 162544 199532 162578 199572
rect 163516 199560 163544 199736
rect 163654 199708 163682 199792
rect 163792 199708 163820 199860
rect 163930 199764 163958 199860
rect 164464 199792 164470 199844
rect 164522 199792 164528 199844
rect 163930 199736 164188 199764
rect 163590 199656 163596 199708
rect 163648 199668 163682 199708
rect 163648 199656 163654 199668
rect 163774 199656 163780 199708
rect 163832 199656 163838 199708
rect 164160 199560 164188 199736
rect 164234 199656 164240 199708
rect 164292 199696 164298 199708
rect 164292 199668 164372 199696
rect 164292 199656 164298 199668
rect 164344 199640 164372 199668
rect 164326 199588 164332 199640
rect 164384 199588 164390 199640
rect 164482 199572 164510 199792
rect 164234 199560 164240 199572
rect 163516 199532 164096 199560
rect 164160 199532 164240 199560
rect 162544 199520 162550 199532
rect 163866 199492 163872 199504
rect 161584 199464 163872 199492
rect 163866 199452 163872 199464
rect 163924 199452 163930 199504
rect 164068 199492 164096 199532
rect 164234 199520 164240 199532
rect 164292 199520 164298 199572
rect 164418 199520 164424 199572
rect 164476 199532 164510 199572
rect 164476 199520 164482 199532
rect 164142 199492 164148 199504
rect 164068 199464 164148 199492
rect 164142 199452 164148 199464
rect 164200 199452 164206 199504
rect 164666 199492 164694 199872
rect 165200 199860 165206 199912
rect 165258 199860 165264 199912
rect 165292 199860 165298 199912
rect 165350 199860 165356 199912
rect 165384 199860 165390 199912
rect 165442 199860 165448 199912
rect 165476 199860 165482 199912
rect 165534 199860 165540 199912
rect 164740 199792 164746 199844
rect 164798 199792 164804 199844
rect 165218 199832 165246 199860
rect 165172 199804 165246 199832
rect 164758 199560 164786 199792
rect 164924 199724 164930 199776
rect 164982 199724 164988 199776
rect 164942 199640 164970 199724
rect 165172 199708 165200 199804
rect 165310 199776 165338 199860
rect 165246 199724 165252 199776
rect 165304 199736 165338 199776
rect 165304 199724 165310 199736
rect 165154 199656 165160 199708
rect 165212 199656 165218 199708
rect 164878 199588 164884 199640
rect 164936 199600 164970 199640
rect 165402 199640 165430 199860
rect 165494 199696 165522 199860
rect 165586 199776 165614 200008
rect 165862 199940 167040 199968
rect 165862 199912 165890 199940
rect 165844 199860 165850 199912
rect 165902 199860 165908 199912
rect 165936 199860 165942 199912
rect 165994 199860 166000 199912
rect 166028 199860 166034 199912
rect 166086 199860 166092 199912
rect 166488 199900 166494 199912
rect 166138 199872 166494 199900
rect 165954 199832 165982 199860
rect 165908 199804 165982 199832
rect 165568 199724 165574 199776
rect 165626 199724 165632 199776
rect 165798 199696 165804 199708
rect 165494 199668 165804 199696
rect 165798 199656 165804 199668
rect 165856 199656 165862 199708
rect 165908 199640 165936 199804
rect 166046 199708 166074 199860
rect 165982 199656 165988 199708
rect 166040 199668 166074 199708
rect 166040 199656 166046 199668
rect 166138 199640 166166 199872
rect 166488 199860 166494 199872
rect 166546 199860 166552 199912
rect 166856 199860 166862 199912
rect 166914 199860 166920 199912
rect 166672 199792 166678 199844
rect 166730 199792 166736 199844
rect 166304 199724 166310 199776
rect 166362 199724 166368 199776
rect 165402 199600 165436 199640
rect 164936 199588 164942 199600
rect 165430 199588 165436 199600
rect 165488 199588 165494 199640
rect 165890 199588 165896 199640
rect 165948 199588 165954 199640
rect 166074 199588 166080 199640
rect 166132 199600 166166 199640
rect 166132 199588 166138 199600
rect 166322 199572 166350 199724
rect 166690 199640 166718 199792
rect 166626 199588 166632 199640
rect 166684 199600 166718 199640
rect 166684 199588 166690 199600
rect 165522 199560 165528 199572
rect 164758 199532 165528 199560
rect 165522 199520 165528 199532
rect 165580 199520 165586 199572
rect 166322 199532 166356 199572
rect 166350 199520 166356 199532
rect 166408 199520 166414 199572
rect 166442 199520 166448 199572
rect 166500 199560 166506 199572
rect 166874 199560 166902 199860
rect 167012 199640 167040 199940
rect 167592 199900 167598 199912
rect 167564 199860 167598 199900
rect 167650 199860 167656 199912
rect 167684 199860 167690 199912
rect 167742 199860 167748 199912
rect 167776 199860 167782 199912
rect 167834 199860 167840 199912
rect 167868 199860 167874 199912
rect 167926 199860 167932 199912
rect 167224 199792 167230 199844
rect 167282 199792 167288 199844
rect 167408 199792 167414 199844
rect 167466 199792 167472 199844
rect 167132 199764 167138 199776
rect 167104 199724 167138 199764
rect 167190 199724 167196 199776
rect 166994 199588 167000 199640
rect 167052 199588 167058 199640
rect 167104 199572 167132 199724
rect 167242 199696 167270 199792
rect 167196 199668 167270 199696
rect 167196 199640 167224 199668
rect 167426 199640 167454 199792
rect 167564 199708 167592 199860
rect 167702 199832 167730 199860
rect 167656 199804 167730 199832
rect 167656 199708 167684 199804
rect 167794 199708 167822 199860
rect 167546 199656 167552 199708
rect 167604 199656 167610 199708
rect 167638 199656 167644 199708
rect 167696 199656 167702 199708
rect 167730 199656 167736 199708
rect 167788 199668 167822 199708
rect 167788 199656 167794 199668
rect 167886 199640 167914 199860
rect 167178 199588 167184 199640
rect 167236 199588 167242 199640
rect 167362 199588 167368 199640
rect 167420 199600 167454 199640
rect 167420 199588 167426 199600
rect 167822 199588 167828 199640
rect 167880 199600 167914 199640
rect 167880 199588 167886 199600
rect 166500 199532 166902 199560
rect 166500 199520 166506 199532
rect 167086 199520 167092 199572
rect 167144 199520 167150 199572
rect 167978 199560 168006 200008
rect 168070 199912 168098 200280
rect 170370 200240 170398 200348
rect 178402 200336 178408 200348
rect 178460 200336 178466 200388
rect 177758 200268 177764 200320
rect 177816 200308 177822 200320
rect 189258 200308 189264 200320
rect 177816 200280 189264 200308
rect 177816 200268 177822 200280
rect 189258 200268 189264 200280
rect 189316 200268 189322 200320
rect 169726 200212 170398 200240
rect 169726 200104 169754 200212
rect 177850 200200 177856 200252
rect 177908 200240 177914 200252
rect 191834 200240 191840 200252
rect 177908 200212 191840 200240
rect 177908 200200 177914 200212
rect 191834 200200 191840 200212
rect 191892 200200 191898 200252
rect 168530 200076 169754 200104
rect 170094 200144 170398 200172
rect 168530 199912 168558 200076
rect 170094 199968 170122 200144
rect 170370 200104 170398 200144
rect 178034 200132 178040 200184
rect 178092 200172 178098 200184
rect 196342 200172 196348 200184
rect 178092 200144 196348 200172
rect 178092 200132 178098 200144
rect 196342 200132 196348 200144
rect 196400 200132 196406 200184
rect 170370 200076 186314 200104
rect 169312 199940 170122 199968
rect 175338 199940 175918 199968
rect 168052 199860 168058 199912
rect 168110 199860 168116 199912
rect 168144 199860 168150 199912
rect 168202 199860 168208 199912
rect 168512 199860 168518 199912
rect 168570 199860 168576 199912
rect 168788 199860 168794 199912
rect 168846 199860 168852 199912
rect 168880 199860 168886 199912
rect 168938 199860 168944 199912
rect 169064 199860 169070 199912
rect 169122 199860 169128 199912
rect 169156 199860 169162 199912
rect 169214 199860 169220 199912
rect 168162 199776 168190 199860
rect 168420 199792 168426 199844
rect 168478 199832 168484 199844
rect 168806 199832 168834 199860
rect 168478 199792 168512 199832
rect 168098 199724 168104 199776
rect 168156 199736 168190 199776
rect 168156 199724 168162 199736
rect 168484 199708 168512 199792
rect 168576 199804 168834 199832
rect 168466 199656 168472 199708
rect 168524 199656 168530 199708
rect 168576 199572 168604 199804
rect 168898 199708 168926 199860
rect 169082 199776 169110 199860
rect 169018 199724 169024 199776
rect 169076 199736 169110 199776
rect 169076 199724 169082 199736
rect 169174 199708 169202 199860
rect 168834 199656 168840 199708
rect 168892 199668 168926 199708
rect 168892 199656 168898 199668
rect 169110 199656 169116 199708
rect 169168 199668 169202 199708
rect 169168 199656 169174 199668
rect 169312 199640 169340 199940
rect 169524 199900 169530 199912
rect 169496 199860 169530 199900
rect 169582 199860 169588 199912
rect 169708 199900 169714 199912
rect 169680 199860 169714 199900
rect 169766 199860 169772 199912
rect 169800 199860 169806 199912
rect 169858 199860 169864 199912
rect 169892 199860 169898 199912
rect 169950 199860 169956 199912
rect 170168 199860 170174 199912
rect 170226 199860 170232 199912
rect 170646 199872 170950 199900
rect 169496 199776 169524 199860
rect 169478 199724 169484 199776
rect 169536 199724 169542 199776
rect 169680 199708 169708 199860
rect 169818 199832 169846 199860
rect 169772 199804 169846 199832
rect 169772 199708 169800 199804
rect 169910 199776 169938 199860
rect 169846 199724 169852 199776
rect 169904 199736 169938 199776
rect 169904 199724 169910 199736
rect 169662 199656 169668 199708
rect 169720 199656 169726 199708
rect 169754 199656 169760 199708
rect 169812 199656 169818 199708
rect 169294 199588 169300 199640
rect 169352 199588 169358 199640
rect 170186 199628 170214 199860
rect 170444 199792 170450 199844
rect 170502 199792 170508 199844
rect 170462 199640 170490 199792
rect 170646 199764 170674 199872
rect 170922 199844 170950 199872
rect 170996 199860 171002 199912
rect 171054 199860 171060 199912
rect 171180 199860 171186 199912
rect 171238 199860 171244 199912
rect 171364 199860 171370 199912
rect 171422 199860 171428 199912
rect 171456 199860 171462 199912
rect 171514 199860 171520 199912
rect 171548 199860 171554 199912
rect 171606 199860 171612 199912
rect 171640 199860 171646 199912
rect 171698 199860 171704 199912
rect 171916 199860 171922 199912
rect 171974 199860 171980 199912
rect 172192 199860 172198 199912
rect 172250 199860 172256 199912
rect 172284 199860 172290 199912
rect 172342 199860 172348 199912
rect 172652 199860 172658 199912
rect 172710 199860 172716 199912
rect 172836 199860 172842 199912
rect 172894 199860 172900 199912
rect 173572 199860 173578 199912
rect 173630 199860 173636 199912
rect 174032 199860 174038 199912
rect 174090 199860 174096 199912
rect 174584 199860 174590 199912
rect 174642 199860 174648 199912
rect 174676 199860 174682 199912
rect 174734 199860 174740 199912
rect 174860 199860 174866 199912
rect 174918 199860 174924 199912
rect 175228 199860 175234 199912
rect 175286 199860 175292 199912
rect 170720 199792 170726 199844
rect 170778 199792 170784 199844
rect 170812 199792 170818 199844
rect 170870 199792 170876 199844
rect 170904 199792 170910 199844
rect 170962 199792 170968 199844
rect 170600 199736 170674 199764
rect 170306 199628 170312 199640
rect 170186 199600 170312 199628
rect 170306 199588 170312 199600
rect 170364 199588 170370 199640
rect 170462 199600 170496 199640
rect 170490 199588 170496 199600
rect 170548 199588 170554 199640
rect 167978 199532 168328 199560
rect 168300 199504 168328 199532
rect 168558 199520 168564 199572
rect 168616 199520 168622 199572
rect 167914 199492 167920 199504
rect 164666 199464 167920 199492
rect 167914 199452 167920 199464
rect 167972 199452 167978 199504
rect 168282 199452 168288 199504
rect 168340 199452 168346 199504
rect 170600 199492 170628 199736
rect 170738 199696 170766 199792
rect 170692 199668 170766 199696
rect 170692 199572 170720 199668
rect 170830 199640 170858 199792
rect 171014 199640 171042 199860
rect 171198 199640 171226 199860
rect 171382 199832 171410 199860
rect 170766 199588 170772 199640
rect 170824 199600 170858 199640
rect 170824 199588 170830 199600
rect 170950 199588 170956 199640
rect 171008 199600 171042 199640
rect 171008 199588 171014 199600
rect 171134 199588 171140 199640
rect 171192 199600 171226 199640
rect 171336 199804 171410 199832
rect 171192 199588 171198 199600
rect 170674 199520 170680 199572
rect 170732 199520 170738 199572
rect 171336 199504 171364 199804
rect 171474 199764 171502 199860
rect 171428 199736 171502 199764
rect 171428 199708 171456 199736
rect 171566 199708 171594 199860
rect 171410 199656 171416 199708
rect 171468 199656 171474 199708
rect 171502 199656 171508 199708
rect 171560 199668 171594 199708
rect 171560 199656 171566 199668
rect 170858 199492 170864 199504
rect 170600 199464 170864 199492
rect 170858 199452 170864 199464
rect 170916 199452 170922 199504
rect 171318 199452 171324 199504
rect 171376 199452 171382 199504
rect 171658 199492 171686 199860
rect 171934 199628 171962 199860
rect 172210 199764 172238 199860
rect 172302 199832 172330 199860
rect 172302 199804 172468 199832
rect 172330 199764 172336 199776
rect 172210 199736 172336 199764
rect 172330 199724 172336 199736
rect 172388 199724 172394 199776
rect 172238 199656 172244 199708
rect 172296 199696 172302 199708
rect 172440 199696 172468 199804
rect 172296 199668 172468 199696
rect 172670 199708 172698 199860
rect 172670 199668 172704 199708
rect 172296 199656 172302 199668
rect 172698 199656 172704 199668
rect 172756 199656 172762 199708
rect 172054 199628 172060 199640
rect 171934 199600 172060 199628
rect 172054 199588 172060 199600
rect 172112 199588 172118 199640
rect 172606 199588 172612 199640
rect 172664 199628 172670 199640
rect 172854 199628 172882 199860
rect 172664 199600 172882 199628
rect 172664 199588 172670 199600
rect 173590 199560 173618 199860
rect 174050 199776 174078 199860
rect 174602 199832 174630 199860
rect 174556 199804 174630 199832
rect 174050 199736 174084 199776
rect 174078 199724 174084 199736
rect 174136 199724 174142 199776
rect 173802 199560 173808 199572
rect 173590 199532 173808 199560
rect 173802 199520 173808 199532
rect 173860 199520 173866 199572
rect 174556 199560 174584 199804
rect 174694 199708 174722 199860
rect 174630 199656 174636 199708
rect 174688 199668 174722 199708
rect 174688 199656 174694 199668
rect 174878 199628 174906 199860
rect 175246 199776 175274 199860
rect 175182 199724 175188 199776
rect 175240 199736 175274 199776
rect 175240 199724 175246 199736
rect 175090 199628 175096 199640
rect 174878 199600 175096 199628
rect 175090 199588 175096 199600
rect 175148 199588 175154 199640
rect 175338 199628 175366 199940
rect 175890 199912 175918 199940
rect 176074 199940 179276 199968
rect 176074 199912 176102 199940
rect 175412 199860 175418 199912
rect 175470 199860 175476 199912
rect 175504 199860 175510 199912
rect 175562 199860 175568 199912
rect 175872 199860 175878 199912
rect 175930 199860 175936 199912
rect 176056 199860 176062 199912
rect 176114 199860 176120 199912
rect 176240 199860 176246 199912
rect 176298 199860 176304 199912
rect 176332 199860 176338 199912
rect 176390 199860 176396 199912
rect 176792 199860 176798 199912
rect 176850 199860 176856 199912
rect 177068 199900 177074 199912
rect 177040 199860 177074 199900
rect 177126 199860 177132 199912
rect 177160 199860 177166 199912
rect 177218 199860 177224 199912
rect 177252 199860 177258 199912
rect 177310 199860 177316 199912
rect 177344 199860 177350 199912
rect 177402 199900 177408 199912
rect 177850 199900 177856 199912
rect 177402 199872 177856 199900
rect 177402 199860 177408 199872
rect 177850 199860 177856 199872
rect 177908 199860 177914 199912
rect 175430 199708 175458 199860
rect 175522 199764 175550 199860
rect 176258 199832 176286 199860
rect 176120 199804 176286 199832
rect 175522 199736 175964 199764
rect 175430 199668 175464 199708
rect 175458 199656 175464 199668
rect 175516 199656 175522 199708
rect 175936 199640 175964 199736
rect 175734 199628 175740 199640
rect 175338 199600 175740 199628
rect 175734 199588 175740 199600
rect 175792 199588 175798 199640
rect 175918 199588 175924 199640
rect 175976 199588 175982 199640
rect 174906 199560 174912 199572
rect 174556 199532 174912 199560
rect 174906 199520 174912 199532
rect 174964 199520 174970 199572
rect 175274 199492 175280 199504
rect 171658 199464 175280 199492
rect 175274 199452 175280 199464
rect 175332 199452 175338 199504
rect 176120 199492 176148 199804
rect 176350 199776 176378 199860
rect 176286 199724 176292 199776
rect 176344 199736 176378 199776
rect 176344 199724 176350 199736
rect 176810 199572 176838 199860
rect 176810 199532 176844 199572
rect 176838 199520 176844 199532
rect 176896 199520 176902 199572
rect 176654 199492 176660 199504
rect 176120 199464 176660 199492
rect 176654 199452 176660 199464
rect 176712 199452 176718 199504
rect 177040 199492 177068 199860
rect 177178 199696 177206 199860
rect 177132 199668 177206 199696
rect 177132 199640 177160 199668
rect 177270 199640 177298 199860
rect 179248 199832 179276 199940
rect 186286 199900 186314 200076
rect 186682 199900 186688 199912
rect 186286 199872 186688 199900
rect 186682 199860 186688 199872
rect 186740 199860 186746 199912
rect 187602 199832 187608 199844
rect 179248 199804 187608 199832
rect 187602 199792 187608 199804
rect 187660 199792 187666 199844
rect 177114 199588 177120 199640
rect 177172 199588 177178 199640
rect 177206 199588 177212 199640
rect 177264 199600 177298 199640
rect 177264 199588 177270 199600
rect 177390 199588 177396 199640
rect 177448 199628 177454 199640
rect 215662 199628 215668 199640
rect 177448 199600 215668 199628
rect 177448 199588 177454 199600
rect 215662 199588 215668 199600
rect 215720 199588 215726 199640
rect 178586 199520 178592 199572
rect 178644 199560 178650 199572
rect 215386 199560 215392 199572
rect 178644 199532 215392 199560
rect 178644 199520 178650 199532
rect 215386 199520 215392 199532
rect 215444 199520 215450 199572
rect 177298 199492 177304 199504
rect 177040 199464 177304 199492
rect 177298 199452 177304 199464
rect 177356 199452 177362 199504
rect 152918 199384 152924 199436
rect 152976 199424 152982 199436
rect 153102 199424 153108 199436
rect 152976 199396 153108 199424
rect 152976 199384 152982 199396
rect 153102 199384 153108 199396
rect 153160 199384 153166 199436
rect 156414 199384 156420 199436
rect 156472 199396 156506 199436
rect 156472 199384 156478 199396
rect 158346 199384 158352 199436
rect 158404 199424 158410 199436
rect 178678 199424 178684 199436
rect 158404 199396 178684 199424
rect 158404 199384 158410 199396
rect 178678 199384 178684 199396
rect 178736 199384 178742 199436
rect 182818 199384 182824 199436
rect 182876 199424 182882 199436
rect 190454 199424 190460 199436
rect 182876 199396 190460 199424
rect 182876 199384 182882 199396
rect 190454 199384 190460 199396
rect 190512 199384 190518 199436
rect 152550 199316 152556 199368
rect 152608 199356 152614 199368
rect 160094 199356 160100 199368
rect 152608 199328 160100 199356
rect 152608 199316 152614 199328
rect 160094 199316 160100 199328
rect 160152 199316 160158 199368
rect 215478 199356 215484 199368
rect 160848 199328 215484 199356
rect 153562 199248 153568 199300
rect 153620 199288 153626 199300
rect 156782 199288 156788 199300
rect 153620 199260 156788 199288
rect 153620 199248 153626 199260
rect 156782 199248 156788 199260
rect 156840 199248 156846 199300
rect 151998 199180 152004 199232
rect 152056 199220 152062 199232
rect 160848 199220 160876 199328
rect 215478 199316 215484 199328
rect 215536 199316 215542 199368
rect 164418 199248 164424 199300
rect 164476 199288 164482 199300
rect 198734 199288 198740 199300
rect 164476 199260 198740 199288
rect 164476 199248 164482 199260
rect 198734 199248 198740 199260
rect 198792 199248 198798 199300
rect 189994 199220 190000 199232
rect 152056 199192 160876 199220
rect 161446 199192 190000 199220
rect 152056 199180 152062 199192
rect 143408 199056 149928 199084
rect 143408 199044 143414 199056
rect 116946 198976 116952 199028
rect 117004 199016 117010 199028
rect 145926 199016 145932 199028
rect 117004 198988 145932 199016
rect 117004 198976 117010 198988
rect 145926 198976 145932 198988
rect 145984 198976 145990 199028
rect 115658 198908 115664 198960
rect 115716 198948 115722 198960
rect 147030 198948 147036 198960
rect 115716 198920 147036 198948
rect 115716 198908 115722 198920
rect 147030 198908 147036 198920
rect 147088 198908 147094 198960
rect 155126 198908 155132 198960
rect 155184 198948 155190 198960
rect 161446 198948 161474 199192
rect 189994 199180 190000 199192
rect 190052 199180 190058 199232
rect 170122 199112 170128 199164
rect 170180 199152 170186 199164
rect 200298 199152 200304 199164
rect 170180 199124 200304 199152
rect 170180 199112 170186 199124
rect 200298 199112 200304 199124
rect 200356 199112 200362 199164
rect 178402 199044 178408 199096
rect 178460 199084 178466 199096
rect 203150 199084 203156 199096
rect 178460 199056 203156 199084
rect 178460 199044 178466 199056
rect 203150 199044 203156 199056
rect 203208 199044 203214 199096
rect 161934 198976 161940 199028
rect 161992 199016 161998 199028
rect 196158 199016 196164 199028
rect 161992 198988 196164 199016
rect 161992 198976 161998 198988
rect 196158 198976 196164 198988
rect 196216 198976 196222 199028
rect 155184 198920 161474 198948
rect 155184 198908 155190 198920
rect 168374 198908 168380 198960
rect 168432 198948 168438 198960
rect 180150 198948 180156 198960
rect 168432 198920 180156 198948
rect 168432 198908 168438 198920
rect 180150 198908 180156 198920
rect 180208 198908 180214 198960
rect 126422 198840 126428 198892
rect 126480 198880 126486 198892
rect 144914 198880 144920 198892
rect 126480 198852 144920 198880
rect 126480 198840 126486 198852
rect 144914 198840 144920 198852
rect 144972 198840 144978 198892
rect 161474 198840 161480 198892
rect 161532 198880 161538 198892
rect 178862 198880 178868 198892
rect 161532 198852 178868 198880
rect 161532 198840 161538 198852
rect 178862 198840 178868 198852
rect 178920 198840 178926 198892
rect 121178 198772 121184 198824
rect 121236 198812 121242 198824
rect 139486 198812 139492 198824
rect 121236 198784 139492 198812
rect 121236 198772 121242 198784
rect 139486 198772 139492 198784
rect 139544 198772 139550 198824
rect 141142 198772 141148 198824
rect 141200 198812 141206 198824
rect 141694 198812 141700 198824
rect 141200 198784 141700 198812
rect 141200 198772 141206 198784
rect 141694 198772 141700 198784
rect 141752 198772 141758 198824
rect 143902 198772 143908 198824
rect 143960 198812 143966 198824
rect 144086 198812 144092 198824
rect 143960 198784 144092 198812
rect 143960 198772 143966 198784
rect 144086 198772 144092 198784
rect 144144 198772 144150 198824
rect 158070 198772 158076 198824
rect 158128 198812 158134 198824
rect 178770 198812 178776 198824
rect 158128 198784 178776 198812
rect 158128 198772 158134 198784
rect 178770 198772 178776 198784
rect 178828 198772 178834 198824
rect 185578 198812 185584 198824
rect 180996 198784 185584 198812
rect 129090 198704 129096 198756
rect 129148 198744 129154 198756
rect 149146 198744 149152 198756
rect 129148 198716 149152 198744
rect 129148 198704 129154 198716
rect 149146 198704 149152 198716
rect 149204 198704 149210 198756
rect 162578 198704 162584 198756
rect 162636 198744 162642 198756
rect 180996 198744 181024 198784
rect 185578 198772 185584 198784
rect 185636 198772 185642 198824
rect 162636 198716 181024 198744
rect 162636 198704 162642 198716
rect 181070 198704 181076 198756
rect 181128 198744 181134 198756
rect 187694 198744 187700 198756
rect 181128 198716 187700 198744
rect 181128 198704 181134 198716
rect 187694 198704 187700 198716
rect 187752 198704 187758 198756
rect 125870 198636 125876 198688
rect 125928 198676 125934 198688
rect 130746 198676 130752 198688
rect 125928 198648 130752 198676
rect 125928 198636 125934 198648
rect 130746 198636 130752 198648
rect 130804 198636 130810 198688
rect 132494 198636 132500 198688
rect 132552 198676 132558 198688
rect 146202 198676 146208 198688
rect 132552 198648 146208 198676
rect 132552 198636 132558 198648
rect 146202 198636 146208 198648
rect 146260 198636 146266 198688
rect 167454 198636 167460 198688
rect 167512 198676 167518 198688
rect 167512 198648 173802 198676
rect 167512 198636 167518 198648
rect 122190 198568 122196 198620
rect 122248 198608 122254 198620
rect 146846 198608 146852 198620
rect 122248 198580 146852 198608
rect 122248 198568 122254 198580
rect 146846 198568 146852 198580
rect 146904 198568 146910 198620
rect 164970 198568 164976 198620
rect 165028 198608 165034 198620
rect 167914 198608 167920 198620
rect 165028 198580 167920 198608
rect 165028 198568 165034 198580
rect 167914 198568 167920 198580
rect 167972 198568 167978 198620
rect 169938 198568 169944 198620
rect 169996 198608 170002 198620
rect 173774 198608 173802 198648
rect 173894 198636 173900 198688
rect 173952 198676 173958 198688
rect 202506 198676 202512 198688
rect 173952 198648 202512 198676
rect 173952 198636 173958 198648
rect 202506 198636 202512 198648
rect 202564 198636 202570 198688
rect 201586 198608 201592 198620
rect 169996 198580 173710 198608
rect 173774 198580 201592 198608
rect 169996 198568 170002 198580
rect 129274 198500 129280 198552
rect 129332 198540 129338 198552
rect 154666 198540 154672 198552
rect 129332 198512 154672 198540
rect 129332 198500 129338 198512
rect 154666 198500 154672 198512
rect 154724 198500 154730 198552
rect 158990 198500 158996 198552
rect 159048 198540 159054 198552
rect 165614 198540 165620 198552
rect 159048 198512 165620 198540
rect 159048 198500 159054 198512
rect 165614 198500 165620 198512
rect 165672 198500 165678 198552
rect 166442 198500 166448 198552
rect 166500 198540 166506 198552
rect 166810 198540 166816 198552
rect 166500 198512 166816 198540
rect 166500 198500 166506 198512
rect 166810 198500 166816 198512
rect 166868 198500 166874 198552
rect 172514 198540 172520 198552
rect 171520 198512 172520 198540
rect 105814 198432 105820 198484
rect 105872 198472 105878 198484
rect 132402 198472 132408 198484
rect 105872 198444 132408 198472
rect 105872 198432 105878 198444
rect 132402 198432 132408 198444
rect 132460 198432 132466 198484
rect 142430 198432 142436 198484
rect 142488 198472 142494 198484
rect 143902 198472 143908 198484
rect 142488 198444 143908 198472
rect 142488 198432 142494 198444
rect 143902 198432 143908 198444
rect 143960 198432 143966 198484
rect 159726 198432 159732 198484
rect 159784 198472 159790 198484
rect 171520 198472 171548 198512
rect 172514 198500 172520 198512
rect 172572 198500 172578 198552
rect 159784 198444 171548 198472
rect 173682 198472 173710 198580
rect 201586 198568 201592 198580
rect 201644 198568 201650 198620
rect 174354 198500 174360 198552
rect 174412 198540 174418 198552
rect 207106 198540 207112 198552
rect 174412 198512 207112 198540
rect 174412 198500 174418 198512
rect 207106 198500 207112 198512
rect 207164 198500 207170 198552
rect 208578 198472 208584 198484
rect 173682 198444 208584 198472
rect 159784 198432 159790 198444
rect 208578 198432 208584 198444
rect 208636 198432 208642 198484
rect 122282 198364 122288 198416
rect 122340 198404 122346 198416
rect 149422 198404 149428 198416
rect 122340 198376 149428 198404
rect 122340 198364 122346 198376
rect 149422 198364 149428 198376
rect 149480 198364 149486 198416
rect 165522 198364 165528 198416
rect 165580 198404 165586 198416
rect 171594 198404 171600 198416
rect 165580 198376 171600 198404
rect 165580 198364 165586 198376
rect 171594 198364 171600 198376
rect 171652 198364 171658 198416
rect 172054 198364 172060 198416
rect 172112 198404 172118 198416
rect 172112 198376 175596 198404
rect 172112 198364 172118 198376
rect 107102 198296 107108 198348
rect 107160 198336 107166 198348
rect 136082 198336 136088 198348
rect 107160 198308 136088 198336
rect 107160 198296 107166 198308
rect 136082 198296 136088 198308
rect 136140 198296 136146 198348
rect 163130 198296 163136 198348
rect 163188 198336 163194 198348
rect 171042 198336 171048 198348
rect 163188 198308 171048 198336
rect 163188 198296 163194 198308
rect 171042 198296 171048 198308
rect 171100 198296 171106 198348
rect 172422 198296 172428 198348
rect 172480 198336 172486 198348
rect 174814 198336 174820 198348
rect 172480 198308 174820 198336
rect 172480 198296 172486 198308
rect 174814 198296 174820 198308
rect 174872 198296 174878 198348
rect 175568 198336 175596 198376
rect 175642 198364 175648 198416
rect 175700 198404 175706 198416
rect 212810 198404 212816 198416
rect 175700 198376 212816 198404
rect 175700 198364 175706 198376
rect 212810 198364 212816 198376
rect 212868 198364 212874 198416
rect 211338 198336 211344 198348
rect 175568 198308 211344 198336
rect 211338 198296 211344 198308
rect 211396 198296 211402 198348
rect 110322 198228 110328 198280
rect 110380 198268 110386 198280
rect 143350 198268 143356 198280
rect 110380 198240 143356 198268
rect 110380 198228 110386 198240
rect 143350 198228 143356 198240
rect 143408 198228 143414 198280
rect 165706 198228 165712 198280
rect 165764 198268 165770 198280
rect 167454 198268 167460 198280
rect 165764 198240 167460 198268
rect 165764 198228 165770 198240
rect 167454 198228 167460 198240
rect 167512 198228 167518 198280
rect 170582 198228 170588 198280
rect 170640 198268 170646 198280
rect 209958 198268 209964 198280
rect 170640 198240 209964 198268
rect 170640 198228 170646 198240
rect 209958 198228 209964 198240
rect 210016 198228 210022 198280
rect 107194 198160 107200 198212
rect 107252 198200 107258 198212
rect 137002 198200 137008 198212
rect 107252 198172 137008 198200
rect 107252 198160 107258 198172
rect 137002 198160 137008 198172
rect 137060 198160 137066 198212
rect 155586 198160 155592 198212
rect 155644 198200 155650 198212
rect 171134 198200 171140 198212
rect 155644 198172 171140 198200
rect 155644 198160 155650 198172
rect 171134 198160 171140 198172
rect 171192 198160 171198 198212
rect 172790 198160 172796 198212
rect 172848 198200 172854 198212
rect 212902 198200 212908 198212
rect 172848 198172 212908 198200
rect 172848 198160 172854 198172
rect 212902 198160 212908 198172
rect 212960 198160 212966 198212
rect 110230 198092 110236 198144
rect 110288 198132 110294 198144
rect 144730 198132 144736 198144
rect 110288 198104 144736 198132
rect 110288 198092 110294 198104
rect 144730 198092 144736 198104
rect 144788 198092 144794 198144
rect 162762 198092 162768 198144
rect 162820 198132 162826 198144
rect 163314 198132 163320 198144
rect 162820 198104 163320 198132
rect 162820 198092 162826 198104
rect 163314 198092 163320 198104
rect 163372 198092 163378 198144
rect 165614 198092 165620 198144
rect 165672 198132 165678 198144
rect 172054 198132 172060 198144
rect 165672 198104 172060 198132
rect 165672 198092 165678 198104
rect 172054 198092 172060 198104
rect 172112 198092 172118 198144
rect 172330 198092 172336 198144
rect 172388 198132 172394 198144
rect 212718 198132 212724 198144
rect 172388 198104 212724 198132
rect 172388 198092 172394 198104
rect 212718 198092 212724 198104
rect 212776 198092 212782 198144
rect 108666 198024 108672 198076
rect 108724 198064 108730 198076
rect 142062 198064 142068 198076
rect 108724 198036 142068 198064
rect 108724 198024 108730 198036
rect 142062 198024 142068 198036
rect 142120 198024 142126 198076
rect 156598 198024 156604 198076
rect 156656 198064 156662 198076
rect 165706 198064 165712 198076
rect 156656 198036 165712 198064
rect 156656 198024 156662 198036
rect 165706 198024 165712 198036
rect 165764 198024 165770 198076
rect 166074 198024 166080 198076
rect 166132 198064 166138 198076
rect 166442 198064 166448 198076
rect 166132 198036 166448 198064
rect 166132 198024 166138 198036
rect 166442 198024 166448 198036
rect 166500 198024 166506 198076
rect 171318 198024 171324 198076
rect 171376 198064 171382 198076
rect 212994 198064 213000 198076
rect 171376 198036 213000 198064
rect 171376 198024 171382 198036
rect 212994 198024 213000 198036
rect 213052 198024 213058 198076
rect 126514 197956 126520 198008
rect 126572 197996 126578 198008
rect 132494 197996 132500 198008
rect 126572 197968 132500 197996
rect 126572 197956 126578 197968
rect 132494 197956 132500 197968
rect 132552 197956 132558 198008
rect 155310 197956 155316 198008
rect 155368 197996 155374 198008
rect 164970 197996 164976 198008
rect 155368 197968 164976 197996
rect 155368 197956 155374 197968
rect 164970 197956 164976 197968
rect 165028 197956 165034 198008
rect 165614 197956 165620 198008
rect 165672 197996 165678 198008
rect 165982 197996 165988 198008
rect 165672 197968 165988 197996
rect 165672 197956 165678 197968
rect 165982 197956 165988 197968
rect 166040 197956 166046 198008
rect 167454 197956 167460 198008
rect 167512 197996 167518 198008
rect 167512 197968 168880 197996
rect 167512 197956 167518 197968
rect 133874 197888 133880 197940
rect 133932 197928 133938 197940
rect 150710 197928 150716 197940
rect 133932 197900 150716 197928
rect 133932 197888 133938 197900
rect 150710 197888 150716 197900
rect 150768 197888 150774 197940
rect 154850 197888 154856 197940
rect 154908 197928 154914 197940
rect 168852 197928 168880 197968
rect 169294 197956 169300 198008
rect 169352 197996 169358 198008
rect 209774 197996 209780 198008
rect 169352 197968 209780 197996
rect 169352 197956 169358 197968
rect 209774 197956 209780 197968
rect 209832 197956 209838 198008
rect 170766 197928 170772 197940
rect 154908 197900 168512 197928
rect 168852 197900 170772 197928
rect 154908 197888 154914 197900
rect 127710 197820 127716 197872
rect 127768 197860 127774 197872
rect 144178 197860 144184 197872
rect 127768 197832 144184 197860
rect 127768 197820 127774 197832
rect 144178 197820 144184 197832
rect 144236 197820 144242 197872
rect 156506 197820 156512 197872
rect 156564 197860 156570 197872
rect 158070 197860 158076 197872
rect 156564 197832 158076 197860
rect 156564 197820 156570 197832
rect 158070 197820 158076 197832
rect 158128 197820 158134 197872
rect 159174 197820 159180 197872
rect 159232 197860 159238 197872
rect 161290 197860 161296 197872
rect 159232 197832 161296 197860
rect 159232 197820 159238 197832
rect 161290 197820 161296 197832
rect 161348 197820 161354 197872
rect 162946 197820 162952 197872
rect 163004 197860 163010 197872
rect 163222 197860 163228 197872
rect 163004 197832 163228 197860
rect 163004 197820 163010 197832
rect 163222 197820 163228 197832
rect 163280 197820 163286 197872
rect 167086 197820 167092 197872
rect 167144 197860 167150 197872
rect 167454 197860 167460 197872
rect 167144 197832 167460 197860
rect 167144 197820 167150 197832
rect 167454 197820 167460 197832
rect 167512 197820 167518 197872
rect 168484 197860 168512 197900
rect 170766 197888 170772 197900
rect 170824 197888 170830 197940
rect 171134 197888 171140 197940
rect 171192 197928 171198 197940
rect 172330 197928 172336 197940
rect 171192 197900 172336 197928
rect 171192 197888 171198 197900
rect 172330 197888 172336 197900
rect 172388 197888 172394 197940
rect 172606 197888 172612 197940
rect 172664 197928 172670 197940
rect 172882 197928 172888 197940
rect 172664 197900 172888 197928
rect 172664 197888 172670 197900
rect 172882 197888 172888 197900
rect 172940 197888 172946 197940
rect 177114 197888 177120 197940
rect 177172 197928 177178 197940
rect 177758 197928 177764 197940
rect 177172 197900 177764 197928
rect 177172 197888 177178 197900
rect 177758 197888 177764 197900
rect 177816 197888 177822 197940
rect 174630 197860 174636 197872
rect 168484 197832 174636 197860
rect 174630 197820 174636 197832
rect 174688 197820 174694 197872
rect 127802 197752 127808 197804
rect 127860 197792 127866 197804
rect 143534 197792 143540 197804
rect 127860 197764 143540 197792
rect 127860 197752 127866 197764
rect 143534 197752 143540 197764
rect 143592 197752 143598 197804
rect 172146 197792 172152 197804
rect 164896 197764 172152 197792
rect 97626 197684 97632 197736
rect 97684 197724 97690 197736
rect 97684 197696 128354 197724
rect 97684 197684 97690 197696
rect 128326 197588 128354 197696
rect 130654 197684 130660 197736
rect 130712 197724 130718 197736
rect 133874 197724 133880 197736
rect 130712 197696 133880 197724
rect 130712 197684 130718 197696
rect 133874 197684 133880 197696
rect 133932 197684 133938 197736
rect 131850 197616 131856 197668
rect 131908 197656 131914 197668
rect 136726 197656 136732 197668
rect 131908 197628 136732 197656
rect 131908 197616 131914 197628
rect 136726 197616 136732 197628
rect 136784 197616 136790 197668
rect 143534 197616 143540 197668
rect 143592 197656 143598 197668
rect 143718 197656 143724 197668
rect 143592 197628 143724 197656
rect 143592 197616 143598 197628
rect 143718 197616 143724 197628
rect 143776 197616 143782 197668
rect 148042 197616 148048 197668
rect 148100 197656 148106 197668
rect 148318 197656 148324 197668
rect 148100 197628 148324 197656
rect 148100 197616 148106 197628
rect 148318 197616 148324 197628
rect 148376 197616 148382 197668
rect 157518 197616 157524 197668
rect 157576 197656 157582 197668
rect 164896 197656 164924 197764
rect 172146 197752 172152 197764
rect 172204 197752 172210 197804
rect 172514 197752 172520 197804
rect 172572 197792 172578 197804
rect 178126 197792 178132 197804
rect 172572 197764 178132 197792
rect 172572 197752 172578 197764
rect 178126 197752 178132 197764
rect 178184 197752 178190 197804
rect 173066 197724 173072 197736
rect 157576 197628 164924 197656
rect 166506 197696 173072 197724
rect 157576 197616 157582 197628
rect 137646 197588 137652 197600
rect 128326 197560 137652 197588
rect 137646 197548 137652 197560
rect 137704 197548 137710 197600
rect 161842 197548 161848 197600
rect 161900 197588 161906 197600
rect 166506 197588 166534 197696
rect 173066 197684 173072 197696
rect 173124 197684 173130 197736
rect 168282 197616 168288 197668
rect 168340 197656 168346 197668
rect 179414 197656 179420 197668
rect 168340 197628 179420 197656
rect 168340 197616 168346 197628
rect 179414 197616 179420 197628
rect 179472 197616 179478 197668
rect 161900 197560 166534 197588
rect 161900 197548 161906 197560
rect 125134 197480 125140 197532
rect 125192 197520 125198 197532
rect 133322 197520 133328 197532
rect 125192 197492 133328 197520
rect 125192 197480 125198 197492
rect 133322 197480 133328 197492
rect 133380 197480 133386 197532
rect 156230 197480 156236 197532
rect 156288 197520 156294 197532
rect 159174 197520 159180 197532
rect 156288 197492 159180 197520
rect 156288 197480 156294 197492
rect 159174 197480 159180 197492
rect 159232 197480 159238 197532
rect 161290 197480 161296 197532
rect 161348 197520 161354 197532
rect 173802 197520 173808 197532
rect 161348 197492 173808 197520
rect 161348 197480 161354 197492
rect 173802 197480 173808 197492
rect 173860 197480 173866 197532
rect 132862 197412 132868 197464
rect 132920 197452 132926 197464
rect 133506 197452 133512 197464
rect 132920 197424 133512 197452
rect 132920 197412 132926 197424
rect 133506 197412 133512 197424
rect 133564 197412 133570 197464
rect 134242 197412 134248 197464
rect 134300 197452 134306 197464
rect 135162 197452 135168 197464
rect 134300 197424 135168 197452
rect 134300 197412 134306 197424
rect 135162 197412 135168 197424
rect 135220 197412 135226 197464
rect 145190 197412 145196 197464
rect 145248 197452 145254 197464
rect 149422 197452 149428 197464
rect 145248 197424 149428 197452
rect 145248 197412 145254 197424
rect 149422 197412 149428 197424
rect 149480 197412 149486 197464
rect 159542 197412 159548 197464
rect 159600 197452 159606 197464
rect 172422 197452 172428 197464
rect 159600 197424 172428 197452
rect 159600 197412 159606 197424
rect 172422 197412 172428 197424
rect 172480 197412 172486 197464
rect 173986 197412 173992 197464
rect 174044 197452 174050 197464
rect 178954 197452 178960 197464
rect 174044 197424 178960 197452
rect 174044 197412 174050 197424
rect 178954 197412 178960 197424
rect 179012 197412 179018 197464
rect 134150 197344 134156 197396
rect 134208 197384 134214 197396
rect 134610 197384 134616 197396
rect 134208 197356 134616 197384
rect 134208 197344 134214 197356
rect 134610 197344 134616 197356
rect 134668 197344 134674 197396
rect 143902 197344 143908 197396
rect 143960 197384 143966 197396
rect 144546 197384 144552 197396
rect 143960 197356 144552 197384
rect 143960 197344 143966 197356
rect 144546 197344 144552 197356
rect 144604 197344 144610 197396
rect 120994 197276 121000 197328
rect 121052 197316 121058 197328
rect 146754 197316 146760 197328
rect 121052 197288 146760 197316
rect 121052 197276 121058 197288
rect 146754 197276 146760 197288
rect 146812 197276 146818 197328
rect 155862 197276 155868 197328
rect 155920 197316 155926 197328
rect 165338 197316 165344 197328
rect 155920 197288 165344 197316
rect 155920 197276 155926 197288
rect 165338 197276 165344 197288
rect 165396 197276 165402 197328
rect 121086 197208 121092 197260
rect 121144 197248 121150 197260
rect 149882 197248 149888 197260
rect 121144 197220 149888 197248
rect 121144 197208 121150 197220
rect 149882 197208 149888 197220
rect 149940 197208 149946 197260
rect 163866 197208 163872 197260
rect 163924 197248 163930 197260
rect 171318 197248 171324 197260
rect 163924 197220 171324 197248
rect 163924 197208 163930 197220
rect 171318 197208 171324 197220
rect 171376 197208 171382 197260
rect 172054 197208 172060 197260
rect 172112 197248 172118 197260
rect 193398 197248 193404 197260
rect 172112 197220 193404 197248
rect 172112 197208 172118 197220
rect 193398 197208 193404 197220
rect 193456 197208 193462 197260
rect 114278 197140 114284 197192
rect 114336 197180 114342 197192
rect 144362 197180 144368 197192
rect 114336 197152 144368 197180
rect 114336 197140 114342 197152
rect 144362 197140 144368 197152
rect 144420 197140 144426 197192
rect 166902 197140 166908 197192
rect 166960 197180 166966 197192
rect 170398 197180 170404 197192
rect 166960 197152 170404 197180
rect 166960 197140 166966 197152
rect 170398 197140 170404 197152
rect 170456 197140 170462 197192
rect 171042 197140 171048 197192
rect 171100 197180 171106 197192
rect 194870 197180 194876 197192
rect 171100 197152 194876 197180
rect 171100 197140 171106 197152
rect 194870 197140 194876 197152
rect 194928 197140 194934 197192
rect 116854 197072 116860 197124
rect 116912 197112 116918 197124
rect 147582 197112 147588 197124
rect 116912 197084 147588 197112
rect 116912 197072 116918 197084
rect 147582 197072 147588 197084
rect 147640 197072 147646 197124
rect 157242 197072 157248 197124
rect 157300 197112 157306 197124
rect 158714 197112 158720 197124
rect 157300 197084 158720 197112
rect 157300 197072 157306 197084
rect 158714 197072 158720 197084
rect 158772 197072 158778 197124
rect 160830 197072 160836 197124
rect 160888 197112 160894 197124
rect 194594 197112 194600 197124
rect 160888 197084 194600 197112
rect 160888 197072 160894 197084
rect 194594 197072 194600 197084
rect 194652 197072 194658 197124
rect 107010 197004 107016 197056
rect 107068 197044 107074 197056
rect 137462 197044 137468 197056
rect 107068 197016 137468 197044
rect 107068 197004 107074 197016
rect 137462 197004 137468 197016
rect 137520 197004 137526 197056
rect 148502 197004 148508 197056
rect 148560 197044 148566 197056
rect 149790 197044 149796 197056
rect 148560 197016 149796 197044
rect 148560 197004 148566 197016
rect 149790 197004 149796 197016
rect 149848 197004 149854 197056
rect 167914 197004 167920 197056
rect 167972 197044 167978 197056
rect 198826 197044 198832 197056
rect 167972 197016 198832 197044
rect 167972 197004 167978 197016
rect 198826 197004 198832 197016
rect 198884 197004 198890 197056
rect 112714 196936 112720 196988
rect 112772 196976 112778 196988
rect 132954 196976 132960 196988
rect 112772 196948 132960 196976
rect 112772 196936 112778 196948
rect 132954 196936 132960 196948
rect 133012 196936 133018 196988
rect 140866 196936 140872 196988
rect 140924 196976 140930 196988
rect 141142 196976 141148 196988
rect 140924 196948 141148 196976
rect 140924 196936 140930 196948
rect 141142 196936 141148 196948
rect 141200 196936 141206 196988
rect 171594 196936 171600 196988
rect 171652 196976 171658 196988
rect 198918 196976 198924 196988
rect 171652 196948 198924 196976
rect 171652 196936 171658 196948
rect 198918 196936 198924 196948
rect 198976 196936 198982 196988
rect 111702 196868 111708 196920
rect 111760 196908 111766 196920
rect 143810 196908 143816 196920
rect 111760 196880 143816 196908
rect 111760 196868 111766 196880
rect 143810 196868 143816 196880
rect 143868 196868 143874 196920
rect 167178 196868 167184 196920
rect 167236 196908 167242 196920
rect 201678 196908 201684 196920
rect 167236 196880 201684 196908
rect 167236 196868 167242 196880
rect 201678 196868 201684 196880
rect 201736 196868 201742 196920
rect 114186 196800 114192 196852
rect 114244 196840 114250 196852
rect 147306 196840 147312 196852
rect 114244 196812 147312 196840
rect 114244 196800 114250 196812
rect 147306 196800 147312 196812
rect 147364 196800 147370 196852
rect 155954 196800 155960 196852
rect 156012 196840 156018 196852
rect 156012 196812 157334 196840
rect 156012 196800 156018 196812
rect 109862 196732 109868 196784
rect 109920 196772 109926 196784
rect 133230 196772 133236 196784
rect 109920 196744 133236 196772
rect 109920 196732 109926 196744
rect 133230 196732 133236 196744
rect 133288 196732 133294 196784
rect 146294 196732 146300 196784
rect 146352 196772 146358 196784
rect 146478 196772 146484 196784
rect 146352 196744 146484 196772
rect 146352 196732 146358 196744
rect 146478 196732 146484 196744
rect 146536 196732 146542 196784
rect 114462 196664 114468 196716
rect 114520 196704 114526 196716
rect 147674 196704 147680 196716
rect 114520 196676 147680 196704
rect 114520 196664 114526 196676
rect 147674 196664 147680 196676
rect 147732 196664 147738 196716
rect 105906 196596 105912 196648
rect 105964 196636 105970 196648
rect 138750 196636 138756 196648
rect 105964 196608 138756 196636
rect 105964 196596 105970 196608
rect 138750 196596 138756 196608
rect 138808 196596 138814 196648
rect 141878 196596 141884 196648
rect 141936 196636 141942 196648
rect 142246 196636 142252 196648
rect 141936 196608 142252 196636
rect 141936 196596 141942 196608
rect 142246 196596 142252 196608
rect 142304 196596 142310 196648
rect 157306 196636 157334 196812
rect 164142 196800 164148 196852
rect 164200 196840 164206 196852
rect 170582 196840 170588 196852
rect 164200 196812 170588 196840
rect 164200 196800 164206 196812
rect 170582 196800 170588 196812
rect 170640 196800 170646 196852
rect 171226 196800 171232 196852
rect 171284 196840 171290 196852
rect 171594 196840 171600 196852
rect 171284 196812 171600 196840
rect 171284 196800 171290 196812
rect 171594 196800 171600 196812
rect 171652 196800 171658 196852
rect 172514 196800 172520 196852
rect 172572 196840 172578 196852
rect 200482 196840 200488 196852
rect 172572 196812 200488 196840
rect 172572 196800 172578 196812
rect 200482 196800 200488 196812
rect 200540 196800 200546 196852
rect 163590 196732 163596 196784
rect 163648 196772 163654 196784
rect 197630 196772 197636 196784
rect 163648 196744 197636 196772
rect 163648 196732 163654 196744
rect 197630 196732 197636 196744
rect 197688 196732 197694 196784
rect 169846 196664 169852 196716
rect 169904 196704 169910 196716
rect 170214 196704 170220 196716
rect 169904 196676 170220 196704
rect 169904 196664 169910 196676
rect 170214 196664 170220 196676
rect 170272 196664 170278 196716
rect 170582 196664 170588 196716
rect 170640 196704 170646 196716
rect 197722 196704 197728 196716
rect 170640 196676 197728 196704
rect 170640 196664 170646 196676
rect 197722 196664 197728 196676
rect 197780 196664 197786 196716
rect 190638 196636 190644 196648
rect 157306 196608 190644 196636
rect 190638 196596 190644 196608
rect 190696 196596 190702 196648
rect 129458 196528 129464 196580
rect 129516 196568 129522 196580
rect 149974 196568 149980 196580
rect 129516 196540 149980 196568
rect 129516 196528 129522 196540
rect 149974 196528 149980 196540
rect 150032 196528 150038 196580
rect 158622 196528 158628 196580
rect 158680 196568 158686 196580
rect 160278 196568 160284 196580
rect 158680 196540 160284 196568
rect 158680 196528 158686 196540
rect 160278 196528 160284 196540
rect 160336 196528 160342 196580
rect 164694 196528 164700 196580
rect 164752 196568 164758 196580
rect 164878 196568 164884 196580
rect 164752 196540 164884 196568
rect 164752 196528 164758 196540
rect 164878 196528 164884 196540
rect 164936 196528 164942 196580
rect 171318 196528 171324 196580
rect 171376 196568 171382 196580
rect 179046 196568 179052 196580
rect 171376 196540 179052 196568
rect 171376 196528 171382 196540
rect 179046 196528 179052 196540
rect 179104 196528 179110 196580
rect 132770 196460 132776 196512
rect 132828 196500 132834 196512
rect 133782 196500 133788 196512
rect 132828 196472 133788 196500
rect 132828 196460 132834 196472
rect 133782 196460 133788 196472
rect 133840 196460 133846 196512
rect 134150 196460 134156 196512
rect 134208 196500 134214 196512
rect 135070 196500 135076 196512
rect 134208 196472 135076 196500
rect 134208 196460 134214 196472
rect 135070 196460 135076 196472
rect 135128 196460 135134 196512
rect 137278 196460 137284 196512
rect 137336 196500 137342 196512
rect 139394 196500 139400 196512
rect 137336 196472 139400 196500
rect 137336 196460 137342 196472
rect 139394 196460 139400 196472
rect 139452 196460 139458 196512
rect 131758 196392 131764 196444
rect 131816 196432 131822 196444
rect 139670 196432 139676 196444
rect 131816 196404 139676 196432
rect 131816 196392 131822 196404
rect 139670 196392 139676 196404
rect 139728 196392 139734 196444
rect 129366 196324 129372 196376
rect 129424 196364 129430 196376
rect 147858 196364 147864 196376
rect 129424 196336 147864 196364
rect 129424 196324 129430 196336
rect 147858 196324 147864 196336
rect 147916 196324 147922 196376
rect 167730 196324 167736 196376
rect 167788 196364 167794 196376
rect 180518 196364 180524 196376
rect 167788 196336 180524 196364
rect 167788 196324 167794 196336
rect 180518 196324 180524 196336
rect 180576 196324 180582 196376
rect 133230 196256 133236 196308
rect 133288 196296 133294 196308
rect 142798 196296 142804 196308
rect 133288 196268 142804 196296
rect 133288 196256 133294 196268
rect 142798 196256 142804 196268
rect 142856 196256 142862 196308
rect 132954 196188 132960 196240
rect 133012 196228 133018 196240
rect 144086 196228 144092 196240
rect 133012 196200 144092 196228
rect 133012 196188 133018 196200
rect 144086 196188 144092 196200
rect 144144 196188 144150 196240
rect 129734 196120 129740 196172
rect 129792 196160 129798 196172
rect 134702 196160 134708 196172
rect 129792 196132 134708 196160
rect 129792 196120 129798 196132
rect 134702 196120 134708 196132
rect 134760 196120 134766 196172
rect 176856 196064 177252 196092
rect 132126 195984 132132 196036
rect 132184 196024 132190 196036
rect 133138 196024 133144 196036
rect 132184 195996 133144 196024
rect 132184 195984 132190 195996
rect 133138 195984 133144 195996
rect 133196 195984 133202 196036
rect 134518 195984 134524 196036
rect 134576 196024 134582 196036
rect 134978 196024 134984 196036
rect 134576 195996 134984 196024
rect 134576 195984 134582 195996
rect 134978 195984 134984 195996
rect 135036 195984 135042 196036
rect 120626 195916 120632 195968
rect 120684 195956 120690 195968
rect 144822 195956 144828 195968
rect 120684 195928 144828 195956
rect 120684 195916 120690 195928
rect 144822 195916 144828 195928
rect 144880 195916 144886 195968
rect 152182 195916 152188 195968
rect 152240 195956 152246 195968
rect 152826 195956 152832 195968
rect 152240 195928 152832 195956
rect 152240 195916 152246 195928
rect 152826 195916 152832 195928
rect 152884 195916 152890 195968
rect 157794 195916 157800 195968
rect 157852 195956 157858 195968
rect 157852 195928 161014 195956
rect 157852 195916 157858 195928
rect 115198 195848 115204 195900
rect 115256 195888 115262 195900
rect 146110 195888 146116 195900
rect 115256 195860 146116 195888
rect 115256 195848 115262 195860
rect 146110 195848 146116 195860
rect 146168 195848 146174 195900
rect 154482 195848 154488 195900
rect 154540 195888 154546 195900
rect 154540 195860 157472 195888
rect 154540 195848 154546 195860
rect 114094 195780 114100 195832
rect 114152 195820 114158 195832
rect 145466 195820 145472 195832
rect 114152 195792 145472 195820
rect 114152 195780 114158 195792
rect 145466 195780 145472 195792
rect 145524 195780 145530 195832
rect 154758 195780 154764 195832
rect 154816 195820 154822 195832
rect 157444 195820 157472 195860
rect 159450 195848 159456 195900
rect 159508 195888 159514 195900
rect 159508 195860 160922 195888
rect 159508 195848 159514 195860
rect 154816 195792 157334 195820
rect 157444 195792 160048 195820
rect 154816 195780 154822 195792
rect 115750 195712 115756 195764
rect 115808 195752 115814 195764
rect 157306 195752 157334 195792
rect 157610 195752 157616 195764
rect 115808 195724 147674 195752
rect 157306 195724 157616 195752
rect 115808 195712 115814 195724
rect 109954 195644 109960 195696
rect 110012 195684 110018 195696
rect 143166 195684 143172 195696
rect 110012 195656 143172 195684
rect 110012 195644 110018 195656
rect 143166 195644 143172 195656
rect 143224 195644 143230 195696
rect 111610 195576 111616 195628
rect 111668 195616 111674 195628
rect 145834 195616 145840 195628
rect 111668 195588 145840 195616
rect 111668 195576 111674 195588
rect 145834 195576 145840 195588
rect 145892 195576 145898 195628
rect 108850 195508 108856 195560
rect 108908 195548 108914 195560
rect 143442 195548 143448 195560
rect 108908 195520 143448 195548
rect 108908 195508 108914 195520
rect 143442 195508 143448 195520
rect 143500 195508 143506 195560
rect 147646 195548 147674 195724
rect 157610 195712 157616 195724
rect 157668 195712 157674 195764
rect 160020 195684 160048 195792
rect 160894 195752 160922 195860
rect 160986 195820 161014 195928
rect 162118 195916 162124 195968
rect 162176 195956 162182 195968
rect 171870 195956 171876 195968
rect 162176 195928 171876 195956
rect 162176 195916 162182 195928
rect 171870 195916 171876 195928
rect 171928 195916 171934 195968
rect 173802 195916 173808 195968
rect 173860 195956 173866 195968
rect 176856 195956 176884 196064
rect 176930 195984 176936 196036
rect 176988 196024 176994 196036
rect 176988 195996 177160 196024
rect 176988 195984 176994 195996
rect 173860 195928 176884 195956
rect 173860 195916 173866 195928
rect 176194 195888 176200 195900
rect 166966 195860 176200 195888
rect 166966 195820 166994 195860
rect 176194 195848 176200 195860
rect 176252 195848 176258 195900
rect 177132 195888 177160 195996
rect 177224 195956 177252 196064
rect 192202 195956 192208 195968
rect 177224 195928 192208 195956
rect 192202 195916 192208 195928
rect 192260 195916 192266 195968
rect 198182 195888 198188 195900
rect 177132 195860 198188 195888
rect 198182 195848 198188 195860
rect 198240 195848 198246 195900
rect 160986 195792 166994 195820
rect 174998 195780 175004 195832
rect 175056 195820 175062 195832
rect 181346 195820 181352 195832
rect 175056 195792 181352 195820
rect 175056 195780 175062 195792
rect 181346 195780 181352 195792
rect 181404 195780 181410 195832
rect 174354 195752 174360 195764
rect 160894 195724 174360 195752
rect 174354 195712 174360 195724
rect 174412 195712 174418 195764
rect 176286 195712 176292 195764
rect 176344 195752 176350 195764
rect 201034 195752 201040 195764
rect 176344 195724 201040 195752
rect 176344 195712 176350 195724
rect 201034 195712 201040 195724
rect 201092 195712 201098 195764
rect 186590 195684 186596 195696
rect 160020 195656 186596 195684
rect 186590 195644 186596 195656
rect 186648 195644 186654 195696
rect 153930 195576 153936 195628
rect 153988 195616 153994 195628
rect 188706 195616 188712 195628
rect 153988 195588 188712 195616
rect 153988 195576 153994 195588
rect 188706 195576 188712 195588
rect 188764 195576 188770 195628
rect 148962 195548 148968 195560
rect 147646 195520 148968 195548
rect 148962 195508 148968 195520
rect 149020 195508 149026 195560
rect 151906 195508 151912 195560
rect 151964 195548 151970 195560
rect 152274 195548 152280 195560
rect 151964 195520 152280 195548
rect 151964 195508 151970 195520
rect 152274 195508 152280 195520
rect 152332 195508 152338 195560
rect 160462 195508 160468 195560
rect 160520 195548 160526 195560
rect 193306 195548 193312 195560
rect 160520 195520 193312 195548
rect 160520 195508 160526 195520
rect 193306 195508 193312 195520
rect 193364 195508 193370 195560
rect 104618 195440 104624 195492
rect 104676 195480 104682 195492
rect 132586 195480 132592 195492
rect 104676 195452 132592 195480
rect 104676 195440 104682 195452
rect 132586 195440 132592 195452
rect 132644 195440 132650 195492
rect 132678 195440 132684 195492
rect 132736 195480 132742 195492
rect 133414 195480 133420 195492
rect 132736 195452 133420 195480
rect 132736 195440 132742 195452
rect 133414 195440 133420 195452
rect 133472 195440 133478 195492
rect 135806 195440 135812 195492
rect 135864 195480 135870 195492
rect 136266 195480 136272 195492
rect 135864 195452 136272 195480
rect 135864 195440 135870 195452
rect 136266 195440 136272 195452
rect 136324 195440 136330 195492
rect 149330 195440 149336 195492
rect 149388 195480 149394 195492
rect 149974 195480 149980 195492
rect 149388 195452 149980 195480
rect 149388 195440 149394 195452
rect 149974 195440 149980 195452
rect 150032 195440 150038 195492
rect 150710 195440 150716 195492
rect 150768 195480 150774 195492
rect 151078 195480 151084 195492
rect 150768 195452 151084 195480
rect 150768 195440 150774 195452
rect 151078 195440 151084 195452
rect 151136 195440 151142 195492
rect 151998 195440 152004 195492
rect 152056 195480 152062 195492
rect 152458 195480 152464 195492
rect 152056 195452 152464 195480
rect 152056 195440 152062 195452
rect 152458 195440 152464 195452
rect 152516 195440 152522 195492
rect 156690 195440 156696 195492
rect 156748 195480 156754 195492
rect 156748 195452 157334 195480
rect 156748 195440 156754 195452
rect 111150 195372 111156 195424
rect 111208 195412 111214 195424
rect 145282 195412 145288 195424
rect 111208 195384 145288 195412
rect 111208 195372 111214 195384
rect 145282 195372 145288 195384
rect 145340 195372 145346 195424
rect 153470 195372 153476 195424
rect 153528 195412 153534 195424
rect 154206 195412 154212 195424
rect 153528 195384 154212 195412
rect 153528 195372 153534 195384
rect 154206 195372 154212 195384
rect 154264 195372 154270 195424
rect 157306 195412 157334 195452
rect 158070 195440 158076 195492
rect 158128 195480 158134 195492
rect 173250 195480 173256 195492
rect 158128 195452 173256 195480
rect 158128 195440 158134 195452
rect 173250 195440 173256 195452
rect 173308 195440 173314 195492
rect 181346 195440 181352 195492
rect 181404 195480 181410 195492
rect 208670 195480 208676 195492
rect 181404 195452 208676 195480
rect 181404 195440 181410 195452
rect 208670 195440 208676 195452
rect 208728 195440 208734 195492
rect 190546 195412 190552 195424
rect 157306 195384 190552 195412
rect 190546 195372 190552 195384
rect 190604 195372 190610 195424
rect 112806 195304 112812 195356
rect 112864 195344 112870 195356
rect 146294 195344 146300 195356
rect 112864 195316 146300 195344
rect 112864 195304 112870 195316
rect 146294 195304 146300 195316
rect 146352 195304 146358 195356
rect 149330 195304 149336 195356
rect 149388 195344 149394 195356
rect 149698 195344 149704 195356
rect 149388 195316 149704 195344
rect 149388 195304 149394 195316
rect 149698 195304 149704 195316
rect 149756 195304 149762 195356
rect 150618 195304 150624 195356
rect 150676 195344 150682 195356
rect 151078 195344 151084 195356
rect 150676 195316 151084 195344
rect 150676 195304 150682 195316
rect 151078 195304 151084 195316
rect 151136 195304 151142 195356
rect 153562 195304 153568 195356
rect 153620 195344 153626 195356
rect 154298 195344 154304 195356
rect 153620 195316 154304 195344
rect 153620 195304 153626 195316
rect 154298 195304 154304 195316
rect 154356 195304 154362 195356
rect 188430 195344 188436 195356
rect 157306 195316 188436 195344
rect 111334 195236 111340 195288
rect 111392 195276 111398 195288
rect 145006 195276 145012 195288
rect 111392 195248 145012 195276
rect 111392 195236 111398 195248
rect 145006 195236 145012 195248
rect 145064 195236 145070 195288
rect 149054 195236 149060 195288
rect 149112 195276 149118 195288
rect 149514 195276 149520 195288
rect 149112 195248 149520 195276
rect 149112 195236 149118 195248
rect 149514 195236 149520 195248
rect 149572 195236 149578 195288
rect 150526 195236 150532 195288
rect 150584 195276 150590 195288
rect 150894 195276 150900 195288
rect 150584 195248 150900 195276
rect 150584 195236 150590 195248
rect 150894 195236 150900 195248
rect 150952 195236 150958 195288
rect 151262 195236 151268 195288
rect 151320 195276 151326 195288
rect 151630 195276 151636 195288
rect 151320 195248 151636 195276
rect 151320 195236 151326 195248
rect 151630 195236 151636 195248
rect 151688 195236 151694 195288
rect 153470 195236 153476 195288
rect 153528 195276 153534 195288
rect 154022 195276 154028 195288
rect 153528 195248 154028 195276
rect 153528 195236 153534 195248
rect 154022 195236 154028 195248
rect 154080 195236 154086 195288
rect 155954 195236 155960 195288
rect 156012 195276 156018 195288
rect 156874 195276 156880 195288
rect 156012 195248 156880 195276
rect 156012 195236 156018 195248
rect 156874 195236 156880 195248
rect 156932 195236 156938 195288
rect 126698 195168 126704 195220
rect 126756 195208 126762 195220
rect 145742 195208 145748 195220
rect 126756 195180 145748 195208
rect 126756 195168 126762 195180
rect 145742 195168 145748 195180
rect 145800 195168 145806 195220
rect 153286 195168 153292 195220
rect 153344 195208 153350 195220
rect 153838 195208 153844 195220
rect 153344 195180 153844 195208
rect 153344 195168 153350 195180
rect 153838 195168 153844 195180
rect 153896 195168 153902 195220
rect 154114 195168 154120 195220
rect 154172 195208 154178 195220
rect 157306 195208 157334 195316
rect 188430 195304 188436 195316
rect 188488 195304 188494 195356
rect 157610 195236 157616 195288
rect 157668 195276 157674 195288
rect 162118 195276 162124 195288
rect 157668 195248 162124 195276
rect 157668 195236 157674 195248
rect 162118 195236 162124 195248
rect 162176 195236 162182 195288
rect 211522 195276 211528 195288
rect 166966 195248 211528 195276
rect 154172 195180 157334 195208
rect 154172 195168 154178 195180
rect 130378 195100 130384 195152
rect 130436 195140 130442 195152
rect 147214 195140 147220 195152
rect 130436 195112 147220 195140
rect 130436 195100 130442 195112
rect 147214 195100 147220 195112
rect 147272 195100 147278 195152
rect 152366 195100 152372 195152
rect 152424 195140 152430 195152
rect 153102 195140 153108 195152
rect 152424 195112 153108 195140
rect 152424 195100 152430 195112
rect 153102 195100 153108 195112
rect 153160 195100 153166 195152
rect 153378 195100 153384 195152
rect 153436 195140 153442 195152
rect 154390 195140 154396 195152
rect 153436 195112 154396 195140
rect 153436 195100 153442 195112
rect 154390 195100 154396 195112
rect 154448 195100 154454 195152
rect 155402 195100 155408 195152
rect 155460 195140 155466 195152
rect 155678 195140 155684 195152
rect 155460 195112 155684 195140
rect 155460 195100 155466 195112
rect 155678 195100 155684 195112
rect 155736 195100 155742 195152
rect 135530 195032 135536 195084
rect 135588 195072 135594 195084
rect 136082 195072 136088 195084
rect 135588 195044 136088 195072
rect 135588 195032 135594 195044
rect 136082 195032 136088 195044
rect 136140 195032 136146 195084
rect 136726 195032 136732 195084
rect 136784 195072 136790 195084
rect 137462 195072 137468 195084
rect 136784 195044 137468 195072
rect 136784 195032 136790 195044
rect 137462 195032 137468 195044
rect 137520 195032 137526 195084
rect 135714 194964 135720 195016
rect 135772 195004 135778 195016
rect 136450 195004 136456 195016
rect 135772 194976 136456 195004
rect 135772 194964 135778 194976
rect 136450 194964 136456 194976
rect 136508 194964 136514 195016
rect 152826 194964 152832 195016
rect 152884 195004 152890 195016
rect 166966 195004 166994 195248
rect 211522 195236 211528 195248
rect 211580 195236 211586 195288
rect 190086 195208 190092 195220
rect 186286 195180 190092 195208
rect 169570 195100 169576 195152
rect 169628 195140 169634 195152
rect 182910 195140 182916 195152
rect 169628 195112 182916 195140
rect 169628 195100 169634 195112
rect 182910 195100 182916 195112
rect 182968 195100 182974 195152
rect 152884 194976 166994 195004
rect 152884 194964 152890 194976
rect 172606 194964 172612 195016
rect 172664 195004 172670 195016
rect 172974 195004 172980 195016
rect 172664 194976 172980 195004
rect 172664 194964 172670 194976
rect 172974 194964 172980 194976
rect 173032 194964 173038 195016
rect 139302 194936 139308 194948
rect 133800 194908 139308 194936
rect 131942 194828 131948 194880
rect 132000 194868 132006 194880
rect 133800 194868 133828 194908
rect 139302 194896 139308 194908
rect 139360 194896 139366 194948
rect 172330 194896 172336 194948
rect 172388 194936 172394 194948
rect 186286 194936 186314 195180
rect 190086 195168 190092 195180
rect 190144 195168 190150 195220
rect 172388 194908 186314 194936
rect 172388 194896 172394 194908
rect 132000 194840 133828 194868
rect 132000 194828 132006 194840
rect 135438 194828 135444 194880
rect 135496 194868 135502 194880
rect 136358 194868 136364 194880
rect 135496 194840 136364 194868
rect 135496 194828 135502 194840
rect 136358 194828 136364 194840
rect 136416 194828 136422 194880
rect 171870 194828 171876 194880
rect 171928 194868 171934 194880
rect 179138 194868 179144 194880
rect 171928 194840 179144 194868
rect 171928 194828 171934 194840
rect 179138 194828 179144 194840
rect 179196 194828 179202 194880
rect 132586 194760 132592 194812
rect 132644 194800 132650 194812
rect 139118 194800 139124 194812
rect 132644 194772 139124 194800
rect 132644 194760 132650 194772
rect 139118 194760 139124 194772
rect 139176 194760 139182 194812
rect 126238 194692 126244 194744
rect 126296 194732 126302 194744
rect 131114 194732 131120 194744
rect 126296 194704 131120 194732
rect 126296 194692 126302 194704
rect 131114 194692 131120 194704
rect 131172 194692 131178 194744
rect 122098 194488 122104 194540
rect 122156 194528 122162 194540
rect 148042 194528 148048 194540
rect 122156 194500 148048 194528
rect 122156 194488 122162 194500
rect 148042 194488 148048 194500
rect 148100 194488 148106 194540
rect 168650 194488 168656 194540
rect 168708 194528 168714 194540
rect 202874 194528 202880 194540
rect 168708 194500 202880 194528
rect 168708 194488 168714 194500
rect 202874 194488 202880 194500
rect 202932 194488 202938 194540
rect 103330 194420 103336 194472
rect 103388 194460 103394 194472
rect 127894 194460 127900 194472
rect 103388 194432 127900 194460
rect 103388 194420 103394 194432
rect 127894 194420 127900 194432
rect 127952 194420 127958 194472
rect 135346 194420 135352 194472
rect 135404 194460 135410 194472
rect 136174 194460 136180 194472
rect 135404 194432 136180 194460
rect 135404 194420 135410 194432
rect 136174 194420 136180 194432
rect 136232 194420 136238 194472
rect 169110 194420 169116 194472
rect 169168 194460 169174 194472
rect 202966 194460 202972 194472
rect 169168 194432 202972 194460
rect 169168 194420 169174 194432
rect 202966 194420 202972 194432
rect 203024 194420 203030 194472
rect 102962 194352 102968 194404
rect 103020 194392 103026 194404
rect 134886 194392 134892 194404
rect 103020 194364 134892 194392
rect 103020 194352 103026 194364
rect 134886 194352 134892 194364
rect 134944 194352 134950 194404
rect 168466 194352 168472 194404
rect 168524 194392 168530 194404
rect 168650 194392 168656 194404
rect 168524 194364 168656 194392
rect 168524 194352 168530 194364
rect 168650 194352 168656 194364
rect 168708 194352 168714 194404
rect 173526 194352 173532 194404
rect 173584 194392 173590 194404
rect 207198 194392 207204 194404
rect 173584 194364 207204 194392
rect 173584 194352 173590 194364
rect 207198 194352 207204 194364
rect 207256 194352 207262 194404
rect 103238 194284 103244 194336
rect 103296 194324 103302 194336
rect 124766 194324 124772 194336
rect 103296 194296 124772 194324
rect 103296 194284 103302 194296
rect 124766 194284 124772 194296
rect 124824 194284 124830 194336
rect 174538 194284 174544 194336
rect 174596 194324 174602 194336
rect 208486 194324 208492 194336
rect 174596 194296 208492 194324
rect 174596 194284 174602 194296
rect 208486 194284 208492 194296
rect 208544 194284 208550 194336
rect 107378 194216 107384 194268
rect 107436 194256 107442 194268
rect 140038 194256 140044 194268
rect 107436 194228 140044 194256
rect 107436 194216 107442 194228
rect 140038 194216 140044 194228
rect 140096 194216 140102 194268
rect 175458 194216 175464 194268
rect 175516 194256 175522 194268
rect 210142 194256 210148 194268
rect 175516 194228 210148 194256
rect 175516 194216 175522 194228
rect 210142 194216 210148 194228
rect 210200 194216 210206 194268
rect 108942 194148 108948 194200
rect 109000 194188 109006 194200
rect 143074 194188 143080 194200
rect 109000 194160 143080 194188
rect 109000 194148 109006 194160
rect 143074 194148 143080 194160
rect 143132 194148 143138 194200
rect 177850 194148 177856 194200
rect 177908 194188 177914 194200
rect 211614 194188 211620 194200
rect 177908 194160 211620 194188
rect 177908 194148 177914 194160
rect 211614 194148 211620 194160
rect 211672 194148 211678 194200
rect 110138 194080 110144 194132
rect 110196 194120 110202 194132
rect 143534 194120 143540 194132
rect 110196 194092 143540 194120
rect 110196 194080 110202 194092
rect 143534 194080 143540 194092
rect 143592 194080 143598 194132
rect 163958 194080 163964 194132
rect 164016 194120 164022 194132
rect 164142 194120 164148 194132
rect 164016 194092 164148 194120
rect 164016 194080 164022 194092
rect 164142 194080 164148 194092
rect 164200 194080 164206 194132
rect 170674 194080 170680 194132
rect 170732 194120 170738 194132
rect 204714 194120 204720 194132
rect 170732 194092 204720 194120
rect 170732 194080 170738 194092
rect 204714 194080 204720 194092
rect 204772 194080 204778 194132
rect 105722 194012 105728 194064
rect 105780 194052 105786 194064
rect 140406 194052 140412 194064
rect 105780 194024 140412 194052
rect 105780 194012 105786 194024
rect 140406 194012 140412 194024
rect 140464 194012 140470 194064
rect 172790 194012 172796 194064
rect 172848 194052 172854 194064
rect 207474 194052 207480 194064
rect 172848 194024 207480 194052
rect 172848 194012 172854 194024
rect 207474 194012 207480 194024
rect 207532 194012 207538 194064
rect 104250 193944 104256 193996
rect 104308 193984 104314 193996
rect 139026 193984 139032 193996
rect 104308 193956 139032 193984
rect 104308 193944 104314 193956
rect 139026 193944 139032 193956
rect 139084 193944 139090 193996
rect 157426 193944 157432 193996
rect 157484 193984 157490 193996
rect 157886 193984 157892 193996
rect 157484 193956 157892 193984
rect 157484 193944 157490 193956
rect 157886 193944 157892 193956
rect 157944 193944 157950 193996
rect 174262 193944 174268 193996
rect 174320 193984 174326 193996
rect 208854 193984 208860 193996
rect 174320 193956 208860 193984
rect 174320 193944 174326 193956
rect 208854 193944 208860 193956
rect 208912 193944 208918 193996
rect 97902 193876 97908 193928
rect 97960 193916 97966 193928
rect 141326 193916 141332 193928
rect 97960 193888 141332 193916
rect 97960 193876 97966 193888
rect 141326 193876 141332 193888
rect 141384 193876 141390 193928
rect 150710 193876 150716 193928
rect 150768 193916 150774 193928
rect 151170 193916 151176 193928
rect 150768 193888 151176 193916
rect 150768 193876 150774 193888
rect 151170 193876 151176 193888
rect 151228 193876 151234 193928
rect 157306 193888 167132 193916
rect 97810 193808 97816 193860
rect 97868 193848 97874 193860
rect 143902 193848 143908 193860
rect 97868 193820 143908 193848
rect 97868 193808 97874 193820
rect 143902 193808 143908 193820
rect 143960 193808 143966 193860
rect 155494 193808 155500 193860
rect 155552 193848 155558 193860
rect 157306 193848 157334 193888
rect 155552 193820 157334 193848
rect 167104 193848 167132 193888
rect 169726 193888 171916 193916
rect 169726 193848 169754 193888
rect 167104 193820 169754 193848
rect 171888 193848 171916 193888
rect 174538 193876 174544 193928
rect 174596 193916 174602 193928
rect 174596 193888 179644 193916
rect 174596 193876 174602 193888
rect 179616 193848 179644 193888
rect 181346 193876 181352 193928
rect 181404 193916 181410 193928
rect 208946 193916 208952 193928
rect 181404 193888 208952 193916
rect 181404 193876 181410 193888
rect 208946 193876 208952 193888
rect 209004 193876 209010 193928
rect 183186 193848 183192 193860
rect 171888 193820 179414 193848
rect 179616 193820 183192 193848
rect 155552 193808 155558 193820
rect 155034 193740 155040 193792
rect 155092 193780 155098 193792
rect 174538 193780 174544 193792
rect 155092 193752 174544 193780
rect 155092 193740 155098 193752
rect 174538 193740 174544 193752
rect 174596 193740 174602 193792
rect 175274 193740 175280 193792
rect 175332 193780 175338 193792
rect 175734 193780 175740 193792
rect 175332 193752 175740 193780
rect 175332 193740 175338 193752
rect 175734 193740 175740 193752
rect 175792 193740 175798 193792
rect 179386 193780 179414 193820
rect 183186 193808 183192 193820
rect 183244 193808 183250 193860
rect 216766 193848 216772 193860
rect 190426 193820 216772 193848
rect 190426 193780 190454 193820
rect 216766 193808 216772 193820
rect 216824 193808 216830 193860
rect 179386 193752 190454 193780
rect 153194 193672 153200 193724
rect 153252 193712 153258 193724
rect 181530 193712 181536 193724
rect 153252 193684 181536 193712
rect 153252 193672 153258 193684
rect 181530 193672 181536 193684
rect 181588 193672 181594 193724
rect 156046 193604 156052 193656
rect 156104 193644 156110 193656
rect 181622 193644 181628 193656
rect 156104 193616 181628 193644
rect 156104 193604 156110 193616
rect 181622 193604 181628 193616
rect 181680 193604 181686 193656
rect 173986 193536 173992 193588
rect 174044 193576 174050 193588
rect 181346 193576 181352 193588
rect 174044 193548 181352 193576
rect 174044 193536 174050 193548
rect 181346 193536 181352 193548
rect 181404 193536 181410 193588
rect 130562 193128 130568 193180
rect 130620 193168 130626 193180
rect 148686 193168 148692 193180
rect 130620 193140 148692 193168
rect 130620 193128 130626 193140
rect 148686 193128 148692 193140
rect 148744 193128 148750 193180
rect 160462 193128 160468 193180
rect 160520 193168 160526 193180
rect 160646 193168 160652 193180
rect 160520 193140 160652 193168
rect 160520 193128 160526 193140
rect 160646 193128 160652 193140
rect 160704 193128 160710 193180
rect 176654 193128 176660 193180
rect 176712 193168 176718 193180
rect 177022 193168 177028 193180
rect 176712 193140 177028 193168
rect 176712 193128 176718 193140
rect 177022 193128 177028 193140
rect 177080 193128 177086 193180
rect 188338 193128 188344 193180
rect 188396 193168 188402 193180
rect 580166 193168 580172 193180
rect 188396 193140 580172 193168
rect 188396 193128 188402 193140
rect 580166 193128 580172 193140
rect 580224 193128 580230 193180
rect 102778 193060 102784 193112
rect 102836 193100 102842 193112
rect 129734 193100 129740 193112
rect 102836 193072 129740 193100
rect 102836 193060 102842 193072
rect 129734 193060 129740 193072
rect 129792 193060 129798 193112
rect 170306 193060 170312 193112
rect 170364 193100 170370 193112
rect 204438 193100 204444 193112
rect 170364 193072 204444 193100
rect 170364 193060 170370 193072
rect 204438 193060 204444 193072
rect 204496 193060 204502 193112
rect 101674 192992 101680 193044
rect 101732 193032 101738 193044
rect 130930 193032 130936 193044
rect 101732 193004 130936 193032
rect 101732 192992 101738 193004
rect 130930 192992 130936 193004
rect 130988 192992 130994 193044
rect 171594 192992 171600 193044
rect 171652 193032 171658 193044
rect 205910 193032 205916 193044
rect 171652 193004 205916 193032
rect 171652 192992 171658 193004
rect 205910 192992 205916 193004
rect 205968 192992 205974 193044
rect 117038 192924 117044 192976
rect 117096 192964 117102 192976
rect 146938 192964 146944 192976
rect 117096 192936 146944 192964
rect 117096 192924 117102 192936
rect 146938 192924 146944 192936
rect 146996 192924 147002 192976
rect 171502 192924 171508 192976
rect 171560 192964 171566 192976
rect 206002 192964 206008 192976
rect 171560 192936 206008 192964
rect 171560 192924 171566 192936
rect 206002 192924 206008 192936
rect 206060 192924 206066 192976
rect 108758 192856 108764 192908
rect 108816 192896 108822 192908
rect 140590 192896 140596 192908
rect 108816 192868 140596 192896
rect 108816 192856 108822 192868
rect 140590 192856 140596 192868
rect 140648 192856 140654 192908
rect 170214 192856 170220 192908
rect 170272 192896 170278 192908
rect 204622 192896 204628 192908
rect 170272 192868 204628 192896
rect 170272 192856 170278 192868
rect 204622 192856 204628 192868
rect 204680 192856 204686 192908
rect 115106 192788 115112 192840
rect 115164 192828 115170 192840
rect 147490 192828 147496 192840
rect 115164 192800 147496 192828
rect 115164 192788 115170 192800
rect 147490 192788 147496 192800
rect 147548 192788 147554 192840
rect 172698 192788 172704 192840
rect 172756 192828 172762 192840
rect 207566 192828 207572 192840
rect 172756 192800 207572 192828
rect 172756 192788 172762 192800
rect 207566 192788 207572 192800
rect 207624 192788 207630 192840
rect 116210 192720 116216 192772
rect 116268 192760 116274 192772
rect 150066 192760 150072 192772
rect 116268 192732 150072 192760
rect 116268 192720 116274 192732
rect 150066 192720 150072 192732
rect 150124 192720 150130 192772
rect 173158 192720 173164 192772
rect 173216 192760 173222 192772
rect 207658 192760 207664 192772
rect 173216 192732 207664 192760
rect 173216 192720 173222 192732
rect 207658 192720 207664 192732
rect 207716 192720 207722 192772
rect 123938 192652 123944 192704
rect 123996 192692 124002 192704
rect 157150 192692 157156 192704
rect 123996 192664 157156 192692
rect 123996 192652 124002 192664
rect 157150 192652 157156 192664
rect 157208 192652 157214 192704
rect 160830 192652 160836 192704
rect 160888 192692 160894 192704
rect 208762 192692 208768 192704
rect 160888 192664 208768 192692
rect 160888 192652 160894 192664
rect 208762 192652 208768 192664
rect 208820 192652 208826 192704
rect 99098 192584 99104 192636
rect 99156 192624 99162 192636
rect 133322 192624 133328 192636
rect 99156 192596 133328 192624
rect 99156 192584 99162 192596
rect 133322 192584 133328 192596
rect 133380 192584 133386 192636
rect 159174 192584 159180 192636
rect 159232 192624 159238 192636
rect 211246 192624 211252 192636
rect 159232 192596 211252 192624
rect 159232 192584 159238 192596
rect 211246 192584 211252 192596
rect 211304 192584 211310 192636
rect 108298 192516 108304 192568
rect 108356 192556 108362 192568
rect 142890 192556 142896 192568
rect 108356 192528 142896 192556
rect 108356 192516 108362 192528
rect 142890 192516 142896 192528
rect 142948 192516 142954 192568
rect 157978 192516 157984 192568
rect 158036 192556 158042 192568
rect 211154 192556 211160 192568
rect 158036 192528 211160 192556
rect 158036 192516 158042 192528
rect 211154 192516 211160 192528
rect 211212 192516 211218 192568
rect 108390 192448 108396 192500
rect 108448 192488 108454 192500
rect 142614 192488 142620 192500
rect 108448 192460 142620 192488
rect 108448 192448 108454 192460
rect 142614 192448 142620 192460
rect 142672 192448 142678 192500
rect 155770 192448 155776 192500
rect 155828 192488 155834 192500
rect 210694 192488 210700 192500
rect 155828 192460 210700 192488
rect 155828 192448 155834 192460
rect 210694 192448 210700 192460
rect 210752 192448 210758 192500
rect 130838 192380 130844 192432
rect 130896 192420 130902 192432
rect 148502 192420 148508 192432
rect 130896 192392 148508 192420
rect 130896 192380 130902 192392
rect 148502 192380 148508 192392
rect 148560 192380 148566 192432
rect 174814 192380 174820 192432
rect 174872 192420 174878 192432
rect 205634 192420 205640 192432
rect 174872 192392 205640 192420
rect 174872 192380 174878 192392
rect 205634 192380 205640 192392
rect 205692 192380 205698 192432
rect 162578 192312 162584 192364
rect 162636 192352 162642 192364
rect 191098 192352 191104 192364
rect 162636 192324 191104 192352
rect 162636 192312 162642 192324
rect 191098 192312 191104 192324
rect 191156 192312 191162 192364
rect 177942 192244 177948 192296
rect 178000 192284 178006 192296
rect 189166 192284 189172 192296
rect 178000 192256 189172 192284
rect 178000 192244 178006 192256
rect 189166 192244 189172 192256
rect 189224 192244 189230 192296
rect 162670 192176 162676 192228
rect 162728 192216 162734 192228
rect 162946 192216 162952 192228
rect 162728 192188 162952 192216
rect 162728 192176 162734 192188
rect 162946 192176 162952 192188
rect 163004 192176 163010 192228
rect 137002 192108 137008 192160
rect 137060 192148 137066 192160
rect 137922 192148 137928 192160
rect 137060 192120 137928 192148
rect 137060 192108 137066 192120
rect 137922 192108 137928 192120
rect 137980 192108 137986 192160
rect 167362 191768 167368 191820
rect 167420 191808 167426 191820
rect 201494 191808 201500 191820
rect 167420 191780 201500 191808
rect 167420 191768 167426 191780
rect 201494 191768 201500 191780
rect 201552 191768 201558 191820
rect 166074 191700 166080 191752
rect 166132 191740 166138 191752
rect 166902 191740 166908 191752
rect 166132 191712 166908 191740
rect 166132 191700 166138 191712
rect 166902 191700 166908 191712
rect 166960 191700 166966 191752
rect 168558 191700 168564 191752
rect 168616 191740 168622 191752
rect 168616 191712 175044 191740
rect 168616 191700 168622 191712
rect 159266 191632 159272 191684
rect 159324 191672 159330 191684
rect 166626 191672 166632 191684
rect 159324 191644 166632 191672
rect 159324 191632 159330 191644
rect 166626 191632 166632 191644
rect 166684 191632 166690 191684
rect 173894 191632 173900 191684
rect 173952 191672 173958 191684
rect 174906 191672 174912 191684
rect 173952 191644 174912 191672
rect 173952 191632 173958 191644
rect 174906 191632 174912 191644
rect 174964 191632 174970 191684
rect 175016 191672 175044 191712
rect 175090 191700 175096 191752
rect 175148 191740 175154 191752
rect 201770 191740 201776 191752
rect 175148 191712 201776 191740
rect 175148 191700 175154 191712
rect 201770 191700 201776 191712
rect 201828 191700 201834 191752
rect 203242 191672 203248 191684
rect 175016 191644 203248 191672
rect 203242 191632 203248 191644
rect 203300 191632 203306 191684
rect 163774 191564 163780 191616
rect 163832 191604 163838 191616
rect 204346 191604 204352 191616
rect 163832 191576 204352 191604
rect 163832 191564 163838 191576
rect 204346 191564 204352 191576
rect 204404 191564 204410 191616
rect 142430 191496 142436 191548
rect 142488 191536 142494 191548
rect 142982 191536 142988 191548
rect 142488 191508 142988 191536
rect 142488 191496 142494 191508
rect 142982 191496 142988 191508
rect 143040 191496 143046 191548
rect 164694 191496 164700 191548
rect 164752 191536 164758 191548
rect 205726 191536 205732 191548
rect 164752 191508 205732 191536
rect 164752 191496 164758 191508
rect 205726 191496 205732 191508
rect 205784 191496 205790 191548
rect 122466 191428 122472 191480
rect 122524 191468 122530 191480
rect 151446 191468 151452 191480
rect 122524 191440 151452 191468
rect 122524 191428 122530 191440
rect 151446 191428 151452 191440
rect 151504 191428 151510 191480
rect 159910 191428 159916 191480
rect 159968 191468 159974 191480
rect 159968 191440 161520 191468
rect 159968 191428 159974 191440
rect 106090 191360 106096 191412
rect 106148 191400 106154 191412
rect 137738 191400 137744 191412
rect 106148 191372 137744 191400
rect 106148 191360 106154 191372
rect 137738 191360 137744 191372
rect 137796 191360 137802 191412
rect 159358 191360 159364 191412
rect 159416 191400 159422 191412
rect 159416 191372 161428 191400
rect 159416 191360 159422 191372
rect 108574 191292 108580 191344
rect 108632 191332 108638 191344
rect 141234 191332 141240 191344
rect 108632 191304 141240 191332
rect 108632 191292 108638 191304
rect 141234 191292 141240 191304
rect 141292 191292 141298 191344
rect 104158 191224 104164 191276
rect 104216 191264 104222 191276
rect 137554 191264 137560 191276
rect 104216 191236 137560 191264
rect 104216 191224 104222 191236
rect 137554 191224 137560 191236
rect 137612 191224 137618 191276
rect 142522 191224 142528 191276
rect 142580 191264 142586 191276
rect 142982 191264 142988 191276
rect 142580 191236 142988 191264
rect 142580 191224 142586 191236
rect 142982 191224 142988 191236
rect 143040 191224 143046 191276
rect 160278 191224 160284 191276
rect 160336 191264 160342 191276
rect 161290 191264 161296 191276
rect 160336 191236 161296 191264
rect 160336 191224 160342 191236
rect 161290 191224 161296 191236
rect 161348 191224 161354 191276
rect 161400 191264 161428 191372
rect 161492 191332 161520 191440
rect 166534 191428 166540 191480
rect 166592 191468 166598 191480
rect 207382 191468 207388 191480
rect 166592 191440 207388 191468
rect 166592 191428 166598 191440
rect 207382 191428 207388 191440
rect 207440 191428 207446 191480
rect 167178 191360 167184 191412
rect 167236 191400 167242 191412
rect 167546 191400 167552 191412
rect 167236 191372 167552 191400
rect 167236 191360 167242 191372
rect 167546 191360 167552 191372
rect 167604 191360 167610 191412
rect 174170 191360 174176 191412
rect 174228 191400 174234 191412
rect 174722 191400 174728 191412
rect 174228 191372 174728 191400
rect 174228 191360 174234 191372
rect 174722 191360 174728 191372
rect 174780 191360 174786 191412
rect 174998 191360 175004 191412
rect 175056 191400 175062 191412
rect 209038 191400 209044 191412
rect 175056 191372 209044 191400
rect 175056 191360 175062 191372
rect 209038 191360 209044 191372
rect 209096 191360 209102 191412
rect 207290 191332 207296 191344
rect 161492 191304 207296 191332
rect 207290 191292 207296 191304
rect 207348 191292 207354 191344
rect 216858 191264 216864 191276
rect 161400 191236 216864 191264
rect 216858 191224 216864 191236
rect 216916 191224 216922 191276
rect 99190 191156 99196 191208
rect 99248 191196 99254 191208
rect 132862 191196 132868 191208
rect 99248 191168 132868 191196
rect 99248 191156 99254 191168
rect 132862 191156 132868 191168
rect 132920 191156 132926 191208
rect 140866 191196 140872 191208
rect 137986 191168 140872 191196
rect 106918 191088 106924 191140
rect 106976 191128 106982 191140
rect 137986 191128 138014 191168
rect 140866 191156 140872 191168
rect 140924 191156 140930 191208
rect 160186 191156 160192 191208
rect 160244 191196 160250 191208
rect 160462 191196 160468 191208
rect 160244 191168 160468 191196
rect 160244 191156 160250 191168
rect 160462 191156 160468 191168
rect 160520 191156 160526 191208
rect 161566 191156 161572 191208
rect 161624 191196 161630 191208
rect 161750 191196 161756 191208
rect 161624 191168 161756 191196
rect 161624 191156 161630 191168
rect 161750 191156 161756 191168
rect 161808 191156 161814 191208
rect 163130 191156 163136 191208
rect 163188 191196 163194 191208
rect 163498 191196 163504 191208
rect 163188 191168 163504 191196
rect 163188 191156 163194 191168
rect 163498 191156 163504 191168
rect 163556 191156 163562 191208
rect 164234 191156 164240 191208
rect 164292 191196 164298 191208
rect 165246 191196 165252 191208
rect 164292 191168 165252 191196
rect 164292 191156 164298 191168
rect 165246 191156 165252 191168
rect 165304 191156 165310 191208
rect 165706 191156 165712 191208
rect 165764 191196 165770 191208
rect 166350 191196 166356 191208
rect 165764 191168 166356 191196
rect 165764 191156 165770 191168
rect 166350 191156 166356 191168
rect 166408 191156 166414 191208
rect 166626 191156 166632 191208
rect 166684 191196 166690 191208
rect 218146 191196 218152 191208
rect 166684 191168 218152 191196
rect 166684 191156 166690 191168
rect 218146 191156 218152 191168
rect 218204 191156 218210 191208
rect 106976 191100 138014 191128
rect 106976 191088 106982 191100
rect 138290 191088 138296 191140
rect 138348 191128 138354 191140
rect 139210 191128 139216 191140
rect 138348 191100 139216 191128
rect 138348 191088 138354 191100
rect 139210 191088 139216 191100
rect 139268 191088 139274 191140
rect 139946 191088 139952 191140
rect 140004 191128 140010 191140
rect 140682 191128 140688 191140
rect 140004 191100 140688 191128
rect 140004 191088 140010 191100
rect 140682 191088 140688 191100
rect 140740 191088 140746 191140
rect 141326 191088 141332 191140
rect 141384 191128 141390 191140
rect 141970 191128 141976 191140
rect 141384 191100 141976 191128
rect 141384 191088 141390 191100
rect 141970 191088 141976 191100
rect 142028 191088 142034 191140
rect 145374 191088 145380 191140
rect 145432 191128 145438 191140
rect 146018 191128 146024 191140
rect 145432 191100 146024 191128
rect 145432 191088 145438 191100
rect 146018 191088 146024 191100
rect 146076 191088 146082 191140
rect 146662 191088 146668 191140
rect 146720 191128 146726 191140
rect 147398 191128 147404 191140
rect 146720 191100 147404 191128
rect 146720 191088 146726 191100
rect 147398 191088 147404 191100
rect 147456 191088 147462 191140
rect 151722 191088 151728 191140
rect 151780 191128 151786 191140
rect 218238 191128 218244 191140
rect 151780 191100 218244 191128
rect 151780 191088 151786 191100
rect 218238 191088 218244 191100
rect 218296 191088 218302 191140
rect 146386 191020 146392 191072
rect 146444 191060 146450 191072
rect 147030 191060 147036 191072
rect 146444 191032 147036 191060
rect 146444 191020 146450 191032
rect 147030 191020 147036 191032
rect 147088 191020 147094 191072
rect 157518 191020 157524 191072
rect 157576 191060 157582 191072
rect 158438 191060 158444 191072
rect 157576 191032 158444 191060
rect 157576 191020 157582 191032
rect 158438 191020 158444 191032
rect 158496 191020 158502 191072
rect 160186 191020 160192 191072
rect 160244 191060 160250 191072
rect 161198 191060 161204 191072
rect 160244 191032 161204 191060
rect 160244 191020 160250 191032
rect 161198 191020 161204 191032
rect 161256 191020 161262 191072
rect 161566 191020 161572 191072
rect 161624 191060 161630 191072
rect 162026 191060 162032 191072
rect 161624 191032 162032 191060
rect 161624 191020 161630 191032
rect 162026 191020 162032 191032
rect 162084 191020 162090 191072
rect 163406 191020 163412 191072
rect 163464 191060 163470 191072
rect 164050 191060 164056 191072
rect 163464 191032 164056 191060
rect 163464 191020 163470 191032
rect 164050 191020 164056 191032
rect 164108 191020 164114 191072
rect 164602 191020 164608 191072
rect 164660 191060 164666 191072
rect 165062 191060 165068 191072
rect 164660 191032 165068 191060
rect 164660 191020 164666 191032
rect 165062 191020 165068 191032
rect 165120 191020 165126 191072
rect 165890 191020 165896 191072
rect 165948 191060 165954 191072
rect 166718 191060 166724 191072
rect 165948 191032 166724 191060
rect 165948 191020 165954 191032
rect 166718 191020 166724 191032
rect 166776 191020 166782 191072
rect 200114 191060 200120 191072
rect 166828 191032 200120 191060
rect 164326 190952 164332 191004
rect 164384 190992 164390 191004
rect 164786 190992 164792 191004
rect 164384 190964 164792 190992
rect 164384 190952 164390 190964
rect 164786 190952 164792 190964
rect 164844 190952 164850 191004
rect 165614 190952 165620 191004
rect 165672 190992 165678 191004
rect 166828 190992 166856 191032
rect 200114 191020 200120 191032
rect 200172 191020 200178 191072
rect 165672 190964 166856 190992
rect 165672 190952 165678 190964
rect 166994 190952 167000 191004
rect 167052 190992 167058 191004
rect 167822 190992 167828 191004
rect 167052 190964 167828 190992
rect 167052 190952 167058 190964
rect 167822 190952 167828 190964
rect 167880 190952 167886 191004
rect 168558 190952 168564 191004
rect 168616 190992 168622 191004
rect 168926 190992 168932 191004
rect 168616 190964 168932 190992
rect 168616 190952 168622 190964
rect 168926 190952 168932 190964
rect 168984 190952 168990 191004
rect 169846 190952 169852 191004
rect 169904 190992 169910 191004
rect 170582 190992 170588 191004
rect 169904 190964 170588 190992
rect 169904 190952 169910 190964
rect 170582 190952 170588 190964
rect 170640 190952 170646 191004
rect 171134 190952 171140 191004
rect 171192 190992 171198 191004
rect 171962 190992 171968 191004
rect 171192 190964 171968 190992
rect 171192 190952 171198 190964
rect 171962 190952 171968 190964
rect 172020 190952 172026 191004
rect 172698 190952 172704 191004
rect 172756 190992 172762 191004
rect 173618 190992 173624 191004
rect 172756 190964 173624 190992
rect 172756 190952 172762 190964
rect 173618 190952 173624 190964
rect 173676 190952 173682 191004
rect 173986 190952 173992 191004
rect 174044 190992 174050 191004
rect 174446 190992 174452 191004
rect 174044 190964 174452 190992
rect 174044 190952 174050 190964
rect 174446 190952 174452 190964
rect 174504 190952 174510 191004
rect 175550 190952 175556 191004
rect 175608 190992 175614 191004
rect 176102 190992 176108 191004
rect 175608 190964 176108 190992
rect 175608 190952 175614 190964
rect 176102 190952 176108 190964
rect 176160 190952 176166 191004
rect 165798 190884 165804 190936
rect 165856 190924 165862 190936
rect 166166 190924 166172 190936
rect 165856 190896 166172 190924
rect 165856 190884 165862 190896
rect 166166 190884 166172 190896
rect 166224 190884 166230 190936
rect 167086 190884 167092 190936
rect 167144 190924 167150 190936
rect 168282 190924 168288 190936
rect 167144 190896 168288 190924
rect 167144 190884 167150 190896
rect 168282 190884 168288 190896
rect 168340 190884 168346 190936
rect 169754 190884 169760 190936
rect 169812 190924 169818 190936
rect 170858 190924 170864 190936
rect 169812 190896 170864 190924
rect 169812 190884 169818 190896
rect 170858 190884 170864 190896
rect 170916 190884 170922 190936
rect 171226 190884 171232 190936
rect 171284 190924 171290 190936
rect 172238 190924 172244 190936
rect 171284 190896 172244 190924
rect 171284 190884 171290 190896
rect 172238 190884 172244 190896
rect 172296 190884 172302 190936
rect 176930 190884 176936 190936
rect 176988 190924 176994 190936
rect 177666 190924 177672 190936
rect 176988 190896 177672 190924
rect 176988 190884 176994 190896
rect 177666 190884 177672 190896
rect 177724 190884 177730 190936
rect 167454 190816 167460 190868
rect 167512 190856 167518 190868
rect 175090 190856 175096 190868
rect 167512 190828 175096 190856
rect 167512 190816 167518 190828
rect 175090 190816 175096 190828
rect 175148 190816 175154 190868
rect 176838 190816 176844 190868
rect 176896 190856 176902 190868
rect 177390 190856 177396 190868
rect 176896 190828 177396 190856
rect 176896 190816 176902 190828
rect 177390 190816 177396 190828
rect 177448 190816 177454 190868
rect 167638 190748 167644 190800
rect 167696 190788 167702 190800
rect 174998 190788 175004 190800
rect 167696 190760 175004 190788
rect 167696 190748 167702 190760
rect 174998 190748 175004 190760
rect 175056 190748 175062 190800
rect 148134 190544 148140 190596
rect 148192 190584 148198 190596
rect 148778 190584 148784 190596
rect 148192 190556 148784 190584
rect 148192 190544 148198 190556
rect 148778 190544 148784 190556
rect 148836 190544 148842 190596
rect 156138 190544 156144 190596
rect 156196 190584 156202 190596
rect 157058 190584 157064 190596
rect 156196 190556 157064 190584
rect 156196 190544 156202 190556
rect 157058 190544 157064 190556
rect 157116 190544 157122 190596
rect 167914 190408 167920 190460
rect 167972 190448 167978 190460
rect 185762 190448 185768 190460
rect 167972 190420 185768 190448
rect 167972 190408 167978 190420
rect 185762 190408 185768 190420
rect 185820 190408 185826 190460
rect 162394 190340 162400 190392
rect 162452 190380 162458 190392
rect 183094 190380 183100 190392
rect 162452 190352 183100 190380
rect 162452 190340 162458 190352
rect 183094 190340 183100 190352
rect 183152 190340 183158 190392
rect 125318 190272 125324 190324
rect 125376 190312 125382 190324
rect 139854 190312 139860 190324
rect 125376 190284 139860 190312
rect 125376 190272 125382 190284
rect 139854 190272 139860 190284
rect 139912 190272 139918 190324
rect 160002 190272 160008 190324
rect 160060 190312 160066 190324
rect 185670 190312 185676 190324
rect 160060 190284 185676 190312
rect 160060 190272 160066 190284
rect 185670 190272 185676 190284
rect 185728 190272 185734 190324
rect 104710 190204 104716 190256
rect 104768 190244 104774 190256
rect 137462 190244 137468 190256
rect 104768 190216 137468 190244
rect 104768 190204 104774 190216
rect 137462 190204 137468 190216
rect 137520 190204 137526 190256
rect 153654 190204 153660 190256
rect 153712 190244 153718 190256
rect 181714 190244 181720 190256
rect 153712 190216 181720 190244
rect 153712 190204 153718 190216
rect 181714 190204 181720 190216
rect 181772 190204 181778 190256
rect 103422 190136 103428 190188
rect 103480 190176 103486 190188
rect 135438 190176 135444 190188
rect 103480 190148 135444 190176
rect 103480 190136 103486 190148
rect 135438 190136 135444 190148
rect 135496 190136 135502 190188
rect 152366 190136 152372 190188
rect 152424 190176 152430 190188
rect 183002 190176 183008 190188
rect 152424 190148 183008 190176
rect 152424 190136 152430 190148
rect 183002 190136 183008 190148
rect 183060 190136 183066 190188
rect 111518 190068 111524 190120
rect 111576 190108 111582 190120
rect 144454 190108 144460 190120
rect 111576 190080 144460 190108
rect 111576 190068 111582 190080
rect 144454 190068 144460 190080
rect 144512 190068 144518 190120
rect 177114 190068 177120 190120
rect 177172 190108 177178 190120
rect 210234 190108 210240 190120
rect 177172 190080 210240 190108
rect 177172 190068 177178 190080
rect 210234 190068 210240 190080
rect 210292 190068 210298 190120
rect 111058 190000 111064 190052
rect 111116 190040 111122 190052
rect 144086 190040 144092 190052
rect 111116 190012 144092 190040
rect 111116 190000 111122 190012
rect 144086 190000 144092 190012
rect 144144 190000 144150 190052
rect 176470 190000 176476 190052
rect 176528 190040 176534 190052
rect 210326 190040 210332 190052
rect 176528 190012 210332 190040
rect 176528 190000 176534 190012
rect 210326 190000 210332 190012
rect 210384 190000 210390 190052
rect 104066 189932 104072 189984
rect 104124 189972 104130 189984
rect 136910 189972 136916 189984
rect 104124 189944 136916 189972
rect 104124 189932 104130 189944
rect 136910 189932 136916 189944
rect 136968 189932 136974 189984
rect 176010 189932 176016 189984
rect 176068 189972 176074 189984
rect 210418 189972 210424 189984
rect 176068 189944 210424 189972
rect 176068 189932 176074 189944
rect 210418 189932 210424 189944
rect 210476 189932 210482 189984
rect 103054 189864 103060 189916
rect 103112 189904 103118 189916
rect 137186 189904 137192 189916
rect 103112 189876 137192 189904
rect 103112 189864 103118 189876
rect 137186 189864 137192 189876
rect 137244 189864 137250 189916
rect 177206 189864 177212 189916
rect 177264 189904 177270 189916
rect 211890 189904 211896 189916
rect 177264 189876 211896 189904
rect 177264 189864 177270 189876
rect 211890 189864 211896 189876
rect 211948 189864 211954 189916
rect 101582 189796 101588 189848
rect 101640 189836 101646 189848
rect 135346 189836 135352 189848
rect 101640 189808 135352 189836
rect 101640 189796 101646 189808
rect 135346 189796 135352 189808
rect 135404 189796 135410 189848
rect 158530 189796 158536 189848
rect 158588 189836 158594 189848
rect 212534 189836 212540 189848
rect 158588 189808 212540 189836
rect 158588 189796 158594 189808
rect 212534 189796 212540 189808
rect 212592 189796 212598 189848
rect 109678 189728 109684 189780
rect 109736 189768 109742 189780
rect 144270 189768 144276 189780
rect 109736 189740 144276 189768
rect 109736 189728 109742 189740
rect 144270 189728 144276 189740
rect 144328 189728 144334 189780
rect 152274 189728 152280 189780
rect 152332 189768 152338 189780
rect 218330 189768 218336 189780
rect 152332 189740 218336 189768
rect 152332 189728 152338 189740
rect 218330 189728 218336 189740
rect 218388 189728 218394 189780
rect 172514 189592 172520 189644
rect 172572 189632 172578 189644
rect 173342 189632 173348 189644
rect 172572 189604 173348 189632
rect 172572 189592 172578 189604
rect 173342 189592 173348 189604
rect 173400 189592 173406 189644
rect 3418 188980 3424 189032
rect 3476 189020 3482 189032
rect 120534 189020 120540 189032
rect 3476 188992 120540 189020
rect 3476 188980 3482 188992
rect 120534 188980 120540 188992
rect 120592 188980 120598 189032
rect 175366 188572 175372 188624
rect 175424 188612 175430 188624
rect 175642 188612 175648 188624
rect 175424 188584 175648 188612
rect 175424 188572 175430 188584
rect 175642 188572 175648 188584
rect 175700 188572 175706 188624
rect 175366 188436 175372 188488
rect 175424 188476 175430 188488
rect 176378 188476 176384 188488
rect 175424 188448 176384 188476
rect 175424 188436 175430 188448
rect 176378 188436 176384 188448
rect 176436 188436 176442 188488
rect 169938 188368 169944 188420
rect 169996 188408 170002 188420
rect 170306 188408 170312 188420
rect 169996 188380 170312 188408
rect 169996 188368 170002 188380
rect 170306 188368 170312 188380
rect 170364 188368 170370 188420
rect 121822 187484 121828 187536
rect 121880 187524 121886 187536
rect 149238 187524 149244 187536
rect 121880 187496 149244 187524
rect 121880 187484 121886 187496
rect 149238 187484 149244 187496
rect 149296 187484 149302 187536
rect 109770 187416 109776 187468
rect 109828 187456 109834 187468
rect 140498 187456 140504 187468
rect 109828 187428 140504 187456
rect 109828 187416 109834 187428
rect 140498 187416 140504 187428
rect 140556 187416 140562 187468
rect 109586 187348 109592 187400
rect 109644 187388 109650 187400
rect 141878 187388 141884 187400
rect 109644 187360 141884 187388
rect 109644 187348 109650 187360
rect 141878 187348 141884 187360
rect 141936 187348 141942 187400
rect 169018 187348 169024 187400
rect 169076 187388 169082 187400
rect 169076 187360 176654 187388
rect 169076 187348 169082 187360
rect 103146 187280 103152 187332
rect 103204 187320 103210 187332
rect 135898 187320 135904 187332
rect 103204 187292 135904 187320
rect 103204 187280 103210 187292
rect 135898 187280 135904 187292
rect 135956 187280 135962 187332
rect 168466 187280 168472 187332
rect 168524 187320 168530 187332
rect 169662 187320 169668 187332
rect 168524 187292 169668 187320
rect 168524 187280 168530 187292
rect 169662 187280 169668 187292
rect 169720 187280 169726 187332
rect 176626 187320 176654 187360
rect 203334 187320 203340 187332
rect 176626 187292 203340 187320
rect 203334 187280 203340 187292
rect 203392 187280 203398 187332
rect 100478 187212 100484 187264
rect 100536 187252 100542 187264
rect 132770 187252 132776 187264
rect 100536 187224 132776 187252
rect 100536 187212 100542 187224
rect 132770 187212 132776 187224
rect 132828 187212 132834 187264
rect 153562 187212 153568 187264
rect 153620 187252 153626 187264
rect 214006 187252 214012 187264
rect 153620 187224 214012 187252
rect 153620 187212 153626 187224
rect 214006 187212 214012 187224
rect 214064 187212 214070 187264
rect 101490 187144 101496 187196
rect 101548 187184 101554 187196
rect 134518 187184 134524 187196
rect 101548 187156 134524 187184
rect 101548 187144 101554 187156
rect 134518 187144 134524 187156
rect 134576 187144 134582 187196
rect 149790 187144 149796 187196
rect 149848 187184 149854 187196
rect 211430 187184 211436 187196
rect 149848 187156 211436 187184
rect 149848 187144 149854 187156
rect 211430 187144 211436 187156
rect 211488 187144 211494 187196
rect 99006 187076 99012 187128
rect 99064 187116 99070 187128
rect 133138 187116 133144 187128
rect 99064 187088 133144 187116
rect 99064 187076 99070 187088
rect 133138 187076 133144 187088
rect 133196 187076 133202 187128
rect 149330 187076 149336 187128
rect 149388 187116 149394 187128
rect 211706 187116 211712 187128
rect 149388 187088 211712 187116
rect 149388 187076 149394 187088
rect 211706 187076 211712 187088
rect 211764 187076 211770 187128
rect 100294 187008 100300 187060
rect 100352 187048 100358 187060
rect 135070 187048 135076 187060
rect 100352 187020 135076 187048
rect 100352 187008 100358 187020
rect 135070 187008 135076 187020
rect 135128 187008 135134 187060
rect 151078 187008 151084 187060
rect 151136 187048 151142 187060
rect 215846 187048 215852 187060
rect 151136 187020 215852 187048
rect 151136 187008 151142 187020
rect 215846 187008 215852 187020
rect 215904 187008 215910 187060
rect 100386 186940 100392 186992
rect 100444 186980 100450 186992
rect 134242 186980 134248 186992
rect 100444 186952 134248 186980
rect 100444 186940 100450 186952
rect 134242 186940 134248 186952
rect 134300 186940 134306 186992
rect 150986 186940 150992 186992
rect 151044 186980 151050 186992
rect 218422 186980 218428 186992
rect 151044 186952 218428 186980
rect 151044 186940 151050 186952
rect 218422 186940 218428 186952
rect 218480 186940 218486 186992
rect 188338 178032 188344 178084
rect 188396 178072 188402 178084
rect 580166 178072 580172 178084
rect 188396 178044 580172 178072
rect 188396 178032 188402 178044
rect 580166 178032 580172 178044
rect 580224 178032 580230 178084
rect 189902 165588 189908 165640
rect 189960 165628 189966 165640
rect 580166 165628 580172 165640
rect 189960 165600 580172 165628
rect 189960 165588 189966 165600
rect 580166 165588 580172 165600
rect 580224 165588 580230 165640
rect 98914 164840 98920 164892
rect 98972 164880 98978 164892
rect 130654 164880 130660 164892
rect 98972 164852 130660 164880
rect 98972 164840 98978 164852
rect 130654 164840 130660 164852
rect 130712 164840 130718 164892
rect 175734 159740 175740 159792
rect 175792 159780 175798 159792
rect 199194 159780 199200 159792
rect 175792 159752 199200 159780
rect 175792 159740 175798 159752
rect 199194 159740 199200 159752
rect 199252 159740 199258 159792
rect 172790 159672 172796 159724
rect 172848 159712 172854 159724
rect 196618 159712 196624 159724
rect 172848 159684 196624 159712
rect 172848 159672 172854 159684
rect 196618 159672 196624 159684
rect 196676 159672 196682 159724
rect 161842 159604 161848 159656
rect 161900 159644 161906 159656
rect 195146 159644 195152 159656
rect 161900 159616 195152 159644
rect 161900 159604 161906 159616
rect 195146 159604 195152 159616
rect 195204 159604 195210 159656
rect 172606 159536 172612 159588
rect 172664 159576 172670 159588
rect 211982 159576 211988 159588
rect 172664 159548 211988 159576
rect 172664 159536 172670 159548
rect 211982 159536 211988 159548
rect 212040 159536 212046 159588
rect 149974 159468 149980 159520
rect 150032 159508 150038 159520
rect 209130 159508 209136 159520
rect 150032 159480 209136 159508
rect 150032 159468 150038 159480
rect 209130 159468 209136 159480
rect 209188 159468 209194 159520
rect 152090 159400 152096 159452
rect 152148 159440 152154 159452
rect 213914 159440 213920 159452
rect 152148 159412 213920 159440
rect 152148 159400 152154 159412
rect 213914 159400 213920 159412
rect 213972 159400 213978 159452
rect 152182 159332 152188 159384
rect 152240 159372 152246 159384
rect 214190 159372 214196 159384
rect 152240 159344 214196 159372
rect 152240 159332 152246 159344
rect 214190 159332 214196 159344
rect 214248 159332 214254 159384
rect 177850 157292 177856 157344
rect 177908 157332 177914 157344
rect 203426 157332 203432 157344
rect 177908 157304 203432 157332
rect 177908 157292 177914 157304
rect 203426 157292 203432 157304
rect 203484 157292 203490 157344
rect 163590 157224 163596 157276
rect 163648 157264 163654 157276
rect 192386 157264 192392 157276
rect 163648 157236 192392 157264
rect 163648 157224 163654 157236
rect 192386 157224 192392 157236
rect 192444 157224 192450 157276
rect 161934 157156 161940 157208
rect 161992 157196 161998 157208
rect 193766 157196 193772 157208
rect 161992 157168 193772 157196
rect 161992 157156 161998 157168
rect 193766 157156 193772 157168
rect 193824 157156 193830 157208
rect 176930 157088 176936 157140
rect 176988 157128 176994 157140
rect 210602 157128 210608 157140
rect 176988 157100 210608 157128
rect 176988 157088 176994 157100
rect 210602 157088 210608 157100
rect 210660 157088 210666 157140
rect 168558 157020 168564 157072
rect 168616 157060 168622 157072
rect 203794 157060 203800 157072
rect 168616 157032 203800 157060
rect 168616 157020 168622 157032
rect 203794 157020 203800 157032
rect 203852 157020 203858 157072
rect 167270 156952 167276 157004
rect 167328 156992 167334 157004
rect 201954 156992 201960 157004
rect 167328 156964 201960 156992
rect 167328 156952 167334 156964
rect 201954 156952 201960 156964
rect 202012 156952 202018 157004
rect 168650 156884 168656 156936
rect 168708 156924 168714 156936
rect 203426 156924 203432 156936
rect 168708 156896 203432 156924
rect 168708 156884 168714 156896
rect 203426 156884 203432 156896
rect 203484 156884 203490 156936
rect 167178 156816 167184 156868
rect 167236 156856 167242 156868
rect 202138 156856 202144 156868
rect 167236 156828 202144 156856
rect 167236 156816 167242 156828
rect 202138 156816 202144 156828
rect 202196 156816 202202 156868
rect 164878 156748 164884 156800
rect 164936 156788 164942 156800
rect 201862 156788 201868 156800
rect 164936 156760 201868 156788
rect 164936 156748 164942 156760
rect 201862 156748 201868 156760
rect 201920 156748 201926 156800
rect 160738 156680 160744 156732
rect 160796 156720 160802 156732
rect 200574 156720 200580 156732
rect 160796 156692 200580 156720
rect 160796 156680 160802 156692
rect 200574 156680 200580 156692
rect 200632 156680 200638 156732
rect 155862 156612 155868 156664
rect 155920 156652 155926 156664
rect 200942 156652 200948 156664
rect 155920 156624 200948 156652
rect 155920 156612 155926 156624
rect 200942 156612 200948 156624
rect 201000 156612 201006 156664
rect 163498 156544 163504 156596
rect 163556 156584 163562 156596
rect 188246 156584 188252 156596
rect 163556 156556 188252 156584
rect 163556 156544 163562 156556
rect 188246 156544 188252 156556
rect 188304 156544 188310 156596
rect 166258 156476 166264 156528
rect 166316 156516 166322 156528
rect 189718 156516 189724 156528
rect 166316 156488 189724 156516
rect 166316 156476 166322 156488
rect 189718 156476 189724 156488
rect 189776 156476 189782 156528
rect 165890 154504 165896 154556
rect 165948 154544 165954 154556
rect 185854 154544 185860 154556
rect 165948 154516 185860 154544
rect 165948 154504 165954 154516
rect 185854 154504 185860 154516
rect 185912 154504 185918 154556
rect 160646 154436 160652 154488
rect 160704 154476 160710 154488
rect 185946 154476 185952 154488
rect 160704 154448 185952 154476
rect 160704 154436 160710 154448
rect 185946 154436 185952 154448
rect 186004 154436 186010 154488
rect 158898 154368 158904 154420
rect 158956 154408 158962 154420
rect 184290 154408 184296 154420
rect 158956 154380 184296 154408
rect 158956 154368 158962 154380
rect 184290 154368 184296 154380
rect 184348 154368 184354 154420
rect 158990 154300 158996 154352
rect 159048 154340 159054 154352
rect 183738 154340 183744 154352
rect 159048 154312 183744 154340
rect 159048 154300 159054 154312
rect 183738 154300 183744 154312
rect 183796 154300 183802 154352
rect 157518 154232 157524 154284
rect 157576 154272 157582 154284
rect 186130 154272 186136 154284
rect 157576 154244 186136 154272
rect 157576 154232 157582 154244
rect 186130 154232 186136 154244
rect 186188 154232 186194 154284
rect 157610 154164 157616 154216
rect 157668 154204 157674 154216
rect 186038 154204 186044 154216
rect 157668 154176 186044 154204
rect 157668 154164 157674 154176
rect 186038 154164 186044 154176
rect 186096 154164 186102 154216
rect 157242 154096 157248 154148
rect 157300 154136 157306 154148
rect 186222 154136 186228 154148
rect 157300 154108 186228 154136
rect 157300 154096 157306 154108
rect 186222 154096 186228 154108
rect 186280 154096 186286 154148
rect 164786 154028 164792 154080
rect 164844 154068 164850 154080
rect 199194 154068 199200 154080
rect 164844 154040 199200 154068
rect 164844 154028 164850 154040
rect 199194 154028 199200 154040
rect 199252 154028 199258 154080
rect 165982 153960 165988 154012
rect 166040 154000 166046 154012
rect 200574 154000 200580 154012
rect 166040 153972 200580 154000
rect 166040 153960 166046 153972
rect 200574 153960 200580 153972
rect 200632 153960 200638 154012
rect 166902 153892 166908 153944
rect 166960 153932 166966 153944
rect 200666 153932 200672 153944
rect 166960 153904 200672 153932
rect 166960 153892 166966 153904
rect 200666 153892 200672 153904
rect 200724 153892 200730 153944
rect 121914 153824 121920 153876
rect 121972 153864 121978 153876
rect 143626 153864 143632 153876
rect 121972 153836 143632 153864
rect 121972 153824 121978 153836
rect 143626 153824 143632 153836
rect 143684 153824 143690 153876
rect 146202 153824 146208 153876
rect 146260 153864 146266 153876
rect 202046 153864 202052 153876
rect 146260 153836 202052 153864
rect 146260 153824 146266 153836
rect 202046 153824 202052 153836
rect 202104 153824 202110 153876
rect 166166 153756 166172 153808
rect 166224 153796 166230 153808
rect 183278 153796 183284 153808
rect 166224 153768 183284 153796
rect 166224 153756 166230 153768
rect 183278 153756 183284 153768
rect 183336 153756 183342 153808
rect 164694 152736 164700 152788
rect 164752 152776 164758 152788
rect 206186 152776 206192 152788
rect 164752 152748 206192 152776
rect 164752 152736 164758 152748
rect 206186 152736 206192 152748
rect 206244 152736 206250 152788
rect 154850 152668 154856 152720
rect 154908 152708 154914 152720
rect 203058 152708 203064 152720
rect 154908 152680 203064 152708
rect 154908 152668 154914 152680
rect 203058 152668 203064 152680
rect 203116 152668 203122 152720
rect 163406 152600 163412 152652
rect 163464 152640 163470 152652
rect 213086 152640 213092 152652
rect 163464 152612 213092 152640
rect 163464 152600 163470 152612
rect 213086 152600 213092 152612
rect 213144 152600 213150 152652
rect 121638 152532 121644 152584
rect 121696 152572 121702 152584
rect 150894 152572 150900 152584
rect 121696 152544 150900 152572
rect 121696 152532 121702 152544
rect 150894 152532 150900 152544
rect 150952 152532 150958 152584
rect 153562 152532 153568 152584
rect 153620 152572 153626 152584
rect 204530 152572 204536 152584
rect 153620 152544 204536 152572
rect 153620 152532 153626 152544
rect 204530 152532 204536 152544
rect 204588 152532 204594 152584
rect 121546 152464 121552 152516
rect 121604 152504 121610 152516
rect 150802 152504 150808 152516
rect 121604 152476 150808 152504
rect 121604 152464 121610 152476
rect 150802 152464 150808 152476
rect 150860 152464 150866 152516
rect 155678 152464 155684 152516
rect 155736 152504 155742 152516
rect 214282 152504 214288 152516
rect 155736 152476 214288 152504
rect 155736 152464 155742 152476
rect 214282 152464 214288 152476
rect 214340 152464 214346 152516
rect 185486 152396 185492 152448
rect 185544 152436 185550 152448
rect 185670 152436 185676 152448
rect 185544 152408 185676 152436
rect 185544 152396 185550 152408
rect 185670 152396 185676 152408
rect 185728 152396 185734 152448
rect 188246 151784 188252 151836
rect 188304 151824 188310 151836
rect 579982 151824 579988 151836
rect 188304 151796 579988 151824
rect 188304 151784 188310 151796
rect 579982 151784 579988 151796
rect 580040 151784 580046 151836
rect 99834 151716 99840 151768
rect 99892 151756 99898 151768
rect 132678 151756 132684 151768
rect 99892 151728 132684 151756
rect 99892 151716 99898 151728
rect 132678 151716 132684 151728
rect 132736 151716 132742 151768
rect 100110 151648 100116 151700
rect 100168 151688 100174 151700
rect 134334 151688 134340 151700
rect 100168 151660 134340 151688
rect 100168 151648 100174 151660
rect 134334 151648 134340 151660
rect 134392 151648 134398 151700
rect 100202 151580 100208 151632
rect 100260 151620 100266 151632
rect 134426 151620 134432 151632
rect 100260 151592 134432 151620
rect 100260 151580 100266 151592
rect 134426 151580 134432 151592
rect 134484 151580 134490 151632
rect 164602 151580 164608 151632
rect 164660 151620 164666 151632
rect 181806 151620 181812 151632
rect 164660 151592 181812 151620
rect 164660 151580 164666 151592
rect 181806 151580 181812 151592
rect 181864 151580 181870 151632
rect 98822 151512 98828 151564
rect 98880 151552 98886 151564
rect 133046 151552 133052 151564
rect 98880 151524 133052 151552
rect 98880 151512 98886 151524
rect 133046 151512 133052 151524
rect 133104 151512 133110 151564
rect 161750 151512 161756 151564
rect 161808 151552 161814 151564
rect 185394 151552 185400 151564
rect 161808 151524 185400 151552
rect 161808 151512 161814 151524
rect 185394 151512 185400 151524
rect 185452 151512 185458 151564
rect 100018 151444 100024 151496
rect 100076 151484 100082 151496
rect 134610 151484 134616 151496
rect 100076 151456 134616 151484
rect 100076 151444 100082 151456
rect 134610 151444 134616 151456
rect 134668 151444 134674 151496
rect 157426 151444 157432 151496
rect 157484 151484 157490 151496
rect 184382 151484 184388 151496
rect 157484 151456 184388 151484
rect 157484 151444 157490 151456
rect 184382 151444 184388 151456
rect 184440 151444 184446 151496
rect 101398 151376 101404 151428
rect 101456 151416 101462 151428
rect 135622 151416 135628 151428
rect 101456 151388 135628 151416
rect 101456 151376 101462 151388
rect 135622 151376 135628 151388
rect 135680 151376 135686 151428
rect 157334 151376 157340 151428
rect 157392 151416 157398 151428
rect 184842 151416 184848 151428
rect 157392 151388 184848 151416
rect 157392 151376 157398 151388
rect 184842 151376 184848 151388
rect 184900 151376 184906 151428
rect 101306 151308 101312 151360
rect 101364 151348 101370 151360
rect 135530 151348 135536 151360
rect 101364 151320 135536 151348
rect 101364 151308 101370 151320
rect 135530 151308 135536 151320
rect 135588 151308 135594 151360
rect 175550 151308 175556 151360
rect 175608 151348 175614 151360
rect 205082 151348 205088 151360
rect 175608 151320 205088 151348
rect 175608 151308 175614 151320
rect 205082 151308 205088 151320
rect 205140 151308 205146 151360
rect 99926 151240 99932 151292
rect 99984 151280 99990 151292
rect 134150 151280 134156 151292
rect 99984 151252 134156 151280
rect 99984 151240 99990 151252
rect 134150 151240 134156 151252
rect 134208 151240 134214 151292
rect 175642 151240 175648 151292
rect 175700 151280 175706 151292
rect 206370 151280 206376 151292
rect 175700 151252 206376 151280
rect 175700 151240 175706 151252
rect 206370 151240 206376 151252
rect 206428 151240 206434 151292
rect 122006 151172 122012 151224
rect 122064 151212 122070 151224
rect 158714 151212 158720 151224
rect 122064 151184 158720 151212
rect 122064 151172 122070 151184
rect 158714 151172 158720 151184
rect 158772 151172 158778 151224
rect 174170 151172 174176 151224
rect 174228 151212 174234 151224
rect 204990 151212 204996 151224
rect 174228 151184 204996 151212
rect 174228 151172 174234 151184
rect 204990 151172 204996 151184
rect 205048 151172 205054 151224
rect 122374 151104 122380 151156
rect 122432 151144 122438 151156
rect 160094 151144 160100 151156
rect 122432 151116 160100 151144
rect 122432 151104 122438 151116
rect 160094 151104 160100 151116
rect 160152 151104 160158 151156
rect 176746 151104 176752 151156
rect 176804 151144 176810 151156
rect 207750 151144 207756 151156
rect 176804 151116 207756 151144
rect 176804 151104 176810 151116
rect 207750 151104 207756 151116
rect 207808 151104 207814 151156
rect 97442 151036 97448 151088
rect 97500 151076 97506 151088
rect 141142 151076 141148 151088
rect 97500 151048 141148 151076
rect 97500 151036 97506 151048
rect 141142 151036 141148 151048
rect 141200 151036 141206 151088
rect 174078 151036 174084 151088
rect 174136 151076 174142 151088
rect 206278 151076 206284 151088
rect 174136 151048 206284 151076
rect 174136 151036 174142 151048
rect 206278 151036 206284 151048
rect 206336 151036 206342 151088
rect 102594 150968 102600 151020
rect 102652 151008 102658 151020
rect 135990 151008 135996 151020
rect 102652 150980 135996 151008
rect 102652 150968 102658 150980
rect 135990 150968 135996 150980
rect 136048 150968 136054 151020
rect 123662 150900 123668 150952
rect 123720 150940 123726 150952
rect 138382 150940 138388 150952
rect 123720 150912 138388 150940
rect 123720 150900 123726 150912
rect 138382 150900 138388 150912
rect 138440 150900 138446 150952
rect 172238 150356 172244 150408
rect 172296 150396 172302 150408
rect 192754 150396 192760 150408
rect 172296 150368 192760 150396
rect 172296 150356 172302 150368
rect 192754 150356 192760 150368
rect 192812 150356 192818 150408
rect 173250 150288 173256 150340
rect 173308 150328 173314 150340
rect 196710 150328 196716 150340
rect 173308 150300 196716 150328
rect 173308 150288 173314 150300
rect 196710 150288 196716 150300
rect 196768 150288 196774 150340
rect 158898 150220 158904 150272
rect 158956 150260 158962 150272
rect 188154 150260 188160 150272
rect 158956 150232 188160 150260
rect 158956 150220 158962 150232
rect 188154 150220 188160 150232
rect 188212 150220 188218 150272
rect 163130 150152 163136 150204
rect 163188 150192 163194 150204
rect 195146 150192 195152 150204
rect 163188 150164 195152 150192
rect 163188 150152 163194 150164
rect 195146 150152 195152 150164
rect 195204 150152 195210 150204
rect 166994 150084 167000 150136
rect 167052 150124 167058 150136
rect 200850 150124 200856 150136
rect 167052 150096 200856 150124
rect 167052 150084 167058 150096
rect 200850 150084 200856 150096
rect 200908 150084 200914 150136
rect 163222 150016 163228 150068
rect 163280 150056 163286 150068
rect 198274 150056 198280 150068
rect 163280 150028 198280 150056
rect 163280 150016 163286 150028
rect 198274 150016 198280 150028
rect 198332 150016 198338 150068
rect 164418 149948 164424 150000
rect 164476 149988 164482 150000
rect 199746 149988 199752 150000
rect 164476 149960 199752 149988
rect 164476 149948 164482 149960
rect 199746 149948 199752 149960
rect 199804 149948 199810 150000
rect 163314 149880 163320 149932
rect 163372 149920 163378 149932
rect 198458 149920 198464 149932
rect 163372 149892 198464 149920
rect 163372 149880 163378 149892
rect 198458 149880 198464 149892
rect 198516 149880 198522 149932
rect 165798 149812 165804 149864
rect 165856 149852 165862 149864
rect 200758 149852 200764 149864
rect 165856 149824 200764 149852
rect 165856 149812 165862 149824
rect 200758 149812 200764 149824
rect 200816 149812 200822 149864
rect 164510 149744 164516 149796
rect 164568 149784 164574 149796
rect 199470 149784 199476 149796
rect 164568 149756 199476 149784
rect 164568 149744 164574 149756
rect 199470 149744 199476 149756
rect 199528 149744 199534 149796
rect 158622 149676 158628 149728
rect 158680 149716 158686 149728
rect 195514 149716 195520 149728
rect 158680 149688 195520 149716
rect 158680 149676 158686 149688
rect 195514 149676 195520 149688
rect 195572 149676 195578 149728
rect 165522 149608 165528 149660
rect 165580 149648 165586 149660
rect 182082 149648 182088 149660
rect 165580 149620 182088 149648
rect 165580 149608 165586 149620
rect 182082 149608 182088 149620
rect 182140 149608 182146 149660
rect 180886 149540 180892 149592
rect 180944 149580 180950 149592
rect 198090 149580 198096 149592
rect 180944 149552 198096 149580
rect 180944 149540 180950 149552
rect 198090 149540 198096 149552
rect 198148 149540 198154 149592
rect 3142 149132 3148 149184
rect 3200 149172 3206 149184
rect 180886 149172 180892 149184
rect 3200 149144 180892 149172
rect 3200 149132 3206 149144
rect 180886 149132 180892 149144
rect 180944 149132 180950 149184
rect 119338 149064 119344 149116
rect 119396 149104 119402 149116
rect 580534 149104 580540 149116
rect 119396 149076 580540 149104
rect 119396 149064 119402 149076
rect 580534 149064 580540 149076
rect 580592 149064 580598 149116
rect 112530 148996 112536 149048
rect 112588 149036 112594 149048
rect 142522 149036 142528 149048
rect 112588 149008 142528 149036
rect 112588 148996 112594 149008
rect 142522 148996 142528 149008
rect 142580 148996 142586 149048
rect 112070 148928 112076 148980
rect 112128 148968 112134 148980
rect 142430 148968 142436 148980
rect 112128 148940 142436 148968
rect 112128 148928 112134 148940
rect 142430 148928 142436 148940
rect 142488 148928 142494 148980
rect 112162 148860 112168 148912
rect 112220 148900 112226 148912
rect 143902 148900 143908 148912
rect 112220 148872 143908 148900
rect 112220 148860 112226 148872
rect 143902 148860 143908 148872
rect 143960 148860 143966 148912
rect 162670 148860 162676 148912
rect 162728 148900 162734 148912
rect 188614 148900 188620 148912
rect 162728 148872 188620 148900
rect 162728 148860 162734 148872
rect 188614 148860 188620 148872
rect 188672 148860 188678 148912
rect 110782 148792 110788 148844
rect 110840 148832 110846 148844
rect 142614 148832 142620 148844
rect 110840 148804 142620 148832
rect 110840 148792 110846 148804
rect 142614 148792 142620 148804
rect 142672 148792 142678 148844
rect 156138 148792 156144 148844
rect 156196 148832 156202 148844
rect 184566 148832 184572 148844
rect 156196 148804 184572 148832
rect 156196 148792 156202 148804
rect 184566 148792 184572 148804
rect 184624 148792 184630 148844
rect 118970 148724 118976 148776
rect 119028 148764 119034 148776
rect 150618 148764 150624 148776
rect 119028 148736 150624 148764
rect 119028 148724 119034 148736
rect 150618 148724 150624 148736
rect 150676 148724 150682 148776
rect 170030 148724 170036 148776
rect 170088 148764 170094 148776
rect 199286 148764 199292 148776
rect 170088 148736 199292 148764
rect 170088 148724 170094 148736
rect 199286 148724 199292 148736
rect 199344 148724 199350 148776
rect 117682 148656 117688 148708
rect 117740 148696 117746 148708
rect 150710 148696 150716 148708
rect 117740 148668 150716 148696
rect 117740 148656 117746 148668
rect 150710 148656 150716 148668
rect 150768 148656 150774 148708
rect 173802 148656 173808 148708
rect 173860 148696 173866 148708
rect 204530 148696 204536 148708
rect 173860 148668 204536 148696
rect 173860 148656 173866 148668
rect 204530 148656 204536 148668
rect 204588 148656 204594 148708
rect 114830 148588 114836 148640
rect 114888 148628 114894 148640
rect 149514 148628 149520 148640
rect 114888 148600 149520 148628
rect 114888 148588 114894 148600
rect 149514 148588 149520 148600
rect 149572 148588 149578 148640
rect 171226 148588 171232 148640
rect 171284 148628 171290 148640
rect 202230 148628 202236 148640
rect 171284 148600 202236 148628
rect 171284 148588 171290 148600
rect 202230 148588 202236 148600
rect 202288 148588 202294 148640
rect 98730 148520 98736 148572
rect 98788 148560 98794 148572
rect 132954 148560 132960 148572
rect 98788 148532 132960 148560
rect 98788 148520 98794 148532
rect 132954 148520 132960 148532
rect 133012 148520 133018 148572
rect 171410 148520 171416 148572
rect 171468 148560 171474 148572
rect 203518 148560 203524 148572
rect 171468 148532 203524 148560
rect 171468 148520 171474 148532
rect 203518 148520 203524 148532
rect 203576 148520 203582 148572
rect 101214 148452 101220 148504
rect 101272 148492 101278 148504
rect 135714 148492 135720 148504
rect 101272 148464 135720 148492
rect 101272 148452 101278 148464
rect 135714 148452 135720 148464
rect 135772 148452 135778 148504
rect 171318 148452 171324 148504
rect 171376 148492 171382 148504
rect 203702 148492 203708 148504
rect 171376 148464 203708 148492
rect 171376 148452 171382 148464
rect 203702 148452 203708 148464
rect 203760 148452 203766 148504
rect 97534 148384 97540 148436
rect 97592 148424 97598 148436
rect 141050 148424 141056 148436
rect 97592 148396 141056 148424
rect 97592 148384 97598 148396
rect 141050 148384 141056 148396
rect 141108 148384 141114 148436
rect 173986 148384 173992 148436
rect 174044 148424 174050 148436
rect 206462 148424 206468 148436
rect 174044 148396 206468 148424
rect 174044 148384 174050 148396
rect 206462 148384 206468 148396
rect 206520 148384 206526 148436
rect 113634 148316 113640 148368
rect 113692 148356 113698 148368
rect 128630 148356 128636 148368
rect 113692 148328 128636 148356
rect 113692 148316 113698 148328
rect 128630 148316 128636 148328
rect 128688 148356 128694 148368
rect 188246 148356 188252 148368
rect 128688 148328 188252 148356
rect 128688 148316 128694 148328
rect 188246 148316 188252 148328
rect 188304 148316 188310 148368
rect 115566 148248 115572 148300
rect 115624 148288 115630 148300
rect 115842 148288 115848 148300
rect 115624 148260 115848 148288
rect 115624 148248 115630 148260
rect 115842 148248 115848 148260
rect 115900 148248 115906 148300
rect 142982 148288 142988 148300
rect 116136 148260 142988 148288
rect 113450 148112 113456 148164
rect 113508 148152 113514 148164
rect 116136 148152 116164 148260
rect 142982 148248 142988 148260
rect 143040 148248 143046 148300
rect 113508 148124 116164 148152
rect 113508 148112 113514 148124
rect 105446 148044 105452 148096
rect 105504 148084 105510 148096
rect 131850 148084 131856 148096
rect 105504 148056 131856 148084
rect 105504 148044 105510 148056
rect 131850 148044 131856 148056
rect 131908 148044 131914 148096
rect 124030 147636 124036 147688
rect 124088 147676 124094 147688
rect 580442 147676 580448 147688
rect 124088 147648 580448 147676
rect 124088 147636 124094 147648
rect 580442 147636 580448 147648
rect 580500 147636 580506 147688
rect 126790 147568 126796 147620
rect 126848 147608 126854 147620
rect 140130 147608 140136 147620
rect 126848 147580 140136 147608
rect 126848 147568 126854 147580
rect 140130 147568 140136 147580
rect 140188 147568 140194 147620
rect 179046 147568 179052 147620
rect 179104 147608 179110 147620
rect 196986 147608 196992 147620
rect 179104 147580 196992 147608
rect 179104 147568 179110 147580
rect 196986 147568 196992 147580
rect 197044 147568 197050 147620
rect 123478 147500 123484 147552
rect 123536 147540 123542 147552
rect 140314 147540 140320 147552
rect 123536 147512 140320 147540
rect 123536 147500 123542 147512
rect 140314 147500 140320 147512
rect 140372 147500 140378 147552
rect 174722 147500 174728 147552
rect 174780 147540 174786 147552
rect 194134 147540 194140 147552
rect 174780 147512 194140 147540
rect 174780 147500 174786 147512
rect 194134 147500 194140 147512
rect 194192 147500 194198 147552
rect 112438 147432 112444 147484
rect 112496 147472 112502 147484
rect 131758 147472 131764 147484
rect 112496 147444 131764 147472
rect 112496 147432 112502 147444
rect 131758 147432 131764 147444
rect 131816 147432 131822 147484
rect 164142 147432 164148 147484
rect 164200 147472 164206 147484
rect 181898 147472 181904 147484
rect 164200 147444 181904 147472
rect 164200 147432 164206 147444
rect 181898 147432 181904 147444
rect 181956 147432 181962 147484
rect 110966 147364 110972 147416
rect 111024 147404 111030 147416
rect 131942 147404 131948 147416
rect 111024 147376 131948 147404
rect 111024 147364 111030 147376
rect 131942 147364 131948 147376
rect 132000 147364 132006 147416
rect 160370 147364 160376 147416
rect 160428 147404 160434 147416
rect 188154 147404 188160 147416
rect 160428 147376 188160 147404
rect 160428 147364 160434 147376
rect 188154 147364 188160 147376
rect 188212 147364 188218 147416
rect 118878 147296 118884 147348
rect 118936 147336 118942 147348
rect 141326 147336 141332 147348
rect 118936 147308 141332 147336
rect 118936 147296 118942 147308
rect 141326 147296 141332 147308
rect 141384 147296 141390 147348
rect 164050 147296 164056 147348
rect 164108 147336 164114 147348
rect 192846 147336 192852 147348
rect 164108 147308 192852 147336
rect 164108 147296 164114 147308
rect 192846 147296 192852 147308
rect 192904 147296 192910 147348
rect 121914 147228 121920 147280
rect 121972 147268 121978 147280
rect 145558 147268 145564 147280
rect 121972 147240 145564 147268
rect 121972 147228 121978 147240
rect 145558 147228 145564 147240
rect 145616 147228 145622 147280
rect 160002 147228 160008 147280
rect 160060 147268 160066 147280
rect 191374 147268 191380 147280
rect 160060 147240 191380 147268
rect 160060 147228 160066 147240
rect 191374 147228 191380 147240
rect 191432 147228 191438 147280
rect 108114 147160 108120 147212
rect 108172 147200 108178 147212
rect 138566 147200 138572 147212
rect 108172 147172 138572 147200
rect 108172 147160 108178 147172
rect 138566 147160 138572 147172
rect 138624 147160 138630 147212
rect 160554 147160 160560 147212
rect 160612 147200 160618 147212
rect 193858 147200 193864 147212
rect 160612 147172 193864 147200
rect 160612 147160 160618 147172
rect 193858 147160 193864 147172
rect 193916 147160 193922 147212
rect 109494 147092 109500 147144
rect 109552 147132 109558 147144
rect 141694 147132 141700 147144
rect 109552 147104 141700 147132
rect 109552 147092 109558 147104
rect 141694 147092 141700 147104
rect 141752 147092 141758 147144
rect 158806 147092 158812 147144
rect 158864 147132 158870 147144
rect 192386 147132 192392 147144
rect 158864 147104 192392 147132
rect 158864 147092 158870 147104
rect 192386 147092 192392 147104
rect 192444 147092 192450 147144
rect 105354 147024 105360 147076
rect 105412 147064 105418 147076
rect 138658 147064 138664 147076
rect 105412 147036 138664 147064
rect 105412 147024 105418 147036
rect 138658 147024 138664 147036
rect 138716 147024 138722 147076
rect 160462 147024 160468 147076
rect 160520 147064 160526 147076
rect 195238 147064 195244 147076
rect 160520 147036 195244 147064
rect 160520 147024 160526 147036
rect 195238 147024 195244 147036
rect 195296 147024 195302 147076
rect 112622 146956 112628 147008
rect 112680 146996 112686 147008
rect 112898 146996 112904 147008
rect 112680 146968 112904 146996
rect 112680 146956 112686 146968
rect 112898 146956 112904 146968
rect 112956 146956 112962 147008
rect 141878 146996 141884 147008
rect 113008 146968 141884 146996
rect 106734 146888 106740 146940
rect 106792 146928 106798 146940
rect 113008 146928 113036 146968
rect 141878 146956 141884 146968
rect 141936 146956 141942 147008
rect 161658 146956 161664 147008
rect 161716 146996 161722 147008
rect 197170 146996 197176 147008
rect 161716 146968 197176 146996
rect 161716 146956 161722 146968
rect 197170 146956 197176 146968
rect 197228 146956 197234 147008
rect 138842 146928 138848 146940
rect 106792 146900 113036 146928
rect 113146 146900 138848 146928
rect 106792 146888 106798 146900
rect 103974 146820 103980 146872
rect 104032 146860 104038 146872
rect 113146 146860 113174 146900
rect 138842 146888 138848 146900
rect 138900 146888 138906 146940
rect 174906 146888 174912 146940
rect 174964 146928 174970 146940
rect 214466 146928 214472 146940
rect 174964 146900 214472 146928
rect 174964 146888 174970 146900
rect 214466 146888 214472 146900
rect 214524 146888 214530 146940
rect 104032 146832 113174 146860
rect 104032 146820 104038 146832
rect 126606 146820 126612 146872
rect 126664 146860 126670 146872
rect 126882 146860 126888 146872
rect 126664 146832 126888 146860
rect 126664 146820 126670 146832
rect 126882 146820 126888 146832
rect 126940 146820 126946 146872
rect 179138 146820 179144 146872
rect 179196 146860 179202 146872
rect 179196 146832 180794 146860
rect 179196 146820 179202 146832
rect 180766 146656 180794 146832
rect 185762 146820 185768 146872
rect 185820 146860 185826 146872
rect 186038 146860 186044 146872
rect 185820 146832 186044 146860
rect 185820 146820 185826 146832
rect 186038 146820 186044 146832
rect 186096 146820 186102 146872
rect 181714 146752 181720 146804
rect 181772 146792 181778 146804
rect 187234 146792 187240 146804
rect 181772 146764 187240 146792
rect 181772 146752 181778 146764
rect 187234 146752 187240 146764
rect 187292 146752 187298 146804
rect 191466 146792 191472 146804
rect 190426 146764 191472 146792
rect 183186 146684 183192 146736
rect 183244 146724 183250 146736
rect 189718 146724 189724 146736
rect 183244 146696 189724 146724
rect 183244 146684 183250 146696
rect 189718 146684 189724 146696
rect 189776 146684 189782 146736
rect 189166 146656 189172 146668
rect 180766 146628 189172 146656
rect 189166 146616 189172 146628
rect 189224 146616 189230 146668
rect 181622 146548 181628 146600
rect 181680 146588 181686 146600
rect 190426 146588 190454 146764
rect 191466 146752 191472 146764
rect 191524 146752 191530 146804
rect 181680 146560 190454 146588
rect 181680 146548 181686 146560
rect 113910 146208 113916 146260
rect 113968 146248 113974 146260
rect 129826 146248 129832 146260
rect 113968 146220 129832 146248
rect 113968 146208 113974 146220
rect 129826 146208 129832 146220
rect 129884 146208 129890 146260
rect 178218 146208 178224 146260
rect 178276 146248 178282 146260
rect 191006 146248 191012 146260
rect 178276 146220 191012 146248
rect 178276 146208 178282 146220
rect 191006 146208 191012 146220
rect 191064 146208 191070 146260
rect 113818 146140 113824 146192
rect 113876 146180 113882 146192
rect 131666 146180 131672 146192
rect 113876 146152 131672 146180
rect 113876 146140 113882 146152
rect 131666 146140 131672 146152
rect 131724 146140 131730 146192
rect 178034 146140 178040 146192
rect 178092 146180 178098 146192
rect 199102 146180 199108 146192
rect 178092 146152 199108 146180
rect 178092 146140 178098 146152
rect 199102 146140 199108 146152
rect 199160 146140 199166 146192
rect 112346 146072 112352 146124
rect 112404 146112 112410 146124
rect 131114 146112 131120 146124
rect 112404 146084 131120 146112
rect 112404 146072 112410 146084
rect 131114 146072 131120 146084
rect 131172 146072 131178 146124
rect 177206 146072 177212 146124
rect 177264 146112 177270 146124
rect 197998 146112 198004 146124
rect 177264 146084 198004 146112
rect 177264 146072 177270 146084
rect 197998 146072 198004 146084
rect 198056 146072 198062 146124
rect 111242 146004 111248 146056
rect 111300 146044 111306 146056
rect 129918 146044 129924 146056
rect 111300 146016 129924 146044
rect 111300 146004 111306 146016
rect 129918 146004 129924 146016
rect 129976 146004 129982 146056
rect 173986 146004 173992 146056
rect 174044 146044 174050 146056
rect 197906 146044 197912 146056
rect 174044 146016 197912 146044
rect 174044 146004 174050 146016
rect 197906 146004 197912 146016
rect 197964 146004 197970 146056
rect 122558 145936 122564 145988
rect 122616 145976 122622 145988
rect 149146 145976 149152 145988
rect 122616 145948 149152 145976
rect 122616 145936 122622 145948
rect 149146 145936 149152 145948
rect 149204 145936 149210 145988
rect 169846 145936 169852 145988
rect 169904 145976 169910 145988
rect 195054 145976 195060 145988
rect 169904 145948 195060 145976
rect 169904 145936 169910 145948
rect 195054 145936 195060 145948
rect 195112 145936 195118 145988
rect 120442 145868 120448 145920
rect 120500 145908 120506 145920
rect 148594 145908 148600 145920
rect 120500 145880 148600 145908
rect 120500 145868 120506 145880
rect 148594 145868 148600 145880
rect 148652 145868 148658 145920
rect 165706 145868 165712 145920
rect 165764 145908 165770 145920
rect 196434 145908 196440 145920
rect 165764 145880 196440 145908
rect 165764 145868 165770 145880
rect 196434 145868 196440 145880
rect 196492 145868 196498 145920
rect 116302 145800 116308 145852
rect 116360 145840 116366 145852
rect 145374 145840 145380 145852
rect 116360 145812 145380 145840
rect 116360 145800 116366 145812
rect 145374 145800 145380 145812
rect 145432 145800 145438 145852
rect 153286 145800 153292 145852
rect 153344 145840 153350 145852
rect 186774 145840 186780 145852
rect 153344 145812 186780 145840
rect 153344 145800 153350 145812
rect 186774 145800 186780 145812
rect 186832 145800 186838 145852
rect 116486 145732 116492 145784
rect 116544 145772 116550 145784
rect 147030 145772 147036 145784
rect 116544 145744 147036 145772
rect 116544 145732 116550 145744
rect 147030 145732 147036 145744
rect 147088 145732 147094 145784
rect 161566 145732 161572 145784
rect 161624 145772 161630 145784
rect 197078 145772 197084 145784
rect 161624 145744 197084 145772
rect 161624 145732 161630 145744
rect 197078 145732 197084 145744
rect 197136 145732 197142 145784
rect 113542 145664 113548 145716
rect 113600 145704 113606 145716
rect 146754 145704 146760 145716
rect 113600 145676 146760 145704
rect 113600 145664 113606 145676
rect 146754 145664 146760 145676
rect 146812 145664 146818 145716
rect 162762 145664 162768 145716
rect 162820 145704 162826 145716
rect 197906 145704 197912 145716
rect 162820 145676 197912 145704
rect 162820 145664 162826 145676
rect 197906 145664 197912 145676
rect 197964 145664 197970 145716
rect 115014 145596 115020 145648
rect 115072 145636 115078 145648
rect 147950 145636 147956 145648
rect 115072 145608 147956 145636
rect 115072 145596 115078 145608
rect 147950 145596 147956 145608
rect 148008 145596 148014 145648
rect 166810 145596 166816 145648
rect 166868 145636 166874 145648
rect 214558 145636 214564 145648
rect 166868 145608 214564 145636
rect 166868 145596 166874 145608
rect 214558 145596 214564 145608
rect 214616 145596 214622 145648
rect 3510 145528 3516 145580
rect 3568 145568 3574 145580
rect 3568 145540 161474 145568
rect 3568 145528 3574 145540
rect 115382 145460 115388 145512
rect 115440 145500 115446 145512
rect 129734 145500 129740 145512
rect 115440 145472 129740 145500
rect 115440 145460 115446 145472
rect 129734 145460 129740 145472
rect 129792 145460 129798 145512
rect 115290 145392 115296 145444
rect 115348 145432 115354 145444
rect 130654 145432 130660 145444
rect 115348 145404 130660 145432
rect 115348 145392 115354 145404
rect 130654 145392 130660 145404
rect 130712 145392 130718 145444
rect 161446 145432 161474 145540
rect 179414 145528 179420 145580
rect 179472 145568 179478 145580
rect 190914 145568 190920 145580
rect 179472 145540 190920 145568
rect 179472 145528 179478 145540
rect 190914 145528 190920 145540
rect 190972 145528 190978 145580
rect 178310 145460 178316 145512
rect 178368 145500 178374 145512
rect 189626 145500 189632 145512
rect 178368 145472 189632 145500
rect 178368 145460 178374 145472
rect 189626 145460 189632 145472
rect 189684 145460 189690 145512
rect 179506 145432 179512 145444
rect 161446 145404 179512 145432
rect 179506 145392 179512 145404
rect 179564 145432 179570 145444
rect 189534 145432 189540 145444
rect 179564 145404 189540 145432
rect 179564 145392 179570 145404
rect 189534 145392 189540 145404
rect 189592 145392 189598 145444
rect 113818 145324 113824 145376
rect 113876 145364 113882 145376
rect 127802 145364 127808 145376
rect 113876 145336 127808 145364
rect 113876 145324 113882 145336
rect 127802 145324 127808 145336
rect 127860 145324 127866 145376
rect 183738 145324 183744 145376
rect 183796 145364 183802 145376
rect 194226 145364 194232 145376
rect 183796 145336 194232 145364
rect 183796 145324 183802 145336
rect 194226 145324 194232 145336
rect 194284 145324 194290 145376
rect 185670 144916 185676 144968
rect 185728 144956 185734 144968
rect 185728 144928 187924 144956
rect 185728 144916 185734 144928
rect 115842 144848 115848 144900
rect 115900 144888 115906 144900
rect 115900 144860 122834 144888
rect 115900 144848 115906 144860
rect 122806 144684 122834 144860
rect 184014 144848 184020 144900
rect 184072 144888 184078 144900
rect 187786 144888 187792 144900
rect 184072 144860 187792 144888
rect 184072 144848 184078 144860
rect 187786 144848 187792 144860
rect 187844 144848 187850 144900
rect 187896 144888 187924 144928
rect 199562 144888 199568 144900
rect 187896 144860 199568 144888
rect 199562 144848 199568 144860
rect 199620 144848 199626 144900
rect 181530 144780 181536 144832
rect 181588 144820 181594 144832
rect 188062 144820 188068 144832
rect 181588 144792 188068 144820
rect 181588 144780 181594 144792
rect 188062 144780 188068 144792
rect 188120 144780 188126 144832
rect 188246 144780 188252 144832
rect 188304 144820 188310 144832
rect 198182 144820 198188 144832
rect 188304 144792 198188 144820
rect 188304 144780 188310 144792
rect 198182 144780 198188 144792
rect 198240 144780 198246 144832
rect 173802 144712 173808 144764
rect 173860 144752 173866 144764
rect 192110 144752 192116 144764
rect 173860 144724 192116 144752
rect 173860 144712 173866 144724
rect 192110 144712 192116 144724
rect 192168 144712 192174 144764
rect 133874 144684 133880 144696
rect 122806 144656 133880 144684
rect 133874 144644 133880 144656
rect 133932 144644 133938 144696
rect 170582 144644 170588 144696
rect 170640 144684 170646 144696
rect 192294 144684 192300 144696
rect 170640 144656 192300 144684
rect 170640 144644 170646 144656
rect 192294 144644 192300 144656
rect 192352 144644 192358 144696
rect 117774 144576 117780 144628
rect 117832 144616 117838 144628
rect 143626 144616 143632 144628
rect 117832 144588 143632 144616
rect 117832 144576 117838 144588
rect 143626 144576 143632 144588
rect 143684 144576 143690 144628
rect 172422 144576 172428 144628
rect 172480 144616 172486 144628
rect 193674 144616 193680 144628
rect 172480 144588 193680 144616
rect 172480 144576 172486 144588
rect 193674 144576 193680 144588
rect 193732 144576 193738 144628
rect 115566 144508 115572 144560
rect 115624 144548 115630 144560
rect 140866 144548 140872 144560
rect 115624 144520 140872 144548
rect 115624 144508 115630 144520
rect 140866 144508 140872 144520
rect 140924 144508 140930 144560
rect 169110 144508 169116 144560
rect 169168 144548 169174 144560
rect 193582 144548 193588 144560
rect 169168 144520 193588 144548
rect 169168 144508 169174 144520
rect 193582 144508 193588 144520
rect 193640 144508 193646 144560
rect 117774 144440 117780 144492
rect 117832 144480 117838 144492
rect 148226 144480 148232 144492
rect 117832 144452 148232 144480
rect 117832 144440 117838 144452
rect 148226 144440 148232 144452
rect 148284 144440 148290 144492
rect 168006 144440 168012 144492
rect 168064 144480 168070 144492
rect 194962 144480 194968 144492
rect 168064 144452 194968 144480
rect 168064 144440 168070 144452
rect 194962 144440 194968 144452
rect 195020 144440 195026 144492
rect 111242 144372 111248 144424
rect 111300 144412 111306 144424
rect 142522 144412 142528 144424
rect 111300 144384 142528 144412
rect 111300 144372 111306 144384
rect 142522 144372 142528 144384
rect 142580 144372 142586 144424
rect 160278 144372 160284 144424
rect 160336 144412 160342 144424
rect 189810 144412 189816 144424
rect 160336 144384 189816 144412
rect 160336 144372 160342 144384
rect 189810 144372 189816 144384
rect 189868 144372 189874 144424
rect 118786 144304 118792 144356
rect 118844 144344 118850 144356
rect 151906 144344 151912 144356
rect 118844 144316 151912 144344
rect 118844 144304 118850 144316
rect 151906 144304 151912 144316
rect 151964 144304 151970 144356
rect 154666 144304 154672 144356
rect 154724 144344 154730 144356
rect 188798 144344 188804 144356
rect 154724 144316 188804 144344
rect 154724 144304 154730 144316
rect 188798 144304 188804 144316
rect 188856 144304 188862 144356
rect 111426 144236 111432 144288
rect 111484 144276 111490 144288
rect 131206 144276 131212 144288
rect 111484 144248 131212 144276
rect 111484 144236 111490 144248
rect 131206 144236 131212 144248
rect 131264 144276 131270 144288
rect 131264 144248 183232 144276
rect 131264 144236 131270 144248
rect 118142 144168 118148 144220
rect 118200 144208 118206 144220
rect 130194 144208 130200 144220
rect 118200 144180 130200 144208
rect 118200 144168 118206 144180
rect 130194 144168 130200 144180
rect 130252 144208 130258 144220
rect 183204 144208 183232 144248
rect 183278 144236 183284 144288
rect 183336 144276 183342 144288
rect 188246 144276 188252 144288
rect 183336 144248 188252 144276
rect 183336 144236 183342 144248
rect 188246 144236 188252 144248
rect 188304 144236 188310 144288
rect 188338 144208 188344 144220
rect 130252 144180 180794 144208
rect 183204 144180 188344 144208
rect 130252 144168 130258 144180
rect 180766 144072 180794 144180
rect 188338 144168 188344 144180
rect 188396 144168 188402 144220
rect 182082 144100 182088 144152
rect 182140 144140 182146 144152
rect 195054 144140 195060 144152
rect 182140 144112 195060 144140
rect 182140 144100 182146 144112
rect 195054 144100 195060 144112
rect 195112 144100 195118 144152
rect 189902 144072 189908 144084
rect 180766 144044 189908 144072
rect 189902 144032 189908 144044
rect 189960 144032 189966 144084
rect 118142 143692 118148 143744
rect 118200 143732 118206 143744
rect 145282 143732 145288 143744
rect 118200 143704 145288 143732
rect 118200 143692 118206 143704
rect 145282 143692 145288 143704
rect 145340 143692 145346 143744
rect 117222 143624 117228 143676
rect 117280 143664 117286 143676
rect 148594 143664 148600 143676
rect 117280 143636 148600 143664
rect 117280 143624 117286 143636
rect 148594 143624 148600 143636
rect 148652 143624 148658 143676
rect 112898 143556 112904 143608
rect 112956 143596 112962 143608
rect 145834 143596 145840 143608
rect 112956 143568 145840 143596
rect 112956 143556 112962 143568
rect 145834 143556 145840 143568
rect 145892 143556 145898 143608
rect 177114 143488 177120 143540
rect 177172 143528 177178 143540
rect 179414 143528 179420 143540
rect 177172 143500 179420 143528
rect 177172 143488 177178 143500
rect 179414 143488 179420 143500
rect 179472 143488 179478 143540
rect 183002 143488 183008 143540
rect 183060 143528 183066 143540
rect 187418 143528 187424 143540
rect 183060 143500 187424 143528
rect 183060 143488 183066 143500
rect 187418 143488 187424 143500
rect 187476 143488 187482 143540
rect 186038 143420 186044 143472
rect 186096 143460 186102 143472
rect 187510 143460 187516 143472
rect 186096 143432 187516 143460
rect 186096 143420 186102 143432
rect 187510 143420 187516 143432
rect 187568 143420 187574 143472
rect 116670 143352 116676 143404
rect 116728 143392 116734 143404
rect 128538 143392 128544 143404
rect 116728 143364 128544 143392
rect 116728 143352 116734 143364
rect 128538 143352 128544 143364
rect 128596 143352 128602 143404
rect 129826 143352 129832 143404
rect 129884 143392 129890 143404
rect 135438 143392 135444 143404
rect 129884 143364 135444 143392
rect 129884 143352 129890 143364
rect 135438 143352 135444 143364
rect 135496 143352 135502 143404
rect 185486 143352 185492 143404
rect 185544 143392 185550 143404
rect 191282 143392 191288 143404
rect 185544 143364 191288 143392
rect 185544 143352 185550 143364
rect 191282 143352 191288 143364
rect 191340 143352 191346 143404
rect 116762 143284 116768 143336
rect 116820 143324 116826 143336
rect 131482 143324 131488 143336
rect 116820 143296 131488 143324
rect 116820 143284 116826 143296
rect 131482 143284 131488 143296
rect 131540 143284 131546 143336
rect 182726 143284 182732 143336
rect 182784 143324 182790 143336
rect 197814 143324 197820 143336
rect 182784 143296 197820 143324
rect 182784 143284 182790 143296
rect 197814 143284 197820 143296
rect 197872 143284 197878 143336
rect 118050 143216 118056 143268
rect 118108 143256 118114 143268
rect 133138 143256 133144 143268
rect 118108 143228 133144 143256
rect 118108 143216 118114 143228
rect 133138 143216 133144 143228
rect 133196 143216 133202 143268
rect 175642 143216 175648 143268
rect 175700 143256 175706 143268
rect 192018 143256 192024 143268
rect 175700 143228 192024 143256
rect 175700 143216 175706 143228
rect 192018 143216 192024 143228
rect 192076 143216 192082 143268
rect 112254 143148 112260 143200
rect 112312 143188 112318 143200
rect 127710 143188 127716 143200
rect 112312 143160 127716 143188
rect 112312 143148 112318 143160
rect 127710 143148 127716 143160
rect 127768 143148 127774 143200
rect 129734 143148 129740 143200
rect 129792 143188 129798 143200
rect 137002 143188 137008 143200
rect 129792 143160 137008 143188
rect 129792 143148 129798 143160
rect 137002 143148 137008 143160
rect 137060 143148 137066 143200
rect 173526 143148 173532 143200
rect 173584 143188 173590 143200
rect 189350 143188 189356 143200
rect 173584 143160 189356 143188
rect 173584 143148 173590 143160
rect 189350 143148 189356 143160
rect 189408 143148 189414 143200
rect 120810 143080 120816 143132
rect 120868 143120 120874 143132
rect 139762 143120 139768 143132
rect 120868 143092 139768 143120
rect 120868 143080 120874 143092
rect 139762 143080 139768 143092
rect 139820 143080 139826 143132
rect 168282 143080 168288 143132
rect 168340 143120 168346 143132
rect 190822 143120 190828 143132
rect 168340 143092 190828 143120
rect 168340 143080 168346 143092
rect 190822 143080 190828 143092
rect 190880 143080 190886 143132
rect 120902 143012 120908 143064
rect 120960 143052 120966 143064
rect 141418 143052 141424 143064
rect 120960 143024 141424 143052
rect 120960 143012 120966 143024
rect 141418 143012 141424 143024
rect 141476 143012 141482 143064
rect 155954 143012 155960 143064
rect 156012 143052 156018 143064
rect 184198 143052 184204 143064
rect 156012 143024 184204 143052
rect 156012 143012 156018 143024
rect 184198 143012 184204 143024
rect 184256 143012 184262 143064
rect 185670 143012 185676 143064
rect 185728 143052 185734 143064
rect 196526 143052 196532 143064
rect 185728 143024 196532 143052
rect 185728 143012 185734 143024
rect 196526 143012 196532 143024
rect 196584 143012 196590 143064
rect 120718 142944 120724 142996
rect 120776 142984 120782 142996
rect 151446 142984 151452 142996
rect 120776 142956 151452 142984
rect 120776 142944 120782 142956
rect 151446 142944 151452 142956
rect 151504 142944 151510 142996
rect 158622 142944 158628 142996
rect 158680 142984 158686 142996
rect 187970 142984 187976 142996
rect 158680 142956 187976 142984
rect 158680 142944 158686 142956
rect 187970 142944 187976 142956
rect 188028 142944 188034 142996
rect 119798 142876 119804 142928
rect 119856 142916 119862 142928
rect 143074 142916 143080 142928
rect 119856 142888 143080 142916
rect 119856 142876 119862 142888
rect 143074 142876 143080 142888
rect 143132 142876 143138 142928
rect 178862 142876 178868 142928
rect 178920 142916 178926 142928
rect 214650 142916 214656 142928
rect 178920 142888 214656 142916
rect 178920 142876 178926 142888
rect 214650 142876 214656 142888
rect 214708 142876 214714 142928
rect 119522 142808 119528 142860
rect 119580 142848 119586 142860
rect 149698 142848 149704 142860
rect 119580 142820 149704 142848
rect 119580 142808 119586 142820
rect 149698 142808 149704 142820
rect 149756 142808 149762 142860
rect 151262 142808 151268 142860
rect 151320 142848 151326 142860
rect 209222 142848 209228 142860
rect 151320 142820 209228 142848
rect 151320 142808 151326 142820
rect 209222 142808 209228 142820
rect 209280 142808 209286 142860
rect 177942 142536 177948 142588
rect 178000 142576 178006 142588
rect 184474 142576 184480 142588
rect 178000 142548 184480 142576
rect 178000 142536 178006 142548
rect 184474 142536 184480 142548
rect 184532 142536 184538 142588
rect 128262 142468 128268 142520
rect 128320 142508 128326 142520
rect 580718 142508 580724 142520
rect 128320 142480 580724 142508
rect 128320 142468 128326 142480
rect 580718 142468 580724 142480
rect 580776 142468 580782 142520
rect 128538 142400 128544 142452
rect 128596 142440 128602 142452
rect 133506 142440 133512 142452
rect 128596 142412 133512 142440
rect 128596 142400 128602 142412
rect 133506 142400 133512 142412
rect 133564 142400 133570 142452
rect 182726 142440 182732 142452
rect 161446 142412 182732 142440
rect 119522 142332 119528 142384
rect 119580 142372 119586 142384
rect 161446 142372 161474 142412
rect 182726 142400 182732 142412
rect 182784 142400 182790 142452
rect 119580 142344 161474 142372
rect 119580 142332 119586 142344
rect 177850 142332 177856 142384
rect 177908 142372 177914 142384
rect 181990 142372 181996 142384
rect 177908 142344 181996 142372
rect 177908 142332 177914 142344
rect 181990 142332 181996 142344
rect 182048 142332 182054 142384
rect 120166 142264 120172 142316
rect 120224 142304 120230 142316
rect 186038 142304 186044 142316
rect 120224 142276 186044 142304
rect 120224 142264 120230 142276
rect 186038 142264 186044 142276
rect 186096 142264 186102 142316
rect 129918 142196 129924 142248
rect 129976 142236 129982 142248
rect 132586 142236 132592 142248
rect 129976 142208 132592 142236
rect 129976 142196 129982 142208
rect 132586 142196 132592 142208
rect 132644 142196 132650 142248
rect 133506 142196 133512 142248
rect 133564 142236 133570 142248
rect 580902 142236 580908 142248
rect 133564 142208 580908 142236
rect 133564 142196 133570 142208
rect 580902 142196 580908 142208
rect 580960 142196 580966 142248
rect 131114 142128 131120 142180
rect 131172 142168 131178 142180
rect 134242 142168 134248 142180
rect 131172 142140 134248 142168
rect 131172 142128 131178 142140
rect 134242 142128 134248 142140
rect 134300 142128 134306 142180
rect 150526 142168 150532 142180
rect 148888 142140 150532 142168
rect 115842 142060 115848 142112
rect 115900 142100 115906 142112
rect 148888 142100 148916 142140
rect 150526 142128 150532 142140
rect 150584 142128 150590 142180
rect 155770 142128 155776 142180
rect 155828 142168 155834 142180
rect 157426 142168 157432 142180
rect 155828 142140 157432 142168
rect 155828 142128 155834 142140
rect 157426 142128 157432 142140
rect 157484 142128 157490 142180
rect 183646 142128 183652 142180
rect 183704 142168 183710 142180
rect 191006 142168 191012 142180
rect 183704 142140 191012 142168
rect 183704 142128 183710 142140
rect 191006 142128 191012 142140
rect 191064 142128 191070 142180
rect 115900 142072 148916 142100
rect 115900 142060 115906 142072
rect 185946 142060 185952 142112
rect 186004 142100 186010 142112
rect 195330 142100 195336 142112
rect 186004 142072 195336 142100
rect 186004 142060 186010 142072
rect 195330 142060 195336 142072
rect 195388 142060 195394 142112
rect 116394 141992 116400 142044
rect 116452 142032 116458 142044
rect 127802 142032 127808 142044
rect 116452 142004 127808 142032
rect 116452 141992 116458 142004
rect 127802 141992 127808 142004
rect 127860 141992 127866 142044
rect 176470 141992 176476 142044
rect 176528 142032 176534 142044
rect 187326 142032 187332 142044
rect 176528 142004 187332 142032
rect 176528 141992 176534 142004
rect 187326 141992 187332 142004
rect 187384 141992 187390 142044
rect 111242 141924 111248 141976
rect 111300 141964 111306 141976
rect 123478 141964 123484 141976
rect 111300 141936 123484 141964
rect 111300 141924 111306 141936
rect 123478 141924 123484 141936
rect 123536 141924 123542 141976
rect 128906 141924 128912 141976
rect 128964 141964 128970 141976
rect 129274 141964 129280 141976
rect 128964 141936 129280 141964
rect 128964 141924 128970 141936
rect 129274 141924 129280 141936
rect 129332 141924 129338 141976
rect 175182 141924 175188 141976
rect 175240 141964 175246 141976
rect 187878 141964 187884 141976
rect 175240 141936 187884 141964
rect 175240 141924 175246 141936
rect 187878 141924 187884 141936
rect 187936 141924 187942 141976
rect 114002 141856 114008 141908
rect 114060 141896 114066 141908
rect 127342 141896 127348 141908
rect 114060 141868 127348 141896
rect 114060 141856 114066 141868
rect 127342 141856 127348 141868
rect 127400 141856 127406 141908
rect 180334 141856 180340 141908
rect 180392 141896 180398 141908
rect 193490 141896 193496 141908
rect 180392 141868 193496 141896
rect 180392 141856 180398 141868
rect 193490 141856 193496 141868
rect 193548 141856 193554 141908
rect 112622 141788 112628 141840
rect 112680 141828 112686 141840
rect 129274 141828 129280 141840
rect 112680 141800 129280 141828
rect 112680 141788 112686 141800
rect 129274 141788 129280 141800
rect 129332 141788 129338 141840
rect 176194 141788 176200 141840
rect 176252 141828 176258 141840
rect 182910 141828 182916 141840
rect 176252 141800 182916 141828
rect 176252 141788 176258 141800
rect 182910 141788 182916 141800
rect 182968 141788 182974 141840
rect 185578 141788 185584 141840
rect 185636 141828 185642 141840
rect 185946 141828 185952 141840
rect 185636 141800 185952 141828
rect 185636 141788 185642 141800
rect 185946 141788 185952 141800
rect 186004 141788 186010 141840
rect 117958 141720 117964 141772
rect 118016 141760 118022 141772
rect 134794 141760 134800 141772
rect 118016 141732 134800 141760
rect 118016 141720 118022 141732
rect 134794 141720 134800 141732
rect 134852 141720 134858 141772
rect 170214 141720 170220 141772
rect 170272 141760 170278 141772
rect 189442 141760 189448 141772
rect 170272 141732 189448 141760
rect 170272 141720 170278 141732
rect 189442 141720 189448 141732
rect 189500 141720 189506 141772
rect 117866 141652 117872 141704
rect 117924 141692 117930 141704
rect 117924 141664 127756 141692
rect 117924 141652 117930 141664
rect 119614 141584 119620 141636
rect 119672 141624 119678 141636
rect 127728 141624 127756 141664
rect 127802 141652 127808 141704
rect 127860 141692 127866 141704
rect 136634 141692 136640 141704
rect 127860 141664 136640 141692
rect 127860 141652 127866 141664
rect 136634 141652 136640 141664
rect 136692 141652 136698 141704
rect 171870 141652 171876 141704
rect 171928 141692 171934 141704
rect 190730 141692 190736 141704
rect 171928 141664 190736 141692
rect 171928 141652 171934 141664
rect 190730 141652 190736 141664
rect 190788 141652 190794 141704
rect 140314 141624 140320 141636
rect 119672 141596 127664 141624
rect 127728 141596 140320 141624
rect 119672 141584 119678 141596
rect 119338 141516 119344 141568
rect 119396 141556 119402 141568
rect 124858 141556 124864 141568
rect 119396 141528 124864 141556
rect 119396 141516 119402 141528
rect 124858 141516 124864 141528
rect 124916 141516 124922 141568
rect 127636 141556 127664 141596
rect 140314 141584 140320 141596
rect 140372 141584 140378 141636
rect 163958 141584 163964 141636
rect 164016 141624 164022 141636
rect 188522 141624 188528 141636
rect 164016 141596 188528 141624
rect 164016 141584 164022 141596
rect 188522 141584 188528 141596
rect 188580 141584 188586 141636
rect 153654 141556 153660 141568
rect 127636 141528 153660 141556
rect 153654 141516 153660 141528
rect 153712 141516 153718 141568
rect 160186 141516 160192 141568
rect 160244 141556 160250 141568
rect 186958 141556 186964 141568
rect 160244 141528 186964 141556
rect 160244 141516 160250 141528
rect 186958 141516 186964 141528
rect 187016 141516 187022 141568
rect 117222 141448 117228 141500
rect 117280 141488 117286 141500
rect 142246 141488 142252 141500
rect 117280 141460 142252 141488
rect 117280 141448 117286 141460
rect 142246 141448 142252 141460
rect 142304 141448 142310 141500
rect 169294 141448 169300 141500
rect 169352 141488 169358 141500
rect 196250 141488 196256 141500
rect 169352 141460 196256 141488
rect 169352 141448 169358 141460
rect 196250 141448 196256 141460
rect 196308 141448 196314 141500
rect 119430 141380 119436 141432
rect 119488 141420 119494 141432
rect 149422 141420 149428 141432
rect 119488 141392 149428 141420
rect 119488 141380 119494 141392
rect 149422 141380 149428 141392
rect 149480 141380 149486 141432
rect 154206 141380 154212 141432
rect 154264 141420 154270 141432
rect 187142 141420 187148 141432
rect 154264 141392 187148 141420
rect 154264 141380 154270 141392
rect 187142 141380 187148 141392
rect 187200 141380 187206 141432
rect 182910 141312 182916 141364
rect 182968 141352 182974 141364
rect 192294 141352 192300 141364
rect 182968 141324 192300 141352
rect 182968 141312 182974 141324
rect 192294 141312 192300 141324
rect 192352 141312 192358 141364
rect 184106 141108 184112 141160
rect 184164 141148 184170 141160
rect 189626 141148 189632 141160
rect 184164 141120 189632 141148
rect 184164 141108 184170 141120
rect 189626 141108 189632 141120
rect 189684 141108 189690 141160
rect 13078 140836 13084 140888
rect 13136 140876 13142 140888
rect 182818 140876 182824 140888
rect 13136 140848 182824 140876
rect 13136 140836 13142 140848
rect 182818 140836 182824 140848
rect 182876 140836 182882 140888
rect 184198 140836 184204 140888
rect 184256 140876 184262 140888
rect 187326 140876 187332 140888
rect 184256 140848 187332 140876
rect 184256 140836 184262 140848
rect 187326 140836 187332 140848
rect 187384 140836 187390 140888
rect 127342 140768 127348 140820
rect 127400 140808 127406 140820
rect 580810 140808 580816 140820
rect 127400 140780 580816 140808
rect 127400 140768 127406 140780
rect 580810 140768 580816 140780
rect 580868 140768 580874 140820
rect 119706 140700 119712 140752
rect 119764 140740 119770 140752
rect 126238 140740 126244 140752
rect 119764 140712 126244 140740
rect 119764 140700 119770 140712
rect 126238 140700 126244 140712
rect 126296 140700 126302 140752
rect 158714 140700 158720 140752
rect 158772 140740 158778 140752
rect 159634 140740 159640 140752
rect 158772 140712 159640 140740
rect 158772 140700 158778 140712
rect 159634 140700 159640 140712
rect 159692 140700 159698 140752
rect 193490 140740 193496 140752
rect 161446 140712 193496 140740
rect 159542 140632 159548 140684
rect 159600 140672 159606 140684
rect 161446 140672 161474 140712
rect 193490 140700 193496 140712
rect 193548 140700 193554 140752
rect 159600 140644 161474 140672
rect 159600 140632 159606 140644
rect 161842 140632 161848 140684
rect 161900 140672 161906 140684
rect 162394 140672 162400 140684
rect 161900 140644 162400 140672
rect 161900 140632 161906 140644
rect 162394 140632 162400 140644
rect 162452 140632 162458 140684
rect 169846 140632 169852 140684
rect 169904 140672 169910 140684
rect 170674 140672 170680 140684
rect 169904 140644 170680 140672
rect 169904 140632 169910 140644
rect 170674 140632 170680 140644
rect 170732 140632 170738 140684
rect 178034 140632 178040 140684
rect 178092 140672 178098 140684
rect 178954 140672 178960 140684
rect 178092 140644 178960 140672
rect 178092 140632 178098 140644
rect 178954 140632 178960 140644
rect 179012 140632 179018 140684
rect 119246 140564 119252 140616
rect 119304 140604 119310 140616
rect 126698 140604 126704 140616
rect 119304 140576 126704 140604
rect 119304 140564 119310 140576
rect 126698 140564 126704 140576
rect 126756 140564 126762 140616
rect 173894 140564 173900 140616
rect 173952 140604 173958 140616
rect 189074 140604 189080 140616
rect 173952 140576 189080 140604
rect 173952 140564 173958 140576
rect 189074 140564 189080 140576
rect 189132 140564 189138 140616
rect 120902 140496 120908 140548
rect 120960 140536 120966 140548
rect 129182 140536 129188 140548
rect 120960 140508 129188 140536
rect 120960 140496 120966 140508
rect 129182 140496 129188 140508
rect 129240 140496 129246 140548
rect 184842 140496 184848 140548
rect 184900 140536 184906 140548
rect 192478 140536 192484 140548
rect 184900 140508 192484 140536
rect 184900 140496 184906 140508
rect 192478 140496 192484 140508
rect 192536 140496 192542 140548
rect 119338 140428 119344 140480
rect 119396 140468 119402 140480
rect 127618 140468 127624 140480
rect 119396 140440 127624 140468
rect 119396 140428 119402 140440
rect 127618 140428 127624 140440
rect 127676 140428 127682 140480
rect 178770 140428 178776 140480
rect 178828 140468 178834 140480
rect 187970 140468 187976 140480
rect 178828 140440 187976 140468
rect 178828 140428 178834 140440
rect 187970 140428 187976 140440
rect 188028 140428 188034 140480
rect 118142 140360 118148 140412
rect 118200 140400 118206 140412
rect 126422 140400 126428 140412
rect 118200 140372 126428 140400
rect 118200 140360 118206 140372
rect 126422 140360 126428 140372
rect 126480 140360 126486 140412
rect 180058 140360 180064 140412
rect 180116 140400 180122 140412
rect 189350 140400 189356 140412
rect 180116 140372 189356 140400
rect 180116 140360 180122 140372
rect 189350 140360 189356 140372
rect 189408 140360 189414 140412
rect 117958 140292 117964 140344
rect 118016 140332 118022 140344
rect 129366 140332 129372 140344
rect 118016 140304 129372 140332
rect 118016 140292 118022 140304
rect 129366 140292 129372 140304
rect 129424 140292 129430 140344
rect 178678 140292 178684 140344
rect 178736 140332 178742 140344
rect 188338 140332 188344 140344
rect 178736 140304 188344 140332
rect 178736 140292 178742 140304
rect 188338 140292 188344 140304
rect 188396 140292 188402 140344
rect 116670 140224 116676 140276
rect 116728 140264 116734 140276
rect 129090 140264 129096 140276
rect 116728 140236 129096 140264
rect 116728 140224 116734 140236
rect 129090 140224 129096 140236
rect 129148 140224 129154 140276
rect 180242 140224 180248 140276
rect 180300 140264 180306 140276
rect 190730 140264 190736 140276
rect 180300 140236 190736 140264
rect 180300 140224 180306 140236
rect 190730 140224 190736 140236
rect 190788 140224 190794 140276
rect 115290 140156 115296 140208
rect 115348 140196 115354 140208
rect 146662 140196 146668 140208
rect 115348 140168 146668 140196
rect 115348 140156 115354 140168
rect 146662 140156 146668 140168
rect 146720 140156 146726 140208
rect 185854 140156 185860 140208
rect 185912 140196 185918 140208
rect 196802 140196 196808 140208
rect 185912 140168 196808 140196
rect 185912 140156 185918 140168
rect 196802 140156 196808 140168
rect 196860 140156 196866 140208
rect 116394 140088 116400 140140
rect 116452 140128 116458 140140
rect 148134 140128 148140 140140
rect 116452 140100 148140 140128
rect 116452 140088 116458 140100
rect 148134 140088 148140 140100
rect 148192 140088 148198 140140
rect 185946 140088 185952 140140
rect 186004 140128 186010 140140
rect 202322 140128 202328 140140
rect 186004 140100 202328 140128
rect 186004 140088 186010 140100
rect 202322 140088 202328 140100
rect 202380 140088 202386 140140
rect 113634 140020 113640 140072
rect 113692 140060 113698 140072
rect 126514 140060 126520 140072
rect 113692 140032 126520 140060
rect 113692 140020 113698 140032
rect 126514 140020 126520 140032
rect 126572 140020 126578 140072
rect 132494 140020 132500 140072
rect 132552 140060 132558 140072
rect 189902 140060 189908 140072
rect 132552 140032 189908 140060
rect 132552 140020 132558 140032
rect 189902 140020 189908 140032
rect 189960 140020 189966 140072
rect 118050 139952 118056 140004
rect 118108 139992 118114 140004
rect 125042 139992 125048 140004
rect 118108 139964 125048 139992
rect 118108 139952 118114 139964
rect 125042 139952 125048 139964
rect 125100 139952 125106 140004
rect 184566 139952 184572 140004
rect 184624 139992 184630 140004
rect 189442 139992 189448 140004
rect 184624 139964 189448 139992
rect 184624 139952 184630 139964
rect 189442 139952 189448 139964
rect 189500 139952 189506 140004
rect 129458 139680 129464 139732
rect 129516 139720 129522 139732
rect 187694 139720 187700 139732
rect 129516 139692 187700 139720
rect 129516 139680 129522 139692
rect 187694 139680 187700 139692
rect 187752 139680 187758 139732
rect 118694 139612 118700 139664
rect 118752 139652 118758 139664
rect 180058 139652 180064 139664
rect 118752 139624 180064 139652
rect 118752 139612 118758 139624
rect 180058 139612 180064 139624
rect 180116 139612 180122 139664
rect 21358 139544 21364 139596
rect 21416 139584 21422 139596
rect 185026 139584 185032 139596
rect 21416 139556 185032 139584
rect 21416 139544 21422 139556
rect 185026 139544 185032 139556
rect 185084 139544 185090 139596
rect 8938 139476 8944 139528
rect 8996 139516 9002 139528
rect 181162 139516 181168 139528
rect 8996 139488 181168 139516
rect 8996 139476 9002 139488
rect 181162 139476 181168 139488
rect 181220 139476 181226 139528
rect 126054 139408 126060 139460
rect 126112 139448 126118 139460
rect 327718 139448 327724 139460
rect 126112 139420 327724 139448
rect 126112 139408 126118 139420
rect 327718 139408 327724 139420
rect 327776 139408 327782 139460
rect 123018 139340 123024 139392
rect 123076 139380 123082 139392
rect 123662 139380 123668 139392
rect 123076 139352 123668 139380
rect 123076 139340 123082 139352
rect 123662 139340 123668 139352
rect 123720 139340 123726 139392
rect 3418 138660 3424 138712
rect 3476 138700 3482 138712
rect 120166 138700 120172 138712
rect 3476 138672 120172 138700
rect 3476 138660 3482 138672
rect 120166 138660 120172 138672
rect 120224 138660 120230 138712
rect 188614 138660 188620 138712
rect 188672 138700 188678 138712
rect 197998 138700 198004 138712
rect 188672 138672 198004 138700
rect 188672 138660 188678 138672
rect 197998 138660 198004 138672
rect 198056 138660 198062 138712
rect 3234 137912 3240 137964
rect 3292 137952 3298 137964
rect 118694 137952 118700 137964
rect 3292 137924 118700 137952
rect 3292 137912 3298 137924
rect 118694 137912 118700 137924
rect 118752 137912 118758 137964
rect 186866 137776 186872 137828
rect 186924 137816 186930 137828
rect 187418 137816 187424 137828
rect 186924 137788 187424 137816
rect 186924 137776 186930 137788
rect 187418 137776 187424 137788
rect 187476 137776 187482 137828
rect 117774 136416 117780 136468
rect 117832 136456 117838 136468
rect 118142 136456 118148 136468
rect 117832 136428 118148 136456
rect 117832 136416 117838 136428
rect 118142 136416 118148 136428
rect 118200 136416 118206 136468
rect 3050 111392 3056 111444
rect 3108 111432 3114 111444
rect 8938 111432 8944 111444
rect 3108 111404 8944 111432
rect 3108 111392 3114 111404
rect 8938 111392 8944 111404
rect 8996 111392 9002 111444
rect 211798 88952 211804 89004
rect 211856 88992 211862 89004
rect 212074 88992 212080 89004
rect 211856 88964 212080 88992
rect 211856 88952 211862 88964
rect 212074 88952 212080 88964
rect 212132 88952 212138 89004
rect 464338 86912 464344 86964
rect 464396 86952 464402 86964
rect 579614 86952 579620 86964
rect 464396 86924 579620 86952
rect 464396 86912 464402 86924
rect 579614 86912 579620 86924
rect 579672 86912 579678 86964
rect 140746 81348 143534 81376
rect 140746 81240 140774 81348
rect 143506 81308 143534 81348
rect 143506 81280 144914 81308
rect 136606 81212 140774 81240
rect 109586 81064 109592 81116
rect 109644 81104 109650 81116
rect 122006 81104 122012 81116
rect 109644 81076 122012 81104
rect 109644 81064 109650 81076
rect 122006 81064 122012 81076
rect 122064 81064 122070 81116
rect 136606 81104 136634 81212
rect 133846 81076 136634 81104
rect 133846 81036 133874 81076
rect 121426 81008 133874 81036
rect 116302 80928 116308 80980
rect 116360 80968 116366 80980
rect 121426 80968 121454 81008
rect 144886 80968 144914 81280
rect 188430 81104 188436 81116
rect 183664 81076 188436 81104
rect 183664 81036 183692 81076
rect 188430 81064 188436 81076
rect 188488 81064 188494 81116
rect 176626 81008 183692 81036
rect 186148 81008 193214 81036
rect 116360 80940 121454 80968
rect 133846 80940 136634 80968
rect 144886 80940 146754 80968
rect 116360 80928 116366 80940
rect 115198 80860 115204 80912
rect 115256 80900 115262 80912
rect 133846 80900 133874 80940
rect 115256 80872 133874 80900
rect 115256 80860 115262 80872
rect 111058 80792 111064 80844
rect 111116 80832 111122 80844
rect 111116 80804 132264 80832
rect 111116 80792 111122 80804
rect 111150 80724 111156 80776
rect 111208 80764 111214 80776
rect 122282 80764 122288 80776
rect 111208 80736 122288 80764
rect 111208 80724 111214 80736
rect 122282 80724 122288 80736
rect 122340 80724 122346 80776
rect 108298 80656 108304 80708
rect 108356 80696 108362 80708
rect 108356 80668 121454 80696
rect 108356 80656 108362 80668
rect 121426 80628 121454 80668
rect 132236 80640 132264 80804
rect 131022 80628 131028 80640
rect 121426 80600 131028 80628
rect 131022 80588 131028 80600
rect 131080 80588 131086 80640
rect 132218 80588 132224 80640
rect 132276 80588 132282 80640
rect 136606 80628 136634 80940
rect 144886 80736 145558 80764
rect 144886 80628 144914 80736
rect 136606 80600 144914 80628
rect 121914 80520 121920 80572
rect 121972 80560 121978 80572
rect 121972 80532 144914 80560
rect 121972 80520 121978 80532
rect 122282 80452 122288 80504
rect 122340 80492 122346 80504
rect 122340 80464 143534 80492
rect 122340 80452 122346 80464
rect 105262 80248 105268 80300
rect 105320 80288 105326 80300
rect 105630 80288 105636 80300
rect 105320 80260 105636 80288
rect 105320 80248 105326 80260
rect 105630 80248 105636 80260
rect 105688 80248 105694 80300
rect 132218 80248 132224 80300
rect 132276 80288 132282 80300
rect 132276 80260 140774 80288
rect 132276 80248 132282 80260
rect 131114 80180 131120 80232
rect 131172 80220 131178 80232
rect 131172 80192 134150 80220
rect 131172 80180 131178 80192
rect 129090 79976 129096 80028
rect 129148 80016 129154 80028
rect 134122 80016 134150 80192
rect 140746 80084 140774 80260
rect 143506 80152 143534 80464
rect 144886 80220 144914 80532
rect 144886 80192 145466 80220
rect 143506 80124 145374 80152
rect 140746 80056 143994 80084
rect 129148 79988 133966 80016
rect 134122 79988 142890 80016
rect 129148 79976 129154 79988
rect 133938 79960 133966 79988
rect 123478 79908 123484 79960
rect 123536 79948 123542 79960
rect 132908 79948 132914 79960
rect 123536 79920 132914 79948
rect 123536 79908 123542 79920
rect 132908 79908 132914 79920
rect 132966 79908 132972 79960
rect 133552 79908 133558 79960
rect 133610 79908 133616 79960
rect 133644 79908 133650 79960
rect 133702 79908 133708 79960
rect 133736 79908 133742 79960
rect 133794 79908 133800 79960
rect 133920 79908 133926 79960
rect 133978 79908 133984 79960
rect 134288 79908 134294 79960
rect 134346 79908 134352 79960
rect 134380 79908 134386 79960
rect 134438 79908 134444 79960
rect 134564 79908 134570 79960
rect 134622 79908 134628 79960
rect 136312 79948 136318 79960
rect 134812 79920 136318 79948
rect 128170 79840 128176 79892
rect 128228 79880 128234 79892
rect 133276 79880 133282 79892
rect 128228 79852 133282 79880
rect 128228 79840 128234 79852
rect 133276 79840 133282 79852
rect 133334 79840 133340 79892
rect 131390 79772 131396 79824
rect 131448 79812 131454 79824
rect 133570 79812 133598 79908
rect 131448 79784 133598 79812
rect 131448 79772 131454 79784
rect 133662 79756 133690 79908
rect 133598 79704 133604 79756
rect 133656 79716 133690 79756
rect 133656 79704 133662 79716
rect 113634 79636 113640 79688
rect 113692 79676 113698 79688
rect 132494 79676 132500 79688
rect 113692 79648 132500 79676
rect 113692 79636 113698 79648
rect 132494 79636 132500 79648
rect 132552 79636 132558 79688
rect 133230 79636 133236 79688
rect 133288 79676 133294 79688
rect 133754 79676 133782 79908
rect 134012 79840 134018 79892
rect 134070 79840 134076 79892
rect 133288 79648 133782 79676
rect 133288 79636 133294 79648
rect 133874 79636 133880 79688
rect 133932 79676 133938 79688
rect 134030 79676 134058 79840
rect 133932 79648 134058 79676
rect 133932 79636 133938 79648
rect 134150 79636 134156 79688
rect 134208 79676 134214 79688
rect 134306 79676 134334 79908
rect 134398 79756 134426 79908
rect 134582 79824 134610 79908
rect 134656 79840 134662 79892
rect 134714 79840 134720 79892
rect 134518 79772 134524 79824
rect 134576 79784 134610 79824
rect 134576 79772 134582 79784
rect 134398 79716 134432 79756
rect 134426 79704 134432 79716
rect 134484 79704 134490 79756
rect 134208 79648 134334 79676
rect 134208 79636 134214 79648
rect 111334 79568 111340 79620
rect 111392 79608 111398 79620
rect 126330 79608 126336 79620
rect 111392 79580 126336 79608
rect 111392 79568 111398 79580
rect 126330 79568 126336 79580
rect 126388 79568 126394 79620
rect 133966 79568 133972 79620
rect 134024 79608 134030 79620
rect 134674 79608 134702 79840
rect 134812 79688 134840 79920
rect 136312 79908 136318 79920
rect 136370 79908 136376 79960
rect 137324 79948 137330 79960
rect 136744 79920 137330 79948
rect 134932 79840 134938 79892
rect 134990 79840 134996 79892
rect 135576 79840 135582 79892
rect 135634 79840 135640 79892
rect 136036 79840 136042 79892
rect 136094 79840 136100 79892
rect 136588 79840 136594 79892
rect 136646 79880 136652 79892
rect 136646 79840 136680 79880
rect 134950 79744 134978 79840
rect 135594 79812 135622 79840
rect 135548 79784 135622 79812
rect 134950 79716 135300 79744
rect 135272 79688 135300 79716
rect 134794 79636 134800 79688
rect 134852 79636 134858 79688
rect 135254 79636 135260 79688
rect 135312 79636 135318 79688
rect 135438 79636 135444 79688
rect 135496 79676 135502 79688
rect 135548 79676 135576 79784
rect 135668 79772 135674 79824
rect 135726 79812 135732 79824
rect 135726 79772 135760 79812
rect 135496 79648 135576 79676
rect 135496 79636 135502 79648
rect 134024 79580 134702 79608
rect 134024 79568 134030 79580
rect 135530 79568 135536 79620
rect 135588 79608 135594 79620
rect 135622 79608 135628 79620
rect 135588 79580 135628 79608
rect 135588 79568 135594 79580
rect 135622 79568 135628 79580
rect 135680 79568 135686 79620
rect 135732 79608 135760 79772
rect 136054 79744 136082 79840
rect 136054 79716 136312 79744
rect 136284 79688 136312 79716
rect 136652 79688 136680 79840
rect 136744 79688 136772 79920
rect 137324 79908 137330 79920
rect 137382 79908 137388 79960
rect 137968 79948 137974 79960
rect 137434 79920 137974 79948
rect 136864 79840 136870 79892
rect 136922 79840 136928 79892
rect 137048 79840 137054 79892
rect 137106 79840 137112 79892
rect 136882 79744 136910 79840
rect 136882 79716 136956 79744
rect 136928 79688 136956 79716
rect 137066 79688 137094 79840
rect 137434 79744 137462 79920
rect 137968 79908 137974 79920
rect 138026 79908 138032 79960
rect 138796 79948 138802 79960
rect 138354 79920 138802 79948
rect 137508 79840 137514 79892
rect 137566 79880 137572 79892
rect 137566 79840 137600 79880
rect 138244 79840 138250 79892
rect 138302 79840 138308 79892
rect 137434 79716 137508 79744
rect 137480 79688 137508 79716
rect 136266 79636 136272 79688
rect 136324 79636 136330 79688
rect 136634 79636 136640 79688
rect 136692 79636 136698 79688
rect 136726 79636 136732 79688
rect 136784 79636 136790 79688
rect 136910 79636 136916 79688
rect 136968 79636 136974 79688
rect 137066 79648 137100 79688
rect 137094 79636 137100 79648
rect 137152 79636 137158 79688
rect 137370 79636 137376 79688
rect 137428 79636 137434 79688
rect 137462 79636 137468 79688
rect 137520 79636 137526 79688
rect 136450 79608 136456 79620
rect 135732 79580 136456 79608
rect 119430 79500 119436 79552
rect 119488 79540 119494 79552
rect 127894 79540 127900 79552
rect 119488 79512 127900 79540
rect 119488 79500 119494 79512
rect 127894 79500 127900 79512
rect 127952 79500 127958 79552
rect 131942 79500 131948 79552
rect 132000 79540 132006 79552
rect 135732 79540 135760 79580
rect 136450 79568 136456 79580
rect 136508 79568 136514 79620
rect 137388 79608 137416 79636
rect 136560 79580 137416 79608
rect 132000 79512 135760 79540
rect 132000 79500 132006 79512
rect 117774 79432 117780 79484
rect 117832 79472 117838 79484
rect 127802 79472 127808 79484
rect 117832 79444 127808 79472
rect 117832 79432 117838 79444
rect 127802 79432 127808 79444
rect 127860 79432 127866 79484
rect 134334 79432 134340 79484
rect 134392 79472 134398 79484
rect 136560 79472 136588 79580
rect 134392 79444 136588 79472
rect 134392 79432 134398 79444
rect 136726 79432 136732 79484
rect 136784 79472 136790 79484
rect 137572 79472 137600 79840
rect 138262 79744 138290 79840
rect 137848 79716 138290 79744
rect 137848 79688 137876 79716
rect 137830 79636 137836 79688
rect 137888 79636 137894 79688
rect 138198 79636 138204 79688
rect 138256 79676 138262 79688
rect 138354 79676 138382 79920
rect 138796 79908 138802 79920
rect 138854 79908 138860 79960
rect 139348 79948 139354 79960
rect 138906 79920 139354 79948
rect 138428 79840 138434 79892
rect 138486 79880 138492 79892
rect 138486 79852 138796 79880
rect 138486 79840 138492 79852
rect 138768 79824 138796 79852
rect 138750 79772 138756 79824
rect 138808 79772 138814 79824
rect 138256 79648 138382 79676
rect 138256 79636 138262 79648
rect 138658 79636 138664 79688
rect 138716 79676 138722 79688
rect 138906 79676 138934 79920
rect 139348 79908 139354 79920
rect 139406 79908 139412 79960
rect 139440 79908 139446 79960
rect 139498 79948 139504 79960
rect 139498 79908 139532 79948
rect 139624 79908 139630 79960
rect 139682 79948 139688 79960
rect 139682 79908 139716 79948
rect 139900 79908 139906 79960
rect 139958 79948 139964 79960
rect 139958 79920 140498 79948
rect 139958 79908 139964 79920
rect 139072 79880 139078 79892
rect 138716 79648 138934 79676
rect 139044 79840 139078 79880
rect 139130 79840 139136 79892
rect 138716 79636 138722 79648
rect 139044 79620 139072 79840
rect 139164 79772 139170 79824
rect 139222 79772 139228 79824
rect 139026 79568 139032 79620
rect 139084 79568 139090 79620
rect 136784 79444 137600 79472
rect 136784 79432 136790 79444
rect 138934 79432 138940 79484
rect 138992 79472 138998 79484
rect 139182 79472 139210 79772
rect 139504 79688 139532 79908
rect 139688 79824 139716 79908
rect 139808 79840 139814 79892
rect 139866 79840 139872 79892
rect 140360 79880 140366 79892
rect 140010 79852 140366 79880
rect 139670 79772 139676 79824
rect 139728 79772 139734 79824
rect 139486 79636 139492 79688
rect 139544 79636 139550 79688
rect 139578 79636 139584 79688
rect 139636 79676 139642 79688
rect 139826 79676 139854 79840
rect 139636 79648 139854 79676
rect 139636 79636 139642 79648
rect 140010 79552 140038 79852
rect 140360 79840 140366 79852
rect 140418 79840 140424 79892
rect 140470 79812 140498 79920
rect 140544 79908 140550 79960
rect 140602 79948 140608 79960
rect 140602 79908 140636 79948
rect 140728 79908 140734 79960
rect 140786 79908 140792 79960
rect 140820 79908 140826 79960
rect 140878 79908 140884 79960
rect 141004 79908 141010 79960
rect 141062 79908 141068 79960
rect 141648 79908 141654 79960
rect 141706 79908 141712 79960
rect 141832 79908 141838 79960
rect 141890 79908 141896 79960
rect 141924 79908 141930 79960
rect 141982 79908 141988 79960
rect 142016 79908 142022 79960
rect 142074 79908 142080 79960
rect 142200 79908 142206 79960
rect 142258 79908 142264 79960
rect 140470 79784 140544 79812
rect 140406 79704 140412 79756
rect 140464 79704 140470 79756
rect 140222 79636 140228 79688
rect 140280 79676 140286 79688
rect 140424 79676 140452 79704
rect 140280 79648 140452 79676
rect 140280 79636 140286 79648
rect 139946 79500 139952 79552
rect 140004 79512 140038 79552
rect 140004 79500 140010 79512
rect 140406 79500 140412 79552
rect 140464 79540 140470 79552
rect 140516 79540 140544 79784
rect 140608 79688 140636 79908
rect 140590 79636 140596 79688
rect 140648 79636 140654 79688
rect 140464 79512 140544 79540
rect 140464 79500 140470 79512
rect 138992 79444 139210 79472
rect 138992 79432 138998 79444
rect 140498 79432 140504 79484
rect 140556 79472 140562 79484
rect 140746 79472 140774 79908
rect 140838 79688 140866 79908
rect 141022 79688 141050 79908
rect 141464 79880 141470 79892
rect 141160 79852 141470 79880
rect 141160 79688 141188 79852
rect 141464 79840 141470 79852
rect 141522 79840 141528 79892
rect 141666 79756 141694 79908
rect 141602 79704 141608 79756
rect 141660 79716 141694 79756
rect 141660 79704 141666 79716
rect 140838 79648 140872 79688
rect 140866 79636 140872 79648
rect 140924 79636 140930 79688
rect 140958 79636 140964 79688
rect 141016 79648 141050 79688
rect 141016 79636 141022 79648
rect 141142 79636 141148 79688
rect 141200 79636 141206 79688
rect 141694 79568 141700 79620
rect 141752 79568 141758 79620
rect 141326 79500 141332 79552
rect 141384 79540 141390 79552
rect 141712 79540 141740 79568
rect 141384 79512 141740 79540
rect 141850 79540 141878 79908
rect 141942 79744 141970 79908
rect 142034 79824 142062 79908
rect 142034 79784 142068 79824
rect 142062 79772 142068 79784
rect 142120 79772 142126 79824
rect 142218 79756 142246 79908
rect 141942 79716 142108 79744
rect 141970 79540 141976 79552
rect 141850 79512 141976 79540
rect 141384 79500 141390 79512
rect 141970 79500 141976 79512
rect 142028 79500 142034 79552
rect 142080 79540 142108 79716
rect 142154 79704 142160 79756
rect 142212 79716 142246 79756
rect 142212 79704 142218 79716
rect 142310 79688 142338 79988
rect 142862 79960 142890 79988
rect 143966 79960 143994 80056
rect 144242 79988 144960 80016
rect 144242 79960 144270 79988
rect 142384 79908 142390 79960
rect 142442 79908 142448 79960
rect 142476 79908 142482 79960
rect 142534 79908 142540 79960
rect 142568 79908 142574 79960
rect 142626 79908 142632 79960
rect 142844 79908 142850 79960
rect 142902 79908 142908 79960
rect 143948 79908 143954 79960
rect 144006 79908 144012 79960
rect 144040 79908 144046 79960
rect 144098 79948 144104 79960
rect 144098 79920 144178 79948
rect 144098 79908 144104 79920
rect 142402 79824 142430 79908
rect 142384 79772 142390 79824
rect 142442 79772 142448 79824
rect 142494 79744 142522 79908
rect 142586 79880 142614 79908
rect 142586 79852 142660 79880
rect 142494 79716 142568 79744
rect 142540 79688 142568 79716
rect 142246 79636 142252 79688
rect 142304 79648 142338 79688
rect 142304 79636 142310 79648
rect 142522 79636 142528 79688
rect 142580 79636 142586 79688
rect 142632 79552 142660 79852
rect 143028 79840 143034 79892
rect 143086 79840 143092 79892
rect 143396 79840 143402 79892
rect 143454 79840 143460 79892
rect 143046 79688 143074 79840
rect 143212 79772 143218 79824
rect 143270 79772 143276 79824
rect 143230 79688 143258 79772
rect 143046 79648 143080 79688
rect 143074 79636 143080 79648
rect 143132 79636 143138 79688
rect 143166 79636 143172 79688
rect 143224 79648 143258 79688
rect 143224 79636 143230 79648
rect 142338 79540 142344 79552
rect 142080 79512 142344 79540
rect 142338 79500 142344 79512
rect 142396 79500 142402 79552
rect 142614 79500 142620 79552
rect 142672 79500 142678 79552
rect 142706 79500 142712 79552
rect 142764 79540 142770 79552
rect 143414 79540 143442 79840
rect 143764 79772 143770 79824
rect 143822 79772 143828 79824
rect 143534 79568 143540 79620
rect 143592 79608 143598 79620
rect 143782 79608 143810 79772
rect 143592 79580 143810 79608
rect 143592 79568 143598 79580
rect 142764 79512 143442 79540
rect 142764 79500 142770 79512
rect 143810 79500 143816 79552
rect 143868 79540 143874 79552
rect 144150 79540 144178 79920
rect 144224 79908 144230 79960
rect 144282 79908 144288 79960
rect 144408 79840 144414 79892
rect 144466 79840 144472 79892
rect 144500 79840 144506 79892
rect 144558 79840 144564 79892
rect 144684 79840 144690 79892
rect 144742 79840 144748 79892
rect 144932 79880 144960 79988
rect 145346 79960 145374 80124
rect 145144 79948 145150 79960
rect 144794 79852 144960 79880
rect 145116 79908 145150 79948
rect 145202 79908 145208 79960
rect 145328 79908 145334 79960
rect 145386 79908 145392 79960
rect 145438 79948 145466 80192
rect 145530 80152 145558 80736
rect 145530 80124 146386 80152
rect 145944 79988 146294 80016
rect 145512 79948 145518 79960
rect 145438 79920 145518 79948
rect 144316 79772 144322 79824
rect 144374 79772 144380 79824
rect 144334 79744 144362 79772
rect 144288 79716 144362 79744
rect 144288 79688 144316 79716
rect 144426 79688 144454 79840
rect 144270 79636 144276 79688
rect 144328 79636 144334 79688
rect 144362 79636 144368 79688
rect 144420 79648 144454 79688
rect 144420 79636 144426 79648
rect 144518 79620 144546 79840
rect 144702 79756 144730 79840
rect 144638 79704 144644 79756
rect 144696 79716 144730 79756
rect 144696 79704 144702 79716
rect 144454 79568 144460 79620
rect 144512 79580 144546 79620
rect 144512 79568 144518 79580
rect 144794 79552 144822 79852
rect 144868 79772 144874 79824
rect 144926 79772 144932 79824
rect 144886 79620 144914 79772
rect 145116 79756 145144 79908
rect 145190 79772 145196 79824
rect 145248 79812 145254 79824
rect 145438 79812 145466 79920
rect 145512 79908 145518 79920
rect 145570 79908 145576 79960
rect 145696 79840 145702 79892
rect 145754 79840 145760 79892
rect 145248 79784 145466 79812
rect 145248 79772 145254 79784
rect 145098 79704 145104 79756
rect 145156 79704 145162 79756
rect 144886 79580 144920 79620
rect 144914 79568 144920 79580
rect 144972 79568 144978 79620
rect 143868 79512 144178 79540
rect 143868 79500 143874 79512
rect 144730 79500 144736 79552
rect 144788 79512 144822 79552
rect 144788 79500 144794 79512
rect 140556 79444 140774 79472
rect 140556 79432 140562 79444
rect 145466 79432 145472 79484
rect 145524 79472 145530 79484
rect 145714 79472 145742 79840
rect 145834 79636 145840 79688
rect 145892 79676 145898 79688
rect 145944 79676 145972 79988
rect 146266 79960 146294 79988
rect 146248 79908 146254 79960
rect 146306 79908 146312 79960
rect 146064 79840 146070 79892
rect 146122 79840 146128 79892
rect 146156 79840 146162 79892
rect 146214 79880 146220 79892
rect 146358 79880 146386 80124
rect 146214 79852 146386 79880
rect 146214 79840 146220 79852
rect 146432 79840 146438 79892
rect 146490 79840 146496 79892
rect 146616 79840 146622 79892
rect 146674 79840 146680 79892
rect 146082 79812 146110 79840
rect 146082 79784 146340 79812
rect 146312 79756 146340 79784
rect 146294 79704 146300 79756
rect 146352 79704 146358 79756
rect 145892 79648 145972 79676
rect 146450 79688 146478 79840
rect 146450 79648 146484 79688
rect 145892 79636 145898 79648
rect 146478 79636 146484 79648
rect 146536 79636 146542 79688
rect 146110 79568 146116 79620
rect 146168 79608 146174 79620
rect 146634 79608 146662 79840
rect 146168 79580 146662 79608
rect 146168 79568 146174 79580
rect 146386 79500 146392 79552
rect 146444 79540 146450 79552
rect 146726 79540 146754 80940
rect 157628 80872 164234 80900
rect 157628 80832 157656 80872
rect 153626 80804 157656 80832
rect 164206 80832 164234 80872
rect 176626 80832 176654 81008
rect 186148 80968 186176 81008
rect 164206 80804 176654 80832
rect 178696 80940 186176 80968
rect 193186 80968 193214 81008
rect 199470 80968 199476 80980
rect 193186 80940 199476 80968
rect 153626 80016 153654 80804
rect 164114 80736 178632 80764
rect 164114 80492 164142 80736
rect 155834 80464 164142 80492
rect 164206 80668 173894 80696
rect 155834 80016 155862 80464
rect 164206 80424 164234 80668
rect 173866 80628 173894 80668
rect 173866 80600 176654 80628
rect 172486 80532 174538 80560
rect 172486 80424 172514 80532
rect 147646 79988 147858 80016
rect 146800 79908 146806 79960
rect 146858 79908 146864 79960
rect 146818 79756 146846 79908
rect 146892 79840 146898 79892
rect 146950 79880 146956 79892
rect 147168 79880 147174 79892
rect 146950 79840 146984 79880
rect 146818 79716 146852 79756
rect 146846 79704 146852 79716
rect 146904 79704 146910 79756
rect 146846 79568 146852 79620
rect 146904 79608 146910 79620
rect 146956 79608 146984 79840
rect 147140 79840 147174 79880
rect 147226 79840 147232 79892
rect 147536 79880 147542 79892
rect 147278 79852 147542 79880
rect 147140 79756 147168 79840
rect 147278 79812 147306 79852
rect 147536 79840 147542 79852
rect 147594 79840 147600 79892
rect 147232 79784 147306 79812
rect 147232 79756 147260 79784
rect 147352 79772 147358 79824
rect 147410 79772 147416 79824
rect 147122 79704 147128 79756
rect 147180 79704 147186 79756
rect 147214 79704 147220 79756
rect 147272 79704 147278 79756
rect 147370 79688 147398 79772
rect 147306 79636 147312 79688
rect 147364 79648 147398 79688
rect 147364 79636 147370 79648
rect 147646 79608 147674 79988
rect 147830 79960 147858 79988
rect 150682 79988 153286 80016
rect 150682 79960 150710 79988
rect 147720 79908 147726 79960
rect 147778 79908 147784 79960
rect 147812 79908 147818 79960
rect 147870 79908 147876 79960
rect 147904 79908 147910 79960
rect 147962 79908 147968 79960
rect 148456 79908 148462 79960
rect 148514 79908 148520 79960
rect 149008 79908 149014 79960
rect 149066 79908 149072 79960
rect 149192 79908 149198 79960
rect 149250 79948 149256 79960
rect 149250 79920 149422 79948
rect 149250 79908 149256 79920
rect 147738 79756 147766 79908
rect 147738 79716 147772 79756
rect 147766 79704 147772 79716
rect 147824 79704 147830 79756
rect 147922 79744 147950 79908
rect 148272 79840 148278 79892
rect 148330 79840 148336 79892
rect 147996 79772 148002 79824
rect 148054 79772 148060 79824
rect 148088 79772 148094 79824
rect 148146 79772 148152 79824
rect 147876 79716 147950 79744
rect 146904 79580 146984 79608
rect 147600 79580 147674 79608
rect 146904 79568 146910 79580
rect 146444 79512 146754 79540
rect 146444 79500 146450 79512
rect 145524 79444 145742 79472
rect 147600 79472 147628 79580
rect 147674 79500 147680 79552
rect 147732 79540 147738 79552
rect 147876 79540 147904 79716
rect 148014 79688 148042 79772
rect 147950 79636 147956 79688
rect 148008 79648 148042 79688
rect 148106 79676 148134 79772
rect 148290 79676 148318 79840
rect 148474 79824 148502 79908
rect 148732 79840 148738 79892
rect 148790 79840 148796 79892
rect 148824 79840 148830 79892
rect 148882 79840 148888 79892
rect 148474 79784 148508 79824
rect 148502 79772 148508 79784
rect 148560 79772 148566 79824
rect 148594 79676 148600 79688
rect 148106 79648 148180 79676
rect 148290 79648 148600 79676
rect 148008 79636 148014 79648
rect 148152 79552 148180 79648
rect 148594 79636 148600 79648
rect 148652 79636 148658 79688
rect 148750 79608 148778 79840
rect 148244 79580 148778 79608
rect 148842 79608 148870 79840
rect 149026 79688 149054 79908
rect 149284 79840 149290 79892
rect 149342 79840 149348 79892
rect 148962 79636 148968 79688
rect 149020 79648 149054 79688
rect 149302 79688 149330 79840
rect 149394 79824 149422 79920
rect 149468 79908 149474 79960
rect 149526 79908 149532 79960
rect 149744 79908 149750 79960
rect 149802 79908 149808 79960
rect 149928 79908 149934 79960
rect 149986 79908 149992 79960
rect 150020 79908 150026 79960
rect 150078 79908 150084 79960
rect 150112 79908 150118 79960
rect 150170 79908 150176 79960
rect 150204 79908 150210 79960
rect 150262 79908 150268 79960
rect 150664 79908 150670 79960
rect 150722 79908 150728 79960
rect 150756 79908 150762 79960
rect 150814 79908 150820 79960
rect 151308 79908 151314 79960
rect 151366 79908 151372 79960
rect 151400 79908 151406 79960
rect 151458 79908 151464 79960
rect 152320 79948 152326 79960
rect 151740 79920 152326 79948
rect 149376 79772 149382 79824
rect 149434 79772 149440 79824
rect 149486 79688 149514 79908
rect 149302 79648 149336 79688
rect 149020 79636 149026 79648
rect 149330 79636 149336 79648
rect 149388 79636 149394 79688
rect 149422 79636 149428 79688
rect 149480 79648 149514 79688
rect 149480 79636 149486 79648
rect 149606 79636 149612 79688
rect 149664 79676 149670 79688
rect 149762 79676 149790 79908
rect 149946 79688 149974 79908
rect 149664 79648 149790 79676
rect 149664 79636 149670 79648
rect 149882 79636 149888 79688
rect 149940 79648 149974 79688
rect 149940 79636 149946 79648
rect 148842 79580 149008 79608
rect 147732 79512 147904 79540
rect 147732 79500 147738 79512
rect 148134 79500 148140 79552
rect 148192 79500 148198 79552
rect 147858 79472 147864 79484
rect 147600 79444 147864 79472
rect 145524 79432 145530 79444
rect 147858 79432 147864 79444
rect 147916 79432 147922 79484
rect 148042 79432 148048 79484
rect 148100 79472 148106 79484
rect 148244 79472 148272 79580
rect 148594 79500 148600 79552
rect 148652 79540 148658 79552
rect 148870 79540 148876 79552
rect 148652 79512 148876 79540
rect 148652 79500 148658 79512
rect 148870 79500 148876 79512
rect 148928 79500 148934 79552
rect 148980 79540 149008 79580
rect 149054 79568 149060 79620
rect 149112 79608 149118 79620
rect 150038 79608 150066 79908
rect 150130 79676 150158 79908
rect 150222 79744 150250 79908
rect 150774 79824 150802 79908
rect 151032 79840 151038 79892
rect 151090 79840 151096 79892
rect 150710 79772 150716 79824
rect 150768 79784 150802 79824
rect 150768 79772 150774 79784
rect 150940 79772 150946 79824
rect 150998 79772 151004 79824
rect 150222 79716 150388 79744
rect 150250 79676 150256 79688
rect 150130 79648 150256 79676
rect 150250 79636 150256 79648
rect 150308 79636 150314 79688
rect 149112 79580 150066 79608
rect 149112 79568 149118 79580
rect 150158 79568 150164 79620
rect 150216 79608 150222 79620
rect 150360 79608 150388 79716
rect 150958 79620 150986 79772
rect 151050 79688 151078 79840
rect 151124 79772 151130 79824
rect 151182 79772 151188 79824
rect 151142 79744 151170 79772
rect 151326 79756 151354 79908
rect 151418 79880 151446 79908
rect 151418 79852 151492 79880
rect 151142 79716 151216 79744
rect 151326 79716 151360 79756
rect 151050 79648 151084 79688
rect 151078 79636 151084 79648
rect 151136 79636 151142 79688
rect 151188 79620 151216 79716
rect 151354 79704 151360 79716
rect 151412 79704 151418 79756
rect 151464 79620 151492 79852
rect 150216 79580 150388 79608
rect 150216 79568 150222 79580
rect 150894 79568 150900 79620
rect 150952 79580 150986 79620
rect 150952 79568 150958 79580
rect 151170 79568 151176 79620
rect 151228 79568 151234 79620
rect 151446 79568 151452 79620
rect 151504 79568 151510 79620
rect 151740 79552 151768 79920
rect 152320 79908 152326 79920
rect 152378 79908 152384 79960
rect 152412 79908 152418 79960
rect 152470 79908 152476 79960
rect 153148 79908 153154 79960
rect 153206 79908 153212 79960
rect 151952 79840 151958 79892
rect 152010 79840 152016 79892
rect 152228 79840 152234 79892
rect 152286 79840 152292 79892
rect 150066 79540 150072 79552
rect 148980 79512 150072 79540
rect 150066 79500 150072 79512
rect 150124 79500 150130 79552
rect 151722 79500 151728 79552
rect 151780 79500 151786 79552
rect 151970 79540 151998 79840
rect 152246 79756 152274 79840
rect 152430 79824 152458 79908
rect 152964 79840 152970 79892
rect 153022 79840 153028 79892
rect 152366 79772 152372 79824
rect 152424 79784 152458 79824
rect 152424 79772 152430 79784
rect 152246 79716 152280 79756
rect 152274 79704 152280 79716
rect 152332 79704 152338 79756
rect 152982 79620 153010 79840
rect 152918 79568 152924 79620
rect 152976 79580 153010 79620
rect 152976 79568 152982 79580
rect 152826 79540 152832 79552
rect 151970 79512 152832 79540
rect 152826 79500 152832 79512
rect 152884 79500 152890 79552
rect 148100 79444 148272 79472
rect 148100 79432 148106 79444
rect 148410 79432 148416 79484
rect 148468 79472 148474 79484
rect 148778 79472 148784 79484
rect 148468 79444 148784 79472
rect 148468 79432 148474 79444
rect 148778 79432 148784 79444
rect 148836 79432 148842 79484
rect 151814 79432 151820 79484
rect 151872 79472 151878 79484
rect 153166 79472 153194 79908
rect 153258 79676 153286 79988
rect 153442 79988 153654 80016
rect 153994 79988 155862 80016
rect 155926 80396 164234 80424
rect 167150 80396 172514 80424
rect 153442 79960 153470 79988
rect 153424 79908 153430 79960
rect 153482 79908 153488 79960
rect 153516 79908 153522 79960
rect 153574 79908 153580 79960
rect 153700 79948 153706 79960
rect 153672 79908 153706 79948
rect 153758 79908 153764 79960
rect 153884 79948 153890 79960
rect 153856 79908 153890 79948
rect 153942 79908 153948 79960
rect 153534 79824 153562 79908
rect 153470 79772 153476 79824
rect 153528 79784 153562 79824
rect 153528 79772 153534 79784
rect 153672 79756 153700 79908
rect 153856 79824 153884 79908
rect 153838 79772 153844 79824
rect 153896 79772 153902 79824
rect 153654 79704 153660 79756
rect 153712 79704 153718 79756
rect 153994 79676 154022 79988
rect 155926 79960 155954 80396
rect 167150 80288 167178 80396
rect 174510 80356 174538 80532
rect 176626 80492 176654 80600
rect 178604 80560 178632 80736
rect 178696 80640 178724 80940
rect 199470 80928 199476 80940
rect 199528 80928 199534 80980
rect 198182 80900 198188 80912
rect 178788 80872 183554 80900
rect 178788 80640 178816 80872
rect 183526 80832 183554 80872
rect 186424 80872 198188 80900
rect 186424 80832 186452 80872
rect 198182 80860 198188 80872
rect 198240 80860 198246 80912
rect 183526 80804 186452 80832
rect 188430 80792 188436 80844
rect 188488 80832 188494 80844
rect 215662 80832 215668 80844
rect 188488 80804 215668 80832
rect 188488 80792 188494 80804
rect 215662 80792 215668 80804
rect 215720 80832 215726 80844
rect 270494 80832 270500 80844
rect 215720 80804 270500 80832
rect 215720 80792 215726 80804
rect 270494 80792 270500 80804
rect 270552 80792 270558 80844
rect 215846 80764 215852 80776
rect 186286 80736 215852 80764
rect 186286 80696 186314 80736
rect 215846 80724 215852 80736
rect 215904 80764 215910 80776
rect 234614 80764 234620 80776
rect 215904 80736 234620 80764
rect 215904 80724 215910 80736
rect 234614 80724 234620 80736
rect 234672 80724 234678 80776
rect 302234 80696 302240 80708
rect 183526 80668 186314 80696
rect 190426 80668 302240 80696
rect 178678 80588 178684 80640
rect 178736 80588 178742 80640
rect 178770 80588 178776 80640
rect 178828 80588 178834 80640
rect 183526 80560 183554 80668
rect 189902 80560 189908 80572
rect 178604 80532 183554 80560
rect 186286 80532 189908 80560
rect 186286 80492 186314 80532
rect 189902 80520 189908 80532
rect 189960 80560 189966 80572
rect 190426 80560 190454 80668
rect 302234 80656 302240 80668
rect 302292 80656 302298 80708
rect 189960 80532 190454 80560
rect 189960 80520 189966 80532
rect 176626 80464 186314 80492
rect 157030 80260 167178 80288
rect 167242 80328 173894 80356
rect 174510 80328 182174 80356
rect 156386 79988 156874 80016
rect 154436 79908 154442 79960
rect 154494 79908 154500 79960
rect 154804 79908 154810 79960
rect 154862 79948 154868 79960
rect 154862 79908 154896 79948
rect 154988 79908 154994 79960
rect 155046 79908 155052 79960
rect 155356 79908 155362 79960
rect 155414 79908 155420 79960
rect 155540 79908 155546 79960
rect 155598 79908 155604 79960
rect 155908 79908 155914 79960
rect 155966 79908 155972 79960
rect 156184 79908 156190 79960
rect 156242 79908 156248 79960
rect 156276 79908 156282 79960
rect 156334 79908 156340 79960
rect 154068 79840 154074 79892
rect 154126 79880 154132 79892
rect 154126 79840 154160 79880
rect 154132 79756 154160 79840
rect 154114 79704 154120 79756
rect 154172 79704 154178 79756
rect 153258 79648 154022 79676
rect 153746 79500 153752 79552
rect 153804 79540 153810 79552
rect 154454 79540 154482 79908
rect 154868 79756 154896 79908
rect 154850 79704 154856 79756
rect 154908 79704 154914 79756
rect 155006 79688 155034 79908
rect 155374 79824 155402 79908
rect 155310 79772 155316 79824
rect 155368 79784 155402 79824
rect 155558 79824 155586 79908
rect 155724 79840 155730 79892
rect 155782 79840 155788 79892
rect 155816 79840 155822 79892
rect 155874 79840 155880 79892
rect 155558 79784 155592 79824
rect 155368 79772 155374 79784
rect 155586 79772 155592 79784
rect 155644 79772 155650 79824
rect 155006 79648 155040 79688
rect 155034 79636 155040 79648
rect 155092 79636 155098 79688
rect 155402 79568 155408 79620
rect 155460 79608 155466 79620
rect 155742 79608 155770 79840
rect 155460 79580 155770 79608
rect 155834 79620 155862 79840
rect 156202 79756 156230 79908
rect 156294 79824 156322 79908
rect 156276 79772 156282 79824
rect 156334 79772 156340 79824
rect 156138 79704 156144 79756
rect 156196 79716 156230 79756
rect 156196 79704 156202 79716
rect 155834 79580 155868 79620
rect 155460 79568 155466 79580
rect 155862 79568 155868 79580
rect 155920 79568 155926 79620
rect 156386 79552 156414 79988
rect 156846 79892 156874 79988
rect 156920 79908 156926 79960
rect 156978 79908 156984 79960
rect 156644 79840 156650 79892
rect 156702 79840 156708 79892
rect 156828 79840 156834 79892
rect 156886 79840 156892 79892
rect 153804 79512 154482 79540
rect 153804 79500 153810 79512
rect 156322 79500 156328 79552
rect 156380 79512 156414 79552
rect 156662 79552 156690 79840
rect 156938 79756 156966 79908
rect 156782 79704 156788 79756
rect 156840 79704 156846 79756
rect 156874 79704 156880 79756
rect 156932 79716 156966 79756
rect 156932 79704 156938 79716
rect 156800 79620 156828 79704
rect 157030 79688 157058 80260
rect 167242 80220 167270 80328
rect 160342 80192 167270 80220
rect 168668 80260 169754 80288
rect 158640 79988 158990 80016
rect 157104 79908 157110 79960
rect 157162 79908 157168 79960
rect 157380 79908 157386 79960
rect 157438 79908 157444 79960
rect 157748 79908 157754 79960
rect 157806 79908 157812 79960
rect 157840 79908 157846 79960
rect 157898 79908 157904 79960
rect 157932 79908 157938 79960
rect 157990 79908 157996 79960
rect 158208 79908 158214 79960
rect 158266 79948 158272 79960
rect 158392 79948 158398 79960
rect 158266 79908 158300 79948
rect 156966 79636 156972 79688
rect 157024 79648 157058 79688
rect 157122 79688 157150 79908
rect 157398 79756 157426 79908
rect 157656 79880 157662 79892
rect 157628 79840 157662 79880
rect 157714 79840 157720 79892
rect 157472 79772 157478 79824
rect 157530 79812 157536 79824
rect 157530 79772 157564 79812
rect 157334 79704 157340 79756
rect 157392 79716 157426 79756
rect 157392 79704 157398 79716
rect 157122 79648 157156 79688
rect 157024 79636 157030 79648
rect 157150 79636 157156 79648
rect 157208 79636 157214 79688
rect 157536 79620 157564 79772
rect 157628 79620 157656 79840
rect 157766 79756 157794 79908
rect 157702 79704 157708 79756
rect 157760 79716 157794 79756
rect 157760 79704 157766 79716
rect 157858 79620 157886 79908
rect 156782 79568 156788 79620
rect 156840 79568 156846 79620
rect 157518 79568 157524 79620
rect 157576 79568 157582 79620
rect 157610 79568 157616 79620
rect 157668 79568 157674 79620
rect 157794 79568 157800 79620
rect 157852 79580 157886 79620
rect 157950 79620 157978 79908
rect 158272 79756 158300 79908
rect 158364 79908 158398 79948
rect 158450 79908 158456 79960
rect 158484 79908 158490 79960
rect 158542 79908 158548 79960
rect 158254 79704 158260 79756
rect 158312 79704 158318 79756
rect 158364 79688 158392 79908
rect 158502 79824 158530 79908
rect 158438 79772 158444 79824
rect 158496 79784 158530 79824
rect 158496 79772 158502 79784
rect 158346 79636 158352 79688
rect 158404 79636 158410 79688
rect 157950 79580 157984 79620
rect 157852 79568 157858 79580
rect 157978 79568 157984 79580
rect 158036 79568 158042 79620
rect 156662 79512 156696 79552
rect 156380 79500 156386 79512
rect 156690 79500 156696 79512
rect 156748 79500 156754 79552
rect 151872 79444 153194 79472
rect 158640 79472 158668 79988
rect 158962 79960 158990 79988
rect 160342 79960 160370 80192
rect 168668 80016 168696 80260
rect 169726 80084 169754 80260
rect 173866 80152 173894 80328
rect 177758 80152 177764 80164
rect 173866 80124 177764 80152
rect 177758 80112 177764 80124
rect 177816 80112 177822 80164
rect 182146 80152 182174 80328
rect 238754 80152 238760 80164
rect 182146 80124 238760 80152
rect 238754 80112 238760 80124
rect 238812 80112 238818 80164
rect 179230 80084 179236 80096
rect 169726 80056 179236 80084
rect 179230 80044 179236 80056
rect 179288 80044 179294 80096
rect 184474 80044 184480 80096
rect 184532 80084 184538 80096
rect 187234 80084 187240 80096
rect 184532 80056 187240 80084
rect 184532 80044 184538 80056
rect 187234 80044 187240 80056
rect 187292 80044 187298 80096
rect 211982 80044 211988 80096
rect 212040 80084 212046 80096
rect 212350 80084 212356 80096
rect 212040 80056 212356 80084
rect 212040 80044 212046 80056
rect 212350 80044 212356 80056
rect 212408 80084 212414 80096
rect 523126 80084 523132 80096
rect 212408 80056 523132 80084
rect 212408 80044 212414 80056
rect 523126 80044 523132 80056
rect 523184 80044 523190 80096
rect 180518 80016 180524 80028
rect 167334 79988 168696 80016
rect 172762 79988 173894 80016
rect 158760 79908 158766 79960
rect 158818 79908 158824 79960
rect 158944 79908 158950 79960
rect 159002 79908 159008 79960
rect 159220 79908 159226 79960
rect 159278 79908 159284 79960
rect 159956 79908 159962 79960
rect 160014 79908 160020 79960
rect 160048 79908 160054 79960
rect 160106 79908 160112 79960
rect 160140 79908 160146 79960
rect 160198 79908 160204 79960
rect 160324 79908 160330 79960
rect 160382 79908 160388 79960
rect 160692 79948 160698 79960
rect 160434 79920 160698 79948
rect 158778 79540 158806 79908
rect 158852 79840 158858 79892
rect 158910 79840 158916 79892
rect 158870 79756 158898 79840
rect 159238 79812 159266 79908
rect 159588 79880 159594 79892
rect 159192 79784 159266 79812
rect 159422 79852 159594 79880
rect 158870 79716 158904 79756
rect 158898 79704 158904 79716
rect 158956 79704 158962 79756
rect 159192 79620 159220 79784
rect 159422 79744 159450 79852
rect 159588 79840 159594 79852
rect 159646 79840 159652 79892
rect 159772 79840 159778 79892
rect 159830 79880 159836 79892
rect 159830 79840 159864 79880
rect 159496 79772 159502 79824
rect 159554 79772 159560 79824
rect 159330 79716 159450 79744
rect 159174 79568 159180 79620
rect 159232 79568 159238 79620
rect 159330 79608 159358 79716
rect 159514 79688 159542 79772
rect 159514 79648 159548 79688
rect 159542 79636 159548 79648
rect 159600 79636 159606 79688
rect 159450 79608 159456 79620
rect 159330 79580 159456 79608
rect 159450 79568 159456 79580
rect 159508 79568 159514 79620
rect 159836 79552 159864 79840
rect 159974 79744 160002 79908
rect 160066 79824 160094 79908
rect 160048 79772 160054 79824
rect 160106 79772 160112 79824
rect 159928 79716 160002 79744
rect 159358 79540 159364 79552
rect 158778 79512 159364 79540
rect 159358 79500 159364 79512
rect 159416 79500 159422 79552
rect 159818 79500 159824 79552
rect 159876 79500 159882 79552
rect 159928 79540 159956 79716
rect 160158 79688 160186 79908
rect 160158 79648 160192 79688
rect 160186 79636 160192 79648
rect 160244 79636 160250 79688
rect 160002 79568 160008 79620
rect 160060 79608 160066 79620
rect 160434 79608 160462 79920
rect 160692 79908 160698 79920
rect 160750 79908 160756 79960
rect 161152 79908 161158 79960
rect 161210 79908 161216 79960
rect 161612 79908 161618 79960
rect 161670 79908 161676 79960
rect 162164 79908 162170 79960
rect 162222 79908 162228 79960
rect 163084 79948 163090 79960
rect 162826 79920 163090 79948
rect 160508 79772 160514 79824
rect 160566 79772 160572 79824
rect 160526 79688 160554 79772
rect 160526 79648 160560 79688
rect 160554 79636 160560 79648
rect 160612 79636 160618 79688
rect 160060 79580 160462 79608
rect 160060 79568 160066 79580
rect 160830 79540 160836 79552
rect 159928 79512 160836 79540
rect 160830 79500 160836 79512
rect 160888 79500 160894 79552
rect 160922 79500 160928 79552
rect 160980 79540 160986 79552
rect 161170 79540 161198 79908
rect 160980 79512 161198 79540
rect 161630 79552 161658 79908
rect 161704 79840 161710 79892
rect 161762 79840 161768 79892
rect 161888 79840 161894 79892
rect 161946 79840 161952 79892
rect 162182 79880 162210 79908
rect 162182 79852 162624 79880
rect 161722 79608 161750 79840
rect 161906 79608 161934 79840
rect 162256 79772 162262 79824
rect 162314 79812 162320 79824
rect 162314 79784 162532 79812
rect 162314 79772 162320 79784
rect 162504 79688 162532 79784
rect 162596 79688 162624 79852
rect 162716 79772 162722 79824
rect 162774 79772 162780 79824
rect 162734 79688 162762 79772
rect 162486 79636 162492 79688
rect 162544 79636 162550 79688
rect 162578 79636 162584 79688
rect 162636 79636 162642 79688
rect 162670 79636 162676 79688
rect 162728 79648 162762 79688
rect 162728 79636 162734 79648
rect 162826 79620 162854 79920
rect 163084 79908 163090 79920
rect 163142 79908 163148 79960
rect 163360 79908 163366 79960
rect 163418 79948 163424 79960
rect 163418 79920 163498 79948
rect 163418 79908 163424 79920
rect 162900 79840 162906 79892
rect 162958 79880 162964 79892
rect 162958 79852 163360 79880
rect 162958 79840 162964 79852
rect 163332 79824 163360 79852
rect 163470 79824 163498 79920
rect 163544 79908 163550 79960
rect 163602 79908 163608 79960
rect 164740 79948 164746 79960
rect 164620 79920 164746 79948
rect 163314 79772 163320 79824
rect 163372 79772 163378 79824
rect 163406 79772 163412 79824
rect 163464 79784 163498 79824
rect 163464 79772 163470 79784
rect 163562 79688 163590 79908
rect 163820 79840 163826 79892
rect 163878 79840 163884 79892
rect 164096 79840 164102 79892
rect 164154 79840 164160 79892
rect 163562 79648 163596 79688
rect 163590 79636 163596 79648
rect 163648 79636 163654 79688
rect 162026 79608 162032 79620
rect 161722 79580 161796 79608
rect 161906 79580 162032 79608
rect 161768 79552 161796 79580
rect 162026 79568 162032 79580
rect 162084 79568 162090 79620
rect 162762 79568 162768 79620
rect 162820 79580 162854 79620
rect 162820 79568 162826 79580
rect 163130 79568 163136 79620
rect 163188 79608 163194 79620
rect 163188 79580 163268 79608
rect 163188 79568 163194 79580
rect 163240 79552 163268 79580
rect 163838 79552 163866 79840
rect 164114 79552 164142 79840
rect 164280 79772 164286 79824
rect 164338 79772 164344 79824
rect 164298 79688 164326 79772
rect 164234 79636 164240 79688
rect 164292 79648 164326 79688
rect 164292 79636 164298 79648
rect 164620 79620 164648 79920
rect 164740 79908 164746 79920
rect 164798 79908 164804 79960
rect 164832 79908 164838 79960
rect 164890 79948 164896 79960
rect 164890 79920 165568 79948
rect 164890 79908 164896 79920
rect 164924 79840 164930 79892
rect 164982 79840 164988 79892
rect 165384 79840 165390 79892
rect 165442 79840 165448 79892
rect 164602 79568 164608 79620
rect 164660 79568 164666 79620
rect 161630 79512 161664 79552
rect 160980 79500 160986 79512
rect 161658 79500 161664 79512
rect 161716 79500 161722 79552
rect 161750 79500 161756 79552
rect 161808 79500 161814 79552
rect 162688 79512 162854 79540
rect 158714 79472 158720 79484
rect 158640 79444 158720 79472
rect 151872 79432 151878 79444
rect 158714 79432 158720 79444
rect 158772 79432 158778 79484
rect 162688 79472 162716 79512
rect 160066 79444 162716 79472
rect 162826 79472 162854 79512
rect 163222 79500 163228 79552
rect 163280 79500 163286 79552
rect 163774 79500 163780 79552
rect 163832 79512 163866 79552
rect 163832 79500 163838 79512
rect 164050 79500 164056 79552
rect 164108 79512 164142 79552
rect 164108 79500 164114 79512
rect 164694 79500 164700 79552
rect 164752 79540 164758 79552
rect 164942 79540 164970 79840
rect 165200 79772 165206 79824
rect 165258 79772 165264 79824
rect 165218 79744 165246 79772
rect 165172 79716 165246 79744
rect 165172 79688 165200 79716
rect 165154 79636 165160 79688
rect 165212 79636 165218 79688
rect 165246 79636 165252 79688
rect 165304 79676 165310 79688
rect 165402 79676 165430 79840
rect 165304 79648 165430 79676
rect 165304 79636 165310 79648
rect 165540 79620 165568 79920
rect 166672 79908 166678 79960
rect 166730 79908 166736 79960
rect 166764 79908 166770 79960
rect 166822 79908 166828 79960
rect 165660 79880 165666 79892
rect 165632 79840 165666 79880
rect 165718 79840 165724 79892
rect 166028 79840 166034 79892
rect 166086 79840 166092 79892
rect 166212 79840 166218 79892
rect 166270 79840 166276 79892
rect 165522 79568 165528 79620
rect 165580 79568 165586 79620
rect 165632 79552 165660 79840
rect 165890 79568 165896 79620
rect 165948 79608 165954 79620
rect 166046 79608 166074 79840
rect 166230 79620 166258 79840
rect 166690 79824 166718 79908
rect 166580 79772 166586 79824
rect 166638 79772 166644 79824
rect 166672 79772 166678 79824
rect 166730 79772 166736 79824
rect 166782 79812 166810 79908
rect 166856 79840 166862 79892
rect 166914 79880 166920 79892
rect 167334 79880 167362 79988
rect 167776 79908 167782 79960
rect 167834 79908 167840 79960
rect 167868 79908 167874 79960
rect 167926 79908 167932 79960
rect 167960 79908 167966 79960
rect 168018 79948 168024 79960
rect 168018 79908 168052 79948
rect 168328 79908 168334 79960
rect 168386 79908 168392 79960
rect 168512 79908 168518 79960
rect 168570 79948 168576 79960
rect 168972 79948 168978 79960
rect 168570 79908 168604 79948
rect 166914 79852 167362 79880
rect 166914 79840 166920 79852
rect 167408 79840 167414 79892
rect 167466 79840 167472 79892
rect 167592 79840 167598 79892
rect 167650 79840 167656 79892
rect 166948 79812 166954 79824
rect 166782 79784 166856 79812
rect 166598 79676 166626 79772
rect 166828 79688 166856 79784
rect 166920 79772 166954 79812
rect 167006 79772 167012 79824
rect 167316 79772 167322 79824
rect 167374 79772 167380 79824
rect 166718 79676 166724 79688
rect 166598 79648 166724 79676
rect 166718 79636 166724 79648
rect 166776 79636 166782 79688
rect 166810 79636 166816 79688
rect 166868 79636 166874 79688
rect 166920 79620 166948 79772
rect 167334 79688 167362 79772
rect 167270 79636 167276 79688
rect 167328 79648 167362 79688
rect 167426 79688 167454 79840
rect 167426 79648 167460 79688
rect 167328 79636 167334 79648
rect 167454 79636 167460 79648
rect 167512 79636 167518 79688
rect 165948 79580 166074 79608
rect 165948 79568 165954 79580
rect 166166 79568 166172 79620
rect 166224 79580 166258 79620
rect 166224 79568 166230 79580
rect 166902 79568 166908 79620
rect 166960 79568 166966 79620
rect 164752 79512 164970 79540
rect 164752 79500 164758 79512
rect 165614 79500 165620 79552
rect 165672 79500 165678 79552
rect 167362 79500 167368 79552
rect 167420 79540 167426 79552
rect 167610 79540 167638 79840
rect 167794 79744 167822 79908
rect 167420 79512 167638 79540
rect 167748 79716 167822 79744
rect 167420 79500 167426 79512
rect 167454 79472 167460 79484
rect 162826 79444 167460 79472
rect 108206 79364 108212 79416
rect 108264 79404 108270 79416
rect 121914 79404 121920 79416
rect 108264 79376 121920 79404
rect 108264 79364 108270 79376
rect 121914 79364 121920 79376
rect 121972 79364 121978 79416
rect 135622 79364 135628 79416
rect 135680 79404 135686 79416
rect 144546 79404 144552 79416
rect 135680 79376 144552 79404
rect 135680 79364 135686 79376
rect 144546 79364 144552 79376
rect 144604 79404 144610 79416
rect 145282 79404 145288 79416
rect 144604 79376 145288 79404
rect 144604 79364 144610 79376
rect 145282 79364 145288 79376
rect 145340 79364 145346 79416
rect 146294 79404 146300 79416
rect 146266 79364 146300 79404
rect 146352 79404 146358 79416
rect 160066 79404 160094 79444
rect 167454 79432 167460 79444
rect 167512 79432 167518 79484
rect 146352 79376 160094 79404
rect 146352 79364 146358 79376
rect 162854 79364 162860 79416
rect 162912 79404 162918 79416
rect 167748 79404 167776 79716
rect 167886 79552 167914 79908
rect 168024 79552 168052 79908
rect 168190 79568 168196 79620
rect 168248 79608 168254 79620
rect 168346 79608 168374 79908
rect 168420 79840 168426 79892
rect 168478 79880 168484 79892
rect 168478 79840 168512 79880
rect 168484 79688 168512 79840
rect 168576 79688 168604 79908
rect 168944 79908 168978 79948
rect 169030 79908 169036 79960
rect 169248 79908 169254 79960
rect 169306 79908 169312 79960
rect 169524 79908 169530 79960
rect 169582 79908 169588 79960
rect 169892 79908 169898 79960
rect 169950 79908 169956 79960
rect 170076 79948 170082 79960
rect 170048 79908 170082 79948
rect 170134 79908 170140 79960
rect 170168 79908 170174 79960
rect 170226 79908 170232 79960
rect 170996 79908 171002 79960
rect 171054 79908 171060 79960
rect 171456 79908 171462 79960
rect 171514 79908 171520 79960
rect 171548 79908 171554 79960
rect 171606 79908 171612 79960
rect 172468 79908 172474 79960
rect 172526 79908 172532 79960
rect 172560 79908 172566 79960
rect 172618 79908 172624 79960
rect 168696 79880 168702 79892
rect 168668 79840 168702 79880
rect 168754 79840 168760 79892
rect 168788 79840 168794 79892
rect 168846 79840 168852 79892
rect 168466 79636 168472 79688
rect 168524 79636 168530 79688
rect 168558 79636 168564 79688
rect 168616 79636 168622 79688
rect 168248 79580 168374 79608
rect 168248 79568 168254 79580
rect 167886 79512 167920 79552
rect 167914 79500 167920 79512
rect 167972 79500 167978 79552
rect 168006 79500 168012 79552
rect 168064 79500 168070 79552
rect 168558 79500 168564 79552
rect 168616 79540 168622 79552
rect 168668 79540 168696 79840
rect 168806 79812 168834 79840
rect 168616 79512 168696 79540
rect 168760 79784 168834 79812
rect 168760 79540 168788 79784
rect 168834 79704 168840 79756
rect 168892 79744 168898 79756
rect 168944 79744 168972 79908
rect 169064 79880 169070 79892
rect 168892 79716 168972 79744
rect 169036 79840 169070 79880
rect 169122 79840 169128 79892
rect 169156 79840 169162 79892
rect 169214 79840 169220 79892
rect 168892 79704 168898 79716
rect 169036 79620 169064 79840
rect 169174 79812 169202 79840
rect 169128 79784 169202 79812
rect 169128 79620 169156 79784
rect 169266 79756 169294 79908
rect 169202 79704 169208 79756
rect 169260 79716 169294 79756
rect 169260 79704 169266 79716
rect 169542 79688 169570 79908
rect 169910 79880 169938 79908
rect 169478 79636 169484 79688
rect 169536 79648 169570 79688
rect 169726 79852 169938 79880
rect 169536 79636 169542 79648
rect 169018 79568 169024 79620
rect 169076 79568 169082 79620
rect 169110 79568 169116 79620
rect 169168 79568 169174 79620
rect 169726 79608 169754 79852
rect 170048 79824 170076 79908
rect 170186 79880 170214 79908
rect 170140 79852 170214 79880
rect 169800 79772 169806 79824
rect 169858 79772 169864 79824
rect 170030 79772 170036 79824
rect 170088 79772 170094 79824
rect 169818 79744 169846 79772
rect 170140 79756 170168 79852
rect 170628 79840 170634 79892
rect 170686 79840 170692 79892
rect 170444 79772 170450 79824
rect 170502 79772 170508 79824
rect 169818 79716 170030 79744
rect 170002 79620 170030 79716
rect 170122 79704 170128 79756
rect 170180 79704 170186 79756
rect 169846 79608 169852 79620
rect 169726 79580 169852 79608
rect 169846 79568 169852 79580
rect 169904 79568 169910 79620
rect 169938 79568 169944 79620
rect 169996 79580 170030 79620
rect 170462 79620 170490 79772
rect 170462 79580 170496 79620
rect 169996 79568 170002 79580
rect 170490 79568 170496 79580
rect 170548 79568 170554 79620
rect 170646 79608 170674 79840
rect 171014 79812 171042 79908
rect 171088 79840 171094 79892
rect 171146 79840 171152 79892
rect 171474 79880 171502 79908
rect 171290 79852 171502 79880
rect 170922 79784 171042 79812
rect 170922 79688 170950 79784
rect 170922 79648 170956 79688
rect 170950 79636 170956 79648
rect 171008 79636 171014 79688
rect 170646 79580 170720 79608
rect 170692 79552 170720 79580
rect 169294 79540 169300 79552
rect 168760 79512 169300 79540
rect 168616 79500 168622 79512
rect 169294 79500 169300 79512
rect 169352 79500 169358 79552
rect 170674 79500 170680 79552
rect 170732 79500 170738 79552
rect 170950 79500 170956 79552
rect 171008 79540 171014 79552
rect 171106 79540 171134 79840
rect 171008 79512 171134 79540
rect 171290 79552 171318 79852
rect 171364 79772 171370 79824
rect 171422 79812 171428 79824
rect 171422 79772 171456 79812
rect 171428 79552 171456 79772
rect 171566 79744 171594 79908
rect 172486 79824 172514 79908
rect 172008 79812 172014 79824
rect 171520 79716 171594 79744
rect 171980 79772 172014 79812
rect 172066 79772 172072 79824
rect 172468 79772 172474 79824
rect 172526 79772 172532 79824
rect 171520 79552 171548 79716
rect 171980 79688 172008 79772
rect 171962 79636 171968 79688
rect 172020 79636 172026 79688
rect 172578 79620 172606 79908
rect 172578 79580 172612 79620
rect 172606 79568 172612 79580
rect 172664 79568 172670 79620
rect 172762 79608 172790 79988
rect 173866 79960 173894 79988
rect 174510 79988 180524 80016
rect 174510 79960 174538 79988
rect 180518 79976 180524 79988
rect 180576 79976 180582 80028
rect 172836 79908 172842 79960
rect 172894 79948 172900 79960
rect 172894 79920 173480 79948
rect 172894 79908 172900 79920
rect 173296 79840 173302 79892
rect 173354 79840 173360 79892
rect 173452 79880 173480 79920
rect 173848 79908 173854 79960
rect 173906 79908 173912 79960
rect 174216 79908 174222 79960
rect 174274 79948 174280 79960
rect 174274 79920 174400 79948
rect 174274 79908 174280 79920
rect 173452 79852 173526 79880
rect 173314 79812 173342 79840
rect 173268 79784 173342 79812
rect 172974 79608 172980 79620
rect 172762 79580 172980 79608
rect 172974 79568 172980 79580
rect 173032 79568 173038 79620
rect 173158 79568 173164 79620
rect 173216 79608 173222 79620
rect 173268 79608 173296 79784
rect 173388 79772 173394 79824
rect 173446 79772 173452 79824
rect 173406 79744 173434 79772
rect 173360 79716 173434 79744
rect 173360 79688 173388 79716
rect 173498 79688 173526 79852
rect 173940 79772 173946 79824
rect 173998 79772 174004 79824
rect 174032 79772 174038 79824
rect 174090 79772 174096 79824
rect 174124 79772 174130 79824
rect 174182 79812 174188 79824
rect 174182 79784 174308 79812
rect 174182 79772 174188 79784
rect 173342 79636 173348 79688
rect 173400 79636 173406 79688
rect 173434 79636 173440 79688
rect 173492 79648 173526 79688
rect 173492 79636 173498 79648
rect 173216 79580 173296 79608
rect 173216 79568 173222 79580
rect 173618 79568 173624 79620
rect 173676 79608 173682 79620
rect 173958 79608 173986 79772
rect 173676 79580 173986 79608
rect 174050 79620 174078 79772
rect 174050 79580 174084 79620
rect 173676 79568 173682 79580
rect 174078 79568 174084 79580
rect 174136 79568 174142 79620
rect 174280 79608 174308 79784
rect 174372 79688 174400 79920
rect 174492 79908 174498 79960
rect 174550 79908 174556 79960
rect 174584 79908 174590 79960
rect 174642 79908 174648 79960
rect 174786 79920 175044 79948
rect 174602 79756 174630 79908
rect 174786 79892 174814 79920
rect 174768 79840 174774 79892
rect 174826 79840 174832 79892
rect 174860 79840 174866 79892
rect 174918 79880 174924 79892
rect 174918 79840 174952 79880
rect 174924 79756 174952 79840
rect 174538 79704 174544 79756
rect 174596 79716 174630 79756
rect 174596 79704 174602 79716
rect 174906 79704 174912 79756
rect 174964 79704 174970 79756
rect 174354 79636 174360 79688
rect 174412 79636 174418 79688
rect 175016 79620 175044 79920
rect 175136 79908 175142 79960
rect 175194 79908 175200 79960
rect 175228 79908 175234 79960
rect 175286 79908 175292 79960
rect 175596 79908 175602 79960
rect 175654 79948 175660 79960
rect 175654 79920 175826 79948
rect 175654 79908 175660 79920
rect 175154 79756 175182 79908
rect 175246 79812 175274 79908
rect 175412 79840 175418 79892
rect 175470 79840 175476 79892
rect 175504 79840 175510 79892
rect 175562 79880 175568 79892
rect 175562 79840 175596 79880
rect 175246 79784 175320 79812
rect 175292 79756 175320 79784
rect 175430 79756 175458 79840
rect 175154 79716 175188 79756
rect 175182 79704 175188 79716
rect 175240 79704 175246 79756
rect 175274 79704 175280 79756
rect 175332 79704 175338 79756
rect 175430 79716 175464 79756
rect 175458 79704 175464 79716
rect 175516 79704 175522 79756
rect 175568 79620 175596 79840
rect 175688 79812 175694 79824
rect 175660 79772 175694 79812
rect 175746 79772 175752 79824
rect 175660 79620 175688 79772
rect 175798 79688 175826 79920
rect 175964 79908 175970 79960
rect 176022 79948 176028 79960
rect 176022 79908 176056 79948
rect 176700 79908 176706 79960
rect 176758 79908 176764 79960
rect 176792 79908 176798 79960
rect 176850 79948 176856 79960
rect 177850 79948 177856 79960
rect 176850 79920 177856 79948
rect 176850 79908 176856 79920
rect 177850 79908 177856 79920
rect 177908 79908 177914 79960
rect 175872 79840 175878 79892
rect 175930 79840 175936 79892
rect 175890 79756 175918 79840
rect 176028 79756 176056 79908
rect 176424 79840 176430 79892
rect 176482 79840 176488 79892
rect 176442 79812 176470 79840
rect 176304 79784 176470 79812
rect 176718 79812 176746 79908
rect 177068 79840 177074 79892
rect 177126 79880 177132 79892
rect 178034 79880 178040 79892
rect 177126 79852 178040 79880
rect 177126 79840 177132 79852
rect 178034 79840 178040 79852
rect 178092 79840 178098 79892
rect 177574 79812 177580 79824
rect 176718 79784 177580 79812
rect 175890 79716 175924 79756
rect 175918 79704 175924 79716
rect 175976 79704 175982 79756
rect 176010 79704 176016 79756
rect 176068 79704 176074 79756
rect 175734 79636 175740 79688
rect 175792 79648 175826 79688
rect 175792 79636 175798 79648
rect 176304 79620 176332 79784
rect 177574 79772 177580 79784
rect 177632 79772 177638 79824
rect 177666 79772 177672 79824
rect 177724 79812 177730 79824
rect 181622 79812 181628 79824
rect 177724 79784 181628 79812
rect 177724 79772 177730 79784
rect 181622 79772 181628 79784
rect 181680 79772 181686 79824
rect 174722 79608 174728 79620
rect 174280 79580 174728 79608
rect 174722 79568 174728 79580
rect 174780 79568 174786 79620
rect 174998 79568 175004 79620
rect 175056 79568 175062 79620
rect 175550 79568 175556 79620
rect 175608 79568 175614 79620
rect 175642 79568 175648 79620
rect 175700 79568 175706 79620
rect 176286 79568 176292 79620
rect 176344 79568 176350 79620
rect 177758 79568 177764 79620
rect 177816 79608 177822 79620
rect 214650 79608 214656 79620
rect 177816 79580 214656 79608
rect 177816 79568 177822 79580
rect 214650 79568 214656 79580
rect 214708 79568 214714 79620
rect 171290 79512 171324 79552
rect 171008 79500 171014 79512
rect 171318 79500 171324 79512
rect 171376 79500 171382 79552
rect 171410 79500 171416 79552
rect 171468 79500 171474 79552
rect 171502 79500 171508 79552
rect 171560 79500 171566 79552
rect 179414 79540 179420 79552
rect 171612 79512 179420 79540
rect 168650 79432 168656 79484
rect 168708 79472 168714 79484
rect 171612 79472 171640 79512
rect 179414 79500 179420 79512
rect 179472 79500 179478 79552
rect 181346 79500 181352 79552
rect 181404 79540 181410 79552
rect 202322 79540 202328 79552
rect 181404 79512 202328 79540
rect 181404 79500 181410 79512
rect 202322 79500 202328 79512
rect 202380 79500 202386 79552
rect 168708 79444 171640 79472
rect 168708 79432 168714 79444
rect 172238 79432 172244 79484
rect 172296 79472 172302 79484
rect 192662 79472 192668 79484
rect 172296 79444 192668 79472
rect 172296 79432 172302 79444
rect 192662 79432 192668 79444
rect 192720 79472 192726 79484
rect 324314 79472 324320 79484
rect 192720 79444 324320 79472
rect 192720 79432 192726 79444
rect 324314 79432 324320 79444
rect 324372 79432 324378 79484
rect 167822 79404 167828 79416
rect 162912 79376 166396 79404
rect 167748 79376 167828 79404
rect 162912 79364 162918 79376
rect 108666 79296 108672 79348
rect 108724 79336 108730 79348
rect 122650 79336 122656 79348
rect 108724 79308 122656 79336
rect 108724 79296 108730 79308
rect 122650 79296 122656 79308
rect 122708 79296 122714 79348
rect 122742 79296 122748 79348
rect 122800 79336 122806 79348
rect 135070 79336 135076 79348
rect 122800 79308 135076 79336
rect 122800 79296 122806 79308
rect 135070 79296 135076 79308
rect 135128 79296 135134 79348
rect 136174 79296 136180 79348
rect 136232 79336 136238 79348
rect 143626 79336 143632 79348
rect 136232 79308 143632 79336
rect 136232 79296 136238 79308
rect 143626 79296 143632 79308
rect 143684 79336 143690 79348
rect 144362 79336 144368 79348
rect 143684 79308 144368 79336
rect 143684 79296 143690 79308
rect 144362 79296 144368 79308
rect 144420 79296 144426 79348
rect 119246 79228 119252 79280
rect 119304 79268 119310 79280
rect 135806 79268 135812 79280
rect 119304 79240 135812 79268
rect 119304 79228 119310 79240
rect 135806 79228 135812 79240
rect 135864 79228 135870 79280
rect 146266 79268 146294 79364
rect 148318 79296 148324 79348
rect 148376 79336 148382 79348
rect 165982 79336 165988 79348
rect 148376 79308 165988 79336
rect 148376 79296 148382 79308
rect 165982 79296 165988 79308
rect 166040 79296 166046 79348
rect 135916 79240 146294 79268
rect 116486 79160 116492 79212
rect 116544 79200 116550 79212
rect 135916 79200 135944 79240
rect 152090 79228 152096 79280
rect 152148 79268 152154 79280
rect 153010 79268 153016 79280
rect 152148 79240 153016 79268
rect 152148 79228 152154 79240
rect 153010 79228 153016 79240
rect 153068 79228 153074 79280
rect 158622 79228 158628 79280
rect 158680 79268 158686 79280
rect 166258 79268 166264 79280
rect 158680 79240 166264 79268
rect 158680 79228 158686 79240
rect 166258 79228 166264 79240
rect 166316 79228 166322 79280
rect 166368 79268 166396 79376
rect 167822 79364 167828 79376
rect 167880 79364 167886 79416
rect 170582 79364 170588 79416
rect 170640 79404 170646 79416
rect 170858 79404 170864 79416
rect 170640 79376 170864 79404
rect 170640 79364 170646 79376
rect 170858 79364 170864 79376
rect 170916 79364 170922 79416
rect 172514 79364 172520 79416
rect 172572 79404 172578 79416
rect 179138 79404 179144 79416
rect 172572 79376 179144 79404
rect 172572 79364 172578 79376
rect 179138 79364 179144 79376
rect 179196 79364 179202 79416
rect 179230 79364 179236 79416
rect 179288 79404 179294 79416
rect 214558 79404 214564 79416
rect 179288 79376 214564 79404
rect 179288 79364 179294 79376
rect 214558 79364 214564 79376
rect 214616 79364 214622 79416
rect 214650 79364 214656 79416
rect 214708 79404 214714 79416
rect 358814 79404 358820 79416
rect 214708 79376 358820 79404
rect 214708 79364 214714 79376
rect 358814 79364 358820 79376
rect 358872 79364 358878 79416
rect 166534 79296 166540 79348
rect 166592 79336 166598 79348
rect 166902 79336 166908 79348
rect 166592 79308 166908 79336
rect 166592 79296 166598 79308
rect 166902 79296 166908 79308
rect 166960 79296 166966 79348
rect 167086 79296 167092 79348
rect 167144 79336 167150 79348
rect 180150 79336 180156 79348
rect 167144 79308 180156 79336
rect 167144 79296 167150 79308
rect 180150 79296 180156 79308
rect 180208 79296 180214 79348
rect 184382 79296 184388 79348
rect 184440 79336 184446 79348
rect 194042 79336 194048 79348
rect 184440 79308 194048 79336
rect 184440 79296 184446 79308
rect 194042 79296 194048 79308
rect 194100 79296 194106 79348
rect 376754 79336 376760 79348
rect 200086 79308 376760 79336
rect 191098 79268 191104 79280
rect 166368 79240 191104 79268
rect 191098 79228 191104 79240
rect 191156 79228 191162 79280
rect 116544 79172 135944 79200
rect 116544 79160 116550 79172
rect 136174 79160 136180 79212
rect 136232 79200 136238 79212
rect 146110 79200 146116 79212
rect 136232 79172 146116 79200
rect 136232 79160 136238 79172
rect 146110 79160 146116 79172
rect 146168 79200 146174 79212
rect 147490 79200 147496 79212
rect 146168 79172 147496 79200
rect 146168 79160 146174 79172
rect 147490 79160 147496 79172
rect 147548 79160 147554 79212
rect 150894 79160 150900 79212
rect 150952 79200 150958 79212
rect 156966 79200 156972 79212
rect 150952 79172 156972 79200
rect 150952 79160 150958 79172
rect 156966 79160 156972 79172
rect 157024 79160 157030 79212
rect 157886 79160 157892 79212
rect 157944 79200 157950 79212
rect 158346 79200 158352 79212
rect 157944 79172 158352 79200
rect 157944 79160 157950 79172
rect 158346 79160 158352 79172
rect 158404 79200 158410 79212
rect 188338 79200 188344 79212
rect 158404 79172 188344 79200
rect 158404 79160 158410 79172
rect 188338 79160 188344 79172
rect 188396 79160 188402 79212
rect 113818 79092 113824 79144
rect 113876 79132 113882 79144
rect 126238 79132 126244 79144
rect 113876 79104 126244 79132
rect 113876 79092 113882 79104
rect 126238 79092 126244 79104
rect 126296 79092 126302 79144
rect 126330 79092 126336 79144
rect 126388 79132 126394 79144
rect 135622 79132 135628 79144
rect 126388 79104 135628 79132
rect 126388 79092 126394 79104
rect 135622 79092 135628 79104
rect 135680 79092 135686 79144
rect 135806 79092 135812 79144
rect 135864 79132 135870 79144
rect 145742 79132 145748 79144
rect 135864 79104 145748 79132
rect 135864 79092 135870 79104
rect 145742 79092 145748 79104
rect 145800 79092 145806 79144
rect 161566 79092 161572 79144
rect 161624 79132 161630 79144
rect 161750 79132 161756 79144
rect 161624 79104 161756 79132
rect 161624 79092 161630 79104
rect 161750 79092 161756 79104
rect 161808 79092 161814 79144
rect 164326 79092 164332 79144
rect 164384 79132 164390 79144
rect 165062 79132 165068 79144
rect 164384 79104 165068 79132
rect 164384 79092 164390 79104
rect 165062 79092 165068 79104
rect 165120 79092 165126 79144
rect 166810 79092 166816 79144
rect 166868 79132 166874 79144
rect 196802 79132 196808 79144
rect 166868 79104 196808 79132
rect 166868 79092 166874 79104
rect 196802 79092 196808 79104
rect 196860 79092 196866 79144
rect 116394 79024 116400 79076
rect 116452 79064 116458 79076
rect 150066 79064 150072 79076
rect 116452 79036 150072 79064
rect 116452 79024 116458 79036
rect 150066 79024 150072 79036
rect 150124 79024 150130 79076
rect 158990 79024 158996 79076
rect 159048 79064 159054 79076
rect 159726 79064 159732 79076
rect 159048 79036 159732 79064
rect 159048 79024 159054 79036
rect 159726 79024 159732 79036
rect 159784 79024 159790 79076
rect 160002 79024 160008 79076
rect 160060 79064 160066 79076
rect 193858 79064 193864 79076
rect 160060 79036 193864 79064
rect 160060 79024 160066 79036
rect 193858 79024 193864 79036
rect 193916 79024 193922 79076
rect 115106 78956 115112 79008
rect 115164 78996 115170 79008
rect 147214 78996 147220 79008
rect 115164 78968 147220 78996
rect 115164 78956 115170 78968
rect 147214 78956 147220 78968
rect 147272 78996 147278 79008
rect 147398 78996 147404 79008
rect 147272 78968 147404 78996
rect 147272 78956 147278 78968
rect 147398 78956 147404 78968
rect 147456 78956 147462 79008
rect 161842 78956 161848 79008
rect 161900 78996 161906 79008
rect 196342 78996 196348 79008
rect 161900 78968 196348 78996
rect 161900 78956 161906 78968
rect 196342 78956 196348 78968
rect 196400 78996 196406 79008
rect 200086 78996 200114 79308
rect 376754 79296 376760 79308
rect 376812 79296 376818 79348
rect 196400 78968 200114 78996
rect 196400 78956 196406 78968
rect 113542 78888 113548 78940
rect 113600 78928 113606 78940
rect 147122 78928 147128 78940
rect 113600 78900 147128 78928
rect 113600 78888 113606 78900
rect 147122 78888 147128 78900
rect 147180 78888 147186 78940
rect 158990 78888 158996 78940
rect 159048 78928 159054 78940
rect 159634 78928 159640 78940
rect 159048 78900 159640 78928
rect 159048 78888 159054 78900
rect 159634 78888 159640 78900
rect 159692 78888 159698 78940
rect 166258 78888 166264 78940
rect 166316 78928 166322 78940
rect 172238 78928 172244 78940
rect 166316 78900 172244 78928
rect 166316 78888 166322 78900
rect 172238 78888 172244 78900
rect 172296 78888 172302 78940
rect 173066 78888 173072 78940
rect 173124 78928 173130 78940
rect 212350 78928 212356 78940
rect 173124 78900 212356 78928
rect 173124 78888 173130 78900
rect 212350 78888 212356 78900
rect 212408 78888 212414 78940
rect 115014 78820 115020 78872
rect 115072 78860 115078 78872
rect 147766 78860 147772 78872
rect 115072 78832 147772 78860
rect 115072 78820 115078 78832
rect 147766 78820 147772 78832
rect 147824 78820 147830 78872
rect 166442 78820 166448 78872
rect 166500 78860 166506 78872
rect 166500 78832 174308 78860
rect 166500 78820 166506 78832
rect 127894 78752 127900 78804
rect 127952 78792 127958 78804
rect 130930 78792 130936 78804
rect 127952 78764 130936 78792
rect 127952 78752 127958 78764
rect 130930 78752 130936 78764
rect 130988 78792 130994 78804
rect 135530 78792 135536 78804
rect 130988 78764 135536 78792
rect 130988 78752 130994 78764
rect 135530 78752 135536 78764
rect 135588 78752 135594 78804
rect 143718 78752 143724 78804
rect 143776 78792 143782 78804
rect 144546 78792 144552 78804
rect 143776 78764 144552 78792
rect 143776 78752 143782 78764
rect 144546 78752 144552 78764
rect 144604 78752 144610 78804
rect 159634 78752 159640 78804
rect 159692 78792 159698 78804
rect 159910 78792 159916 78804
rect 159692 78764 159916 78792
rect 159692 78752 159698 78764
rect 159910 78752 159916 78764
rect 159968 78752 159974 78804
rect 160370 78752 160376 78804
rect 160428 78792 160434 78804
rect 161198 78792 161204 78804
rect 160428 78764 161204 78792
rect 160428 78752 160434 78764
rect 161198 78752 161204 78764
rect 161256 78752 161262 78804
rect 127802 78684 127808 78736
rect 127860 78724 127866 78736
rect 131022 78724 131028 78736
rect 127860 78696 131028 78724
rect 127860 78684 127866 78696
rect 131022 78684 131028 78696
rect 131080 78724 131086 78736
rect 145006 78724 145012 78736
rect 131080 78696 145012 78724
rect 131080 78684 131086 78696
rect 145006 78684 145012 78696
rect 145064 78684 145070 78736
rect 153194 78684 153200 78736
rect 153252 78724 153258 78736
rect 153930 78724 153936 78736
rect 153252 78696 153936 78724
rect 153252 78684 153258 78696
rect 153930 78684 153936 78696
rect 153988 78684 153994 78736
rect 169938 78684 169944 78736
rect 169996 78724 170002 78736
rect 170582 78724 170588 78736
rect 169996 78696 170588 78724
rect 169996 78684 170002 78696
rect 170582 78684 170588 78696
rect 170640 78684 170646 78736
rect 171042 78684 171048 78736
rect 171100 78724 171106 78736
rect 171686 78724 171692 78736
rect 171100 78696 171692 78724
rect 171100 78684 171106 78696
rect 171686 78684 171692 78696
rect 171744 78684 171750 78736
rect 171962 78684 171968 78736
rect 172020 78724 172026 78736
rect 172238 78724 172244 78736
rect 172020 78696 172244 78724
rect 172020 78684 172026 78696
rect 172238 78684 172244 78696
rect 172296 78684 172302 78736
rect 172422 78684 172428 78736
rect 172480 78724 172486 78736
rect 173342 78724 173348 78736
rect 172480 78696 173348 78724
rect 172480 78684 172486 78696
rect 173342 78684 173348 78696
rect 173400 78684 173406 78736
rect 174280 78724 174308 78832
rect 175366 78820 175372 78872
rect 175424 78860 175430 78872
rect 176010 78860 176016 78872
rect 175424 78832 176016 78860
rect 175424 78820 175430 78832
rect 176010 78820 176016 78832
rect 176068 78860 176074 78872
rect 176068 78832 190454 78860
rect 176068 78820 176074 78832
rect 174538 78752 174544 78804
rect 174596 78792 174602 78804
rect 190426 78792 190454 78832
rect 210418 78792 210424 78804
rect 174596 78764 186314 78792
rect 190426 78764 210424 78792
rect 174596 78752 174602 78764
rect 178770 78724 178776 78736
rect 174280 78696 178776 78724
rect 178770 78684 178776 78696
rect 178828 78684 178834 78736
rect 186286 78724 186314 78764
rect 210418 78752 210424 78764
rect 210476 78752 210482 78804
rect 212442 78752 212448 78804
rect 212500 78792 212506 78804
rect 480254 78792 480260 78804
rect 212500 78764 480260 78792
rect 212500 78752 212506 78764
rect 480254 78752 480260 78764
rect 480312 78752 480318 78804
rect 201034 78724 201040 78736
rect 186286 78696 201040 78724
rect 201034 78684 201040 78696
rect 201092 78724 201098 78736
rect 539686 78724 539692 78736
rect 201092 78696 539692 78724
rect 201092 78684 201098 78696
rect 539686 78684 539692 78696
rect 539744 78684 539750 78736
rect 106826 78616 106832 78668
rect 106884 78656 106890 78668
rect 107562 78656 107568 78668
rect 106884 78628 107568 78656
rect 106884 78616 106890 78628
rect 107562 78616 107568 78628
rect 107620 78616 107626 78668
rect 135622 78616 135628 78668
rect 135680 78656 135686 78668
rect 142430 78656 142436 78668
rect 135680 78628 142436 78656
rect 135680 78616 135686 78628
rect 142430 78616 142436 78628
rect 142488 78616 142494 78668
rect 153470 78616 153476 78668
rect 153528 78656 153534 78668
rect 153654 78656 153660 78668
rect 153528 78628 153660 78656
rect 153528 78616 153534 78628
rect 153654 78616 153660 78628
rect 153712 78616 153718 78668
rect 157426 78616 157432 78668
rect 157484 78656 157490 78668
rect 157610 78656 157616 78668
rect 157484 78628 157616 78656
rect 157484 78616 157490 78628
rect 157610 78616 157616 78628
rect 157668 78616 157674 78668
rect 158806 78616 158812 78668
rect 158864 78656 158870 78668
rect 159082 78656 159088 78668
rect 158864 78628 159088 78656
rect 158864 78616 158870 78628
rect 159082 78616 159088 78628
rect 159140 78616 159146 78668
rect 160830 78616 160836 78668
rect 160888 78656 160894 78668
rect 162210 78656 162216 78668
rect 160888 78628 162216 78656
rect 160888 78616 160894 78628
rect 162210 78616 162216 78628
rect 162268 78616 162274 78668
rect 168650 78616 168656 78668
rect 168708 78656 168714 78668
rect 169202 78656 169208 78668
rect 168708 78628 169208 78656
rect 168708 78616 168714 78628
rect 169202 78616 169208 78628
rect 169260 78616 169266 78668
rect 169662 78616 169668 78668
rect 169720 78656 169726 78668
rect 169720 78628 176654 78656
rect 169720 78616 169726 78628
rect 98914 78548 98920 78600
rect 98972 78588 98978 78600
rect 150618 78588 150624 78600
rect 98972 78560 150624 78588
rect 98972 78548 98978 78560
rect 150618 78548 150624 78560
rect 150676 78588 150682 78600
rect 151170 78588 151176 78600
rect 150676 78560 151176 78588
rect 150676 78548 150682 78560
rect 151170 78548 151176 78560
rect 151228 78548 151234 78600
rect 176626 78588 176654 78628
rect 176838 78616 176844 78668
rect 176896 78656 176902 78668
rect 177574 78656 177580 78668
rect 176896 78628 177580 78656
rect 176896 78616 176902 78628
rect 177574 78616 177580 78628
rect 177632 78616 177638 78668
rect 212074 78588 212080 78600
rect 176626 78560 212080 78588
rect 212074 78548 212080 78560
rect 212132 78588 212138 78600
rect 212442 78588 212448 78600
rect 212132 78560 212448 78588
rect 212132 78548 212138 78560
rect 212442 78548 212448 78560
rect 212500 78548 212506 78600
rect 103974 78480 103980 78532
rect 104032 78520 104038 78532
rect 104342 78520 104348 78532
rect 104032 78492 104348 78520
rect 104032 78480 104038 78492
rect 104342 78480 104348 78492
rect 104400 78480 104406 78532
rect 132494 78480 132500 78532
rect 132552 78520 132558 78532
rect 136174 78520 136180 78532
rect 132552 78492 136180 78520
rect 132552 78480 132558 78492
rect 136174 78480 136180 78492
rect 136232 78480 136238 78532
rect 152182 78480 152188 78532
rect 152240 78520 152246 78532
rect 153470 78520 153476 78532
rect 152240 78492 153476 78520
rect 152240 78480 152246 78492
rect 153470 78480 153476 78492
rect 153528 78480 153534 78532
rect 158898 78480 158904 78532
rect 158956 78520 158962 78532
rect 163406 78520 163412 78532
rect 158956 78492 163412 78520
rect 158956 78480 158962 78492
rect 163406 78480 163412 78492
rect 163464 78480 163470 78532
rect 164878 78480 164884 78532
rect 164936 78520 164942 78532
rect 178678 78520 178684 78532
rect 164936 78492 178684 78520
rect 164936 78480 164942 78492
rect 178678 78480 178684 78492
rect 178736 78480 178742 78532
rect 205818 78480 205824 78532
rect 205876 78520 205882 78532
rect 205876 78492 205956 78520
rect 205876 78480 205882 78492
rect 110414 78412 110420 78464
rect 110472 78452 110478 78464
rect 110874 78452 110880 78464
rect 110472 78424 110880 78452
rect 110472 78412 110478 78424
rect 110874 78412 110880 78424
rect 110932 78452 110938 78464
rect 140958 78452 140964 78464
rect 110932 78424 140964 78452
rect 110932 78412 110938 78424
rect 140958 78412 140964 78424
rect 141016 78412 141022 78464
rect 157150 78412 157156 78464
rect 157208 78452 157214 78464
rect 161290 78452 161296 78464
rect 157208 78424 161296 78452
rect 157208 78412 157214 78424
rect 161290 78412 161296 78424
rect 161348 78412 161354 78464
rect 181438 78412 181444 78464
rect 181496 78452 181502 78464
rect 202138 78452 202144 78464
rect 181496 78424 202144 78452
rect 181496 78412 181502 78424
rect 202138 78412 202144 78424
rect 202196 78412 202202 78464
rect 105630 78344 105636 78396
rect 105688 78384 105694 78396
rect 136634 78384 136640 78396
rect 105688 78356 136640 78384
rect 105688 78344 105694 78356
rect 136634 78344 136640 78356
rect 136692 78344 136698 78396
rect 168742 78344 168748 78396
rect 168800 78384 168806 78396
rect 203150 78384 203156 78396
rect 168800 78356 203156 78384
rect 168800 78344 168806 78356
rect 203150 78344 203156 78356
rect 203208 78384 203214 78396
rect 204162 78384 204168 78396
rect 203208 78356 204168 78384
rect 203208 78344 203214 78356
rect 204162 78344 204168 78356
rect 204220 78344 204226 78396
rect 205928 78328 205956 78492
rect 207474 78344 207480 78396
rect 207532 78384 207538 78396
rect 207934 78384 207940 78396
rect 207532 78356 207940 78384
rect 207532 78344 207538 78356
rect 207934 78344 207940 78356
rect 207992 78344 207998 78396
rect 60734 78276 60740 78328
rect 60792 78316 60798 78328
rect 107194 78316 107200 78328
rect 60792 78288 107200 78316
rect 60792 78276 60798 78288
rect 107194 78276 107200 78288
rect 107252 78316 107258 78328
rect 133690 78316 133696 78328
rect 107252 78288 133696 78316
rect 107252 78276 107258 78288
rect 133690 78276 133696 78288
rect 133748 78276 133754 78328
rect 136910 78316 136916 78328
rect 133984 78288 136916 78316
rect 75914 78208 75920 78260
rect 75972 78248 75978 78260
rect 104434 78248 104440 78260
rect 75972 78220 104440 78248
rect 75972 78208 75978 78220
rect 104434 78208 104440 78220
rect 104492 78208 104498 78260
rect 133984 78248 134012 78288
rect 136910 78276 136916 78288
rect 136968 78276 136974 78328
rect 165706 78276 165712 78328
rect 165764 78316 165770 78328
rect 166442 78316 166448 78328
rect 165764 78288 166448 78316
rect 165764 78276 165770 78288
rect 166442 78276 166448 78288
rect 166500 78276 166506 78328
rect 169018 78276 169024 78328
rect 169076 78316 169082 78328
rect 203334 78316 203340 78328
rect 169076 78288 203340 78316
rect 169076 78276 169082 78288
rect 203334 78276 203340 78288
rect 203392 78316 203398 78328
rect 204070 78316 204076 78328
rect 203392 78288 204076 78316
rect 203392 78276 203398 78288
rect 204070 78276 204076 78288
rect 204128 78276 204134 78328
rect 205910 78276 205916 78328
rect 205968 78276 205974 78328
rect 107948 78220 134012 78248
rect 57974 78072 57980 78124
rect 58032 78112 58038 78124
rect 107286 78112 107292 78124
rect 58032 78084 107292 78112
rect 58032 78072 58038 78084
rect 107286 78072 107292 78084
rect 107344 78112 107350 78124
rect 107948 78112 107976 78220
rect 135070 78208 135076 78260
rect 135128 78248 135134 78260
rect 149606 78248 149612 78260
rect 135128 78220 149612 78248
rect 135128 78208 135134 78220
rect 149606 78208 149612 78220
rect 149664 78248 149670 78260
rect 153010 78248 153016 78260
rect 149664 78220 153016 78248
rect 149664 78208 149670 78220
rect 153010 78208 153016 78220
rect 153068 78208 153074 78260
rect 163222 78208 163228 78260
rect 163280 78248 163286 78260
rect 166626 78248 166632 78260
rect 163280 78220 166632 78248
rect 163280 78208 163286 78220
rect 166626 78208 166632 78220
rect 166684 78208 166690 78260
rect 168006 78208 168012 78260
rect 168064 78248 168070 78260
rect 199010 78248 199016 78260
rect 168064 78220 199016 78248
rect 168064 78208 168070 78220
rect 199010 78208 199016 78220
rect 199068 78208 199074 78260
rect 136266 78180 136272 78192
rect 107344 78084 107976 78112
rect 108040 78152 136272 78180
rect 107344 78072 107350 78084
rect 53834 78004 53840 78056
rect 53892 78044 53898 78056
rect 105630 78044 105636 78056
rect 53892 78016 105636 78044
rect 53892 78004 53898 78016
rect 105630 78004 105636 78016
rect 105688 78004 105694 78056
rect 46934 77936 46940 77988
rect 46992 77976 46998 77988
rect 107102 77976 107108 77988
rect 46992 77948 107108 77976
rect 46992 77936 46998 77948
rect 107102 77936 107108 77948
rect 107160 77976 107166 77988
rect 108040 77976 108068 78152
rect 136266 78140 136272 78152
rect 136324 78140 136330 78192
rect 165798 78140 165804 78192
rect 165856 78180 165862 78192
rect 171870 78180 171876 78192
rect 165856 78152 171876 78180
rect 165856 78140 165862 78152
rect 171870 78140 171876 78152
rect 171928 78140 171934 78192
rect 175458 78140 175464 78192
rect 175516 78180 175522 78192
rect 176378 78180 176384 78192
rect 175516 78152 176384 78180
rect 175516 78140 175522 78152
rect 176378 78140 176384 78152
rect 176436 78140 176442 78192
rect 180702 78140 180708 78192
rect 180760 78180 180766 78192
rect 207842 78180 207848 78192
rect 180760 78152 207848 78180
rect 180760 78140 180766 78152
rect 207842 78140 207848 78152
rect 207900 78140 207906 78192
rect 122098 78072 122104 78124
rect 122156 78112 122162 78124
rect 148686 78112 148692 78124
rect 122156 78084 148692 78112
rect 122156 78072 122162 78084
rect 148686 78072 148692 78084
rect 148744 78072 148750 78124
rect 164050 78072 164056 78124
rect 164108 78112 164114 78124
rect 178770 78112 178776 78124
rect 164108 78084 178776 78112
rect 164108 78072 164114 78084
rect 178770 78072 178776 78084
rect 178828 78072 178834 78124
rect 179138 78072 179144 78124
rect 179196 78112 179202 78124
rect 197906 78112 197912 78124
rect 179196 78084 197912 78112
rect 179196 78072 179202 78084
rect 197906 78072 197912 78084
rect 197964 78072 197970 78124
rect 199010 78072 199016 78124
rect 199068 78112 199074 78124
rect 199562 78112 199568 78124
rect 199068 78084 199568 78112
rect 199068 78072 199074 78084
rect 199562 78072 199568 78084
rect 199620 78112 199626 78124
rect 456794 78112 456800 78124
rect 199620 78084 456800 78112
rect 199620 78072 199626 78084
rect 456794 78072 456800 78084
rect 456852 78072 456858 78124
rect 129826 78044 129832 78056
rect 107160 77948 108068 77976
rect 108132 78016 129832 78044
rect 107160 77936 107166 77948
rect 107010 77868 107016 77920
rect 107068 77908 107074 77920
rect 108132 77908 108160 78016
rect 129826 78004 129832 78016
rect 129884 78044 129890 78056
rect 134334 78044 134340 78056
rect 129884 78016 134340 78044
rect 129884 78004 129890 78016
rect 134334 78004 134340 78016
rect 134392 78004 134398 78056
rect 163590 78004 163596 78056
rect 163648 78044 163654 78056
rect 179322 78044 179328 78056
rect 163648 78016 179328 78044
rect 163648 78004 163654 78016
rect 179322 78004 179328 78016
rect 179380 78044 179386 78056
rect 195146 78044 195152 78056
rect 179380 78016 195152 78044
rect 179380 78004 179386 78016
rect 195146 78004 195152 78016
rect 195204 78004 195210 78056
rect 204162 78004 204168 78056
rect 204220 78044 204226 78056
rect 465166 78044 465172 78056
rect 204220 78016 465172 78044
rect 204220 78004 204226 78016
rect 465166 78004 465172 78016
rect 465224 78004 465230 78056
rect 108390 77936 108396 77988
rect 108448 77976 108454 77988
rect 108448 77948 118694 77976
rect 108448 77936 108454 77948
rect 107068 77880 108160 77908
rect 107068 77868 107074 77880
rect 118666 77704 118694 77948
rect 159726 77936 159732 77988
rect 159784 77976 159790 77988
rect 159910 77976 159916 77988
rect 159784 77948 159916 77976
rect 159784 77936 159790 77948
rect 159910 77936 159916 77948
rect 159968 77936 159974 77988
rect 160186 77936 160192 77988
rect 160244 77976 160250 77988
rect 162302 77976 162308 77988
rect 160244 77948 162308 77976
rect 160244 77936 160250 77948
rect 162302 77936 162308 77948
rect 162360 77936 162366 77988
rect 165798 77936 165804 77988
rect 165856 77976 165862 77988
rect 166534 77976 166540 77988
rect 165856 77948 166540 77976
rect 165856 77936 165862 77948
rect 166534 77936 166540 77948
rect 166592 77936 166598 77988
rect 167546 77936 167552 77988
rect 167604 77976 167610 77988
rect 168098 77976 168104 77988
rect 167604 77948 168104 77976
rect 167604 77936 167610 77948
rect 168098 77936 168104 77948
rect 168156 77936 168162 77988
rect 180518 77976 180524 77988
rect 171796 77948 180524 77976
rect 121914 77868 121920 77920
rect 121972 77908 121978 77920
rect 122098 77908 122104 77920
rect 121972 77880 122104 77908
rect 121972 77868 121978 77880
rect 122098 77868 122104 77880
rect 122156 77908 122162 77920
rect 132310 77908 132316 77920
rect 122156 77880 132316 77908
rect 122156 77868 122162 77880
rect 132310 77868 132316 77880
rect 132368 77868 132374 77920
rect 161658 77868 161664 77920
rect 161716 77908 161722 77920
rect 164050 77908 164056 77920
rect 161716 77880 164056 77908
rect 161716 77868 161722 77880
rect 164050 77868 164056 77880
rect 164108 77868 164114 77920
rect 165154 77868 165160 77920
rect 165212 77908 165218 77920
rect 171796 77908 171824 77948
rect 180518 77936 180524 77948
rect 180576 77976 180582 77988
rect 180702 77976 180708 77988
rect 180576 77948 180708 77976
rect 180576 77936 180582 77948
rect 180702 77936 180708 77948
rect 180760 77936 180766 77988
rect 200942 77976 200948 77988
rect 186286 77948 200948 77976
rect 165212 77880 171824 77908
rect 165212 77868 165218 77880
rect 171870 77868 171876 77920
rect 171928 77908 171934 77920
rect 181898 77908 181904 77920
rect 171928 77880 181904 77908
rect 171928 77868 171934 77880
rect 181898 77868 181904 77880
rect 181956 77908 181962 77920
rect 186286 77908 186314 77948
rect 200942 77936 200948 77948
rect 201000 77936 201006 77988
rect 204070 77936 204076 77988
rect 204128 77976 204134 77988
rect 471974 77976 471980 77988
rect 204128 77948 471980 77976
rect 204128 77936 204134 77948
rect 471974 77936 471980 77948
rect 472032 77936 472038 77988
rect 181956 77880 186314 77908
rect 181956 77868 181962 77880
rect 166350 77800 166356 77852
rect 166408 77840 166414 77852
rect 180702 77840 180708 77852
rect 166408 77812 180708 77840
rect 166408 77800 166414 77812
rect 180702 77800 180708 77812
rect 180760 77800 180766 77852
rect 125594 77732 125600 77784
rect 125652 77772 125658 77784
rect 139670 77772 139676 77784
rect 125652 77744 139676 77772
rect 125652 77732 125658 77744
rect 139670 77732 139676 77744
rect 139728 77732 139734 77784
rect 167638 77732 167644 77784
rect 167696 77772 167702 77784
rect 181622 77772 181628 77784
rect 167696 77744 181628 77772
rect 167696 77732 167702 77744
rect 181622 77732 181628 77744
rect 181680 77732 181686 77784
rect 131298 77704 131304 77716
rect 118666 77676 131304 77704
rect 131298 77664 131304 77676
rect 131356 77704 131362 77716
rect 142522 77704 142528 77716
rect 131356 77676 142528 77704
rect 131356 77664 131362 77676
rect 142522 77664 142528 77676
rect 142580 77664 142586 77716
rect 163038 77664 163044 77716
rect 163096 77704 163102 77716
rect 172514 77704 172520 77716
rect 163096 77676 172520 77704
rect 163096 77664 163102 77676
rect 172514 77664 172520 77676
rect 172572 77664 172578 77716
rect 178034 77664 178040 77716
rect 178092 77704 178098 77716
rect 211890 77704 211896 77716
rect 178092 77676 211896 77704
rect 178092 77664 178098 77676
rect 211890 77664 211896 77676
rect 211948 77664 211954 77716
rect 104434 77596 104440 77648
rect 104492 77636 104498 77648
rect 137830 77636 137836 77648
rect 104492 77608 137836 77636
rect 104492 77596 104498 77608
rect 137830 77596 137836 77608
rect 137888 77596 137894 77648
rect 149330 77596 149336 77648
rect 149388 77636 149394 77648
rect 209130 77636 209136 77648
rect 149388 77608 209136 77636
rect 149388 77596 149394 77608
rect 209130 77596 209136 77608
rect 209188 77596 209194 77648
rect 107562 77528 107568 77580
rect 107620 77568 107626 77580
rect 141234 77568 141240 77580
rect 107620 77540 141240 77568
rect 107620 77528 107626 77540
rect 141234 77528 141240 77540
rect 141292 77528 141298 77580
rect 154666 77528 154672 77580
rect 154724 77568 154730 77580
rect 155034 77568 155040 77580
rect 154724 77540 155040 77568
rect 154724 77528 154730 77540
rect 155034 77528 155040 77540
rect 155092 77528 155098 77580
rect 167638 77528 167644 77580
rect 167696 77568 167702 77580
rect 167822 77568 167828 77580
rect 167696 77540 167828 77568
rect 167696 77528 167702 77540
rect 167822 77528 167828 77540
rect 167880 77528 167886 77580
rect 174722 77528 174728 77580
rect 174780 77568 174786 77580
rect 177574 77568 177580 77580
rect 174780 77540 177580 77568
rect 174780 77528 174786 77540
rect 177574 77528 177580 77540
rect 177632 77528 177638 77580
rect 118878 77460 118884 77512
rect 118936 77500 118942 77512
rect 131666 77500 131672 77512
rect 118936 77472 131672 77500
rect 118936 77460 118942 77472
rect 131666 77460 131672 77472
rect 131724 77500 131730 77512
rect 134518 77500 134524 77512
rect 131724 77472 134524 77500
rect 131724 77460 131730 77472
rect 134518 77460 134524 77472
rect 134576 77460 134582 77512
rect 175458 77460 175464 77512
rect 175516 77500 175522 77512
rect 176654 77500 176660 77512
rect 175516 77472 176660 77500
rect 175516 77460 175522 77472
rect 176654 77460 176660 77472
rect 176712 77460 176718 77512
rect 122006 77392 122012 77444
rect 122064 77432 122070 77444
rect 124858 77432 124864 77444
rect 122064 77404 124864 77432
rect 122064 77392 122070 77404
rect 124858 77392 124864 77404
rect 124916 77392 124922 77444
rect 142982 77392 142988 77444
rect 143040 77432 143046 77444
rect 143258 77432 143264 77444
rect 143040 77404 143264 77432
rect 143040 77392 143046 77404
rect 143258 77392 143264 77404
rect 143316 77392 143322 77444
rect 162118 77392 162124 77444
rect 162176 77432 162182 77444
rect 162854 77432 162860 77444
rect 162176 77404 162860 77432
rect 162176 77392 162182 77404
rect 162854 77392 162860 77404
rect 162912 77392 162918 77444
rect 173986 77392 173992 77444
rect 174044 77432 174050 77444
rect 174998 77432 175004 77444
rect 174044 77404 175004 77432
rect 174044 77392 174050 77404
rect 174998 77392 175004 77404
rect 175056 77392 175062 77444
rect 176286 77392 176292 77444
rect 176344 77432 176350 77444
rect 176562 77432 176568 77444
rect 176344 77404 176568 77432
rect 176344 77392 176350 77404
rect 176562 77392 176568 77404
rect 176620 77392 176626 77444
rect 161106 77324 161112 77376
rect 161164 77364 161170 77376
rect 161164 77336 164234 77364
rect 161164 77324 161170 77336
rect 153194 77256 153200 77308
rect 153252 77296 153258 77308
rect 154022 77296 154028 77308
rect 153252 77268 154028 77296
rect 153252 77256 153258 77268
rect 154022 77256 154028 77268
rect 154080 77256 154086 77308
rect 156690 77256 156696 77308
rect 156748 77296 156754 77308
rect 157150 77296 157156 77308
rect 156748 77268 157156 77296
rect 156748 77256 156754 77268
rect 157150 77256 157156 77268
rect 157208 77256 157214 77308
rect 161842 77256 161848 77308
rect 161900 77296 161906 77308
rect 162670 77296 162676 77308
rect 161900 77268 162676 77296
rect 161900 77256 161906 77268
rect 162670 77256 162676 77268
rect 162728 77256 162734 77308
rect 164206 77296 164234 77336
rect 167362 77324 167368 77376
rect 167420 77364 167426 77376
rect 181438 77364 181444 77376
rect 167420 77336 181444 77364
rect 167420 77324 167426 77336
rect 181438 77324 181444 77336
rect 181496 77324 181502 77376
rect 166442 77296 166448 77308
rect 164206 77268 166448 77296
rect 166442 77256 166448 77268
rect 166500 77256 166506 77308
rect 172882 77256 172888 77308
rect 172940 77296 172946 77308
rect 177482 77296 177488 77308
rect 172940 77268 177488 77296
rect 172940 77256 172946 77268
rect 177482 77256 177488 77268
rect 177540 77256 177546 77308
rect 97626 77188 97632 77240
rect 97684 77228 97690 77240
rect 137646 77228 137652 77240
rect 97684 77200 137652 77228
rect 97684 77188 97690 77200
rect 137646 77188 137652 77200
rect 137704 77188 137710 77240
rect 151722 77188 151728 77240
rect 151780 77228 151786 77240
rect 151906 77228 151912 77240
rect 151780 77200 151912 77228
rect 151780 77188 151786 77200
rect 151906 77188 151912 77200
rect 151964 77188 151970 77240
rect 162118 77188 162124 77240
rect 162176 77228 162182 77240
rect 213914 77228 213920 77240
rect 162176 77200 213920 77228
rect 162176 77188 162182 77200
rect 213914 77188 213920 77200
rect 213972 77228 213978 77240
rect 213972 77200 219434 77228
rect 213972 77188 213978 77200
rect 113726 77120 113732 77172
rect 113784 77160 113790 77172
rect 146662 77160 146668 77172
rect 113784 77132 146668 77160
rect 113784 77120 113790 77132
rect 146662 77120 146668 77132
rect 146720 77160 146726 77172
rect 148502 77160 148508 77172
rect 146720 77132 148508 77160
rect 146720 77120 146726 77132
rect 148502 77120 148508 77132
rect 148560 77120 148566 77172
rect 154850 77120 154856 77172
rect 154908 77160 154914 77172
rect 155218 77160 155224 77172
rect 154908 77132 155224 77160
rect 154908 77120 154914 77132
rect 155218 77120 155224 77132
rect 155276 77120 155282 77172
rect 155494 77120 155500 77172
rect 155552 77160 155558 77172
rect 214282 77160 214288 77172
rect 155552 77132 214288 77160
rect 155552 77120 155558 77132
rect 214282 77120 214288 77132
rect 214340 77160 214346 77172
rect 214558 77160 214564 77172
rect 214340 77132 214564 77160
rect 214340 77120 214346 77132
rect 214558 77120 214564 77132
rect 214616 77120 214622 77172
rect 104158 77052 104164 77104
rect 104216 77092 104222 77104
rect 104434 77092 104440 77104
rect 104216 77064 104440 77092
rect 104216 77052 104222 77064
rect 104434 77052 104440 77064
rect 104492 77092 104498 77104
rect 136726 77092 136732 77104
rect 104492 77064 136732 77092
rect 104492 77052 104498 77064
rect 136726 77052 136732 77064
rect 136784 77052 136790 77104
rect 158070 77052 158076 77104
rect 158128 77092 158134 77104
rect 158128 77064 209774 77092
rect 158128 77052 158134 77064
rect 104066 76984 104072 77036
rect 104124 77024 104130 77036
rect 104342 77024 104348 77036
rect 104124 76996 104348 77024
rect 104124 76984 104130 76996
rect 104342 76984 104348 76996
rect 104400 77024 104406 77036
rect 137002 77024 137008 77036
rect 104400 76996 137008 77024
rect 104400 76984 104406 76996
rect 137002 76984 137008 76996
rect 137060 76984 137066 77036
rect 138290 76984 138296 77036
rect 138348 77024 138354 77036
rect 138566 77024 138572 77036
rect 138348 76996 138572 77024
rect 138348 76984 138354 76996
rect 138566 76984 138572 76996
rect 138624 76984 138630 77036
rect 154666 76984 154672 77036
rect 154724 77024 154730 77036
rect 155494 77024 155500 77036
rect 154724 76996 155500 77024
rect 154724 76984 154730 76996
rect 155494 76984 155500 76996
rect 155552 76984 155558 77036
rect 160830 76984 160836 77036
rect 160888 77024 160894 77036
rect 195330 77024 195336 77036
rect 160888 76996 195336 77024
rect 160888 76984 160894 76996
rect 195330 76984 195336 76996
rect 195388 76984 195394 77036
rect 114186 76916 114192 76968
rect 114244 76956 114250 76968
rect 142890 76956 142896 76968
rect 114244 76928 142896 76956
rect 114244 76916 114250 76928
rect 142890 76916 142896 76928
rect 142948 76916 142954 76968
rect 147030 76956 147036 76968
rect 143000 76928 147036 76956
rect 115658 76848 115664 76900
rect 115716 76888 115722 76900
rect 143000 76888 143028 76928
rect 147030 76916 147036 76928
rect 147088 76916 147094 76968
rect 162486 76916 162492 76968
rect 162544 76956 162550 76968
rect 162854 76956 162860 76968
rect 162544 76928 162860 76956
rect 162544 76916 162550 76928
rect 162854 76916 162860 76928
rect 162912 76916 162918 76968
rect 168190 76916 168196 76968
rect 168248 76956 168254 76968
rect 168248 76928 174584 76956
rect 168248 76916 168254 76928
rect 145650 76888 145656 76900
rect 115716 76860 143028 76888
rect 143092 76860 145656 76888
rect 115716 76848 115722 76860
rect 114094 76780 114100 76832
rect 114152 76820 114158 76832
rect 143092 76820 143120 76860
rect 145650 76848 145656 76860
rect 145708 76848 145714 76900
rect 159634 76848 159640 76900
rect 159692 76888 159698 76900
rect 174556 76888 174584 76928
rect 175642 76916 175648 76968
rect 175700 76956 175706 76968
rect 175826 76956 175832 76968
rect 175700 76928 175832 76956
rect 175700 76916 175706 76928
rect 175826 76916 175832 76928
rect 175884 76916 175890 76968
rect 175918 76916 175924 76968
rect 175976 76956 175982 76968
rect 207658 76956 207664 76968
rect 175976 76928 207664 76956
rect 175976 76916 175982 76928
rect 207658 76916 207664 76928
rect 207716 76916 207722 76968
rect 190822 76888 190828 76900
rect 159692 76860 166994 76888
rect 174556 76860 190828 76888
rect 159692 76848 159698 76860
rect 114152 76792 143120 76820
rect 114152 76780 114158 76792
rect 143994 76780 144000 76832
rect 144052 76820 144058 76832
rect 147030 76820 147036 76832
rect 144052 76792 147036 76820
rect 144052 76780 144058 76792
rect 147030 76780 147036 76792
rect 147088 76780 147094 76832
rect 166966 76820 166994 76860
rect 190822 76848 190828 76860
rect 190880 76848 190886 76900
rect 192386 76820 192392 76832
rect 166966 76792 192392 76820
rect 192386 76780 192392 76792
rect 192444 76820 192450 76832
rect 209746 76820 209774 77064
rect 219406 76888 219434 77200
rect 253934 76888 253940 76900
rect 219406 76860 253940 76888
rect 253934 76848 253940 76860
rect 253992 76848 253998 76900
rect 214466 76820 214472 76832
rect 192444 76792 200114 76820
rect 209746 76792 214472 76820
rect 192444 76780 192450 76792
rect 117958 76712 117964 76764
rect 118016 76752 118022 76764
rect 147950 76752 147956 76764
rect 118016 76724 147956 76752
rect 118016 76712 118022 76724
rect 147950 76712 147956 76724
rect 148008 76752 148014 76764
rect 148686 76752 148692 76764
rect 148008 76724 148692 76752
rect 148008 76712 148014 76724
rect 148686 76712 148692 76724
rect 148744 76712 148750 76764
rect 153470 76712 153476 76764
rect 153528 76752 153534 76764
rect 162118 76752 162124 76764
rect 153528 76724 162124 76752
rect 153528 76712 153534 76724
rect 162118 76712 162124 76724
rect 162176 76712 162182 76764
rect 162302 76712 162308 76764
rect 162360 76752 162366 76764
rect 162360 76724 190454 76752
rect 162360 76712 162366 76724
rect 67634 76644 67640 76696
rect 67692 76684 67698 76696
rect 97626 76684 97632 76696
rect 67692 76656 97632 76684
rect 67692 76644 67698 76656
rect 97626 76644 97632 76656
rect 97684 76644 97690 76696
rect 114002 76644 114008 76696
rect 114060 76684 114066 76696
rect 114060 76656 131114 76684
rect 114060 76644 114066 76656
rect 66254 76576 66260 76628
rect 66312 76616 66318 76628
rect 104434 76616 104440 76628
rect 66312 76588 104440 76616
rect 66312 76576 66318 76588
rect 104434 76576 104440 76588
rect 104492 76576 104498 76628
rect 114278 76576 114284 76628
rect 114336 76616 114342 76628
rect 126238 76616 126244 76628
rect 114336 76588 126244 76616
rect 114336 76576 114342 76588
rect 126238 76576 126244 76588
rect 126296 76576 126302 76628
rect 131086 76616 131114 76656
rect 133874 76644 133880 76696
rect 133932 76684 133938 76696
rect 134150 76684 134156 76696
rect 133932 76656 134156 76684
rect 133932 76644 133938 76656
rect 134150 76644 134156 76656
rect 134208 76644 134214 76696
rect 137554 76684 137560 76696
rect 134444 76656 137560 76684
rect 134444 76616 134472 76656
rect 137554 76644 137560 76656
rect 137612 76644 137618 76696
rect 143534 76644 143540 76696
rect 143592 76684 143598 76696
rect 144086 76684 144092 76696
rect 143592 76656 144092 76684
rect 143592 76644 143598 76656
rect 144086 76644 144092 76656
rect 144144 76644 144150 76696
rect 147214 76644 147220 76696
rect 147272 76684 147278 76696
rect 180058 76684 180064 76696
rect 147272 76656 180064 76684
rect 147272 76644 147278 76656
rect 180058 76644 180064 76656
rect 180116 76644 180122 76696
rect 131086 76588 134472 76616
rect 135346 76576 135352 76628
rect 135404 76616 135410 76628
rect 135530 76616 135536 76628
rect 135404 76588 135536 76616
rect 135404 76576 135410 76588
rect 135530 76576 135536 76588
rect 135588 76576 135594 76628
rect 135898 76576 135904 76628
rect 135956 76616 135962 76628
rect 136358 76616 136364 76628
rect 135956 76588 136364 76616
rect 135956 76576 135962 76588
rect 136358 76576 136364 76588
rect 136416 76576 136422 76628
rect 137002 76576 137008 76628
rect 137060 76616 137066 76628
rect 137738 76616 137744 76628
rect 137060 76588 137744 76616
rect 137060 76576 137066 76588
rect 137738 76576 137744 76588
rect 137796 76576 137802 76628
rect 138106 76576 138112 76628
rect 138164 76616 138170 76628
rect 138290 76616 138296 76628
rect 138164 76588 138296 76616
rect 138164 76576 138170 76588
rect 138290 76576 138296 76588
rect 138348 76576 138354 76628
rect 140038 76576 140044 76628
rect 140096 76616 140102 76628
rect 140406 76616 140412 76628
rect 140096 76588 140412 76616
rect 140096 76576 140102 76588
rect 140406 76576 140412 76588
rect 140464 76576 140470 76628
rect 142890 76576 142896 76628
rect 142948 76616 142954 76628
rect 146754 76616 146760 76628
rect 142948 76588 146760 76616
rect 142948 76576 142954 76588
rect 146754 76576 146760 76588
rect 146812 76616 146818 76628
rect 146812 76588 149054 76616
rect 146812 76576 146818 76588
rect 59354 76508 59360 76560
rect 59412 76548 59418 76560
rect 104342 76548 104348 76560
rect 59412 76520 104348 76548
rect 59412 76508 59418 76520
rect 104342 76508 104348 76520
rect 104400 76508 104406 76560
rect 112714 76508 112720 76560
rect 112772 76548 112778 76560
rect 143810 76548 143816 76560
rect 112772 76520 143816 76548
rect 112772 76508 112778 76520
rect 143810 76508 143816 76520
rect 143868 76508 143874 76560
rect 149026 76548 149054 76588
rect 150066 76576 150072 76628
rect 150124 76616 150130 76628
rect 182818 76616 182824 76628
rect 150124 76588 182824 76616
rect 150124 76576 150130 76588
rect 182818 76576 182824 76588
rect 182876 76576 182882 76628
rect 190426 76616 190454 76724
rect 200086 76684 200114 76792
rect 214466 76780 214472 76792
rect 214524 76820 214530 76832
rect 289814 76820 289820 76832
rect 214524 76792 289820 76820
rect 214524 76780 214530 76792
rect 289814 76780 289820 76792
rect 289872 76780 289878 76832
rect 214558 76712 214564 76764
rect 214616 76752 214622 76764
rect 296714 76752 296720 76764
rect 214616 76724 296720 76752
rect 214616 76712 214622 76724
rect 296714 76712 296720 76724
rect 296772 76712 296778 76764
rect 353294 76684 353300 76696
rect 200086 76656 353300 76684
rect 353294 76644 353300 76656
rect 353352 76644 353358 76696
rect 195238 76616 195244 76628
rect 190426 76588 195244 76616
rect 195238 76576 195244 76588
rect 195296 76616 195302 76628
rect 357526 76616 357532 76628
rect 195296 76588 357532 76616
rect 195296 76576 195302 76588
rect 357526 76576 357532 76588
rect 357584 76576 357590 76628
rect 184934 76548 184940 76560
rect 149026 76520 184940 76548
rect 184934 76508 184940 76520
rect 184992 76508 184998 76560
rect 195330 76508 195336 76560
rect 195388 76548 195394 76560
rect 367094 76548 367100 76560
rect 195388 76520 367100 76548
rect 195388 76508 195394 76520
rect 367094 76508 367100 76520
rect 367152 76508 367158 76560
rect 112438 76440 112444 76492
rect 112496 76480 112502 76492
rect 126974 76480 126980 76492
rect 112496 76452 126980 76480
rect 112496 76440 112502 76452
rect 126974 76440 126980 76452
rect 127032 76440 127038 76492
rect 134334 76440 134340 76492
rect 134392 76480 134398 76492
rect 134886 76480 134892 76492
rect 134392 76452 134892 76480
rect 134392 76440 134398 76452
rect 134886 76440 134892 76452
rect 134944 76440 134950 76492
rect 135714 76440 135720 76492
rect 135772 76480 135778 76492
rect 136542 76480 136548 76492
rect 135772 76452 136548 76480
rect 135772 76440 135778 76452
rect 136542 76440 136548 76452
rect 136600 76440 136606 76492
rect 139394 76440 139400 76492
rect 139452 76480 139458 76492
rect 141878 76480 141884 76492
rect 139452 76452 141884 76480
rect 139452 76440 139458 76452
rect 141878 76440 141884 76452
rect 141936 76440 141942 76492
rect 164326 76440 164332 76492
rect 164384 76480 164390 76492
rect 164878 76480 164884 76492
rect 164384 76452 164884 76480
rect 164384 76440 164390 76452
rect 164878 76440 164884 76452
rect 164936 76440 164942 76492
rect 170582 76440 170588 76492
rect 170640 76480 170646 76492
rect 199286 76480 199292 76492
rect 170640 76452 199292 76480
rect 170640 76440 170646 76452
rect 199286 76440 199292 76452
rect 199344 76440 199350 76492
rect 129642 76372 129648 76424
rect 129700 76412 129706 76424
rect 142154 76412 142160 76424
rect 129700 76384 142160 76412
rect 129700 76372 129706 76384
rect 142154 76372 142160 76384
rect 142212 76372 142218 76424
rect 154574 76372 154580 76424
rect 154632 76412 154638 76424
rect 155126 76412 155132 76424
rect 154632 76384 155132 76412
rect 154632 76372 154638 76384
rect 155126 76372 155132 76384
rect 155184 76372 155190 76424
rect 163958 76372 163964 76424
rect 164016 76412 164022 76424
rect 165062 76412 165068 76424
rect 164016 76384 165068 76412
rect 164016 76372 164022 76384
rect 165062 76372 165068 76384
rect 165120 76412 165126 76424
rect 192846 76412 192852 76424
rect 165120 76384 192852 76412
rect 165120 76372 165126 76384
rect 192846 76372 192852 76384
rect 192904 76372 192910 76424
rect 134242 76304 134248 76356
rect 134300 76344 134306 76356
rect 135162 76344 135168 76356
rect 134300 76316 135168 76344
rect 134300 76304 134306 76316
rect 135162 76304 135168 76316
rect 135220 76304 135226 76356
rect 139762 76304 139768 76356
rect 139820 76344 139826 76356
rect 140222 76344 140228 76356
rect 139820 76316 140228 76344
rect 139820 76304 139826 76316
rect 140222 76304 140228 76316
rect 140280 76304 140286 76356
rect 141694 76304 141700 76356
rect 141752 76344 141758 76356
rect 146018 76344 146024 76356
rect 141752 76316 146024 76344
rect 141752 76304 141758 76316
rect 146018 76304 146024 76316
rect 146076 76304 146082 76356
rect 173342 76304 173348 76356
rect 173400 76344 173406 76356
rect 173802 76344 173808 76356
rect 173400 76316 173808 76344
rect 173400 76304 173406 76316
rect 173802 76304 173808 76316
rect 173860 76304 173866 76356
rect 174078 76304 174084 76356
rect 174136 76344 174142 76356
rect 174630 76344 174636 76356
rect 174136 76316 174636 76344
rect 174136 76304 174142 76316
rect 174630 76304 174636 76316
rect 174688 76304 174694 76356
rect 181622 76304 181628 76356
rect 181680 76344 181686 76356
rect 181898 76344 181904 76356
rect 181680 76316 181904 76344
rect 181680 76304 181686 76316
rect 181898 76304 181904 76316
rect 181956 76344 181962 76356
rect 201494 76344 201500 76356
rect 181956 76316 201500 76344
rect 181956 76304 181962 76316
rect 201494 76304 201500 76316
rect 201552 76304 201558 76356
rect 139670 76236 139676 76288
rect 139728 76276 139734 76288
rect 140590 76276 140596 76288
rect 139728 76248 140596 76276
rect 139728 76236 139734 76248
rect 140590 76236 140596 76248
rect 140648 76236 140654 76288
rect 180426 76236 180432 76288
rect 180484 76276 180490 76288
rect 180702 76276 180708 76288
rect 180484 76248 180708 76276
rect 180484 76236 180490 76248
rect 180702 76236 180708 76248
rect 180760 76276 180766 76288
rect 214374 76276 214380 76288
rect 180760 76248 214380 76276
rect 180760 76236 180766 76248
rect 214374 76236 214380 76248
rect 214432 76236 214438 76288
rect 126238 76168 126244 76220
rect 126296 76208 126302 76220
rect 140314 76208 140320 76220
rect 126296 76180 140320 76208
rect 126296 76168 126302 76180
rect 140314 76168 140320 76180
rect 140372 76168 140378 76220
rect 140958 76168 140964 76220
rect 141016 76208 141022 76220
rect 141418 76208 141424 76220
rect 141016 76180 141424 76208
rect 141016 76168 141022 76180
rect 141418 76168 141424 76180
rect 141476 76168 141482 76220
rect 156046 76168 156052 76220
rect 156104 76208 156110 76220
rect 161014 76208 161020 76220
rect 156104 76180 161020 76208
rect 156104 76168 156110 76180
rect 161014 76168 161020 76180
rect 161072 76168 161078 76220
rect 162118 76168 162124 76220
rect 162176 76208 162182 76220
rect 162946 76208 162952 76220
rect 162176 76180 162952 76208
rect 162176 76168 162182 76180
rect 162946 76168 162952 76180
rect 163004 76168 163010 76220
rect 174354 76168 174360 76220
rect 174412 76208 174418 76220
rect 174998 76208 175004 76220
rect 174412 76180 175004 76208
rect 174412 76168 174418 76180
rect 174998 76168 175004 76180
rect 175056 76168 175062 76220
rect 126974 76100 126980 76152
rect 127032 76140 127038 76152
rect 141970 76140 141976 76152
rect 127032 76112 141976 76140
rect 127032 76100 127038 76112
rect 141970 76100 141976 76112
rect 142028 76100 142034 76152
rect 144178 76100 144184 76152
rect 144236 76140 144242 76152
rect 144914 76140 144920 76152
rect 144236 76112 144920 76140
rect 144236 76100 144242 76112
rect 144914 76100 144920 76112
rect 144972 76100 144978 76152
rect 172790 76100 172796 76152
rect 172848 76140 172854 76152
rect 177206 76140 177212 76152
rect 172848 76112 177212 76140
rect 172848 76100 172854 76112
rect 177206 76100 177212 76112
rect 177264 76100 177270 76152
rect 139486 76032 139492 76084
rect 139544 76072 139550 76084
rect 140222 76072 140228 76084
rect 139544 76044 140228 76072
rect 139544 76032 139550 76044
rect 140222 76032 140228 76044
rect 140280 76032 140286 76084
rect 162578 76032 162584 76084
rect 162636 76072 162642 76084
rect 168006 76072 168012 76084
rect 162636 76044 168012 76072
rect 162636 76032 162642 76044
rect 168006 76032 168012 76044
rect 168064 76032 168070 76084
rect 172698 76032 172704 76084
rect 172756 76072 172762 76084
rect 178402 76072 178408 76084
rect 172756 76044 178408 76072
rect 172756 76032 172762 76044
rect 178402 76032 178408 76044
rect 178460 76032 178466 76084
rect 173526 75964 173532 76016
rect 173584 76004 173590 76016
rect 173710 76004 173716 76016
rect 173584 75976 173716 76004
rect 173584 75964 173590 75976
rect 173710 75964 173716 75976
rect 173768 75964 173774 76016
rect 167822 75896 167828 75948
rect 167880 75936 167886 75948
rect 168190 75936 168196 75948
rect 167880 75908 168196 75936
rect 167880 75896 167886 75908
rect 168190 75896 168196 75908
rect 168248 75896 168254 75948
rect 108574 75828 108580 75880
rect 108632 75868 108638 75880
rect 113174 75868 113180 75880
rect 108632 75840 113180 75868
rect 108632 75828 108638 75840
rect 113174 75828 113180 75840
rect 113232 75868 113238 75880
rect 114278 75868 114284 75880
rect 113232 75840 114284 75868
rect 113232 75828 113238 75840
rect 114278 75828 114284 75840
rect 114336 75828 114342 75880
rect 123938 75828 123944 75880
rect 123996 75868 124002 75880
rect 148226 75868 148232 75880
rect 123996 75840 148232 75868
rect 123996 75828 124002 75840
rect 148226 75828 148232 75840
rect 148284 75868 148290 75880
rect 148284 75840 151814 75868
rect 148284 75828 148290 75840
rect 112806 75760 112812 75812
rect 112864 75800 112870 75812
rect 146202 75800 146208 75812
rect 112864 75772 146208 75800
rect 112864 75760 112870 75772
rect 146202 75760 146208 75772
rect 146260 75800 146266 75812
rect 146478 75800 146484 75812
rect 146260 75772 146484 75800
rect 146260 75760 146266 75772
rect 146478 75760 146484 75772
rect 146536 75760 146542 75812
rect 102870 75692 102876 75744
rect 102928 75732 102934 75744
rect 135162 75732 135168 75744
rect 102928 75704 135168 75732
rect 102928 75692 102934 75704
rect 135162 75692 135168 75704
rect 135220 75692 135226 75744
rect 136726 75692 136732 75744
rect 136784 75732 136790 75744
rect 138014 75732 138020 75744
rect 136784 75704 138020 75732
rect 136784 75692 136790 75704
rect 138014 75692 138020 75704
rect 138072 75692 138078 75744
rect 151786 75732 151814 75840
rect 171502 75828 171508 75880
rect 171560 75868 171566 75880
rect 172054 75868 172060 75880
rect 171560 75840 172060 75868
rect 171560 75828 171566 75840
rect 172054 75828 172060 75840
rect 172112 75868 172118 75880
rect 175826 75868 175832 75880
rect 172112 75840 175832 75868
rect 172112 75828 172118 75840
rect 175826 75828 175832 75840
rect 175884 75828 175890 75880
rect 176654 75828 176660 75880
rect 176712 75868 176718 75880
rect 185026 75868 185032 75880
rect 176712 75840 185032 75868
rect 176712 75828 176718 75840
rect 185026 75828 185032 75840
rect 185084 75828 185090 75880
rect 185118 75828 185124 75880
rect 185176 75868 185182 75880
rect 212902 75868 212908 75880
rect 185176 75840 212908 75868
rect 185176 75828 185182 75840
rect 212902 75828 212908 75840
rect 212960 75828 212966 75880
rect 172330 75760 172336 75812
rect 172388 75800 172394 75812
rect 206370 75800 206376 75812
rect 172388 75772 206376 75800
rect 172388 75760 172394 75772
rect 206370 75760 206376 75772
rect 206428 75760 206434 75812
rect 159542 75732 159548 75744
rect 151786 75704 159548 75732
rect 159542 75692 159548 75704
rect 159600 75692 159606 75744
rect 171226 75692 171232 75744
rect 171284 75732 171290 75744
rect 205818 75732 205824 75744
rect 171284 75704 205824 75732
rect 171284 75692 171290 75704
rect 205818 75692 205824 75704
rect 205876 75692 205882 75744
rect 116854 75624 116860 75676
rect 116912 75664 116918 75676
rect 147306 75664 147312 75676
rect 116912 75636 147312 75664
rect 116912 75624 116918 75636
rect 147306 75624 147312 75636
rect 147364 75624 147370 75676
rect 175826 75624 175832 75676
rect 175884 75664 175890 75676
rect 206002 75664 206008 75676
rect 175884 75636 206008 75664
rect 175884 75624 175890 75636
rect 206002 75624 206008 75636
rect 206060 75624 206066 75676
rect 114186 75556 114192 75608
rect 114244 75596 114250 75608
rect 144270 75596 144276 75608
rect 114244 75568 144276 75596
rect 114244 75556 114250 75568
rect 144270 75556 144276 75568
rect 144328 75556 144334 75608
rect 159744 75568 161520 75596
rect 117130 75488 117136 75540
rect 117188 75528 117194 75540
rect 145558 75528 145564 75540
rect 117188 75500 145564 75528
rect 117188 75488 117194 75500
rect 145558 75488 145564 75500
rect 145616 75488 145622 75540
rect 157058 75488 157064 75540
rect 157116 75528 157122 75540
rect 159082 75528 159088 75540
rect 157116 75500 159088 75528
rect 157116 75488 157122 75500
rect 159082 75488 159088 75500
rect 159140 75488 159146 75540
rect 159744 75472 159772 75568
rect 160370 75488 160376 75540
rect 160428 75528 160434 75540
rect 161382 75528 161388 75540
rect 160428 75500 161388 75528
rect 160428 75488 160434 75500
rect 161382 75488 161388 75500
rect 161440 75488 161446 75540
rect 161492 75528 161520 75568
rect 171778 75556 171784 75608
rect 171836 75596 171842 75608
rect 205910 75596 205916 75608
rect 171836 75568 205916 75596
rect 171836 75556 171842 75568
rect 205910 75556 205916 75568
rect 205968 75556 205974 75608
rect 192202 75528 192208 75540
rect 161492 75500 192208 75528
rect 192202 75488 192208 75500
rect 192260 75488 192266 75540
rect 118418 75420 118424 75472
rect 118476 75460 118482 75472
rect 135254 75460 135260 75472
rect 118476 75432 135260 75460
rect 118476 75420 118482 75432
rect 135254 75420 135260 75432
rect 135312 75420 135318 75472
rect 157334 75420 157340 75472
rect 157392 75460 157398 75472
rect 157610 75460 157616 75472
rect 157392 75432 157616 75460
rect 157392 75420 157398 75432
rect 157610 75420 157616 75432
rect 157668 75420 157674 75472
rect 158806 75420 158812 75472
rect 158864 75460 158870 75472
rect 159726 75460 159732 75472
rect 158864 75432 159732 75460
rect 158864 75420 158870 75432
rect 159726 75420 159732 75432
rect 159784 75420 159790 75472
rect 160186 75420 160192 75472
rect 160244 75460 160250 75472
rect 160738 75460 160744 75472
rect 160244 75432 160744 75460
rect 160244 75420 160250 75432
rect 160738 75420 160744 75432
rect 160796 75420 160802 75472
rect 161566 75420 161572 75472
rect 161624 75460 161630 75472
rect 162394 75460 162400 75472
rect 161624 75432 162400 75460
rect 161624 75420 161630 75432
rect 162394 75420 162400 75432
rect 162452 75420 162458 75472
rect 163038 75420 163044 75472
rect 163096 75460 163102 75472
rect 163774 75460 163780 75472
rect 163096 75432 163780 75460
rect 163096 75420 163102 75432
rect 163774 75420 163780 75432
rect 163832 75420 163838 75472
rect 168466 75420 168472 75472
rect 168524 75460 168530 75472
rect 169018 75460 169024 75472
rect 168524 75432 169024 75460
rect 168524 75420 168530 75432
rect 169018 75420 169024 75432
rect 169076 75420 169082 75472
rect 178402 75420 178408 75472
rect 178460 75460 178466 75472
rect 207474 75460 207480 75472
rect 178460 75432 207480 75460
rect 178460 75420 178466 75432
rect 207474 75420 207480 75432
rect 207532 75420 207538 75472
rect 120994 75352 121000 75404
rect 121052 75392 121058 75404
rect 136174 75392 136180 75404
rect 121052 75364 136180 75392
rect 121052 75352 121058 75364
rect 136174 75352 136180 75364
rect 136232 75352 136238 75404
rect 141786 75392 141792 75404
rect 140746 75364 141792 75392
rect 121178 75284 121184 75336
rect 121236 75324 121242 75336
rect 131114 75324 131120 75336
rect 121236 75296 131120 75324
rect 121236 75284 121242 75296
rect 131114 75284 131120 75296
rect 131172 75284 131178 75336
rect 85574 75216 85580 75268
rect 85632 75256 85638 75268
rect 103882 75256 103888 75268
rect 85632 75228 103888 75256
rect 85632 75216 85638 75228
rect 103882 75216 103888 75228
rect 103940 75256 103946 75268
rect 104434 75256 104440 75268
rect 103940 75228 104440 75256
rect 103940 75216 103946 75228
rect 104434 75216 104440 75228
rect 104492 75216 104498 75268
rect 106918 75216 106924 75268
rect 106976 75256 106982 75268
rect 131482 75256 131488 75268
rect 106976 75228 131488 75256
rect 106976 75216 106982 75228
rect 131482 75216 131488 75228
rect 131540 75256 131546 75268
rect 140746 75256 140774 75364
rect 141786 75352 141792 75364
rect 141844 75352 141850 75404
rect 153010 75352 153016 75404
rect 153068 75392 153074 75404
rect 216674 75392 216680 75404
rect 153068 75364 216680 75392
rect 153068 75352 153074 75364
rect 216674 75352 216680 75364
rect 216732 75352 216738 75404
rect 148502 75284 148508 75336
rect 148560 75324 148566 75336
rect 157058 75324 157064 75336
rect 148560 75296 157064 75324
rect 148560 75284 148566 75296
rect 157058 75284 157064 75296
rect 157116 75284 157122 75336
rect 159082 75284 159088 75336
rect 159140 75324 159146 75336
rect 176654 75324 176660 75336
rect 159140 75296 176660 75324
rect 159140 75284 159146 75296
rect 176654 75284 176660 75296
rect 176712 75284 176718 75336
rect 176746 75284 176752 75336
rect 176804 75324 176810 75336
rect 177022 75324 177028 75336
rect 176804 75296 177028 75324
rect 176804 75284 176810 75296
rect 177022 75284 177028 75296
rect 177080 75284 177086 75336
rect 177206 75284 177212 75336
rect 177264 75324 177270 75336
rect 177758 75324 177764 75336
rect 177264 75296 177764 75324
rect 177264 75284 177270 75296
rect 177758 75284 177764 75296
rect 177816 75324 177822 75336
rect 185118 75324 185124 75336
rect 177816 75296 185124 75324
rect 177816 75284 177822 75296
rect 185118 75284 185124 75296
rect 185176 75284 185182 75336
rect 205818 75284 205824 75336
rect 205876 75324 205882 75336
rect 478138 75324 478144 75336
rect 205876 75296 478144 75324
rect 205876 75284 205882 75296
rect 478138 75284 478144 75296
rect 478196 75284 478202 75336
rect 131540 75228 140774 75256
rect 131540 75216 131546 75228
rect 145466 75216 145472 75268
rect 145524 75256 145530 75268
rect 147214 75256 147220 75268
rect 145524 75228 147220 75256
rect 145524 75216 145530 75228
rect 147214 75216 147220 75228
rect 147272 75216 147278 75268
rect 147398 75216 147404 75268
rect 147456 75256 147462 75268
rect 193858 75256 193864 75268
rect 147456 75228 157104 75256
rect 147456 75216 147462 75228
rect 99190 75148 99196 75200
rect 99248 75188 99254 75200
rect 131390 75188 131396 75200
rect 99248 75160 131396 75188
rect 99248 75148 99254 75160
rect 131390 75148 131396 75160
rect 131448 75148 131454 75200
rect 131574 75148 131580 75200
rect 131632 75188 131638 75200
rect 133138 75188 133144 75200
rect 131632 75160 133144 75188
rect 131632 75148 131638 75160
rect 133138 75148 133144 75160
rect 133196 75148 133202 75200
rect 136174 75148 136180 75200
rect 136232 75188 136238 75200
rect 146570 75188 146576 75200
rect 136232 75160 146576 75188
rect 136232 75148 136238 75160
rect 146570 75148 146576 75160
rect 146628 75148 146634 75200
rect 152090 75148 152096 75200
rect 152148 75188 152154 75200
rect 152918 75188 152924 75200
rect 152148 75160 152924 75188
rect 152148 75148 152154 75160
rect 152918 75148 152924 75160
rect 152976 75148 152982 75200
rect 154022 75148 154028 75200
rect 154080 75188 154086 75200
rect 154390 75188 154396 75200
rect 154080 75160 154396 75188
rect 154080 75148 154086 75160
rect 154390 75148 154396 75160
rect 154448 75148 154454 75200
rect 157076 75188 157104 75228
rect 157260 75228 193864 75256
rect 157260 75188 157288 75228
rect 193858 75216 193864 75228
rect 193916 75216 193922 75268
rect 205910 75216 205916 75268
rect 205968 75256 205974 75268
rect 506474 75256 506480 75268
rect 205968 75228 506480 75256
rect 205968 75216 205974 75228
rect 506474 75216 506480 75228
rect 506532 75216 506538 75268
rect 157076 75160 157288 75188
rect 159542 75148 159548 75200
rect 159600 75188 159606 75200
rect 201494 75188 201500 75200
rect 159600 75160 201500 75188
rect 159600 75148 159606 75160
rect 201494 75148 201500 75160
rect 201552 75148 201558 75200
rect 207474 75148 207480 75200
rect 207532 75188 207538 75200
rect 517514 75188 517520 75200
rect 207532 75160 517520 75188
rect 207532 75148 207538 75160
rect 517514 75148 517520 75160
rect 517572 75148 517578 75200
rect 120626 75080 120632 75132
rect 120684 75120 120690 75132
rect 144178 75120 144184 75132
rect 120684 75092 144184 75120
rect 120684 75080 120690 75092
rect 144178 75080 144184 75092
rect 144236 75080 144242 75132
rect 151814 75080 151820 75132
rect 151872 75120 151878 75132
rect 152458 75120 152464 75132
rect 151872 75092 152464 75120
rect 151872 75080 151878 75092
rect 152458 75080 152464 75092
rect 152516 75080 152522 75132
rect 156046 75080 156052 75132
rect 156104 75120 156110 75132
rect 157242 75120 157248 75132
rect 156104 75092 157248 75120
rect 156104 75080 156110 75092
rect 157242 75080 157248 75092
rect 157300 75080 157306 75132
rect 157426 75080 157432 75132
rect 157484 75120 157490 75132
rect 158162 75120 158168 75132
rect 157484 75092 158168 75120
rect 157484 75080 157490 75092
rect 158162 75080 158168 75092
rect 158220 75080 158226 75132
rect 158806 75080 158812 75132
rect 158864 75120 158870 75132
rect 159818 75120 159824 75132
rect 158864 75092 159824 75120
rect 158864 75080 158870 75092
rect 159818 75080 159824 75092
rect 159876 75080 159882 75132
rect 160370 75080 160376 75132
rect 160428 75120 160434 75132
rect 160554 75120 160560 75132
rect 160428 75092 160560 75120
rect 160428 75080 160434 75092
rect 160554 75080 160560 75092
rect 160612 75080 160618 75132
rect 161658 75080 161664 75132
rect 161716 75120 161722 75132
rect 162026 75120 162032 75132
rect 161716 75092 162032 75120
rect 161716 75080 161722 75092
rect 162026 75080 162032 75092
rect 162084 75080 162090 75132
rect 162946 75080 162952 75132
rect 163004 75120 163010 75132
rect 163314 75120 163320 75132
rect 163004 75092 163320 75120
rect 163004 75080 163010 75092
rect 163314 75080 163320 75092
rect 163372 75080 163378 75132
rect 164326 75080 164332 75132
rect 164384 75120 164390 75132
rect 164510 75120 164516 75132
rect 164384 75092 164516 75120
rect 164384 75080 164390 75092
rect 164510 75080 164516 75092
rect 164568 75080 164574 75132
rect 165982 75080 165988 75132
rect 166040 75120 166046 75132
rect 166166 75120 166172 75132
rect 166040 75092 166172 75120
rect 166040 75080 166046 75092
rect 166166 75080 166172 75092
rect 166224 75080 166230 75132
rect 168926 75080 168932 75132
rect 168984 75120 168990 75132
rect 169478 75120 169484 75132
rect 168984 75092 169484 75120
rect 168984 75080 168990 75092
rect 169478 75080 169484 75092
rect 169536 75080 169542 75132
rect 174998 75080 175004 75132
rect 175056 75120 175062 75132
rect 206278 75120 206284 75132
rect 175056 75092 206284 75120
rect 175056 75080 175062 75092
rect 206278 75080 206284 75092
rect 206336 75080 206342 75132
rect 104434 75012 104440 75064
rect 104492 75052 104498 75064
rect 138842 75052 138848 75064
rect 104492 75024 138848 75052
rect 104492 75012 104498 75024
rect 138842 75012 138848 75024
rect 138900 75012 138906 75064
rect 146202 75012 146208 75064
rect 146260 75052 146266 75064
rect 180794 75052 180800 75064
rect 146260 75024 180800 75052
rect 146260 75012 146266 75024
rect 180794 75012 180800 75024
rect 180852 75012 180858 75064
rect 108482 74944 108488 74996
rect 108540 74984 108546 74996
rect 125594 74984 125600 74996
rect 108540 74956 125600 74984
rect 108540 74944 108546 74956
rect 125594 74944 125600 74956
rect 125652 74944 125658 74996
rect 165614 74944 165620 74996
rect 165672 74984 165678 74996
rect 166166 74984 166172 74996
rect 165672 74956 166172 74984
rect 165672 74944 165678 74956
rect 166166 74944 166172 74956
rect 166224 74944 166230 74996
rect 168742 74944 168748 74996
rect 168800 74984 168806 74996
rect 169110 74984 169116 74996
rect 168800 74956 169116 74984
rect 168800 74944 168806 74956
rect 169110 74944 169116 74956
rect 169168 74944 169174 74996
rect 176654 74944 176660 74996
rect 176712 74984 176718 74996
rect 177298 74984 177304 74996
rect 176712 74956 177304 74984
rect 176712 74944 176718 74956
rect 177298 74944 177304 74956
rect 177356 74944 177362 74996
rect 135254 74876 135260 74928
rect 135312 74916 135318 74928
rect 145466 74916 145472 74928
rect 135312 74888 145472 74916
rect 135312 74876 135318 74888
rect 145466 74876 145472 74888
rect 145524 74876 145530 74928
rect 164602 74876 164608 74928
rect 164660 74916 164666 74928
rect 165246 74916 165252 74928
rect 164660 74888 165252 74916
rect 164660 74876 164666 74888
rect 165246 74876 165252 74888
rect 165304 74876 165310 74928
rect 168466 74876 168472 74928
rect 168524 74916 168530 74928
rect 169294 74916 169300 74928
rect 168524 74888 169300 74916
rect 168524 74876 168530 74888
rect 169294 74876 169300 74888
rect 169352 74876 169358 74928
rect 165614 74808 165620 74860
rect 165672 74848 165678 74860
rect 166902 74848 166908 74860
rect 165672 74820 166908 74848
rect 165672 74808 165678 74820
rect 166902 74808 166908 74820
rect 166960 74808 166966 74860
rect 138474 74672 138480 74724
rect 138532 74712 138538 74724
rect 139302 74712 139308 74724
rect 138532 74684 139308 74712
rect 138532 74672 138538 74684
rect 139302 74672 139308 74684
rect 139360 74672 139366 74724
rect 131114 74536 131120 74588
rect 131172 74576 131178 74588
rect 134794 74576 134800 74588
rect 131172 74548 134800 74576
rect 131172 74536 131178 74548
rect 134794 74536 134800 74548
rect 134852 74536 134858 74588
rect 206370 74536 206376 74588
rect 206428 74576 206434 74588
rect 511258 74576 511264 74588
rect 206428 74548 511264 74576
rect 206428 74536 206434 74548
rect 511258 74536 511264 74548
rect 511316 74536 511322 74588
rect 104250 74468 104256 74520
rect 104308 74508 104314 74520
rect 138658 74508 138664 74520
rect 104308 74480 138664 74508
rect 104308 74468 104314 74480
rect 138658 74468 138664 74480
rect 138716 74468 138722 74520
rect 142154 74468 142160 74520
rect 142212 74508 142218 74520
rect 143258 74508 143264 74520
rect 142212 74480 143264 74508
rect 142212 74468 142218 74480
rect 143258 74468 143264 74480
rect 143316 74468 143322 74520
rect 152274 74468 152280 74520
rect 152332 74508 152338 74520
rect 211522 74508 211528 74520
rect 152332 74480 211528 74508
rect 152332 74468 152338 74480
rect 211522 74468 211528 74480
rect 211580 74468 211586 74520
rect 109678 74400 109684 74452
rect 109736 74440 109742 74452
rect 142338 74440 142344 74452
rect 109736 74412 142344 74440
rect 109736 74400 109742 74412
rect 142338 74400 142344 74412
rect 142396 74400 142402 74452
rect 142798 74400 142804 74452
rect 142856 74440 142862 74452
rect 143442 74440 143448 74452
rect 142856 74412 143448 74440
rect 142856 74400 142862 74412
rect 143442 74400 143448 74412
rect 143500 74400 143506 74452
rect 145374 74400 145380 74452
rect 145432 74440 145438 74452
rect 146018 74440 146024 74452
rect 145432 74412 146024 74440
rect 145432 74400 145438 74412
rect 146018 74400 146024 74412
rect 146076 74400 146082 74452
rect 171318 74400 171324 74452
rect 171376 74440 171382 74452
rect 172238 74440 172244 74452
rect 171376 74412 172244 74440
rect 171376 74400 171382 74412
rect 172238 74400 172244 74412
rect 172296 74400 172302 74452
rect 204714 74440 204720 74452
rect 176626 74412 204720 74440
rect 100386 74332 100392 74384
rect 100444 74372 100450 74384
rect 129090 74372 129096 74384
rect 100444 74344 129096 74372
rect 100444 74332 100450 74344
rect 129090 74332 129096 74344
rect 129148 74332 129154 74384
rect 170858 74332 170864 74384
rect 170916 74372 170922 74384
rect 176626 74372 176654 74412
rect 204714 74400 204720 74412
rect 204772 74400 204778 74452
rect 170916 74344 176654 74372
rect 170916 74332 170922 74344
rect 177390 74332 177396 74384
rect 177448 74372 177454 74384
rect 211614 74372 211620 74384
rect 177448 74344 211620 74372
rect 177448 74332 177454 74344
rect 211614 74332 211620 74344
rect 211672 74332 211678 74384
rect 116670 74264 116676 74316
rect 116728 74304 116734 74316
rect 149698 74304 149704 74316
rect 116728 74276 149704 74304
rect 116728 74264 116734 74276
rect 149698 74264 149704 74276
rect 149756 74304 149762 74316
rect 149974 74304 149980 74316
rect 149756 74276 149980 74304
rect 149756 74264 149762 74276
rect 149974 74264 149980 74276
rect 150032 74264 150038 74316
rect 153378 74264 153384 74316
rect 153436 74304 153442 74316
rect 188062 74304 188068 74316
rect 153436 74276 188068 74304
rect 153436 74264 153442 74276
rect 188062 74264 188068 74276
rect 188120 74264 188126 74316
rect 109862 74196 109868 74248
rect 109920 74236 109926 74248
rect 142798 74236 142804 74248
rect 109920 74208 142804 74236
rect 109920 74196 109926 74208
rect 142798 74196 142804 74208
rect 142856 74196 142862 74248
rect 143442 74196 143448 74248
rect 143500 74236 143506 74248
rect 143810 74236 143816 74248
rect 143500 74208 143816 74236
rect 143500 74196 143506 74208
rect 143810 74196 143816 74208
rect 143868 74196 143874 74248
rect 153654 74196 153660 74248
rect 153712 74236 153718 74248
rect 154206 74236 154212 74248
rect 153712 74208 154212 74236
rect 153712 74196 153718 74208
rect 154206 74196 154212 74208
rect 154264 74236 154270 74248
rect 187142 74236 187148 74248
rect 154264 74208 187148 74236
rect 154264 74196 154270 74208
rect 187142 74196 187148 74208
rect 187200 74196 187206 74248
rect 111702 74128 111708 74180
rect 111760 74168 111766 74180
rect 144086 74168 144092 74180
rect 111760 74140 144092 74168
rect 111760 74128 111766 74140
rect 144086 74128 144092 74140
rect 144144 74128 144150 74180
rect 172238 74128 172244 74180
rect 172296 74168 172302 74180
rect 203702 74168 203708 74180
rect 172296 74140 203708 74168
rect 172296 74128 172302 74140
rect 203702 74128 203708 74140
rect 203760 74128 203766 74180
rect 108758 74060 108764 74112
rect 108816 74100 108822 74112
rect 140498 74100 140504 74112
rect 108816 74072 140504 74100
rect 108816 74060 108822 74072
rect 140498 74060 140504 74072
rect 140556 74060 140562 74112
rect 171686 74060 171692 74112
rect 171744 74100 171750 74112
rect 203610 74100 203616 74112
rect 171744 74072 203616 74100
rect 171744 74060 171750 74072
rect 203610 74060 203616 74072
rect 203668 74060 203674 74112
rect 119890 73992 119896 74044
rect 119948 74032 119954 74044
rect 151722 74032 151728 74044
rect 119948 74004 151728 74032
rect 119948 73992 119954 74004
rect 151722 73992 151728 74004
rect 151780 73992 151786 74044
rect 163406 73992 163412 74044
rect 163464 74032 163470 74044
rect 193766 74032 193772 74044
rect 163464 74004 193772 74032
rect 163464 73992 163470 74004
rect 193766 73992 193772 74004
rect 193824 73992 193830 74044
rect 89714 73924 89720 73976
rect 89772 73964 89778 73976
rect 104250 73964 104256 73976
rect 89772 73936 104256 73964
rect 89772 73924 89778 73936
rect 104250 73924 104256 73936
rect 104308 73924 104314 73976
rect 121270 73924 121276 73976
rect 121328 73964 121334 73976
rect 152182 73964 152188 73976
rect 121328 73936 152188 73964
rect 121328 73924 121334 73936
rect 152182 73924 152188 73936
rect 152240 73924 152246 73976
rect 161382 73924 161388 73976
rect 161440 73964 161446 73976
rect 186958 73964 186964 73976
rect 161440 73936 186964 73964
rect 161440 73924 161446 73936
rect 186958 73924 186964 73936
rect 187016 73924 187022 73976
rect 211522 73924 211528 73976
rect 211580 73964 211586 73976
rect 255314 73964 255320 73976
rect 211580 73936 255320 73964
rect 211580 73924 211586 73936
rect 255314 73924 255320 73936
rect 255372 73924 255378 73976
rect 22738 73856 22744 73908
rect 22796 73896 22802 73908
rect 100386 73896 100392 73908
rect 22796 73868 100392 73896
rect 22796 73856 22802 73868
rect 100386 73856 100392 73868
rect 100444 73856 100450 73908
rect 112990 73856 112996 73908
rect 113048 73896 113054 73908
rect 142154 73896 142160 73908
rect 113048 73868 142160 73896
rect 113048 73856 113054 73868
rect 142154 73856 142160 73868
rect 142212 73856 142218 73908
rect 146386 73856 146392 73908
rect 146444 73896 146450 73908
rect 146938 73896 146944 73908
rect 146444 73868 146944 73896
rect 146444 73856 146450 73868
rect 146938 73856 146944 73868
rect 146996 73856 147002 73908
rect 188062 73856 188068 73908
rect 188120 73896 188126 73908
rect 269114 73896 269120 73908
rect 188120 73868 269120 73896
rect 188120 73856 188126 73868
rect 269114 73856 269120 73868
rect 269172 73856 269178 73908
rect 8938 73788 8944 73840
rect 8996 73828 9002 73840
rect 105814 73828 105820 73840
rect 8996 73800 105820 73828
rect 8996 73788 9002 73800
rect 105814 73788 105820 73800
rect 105872 73788 105878 73840
rect 106826 73788 106832 73840
rect 106884 73828 106890 73840
rect 131114 73828 131120 73840
rect 106884 73800 131120 73828
rect 106884 73788 106890 73800
rect 131114 73788 131120 73800
rect 131172 73788 131178 73840
rect 131206 73788 131212 73840
rect 131264 73828 131270 73840
rect 145098 73828 145104 73840
rect 131264 73800 145104 73828
rect 131264 73788 131270 73800
rect 145098 73788 145104 73800
rect 145156 73828 145162 73840
rect 145156 73800 147674 73828
rect 145156 73788 145162 73800
rect 111794 73720 111800 73772
rect 111852 73760 111858 73772
rect 140682 73760 140688 73772
rect 111852 73732 140688 73760
rect 111852 73720 111858 73732
rect 140682 73720 140688 73732
rect 140740 73720 140746 73772
rect 147646 73760 147674 73800
rect 175090 73788 175096 73840
rect 175148 73828 175154 73840
rect 189074 73828 189080 73840
rect 175148 73800 189080 73828
rect 175148 73788 175154 73800
rect 189074 73788 189080 73800
rect 189132 73788 189138 73840
rect 193766 73788 193772 73840
rect 193824 73828 193830 73840
rect 340874 73828 340880 73840
rect 193824 73800 340880 73828
rect 193824 73788 193830 73800
rect 340874 73788 340880 73800
rect 340932 73788 340938 73840
rect 152458 73760 152464 73772
rect 147646 73732 152464 73760
rect 152458 73720 152464 73732
rect 152516 73720 152522 73772
rect 170766 73720 170772 73772
rect 170824 73760 170830 73772
rect 196894 73760 196900 73772
rect 170824 73732 196900 73760
rect 170824 73720 170830 73732
rect 196894 73720 196900 73732
rect 196952 73720 196958 73772
rect 105814 73584 105820 73636
rect 105872 73624 105878 73636
rect 132402 73624 132408 73636
rect 105872 73596 132408 73624
rect 105872 73584 105878 73596
rect 132402 73584 132408 73596
rect 132460 73584 132466 73636
rect 145006 73584 145012 73636
rect 145064 73624 145070 73636
rect 145742 73624 145748 73636
rect 145064 73596 145748 73624
rect 145064 73584 145070 73596
rect 145742 73584 145748 73596
rect 145800 73584 145806 73636
rect 131298 73516 131304 73568
rect 131356 73556 131362 73568
rect 131666 73556 131672 73568
rect 131356 73528 131672 73556
rect 131356 73516 131362 73528
rect 131666 73516 131672 73528
rect 131724 73516 131730 73568
rect 135622 73516 135628 73568
rect 135680 73556 135686 73568
rect 136082 73556 136088 73568
rect 135680 73528 136088 73556
rect 135680 73516 135686 73528
rect 136082 73516 136088 73528
rect 136140 73516 136146 73568
rect 107654 73176 107660 73228
rect 107712 73216 107718 73228
rect 108758 73216 108764 73228
rect 107712 73188 108764 73216
rect 107712 73176 107718 73188
rect 108758 73176 108764 73188
rect 108816 73176 108822 73228
rect 142338 73176 142344 73228
rect 142396 73216 142402 73228
rect 144730 73216 144736 73228
rect 142396 73188 144736 73216
rect 142396 73176 142402 73188
rect 144730 73176 144736 73188
rect 144788 73216 144794 73228
rect 149698 73216 149704 73228
rect 144788 73188 149704 73216
rect 144788 73176 144794 73188
rect 149698 73176 149704 73188
rect 149756 73176 149762 73228
rect 97718 73108 97724 73160
rect 97776 73148 97782 73160
rect 151262 73148 151268 73160
rect 97776 73120 151268 73148
rect 97776 73108 97782 73120
rect 151262 73108 151268 73120
rect 151320 73108 151326 73160
rect 153746 73108 153752 73160
rect 153804 73148 153810 73160
rect 154390 73148 154396 73160
rect 153804 73120 154396 73148
rect 153804 73108 153810 73120
rect 154390 73108 154396 73120
rect 154448 73108 154454 73160
rect 155678 73108 155684 73160
rect 155736 73148 155742 73160
rect 216766 73148 216772 73160
rect 155736 73120 216772 73148
rect 155736 73108 155742 73120
rect 216766 73108 216772 73120
rect 216824 73108 216830 73160
rect 327718 73108 327724 73160
rect 327776 73148 327782 73160
rect 580166 73148 580172 73160
rect 327776 73120 580172 73148
rect 327776 73108 327782 73120
rect 580166 73108 580172 73120
rect 580224 73108 580230 73160
rect 122466 73040 122472 73092
rect 122524 73080 122530 73092
rect 151078 73080 151084 73092
rect 122524 73052 151084 73080
rect 122524 73040 122530 73052
rect 151078 73040 151084 73052
rect 151136 73080 151142 73092
rect 151446 73080 151452 73092
rect 151136 73052 151452 73080
rect 151136 73040 151142 73052
rect 151446 73040 151452 73052
rect 151504 73040 151510 73092
rect 161474 73040 161480 73092
rect 161532 73080 161538 73092
rect 162670 73080 162676 73092
rect 161532 73052 162676 73080
rect 161532 73040 161538 73052
rect 162670 73040 162676 73052
rect 162728 73040 162734 73092
rect 163222 73040 163228 73092
rect 163280 73080 163286 73092
rect 197998 73080 198004 73092
rect 163280 73052 198004 73080
rect 163280 73040 163286 73052
rect 197998 73040 198004 73052
rect 198056 73040 198062 73092
rect 98822 72972 98828 73024
rect 98880 73012 98886 73024
rect 133782 73012 133788 73024
rect 98880 72984 133788 73012
rect 98880 72972 98886 72984
rect 133782 72972 133788 72984
rect 133840 72972 133846 73024
rect 142338 72972 142344 73024
rect 142396 73012 142402 73024
rect 143166 73012 143172 73024
rect 142396 72984 143172 73012
rect 142396 72972 142402 72984
rect 143166 72972 143172 72984
rect 143224 72972 143230 73024
rect 153102 72972 153108 73024
rect 153160 73012 153166 73024
rect 186866 73012 186872 73024
rect 153160 72984 186872 73012
rect 153160 72972 153166 72984
rect 186866 72972 186872 72984
rect 186924 72972 186930 73024
rect 99006 72904 99012 72956
rect 99064 72944 99070 72956
rect 132954 72944 132960 72956
rect 99064 72916 132960 72944
rect 99064 72904 99070 72916
rect 132954 72904 132960 72916
rect 133012 72904 133018 72956
rect 157150 72904 157156 72956
rect 157208 72944 157214 72956
rect 191190 72944 191196 72956
rect 157208 72916 191196 72944
rect 157208 72904 157214 72916
rect 191190 72904 191196 72916
rect 191248 72944 191254 72956
rect 191742 72944 191748 72956
rect 191248 72916 191748 72944
rect 191248 72904 191254 72916
rect 191742 72904 191748 72916
rect 191800 72904 191806 72956
rect 96614 72836 96620 72888
rect 96672 72876 96678 72888
rect 105906 72876 105912 72888
rect 96672 72848 105912 72876
rect 96672 72836 96678 72848
rect 105906 72836 105912 72848
rect 105964 72876 105970 72888
rect 140038 72876 140044 72888
rect 105964 72848 140044 72876
rect 105964 72836 105970 72848
rect 140038 72836 140044 72848
rect 140096 72836 140102 72888
rect 161474 72836 161480 72888
rect 161532 72876 161538 72888
rect 162118 72876 162124 72888
rect 161532 72848 162124 72876
rect 161532 72836 161538 72848
rect 162118 72836 162124 72848
rect 162176 72836 162182 72888
rect 163222 72836 163228 72888
rect 163280 72876 163286 72888
rect 163866 72876 163872 72888
rect 163280 72848 163872 72876
rect 163280 72836 163286 72848
rect 163866 72836 163872 72848
rect 163924 72836 163930 72888
rect 169846 72836 169852 72888
rect 169904 72876 169910 72888
rect 171042 72876 171048 72888
rect 169904 72848 171048 72876
rect 169904 72836 169910 72848
rect 171042 72836 171048 72848
rect 171100 72876 171106 72888
rect 204622 72876 204628 72888
rect 171100 72848 204628 72876
rect 171100 72836 171106 72848
rect 204622 72836 204628 72848
rect 204680 72836 204686 72888
rect 216766 72836 216772 72888
rect 216824 72876 216830 72888
rect 220078 72876 220084 72888
rect 216824 72848 220084 72876
rect 216824 72836 216830 72848
rect 220078 72836 220084 72848
rect 220136 72836 220142 72888
rect 118602 72768 118608 72820
rect 118660 72808 118666 72820
rect 150986 72808 150992 72820
rect 118660 72780 150992 72808
rect 118660 72768 118666 72780
rect 150986 72768 150992 72780
rect 151044 72768 151050 72820
rect 162670 72768 162676 72820
rect 162728 72808 162734 72820
rect 181346 72808 181352 72820
rect 162728 72780 181352 72808
rect 162728 72768 162734 72780
rect 181346 72768 181352 72780
rect 181404 72768 181410 72820
rect 191742 72768 191748 72820
rect 191800 72808 191806 72820
rect 287698 72808 287704 72820
rect 191800 72780 287704 72808
rect 191800 72768 191806 72780
rect 287698 72768 287704 72780
rect 287756 72768 287762 72820
rect 114922 72700 114928 72752
rect 114980 72740 114986 72752
rect 147674 72740 147680 72752
rect 114980 72712 147680 72740
rect 114980 72700 114986 72712
rect 147674 72700 147680 72712
rect 147732 72740 147738 72752
rect 148870 72740 148876 72752
rect 147732 72712 148876 72740
rect 147732 72700 147738 72712
rect 148870 72700 148876 72712
rect 148928 72700 148934 72752
rect 154390 72700 154396 72752
rect 154448 72740 154454 72752
rect 187326 72740 187332 72752
rect 154448 72712 187332 72740
rect 154448 72700 154454 72712
rect 187326 72700 187332 72712
rect 187384 72700 187390 72752
rect 191650 72700 191656 72752
rect 191708 72740 191714 72752
rect 304994 72740 305000 72752
rect 191708 72712 305000 72740
rect 191708 72700 191714 72712
rect 304994 72700 305000 72712
rect 305052 72700 305058 72752
rect 109954 72632 109960 72684
rect 110012 72672 110018 72684
rect 142338 72672 142344 72684
rect 110012 72644 142344 72672
rect 110012 72632 110018 72644
rect 142338 72632 142344 72644
rect 142396 72632 142402 72684
rect 150986 72632 150992 72684
rect 151044 72672 151050 72684
rect 151630 72672 151636 72684
rect 151044 72644 151636 72672
rect 151044 72632 151050 72644
rect 151630 72632 151636 72644
rect 151688 72632 151694 72684
rect 157518 72632 157524 72684
rect 157576 72672 157582 72684
rect 192754 72672 192760 72684
rect 157576 72644 192760 72672
rect 157576 72632 157582 72644
rect 192754 72632 192760 72644
rect 192812 72672 192818 72684
rect 322934 72672 322940 72684
rect 192812 72644 322940 72672
rect 192812 72632 192818 72644
rect 322934 72632 322940 72644
rect 322992 72632 322998 72684
rect 108298 72564 108304 72616
rect 108356 72604 108362 72616
rect 138382 72604 138388 72616
rect 108356 72576 138388 72604
rect 108356 72564 108362 72576
rect 138382 72564 138388 72576
rect 138440 72564 138446 72616
rect 156782 72564 156788 72616
rect 156840 72604 156846 72616
rect 157058 72604 157064 72616
rect 156840 72576 157064 72604
rect 156840 72564 156846 72576
rect 157058 72564 157064 72576
rect 157116 72564 157122 72616
rect 157702 72564 157708 72616
rect 157760 72604 157766 72616
rect 192294 72604 192300 72616
rect 157760 72576 192300 72604
rect 157760 72564 157766 72576
rect 192294 72564 192300 72576
rect 192352 72604 192358 72616
rect 323578 72604 323584 72616
rect 192352 72576 323584 72604
rect 192352 72564 192358 72576
rect 323578 72564 323584 72576
rect 323636 72564 323642 72616
rect 21450 72496 21456 72548
rect 21508 72536 21514 72548
rect 98822 72536 98828 72548
rect 21508 72508 98828 72536
rect 21508 72496 21514 72508
rect 98822 72496 98828 72508
rect 98880 72496 98886 72548
rect 121086 72496 121092 72548
rect 121144 72536 121150 72548
rect 149790 72536 149796 72548
rect 121144 72508 149796 72536
rect 121144 72496 121150 72508
rect 149790 72496 149796 72508
rect 149848 72496 149854 72548
rect 159174 72496 159180 72548
rect 159232 72536 159238 72548
rect 194134 72536 194140 72548
rect 159232 72508 194140 72536
rect 159232 72496 159238 72508
rect 194134 72496 194140 72508
rect 194192 72536 194198 72548
rect 342898 72536 342904 72548
rect 194192 72508 342904 72536
rect 194192 72496 194198 72508
rect 342898 72496 342904 72508
rect 342956 72496 342962 72548
rect 9674 72428 9680 72480
rect 9732 72468 9738 72480
rect 98730 72468 98736 72480
rect 9732 72440 98736 72468
rect 9732 72428 9738 72440
rect 98730 72428 98736 72440
rect 98788 72428 98794 72480
rect 119062 72428 119068 72480
rect 119120 72468 119126 72480
rect 148134 72468 148140 72480
rect 119120 72440 148140 72468
rect 119120 72428 119126 72440
rect 148134 72428 148140 72440
rect 148192 72428 148198 72480
rect 161014 72428 161020 72480
rect 161072 72468 161078 72480
rect 191650 72468 191656 72480
rect 161072 72440 191656 72468
rect 161072 72428 161078 72440
rect 191650 72428 191656 72440
rect 191708 72428 191714 72480
rect 197998 72428 198004 72480
rect 198056 72468 198062 72480
rect 396718 72468 396724 72480
rect 198056 72440 396724 72468
rect 198056 72428 198062 72440
rect 396718 72428 396724 72440
rect 396776 72428 396782 72480
rect 110966 72360 110972 72412
rect 111024 72400 111030 72412
rect 138106 72400 138112 72412
rect 111024 72372 138112 72400
rect 111024 72360 111030 72372
rect 138106 72360 138112 72372
rect 138164 72400 138170 72412
rect 138934 72400 138940 72412
rect 138164 72372 138940 72400
rect 138164 72360 138170 72372
rect 138934 72360 138940 72372
rect 138992 72360 138998 72412
rect 180518 72400 180524 72412
rect 176626 72372 180524 72400
rect 121362 72292 121368 72344
rect 121420 72332 121426 72344
rect 129918 72332 129924 72344
rect 121420 72304 129924 72332
rect 121420 72292 121426 72304
rect 129918 72292 129924 72304
rect 129976 72332 129982 72344
rect 141510 72332 141516 72344
rect 129976 72304 141516 72332
rect 129976 72292 129982 72304
rect 141510 72292 141516 72304
rect 141568 72292 141574 72344
rect 170306 72292 170312 72344
rect 170364 72332 170370 72344
rect 176626 72332 176654 72372
rect 180518 72360 180524 72372
rect 180576 72400 180582 72412
rect 207106 72400 207112 72412
rect 180576 72372 207112 72400
rect 180576 72360 180582 72372
rect 207106 72360 207112 72372
rect 207164 72360 207170 72412
rect 170364 72304 176654 72332
rect 170364 72292 170370 72304
rect 98730 72224 98736 72276
rect 98788 72264 98794 72276
rect 128630 72264 128636 72276
rect 98788 72236 128636 72264
rect 98788 72224 98794 72236
rect 128630 72224 128636 72236
rect 128688 72224 128694 72276
rect 159910 72224 159916 72276
rect 159968 72264 159974 72276
rect 194226 72264 194232 72276
rect 159968 72236 194232 72264
rect 159968 72224 159974 72236
rect 194226 72224 194232 72236
rect 194284 72224 194290 72276
rect 132862 72020 132868 72072
rect 132920 72060 132926 72072
rect 133506 72060 133512 72072
rect 132920 72032 133512 72060
rect 132920 72020 132926 72032
rect 133506 72020 133512 72032
rect 133564 72020 133570 72072
rect 149790 71952 149796 72004
rect 149848 71992 149854 72004
rect 150250 71992 150256 72004
rect 149848 71964 150256 71992
rect 149848 71952 149854 71964
rect 150250 71952 150256 71964
rect 150308 71952 150314 72004
rect 3510 71680 3516 71732
rect 3568 71720 3574 71732
rect 13078 71720 13084 71732
rect 3568 71692 13084 71720
rect 3568 71680 3574 71692
rect 13078 71680 13084 71692
rect 13136 71680 13142 71732
rect 119706 71680 119712 71732
rect 119764 71720 119770 71732
rect 128446 71720 128452 71732
rect 119764 71692 128452 71720
rect 119764 71680 119770 71692
rect 128446 71680 128452 71692
rect 128504 71720 128510 71732
rect 129642 71720 129648 71732
rect 128504 71692 129648 71720
rect 128504 71680 128510 71692
rect 129642 71680 129648 71692
rect 129700 71680 129706 71732
rect 135346 71680 135352 71732
rect 135404 71720 135410 71732
rect 137462 71720 137468 71732
rect 135404 71692 137468 71720
rect 135404 71680 135410 71692
rect 137462 71680 137468 71692
rect 137520 71680 137526 71732
rect 142430 71680 142436 71732
rect 142488 71720 142494 71732
rect 142982 71720 142988 71732
rect 142488 71692 142988 71720
rect 142488 71680 142494 71692
rect 142982 71680 142988 71692
rect 143040 71680 143046 71732
rect 144086 71680 144092 71732
rect 144144 71720 144150 71732
rect 146294 71720 146300 71732
rect 144144 71692 146300 71720
rect 144144 71680 144150 71692
rect 146294 71680 146300 71692
rect 146352 71680 146358 71732
rect 149330 71680 149336 71732
rect 149388 71720 149394 71732
rect 150158 71720 150164 71732
rect 149388 71692 150164 71720
rect 149388 71680 149394 71692
rect 150158 71680 150164 71692
rect 150216 71680 150222 71732
rect 150710 71680 150716 71732
rect 150768 71720 150774 71732
rect 151446 71720 151452 71732
rect 150768 71692 151452 71720
rect 150768 71680 150774 71692
rect 151446 71680 151452 71692
rect 151504 71680 151510 71732
rect 157978 71680 157984 71732
rect 158036 71720 158042 71732
rect 158530 71720 158536 71732
rect 158036 71692 158536 71720
rect 158036 71680 158042 71692
rect 158530 71680 158536 71692
rect 158588 71680 158594 71732
rect 159358 71680 159364 71732
rect 159416 71720 159422 71732
rect 159542 71720 159548 71732
rect 159416 71692 159548 71720
rect 159416 71680 159422 71692
rect 159542 71680 159548 71692
rect 159600 71680 159606 71732
rect 164234 71680 164240 71732
rect 164292 71720 164298 71732
rect 165062 71720 165068 71732
rect 164292 71692 165068 71720
rect 164292 71680 164298 71692
rect 165062 71680 165068 71692
rect 165120 71680 165126 71732
rect 165522 71680 165528 71732
rect 165580 71720 165586 71732
rect 206186 71720 206192 71732
rect 165580 71692 206192 71720
rect 165580 71680 165586 71692
rect 206186 71680 206192 71692
rect 206244 71680 206250 71732
rect 105722 71612 105728 71664
rect 105780 71652 105786 71664
rect 139762 71652 139768 71664
rect 105780 71624 139768 71652
rect 105780 71612 105786 71624
rect 139762 71612 139768 71624
rect 139820 71612 139826 71664
rect 140774 71612 140780 71664
rect 140832 71652 140838 71664
rect 143350 71652 143356 71664
rect 140832 71624 143356 71652
rect 140832 71612 140838 71624
rect 143350 71612 143356 71624
rect 143408 71612 143414 71664
rect 157334 71612 157340 71664
rect 157392 71652 157398 71664
rect 158254 71652 158260 71664
rect 157392 71624 158260 71652
rect 157392 71612 157398 71624
rect 158254 71612 158260 71624
rect 158312 71612 158318 71664
rect 159560 71652 159588 71680
rect 159560 71624 165016 71652
rect 118050 71544 118056 71596
rect 118108 71584 118114 71596
rect 149330 71584 149336 71596
rect 118108 71556 149336 71584
rect 118108 71544 118114 71556
rect 149330 71544 149336 71556
rect 149388 71544 149394 71596
rect 150434 71544 150440 71596
rect 150492 71584 150498 71596
rect 151538 71584 151544 71596
rect 150492 71556 151544 71584
rect 150492 71544 150498 71556
rect 151538 71544 151544 71556
rect 151596 71544 151602 71596
rect 157610 71544 157616 71596
rect 157668 71584 157674 71596
rect 158438 71584 158444 71596
rect 157668 71556 158444 71584
rect 157668 71544 157674 71556
rect 158438 71544 158444 71556
rect 158496 71544 158502 71596
rect 164234 71544 164240 71596
rect 164292 71584 164298 71596
rect 164878 71584 164884 71596
rect 164292 71556 164884 71584
rect 164292 71544 164298 71556
rect 164878 71544 164884 71556
rect 164936 71544 164942 71596
rect 164988 71584 165016 71624
rect 166810 71612 166816 71664
rect 166868 71652 166874 71664
rect 207382 71652 207388 71664
rect 166868 71624 207388 71652
rect 166868 71612 166874 71624
rect 207382 71612 207388 71624
rect 207440 71612 207446 71664
rect 193950 71584 193956 71596
rect 164988 71556 193956 71584
rect 193950 71544 193956 71556
rect 194008 71544 194014 71596
rect 104250 71476 104256 71528
rect 104308 71516 104314 71528
rect 104526 71516 104532 71528
rect 104308 71488 104532 71516
rect 104308 71476 104314 71488
rect 104526 71476 104532 71488
rect 104584 71516 104590 71528
rect 135346 71516 135352 71528
rect 104584 71488 135352 71516
rect 104584 71476 104590 71488
rect 135346 71476 135352 71488
rect 135404 71476 135410 71528
rect 149146 71476 149152 71528
rect 149204 71516 149210 71528
rect 150158 71516 150164 71528
rect 149204 71488 150164 71516
rect 149204 71476 149210 71488
rect 150158 71476 150164 71488
rect 150216 71476 150222 71528
rect 157334 71476 157340 71528
rect 157392 71516 157398 71528
rect 157886 71516 157892 71528
rect 157392 71488 157892 71516
rect 157392 71476 157398 71488
rect 157886 71476 157892 71488
rect 157944 71476 157950 71528
rect 158346 71476 158352 71528
rect 158404 71516 158410 71528
rect 192570 71516 192576 71528
rect 158404 71488 192576 71516
rect 158404 71476 158410 71488
rect 192570 71476 192576 71488
rect 192628 71476 192634 71528
rect 105998 71448 106004 71460
rect 103486 71420 106004 71448
rect 84838 71068 84844 71120
rect 84896 71108 84902 71120
rect 103486 71108 103514 71420
rect 105998 71408 106004 71420
rect 106056 71448 106062 71460
rect 138198 71448 138204 71460
rect 106056 71420 138204 71448
rect 106056 71408 106062 71420
rect 138198 71408 138204 71420
rect 138256 71408 138262 71460
rect 162486 71408 162492 71460
rect 162544 71448 162550 71460
rect 197078 71448 197084 71460
rect 162544 71420 197084 71448
rect 162544 71408 162550 71420
rect 197078 71408 197084 71420
rect 197136 71408 197142 71460
rect 120902 71340 120908 71392
rect 120960 71380 120966 71392
rect 151998 71380 152004 71392
rect 120960 71352 152004 71380
rect 120960 71340 120966 71352
rect 151998 71340 152004 71352
rect 152056 71340 152062 71392
rect 158438 71340 158444 71392
rect 158496 71380 158502 71392
rect 192478 71380 192484 71392
rect 158496 71352 192484 71380
rect 158496 71340 158502 71352
rect 192478 71340 192484 71352
rect 192536 71340 192542 71392
rect 117590 71272 117596 71324
rect 117648 71312 117654 71324
rect 149422 71312 149428 71324
rect 117648 71284 149428 71312
rect 117648 71272 117654 71284
rect 149422 71272 149428 71284
rect 149480 71272 149486 71324
rect 165062 71272 165068 71324
rect 165120 71312 165126 71324
rect 199194 71312 199200 71324
rect 165120 71284 199200 71312
rect 165120 71272 165126 71284
rect 199194 71272 199200 71284
rect 199252 71272 199258 71324
rect 112530 71204 112536 71256
rect 112588 71244 112594 71256
rect 142430 71244 142436 71256
rect 112588 71216 142436 71244
rect 112588 71204 112594 71216
rect 142430 71204 142436 71216
rect 142488 71204 142494 71256
rect 158254 71204 158260 71256
rect 158312 71244 158318 71256
rect 191006 71244 191012 71256
rect 158312 71216 191012 71244
rect 158312 71204 158318 71216
rect 191006 71204 191012 71216
rect 191064 71204 191070 71256
rect 135254 71136 135260 71188
rect 135312 71176 135318 71188
rect 135714 71176 135720 71188
rect 135312 71148 135720 71176
rect 135312 71136 135318 71148
rect 135714 71136 135720 71148
rect 135772 71136 135778 71188
rect 146570 71136 146576 71188
rect 146628 71176 146634 71188
rect 181438 71176 181444 71188
rect 146628 71148 181444 71176
rect 146628 71136 146634 71148
rect 181438 71136 181444 71148
rect 181496 71136 181502 71188
rect 181806 71136 181812 71188
rect 181864 71176 181870 71188
rect 203242 71176 203248 71188
rect 181864 71148 203248 71176
rect 181864 71136 181870 71148
rect 203242 71136 203248 71148
rect 203300 71136 203306 71188
rect 84896 71080 103514 71108
rect 84896 71068 84902 71080
rect 114370 71068 114376 71120
rect 114428 71108 114434 71120
rect 128354 71108 128360 71120
rect 114428 71080 128360 71108
rect 114428 71068 114434 71080
rect 128354 71068 128360 71080
rect 128412 71108 128418 71120
rect 141234 71108 141240 71120
rect 128412 71080 141240 71108
rect 128412 71068 128418 71080
rect 141234 71068 141240 71080
rect 141292 71068 141298 71120
rect 147122 71068 147128 71120
rect 147180 71108 147186 71120
rect 184290 71108 184296 71120
rect 147180 71080 184296 71108
rect 147180 71068 147186 71080
rect 184290 71068 184296 71080
rect 184348 71068 184354 71120
rect 71774 71000 71780 71052
rect 71832 71040 71838 71052
rect 104250 71040 104256 71052
rect 71832 71012 104256 71040
rect 71832 71000 71838 71012
rect 104250 71000 104256 71012
rect 104308 71000 104314 71052
rect 110782 71000 110788 71052
rect 110840 71040 110846 71052
rect 140774 71040 140780 71052
rect 110840 71012 140780 71040
rect 110840 71000 110846 71012
rect 140774 71000 140780 71012
rect 140832 71000 140838 71052
rect 148870 71000 148876 71052
rect 148928 71040 148934 71052
rect 200850 71040 200856 71052
rect 148928 71012 200856 71040
rect 148928 71000 148934 71012
rect 200850 71000 200856 71012
rect 200908 71000 200914 71052
rect 121546 70932 121552 70984
rect 121604 70972 121610 70984
rect 151446 70972 151452 70984
rect 121604 70944 151452 70972
rect 121604 70932 121610 70944
rect 151446 70932 151452 70944
rect 151504 70932 151510 70984
rect 156322 70932 156328 70984
rect 156380 70972 156386 70984
rect 157242 70972 157248 70984
rect 156380 70944 157248 70972
rect 156380 70932 156386 70944
rect 157242 70932 157248 70944
rect 157300 70972 157306 70984
rect 187694 70972 187700 70984
rect 157300 70944 187700 70972
rect 157300 70932 157306 70944
rect 187694 70932 187700 70944
rect 187752 70932 187758 70984
rect 117222 70864 117228 70916
rect 117280 70904 117286 70916
rect 140958 70904 140964 70916
rect 117280 70876 140964 70904
rect 117280 70864 117286 70876
rect 140958 70864 140964 70876
rect 141016 70864 141022 70916
rect 151998 70864 152004 70916
rect 152056 70904 152062 70916
rect 152918 70904 152924 70916
rect 152056 70876 152924 70904
rect 152056 70864 152062 70876
rect 152918 70864 152924 70876
rect 152976 70864 152982 70916
rect 158530 70864 158536 70916
rect 158588 70904 158594 70916
rect 188246 70904 188252 70916
rect 158588 70876 188252 70904
rect 158588 70864 158594 70876
rect 188246 70864 188252 70876
rect 188304 70864 188310 70916
rect 114830 70796 114836 70848
rect 114888 70836 114894 70848
rect 149146 70836 149152 70848
rect 114888 70808 149152 70836
rect 114888 70796 114894 70808
rect 149146 70796 149152 70808
rect 149204 70796 149210 70848
rect 150434 70836 150440 70848
rect 149348 70808 150440 70836
rect 121638 70728 121644 70780
rect 121696 70768 121702 70780
rect 149348 70768 149376 70808
rect 150434 70796 150440 70808
rect 150492 70796 150498 70848
rect 158622 70796 158628 70848
rect 158680 70836 158686 70848
rect 187050 70836 187056 70848
rect 158680 70808 187056 70836
rect 158680 70796 158686 70808
rect 187050 70796 187056 70808
rect 187108 70796 187114 70848
rect 121696 70740 149376 70768
rect 121696 70728 121702 70740
rect 149422 70728 149428 70780
rect 149480 70768 149486 70780
rect 150066 70768 150072 70780
rect 149480 70740 150072 70768
rect 149480 70728 149486 70740
rect 150066 70728 150072 70740
rect 150124 70728 150130 70780
rect 167362 70728 167368 70780
rect 167420 70768 167426 70780
rect 167730 70768 167736 70780
rect 167420 70740 167736 70768
rect 167420 70728 167426 70740
rect 167730 70728 167736 70740
rect 167788 70728 167794 70780
rect 171226 70728 171232 70780
rect 171284 70768 171290 70780
rect 171962 70768 171968 70780
rect 171284 70740 171968 70768
rect 171284 70728 171290 70740
rect 171962 70728 171968 70740
rect 172020 70728 172026 70780
rect 174998 70728 175004 70780
rect 175056 70768 175062 70780
rect 175182 70768 175188 70780
rect 175056 70740 175188 70768
rect 175056 70728 175062 70740
rect 175182 70728 175188 70740
rect 175240 70728 175246 70780
rect 103514 70388 103520 70440
rect 103572 70428 103578 70440
rect 105722 70428 105728 70440
rect 103572 70400 105728 70428
rect 103572 70388 103578 70400
rect 105722 70388 105728 70400
rect 105780 70388 105786 70440
rect 100110 70320 100116 70372
rect 100168 70360 100174 70372
rect 134334 70360 134340 70372
rect 100168 70332 134340 70360
rect 100168 70320 100174 70332
rect 134334 70320 134340 70332
rect 134392 70320 134398 70372
rect 165338 70320 165344 70372
rect 165396 70360 165402 70372
rect 205726 70360 205732 70372
rect 165396 70332 205732 70360
rect 165396 70320 165402 70332
rect 205726 70320 205732 70332
rect 205784 70320 205790 70372
rect 209130 70320 209136 70372
rect 209188 70360 209194 70372
rect 210418 70360 210424 70372
rect 209188 70332 210424 70360
rect 209188 70320 209194 70332
rect 210418 70320 210424 70332
rect 210476 70320 210482 70372
rect 100754 70252 100760 70304
rect 100812 70292 100818 70304
rect 101306 70292 101312 70304
rect 100812 70264 101312 70292
rect 100812 70252 100818 70264
rect 101306 70252 101312 70264
rect 101364 70292 101370 70304
rect 135990 70292 135996 70304
rect 101364 70264 135996 70292
rect 101364 70252 101370 70264
rect 135990 70252 135996 70264
rect 136048 70252 136054 70304
rect 162394 70252 162400 70304
rect 162452 70292 162458 70304
rect 196618 70292 196624 70304
rect 162452 70264 196624 70292
rect 162452 70252 162458 70264
rect 196618 70252 196624 70264
rect 196676 70252 196682 70304
rect 104618 70184 104624 70236
rect 104676 70224 104682 70236
rect 138750 70224 138756 70236
rect 104676 70196 138756 70224
rect 104676 70184 104682 70196
rect 138750 70184 138756 70196
rect 138808 70184 138814 70236
rect 163866 70184 163872 70236
rect 163924 70224 163930 70236
rect 198274 70224 198280 70236
rect 163924 70196 198280 70224
rect 163924 70184 163930 70196
rect 198274 70184 198280 70196
rect 198332 70184 198338 70236
rect 97902 70116 97908 70168
rect 97960 70156 97966 70168
rect 115934 70156 115940 70168
rect 97960 70128 115940 70156
rect 97960 70116 97966 70128
rect 115934 70116 115940 70128
rect 115992 70156 115998 70168
rect 117222 70156 117228 70168
rect 115992 70128 117228 70156
rect 115992 70116 115998 70128
rect 117222 70116 117228 70128
rect 117280 70116 117286 70168
rect 117682 70116 117688 70168
rect 117740 70156 117746 70168
rect 151354 70156 151360 70168
rect 117740 70128 151360 70156
rect 117740 70116 117746 70128
rect 151354 70116 151360 70128
rect 151412 70116 151418 70168
rect 162578 70116 162584 70168
rect 162636 70156 162642 70168
rect 197170 70156 197176 70168
rect 162636 70128 197176 70156
rect 162636 70116 162642 70128
rect 197170 70116 197176 70128
rect 197228 70116 197234 70168
rect 118786 70048 118792 70100
rect 118844 70088 118850 70100
rect 151814 70088 151820 70100
rect 118844 70060 151820 70088
rect 118844 70048 118850 70060
rect 151814 70048 151820 70060
rect 151872 70048 151878 70100
rect 171226 70048 171232 70100
rect 171284 70088 171290 70100
rect 172146 70088 172152 70100
rect 171284 70060 172152 70088
rect 171284 70048 171290 70060
rect 172146 70048 172152 70060
rect 172204 70088 172210 70100
rect 205634 70088 205640 70100
rect 172204 70060 205640 70088
rect 172204 70048 172210 70060
rect 205634 70048 205640 70060
rect 205692 70048 205698 70100
rect 107378 69980 107384 70032
rect 107436 70020 107442 70032
rect 140130 70020 140136 70032
rect 107436 69992 140136 70020
rect 107436 69980 107442 69992
rect 140130 69980 140136 69992
rect 140188 69980 140194 70032
rect 161750 69980 161756 70032
rect 161808 70020 161814 70032
rect 162394 70020 162400 70032
rect 161808 69992 162400 70020
rect 161808 69980 161814 69992
rect 162394 69980 162400 69992
rect 162452 69980 162458 70032
rect 164694 69980 164700 70032
rect 164752 70020 164758 70032
rect 165338 70020 165344 70032
rect 164752 69992 165344 70020
rect 164752 69980 164758 69992
rect 165338 69980 165344 69992
rect 165396 69980 165402 70032
rect 169018 69980 169024 70032
rect 169076 70020 169082 70032
rect 169478 70020 169484 70032
rect 169076 69992 169484 70020
rect 169076 69980 169082 69992
rect 169478 69980 169484 69992
rect 169536 70020 169542 70032
rect 203426 70020 203432 70032
rect 169536 69992 203432 70020
rect 169536 69980 169542 69992
rect 203426 69980 203432 69992
rect 203484 69980 203490 70032
rect 102134 69912 102140 69964
rect 102192 69952 102198 69964
rect 102962 69952 102968 69964
rect 102192 69924 102968 69952
rect 102192 69912 102198 69924
rect 102962 69912 102968 69924
rect 103020 69952 103026 69964
rect 134886 69952 134892 69964
rect 103020 69924 134892 69952
rect 103020 69912 103026 69924
rect 134886 69912 134892 69924
rect 134944 69912 134950 69964
rect 161934 69912 161940 69964
rect 161992 69952 161998 69964
rect 162578 69952 162584 69964
rect 161992 69924 162584 69952
rect 161992 69912 161998 69924
rect 162578 69912 162584 69924
rect 162636 69912 162642 69964
rect 163130 69912 163136 69964
rect 163188 69952 163194 69964
rect 163866 69952 163872 69964
rect 163188 69924 163872 69952
rect 163188 69912 163194 69924
rect 163866 69912 163872 69924
rect 163924 69912 163930 69964
rect 164786 69912 164792 69964
rect 164844 69952 164850 69964
rect 165522 69952 165528 69964
rect 164844 69924 165528 69952
rect 164844 69912 164850 69924
rect 165522 69912 165528 69924
rect 165580 69952 165586 69964
rect 199746 69952 199752 69964
rect 165580 69924 199752 69952
rect 165580 69912 165586 69924
rect 199746 69912 199752 69924
rect 199804 69912 199810 69964
rect 112162 69844 112168 69896
rect 112220 69884 112226 69896
rect 143534 69884 143540 69896
rect 112220 69856 143540 69884
rect 112220 69844 112226 69856
rect 143534 69844 143540 69856
rect 143592 69884 143598 69896
rect 144454 69884 144460 69896
rect 143592 69856 144460 69884
rect 143592 69844 143598 69856
rect 144454 69844 144460 69856
rect 144512 69844 144518 69896
rect 159082 69844 159088 69896
rect 159140 69884 159146 69896
rect 159910 69884 159916 69896
rect 159140 69856 159916 69884
rect 159140 69844 159146 69856
rect 159910 69844 159916 69856
rect 159968 69884 159974 69896
rect 191374 69884 191380 69896
rect 159968 69856 191380 69884
rect 159968 69844 159974 69856
rect 191374 69844 191380 69856
rect 191432 69844 191438 69896
rect 85666 69776 85672 69828
rect 85724 69816 85730 69828
rect 104618 69816 104624 69828
rect 85724 69788 104624 69816
rect 85724 69776 85730 69788
rect 104618 69776 104624 69788
rect 104676 69776 104682 69828
rect 112070 69776 112076 69828
rect 112128 69816 112134 69828
rect 142522 69816 142528 69828
rect 112128 69788 142528 69816
rect 112128 69776 112134 69788
rect 142522 69776 142528 69788
rect 142580 69816 142586 69828
rect 143074 69816 143080 69828
rect 142580 69788 143080 69816
rect 142580 69776 142586 69788
rect 143074 69776 143080 69788
rect 143132 69776 143138 69828
rect 154482 69776 154488 69828
rect 154540 69816 154546 69828
rect 184474 69816 184480 69828
rect 154540 69788 184480 69816
rect 154540 69776 154546 69788
rect 184474 69776 184480 69788
rect 184532 69776 184538 69828
rect 45554 69708 45560 69760
rect 45612 69748 45618 69760
rect 100754 69748 100760 69760
rect 45612 69720 100760 69748
rect 45612 69708 45618 69720
rect 100754 69708 100760 69720
rect 100812 69708 100818 69760
rect 102778 69708 102784 69760
rect 102836 69748 102842 69760
rect 107378 69748 107384 69760
rect 102836 69720 107384 69748
rect 102836 69708 102842 69720
rect 107378 69708 107384 69720
rect 107436 69708 107442 69760
rect 113082 69708 113088 69760
rect 113140 69748 113146 69760
rect 139394 69748 139400 69760
rect 113140 69720 139400 69748
rect 113140 69708 113146 69720
rect 139394 69708 139400 69720
rect 139452 69708 139458 69760
rect 158990 69708 158996 69760
rect 159048 69748 159054 69760
rect 159634 69748 159640 69760
rect 159048 69720 159640 69748
rect 159048 69708 159054 69720
rect 159634 69708 159640 69720
rect 159692 69748 159698 69760
rect 189626 69748 189632 69760
rect 159692 69720 189632 69748
rect 159692 69708 159698 69720
rect 189626 69708 189632 69720
rect 189684 69708 189690 69760
rect 201678 69708 201684 69760
rect 201736 69748 201742 69760
rect 201862 69748 201868 69760
rect 201736 69720 201868 69748
rect 201736 69708 201742 69720
rect 201862 69708 201868 69720
rect 201920 69708 201926 69760
rect 35158 69640 35164 69692
rect 35216 69680 35222 69692
rect 102134 69680 102140 69692
rect 35216 69652 102140 69680
rect 35216 69640 35222 69652
rect 102134 69640 102140 69652
rect 102192 69640 102198 69692
rect 147582 69640 147588 69692
rect 147640 69680 147646 69692
rect 183554 69680 183560 69692
rect 147640 69652 183560 69680
rect 147640 69640 147646 69652
rect 183554 69640 183560 69652
rect 183612 69640 183618 69692
rect 210510 69680 210516 69692
rect 200086 69652 210516 69680
rect 153562 69572 153568 69624
rect 153620 69612 153626 69624
rect 154482 69612 154488 69624
rect 153620 69584 154488 69612
rect 153620 69572 153626 69584
rect 154482 69572 154488 69584
rect 154540 69572 154546 69624
rect 160462 69572 160468 69624
rect 160520 69612 160526 69624
rect 161106 69612 161112 69624
rect 160520 69584 161112 69612
rect 160520 69572 160526 69584
rect 161106 69572 161112 69584
rect 161164 69612 161170 69624
rect 188154 69612 188160 69624
rect 161164 69584 188160 69612
rect 161164 69572 161170 69584
rect 188154 69572 188160 69584
rect 188212 69572 188218 69624
rect 162302 69504 162308 69556
rect 162360 69544 162366 69556
rect 185394 69544 185400 69556
rect 162360 69516 185400 69544
rect 162360 69504 162366 69516
rect 185394 69504 185400 69516
rect 185452 69504 185458 69556
rect 180150 69436 180156 69488
rect 180208 69476 180214 69488
rect 197262 69476 197268 69488
rect 180208 69448 197268 69476
rect 180208 69436 180214 69448
rect 197262 69436 197268 69448
rect 197320 69476 197326 69488
rect 200086 69476 200114 69652
rect 210510 69640 210516 69652
rect 210568 69640 210574 69692
rect 197320 69448 200114 69476
rect 197320 69436 197326 69448
rect 151814 69028 151820 69080
rect 151872 69068 151878 69080
rect 152550 69068 152556 69080
rect 151872 69040 152556 69068
rect 151872 69028 151878 69040
rect 152550 69028 152556 69040
rect 152608 69028 152614 69080
rect 185394 69028 185400 69080
rect 185452 69068 185458 69080
rect 354674 69068 354680 69080
rect 185452 69040 354680 69068
rect 185452 69028 185458 69040
rect 354674 69028 354680 69040
rect 354732 69028 354738 69080
rect 107562 68960 107568 69012
rect 107620 69000 107626 69012
rect 114554 69000 114560 69012
rect 107620 68972 114560 69000
rect 107620 68960 107626 68972
rect 114554 68960 114560 68972
rect 114612 68960 114618 69012
rect 117976 68972 138014 69000
rect 110322 68892 110328 68944
rect 110380 68932 110386 68944
rect 117976 68932 118004 68972
rect 132034 68932 132040 68944
rect 110380 68904 118004 68932
rect 118068 68904 132040 68932
rect 110380 68892 110386 68904
rect 110138 68824 110144 68876
rect 110196 68864 110202 68876
rect 118068 68864 118096 68904
rect 132034 68892 132040 68904
rect 132092 68892 132098 68944
rect 137986 68932 138014 68972
rect 141510 68960 141516 69012
rect 141568 69000 141574 69012
rect 142154 69000 142160 69012
rect 141568 68972 142160 69000
rect 141568 68960 141574 68972
rect 142154 68960 142160 68972
rect 142212 68960 142218 69012
rect 158898 68960 158904 69012
rect 158956 69000 158962 69012
rect 159726 69000 159732 69012
rect 158956 68972 159732 69000
rect 158956 68960 158962 68972
rect 159726 68960 159732 68972
rect 159784 69000 159790 69012
rect 207290 69000 207296 69012
rect 159784 68972 207296 69000
rect 159784 68960 159790 68972
rect 207290 68960 207296 68972
rect 207348 68960 207354 69012
rect 143994 68932 144000 68944
rect 137986 68904 144000 68932
rect 143994 68892 144000 68904
rect 144052 68932 144058 68944
rect 144454 68932 144460 68944
rect 144052 68904 144460 68932
rect 144052 68892 144058 68904
rect 144454 68892 144460 68904
rect 144512 68892 144518 68944
rect 166074 68892 166080 68944
rect 166132 68932 166138 68944
rect 166810 68932 166816 68944
rect 166132 68904 166816 68932
rect 166132 68892 166138 68904
rect 166810 68892 166816 68904
rect 166868 68892 166874 68944
rect 177574 68892 177580 68944
rect 177632 68932 177638 68944
rect 212810 68932 212816 68944
rect 177632 68904 212816 68932
rect 177632 68892 177638 68904
rect 212810 68892 212816 68904
rect 212868 68932 212874 68944
rect 213822 68932 213828 68944
rect 212868 68904 213828 68932
rect 212868 68892 212874 68904
rect 213822 68892 213828 68904
rect 213880 68892 213886 68944
rect 110196 68836 118096 68864
rect 110196 68824 110202 68836
rect 121730 68824 121736 68876
rect 121788 68864 121794 68876
rect 132218 68864 132224 68876
rect 121788 68836 132224 68864
rect 121788 68824 121794 68836
rect 132218 68824 132224 68836
rect 132276 68824 132282 68876
rect 132402 68824 132408 68876
rect 132460 68864 132466 68876
rect 156046 68864 156052 68876
rect 132460 68836 156052 68864
rect 132460 68824 132466 68836
rect 156046 68824 156052 68836
rect 156104 68824 156110 68876
rect 165982 68824 165988 68876
rect 166040 68864 166046 68876
rect 166902 68864 166908 68876
rect 166040 68836 166908 68864
rect 166040 68824 166046 68836
rect 166902 68824 166908 68836
rect 166960 68824 166966 68876
rect 166994 68824 167000 68876
rect 167052 68864 167058 68876
rect 167914 68864 167920 68876
rect 167052 68836 167920 68864
rect 167052 68824 167058 68836
rect 167914 68824 167920 68836
rect 167972 68864 167978 68876
rect 202046 68864 202052 68876
rect 167972 68836 202052 68864
rect 167972 68824 167978 68836
rect 202046 68824 202052 68836
rect 202104 68824 202110 68876
rect 101582 68796 101588 68808
rect 84166 68768 101588 68796
rect 48314 68416 48320 68468
rect 48372 68456 48378 68468
rect 84166 68456 84194 68768
rect 101582 68756 101588 68768
rect 101640 68796 101646 68808
rect 131942 68796 131948 68808
rect 101640 68768 131948 68796
rect 101640 68756 101646 68768
rect 131942 68756 131948 68768
rect 132000 68756 132006 68808
rect 132034 68756 132040 68808
rect 132092 68796 132098 68808
rect 144270 68796 144276 68808
rect 132092 68768 144276 68796
rect 132092 68756 132098 68768
rect 144270 68756 144276 68768
rect 144328 68796 144334 68808
rect 144546 68796 144552 68808
rect 144328 68768 144552 68796
rect 144328 68756 144334 68768
rect 144546 68756 144552 68768
rect 144604 68756 144610 68808
rect 167086 68756 167092 68808
rect 167144 68796 167150 68808
rect 168006 68796 168012 68808
rect 167144 68768 168012 68796
rect 167144 68756 167150 68768
rect 168006 68756 168012 68768
rect 168064 68796 168070 68808
rect 201954 68796 201960 68808
rect 168064 68768 201960 68796
rect 168064 68756 168070 68768
rect 201954 68756 201960 68768
rect 202012 68756 202018 68808
rect 108850 68688 108856 68740
rect 108908 68728 108914 68740
rect 142706 68728 142712 68740
rect 108908 68700 142712 68728
rect 108908 68688 108914 68700
rect 142706 68688 142712 68700
rect 142764 68688 142770 68740
rect 166902 68688 166908 68740
rect 166960 68728 166966 68740
rect 200758 68728 200764 68740
rect 166960 68700 200764 68728
rect 166960 68688 166966 68700
rect 200758 68688 200764 68700
rect 200816 68688 200822 68740
rect 134426 68660 134432 68672
rect 48372 68428 84194 68456
rect 103486 68632 134432 68660
rect 48372 68416 48378 68428
rect 26234 68348 26240 68400
rect 26292 68388 26298 68400
rect 101674 68388 101680 68400
rect 26292 68360 101680 68388
rect 26292 68348 26298 68360
rect 101674 68348 101680 68360
rect 101732 68388 101738 68400
rect 103486 68388 103514 68632
rect 134426 68620 134432 68632
rect 134484 68620 134490 68672
rect 142154 68620 142160 68672
rect 142212 68660 142218 68672
rect 142338 68660 142344 68672
rect 142212 68632 142344 68660
rect 142212 68620 142218 68632
rect 142338 68620 142344 68632
rect 142396 68620 142402 68672
rect 153286 68620 153292 68672
rect 153344 68660 153350 68672
rect 154298 68660 154304 68672
rect 153344 68632 154304 68660
rect 153344 68620 153350 68632
rect 154298 68620 154304 68632
rect 154356 68620 154362 68672
rect 166810 68620 166816 68672
rect 166868 68660 166874 68672
rect 200666 68660 200672 68672
rect 166868 68632 200672 68660
rect 166868 68620 166874 68632
rect 200666 68620 200672 68632
rect 200724 68620 200730 68672
rect 106918 68552 106924 68604
rect 106976 68592 106982 68604
rect 109770 68592 109776 68604
rect 106976 68564 109776 68592
rect 106976 68552 106982 68564
rect 109770 68552 109776 68564
rect 109828 68592 109834 68604
rect 139670 68592 139676 68604
rect 109828 68564 139676 68592
rect 109828 68552 109834 68564
rect 139670 68552 139676 68564
rect 139728 68552 139734 68604
rect 169846 68552 169852 68604
rect 169904 68592 169910 68604
rect 170950 68592 170956 68604
rect 169904 68564 170956 68592
rect 169904 68552 169910 68564
rect 170950 68552 170956 68564
rect 171008 68592 171014 68604
rect 204438 68592 204444 68604
rect 171008 68564 204444 68592
rect 171008 68552 171014 68564
rect 204438 68552 204444 68564
rect 204496 68552 204502 68604
rect 133598 68524 133604 68536
rect 101732 68360 103514 68388
rect 113146 68496 133604 68524
rect 101732 68348 101738 68360
rect 18598 68280 18604 68332
rect 18656 68320 18662 68332
rect 101766 68320 101772 68332
rect 18656 68292 101772 68320
rect 18656 68280 18662 68292
rect 101766 68280 101772 68292
rect 101824 68320 101830 68332
rect 113146 68320 113174 68496
rect 133598 68484 133604 68496
rect 133656 68484 133662 68536
rect 142430 68484 142436 68536
rect 142488 68484 142494 68536
rect 186314 68484 186320 68536
rect 186372 68524 186378 68536
rect 186682 68524 186688 68536
rect 186372 68496 186688 68524
rect 186372 68484 186378 68496
rect 186682 68484 186688 68496
rect 186740 68524 186746 68536
rect 252554 68524 252560 68536
rect 186740 68496 252560 68524
rect 186740 68484 186746 68496
rect 252554 68484 252560 68496
rect 252612 68484 252618 68536
rect 131942 68416 131948 68468
rect 132000 68456 132006 68468
rect 135622 68456 135628 68468
rect 132000 68428 135628 68456
rect 132000 68416 132006 68428
rect 135622 68416 135628 68428
rect 135680 68416 135686 68468
rect 101824 68292 113174 68320
rect 101824 68280 101830 68292
rect 142448 68264 142476 68484
rect 166166 68416 166172 68468
rect 166224 68456 166230 68468
rect 200574 68456 200580 68468
rect 166224 68428 200580 68456
rect 166224 68416 166230 68428
rect 200574 68416 200580 68428
rect 200632 68456 200638 68468
rect 427814 68456 427820 68468
rect 200632 68428 427820 68456
rect 200632 68416 200638 68428
rect 427814 68416 427820 68428
rect 427872 68416 427878 68468
rect 164602 68348 164608 68400
rect 164660 68388 164666 68400
rect 195054 68388 195060 68400
rect 164660 68360 195060 68388
rect 164660 68348 164666 68360
rect 195054 68348 195060 68360
rect 195112 68388 195118 68400
rect 423674 68388 423680 68400
rect 195112 68360 423680 68388
rect 195112 68348 195118 68360
rect 423674 68348 423680 68360
rect 423732 68348 423738 68400
rect 147306 68280 147312 68332
rect 147364 68320 147370 68332
rect 189718 68320 189724 68332
rect 147364 68292 189724 68320
rect 147364 68280 147370 68292
rect 189718 68280 189724 68292
rect 189776 68280 189782 68332
rect 213822 68280 213828 68332
rect 213880 68320 213886 68332
rect 536834 68320 536840 68332
rect 213880 68292 536840 68320
rect 213880 68280 213886 68292
rect 536834 68280 536840 68292
rect 536892 68280 536898 68332
rect 142430 68212 142436 68264
rect 142488 68212 142494 68264
rect 168834 68212 168840 68264
rect 168892 68252 168898 68264
rect 169570 68252 169576 68264
rect 168892 68224 169576 68252
rect 168892 68212 168898 68224
rect 169570 68212 169576 68224
rect 169628 68252 169634 68264
rect 203794 68252 203800 68264
rect 169628 68224 203800 68252
rect 169628 68212 169634 68224
rect 203794 68212 203800 68224
rect 203852 68212 203858 68264
rect 168926 68144 168932 68196
rect 168984 68184 168990 68196
rect 169662 68184 169668 68196
rect 168984 68156 169668 68184
rect 168984 68144 168990 68156
rect 169662 68144 169668 68156
rect 169720 68184 169726 68196
rect 199378 68184 199384 68196
rect 169720 68156 199384 68184
rect 169720 68144 169726 68156
rect 199378 68144 199384 68156
rect 199436 68144 199442 68196
rect 152734 68076 152740 68128
rect 152792 68116 152798 68128
rect 186314 68116 186320 68128
rect 152792 68088 186320 68116
rect 152792 68076 152798 68088
rect 186314 68076 186320 68088
rect 186372 68076 186378 68128
rect 154298 68008 154304 68060
rect 154356 68048 154362 68060
rect 186774 68048 186780 68060
rect 154356 68020 186780 68048
rect 154356 68008 154362 68020
rect 186774 68008 186780 68020
rect 186832 68008 186838 68060
rect 156046 67600 156052 67652
rect 156104 67640 156110 67652
rect 156782 67640 156788 67652
rect 156104 67612 156788 67640
rect 156104 67600 156110 67612
rect 156782 67600 156788 67612
rect 156840 67600 156846 67652
rect 114462 67532 114468 67584
rect 114520 67572 114526 67584
rect 147950 67572 147956 67584
rect 114520 67544 147956 67572
rect 114520 67532 114526 67544
rect 147950 67532 147956 67544
rect 148008 67532 148014 67584
rect 161290 67532 161296 67584
rect 161348 67572 161354 67584
rect 189074 67572 189080 67584
rect 161348 67544 189080 67572
rect 161348 67532 161354 67544
rect 189074 67532 189080 67544
rect 189132 67572 189138 67584
rect 189442 67572 189448 67584
rect 189132 67544 189448 67572
rect 189132 67532 189138 67544
rect 189442 67532 189448 67544
rect 189500 67532 189506 67584
rect 108942 67464 108948 67516
rect 109000 67504 109006 67516
rect 142614 67504 142620 67516
rect 109000 67476 142620 67504
rect 109000 67464 109006 67476
rect 142614 67464 142620 67476
rect 142672 67464 142678 67516
rect 160278 67464 160284 67516
rect 160336 67504 160342 67516
rect 160922 67504 160928 67516
rect 160336 67476 160928 67504
rect 160336 67464 160342 67476
rect 160922 67464 160928 67476
rect 160980 67504 160986 67516
rect 195514 67504 195520 67516
rect 160980 67476 195520 67504
rect 160980 67464 160986 67476
rect 195514 67464 195520 67476
rect 195572 67464 195578 67516
rect 115382 67396 115388 67448
rect 115440 67436 115446 67448
rect 148502 67436 148508 67448
rect 115440 67408 148508 67436
rect 115440 67396 115446 67408
rect 148502 67396 148508 67408
rect 148560 67436 148566 67448
rect 148778 67436 148784 67448
rect 148560 67408 148784 67436
rect 148560 67396 148566 67408
rect 148778 67396 148784 67408
rect 148836 67396 148842 67448
rect 174354 67396 174360 67448
rect 174412 67436 174418 67448
rect 174998 67436 175004 67448
rect 174412 67408 175004 67436
rect 174412 67396 174418 67408
rect 174998 67396 175004 67408
rect 175056 67396 175062 67448
rect 176286 67396 176292 67448
rect 176344 67436 176350 67448
rect 208854 67436 208860 67448
rect 176344 67408 208860 67436
rect 176344 67396 176350 67408
rect 208854 67396 208860 67408
rect 208912 67396 208918 67448
rect 116210 67328 116216 67380
rect 116268 67368 116274 67380
rect 149054 67368 149060 67380
rect 116268 67340 149060 67368
rect 116268 67328 116274 67340
rect 149054 67328 149060 67340
rect 149112 67368 149118 67380
rect 149882 67368 149888 67380
rect 149112 67340 149888 67368
rect 149112 67328 149118 67340
rect 149882 67328 149888 67340
rect 149940 67328 149946 67380
rect 155034 67328 155040 67380
rect 155092 67368 155098 67380
rect 155862 67368 155868 67380
rect 155092 67340 155868 67368
rect 155092 67328 155098 67340
rect 155862 67328 155868 67340
rect 155920 67368 155926 67380
rect 189166 67368 189172 67380
rect 155920 67340 189172 67368
rect 155920 67328 155926 67340
rect 189166 67328 189172 67340
rect 189224 67328 189230 67380
rect 103238 67260 103244 67312
rect 103296 67300 103302 67312
rect 135806 67300 135812 67312
rect 103296 67272 135812 67300
rect 103296 67260 103302 67272
rect 40034 66920 40040 66972
rect 40092 66960 40098 66972
rect 103486 66960 103514 67272
rect 135806 67260 135812 67272
rect 135864 67260 135870 67312
rect 174262 67260 174268 67312
rect 174320 67300 174326 67312
rect 174906 67300 174912 67312
rect 174320 67272 174912 67300
rect 174320 67260 174326 67272
rect 174906 67260 174912 67272
rect 174964 67260 174970 67312
rect 174998 67260 175004 67312
rect 175056 67300 175062 67312
rect 208670 67300 208676 67312
rect 175056 67272 208676 67300
rect 175056 67260 175062 67272
rect 208670 67260 208676 67272
rect 208728 67260 208734 67312
rect 109034 67192 109040 67244
rect 109092 67232 109098 67244
rect 138566 67232 138572 67244
rect 109092 67204 138572 67232
rect 109092 67192 109098 67204
rect 138566 67192 138572 67204
rect 138624 67192 138630 67244
rect 164050 67192 164056 67244
rect 164108 67232 164114 67244
rect 196986 67232 196992 67244
rect 164108 67204 196992 67232
rect 164108 67192 164114 67204
rect 196986 67192 196992 67204
rect 197044 67192 197050 67244
rect 174170 67124 174176 67176
rect 174228 67164 174234 67176
rect 174814 67164 174820 67176
rect 174228 67136 174820 67164
rect 174228 67124 174234 67136
rect 174814 67124 174820 67136
rect 174872 67124 174878 67176
rect 175550 67124 175556 67176
rect 175608 67164 175614 67176
rect 201678 67164 201684 67176
rect 175608 67136 201684 67164
rect 175608 67124 175614 67136
rect 201678 67124 201684 67136
rect 201736 67164 201742 67176
rect 202782 67164 202788 67176
rect 201736 67136 202788 67164
rect 201736 67124 201742 67136
rect 202782 67124 202788 67136
rect 202840 67124 202846 67176
rect 172882 67056 172888 67108
rect 172940 67096 172946 67108
rect 199194 67096 199200 67108
rect 172940 67068 199200 67096
rect 172940 67056 172946 67068
rect 199194 67056 199200 67068
rect 199252 67056 199258 67108
rect 169754 66988 169760 67040
rect 169812 67028 169818 67040
rect 193398 67028 193404 67040
rect 169812 67000 193404 67028
rect 169812 66988 169818 67000
rect 193398 66988 193404 67000
rect 193456 67028 193462 67040
rect 194502 67028 194508 67040
rect 193456 67000 194508 67028
rect 193456 66988 193462 67000
rect 194502 66988 194508 67000
rect 194560 66988 194566 67040
rect 40092 66932 103514 66960
rect 40092 66920 40098 66932
rect 168098 66920 168104 66972
rect 168156 66960 168162 66972
rect 184382 66960 184388 66972
rect 168156 66932 184388 66960
rect 168156 66920 168162 66932
rect 184382 66920 184388 66932
rect 184440 66920 184446 66972
rect 97442 66852 97448 66904
rect 97500 66892 97506 66904
rect 113174 66892 113180 66904
rect 97500 66864 113180 66892
rect 97500 66852 97506 66864
rect 113174 66852 113180 66864
rect 113232 66892 113238 66904
rect 141050 66892 141056 66904
rect 113232 66864 141056 66892
rect 113232 66852 113238 66864
rect 141050 66852 141056 66864
rect 141108 66852 141114 66904
rect 174906 66852 174912 66904
rect 174964 66892 174970 66904
rect 176286 66892 176292 66904
rect 174964 66864 176292 66892
rect 174964 66852 174970 66864
rect 176286 66852 176292 66864
rect 176344 66852 176350 66904
rect 189074 66852 189080 66904
rect 189132 66892 189138 66904
rect 317414 66892 317420 66904
rect 189132 66864 317420 66892
rect 189132 66852 189138 66864
rect 317414 66852 317420 66864
rect 317472 66852 317478 66904
rect 174814 66784 174820 66836
rect 174872 66824 174878 66836
rect 208946 66824 208952 66836
rect 174872 66796 208952 66824
rect 174872 66784 174878 66796
rect 208946 66784 208952 66796
rect 209004 66784 209010 66836
rect 194502 66376 194508 66428
rect 194560 66416 194566 66428
rect 494054 66416 494060 66428
rect 194560 66388 494060 66416
rect 194560 66376 194566 66388
rect 494054 66376 494060 66388
rect 494112 66376 494118 66428
rect 199194 66308 199200 66360
rect 199252 66348 199258 66360
rect 529934 66348 529940 66360
rect 199252 66320 529940 66348
rect 199252 66308 199258 66320
rect 529934 66308 529940 66320
rect 529992 66308 529998 66360
rect 202782 66240 202788 66292
rect 202840 66280 202846 66292
rect 554038 66280 554044 66292
rect 202840 66252 554044 66280
rect 202840 66240 202846 66252
rect 554038 66240 554044 66252
rect 554096 66240 554102 66292
rect 121822 66172 121828 66224
rect 121880 66212 121886 66224
rect 155954 66212 155960 66224
rect 121880 66184 155960 66212
rect 121880 66172 121886 66184
rect 155954 66172 155960 66184
rect 156012 66172 156018 66224
rect 160186 66172 160192 66224
rect 160244 66212 160250 66224
rect 161290 66212 161296 66224
rect 160244 66184 161296 66212
rect 160244 66172 160250 66184
rect 161290 66172 161296 66184
rect 161348 66212 161354 66224
rect 208762 66212 208768 66224
rect 161348 66184 208768 66212
rect 161348 66172 161354 66184
rect 208762 66172 208768 66184
rect 208820 66172 208826 66224
rect 101398 66104 101404 66156
rect 101456 66144 101462 66156
rect 135530 66144 135536 66156
rect 101456 66116 135536 66144
rect 101456 66104 101462 66116
rect 135530 66104 135536 66116
rect 135588 66104 135594 66156
rect 138106 66104 138112 66156
rect 138164 66144 138170 66156
rect 138658 66144 138664 66156
rect 138164 66116 138664 66144
rect 138164 66104 138170 66116
rect 138658 66104 138664 66116
rect 138716 66104 138722 66156
rect 163038 66104 163044 66156
rect 163096 66144 163102 66156
rect 163774 66144 163780 66156
rect 163096 66116 163780 66144
rect 163096 66104 163102 66116
rect 163774 66104 163780 66116
rect 163832 66144 163838 66156
rect 204346 66144 204352 66156
rect 163832 66116 204352 66144
rect 163832 66104 163838 66116
rect 204346 66104 204352 66116
rect 204404 66104 204410 66156
rect 108298 66036 108304 66088
rect 108356 66076 108362 66088
rect 140222 66076 140228 66088
rect 108356 66048 140228 66076
rect 108356 66036 108362 66048
rect 140222 66036 140228 66048
rect 140280 66036 140286 66088
rect 154850 66036 154856 66088
rect 154908 66076 154914 66088
rect 189074 66076 189080 66088
rect 154908 66048 189080 66076
rect 154908 66036 154914 66048
rect 189074 66036 189080 66048
rect 189132 66036 189138 66088
rect 204162 66036 204168 66088
rect 204220 66076 204226 66088
rect 211430 66076 211436 66088
rect 204220 66048 211436 66076
rect 204220 66036 204226 66048
rect 211430 66036 211436 66048
rect 211488 66036 211494 66088
rect 102134 65968 102140 66020
rect 102192 66008 102198 66020
rect 103330 66008 103336 66020
rect 102192 65980 103336 66008
rect 102192 65968 102198 65980
rect 103330 65968 103336 65980
rect 103388 66008 103394 66020
rect 134242 66008 134248 66020
rect 103388 65980 134248 66008
rect 103388 65968 103394 65980
rect 134242 65968 134248 65980
rect 134300 65968 134306 66020
rect 164510 65968 164516 66020
rect 164568 66008 164574 66020
rect 198918 66008 198924 66020
rect 164568 65980 198924 66008
rect 164568 65968 164574 65980
rect 198918 65968 198924 65980
rect 198976 65968 198982 66020
rect 108114 65900 108120 65952
rect 108172 65940 108178 65952
rect 138106 65940 138112 65952
rect 108172 65912 138112 65940
rect 108172 65900 108178 65912
rect 138106 65900 138112 65912
rect 138164 65900 138170 65952
rect 158806 65900 158812 65952
rect 158864 65940 158870 65952
rect 191926 65940 191932 65952
rect 158864 65912 191932 65940
rect 158864 65900 158870 65912
rect 191926 65900 191932 65912
rect 191984 65940 191990 65952
rect 193030 65940 193036 65952
rect 191984 65912 193036 65940
rect 191984 65900 191990 65912
rect 193030 65900 193036 65912
rect 193088 65900 193094 65952
rect 104618 65832 104624 65884
rect 104676 65872 104682 65884
rect 133046 65872 133052 65884
rect 104676 65844 133052 65872
rect 104676 65832 104682 65844
rect 133046 65832 133052 65844
rect 133104 65832 133110 65884
rect 172790 65832 172796 65884
rect 172848 65872 172854 65884
rect 196158 65872 196164 65884
rect 172848 65844 196164 65872
rect 172848 65832 172854 65844
rect 196158 65832 196164 65844
rect 196216 65832 196222 65884
rect 111242 65764 111248 65816
rect 111300 65804 111306 65816
rect 139946 65804 139952 65816
rect 111300 65776 139952 65804
rect 111300 65764 111306 65776
rect 139946 65764 139952 65776
rect 140004 65764 140010 65816
rect 155954 65764 155960 65816
rect 156012 65804 156018 65816
rect 156782 65804 156788 65816
rect 156012 65776 156788 65804
rect 156012 65764 156018 65776
rect 156782 65764 156788 65776
rect 156840 65764 156846 65816
rect 148134 65696 148140 65748
rect 148192 65736 148198 65748
rect 207658 65736 207664 65748
rect 148192 65708 207664 65736
rect 148192 65696 148198 65708
rect 207658 65696 207664 65708
rect 207716 65696 207722 65748
rect 189074 65628 189080 65680
rect 189132 65668 189138 65680
rect 295334 65668 295340 65680
rect 189132 65640 295340 65668
rect 189132 65628 189138 65640
rect 295334 65628 295340 65640
rect 295392 65628 295398 65680
rect 193030 65560 193036 65612
rect 193088 65600 193094 65612
rect 351914 65600 351920 65612
rect 193088 65572 351920 65600
rect 193088 65560 193094 65572
rect 351914 65560 351920 65572
rect 351972 65560 351978 65612
rect 35986 65492 35992 65544
rect 36044 65532 36050 65544
rect 102134 65532 102140 65544
rect 36044 65504 102140 65532
rect 36044 65492 36050 65504
rect 102134 65492 102140 65504
rect 102192 65492 102198 65544
rect 109494 65492 109500 65544
rect 109552 65532 109558 65544
rect 117314 65532 117320 65544
rect 109552 65504 117320 65532
rect 109552 65492 109558 65504
rect 117314 65492 117320 65504
rect 117372 65532 117378 65544
rect 141142 65532 141148 65544
rect 117372 65504 141148 65532
rect 117372 65492 117378 65504
rect 141142 65492 141148 65504
rect 141200 65492 141206 65544
rect 198918 65492 198924 65544
rect 198976 65532 198982 65544
rect 414658 65532 414664 65544
rect 198976 65504 414664 65532
rect 198976 65492 198982 65504
rect 414658 65492 414664 65504
rect 414716 65492 414722 65544
rect 196158 64880 196164 64932
rect 196216 64920 196222 64932
rect 525794 64920 525800 64932
rect 196216 64892 525800 64920
rect 196216 64880 196222 64892
rect 525794 64880 525800 64892
rect 525852 64880 525858 64932
rect 103054 64812 103060 64864
rect 103112 64852 103118 64864
rect 137278 64852 137284 64864
rect 103112 64824 137284 64852
rect 103112 64812 103118 64824
rect 137278 64812 137284 64824
rect 137336 64812 137342 64864
rect 164418 64812 164424 64864
rect 164476 64852 164482 64864
rect 199654 64852 199660 64864
rect 164476 64824 199660 64852
rect 164476 64812 164482 64824
rect 199654 64812 199660 64824
rect 199712 64812 199718 64864
rect 104710 64744 104716 64796
rect 104768 64784 104774 64796
rect 136818 64784 136824 64796
rect 104768 64756 136824 64784
rect 104768 64744 104774 64756
rect 136818 64744 136824 64756
rect 136876 64744 136882 64796
rect 156138 64744 156144 64796
rect 156196 64784 156202 64796
rect 190638 64784 190644 64796
rect 156196 64756 190644 64784
rect 156196 64744 156202 64756
rect 190638 64744 190644 64756
rect 190696 64784 190702 64796
rect 191742 64784 191748 64796
rect 190696 64756 191748 64784
rect 190696 64744 190702 64756
rect 191742 64744 191748 64756
rect 191800 64744 191806 64796
rect 111242 64676 111248 64728
rect 111300 64716 111306 64728
rect 139854 64716 139860 64728
rect 111300 64688 139860 64716
rect 111300 64676 111306 64688
rect 139854 64676 139860 64688
rect 139912 64676 139918 64728
rect 165890 64676 165896 64728
rect 165948 64716 165954 64728
rect 200114 64716 200120 64728
rect 165948 64688 200120 64716
rect 165948 64676 165954 64688
rect 200114 64676 200120 64688
rect 200172 64676 200178 64728
rect 168742 64608 168748 64660
rect 168800 64648 168806 64660
rect 202966 64648 202972 64660
rect 168800 64620 202972 64648
rect 168800 64608 168806 64620
rect 202966 64608 202972 64620
rect 203024 64608 203030 64660
rect 174078 64540 174084 64592
rect 174136 64580 174142 64592
rect 198918 64580 198924 64592
rect 174136 64552 198924 64580
rect 174136 64540 174142 64552
rect 198918 64540 198924 64552
rect 198976 64540 198982 64592
rect 161566 64472 161572 64524
rect 161624 64512 161630 64524
rect 162302 64512 162308 64524
rect 161624 64484 162308 64512
rect 161624 64472 161630 64484
rect 162302 64472 162308 64484
rect 162360 64512 162366 64524
rect 185670 64512 185676 64524
rect 162360 64484 185676 64512
rect 162360 64472 162366 64484
rect 185670 64472 185676 64484
rect 185728 64472 185734 64524
rect 62114 64200 62120 64252
rect 62172 64240 62178 64252
rect 103054 64240 103060 64252
rect 62172 64212 103060 64240
rect 62172 64200 62178 64212
rect 103054 64200 103060 64212
rect 103112 64200 103118 64252
rect 191742 64200 191748 64252
rect 191800 64240 191806 64252
rect 306374 64240 306380 64252
rect 191800 64212 306380 64240
rect 191800 64200 191806 64212
rect 306374 64200 306380 64212
rect 306432 64200 306438 64252
rect 57238 64132 57244 64184
rect 57296 64172 57302 64184
rect 104710 64172 104716 64184
rect 57296 64144 104716 64172
rect 57296 64132 57302 64144
rect 104710 64132 104716 64144
rect 104768 64132 104774 64184
rect 106734 64132 106740 64184
rect 106792 64172 106798 64184
rect 120074 64172 120080 64184
rect 106792 64144 120080 64172
rect 106792 64132 106798 64144
rect 120074 64132 120080 64144
rect 120132 64172 120138 64184
rect 141234 64172 141240 64184
rect 120132 64144 141240 64172
rect 120132 64132 120138 64144
rect 141234 64132 141240 64144
rect 141292 64132 141298 64184
rect 146386 64132 146392 64184
rect 146444 64172 146450 64184
rect 185578 64172 185584 64184
rect 146444 64144 185584 64172
rect 146444 64132 146450 64144
rect 185578 64132 185584 64144
rect 185636 64132 185642 64184
rect 202966 64132 202972 64184
rect 203024 64172 203030 64184
rect 472618 64172 472624 64184
rect 203024 64144 472624 64172
rect 203024 64132 203030 64144
rect 472618 64132 472624 64144
rect 472676 64132 472682 64184
rect 164418 63860 164424 63912
rect 164476 63900 164482 63912
rect 165246 63900 165252 63912
rect 164476 63872 165252 63900
rect 164476 63860 164482 63872
rect 165246 63860 165252 63872
rect 165304 63860 165310 63912
rect 165890 63860 165896 63912
rect 165948 63900 165954 63912
rect 166626 63900 166632 63912
rect 165948 63872 166632 63900
rect 165948 63860 165954 63872
rect 166626 63860 166632 63872
rect 166684 63860 166690 63912
rect 144454 63520 144460 63572
rect 144512 63560 144518 63572
rect 147214 63560 147220 63572
rect 144512 63532 147220 63560
rect 144512 63520 144518 63532
rect 147214 63520 147220 63532
rect 147272 63520 147278 63572
rect 198918 63520 198924 63572
rect 198976 63560 198982 63572
rect 543734 63560 543740 63572
rect 198976 63532 543740 63560
rect 198976 63520 198982 63532
rect 543734 63520 543740 63532
rect 543792 63520 543798 63572
rect 106090 63452 106096 63504
rect 106148 63492 106154 63504
rect 137002 63492 137008 63504
rect 106148 63464 137008 63492
rect 106148 63452 106154 63464
rect 137002 63452 137008 63464
rect 137060 63452 137066 63504
rect 164326 63452 164332 63504
rect 164384 63492 164390 63504
rect 198734 63492 198740 63504
rect 164384 63464 198740 63492
rect 164384 63452 164390 63464
rect 198734 63452 198740 63464
rect 198792 63452 198798 63504
rect 115106 63384 115112 63436
rect 115164 63424 115170 63436
rect 138474 63424 138480 63436
rect 115164 63396 138480 63424
rect 115164 63384 115170 63396
rect 138474 63384 138480 63396
rect 138532 63384 138538 63436
rect 154758 63384 154764 63436
rect 154816 63424 154822 63436
rect 189074 63424 189080 63436
rect 154816 63396 189080 63424
rect 154816 63384 154822 63396
rect 189074 63384 189080 63396
rect 189132 63384 189138 63436
rect 166442 63316 166448 63368
rect 166500 63356 166506 63368
rect 187234 63356 187240 63368
rect 166500 63328 187240 63356
rect 166500 63316 166506 63328
rect 187234 63316 187240 63328
rect 187292 63316 187298 63368
rect 144362 63180 144368 63232
rect 144420 63220 144426 63232
rect 148318 63220 148324 63232
rect 144420 63192 148324 63220
rect 144420 63180 144426 63192
rect 148318 63180 148324 63192
rect 148376 63180 148382 63232
rect 150802 62908 150808 62960
rect 150860 62948 150866 62960
rect 245654 62948 245660 62960
rect 150860 62920 245660 62948
rect 150860 62908 150866 62920
rect 245654 62908 245660 62920
rect 245712 62908 245718 62960
rect 189074 62840 189080 62892
rect 189132 62880 189138 62892
rect 189994 62880 190000 62892
rect 189132 62852 190000 62880
rect 189132 62840 189138 62852
rect 189994 62840 190000 62852
rect 190052 62880 190058 62892
rect 292574 62880 292580 62892
rect 190052 62852 292580 62880
rect 190052 62840 190058 62852
rect 292574 62840 292580 62852
rect 292632 62840 292638 62892
rect 69014 62772 69020 62824
rect 69072 62812 69078 62824
rect 106090 62812 106096 62824
rect 69072 62784 106096 62812
rect 69072 62772 69078 62784
rect 106090 62772 106096 62784
rect 106148 62772 106154 62824
rect 198734 62772 198740 62824
rect 198792 62812 198798 62824
rect 412634 62812 412640 62824
rect 198792 62784 412640 62812
rect 198792 62772 198798 62784
rect 412634 62772 412640 62784
rect 412692 62772 412698 62824
rect 138658 62568 138664 62620
rect 138716 62608 138722 62620
rect 142430 62608 142436 62620
rect 138716 62580 142436 62608
rect 138716 62568 138722 62580
rect 142430 62568 142436 62580
rect 142488 62568 142494 62620
rect 187234 62092 187240 62144
rect 187292 62132 187298 62144
rect 368474 62132 368480 62144
rect 187292 62104 368480 62132
rect 187292 62092 187298 62104
rect 368474 62092 368480 62104
rect 368532 62092 368538 62144
rect 102134 62024 102140 62076
rect 102192 62064 102198 62076
rect 103146 62064 103152 62076
rect 102192 62036 103152 62064
rect 102192 62024 102198 62036
rect 103146 62024 103152 62036
rect 103204 62064 103210 62076
rect 135438 62064 135444 62076
rect 103204 62036 135444 62064
rect 103204 62024 103210 62036
rect 135438 62024 135444 62036
rect 135496 62024 135502 62076
rect 162946 62024 162952 62076
rect 163004 62064 163010 62076
rect 197722 62064 197728 62076
rect 163004 62036 197728 62064
rect 163004 62024 163010 62036
rect 197722 62024 197728 62036
rect 197780 62064 197786 62076
rect 198182 62064 198188 62076
rect 197780 62036 198188 62064
rect 197780 62024 197786 62036
rect 198182 62024 198188 62036
rect 198240 62024 198246 62076
rect 153194 61956 153200 62008
rect 153252 61996 153258 62008
rect 187878 61996 187884 62008
rect 153252 61968 187884 61996
rect 153252 61956 153258 61968
rect 187878 61956 187884 61968
rect 187936 61956 187942 62008
rect 157058 61888 157064 61940
rect 157116 61928 157122 61940
rect 190546 61928 190552 61940
rect 157116 61900 190552 61928
rect 157116 61888 157122 61900
rect 190546 61888 190552 61900
rect 190604 61928 190610 61940
rect 191742 61928 191748 61940
rect 190604 61900 191748 61928
rect 190604 61888 190610 61900
rect 191742 61888 191748 61900
rect 191800 61888 191806 61940
rect 172698 61820 172704 61872
rect 172756 61860 172762 61872
rect 202138 61860 202144 61872
rect 172756 61832 202144 61860
rect 172756 61820 172762 61832
rect 202138 61820 202144 61832
rect 202196 61860 202202 61872
rect 202782 61860 202788 61872
rect 202196 61832 202788 61860
rect 202196 61820 202202 61832
rect 202782 61820 202788 61832
rect 202840 61820 202846 61872
rect 187878 61480 187884 61532
rect 187936 61520 187942 61532
rect 188706 61520 188712 61532
rect 187936 61492 188712 61520
rect 187936 61480 187942 61492
rect 188706 61480 188712 61492
rect 188764 61520 188770 61532
rect 277394 61520 277400 61532
rect 188764 61492 277400 61520
rect 188764 61480 188770 61492
rect 277394 61480 277400 61492
rect 277452 61480 277458 61532
rect 191742 61412 191748 61464
rect 191800 61452 191806 61464
rect 313274 61452 313280 61464
rect 191800 61424 313280 61452
rect 191800 61412 191806 61424
rect 313274 61412 313280 61424
rect 313332 61412 313338 61464
rect 43438 61344 43444 61396
rect 43496 61384 43502 61396
rect 102134 61384 102140 61396
rect 43496 61356 102140 61384
rect 43496 61344 43502 61356
rect 102134 61344 102140 61356
rect 102192 61344 102198 61396
rect 147766 61344 147772 61396
rect 147824 61384 147830 61396
rect 197446 61384 197452 61396
rect 147824 61356 197452 61384
rect 147824 61344 147830 61356
rect 197446 61344 197452 61356
rect 197504 61344 197510 61396
rect 198182 61344 198188 61396
rect 198240 61384 198246 61396
rect 398834 61384 398840 61396
rect 198240 61356 398840 61384
rect 198240 61344 198246 61356
rect 398834 61344 398840 61356
rect 398892 61344 398898 61396
rect 202782 60732 202788 60784
rect 202840 60772 202846 60784
rect 527818 60772 527824 60784
rect 202840 60744 527824 60772
rect 202840 60732 202846 60744
rect 527818 60732 527824 60744
rect 527876 60732 527882 60784
rect 102134 60664 102140 60716
rect 102192 60704 102198 60716
rect 103422 60704 103428 60716
rect 102192 60676 103428 60704
rect 102192 60664 102198 60676
rect 103422 60664 103428 60676
rect 103480 60704 103486 60716
rect 135898 60704 135904 60716
rect 103480 60676 135904 60704
rect 103480 60664 103486 60676
rect 135898 60664 135904 60676
rect 135956 60664 135962 60716
rect 158714 60664 158720 60716
rect 158772 60704 158778 60716
rect 193490 60704 193496 60716
rect 158772 60676 193496 60704
rect 158772 60664 158778 60676
rect 193490 60664 193496 60676
rect 193548 60704 193554 60716
rect 194502 60704 194508 60716
rect 193548 60676 194508 60704
rect 193548 60664 193554 60676
rect 194502 60664 194508 60676
rect 194560 60664 194566 60716
rect 162854 60596 162860 60648
rect 162912 60636 162918 60648
rect 197722 60636 197728 60648
rect 162912 60608 197728 60636
rect 162912 60596 162918 60608
rect 197722 60596 197728 60608
rect 197780 60596 197786 60648
rect 154666 60528 154672 60580
rect 154724 60568 154730 60580
rect 189074 60568 189080 60580
rect 154724 60540 189080 60568
rect 154724 60528 154730 60540
rect 189074 60528 189080 60540
rect 189132 60528 189138 60580
rect 166534 60460 166540 60512
rect 166592 60500 166598 60512
rect 197814 60500 197820 60512
rect 166592 60472 197820 60500
rect 166592 60460 166598 60472
rect 197814 60460 197820 60472
rect 197872 60460 197878 60512
rect 147950 60324 147956 60376
rect 148008 60364 148014 60376
rect 198734 60364 198740 60376
rect 148008 60336 198740 60364
rect 148008 60324 148014 60336
rect 198734 60324 198740 60336
rect 198792 60324 198798 60376
rect 149606 60256 149612 60308
rect 149664 60296 149670 60308
rect 231854 60296 231860 60308
rect 149664 60268 231860 60296
rect 149664 60256 149670 60268
rect 231854 60256 231860 60268
rect 231912 60256 231918 60308
rect 145282 60188 145288 60240
rect 145340 60228 145346 60240
rect 148410 60228 148416 60240
rect 145340 60200 148416 60228
rect 145340 60188 145346 60200
rect 148410 60188 148416 60200
rect 148468 60188 148474 60240
rect 189074 60188 189080 60240
rect 189132 60228 189138 60240
rect 190086 60228 190092 60240
rect 189132 60200 190092 60228
rect 189132 60188 189138 60200
rect 190086 60188 190092 60200
rect 190144 60228 190150 60240
rect 299474 60228 299480 60240
rect 190144 60200 299480 60228
rect 190144 60188 190150 60200
rect 299474 60188 299480 60200
rect 299532 60188 299538 60240
rect 194502 60120 194508 60172
rect 194560 60160 194566 60172
rect 340966 60160 340972 60172
rect 194560 60132 340972 60160
rect 194560 60120 194566 60132
rect 340966 60120 340972 60132
rect 341024 60120 341030 60172
rect 197722 60052 197728 60104
rect 197780 60092 197786 60104
rect 198366 60092 198372 60104
rect 197780 60064 198372 60092
rect 197780 60052 197786 60064
rect 198366 60052 198372 60064
rect 198424 60092 198430 60104
rect 394694 60092 394700 60104
rect 198424 60064 394700 60092
rect 198424 60052 198430 60064
rect 394694 60052 394700 60064
rect 394752 60052 394758 60104
rect 52546 59984 52552 60036
rect 52604 60024 52610 60036
rect 102134 60024 102140 60036
rect 52604 59996 102140 60024
rect 52604 59984 52610 59996
rect 102134 59984 102140 59996
rect 102192 59984 102198 60036
rect 197814 59984 197820 60036
rect 197872 60024 197878 60036
rect 198458 60024 198464 60036
rect 197872 59996 198464 60024
rect 197872 59984 197878 59996
rect 198458 59984 198464 59996
rect 198516 60024 198522 60036
rect 396074 60024 396080 60036
rect 198516 59996 396080 60024
rect 198516 59984 198522 59996
rect 396074 59984 396080 59996
rect 396132 59984 396138 60036
rect 157518 59304 157524 59356
rect 157576 59344 157582 59356
rect 191926 59344 191932 59356
rect 157576 59316 191932 59344
rect 157576 59304 157582 59316
rect 191926 59304 191932 59316
rect 191984 59344 191990 59356
rect 193030 59344 193036 59356
rect 191984 59316 193036 59344
rect 191984 59304 191990 59316
rect 193030 59304 193036 59316
rect 193088 59304 193094 59356
rect 139394 58760 139400 58812
rect 139452 58800 139458 58812
rect 142154 58800 142160 58812
rect 139452 58772 142160 58800
rect 139452 58760 139458 58772
rect 142154 58760 142160 58772
rect 142212 58760 142218 58812
rect 151722 58692 151728 58744
rect 151780 58732 151786 58744
rect 249794 58732 249800 58744
rect 151780 58704 249800 58732
rect 151780 58692 151786 58704
rect 249794 58692 249800 58704
rect 249852 58692 249858 58744
rect 193030 58624 193036 58676
rect 193088 58664 193094 58676
rect 327074 58664 327080 58676
rect 193088 58636 327080 58664
rect 193088 58624 193094 58636
rect 327074 58624 327080 58636
rect 327132 58624 327138 58676
rect 168650 57876 168656 57928
rect 168708 57916 168714 57928
rect 203242 57916 203248 57928
rect 168708 57888 203248 57916
rect 168708 57876 168714 57888
rect 203242 57876 203248 57888
rect 203300 57916 203306 57928
rect 204070 57916 204076 57928
rect 203300 57888 204076 57916
rect 203300 57876 203306 57888
rect 204070 57876 204076 57888
rect 204128 57876 204134 57928
rect 173986 57808 173992 57860
rect 174044 57848 174050 57860
rect 204990 57848 204996 57860
rect 174044 57820 204996 57848
rect 174044 57808 174050 57820
rect 204990 57808 204996 57820
rect 205048 57808 205054 57860
rect 176930 57740 176936 57792
rect 176988 57780 176994 57792
rect 197998 57780 198004 57792
rect 176988 57752 198004 57780
rect 176988 57740 176994 57752
rect 197998 57740 198004 57752
rect 198056 57740 198062 57792
rect 152366 57264 152372 57316
rect 152424 57304 152430 57316
rect 263594 57304 263600 57316
rect 152424 57276 263600 57304
rect 152424 57264 152430 57276
rect 263594 57264 263600 57276
rect 263652 57264 263658 57316
rect 145650 57196 145656 57248
rect 145708 57236 145714 57248
rect 169754 57236 169760 57248
rect 145708 57208 169760 57236
rect 145708 57196 145714 57208
rect 169754 57196 169760 57208
rect 169812 57196 169818 57248
rect 204990 57196 204996 57248
rect 205048 57236 205054 57248
rect 545114 57236 545120 57248
rect 205048 57208 545120 57236
rect 205048 57196 205054 57208
rect 545114 57196 545120 57208
rect 545172 57196 545178 57248
rect 204070 56652 204076 56704
rect 204128 56692 204134 56704
rect 473446 56692 473452 56704
rect 204128 56664 473452 56692
rect 204128 56652 204134 56664
rect 473446 56652 473452 56664
rect 473504 56652 473510 56704
rect 197998 56584 198004 56636
rect 198056 56624 198062 56636
rect 567838 56624 567844 56636
rect 198056 56596 567844 56624
rect 198056 56584 198062 56596
rect 567838 56584 567844 56596
rect 567896 56584 567902 56636
rect 104434 56516 104440 56568
rect 104492 56556 104498 56568
rect 137094 56556 137100 56568
rect 104492 56528 137100 56556
rect 104492 56516 104498 56528
rect 137094 56516 137100 56528
rect 137152 56516 137158 56568
rect 157426 56516 157432 56568
rect 157484 56556 157490 56568
rect 187970 56556 187976 56568
rect 157484 56528 187976 56556
rect 157484 56516 157490 56528
rect 187970 56516 187976 56528
rect 188028 56516 188034 56568
rect 149422 55904 149428 55956
rect 149480 55944 149486 55956
rect 229094 55944 229100 55956
rect 149480 55916 229100 55944
rect 149480 55904 149486 55916
rect 229094 55904 229100 55916
rect 229152 55904 229158 55956
rect 187970 55836 187976 55888
rect 188028 55876 188034 55888
rect 331214 55876 331220 55888
rect 188028 55848 331220 55876
rect 188028 55836 188034 55848
rect 331214 55836 331220 55848
rect 331272 55836 331278 55888
rect 136634 55224 136640 55276
rect 136692 55264 136698 55276
rect 142338 55264 142344 55276
rect 136692 55236 142344 55264
rect 136692 55224 136698 55236
rect 142338 55224 142344 55236
rect 142396 55224 142402 55276
rect 156966 55156 156972 55208
rect 157024 55196 157030 55208
rect 189350 55196 189356 55208
rect 157024 55168 189356 55196
rect 157024 55156 157030 55168
rect 189350 55156 189356 55168
rect 189408 55156 189414 55208
rect 150434 54544 150440 54596
rect 150492 54584 150498 54596
rect 239398 54584 239404 54596
rect 150492 54556 239404 54584
rect 150492 54544 150498 54556
rect 239398 54544 239404 54556
rect 239456 54544 239462 54596
rect 189350 54476 189356 54528
rect 189408 54516 189414 54528
rect 315298 54516 315304 54528
rect 189408 54488 315304 54516
rect 189408 54476 189414 54488
rect 315298 54476 315304 54488
rect 315356 54476 315362 54528
rect 163498 53728 163504 53780
rect 163556 53768 163562 53780
rect 194318 53768 194324 53780
rect 163556 53740 194324 53768
rect 163556 53728 163562 53740
rect 194318 53728 194324 53740
rect 194376 53728 194382 53780
rect 148686 53184 148692 53236
rect 148744 53224 148750 53236
rect 201586 53224 201592 53236
rect 148744 53196 201592 53224
rect 148744 53184 148750 53196
rect 201586 53184 201592 53196
rect 201644 53184 201650 53236
rect 153010 53116 153016 53168
rect 153068 53156 153074 53168
rect 267734 53156 267740 53168
rect 153068 53128 267740 53156
rect 153068 53116 153074 53128
rect 267734 53116 267740 53128
rect 267792 53116 267798 53168
rect 194318 53048 194324 53100
rect 194376 53088 194382 53100
rect 389174 53088 389180 53100
rect 194376 53060 389180 53088
rect 194376 53048 194382 53060
rect 389174 53048 389180 53060
rect 389232 53048 389238 53100
rect 99466 52368 99472 52420
rect 99524 52408 99530 52420
rect 100478 52408 100484 52420
rect 99524 52380 100484 52408
rect 99524 52368 99530 52380
rect 100478 52368 100484 52380
rect 100536 52408 100542 52420
rect 133138 52408 133144 52420
rect 100536 52380 133144 52408
rect 100536 52368 100542 52380
rect 133138 52368 133144 52380
rect 133196 52368 133202 52420
rect 168374 52368 168380 52420
rect 168432 52408 168438 52420
rect 202874 52408 202880 52420
rect 168432 52380 202880 52408
rect 168432 52368 168438 52380
rect 202874 52368 202880 52380
rect 202932 52408 202938 52420
rect 204070 52408 204076 52420
rect 202932 52380 204076 52408
rect 202932 52368 202938 52380
rect 204070 52368 204076 52380
rect 204128 52368 204134 52420
rect 150250 51756 150256 51808
rect 150308 51796 150314 51808
rect 224954 51796 224960 51808
rect 150308 51768 224960 51796
rect 150308 51756 150314 51768
rect 224954 51756 224960 51768
rect 225012 51756 225018 51808
rect 17954 51688 17960 51740
rect 18012 51728 18018 51740
rect 99466 51728 99472 51740
rect 18012 51700 99472 51728
rect 18012 51688 18018 51700
rect 99466 51688 99472 51700
rect 99524 51688 99530 51740
rect 204070 51688 204076 51740
rect 204128 51728 204134 51740
rect 464338 51728 464344 51740
rect 204128 51700 464344 51728
rect 204128 51688 204134 51700
rect 464338 51688 464344 51700
rect 464396 51688 464402 51740
rect 176838 51008 176844 51060
rect 176896 51048 176902 51060
rect 207106 51048 207112 51060
rect 176896 51020 207112 51048
rect 176896 51008 176902 51020
rect 207106 51008 207112 51020
rect 207164 51048 207170 51060
rect 207750 51048 207756 51060
rect 207164 51020 207756 51048
rect 207164 51008 207170 51020
rect 207750 51008 207756 51020
rect 207808 51008 207814 51060
rect 207106 50328 207112 50380
rect 207164 50368 207170 50380
rect 569954 50368 569960 50380
rect 207164 50340 569960 50368
rect 207164 50328 207170 50340
rect 569954 50328 569960 50340
rect 570012 50328 570018 50380
rect 172606 49648 172612 49700
rect 172664 49688 172670 49700
rect 204898 49688 204904 49700
rect 172664 49660 204904 49688
rect 172664 49648 172670 49660
rect 204898 49648 204904 49660
rect 204956 49648 204962 49700
rect 148594 49104 148600 49156
rect 148652 49144 148658 49156
rect 204254 49144 204260 49156
rect 148652 49116 204260 49144
rect 148652 49104 148658 49116
rect 204254 49104 204260 49116
rect 204312 49104 204318 49156
rect 167638 49036 167644 49088
rect 167696 49076 167702 49088
rect 455414 49076 455420 49088
rect 167696 49048 455420 49076
rect 167696 49036 167702 49048
rect 455414 49036 455420 49048
rect 455472 49036 455478 49088
rect 145190 48968 145196 49020
rect 145248 49008 145254 49020
rect 168650 49008 168656 49020
rect 145248 48980 168656 49008
rect 145248 48968 145254 48980
rect 168650 48968 168656 48980
rect 168708 48968 168714 49020
rect 204898 48968 204904 49020
rect 204956 49008 204962 49020
rect 516134 49008 516140 49020
rect 204956 48980 516140 49008
rect 204956 48968 204962 48980
rect 516134 48968 516140 48980
rect 516192 48968 516198 49020
rect 168558 48220 168564 48272
rect 168616 48260 168622 48272
rect 203058 48260 203064 48272
rect 168616 48232 203064 48260
rect 168616 48220 168622 48232
rect 203058 48220 203064 48232
rect 203116 48260 203122 48272
rect 204070 48260 204076 48272
rect 203116 48232 204076 48260
rect 203116 48220 203122 48232
rect 204070 48220 204076 48232
rect 204128 48220 204134 48272
rect 150158 47608 150164 47660
rect 150216 47648 150222 47660
rect 215294 47648 215300 47660
rect 150216 47620 215300 47648
rect 150216 47608 150222 47620
rect 215294 47608 215300 47620
rect 215352 47608 215358 47660
rect 149514 47540 149520 47592
rect 149572 47580 149578 47592
rect 218146 47580 218152 47592
rect 149572 47552 218152 47580
rect 149572 47540 149578 47552
rect 218146 47540 218152 47552
rect 218204 47540 218210 47592
rect 204070 46928 204076 46980
rect 204128 46968 204134 46980
rect 466454 46968 466460 46980
rect 204128 46940 466460 46968
rect 204128 46928 204134 46940
rect 466454 46928 466460 46940
rect 466512 46928 466518 46980
rect 176746 46860 176752 46912
rect 176804 46900 176810 46912
rect 207106 46900 207112 46912
rect 176804 46872 207112 46900
rect 176804 46860 176810 46872
rect 207106 46860 207112 46872
rect 207164 46860 207170 46912
rect 150066 46248 150072 46300
rect 150124 46288 150130 46300
rect 219434 46288 219440 46300
rect 150124 46260 219440 46288
rect 150124 46248 150130 46260
rect 219434 46248 219440 46260
rect 219492 46248 219498 46300
rect 155310 46180 155316 46232
rect 155368 46220 155374 46232
rect 285674 46220 285680 46232
rect 155368 46192 285680 46220
rect 155368 46180 155374 46192
rect 285674 46180 285680 46192
rect 285732 46180 285738 46232
rect 135346 45568 135352 45620
rect 135404 45608 135410 45620
rect 142246 45608 142252 45620
rect 135404 45580 142252 45608
rect 135404 45568 135410 45580
rect 142246 45568 142252 45580
rect 142304 45568 142310 45620
rect 207842 45568 207848 45620
rect 207900 45608 207906 45620
rect 571978 45608 571984 45620
rect 207900 45580 571984 45608
rect 207900 45568 207906 45580
rect 571978 45568 571984 45580
rect 572036 45568 572042 45620
rect 151630 44888 151636 44940
rect 151688 44928 151694 44940
rect 242894 44928 242900 44940
rect 151688 44900 242900 44928
rect 151688 44888 151694 44900
rect 242894 44888 242900 44900
rect 242952 44888 242958 44940
rect 161474 44820 161480 44872
rect 161532 44860 161538 44872
rect 390554 44860 390560 44872
rect 161532 44832 390560 44860
rect 161532 44820 161538 44832
rect 390554 44820 390560 44832
rect 390612 44820 390618 44872
rect 176654 44072 176660 44124
rect 176712 44112 176718 44124
rect 207014 44112 207020 44124
rect 176712 44084 207020 44112
rect 176712 44072 176718 44084
rect 207014 44072 207020 44084
rect 207072 44072 207078 44124
rect 167454 43392 167460 43444
rect 167512 43432 167518 43444
rect 458174 43432 458180 43444
rect 167512 43404 458180 43432
rect 167512 43392 167518 43404
rect 458174 43392 458180 43404
rect 458232 43392 458238 43444
rect 207014 42780 207020 42832
rect 207072 42820 207078 42832
rect 576854 42820 576860 42832
rect 207072 42792 576860 42820
rect 207072 42780 207078 42792
rect 576854 42780 576860 42792
rect 576912 42780 576918 42832
rect 158254 42236 158260 42288
rect 158312 42276 158318 42288
rect 324406 42276 324412 42288
rect 158312 42248 324412 42276
rect 158312 42236 158318 42248
rect 324406 42236 324412 42248
rect 324464 42236 324470 42288
rect 164234 42168 164240 42220
rect 164292 42208 164298 42220
rect 426434 42208 426440 42220
rect 164292 42180 426440 42208
rect 164292 42168 164298 42180
rect 426434 42168 426440 42180
rect 426492 42168 426498 42220
rect 167730 42100 167736 42152
rect 167788 42140 167794 42152
rect 452654 42140 452660 42152
rect 167788 42112 452660 42140
rect 167788 42100 167794 42112
rect 452654 42100 452660 42112
rect 452712 42100 452718 42152
rect 70394 42032 70400 42084
rect 70452 42072 70458 42084
rect 136726 42072 136732 42084
rect 70452 42044 136732 42072
rect 70452 42032 70458 42044
rect 136726 42032 136732 42044
rect 136784 42032 136790 42084
rect 170490 42032 170496 42084
rect 170548 42072 170554 42084
rect 495434 42072 495440 42084
rect 170548 42044 495440 42072
rect 170548 42032 170554 42044
rect 495434 42032 495440 42044
rect 495492 42032 495498 42084
rect 154574 41352 154580 41404
rect 154632 41392 154638 41404
rect 187786 41392 187792 41404
rect 154632 41364 187792 41392
rect 154632 41352 154638 41364
rect 187786 41352 187792 41364
rect 187844 41352 187850 41404
rect 151538 41012 151544 41064
rect 151596 41052 151602 41064
rect 233234 41052 233240 41064
rect 151596 41024 233240 41052
rect 151596 41012 151602 41024
rect 233234 41012 233240 41024
rect 233292 41012 233298 41064
rect 187786 40944 187792 40996
rect 187844 40984 187850 40996
rect 188798 40984 188804 40996
rect 187844 40956 188804 40984
rect 187844 40944 187850 40956
rect 188798 40944 188804 40956
rect 188856 40984 188862 40996
rect 292666 40984 292672 40996
rect 188856 40956 292672 40984
rect 188856 40944 188862 40956
rect 292666 40944 292672 40956
rect 292724 40944 292730 40996
rect 157334 40876 157340 40928
rect 157392 40916 157398 40928
rect 333974 40916 333980 40928
rect 157392 40888 333980 40916
rect 157392 40876 157398 40888
rect 333974 40876 333980 40888
rect 334032 40876 334038 40928
rect 165798 40808 165804 40860
rect 165856 40848 165862 40860
rect 444374 40848 444380 40860
rect 165856 40820 444380 40848
rect 165856 40808 165862 40820
rect 444374 40808 444380 40820
rect 444432 40808 444438 40860
rect 171962 40740 171968 40792
rect 172020 40780 172026 40792
rect 498286 40780 498292 40792
rect 172020 40752 498292 40780
rect 172020 40740 172026 40752
rect 498286 40740 498292 40752
rect 498344 40740 498350 40792
rect 74534 40672 74540 40724
rect 74592 40712 74598 40724
rect 138290 40712 138296 40724
rect 74592 40684 138296 40712
rect 74592 40672 74598 40684
rect 138290 40672 138296 40684
rect 138348 40672 138354 40724
rect 174814 40672 174820 40724
rect 174872 40712 174878 40724
rect 535454 40712 535460 40724
rect 174872 40684 535460 40712
rect 174872 40672 174878 40684
rect 535454 40672 535460 40684
rect 535512 40672 535518 40724
rect 153102 39516 153108 39568
rect 153160 39556 153166 39568
rect 266354 39556 266360 39568
rect 153160 39528 266360 39556
rect 153160 39516 153166 39528
rect 266354 39516 266360 39528
rect 266412 39516 266418 39568
rect 165062 39448 165068 39500
rect 165120 39488 165126 39500
rect 409874 39488 409880 39500
rect 165120 39460 409880 39488
rect 165120 39448 165126 39460
rect 409874 39448 409880 39460
rect 409932 39448 409938 39500
rect 167822 39380 167828 39432
rect 167880 39420 167886 39432
rect 462314 39420 462320 39432
rect 167880 39392 462320 39420
rect 167880 39380 167886 39392
rect 462314 39380 462320 39392
rect 462372 39380 462378 39432
rect 77386 39312 77392 39364
rect 77444 39352 77450 39364
rect 138106 39352 138112 39364
rect 77444 39324 138112 39352
rect 77444 39312 77450 39324
rect 138106 39312 138112 39324
rect 138164 39312 138170 39364
rect 176286 39312 176292 39364
rect 176344 39352 176350 39364
rect 562318 39352 562324 39364
rect 176344 39324 562324 39352
rect 176344 39312 176350 39324
rect 562318 39312 562324 39324
rect 562376 39312 562382 39364
rect 156874 38088 156880 38140
rect 156932 38128 156938 38140
rect 318794 38128 318800 38140
rect 156932 38100 318800 38128
rect 156932 38088 156938 38100
rect 318794 38088 318800 38100
rect 318852 38088 318858 38140
rect 169478 38020 169484 38072
rect 169536 38060 169542 38072
rect 463694 38060 463700 38072
rect 169536 38032 463700 38060
rect 169536 38020 169542 38032
rect 463694 38020 463700 38032
rect 463752 38020 463758 38072
rect 168466 37952 168472 38004
rect 168524 37992 168530 38004
rect 476114 37992 476120 38004
rect 168524 37964 476120 37992
rect 168524 37952 168530 37964
rect 476114 37952 476120 37964
rect 476172 37952 476178 38004
rect 13814 37884 13820 37936
rect 13872 37924 13878 37936
rect 132862 37924 132868 37936
rect 13872 37896 132868 37924
rect 13872 37884 13878 37896
rect 132862 37884 132868 37896
rect 132920 37884 132926 37936
rect 172514 37884 172520 37936
rect 172572 37924 172578 37936
rect 525058 37924 525064 37936
rect 172572 37896 525064 37924
rect 172572 37884 172578 37896
rect 525058 37884 525064 37896
rect 525116 37884 525122 37936
rect 148502 36796 148508 36848
rect 148560 36836 148566 36848
rect 205634 36836 205640 36848
rect 148560 36808 205640 36836
rect 148560 36796 148566 36808
rect 205634 36796 205640 36808
rect 205692 36796 205698 36848
rect 153654 36728 153660 36780
rect 153712 36768 153718 36780
rect 267826 36768 267832 36780
rect 153712 36740 267832 36768
rect 153712 36728 153718 36740
rect 267826 36728 267832 36740
rect 267884 36728 267890 36780
rect 160922 36660 160928 36712
rect 160980 36700 160986 36712
rect 356698 36700 356704 36712
rect 160980 36672 356704 36700
rect 160980 36660 160986 36672
rect 356698 36660 356704 36672
rect 356756 36660 356762 36712
rect 170674 36592 170680 36644
rect 170732 36632 170738 36644
rect 481634 36632 481640 36644
rect 170732 36604 481640 36632
rect 170732 36592 170738 36604
rect 481634 36592 481640 36604
rect 481692 36592 481698 36644
rect 23474 36524 23480 36576
rect 23532 36564 23538 36576
rect 134058 36564 134064 36576
rect 23532 36536 134064 36564
rect 23532 36524 23538 36536
rect 134058 36524 134064 36536
rect 134116 36524 134122 36576
rect 172054 36524 172060 36576
rect 172112 36564 172118 36576
rect 503714 36564 503720 36576
rect 172112 36536 503720 36564
rect 172112 36524 172118 36536
rect 503714 36524 503720 36536
rect 503772 36524 503778 36576
rect 156782 35368 156788 35420
rect 156840 35408 156846 35420
rect 303614 35408 303620 35420
rect 156840 35380 303620 35408
rect 156840 35368 156846 35380
rect 303614 35368 303620 35380
rect 303672 35368 303678 35420
rect 170582 35300 170588 35352
rect 170640 35340 170646 35352
rect 488534 35340 488540 35352
rect 170640 35312 488540 35340
rect 170640 35300 170646 35312
rect 488534 35300 488540 35312
rect 488592 35300 488598 35352
rect 174906 35232 174912 35284
rect 174964 35272 174970 35284
rect 538858 35272 538864 35284
rect 174964 35244 538864 35272
rect 174964 35232 174970 35244
rect 538858 35232 538864 35244
rect 538916 35232 538922 35284
rect 31754 35164 31760 35216
rect 31812 35204 31818 35216
rect 134150 35204 134156 35216
rect 31812 35176 134156 35204
rect 31812 35164 31818 35176
rect 134150 35164 134156 35176
rect 134208 35164 134214 35216
rect 176378 35164 176384 35216
rect 176436 35204 176442 35216
rect 552014 35204 552020 35216
rect 176436 35176 552020 35204
rect 176436 35164 176442 35176
rect 552014 35164 552020 35176
rect 552072 35164 552078 35216
rect 151446 34076 151452 34128
rect 151504 34116 151510 34128
rect 235994 34116 236000 34128
rect 151504 34088 236000 34116
rect 151504 34076 151510 34088
rect 235994 34076 236000 34088
rect 236052 34076 236058 34128
rect 152918 34008 152924 34060
rect 152976 34048 152982 34060
rect 251174 34048 251180 34060
rect 152976 34020 251180 34048
rect 152976 34008 152982 34020
rect 251174 34008 251180 34020
rect 251232 34008 251238 34060
rect 159542 33940 159548 33992
rect 159600 33980 159606 33992
rect 339494 33980 339500 33992
rect 159600 33952 339500 33980
rect 159600 33940 159606 33952
rect 339494 33940 339500 33952
rect 339552 33940 339558 33992
rect 166626 33872 166632 33924
rect 166684 33912 166690 33924
rect 431954 33912 431960 33924
rect 166684 33884 431960 33912
rect 166684 33872 166690 33884
rect 431954 33872 431960 33884
rect 432012 33872 432018 33924
rect 175642 33804 175648 33856
rect 175700 33844 175706 33856
rect 558914 33844 558920 33856
rect 175700 33816 558920 33844
rect 175700 33804 175706 33816
rect 558914 33804 558920 33816
rect 558972 33804 558978 33856
rect 38654 33736 38660 33788
rect 38712 33776 38718 33788
rect 135530 33776 135536 33788
rect 38712 33748 135536 33776
rect 38712 33736 38718 33748
rect 135530 33736 135536 33748
rect 135588 33736 135594 33788
rect 177666 33736 177672 33788
rect 177724 33776 177730 33788
rect 578234 33776 578240 33788
rect 177724 33748 578240 33776
rect 177724 33736 177730 33748
rect 578234 33736 578240 33748
rect 578292 33736 578298 33788
rect 148962 32648 148968 32700
rect 149020 32688 149026 32700
rect 208394 32688 208400 32700
rect 149020 32660 208400 32688
rect 149020 32648 149026 32660
rect 208394 32648 208400 32660
rect 208452 32648 208458 32700
rect 151354 32580 151360 32632
rect 151412 32620 151418 32632
rect 242986 32620 242992 32632
rect 151412 32592 242992 32620
rect 151412 32580 151418 32592
rect 242986 32580 242992 32592
rect 243044 32580 243050 32632
rect 158346 32512 158352 32564
rect 158404 32552 158410 32564
rect 332686 32552 332692 32564
rect 158404 32524 332692 32552
rect 158404 32512 158410 32524
rect 332686 32512 332692 32524
rect 332744 32512 332750 32564
rect 161014 32444 161020 32496
rect 161072 32484 161078 32496
rect 372614 32484 372620 32496
rect 161072 32456 372620 32484
rect 161072 32444 161078 32456
rect 372614 32444 372620 32456
rect 372672 32444 372678 32496
rect 165706 32376 165712 32428
rect 165764 32416 165770 32428
rect 438854 32416 438860 32428
rect 165764 32388 438860 32416
rect 165764 32376 165770 32388
rect 438854 32376 438860 32388
rect 438912 32376 438918 32428
rect 149974 31288 149980 31340
rect 150032 31328 150038 31340
rect 222194 31328 222200 31340
rect 150032 31300 222200 31328
rect 150032 31288 150038 31300
rect 222194 31288 222200 31300
rect 222252 31288 222258 31340
rect 152274 31220 152280 31272
rect 152332 31260 152338 31272
rect 264974 31260 264980 31272
rect 152332 31232 264980 31260
rect 152332 31220 152338 31232
rect 264974 31220 264980 31232
rect 265032 31220 265038 31272
rect 159634 31152 159640 31204
rect 159692 31192 159698 31204
rect 346394 31192 346400 31204
rect 159692 31164 346400 31192
rect 159692 31152 159698 31164
rect 346394 31152 346400 31164
rect 346452 31152 346458 31204
rect 162210 31084 162216 31136
rect 162268 31124 162274 31136
rect 390646 31124 390652 31136
rect 162268 31096 390652 31124
rect 162268 31084 162274 31096
rect 390646 31084 390652 31096
rect 390704 31084 390710 31136
rect 42794 31016 42800 31068
rect 42852 31056 42858 31068
rect 136542 31056 136548 31068
rect 42852 31028 136548 31056
rect 42852 31016 42858 31028
rect 136542 31016 136548 31028
rect 136600 31016 136606 31068
rect 145558 31016 145564 31068
rect 145616 31056 145622 31068
rect 164878 31056 164884 31068
rect 145616 31028 164884 31056
rect 145616 31016 145622 31028
rect 164878 31016 164884 31028
rect 164936 31016 164942 31068
rect 169570 31016 169576 31068
rect 169628 31056 169634 31068
rect 470594 31056 470600 31068
rect 169628 31028 470600 31056
rect 169628 31016 169634 31028
rect 470594 31016 470600 31028
rect 470652 31016 470658 31068
rect 144270 30268 144276 30320
rect 144328 30308 144334 30320
rect 145098 30308 145104 30320
rect 144328 30280 145104 30308
rect 144328 30268 144334 30280
rect 145098 30268 145104 30280
rect 145156 30268 145162 30320
rect 155218 29860 155224 29912
rect 155276 29900 155282 29912
rect 299566 29900 299572 29912
rect 155276 29872 299572 29900
rect 155276 29860 155282 29872
rect 299566 29860 299572 29872
rect 299624 29860 299630 29912
rect 163958 29792 163964 29844
rect 164016 29832 164022 29844
rect 398926 29832 398932 29844
rect 164016 29804 398932 29832
rect 164016 29792 164022 29804
rect 398926 29792 398932 29804
rect 398984 29792 398990 29844
rect 170766 29724 170772 29776
rect 170824 29764 170830 29776
rect 491294 29764 491300 29776
rect 170824 29736 491300 29764
rect 170824 29724 170830 29736
rect 491294 29724 491300 29736
rect 491352 29724 491358 29776
rect 145926 29656 145932 29708
rect 145984 29696 145990 29708
rect 175918 29696 175924 29708
rect 145984 29668 175924 29696
rect 145984 29656 145990 29668
rect 175918 29656 175924 29668
rect 175976 29656 175982 29708
rect 176470 29656 176476 29708
rect 176528 29696 176534 29708
rect 553394 29696 553400 29708
rect 176528 29668 553400 29696
rect 176528 29656 176534 29668
rect 553394 29656 553400 29668
rect 553452 29656 553458 29708
rect 175458 29588 175464 29640
rect 175516 29628 175522 29640
rect 567930 29628 567936 29640
rect 175516 29600 567936 29628
rect 175516 29588 175522 29600
rect 567930 29588 567936 29600
rect 567988 29588 567994 29640
rect 158438 28432 158444 28484
rect 158496 28472 158502 28484
rect 321554 28472 321560 28484
rect 158496 28444 321560 28472
rect 158496 28432 158502 28444
rect 321554 28432 321560 28444
rect 321612 28432 321618 28484
rect 165154 28364 165160 28416
rect 165212 28404 165218 28416
rect 420914 28404 420920 28416
rect 165212 28376 420920 28404
rect 165212 28364 165218 28376
rect 420914 28364 420920 28376
rect 420972 28364 420978 28416
rect 172238 28296 172244 28348
rect 172296 28336 172302 28348
rect 502334 28336 502340 28348
rect 172296 28308 502340 28336
rect 172296 28296 172302 28308
rect 502334 28296 502340 28308
rect 502392 28296 502398 28348
rect 177758 28228 177764 28280
rect 177816 28268 177822 28280
rect 518894 28268 518900 28280
rect 177816 28240 518900 28268
rect 177816 28228 177822 28240
rect 518894 28228 518900 28240
rect 518952 28228 518958 28280
rect 154206 27140 154212 27192
rect 154264 27180 154270 27192
rect 271874 27180 271880 27192
rect 154264 27152 271880 27180
rect 154264 27140 154270 27152
rect 271874 27140 271880 27152
rect 271932 27140 271938 27192
rect 161106 27072 161112 27124
rect 161164 27112 161170 27124
rect 360194 27112 360200 27124
rect 161164 27084 360200 27112
rect 161164 27072 161170 27084
rect 360194 27072 360200 27084
rect 360252 27072 360258 27124
rect 162302 27004 162308 27056
rect 162360 27044 162366 27056
rect 386414 27044 386420 27056
rect 162360 27016 386420 27044
rect 162360 27004 162366 27016
rect 386414 27004 386420 27016
rect 386472 27004 386478 27056
rect 170858 26936 170864 26988
rect 170916 26976 170922 26988
rect 492674 26976 492680 26988
rect 170916 26948 492680 26976
rect 170916 26936 170922 26948
rect 492674 26936 492680 26948
rect 492732 26936 492738 26988
rect 46198 26868 46204 26920
rect 46256 26908 46262 26920
rect 135714 26908 135720 26920
rect 46256 26880 135720 26908
rect 46256 26868 46262 26880
rect 135714 26868 135720 26880
rect 135772 26868 135778 26920
rect 172330 26868 172336 26920
rect 172388 26908 172394 26920
rect 506566 26908 506572 26920
rect 172388 26880 506572 26908
rect 172388 26868 172394 26880
rect 506566 26868 506572 26880
rect 506624 26868 506630 26920
rect 154022 25712 154028 25764
rect 154080 25752 154086 25764
rect 278774 25752 278780 25764
rect 154080 25724 278780 25752
rect 154080 25712 154086 25724
rect 278774 25712 278780 25724
rect 278832 25712 278838 25764
rect 162394 25644 162400 25696
rect 162452 25684 162458 25696
rect 374086 25684 374092 25696
rect 162452 25656 374092 25684
rect 162452 25644 162458 25656
rect 374086 25644 374092 25656
rect 374144 25644 374150 25696
rect 172422 25576 172428 25628
rect 172480 25616 172486 25628
rect 509234 25616 509240 25628
rect 172480 25588 509240 25616
rect 172480 25576 172486 25588
rect 509234 25576 509240 25588
rect 509292 25576 509298 25628
rect 145006 25508 145012 25560
rect 145064 25548 145070 25560
rect 171778 25548 171784 25560
rect 145064 25520 171784 25548
rect 145064 25508 145070 25520
rect 171778 25508 171784 25520
rect 171836 25508 171842 25560
rect 172146 25508 172152 25560
rect 172204 25548 172210 25560
rect 510614 25548 510620 25560
rect 172204 25520 510620 25548
rect 172204 25508 172210 25520
rect 510614 25508 510620 25520
rect 510672 25508 510678 25560
rect 163866 24216 163872 24268
rect 163924 24256 163930 24268
rect 391934 24256 391940 24268
rect 163924 24228 391940 24256
rect 163924 24216 163930 24228
rect 391934 24216 391940 24228
rect 391992 24216 391998 24268
rect 171134 24148 171140 24200
rect 171192 24188 171198 24200
rect 513374 24188 513380 24200
rect 171192 24160 513380 24188
rect 171192 24148 171198 24160
rect 513374 24148 513380 24160
rect 513432 24148 513438 24200
rect 173618 24080 173624 24132
rect 173676 24120 173682 24132
rect 531406 24120 531412 24132
rect 173676 24092 531412 24120
rect 173676 24080 173682 24092
rect 531406 24080 531412 24092
rect 531464 24080 531470 24132
rect 153838 22992 153844 23044
rect 153896 23032 153902 23044
rect 282914 23032 282920 23044
rect 153896 23004 282920 23032
rect 153896 22992 153902 23004
rect 282914 22992 282920 23004
rect 282972 22992 282978 23044
rect 162486 22924 162492 22976
rect 162544 22964 162550 22976
rect 382274 22964 382280 22976
rect 162544 22936 382280 22964
rect 162544 22924 162550 22936
rect 382274 22924 382280 22936
rect 382332 22924 382338 22976
rect 163774 22856 163780 22908
rect 163832 22896 163838 22908
rect 404354 22896 404360 22908
rect 163832 22868 404360 22896
rect 163832 22856 163838 22868
rect 404354 22856 404360 22868
rect 404412 22856 404418 22908
rect 173710 22788 173716 22840
rect 173768 22828 173774 22840
rect 520274 22828 520280 22840
rect 173768 22800 520280 22828
rect 173768 22788 173774 22800
rect 520274 22788 520280 22800
rect 520332 22788 520338 22840
rect 173802 22720 173808 22772
rect 173860 22760 173866 22772
rect 524414 22760 524420 22772
rect 173860 22732 524420 22760
rect 173860 22720 173866 22732
rect 524414 22720 524420 22732
rect 524472 22720 524478 22772
rect 159726 21428 159732 21480
rect 159784 21468 159790 21480
rect 350534 21468 350540 21480
rect 159784 21440 350540 21468
rect 159784 21428 159790 21440
rect 350534 21428 350540 21440
rect 350592 21428 350598 21480
rect 165338 21360 165344 21412
rect 165396 21400 165402 21412
rect 418154 21400 418160 21412
rect 165396 21372 418160 21400
rect 165396 21360 165402 21372
rect 418154 21360 418160 21372
rect 418212 21360 418218 21412
rect 155862 20068 155868 20120
rect 155920 20108 155926 20120
rect 287054 20108 287060 20120
rect 155920 20080 287060 20108
rect 155920 20068 155926 20080
rect 287054 20068 287060 20080
rect 287112 20068 287118 20120
rect 155770 20000 155776 20052
rect 155828 20040 155834 20052
rect 291194 20040 291200 20052
rect 155828 20012 291200 20040
rect 155828 20000 155834 20012
rect 291194 20000 291200 20012
rect 291252 20000 291258 20052
rect 143626 19932 143632 19984
rect 143684 19972 143690 19984
rect 154574 19972 154580 19984
rect 143684 19944 154580 19972
rect 143684 19932 143690 19944
rect 154574 19932 154580 19944
rect 154632 19932 154638 19984
rect 161198 19932 161204 19984
rect 161256 19972 161262 19984
rect 361574 19972 361580 19984
rect 161256 19944 361580 19972
rect 161256 19932 161262 19944
rect 361574 19932 361580 19944
rect 361632 19932 361638 19984
rect 152826 18844 152832 18896
rect 152884 18884 152890 18896
rect 251266 18884 251272 18896
rect 152884 18856 251272 18884
rect 152884 18844 152890 18856
rect 251266 18844 251272 18856
rect 251324 18844 251330 18896
rect 159818 18776 159824 18828
rect 159876 18816 159882 18828
rect 345014 18816 345020 18828
rect 159876 18788 345020 18816
rect 159876 18776 159882 18788
rect 345014 18776 345020 18788
rect 345072 18776 345078 18828
rect 165246 18708 165252 18760
rect 165304 18748 165310 18760
rect 411254 18748 411260 18760
rect 165304 18720 411260 18748
rect 165304 18708 165310 18720
rect 411254 18708 411260 18720
rect 411312 18708 411318 18760
rect 177850 18640 177856 18692
rect 177908 18680 177914 18692
rect 571334 18680 571340 18692
rect 177908 18652 571340 18680
rect 177908 18640 177914 18652
rect 571334 18640 571340 18652
rect 571392 18640 571398 18692
rect 177942 18572 177948 18624
rect 178000 18612 178006 18624
rect 574094 18612 574100 18624
rect 178000 18584 574100 18612
rect 178000 18572 178006 18584
rect 574094 18572 574100 18584
rect 574152 18572 574158 18624
rect 152642 17416 152648 17468
rect 152700 17456 152706 17468
rect 259546 17456 259552 17468
rect 152700 17428 259552 17456
rect 152700 17416 152706 17428
rect 259546 17416 259552 17428
rect 259604 17416 259610 17468
rect 167914 17348 167920 17400
rect 167972 17388 167978 17400
rect 445754 17388 445760 17400
rect 167972 17360 445760 17388
rect 167972 17348 167978 17360
rect 445754 17348 445760 17360
rect 445812 17348 445818 17400
rect 168006 17280 168012 17332
rect 168064 17320 168070 17332
rect 448606 17320 448612 17332
rect 168064 17292 448612 17320
rect 168064 17280 168070 17292
rect 448606 17280 448612 17292
rect 448664 17280 448670 17332
rect 146018 17212 146024 17264
rect 146076 17252 146082 17264
rect 166994 17252 167000 17264
rect 146076 17224 167000 17252
rect 146076 17212 146082 17224
rect 166994 17212 167000 17224
rect 167052 17212 167058 17264
rect 169662 17212 169668 17264
rect 169720 17252 169726 17264
rect 477494 17252 477500 17264
rect 169720 17224 477500 17252
rect 169720 17212 169726 17224
rect 477494 17212 477500 17224
rect 477552 17212 477558 17264
rect 154390 16124 154396 16176
rect 154448 16164 154454 16176
rect 284386 16164 284392 16176
rect 154448 16136 284392 16164
rect 154448 16124 154454 16136
rect 284386 16124 284392 16136
rect 284444 16124 284450 16176
rect 160094 16056 160100 16108
rect 160152 16096 160158 16108
rect 364610 16096 364616 16108
rect 160152 16068 364616 16096
rect 160152 16056 160158 16068
rect 364610 16056 364616 16068
rect 364668 16056 364674 16108
rect 165430 15988 165436 16040
rect 165488 16028 165494 16040
rect 417418 16028 417424 16040
rect 165488 16000 417424 16028
rect 165488 15988 165494 16000
rect 417418 15988 417424 16000
rect 417476 15988 417482 16040
rect 166718 15920 166724 15972
rect 166776 15960 166782 15972
rect 440326 15960 440332 15972
rect 166776 15932 440332 15960
rect 166776 15920 166782 15932
rect 440326 15920 440332 15932
rect 440384 15920 440390 15972
rect 174998 15852 175004 15904
rect 175056 15892 175062 15904
rect 546494 15892 546500 15904
rect 175056 15864 546500 15892
rect 175056 15852 175062 15864
rect 546494 15852 546500 15864
rect 546552 15852 546558 15904
rect 154298 14696 154304 14748
rect 154356 14736 154362 14748
rect 276014 14736 276020 14748
rect 154356 14708 276020 14736
rect 154356 14696 154362 14708
rect 276014 14696 276020 14708
rect 276072 14696 276078 14748
rect 157242 14628 157248 14680
rect 157300 14668 157306 14680
rect 314654 14668 314660 14680
rect 157300 14640 314660 14668
rect 157300 14628 157306 14640
rect 314654 14628 314660 14640
rect 314712 14628 314718 14680
rect 168098 14560 168104 14612
rect 168156 14600 168162 14612
rect 382366 14600 382372 14612
rect 168156 14572 382372 14600
rect 168156 14560 168162 14572
rect 382366 14560 382372 14572
rect 382424 14560 382430 14612
rect 162670 14492 162676 14544
rect 162728 14532 162734 14544
rect 385954 14532 385960 14544
rect 162728 14504 385960 14532
rect 162728 14492 162734 14504
rect 385954 14492 385960 14504
rect 386012 14492 386018 14544
rect 170950 14424 170956 14476
rect 171008 14464 171014 14476
rect 486418 14464 486424 14476
rect 171008 14436 486424 14464
rect 171008 14424 171014 14436
rect 486418 14424 486424 14436
rect 486476 14424 486482 14476
rect 152550 13336 152556 13388
rect 152608 13376 152614 13388
rect 258258 13376 258264 13388
rect 152608 13348 258264 13376
rect 152608 13336 152614 13348
rect 258258 13336 258264 13348
rect 258316 13336 258322 13388
rect 156690 13268 156696 13320
rect 156748 13308 156754 13320
rect 307938 13308 307944 13320
rect 156748 13280 307944 13308
rect 156748 13268 156754 13280
rect 307938 13268 307944 13280
rect 307996 13268 308002 13320
rect 164050 13200 164056 13252
rect 164108 13240 164114 13252
rect 376018 13240 376024 13252
rect 164108 13212 376024 13240
rect 164108 13200 164114 13212
rect 376018 13200 376024 13212
rect 376076 13200 376082 13252
rect 162578 13132 162584 13184
rect 162636 13172 162642 13184
rect 378410 13172 378416 13184
rect 162636 13144 378416 13172
rect 162636 13132 162642 13144
rect 378410 13132 378416 13144
rect 378468 13132 378474 13184
rect 171042 13064 171048 13116
rect 171100 13104 171106 13116
rect 482186 13104 482192 13116
rect 171100 13076 482192 13104
rect 171100 13064 171106 13076
rect 482186 13064 482192 13076
rect 482244 13064 482250 13116
rect 149790 11976 149796 12028
rect 149848 12016 149854 12028
rect 226334 12016 226340 12028
rect 149848 11988 226340 12016
rect 149848 11976 149854 11988
rect 226334 11976 226340 11988
rect 226392 11976 226398 12028
rect 158530 11908 158536 11960
rect 158588 11948 158594 11960
rect 328730 11948 328736 11960
rect 158588 11920 328736 11948
rect 158588 11908 158594 11920
rect 328730 11908 328736 11920
rect 328788 11908 328794 11960
rect 164142 11840 164148 11892
rect 164200 11880 164206 11892
rect 407206 11880 407212 11892
rect 164200 11852 407212 11880
rect 164200 11840 164206 11852
rect 407206 11840 407212 11852
rect 407264 11840 407270 11892
rect 168190 11772 168196 11824
rect 168248 11812 168254 11824
rect 454034 11812 454040 11824
rect 168248 11784 454040 11812
rect 168248 11772 168254 11784
rect 454034 11772 454040 11784
rect 454092 11772 454098 11824
rect 175366 11704 175372 11756
rect 175424 11744 175430 11756
rect 560386 11744 560392 11756
rect 175424 11716 560392 11744
rect 175424 11704 175430 11716
rect 560386 11704 560392 11716
rect 560444 11704 560450 11756
rect 184934 11636 184940 11688
rect 184992 11676 184998 11688
rect 186130 11676 186136 11688
rect 184992 11648 186136 11676
rect 184992 11636 184998 11648
rect 186130 11636 186136 11648
rect 186188 11636 186194 11688
rect 201494 11636 201500 11688
rect 201552 11676 201558 11688
rect 202690 11676 202696 11688
rect 201552 11648 202696 11676
rect 201552 11636 201558 11648
rect 202690 11636 202696 11648
rect 202748 11636 202754 11688
rect 234614 11636 234620 11688
rect 234672 11676 234678 11688
rect 235810 11676 235816 11688
rect 234672 11648 235816 11676
rect 234672 11636 234678 11648
rect 235810 11636 235816 11648
rect 235868 11636 235874 11688
rect 151170 10548 151176 10600
rect 151228 10588 151234 10600
rect 234614 10588 234620 10600
rect 151228 10560 234620 10588
rect 151228 10548 151234 10560
rect 234614 10548 234620 10560
rect 234672 10548 234678 10600
rect 158622 10480 158628 10532
rect 158680 10520 158686 10532
rect 336274 10520 336280 10532
rect 158680 10492 336280 10520
rect 158680 10480 158686 10492
rect 336274 10480 336280 10492
rect 336332 10480 336338 10532
rect 161290 10412 161296 10464
rect 161348 10452 161354 10464
rect 365806 10452 365812 10464
rect 161348 10424 365812 10452
rect 161348 10412 161354 10424
rect 365806 10412 365812 10424
rect 365864 10412 365870 10464
rect 166810 10344 166816 10396
rect 166868 10384 166874 10396
rect 432046 10384 432052 10396
rect 166868 10356 432052 10384
rect 166868 10344 166874 10356
rect 432046 10344 432052 10356
rect 432104 10344 432110 10396
rect 30098 10276 30104 10328
rect 30156 10316 30162 10328
rect 133966 10316 133972 10328
rect 30156 10288 133972 10316
rect 30156 10276 30162 10288
rect 133966 10276 133972 10288
rect 134024 10276 134030 10328
rect 175090 10276 175096 10328
rect 175148 10316 175154 10328
rect 548610 10316 548616 10328
rect 175148 10288 548616 10316
rect 175148 10276 175154 10288
rect 548610 10276 548616 10288
rect 548668 10276 548674 10328
rect 149882 9188 149888 9240
rect 149940 9228 149946 9240
rect 227530 9228 227536 9240
rect 149940 9200 227536 9228
rect 149940 9188 149946 9200
rect 227530 9188 227536 9200
rect 227588 9188 227594 9240
rect 156598 9120 156604 9172
rect 156656 9160 156662 9172
rect 316218 9160 316224 9172
rect 156656 9132 316224 9160
rect 156656 9120 156662 9132
rect 316218 9120 316224 9132
rect 316276 9120 316282 9172
rect 165522 9052 165528 9104
rect 165580 9092 165586 9104
rect 414290 9092 414296 9104
rect 165580 9064 414296 9092
rect 165580 9052 165586 9064
rect 414290 9052 414296 9064
rect 414348 9052 414354 9104
rect 184198 8984 184204 9036
rect 184256 9024 184262 9036
rect 562042 9024 562048 9036
rect 184256 8996 562048 9024
rect 184256 8984 184262 8996
rect 562042 8984 562048 8996
rect 562100 8984 562106 9036
rect 6454 8916 6460 8968
rect 6512 8956 6518 8968
rect 132586 8956 132592 8968
rect 6512 8928 132592 8956
rect 6512 8916 6518 8928
rect 132586 8916 132592 8928
rect 132644 8916 132650 8968
rect 175274 8916 175280 8968
rect 175332 8956 175338 8968
rect 556154 8956 556160 8968
rect 175332 8928 556160 8956
rect 175332 8916 175338 8928
rect 556154 8916 556160 8928
rect 556212 8916 556218 8968
rect 151262 7828 151268 7880
rect 151320 7868 151326 7880
rect 241698 7868 241704 7880
rect 151320 7840 241704 7868
rect 151320 7828 151326 7840
rect 241698 7828 241704 7840
rect 241756 7828 241762 7880
rect 160002 7760 160008 7812
rect 160060 7800 160066 7812
rect 343358 7800 343364 7812
rect 160060 7772 343364 7800
rect 160060 7760 160066 7772
rect 343358 7760 343364 7772
rect 343416 7760 343422 7812
rect 162762 7692 162768 7744
rect 162820 7732 162826 7744
rect 379974 7732 379980 7744
rect 162820 7704 379980 7732
rect 162820 7692 162826 7704
rect 379974 7692 379980 7704
rect 380032 7692 380038 7744
rect 166902 7624 166908 7676
rect 166960 7664 166966 7676
rect 435542 7664 435548 7676
rect 166960 7636 435548 7664
rect 166960 7624 166966 7636
rect 435542 7624 435548 7636
rect 435600 7624 435606 7676
rect 103330 7556 103336 7608
rect 103388 7596 103394 7608
rect 139578 7596 139584 7608
rect 103388 7568 139584 7596
rect 103388 7556 103394 7568
rect 139578 7556 139584 7568
rect 139636 7556 139642 7608
rect 175182 7556 175188 7608
rect 175240 7596 175246 7608
rect 538398 7596 538404 7608
rect 175240 7568 538404 7596
rect 175240 7556 175246 7568
rect 538398 7556 538404 7568
rect 538456 7556 538462 7608
rect 3418 6808 3424 6860
rect 3476 6848 3482 6860
rect 21358 6848 21364 6860
rect 3476 6820 21364 6848
rect 3476 6808 3482 6820
rect 21358 6808 21364 6820
rect 21416 6808 21422 6860
rect 154482 6740 154488 6792
rect 154540 6780 154546 6792
rect 273622 6780 273628 6792
rect 154540 6752 273628 6780
rect 154540 6740 154546 6752
rect 273622 6740 273628 6752
rect 273680 6740 273686 6792
rect 159910 6672 159916 6724
rect 159968 6712 159974 6724
rect 350442 6712 350448 6724
rect 159968 6684 350448 6712
rect 159968 6672 159974 6684
rect 350442 6672 350448 6684
rect 350500 6672 350506 6724
rect 180702 6604 180708 6656
rect 180760 6644 180766 6656
rect 422570 6644 422576 6656
rect 180760 6616 422576 6644
rect 180760 6604 180766 6616
rect 422570 6604 422576 6616
rect 422628 6604 422634 6656
rect 181990 6536 181996 6588
rect 182048 6576 182054 6588
rect 429654 6576 429660 6588
rect 182048 6548 429660 6576
rect 182048 6536 182054 6548
rect 429654 6536 429660 6548
rect 429712 6536 429718 6588
rect 180610 6468 180616 6520
rect 180668 6508 180674 6520
rect 436738 6508 436744 6520
rect 180668 6480 436744 6508
rect 180668 6468 180674 6480
rect 436738 6468 436744 6480
rect 436796 6468 436802 6520
rect 179138 6400 179144 6452
rect 179196 6440 179202 6452
rect 443822 6440 443828 6452
rect 179196 6412 443828 6440
rect 179196 6400 179202 6412
rect 443822 6400 443828 6412
rect 443880 6400 443886 6452
rect 181898 6332 181904 6384
rect 181956 6372 181962 6384
rect 450906 6372 450912 6384
rect 181956 6344 450912 6372
rect 181956 6332 181962 6344
rect 450906 6332 450912 6344
rect 450964 6332 450970 6384
rect 165614 6264 165620 6316
rect 165672 6304 165678 6316
rect 442626 6304 442632 6316
rect 165672 6276 442632 6304
rect 165672 6264 165678 6276
rect 442626 6264 442632 6276
rect 442684 6264 442690 6316
rect 176562 6196 176568 6248
rect 176620 6236 176626 6248
rect 563238 6236 563244 6248
rect 176620 6208 563244 6236
rect 176620 6196 176626 6208
rect 563238 6196 563244 6208
rect 563296 6196 563302 6248
rect 87966 6128 87972 6180
rect 88024 6168 88030 6180
rect 138198 6168 138204 6180
rect 88024 6140 138204 6168
rect 88024 6128 88030 6140
rect 138198 6128 138204 6140
rect 138256 6128 138262 6180
rect 144178 6128 144184 6180
rect 144236 6168 144242 6180
rect 161290 6168 161296 6180
rect 144236 6140 161296 6168
rect 144236 6128 144242 6140
rect 161290 6128 161296 6140
rect 161348 6128 161354 6180
rect 182082 6128 182088 6180
rect 182140 6168 182146 6180
rect 583386 6168 583392 6180
rect 182140 6140 583392 6168
rect 182140 6128 182146 6140
rect 583386 6128 583392 6140
rect 583444 6128 583450 6180
rect 143534 5652 143540 5704
rect 143592 5692 143598 5704
rect 144730 5692 144736 5704
rect 143592 5664 144736 5692
rect 143592 5652 143598 5664
rect 144730 5652 144736 5664
rect 144788 5652 144794 5704
rect 138842 5516 138848 5568
rect 138900 5556 138906 5568
rect 142522 5556 142528 5568
rect 138900 5528 142528 5556
rect 138900 5516 138906 5528
rect 142522 5516 142528 5528
rect 142580 5516 142586 5568
rect 142798 5516 142804 5568
rect 142856 5556 142862 5568
rect 143534 5556 143540 5568
rect 142856 5528 143540 5556
rect 142856 5516 142862 5528
rect 143534 5516 143540 5528
rect 143592 5516 143598 5568
rect 151078 4972 151084 5024
rect 151136 5012 151142 5024
rect 245194 5012 245200 5024
rect 151136 4984 245200 5012
rect 151136 4972 151142 4984
rect 245194 4972 245200 4984
rect 245252 4972 245258 5024
rect 161382 4904 161388 4956
rect 161440 4944 161446 4956
rect 371694 4944 371700 4956
rect 161440 4916 371700 4944
rect 161440 4904 161446 4916
rect 371694 4904 371700 4916
rect 371752 4904 371758 4956
rect 168282 4836 168288 4888
rect 168340 4876 168346 4888
rect 456886 4876 456892 4888
rect 168340 4848 456892 4876
rect 168340 4836 168346 4848
rect 456886 4836 456892 4848
rect 456944 4836 456950 4888
rect 25314 4768 25320 4820
rect 25372 4808 25378 4820
rect 133874 4808 133880 4820
rect 25372 4780 133880 4808
rect 25372 4768 25378 4780
rect 133874 4768 133880 4780
rect 133932 4768 133938 4820
rect 173894 4768 173900 4820
rect 173952 4808 173958 4820
rect 541986 4808 541992 4820
rect 173952 4780 541992 4808
rect 173952 4768 173958 4780
rect 541986 4768 541992 4780
rect 542044 4768 542050 4820
rect 566 4088 572 4140
rect 624 4128 630 4140
rect 7558 4128 7564 4140
rect 624 4100 7564 4128
rect 624 4088 630 4100
rect 7558 4088 7564 4100
rect 7616 4088 7622 4140
rect 73798 4088 73804 4140
rect 73856 4128 73862 4140
rect 75178 4128 75184 4140
rect 73856 4100 75184 4128
rect 73856 4088 73862 4100
rect 75178 4088 75184 4100
rect 75236 4088 75242 4140
rect 83274 4088 83280 4140
rect 83332 4128 83338 4140
rect 84838 4128 84844 4140
rect 83332 4100 84844 4128
rect 83332 4088 83338 4100
rect 84838 4088 84844 4100
rect 84896 4088 84902 4140
rect 112806 4088 112812 4140
rect 112864 4128 112870 4140
rect 113266 4128 113272 4140
rect 112864 4100 113272 4128
rect 112864 4088 112870 4100
rect 113266 4088 113272 4100
rect 113324 4088 113330 4140
rect 148318 4088 148324 4140
rect 148376 4128 148382 4140
rect 154206 4128 154212 4140
rect 148376 4100 154212 4128
rect 148376 4088 148382 4100
rect 154206 4088 154212 4100
rect 154264 4088 154270 4140
rect 181806 4088 181812 4140
rect 181864 4128 181870 4140
rect 187418 4128 187424 4140
rect 181864 4100 187424 4128
rect 181864 4088 181870 4100
rect 187418 4088 187424 4100
rect 187476 4088 187482 4140
rect 188338 4088 188344 4140
rect 188396 4128 188402 4140
rect 196802 4128 196808 4140
rect 188396 4100 196808 4128
rect 188396 4088 188402 4100
rect 196802 4088 196808 4100
rect 196860 4088 196866 4140
rect 197262 4088 197268 4140
rect 197320 4128 197326 4140
rect 203886 4128 203892 4140
rect 197320 4100 203892 4128
rect 197320 4088 197326 4100
rect 203886 4088 203892 4100
rect 203944 4088 203950 4140
rect 207658 4088 207664 4140
rect 207716 4128 207722 4140
rect 210970 4128 210976 4140
rect 207716 4100 210976 4128
rect 207716 4088 207722 4100
rect 210970 4088 210976 4100
rect 211028 4088 211034 4140
rect 211798 4088 211804 4140
rect 211856 4128 211862 4140
rect 223942 4128 223948 4140
rect 211856 4100 223948 4128
rect 211856 4088 211862 4100
rect 223942 4088 223948 4100
rect 224000 4088 224006 4140
rect 242158 4088 242164 4140
rect 242216 4128 242222 4140
rect 260650 4128 260656 4140
rect 242216 4100 260656 4128
rect 242216 4088 242222 4100
rect 260650 4088 260656 4100
rect 260708 4088 260714 4140
rect 315298 4088 315304 4140
rect 315356 4128 315362 4140
rect 317322 4128 317328 4140
rect 315356 4100 317328 4128
rect 315356 4088 315362 4100
rect 317322 4088 317328 4100
rect 317380 4088 317386 4140
rect 323578 4088 323584 4140
rect 323636 4128 323642 4140
rect 326798 4128 326804 4140
rect 323636 4100 326804 4128
rect 323636 4088 323642 4100
rect 326798 4088 326804 4100
rect 326856 4088 326862 4140
rect 450538 4088 450544 4140
rect 450596 4128 450602 4140
rect 452102 4128 452108 4140
rect 450596 4100 452108 4128
rect 450596 4088 450602 4100
rect 452102 4088 452108 4100
rect 452160 4088 452166 4140
rect 180058 4020 180064 4072
rect 180116 4060 180122 4072
rect 189810 4060 189816 4072
rect 180116 4032 189816 4060
rect 180116 4020 180122 4032
rect 189810 4020 189816 4032
rect 189868 4020 189874 4072
rect 193858 4020 193864 4072
rect 193916 4060 193922 4072
rect 195606 4060 195612 4072
rect 193916 4032 195612 4060
rect 193916 4020 193922 4032
rect 195606 4020 195612 4032
rect 195664 4020 195670 4072
rect 195698 4020 195704 4072
rect 195756 4060 195762 4072
rect 247586 4060 247592 4072
rect 195756 4032 247592 4060
rect 195756 4020 195762 4032
rect 247586 4020 247592 4032
rect 247644 4020 247650 4072
rect 284294 4020 284300 4072
rect 284352 4060 284358 4072
rect 285030 4060 285036 4072
rect 284352 4032 285036 4060
rect 284352 4020 284358 4032
rect 285030 4020 285036 4032
rect 285088 4020 285094 4072
rect 287698 4020 287704 4072
rect 287756 4060 287762 4072
rect 312630 4060 312636 4072
rect 287756 4032 312636 4060
rect 287756 4020 287762 4032
rect 312630 4020 312636 4032
rect 312688 4020 312694 4072
rect 566458 4020 566464 4072
rect 566516 4060 566522 4072
rect 568022 4060 568028 4072
rect 566516 4032 568028 4060
rect 566516 4020 566522 4032
rect 568022 4020 568028 4032
rect 568080 4020 568086 4072
rect 146938 3952 146944 4004
rect 146996 3992 147002 4004
rect 148502 3992 148508 4004
rect 146996 3964 148508 3992
rect 146996 3952 147002 3964
rect 148502 3952 148508 3964
rect 148560 3952 148566 4004
rect 149698 3952 149704 4004
rect 149756 3992 149762 4004
rect 153010 3992 153016 4004
rect 149756 3964 153016 3992
rect 149756 3952 149762 3964
rect 153010 3952 153016 3964
rect 153068 3952 153074 4004
rect 182818 3952 182824 4004
rect 182876 3992 182882 4004
rect 212166 3992 212172 4004
rect 182876 3964 212172 3992
rect 182876 3952 182882 3964
rect 212166 3952 212172 3964
rect 212224 3952 212230 4004
rect 220078 3952 220084 4004
rect 220136 3992 220142 4004
rect 298462 3992 298468 4004
rect 220136 3964 298468 3992
rect 220136 3952 220142 3964
rect 298462 3952 298468 3964
rect 298520 3952 298526 4004
rect 299566 3952 299572 4004
rect 299624 3992 299630 4004
rect 300762 3992 300768 4004
rect 299624 3964 300768 3992
rect 299624 3952 299630 3964
rect 300762 3952 300768 3964
rect 300820 3952 300826 4004
rect 147122 3884 147128 3936
rect 147180 3924 147186 3936
rect 149606 3924 149612 3936
rect 147180 3896 149612 3924
rect 147180 3884 147186 3896
rect 149606 3884 149612 3896
rect 149664 3884 149670 3936
rect 179230 3884 179236 3936
rect 179288 3924 179294 3936
rect 394234 3924 394240 3936
rect 179288 3896 394240 3924
rect 179288 3884 179294 3896
rect 394234 3884 394240 3896
rect 394292 3884 394298 3936
rect 44266 3816 44272 3868
rect 44324 3856 44330 3868
rect 46198 3856 46204 3868
rect 44324 3828 46204 3856
rect 44324 3816 44330 3828
rect 46198 3816 46204 3828
rect 46256 3816 46262 3868
rect 148410 3816 148416 3868
rect 148468 3856 148474 3868
rect 163682 3856 163688 3868
rect 148468 3828 163688 3856
rect 148468 3816 148474 3828
rect 163682 3816 163688 3828
rect 163740 3816 163746 3868
rect 179322 3816 179328 3868
rect 179380 3856 179386 3868
rect 401318 3856 401324 3868
rect 179380 3828 401324 3856
rect 179380 3816 179386 3828
rect 401318 3816 401324 3828
rect 401376 3816 401382 3868
rect 122282 3748 122288 3800
rect 122340 3788 122346 3800
rect 127066 3788 127072 3800
rect 122340 3760 127072 3788
rect 122340 3748 122346 3760
rect 127066 3748 127072 3760
rect 127124 3748 127130 3800
rect 130838 3748 130844 3800
rect 130896 3788 130902 3800
rect 151814 3788 151820 3800
rect 130896 3760 151820 3788
rect 130896 3748 130902 3760
rect 151814 3748 151820 3760
rect 151872 3748 151878 3800
rect 152458 3748 152464 3800
rect 152516 3788 152522 3800
rect 164510 3788 164516 3800
rect 152516 3760 164516 3788
rect 152516 3748 152522 3760
rect 164510 3748 164516 3760
rect 164568 3748 164574 3800
rect 178770 3748 178776 3800
rect 178828 3788 178834 3800
rect 408402 3788 408408 3800
rect 178828 3760 408408 3788
rect 178828 3748 178834 3760
rect 408402 3748 408408 3760
rect 408460 3748 408466 3800
rect 119890 3680 119896 3732
rect 119948 3720 119954 3732
rect 131482 3720 131488 3732
rect 119948 3692 131488 3720
rect 119948 3680 119954 3692
rect 131482 3680 131488 3692
rect 131540 3680 131546 3732
rect 147030 3680 147036 3732
rect 147088 3720 147094 3732
rect 149514 3720 149520 3732
rect 147088 3692 149520 3720
rect 147088 3680 147094 3692
rect 149514 3680 149520 3692
rect 149572 3680 149578 3732
rect 149606 3680 149612 3732
rect 149664 3720 149670 3732
rect 171962 3720 171968 3732
rect 149664 3692 171968 3720
rect 149664 3680 149670 3692
rect 171962 3680 171968 3692
rect 172020 3680 172026 3732
rect 178678 3680 178684 3732
rect 178736 3720 178742 3732
rect 415486 3720 415492 3732
rect 178736 3692 415492 3720
rect 178736 3680 178742 3692
rect 415486 3680 415492 3692
rect 415544 3680 415550 3732
rect 454678 3680 454684 3732
rect 454736 3720 454742 3732
rect 497090 3720 497096 3732
rect 454736 3692 497096 3720
rect 454736 3680 454742 3692
rect 497090 3680 497096 3692
rect 497148 3680 497154 3732
rect 51350 3612 51356 3664
rect 51408 3652 51414 3664
rect 54478 3652 54484 3664
rect 51408 3624 54484 3652
rect 51408 3612 51414 3624
rect 54478 3612 54484 3624
rect 54536 3612 54542 3664
rect 65518 3612 65524 3664
rect 65576 3652 65582 3664
rect 65576 3624 74534 3652
rect 65576 3612 65582 3624
rect 17034 3544 17040 3596
rect 17092 3584 17098 3596
rect 18598 3584 18604 3596
rect 17092 3556 18604 3584
rect 17092 3544 17098 3556
rect 18598 3544 18604 3556
rect 18656 3544 18662 3596
rect 19426 3544 19432 3596
rect 19484 3584 19490 3596
rect 21450 3584 21456 3596
rect 19484 3556 21456 3584
rect 19484 3544 19490 3556
rect 21450 3544 21456 3556
rect 21508 3544 21514 3596
rect 27614 3544 27620 3596
rect 27672 3584 27678 3596
rect 28534 3584 28540 3596
rect 27672 3556 28540 3584
rect 27672 3544 27678 3556
rect 28534 3544 28540 3556
rect 28592 3544 28598 3596
rect 52454 3544 52460 3596
rect 52512 3584 52518 3596
rect 53374 3584 53380 3596
rect 52512 3556 53380 3584
rect 52512 3544 52518 3556
rect 53374 3544 53380 3556
rect 53432 3544 53438 3596
rect 56042 3544 56048 3596
rect 56100 3584 56106 3596
rect 57238 3584 57244 3596
rect 56100 3556 57244 3584
rect 56100 3544 56106 3556
rect 57238 3544 57244 3556
rect 57296 3544 57302 3596
rect 60734 3544 60740 3596
rect 60792 3584 60798 3596
rect 61654 3584 61660 3596
rect 60792 3556 61660 3584
rect 60792 3544 60798 3556
rect 61654 3544 61660 3556
rect 61712 3544 61718 3596
rect 69106 3544 69112 3596
rect 69164 3584 69170 3596
rect 71038 3584 71044 3596
rect 69164 3556 71044 3584
rect 69164 3544 69170 3556
rect 71038 3544 71044 3556
rect 71096 3544 71102 3596
rect 74506 3584 74534 3624
rect 93946 3612 93952 3664
rect 94004 3652 94010 3664
rect 125594 3652 125600 3664
rect 94004 3624 125600 3652
rect 94004 3612 94010 3624
rect 125594 3612 125600 3624
rect 125652 3612 125658 3664
rect 129826 3652 129832 3664
rect 125796 3624 129832 3652
rect 125796 3584 125824 3624
rect 129826 3612 129832 3624
rect 129884 3612 129890 3664
rect 131022 3612 131028 3664
rect 131080 3652 131086 3664
rect 162486 3652 162492 3664
rect 131080 3624 162492 3652
rect 131080 3612 131086 3624
rect 162486 3612 162492 3624
rect 162544 3612 162550 3664
rect 179046 3612 179052 3664
rect 179104 3652 179110 3664
rect 461578 3652 461584 3664
rect 179104 3624 461584 3652
rect 179104 3612 179110 3624
rect 461578 3612 461584 3624
rect 461636 3612 461642 3664
rect 74506 3556 125824 3584
rect 125870 3544 125876 3596
rect 125928 3584 125934 3596
rect 129918 3584 129924 3596
rect 125928 3556 129924 3584
rect 125928 3544 125934 3556
rect 129918 3544 129924 3556
rect 129976 3544 129982 3596
rect 130930 3544 130936 3596
rect 130988 3584 130994 3596
rect 166074 3584 166080 3596
rect 130988 3556 166080 3584
rect 130988 3544 130994 3556
rect 166074 3544 166080 3556
rect 166132 3544 166138 3596
rect 170398 3544 170404 3596
rect 170456 3584 170462 3596
rect 174262 3584 174268 3596
rect 170456 3556 174268 3584
rect 170456 3544 170462 3556
rect 174262 3544 174268 3556
rect 174320 3544 174326 3596
rect 185578 3544 185584 3596
rect 185636 3584 185642 3596
rect 187326 3584 187332 3596
rect 185636 3556 187332 3584
rect 185636 3544 185642 3556
rect 187326 3544 187332 3556
rect 187384 3544 187390 3596
rect 187418 3544 187424 3596
rect 187476 3584 187482 3596
rect 468294 3584 468300 3596
rect 187476 3556 468300 3584
rect 187476 3544 187482 3556
rect 468294 3544 468300 3556
rect 468352 3544 468358 3596
rect 468478 3544 468484 3596
rect 468536 3584 468542 3596
rect 469858 3584 469864 3596
rect 468536 3556 469864 3584
rect 468536 3544 468542 3556
rect 469858 3544 469864 3556
rect 469916 3544 469922 3596
rect 470566 3556 478184 3584
rect 15930 3476 15936 3528
rect 15988 3516 15994 3528
rect 15988 3488 123432 3516
rect 15988 3476 15994 3488
rect 1670 3408 1676 3460
rect 1728 3448 1734 3460
rect 8938 3448 8944 3460
rect 1728 3420 8944 3448
rect 1728 3408 1734 3420
rect 8938 3408 8944 3420
rect 8996 3408 9002 3460
rect 11146 3408 11152 3460
rect 11204 3448 11210 3460
rect 11204 3420 122834 3448
rect 11204 3408 11210 3420
rect 91554 3340 91560 3392
rect 91612 3380 91618 3392
rect 93118 3380 93124 3392
rect 91612 3352 93124 3380
rect 91612 3340 91618 3352
rect 93118 3340 93124 3352
rect 93176 3340 93182 3392
rect 101030 3340 101036 3392
rect 101088 3380 101094 3392
rect 102778 3380 102784 3392
rect 101088 3352 102784 3380
rect 101088 3340 101094 3352
rect 102778 3340 102784 3352
rect 102836 3340 102842 3392
rect 105722 3340 105728 3392
rect 105780 3380 105786 3392
rect 106918 3380 106924 3392
rect 105780 3352 106924 3380
rect 105780 3340 105786 3352
rect 106918 3340 106924 3352
rect 106976 3340 106982 3392
rect 110414 3340 110420 3392
rect 110472 3380 110478 3392
rect 111610 3380 111616 3392
rect 110472 3352 111616 3380
rect 110472 3340 110478 3352
rect 111610 3340 111616 3352
rect 111668 3340 111674 3392
rect 109310 3272 109316 3324
rect 109368 3312 109374 3324
rect 112438 3312 112444 3324
rect 109368 3284 112444 3312
rect 109368 3272 109374 3284
rect 112438 3272 112444 3284
rect 112496 3272 112502 3324
rect 122806 3312 122834 3420
rect 123404 3380 123432 3488
rect 123478 3476 123484 3528
rect 123536 3516 123542 3528
rect 124858 3516 124864 3528
rect 123536 3488 124864 3516
rect 123536 3476 123542 3488
rect 124858 3476 124864 3488
rect 124916 3476 124922 3528
rect 126974 3476 126980 3528
rect 127032 3516 127038 3528
rect 128446 3516 128452 3528
rect 127032 3488 128452 3516
rect 127032 3476 127038 3488
rect 128446 3476 128452 3488
rect 128504 3476 128510 3528
rect 136450 3476 136456 3528
rect 136508 3516 136514 3528
rect 141510 3516 141516 3528
rect 136508 3488 141516 3516
rect 136508 3476 136514 3488
rect 141510 3476 141516 3488
rect 141568 3476 141574 3528
rect 147214 3476 147220 3528
rect 147272 3516 147278 3528
rect 148318 3516 148324 3528
rect 147272 3488 148324 3516
rect 147272 3476 147278 3488
rect 148318 3476 148324 3488
rect 148376 3476 148382 3528
rect 148502 3476 148508 3528
rect 148560 3516 148566 3528
rect 148560 3488 171640 3516
rect 148560 3476 148566 3488
rect 124674 3408 124680 3460
rect 124732 3448 124738 3460
rect 131298 3448 131304 3460
rect 124732 3420 131304 3448
rect 124732 3408 124738 3420
rect 131298 3408 131304 3420
rect 131356 3408 131362 3460
rect 141418 3408 141424 3460
rect 141476 3448 141482 3460
rect 141476 3420 161474 3448
rect 141476 3408 141482 3420
rect 131390 3380 131396 3392
rect 123404 3352 131396 3380
rect 131390 3340 131396 3352
rect 131448 3340 131454 3392
rect 143442 3340 143448 3392
rect 143500 3380 143506 3392
rect 150618 3380 150624 3392
rect 143500 3352 150624 3380
rect 143500 3340 143506 3352
rect 150618 3340 150624 3352
rect 150676 3340 150682 3392
rect 157978 3340 157984 3392
rect 158036 3380 158042 3392
rect 158898 3380 158904 3392
rect 158036 3352 158904 3380
rect 158036 3340 158042 3352
rect 158898 3340 158904 3352
rect 158956 3340 158962 3392
rect 131574 3312 131580 3324
rect 122806 3284 131580 3312
rect 131574 3272 131580 3284
rect 131632 3272 131638 3324
rect 161446 3312 161474 3420
rect 171612 3380 171640 3488
rect 171778 3476 171784 3528
rect 171836 3516 171842 3528
rect 173158 3516 173164 3528
rect 171836 3488 173164 3516
rect 171836 3476 171842 3488
rect 173158 3476 173164 3488
rect 173216 3476 173222 3528
rect 178954 3476 178960 3528
rect 179012 3516 179018 3528
rect 470566 3516 470594 3556
rect 179012 3488 470594 3516
rect 179012 3476 179018 3488
rect 472618 3476 472624 3528
rect 472676 3516 472682 3528
rect 473446 3516 473452 3528
rect 472676 3488 473452 3516
rect 472676 3476 472682 3488
rect 473446 3476 473452 3488
rect 473504 3476 473510 3528
rect 478156 3516 478184 3556
rect 478230 3544 478236 3596
rect 478288 3584 478294 3596
rect 500586 3584 500592 3596
rect 478288 3556 500592 3584
rect 478288 3544 478294 3556
rect 500586 3544 500592 3556
rect 500644 3544 500650 3596
rect 525058 3544 525064 3596
rect 525116 3584 525122 3596
rect 527818 3584 527824 3596
rect 525116 3556 527824 3584
rect 525116 3544 525122 3556
rect 527818 3544 527824 3556
rect 527876 3544 527882 3596
rect 560938 3544 560944 3596
rect 560996 3584 561002 3596
rect 564434 3584 564440 3596
rect 560996 3556 564440 3584
rect 560996 3544 561002 3556
rect 564434 3544 564440 3556
rect 564492 3544 564498 3596
rect 574738 3544 574744 3596
rect 574796 3584 574802 3596
rect 576302 3584 576308 3596
rect 574796 3556 576308 3584
rect 574796 3544 574802 3556
rect 576302 3544 576308 3556
rect 576360 3544 576366 3596
rect 479334 3516 479340 3528
rect 478156 3488 479340 3516
rect 479334 3476 479340 3488
rect 479392 3476 479398 3528
rect 506474 3476 506480 3528
rect 506532 3516 506538 3528
rect 507302 3516 507308 3528
rect 506532 3488 507308 3516
rect 506532 3476 506538 3488
rect 507302 3476 507308 3488
rect 507360 3476 507366 3528
rect 514018 3476 514024 3528
rect 514076 3516 514082 3528
rect 515950 3516 515956 3528
rect 514076 3488 515956 3516
rect 514076 3476 514082 3488
rect 515950 3476 515956 3488
rect 516008 3476 516014 3528
rect 538858 3476 538864 3528
rect 538916 3516 538922 3528
rect 539594 3516 539600 3528
rect 538916 3488 539600 3516
rect 538916 3476 538922 3488
rect 539594 3476 539600 3488
rect 539652 3476 539658 3528
rect 549898 3476 549904 3528
rect 549956 3516 549962 3528
rect 551462 3516 551468 3528
rect 549956 3488 551468 3516
rect 549956 3476 549962 3488
rect 551462 3476 551468 3488
rect 551520 3476 551526 3528
rect 554038 3476 554044 3528
rect 554096 3516 554102 3528
rect 554958 3516 554964 3528
rect 554096 3488 554964 3516
rect 554096 3476 554102 3488
rect 554958 3476 554964 3488
rect 555016 3476 555022 3528
rect 563698 3476 563704 3528
rect 563756 3516 563762 3528
rect 565630 3516 565636 3528
rect 563756 3488 565636 3516
rect 563756 3476 563762 3488
rect 565630 3476 565636 3488
rect 565688 3476 565694 3528
rect 567930 3476 567936 3528
rect 567988 3516 567994 3528
rect 569126 3516 569132 3528
rect 567988 3488 569132 3516
rect 567988 3476 567994 3488
rect 569126 3476 569132 3488
rect 569184 3476 569190 3528
rect 180518 3408 180524 3460
rect 180576 3448 180582 3460
rect 487614 3448 487620 3460
rect 180576 3420 487620 3448
rect 180576 3408 180582 3420
rect 487614 3408 487620 3420
rect 487672 3408 487678 3460
rect 511350 3408 511356 3460
rect 511408 3448 511414 3460
rect 514754 3448 514760 3460
rect 511408 3420 514760 3448
rect 511408 3408 511414 3420
rect 514754 3408 514760 3420
rect 514812 3408 514818 3460
rect 527910 3408 527916 3460
rect 527968 3448 527974 3460
rect 533706 3448 533712 3460
rect 527968 3420 533712 3448
rect 527968 3408 527974 3420
rect 533706 3408 533712 3420
rect 533764 3408 533770 3460
rect 567838 3408 567844 3460
rect 567896 3448 567902 3460
rect 572714 3448 572720 3460
rect 567896 3420 572720 3448
rect 567896 3408 567902 3420
rect 572714 3408 572720 3420
rect 572772 3408 572778 3460
rect 176654 3380 176660 3392
rect 171612 3352 176660 3380
rect 176654 3340 176660 3352
rect 176712 3340 176718 3392
rect 184290 3340 184296 3392
rect 184348 3380 184354 3392
rect 189718 3380 189724 3392
rect 184348 3352 189724 3380
rect 184348 3340 184354 3352
rect 189718 3340 189724 3352
rect 189776 3340 189782 3392
rect 189810 3340 189816 3392
rect 189868 3380 189874 3392
rect 190822 3380 190828 3392
rect 189868 3352 190828 3380
rect 189868 3340 189874 3352
rect 190822 3340 190828 3352
rect 190880 3340 190886 3392
rect 193122 3340 193128 3392
rect 193180 3380 193186 3392
rect 195698 3380 195704 3392
rect 193180 3352 195704 3380
rect 193180 3340 193186 3352
rect 195698 3340 195704 3352
rect 195756 3340 195762 3392
rect 204162 3340 204168 3392
rect 204220 3380 204226 3392
rect 207382 3380 207388 3392
rect 204220 3352 207388 3380
rect 204220 3340 204226 3352
rect 207382 3340 207388 3352
rect 207440 3340 207446 3392
rect 239398 3340 239404 3392
rect 239456 3380 239462 3392
rect 240502 3380 240508 3392
rect 239456 3352 240508 3380
rect 239456 3340 239462 3352
rect 240502 3340 240508 3352
rect 240560 3340 240566 3392
rect 261478 3340 261484 3392
rect 261536 3380 261542 3392
rect 262950 3380 262956 3392
rect 261536 3352 262956 3380
rect 261536 3340 261542 3352
rect 262950 3340 262956 3352
rect 263008 3340 263014 3392
rect 275278 3340 275284 3392
rect 275336 3380 275342 3392
rect 277118 3380 277124 3392
rect 275336 3352 277124 3380
rect 275336 3340 275342 3352
rect 277118 3340 277124 3352
rect 277176 3340 277182 3392
rect 279418 3340 279424 3392
rect 279476 3380 279482 3392
rect 280706 3380 280712 3392
rect 279476 3352 280712 3380
rect 279476 3340 279482 3352
rect 280706 3340 280712 3352
rect 280764 3340 280770 3392
rect 307018 3340 307024 3392
rect 307076 3380 307082 3392
rect 309042 3380 309048 3392
rect 307076 3352 309048 3380
rect 307076 3340 307082 3352
rect 309042 3340 309048 3352
rect 309100 3340 309106 3392
rect 324406 3340 324412 3392
rect 324464 3380 324470 3392
rect 325602 3380 325608 3392
rect 324464 3352 325608 3380
rect 324464 3340 324470 3352
rect 325602 3340 325608 3352
rect 325660 3340 325666 3392
rect 329098 3340 329104 3392
rect 329156 3380 329162 3392
rect 330386 3380 330392 3392
rect 329156 3352 330392 3380
rect 329156 3340 329162 3352
rect 330386 3340 330392 3352
rect 330444 3340 330450 3392
rect 340966 3340 340972 3392
rect 341024 3380 341030 3392
rect 342162 3380 342168 3392
rect 341024 3352 342168 3380
rect 341024 3340 341030 3352
rect 342162 3340 342168 3352
rect 342220 3340 342226 3392
rect 342898 3340 342904 3392
rect 342956 3380 342962 3392
rect 344554 3380 344560 3392
rect 342956 3352 344560 3380
rect 342956 3340 342962 3352
rect 344554 3340 344560 3352
rect 344612 3340 344618 3392
rect 356698 3340 356704 3392
rect 356756 3380 356762 3392
rect 358722 3380 358728 3392
rect 356756 3352 358728 3380
rect 356756 3340 356762 3352
rect 358722 3340 358728 3352
rect 358780 3340 358786 3392
rect 364978 3340 364984 3392
rect 365036 3380 365042 3392
rect 367002 3380 367008 3392
rect 365036 3352 367008 3380
rect 365036 3340 365042 3352
rect 367002 3340 367008 3352
rect 367060 3340 367066 3392
rect 374086 3340 374092 3392
rect 374144 3380 374150 3392
rect 375282 3380 375288 3392
rect 374144 3352 375288 3380
rect 374144 3340 374150 3352
rect 375282 3340 375288 3352
rect 375340 3340 375346 3392
rect 382366 3340 382372 3392
rect 382424 3380 382430 3392
rect 383562 3380 383568 3392
rect 382424 3352 383568 3380
rect 382424 3340 382430 3352
rect 383562 3340 383568 3352
rect 383620 3340 383626 3392
rect 390554 3340 390560 3392
rect 390612 3380 390618 3392
rect 391842 3380 391848 3392
rect 390612 3352 391848 3380
rect 390612 3340 390618 3352
rect 391842 3340 391848 3352
rect 391900 3340 391906 3392
rect 398926 3340 398932 3392
rect 398984 3380 398990 3392
rect 400122 3380 400128 3392
rect 398984 3352 400128 3380
rect 398984 3340 398990 3352
rect 400122 3340 400128 3352
rect 400180 3340 400186 3392
rect 400858 3340 400864 3392
rect 400916 3380 400922 3392
rect 402514 3380 402520 3392
rect 400916 3352 402520 3380
rect 400916 3340 400922 3352
rect 402514 3340 402520 3352
rect 402572 3340 402578 3392
rect 414658 3340 414664 3392
rect 414716 3380 414722 3392
rect 416682 3380 416688 3392
rect 414716 3352 416688 3380
rect 414716 3340 414722 3352
rect 416682 3340 416688 3352
rect 416740 3340 416746 3392
rect 418798 3340 418804 3392
rect 418856 3380 418862 3392
rect 420178 3380 420184 3392
rect 418856 3352 420184 3380
rect 418856 3340 418862 3352
rect 420178 3340 420184 3352
rect 420236 3340 420242 3392
rect 423674 3340 423680 3392
rect 423732 3380 423738 3392
rect 424962 3380 424968 3392
rect 423732 3352 424968 3380
rect 423732 3340 423738 3352
rect 424962 3340 424968 3352
rect 425020 3340 425026 3392
rect 432598 3340 432604 3392
rect 432656 3380 432662 3392
rect 434438 3380 434444 3392
rect 432656 3352 434444 3380
rect 432656 3340 432662 3352
rect 434438 3340 434444 3352
rect 434496 3340 434502 3392
rect 440234 3340 440240 3392
rect 440292 3380 440298 3392
rect 441522 3380 441528 3392
rect 440292 3352 441528 3380
rect 440292 3340 440298 3352
rect 441522 3340 441528 3352
rect 441580 3340 441586 3392
rect 446398 3340 446404 3392
rect 446456 3380 446462 3392
rect 447410 3380 447416 3392
rect 446456 3352 447416 3380
rect 446456 3340 446462 3352
rect 447410 3340 447416 3352
rect 447468 3340 447474 3392
rect 448606 3340 448612 3392
rect 448664 3380 448670 3392
rect 449802 3380 449808 3392
rect 448664 3352 449808 3380
rect 448664 3340 448670 3352
rect 449802 3340 449808 3352
rect 449860 3340 449866 3392
rect 456794 3340 456800 3392
rect 456852 3380 456858 3392
rect 458082 3380 458088 3392
rect 456852 3352 458088 3380
rect 456852 3340 456858 3352
rect 458082 3340 458088 3352
rect 458140 3340 458146 3392
rect 482278 3340 482284 3392
rect 482336 3380 482342 3392
rect 484026 3380 484032 3392
rect 482336 3352 484032 3380
rect 482336 3340 482342 3352
rect 484026 3340 484032 3352
rect 484084 3340 484090 3392
rect 534718 3340 534724 3392
rect 534776 3380 534782 3392
rect 550266 3380 550272 3392
rect 534776 3352 550272 3380
rect 534776 3340 534782 3352
rect 550266 3340 550272 3352
rect 550324 3340 550330 3392
rect 175458 3312 175464 3324
rect 161446 3284 175464 3312
rect 175458 3272 175464 3284
rect 175516 3272 175522 3324
rect 189902 3272 189908 3324
rect 189960 3312 189966 3324
rect 193214 3312 193220 3324
rect 189960 3284 193220 3312
rect 189960 3272 189966 3284
rect 193214 3272 193220 3284
rect 193272 3272 193278 3324
rect 210418 3272 210424 3324
rect 210476 3312 210482 3324
rect 218054 3312 218060 3324
rect 210476 3284 218060 3312
rect 210476 3272 210482 3284
rect 218054 3272 218060 3284
rect 218112 3272 218118 3324
rect 224218 3272 224224 3324
rect 224276 3312 224282 3324
rect 231026 3312 231032 3324
rect 224276 3284 231032 3312
rect 224276 3272 224282 3284
rect 231026 3272 231032 3284
rect 231084 3272 231090 3324
rect 260098 3272 260104 3324
rect 260156 3312 260162 3324
rect 261754 3312 261760 3324
rect 260156 3284 261760 3312
rect 260156 3272 260162 3284
rect 261754 3272 261760 3284
rect 261812 3272 261818 3324
rect 396718 3272 396724 3324
rect 396776 3312 396782 3324
rect 397730 3312 397736 3324
rect 396776 3284 397736 3312
rect 396776 3272 396782 3284
rect 397730 3272 397736 3284
rect 397788 3272 397794 3324
rect 431954 3272 431960 3324
rect 432012 3312 432018 3324
rect 433242 3312 433248 3324
rect 432012 3284 433248 3312
rect 432012 3272 432018 3284
rect 433242 3272 433248 3284
rect 433300 3272 433306 3324
rect 520918 3272 520924 3324
rect 520976 3312 520982 3324
rect 524230 3312 524236 3324
rect 520976 3284 524236 3312
rect 520976 3272 520982 3284
rect 524230 3272 524236 3284
rect 524288 3272 524294 3324
rect 562318 3272 562324 3324
rect 562376 3312 562382 3324
rect 566826 3312 566832 3324
rect 562376 3284 566832 3312
rect 562376 3272 562382 3284
rect 566826 3272 566832 3284
rect 566884 3272 566890 3324
rect 571978 3272 571984 3324
rect 572036 3312 572042 3324
rect 573910 3312 573916 3324
rect 572036 3284 573916 3312
rect 572036 3272 572042 3284
rect 573910 3272 573916 3284
rect 573968 3272 573974 3324
rect 134150 3204 134156 3256
rect 134208 3244 134214 3256
rect 138658 3244 138664 3256
rect 134208 3216 138664 3244
rect 134208 3204 134214 3216
rect 138658 3204 138664 3216
rect 138716 3204 138722 3256
rect 33594 3136 33600 3188
rect 33652 3176 33658 3188
rect 35158 3176 35164 3188
rect 33652 3148 35164 3176
rect 33652 3136 33658 3148
rect 35158 3136 35164 3148
rect 35216 3136 35222 3188
rect 38378 3136 38384 3188
rect 38436 3176 38442 3188
rect 39298 3176 39304 3188
rect 38436 3148 39304 3176
rect 38436 3136 38442 3148
rect 39298 3136 39304 3148
rect 39356 3136 39362 3188
rect 41874 3136 41880 3188
rect 41932 3176 41938 3188
rect 43438 3176 43444 3188
rect 41932 3148 43444 3176
rect 41932 3136 41938 3148
rect 43438 3136 43444 3148
rect 43496 3136 43502 3188
rect 118786 3136 118792 3188
rect 118844 3176 118850 3188
rect 122098 3176 122104 3188
rect 118844 3148 122104 3176
rect 118844 3136 118850 3148
rect 122098 3136 122104 3148
rect 122156 3136 122162 3188
rect 164878 3136 164884 3188
rect 164936 3176 164942 3188
rect 168374 3176 168380 3188
rect 164936 3148 168380 3176
rect 164936 3136 164942 3148
rect 168374 3136 168380 3148
rect 168432 3136 168438 3188
rect 12342 3068 12348 3120
rect 12400 3108 12406 3120
rect 17218 3108 17224 3120
rect 12400 3080 17224 3108
rect 12400 3068 12406 3080
rect 17218 3068 17224 3080
rect 17276 3068 17282 3120
rect 382918 3068 382924 3120
rect 382976 3108 382982 3120
rect 384758 3108 384764 3120
rect 382976 3080 384764 3108
rect 382976 3068 382982 3080
rect 384758 3068 384764 3080
rect 384816 3068 384822 3120
rect 20622 3000 20628 3052
rect 20680 3040 20686 3052
rect 22738 3040 22744 3052
rect 20680 3012 22744 3040
rect 20680 3000 20686 3012
rect 22738 3000 22744 3012
rect 22796 3000 22802 3052
rect 175918 3000 175924 3052
rect 175976 3040 175982 3052
rect 177850 3040 177856 3052
rect 175976 3012 177856 3040
rect 175976 3000 175982 3012
rect 177850 3000 177856 3012
rect 177908 3000 177914 3052
rect 464338 3000 464344 3052
rect 464396 3040 464402 3052
rect 466270 3040 466276 3052
rect 464396 3012 466276 3040
rect 464396 3000 464402 3012
rect 466270 3000 466276 3012
rect 466328 3000 466334 3052
rect 132954 2932 132960 2984
rect 133012 2972 133018 2984
rect 139486 2972 139492 2984
rect 133012 2944 139492 2972
rect 133012 2932 133018 2944
rect 139486 2932 139492 2944
rect 139544 2932 139550 2984
rect 23014 2864 23020 2916
rect 23072 2904 23078 2916
rect 25498 2904 25504 2916
rect 23072 2876 25504 2904
rect 23072 2864 23078 2876
rect 25498 2864 25504 2876
rect 25556 2864 25562 2916
rect 128170 2864 128176 2916
rect 128228 2904 128234 2916
rect 128998 2904 129004 2916
rect 128228 2876 129004 2904
rect 128228 2864 128234 2876
rect 128998 2864 129004 2876
rect 129056 2864 129062 2916
rect 181438 2864 181444 2916
rect 181496 2904 181502 2916
rect 182542 2904 182548 2916
rect 181496 2876 182548 2904
rect 181496 2864 181502 2876
rect 182542 2864 182548 2876
rect 182600 2864 182606 2916
rect 332594 1096 332600 1148
rect 332652 1136 332658 1148
rect 333882 1136 333888 1148
rect 332652 1108 333888 1136
rect 332652 1096 332658 1108
rect 333882 1096 333888 1108
rect 333940 1096 333946 1148
<< via1 >>
rect 71780 702992 71832 703044
rect 72976 702992 73028 703044
rect 137836 700816 137888 700868
rect 157340 700816 157392 700868
rect 155960 700748 156012 700800
rect 202788 700748 202840 700800
rect 89168 700680 89220 700732
rect 160744 700680 160796 700732
rect 154580 700612 154632 700664
rect 267648 700612 267700 700664
rect 24308 700544 24360 700596
rect 162216 700544 162268 700596
rect 8116 700476 8168 700528
rect 162124 700476 162176 700528
rect 153292 700408 153344 700460
rect 332508 700408 332560 700460
rect 153108 700340 153160 700392
rect 413652 700340 413704 700392
rect 148324 700272 148376 700324
rect 543464 700272 543516 700324
rect 543004 700204 543056 700256
rect 559656 700272 559708 700324
rect 105452 699660 105504 699712
rect 106924 699660 106976 699712
rect 396724 699660 396776 699712
rect 397460 699660 397512 699712
rect 428464 699660 428516 699712
rect 429844 699660 429896 699712
rect 146300 696940 146352 696992
rect 580172 696940 580224 696992
rect 3424 683204 3476 683256
rect 162308 683204 162360 683256
rect 146944 683136 146996 683188
rect 580172 683136 580224 683188
rect 3516 670692 3568 670744
rect 163504 670692 163556 670744
rect 185584 670692 185636 670744
rect 580172 670692 580224 670744
rect 149060 660288 149112 660340
rect 462320 660288 462372 660340
rect 3424 656888 3476 656940
rect 163596 656888 163648 656940
rect 184204 643084 184256 643136
rect 580172 643084 580224 643136
rect 3424 632068 3476 632120
rect 164240 632068 164292 632120
rect 203524 630640 203576 630692
rect 580172 630640 580224 630692
rect 3148 618264 3200 618316
rect 164884 618264 164936 618316
rect 143632 616836 143684 616888
rect 580172 616836 580224 616888
rect 3240 605820 3292 605872
rect 164976 605820 165028 605872
rect 142160 590656 142212 590708
rect 579804 590656 579856 590708
rect 3332 579640 3384 579692
rect 165620 579640 165672 579692
rect 144184 576852 144236 576904
rect 580172 576852 580224 576904
rect 3424 565836 3476 565888
rect 167644 565836 167696 565888
rect 142804 563048 142856 563100
rect 579804 563048 579856 563100
rect 3424 553392 3476 553444
rect 166264 553392 166316 553444
rect 178684 536800 178736 536852
rect 580172 536800 580224 536852
rect 3424 527144 3476 527196
rect 167000 527144 167052 527196
rect 142896 524424 142948 524476
rect 580172 524424 580224 524476
rect 3424 514768 3476 514820
rect 8944 514768 8996 514820
rect 181444 510620 181496 510672
rect 580172 510620 580224 510672
rect 3056 500964 3108 501016
rect 167736 500964 167788 501016
rect 139400 484372 139452 484424
rect 580172 484372 580224 484424
rect 140044 470568 140096 470620
rect 579988 470568 580040 470620
rect 3516 462340 3568 462392
rect 170404 462340 170456 462392
rect 180064 456764 180116 456816
rect 580172 456764 580224 456816
rect 3148 448536 3200 448588
rect 170496 448536 170548 448588
rect 157432 447788 157484 447840
rect 169760 447788 169812 447840
rect 138664 430584 138716 430636
rect 580172 430584 580224 430636
rect 3516 422288 3568 422340
rect 169760 422288 169812 422340
rect 138756 418140 138808 418192
rect 580172 418140 580224 418192
rect 2872 409844 2924 409896
rect 171784 409844 171836 409896
rect 199384 404336 199436 404388
rect 580172 404336 580224 404388
rect 3516 397468 3568 397520
rect 171140 397468 171192 397520
rect 182824 378156 182876 378208
rect 580172 378156 580224 378208
rect 2780 371288 2832 371340
rect 4804 371288 4856 371340
rect 3148 357416 3200 357468
rect 10324 357416 10376 357468
rect 135260 351908 135312 351960
rect 580172 351908 580224 351960
rect 3516 345176 3568 345228
rect 7564 345176 7616 345228
rect 134524 324300 134576 324352
rect 580172 324300 580224 324352
rect 3332 318792 3384 318844
rect 173900 318792 173952 318844
rect 135904 311856 135956 311908
rect 579988 311856 580040 311908
rect 3516 304988 3568 305040
rect 175924 304988 175976 305040
rect 134616 298120 134668 298172
rect 580172 298120 580224 298172
rect 3516 292544 3568 292596
rect 174544 292544 174596 292596
rect 10324 289076 10376 289128
rect 173164 289076 173216 289128
rect 145564 287648 145616 287700
rect 203524 287648 203576 287700
rect 137284 286288 137336 286340
rect 182824 286288 182876 286340
rect 186320 284928 186372 284980
rect 187148 284928 187200 284980
rect 396724 284928 396776 284980
rect 150440 284316 150492 284368
rect 186320 284316 186372 284368
rect 147956 283568 148008 283620
rect 527180 283568 527232 283620
rect 145104 282140 145156 282192
rect 184204 282140 184256 282192
rect 140780 280780 140832 280832
rect 178684 280780 178736 280832
rect 40040 279420 40092 279472
rect 160100 279420 160152 279472
rect 204168 276632 204220 276684
rect 299480 276632 299532 276684
rect 153384 276020 153436 276072
rect 203064 276020 203116 276072
rect 204168 276020 204220 276072
rect 204812 275272 204864 275324
rect 364340 275272 364392 275324
rect 151820 274660 151872 274712
rect 204536 274660 204588 274712
rect 204812 274660 204864 274712
rect 8944 273980 8996 274032
rect 169024 273980 169076 274032
rect 151084 273912 151136 273964
rect 428464 273912 428516 273964
rect 133144 271872 133196 271924
rect 580172 271872 580224 271924
rect 7564 271192 7616 271244
rect 173256 271192 173308 271244
rect 149152 271124 149204 271176
rect 494060 271124 494112 271176
rect 71780 269764 71832 269816
rect 121460 269764 121512 269816
rect 147772 269764 147824 269816
rect 543004 269764 543056 269816
rect 121460 269084 121512 269136
rect 122380 269084 122432 269136
rect 158720 269084 158772 269136
rect 146208 268404 146260 268456
rect 185584 268404 185636 268456
rect 4804 268336 4856 268388
rect 172704 268336 172756 268388
rect 137836 266976 137888 267028
rect 199384 266976 199436 267028
rect 3056 266364 3108 266416
rect 175924 266364 175976 266416
rect 174544 265752 174596 265804
rect 141700 265684 141752 265736
rect 181444 265684 181496 265736
rect 3424 265616 3476 265668
rect 169208 265616 169260 265668
rect 192024 265616 192076 265668
rect 173256 265548 173308 265600
rect 192116 265548 192168 265600
rect 175832 265480 175884 265532
rect 199200 265480 199252 265532
rect 170404 265412 170456 265464
rect 170680 265412 170732 265464
rect 195060 265412 195112 265464
rect 171784 265344 171836 265396
rect 196624 265344 196676 265396
rect 167828 265276 167880 265328
rect 193588 265276 193640 265328
rect 162308 265208 162360 265260
rect 188252 265208 188304 265260
rect 169116 265140 169168 265192
rect 196256 265140 196308 265192
rect 167460 265072 167512 265124
rect 194968 265072 195020 265124
rect 164884 265004 164936 265056
rect 165344 265004 165396 265056
rect 196440 265004 196492 265056
rect 152188 264936 152240 264988
rect 153108 264936 153160 264988
rect 187516 264936 187568 264988
rect 120816 264256 120868 264308
rect 139492 264256 139544 264308
rect 106924 264188 106976 264240
rect 121460 264188 121512 264240
rect 180064 264188 180116 264240
rect 118240 264120 118292 264172
rect 134248 264120 134300 264172
rect 134616 264120 134668 264172
rect 115572 264052 115624 264104
rect 133144 264052 133196 264104
rect 120908 263984 120960 264036
rect 141148 263984 141200 264036
rect 141700 263984 141752 264036
rect 115388 263916 115440 263968
rect 137192 263916 137244 263968
rect 119804 263848 119856 263900
rect 142620 263848 142672 263900
rect 122564 263780 122616 263832
rect 148508 263780 148560 263832
rect 119712 263712 119764 263764
rect 146208 263712 146260 263764
rect 120724 263644 120776 263696
rect 151084 263644 151136 263696
rect 172704 263644 172756 263696
rect 189356 263644 189408 263696
rect 121460 263576 121512 263628
rect 122012 263576 122064 263628
rect 159088 263576 159140 263628
rect 173164 263576 173216 263628
rect 173716 263576 173768 263628
rect 197912 263576 197964 263628
rect 137468 263508 137520 263560
rect 580264 263508 580316 263560
rect 150440 263440 150492 263492
rect 151360 263440 151412 263492
rect 193128 263440 193180 263492
rect 218060 263440 218112 263492
rect 163412 263236 163464 263288
rect 163596 263236 163648 263288
rect 170220 263032 170272 263084
rect 170496 263032 170548 263084
rect 192300 263032 192352 263084
rect 116768 262964 116820 263016
rect 131120 262964 131172 263016
rect 132040 262964 132092 263016
rect 580356 262964 580408 263016
rect 3424 262896 3476 262948
rect 178500 262896 178552 262948
rect 179236 262896 179288 262948
rect 189540 262896 189592 262948
rect 113824 262828 113876 262880
rect 131764 262828 131816 262880
rect 580448 262828 580500 262880
rect 113916 262760 113968 262812
rect 134524 262760 134576 262812
rect 134800 262760 134852 262812
rect 163412 262760 163464 262812
rect 192392 262760 192444 262812
rect 116676 262692 116728 262744
rect 127716 262692 127768 262744
rect 162032 262692 162084 262744
rect 193772 262692 193824 262744
rect 115296 262624 115348 262676
rect 129832 262624 129884 262676
rect 153200 262624 153252 262676
rect 158720 262624 158772 262676
rect 162216 262624 162268 262676
rect 195152 262624 195204 262676
rect 112904 262556 112956 262608
rect 128728 262556 128780 262608
rect 157156 262556 157208 262608
rect 192484 262556 192536 262608
rect 193128 262556 193180 262608
rect 121920 262488 121972 262540
rect 144184 262488 144236 262540
rect 160744 262488 160796 262540
rect 200580 262488 200632 262540
rect 3516 262420 3568 262472
rect 176752 262420 176804 262472
rect 180156 262420 180208 262472
rect 193496 262420 193548 262472
rect 118148 262352 118200 262404
rect 129280 262352 129332 262404
rect 182916 262352 182968 262404
rect 184572 262284 184624 262336
rect 189172 262284 189224 262336
rect 190460 262284 190512 262336
rect 122472 262216 122524 262268
rect 125968 262216 126020 262268
rect 181260 262216 181312 262268
rect 187792 262216 187844 262268
rect 129832 261400 129884 261452
rect 188344 261400 188396 261452
rect 176752 261332 176804 261384
rect 198004 261332 198056 261384
rect 131120 261264 131172 261316
rect 471244 261264 471296 261316
rect 184020 261196 184072 261248
rect 199016 261196 199068 261248
rect 118056 261128 118108 261180
rect 132868 261128 132920 261180
rect 180524 261128 180576 261180
rect 198096 261128 198148 261180
rect 111248 261060 111300 261112
rect 132040 261060 132092 261112
rect 178500 261060 178552 261112
rect 199108 261060 199160 261112
rect 111432 260992 111484 261044
rect 130384 260992 130436 261044
rect 181996 260992 182048 261044
rect 197820 260992 197872 261044
rect 4804 260924 4856 260976
rect 176200 260924 176252 260976
rect 190920 260924 190972 260976
rect 112628 260856 112680 260908
rect 133972 260856 134024 260908
rect 177580 260856 177632 260908
rect 191012 260856 191064 260908
rect 119344 260788 119396 260840
rect 124312 260788 124364 260840
rect 173900 260380 173952 260432
rect 185584 260380 185636 260432
rect 190736 260380 190788 260432
rect 187884 260312 187936 260364
rect 116584 260176 116636 260228
rect 135260 260176 135312 260228
rect 136226 260176 136278 260228
rect 157340 260176 157392 260228
rect 158306 260176 158358 260228
rect 167000 260176 167052 260228
rect 167690 260176 167742 260228
rect 169760 260176 169812 260228
rect 171002 260176 171054 260228
rect 175924 260244 175976 260296
rect 176108 260176 176160 260228
rect 178408 260244 178460 260296
rect 189632 260244 189684 260296
rect 187332 260176 187384 260228
rect 132914 260108 132966 260160
rect 485044 260108 485096 260160
rect 114008 260040 114060 260092
rect 126842 260040 126894 260092
rect 171002 260040 171054 260092
rect 185584 260040 185636 260092
rect 185676 260040 185728 260092
rect 190828 260040 190880 260092
rect 113640 259972 113692 260024
rect 128360 259972 128412 260024
rect 117872 259904 117924 259956
rect 142160 259904 142212 259956
rect 143080 259904 143132 259956
rect 119436 259836 119488 259888
rect 146300 259836 146352 259888
rect 169484 259836 169536 259888
rect 189448 259972 189500 260024
rect 171692 259904 171744 259956
rect 176108 259836 176160 259888
rect 185676 259836 185728 259888
rect 119528 259768 119580 259820
rect 149152 259768 149204 259820
rect 158076 259768 158128 259820
rect 187976 259768 188028 259820
rect 193680 259904 193732 259956
rect 119620 259700 119672 259752
rect 153200 259700 153252 259752
rect 158628 259700 158680 259752
rect 188160 259700 188212 259752
rect 134340 259632 134392 259684
rect 187700 259632 187752 259684
rect 120540 259564 120592 259616
rect 178040 259564 178092 259616
rect 181812 259564 181864 259616
rect 203432 259564 203484 259616
rect 7564 259496 7616 259548
rect 177304 259496 177356 259548
rect 183468 259496 183520 259548
rect 206100 259496 206152 259548
rect 117964 259428 118016 259480
rect 139400 259428 139452 259480
rect 139768 259428 139820 259480
rect 184940 259428 184992 259480
rect 196532 259428 196584 259480
rect 187700 259360 187752 259412
rect 580172 259360 580224 259412
rect 187792 258476 187844 258528
rect 188068 258476 188120 258528
rect 485044 245556 485096 245608
rect 580172 245556 580224 245608
rect 2780 241204 2832 241256
rect 4804 241204 4856 241256
rect 3516 215092 3568 215144
rect 7564 215092 7616 215144
rect 471244 206932 471296 206984
rect 579804 206932 579856 206984
rect 104440 200540 104492 200592
rect 130844 200676 130896 200728
rect 119068 200472 119120 200524
rect 132040 200676 132092 200728
rect 132132 200676 132184 200728
rect 132224 200676 132276 200728
rect 131120 200608 131172 200660
rect 132040 200540 132092 200592
rect 132224 200540 132276 200592
rect 113088 200404 113140 200456
rect 112996 200336 113048 200388
rect 119896 200268 119948 200320
rect 132132 200268 132184 200320
rect 118608 200200 118660 200252
rect 130844 200064 130896 200116
rect 102876 199656 102928 199708
rect 106004 199588 106056 199640
rect 132914 199860 132966 199912
rect 133006 199860 133058 199912
rect 126060 199724 126112 199776
rect 130752 199656 130804 199708
rect 130660 199588 130712 199640
rect 133282 199860 133334 199912
rect 133466 199860 133518 199912
rect 133650 199860 133702 199912
rect 133742 199860 133794 199912
rect 133926 199860 133978 199912
rect 134202 199860 134254 199912
rect 134478 199860 134530 199912
rect 134754 199860 134806 199912
rect 135030 199860 135082 199912
rect 135122 199860 135174 199912
rect 135214 199860 135266 199912
rect 135306 199860 135358 199912
rect 135398 199860 135450 199912
rect 133650 199724 133702 199776
rect 134018 199792 134070 199844
rect 133880 199724 133932 199776
rect 133788 199656 133840 199708
rect 133420 199588 133472 199640
rect 133604 199588 133656 199640
rect 134156 199656 134208 199708
rect 134432 199656 134484 199708
rect 134800 199656 134852 199708
rect 135076 199724 135128 199776
rect 135766 199860 135818 199912
rect 136042 199860 136094 199912
rect 136134 199860 136186 199912
rect 136318 199792 136370 199844
rect 135490 199724 135542 199776
rect 136088 199724 136140 199776
rect 134984 199588 135036 199640
rect 135168 199588 135220 199640
rect 135306 199588 135358 199640
rect 135444 199588 135496 199640
rect 136180 199588 136232 199640
rect 136594 199860 136646 199912
rect 136686 199860 136738 199912
rect 136778 199860 136830 199912
rect 137238 199860 137290 199912
rect 137330 199860 137382 199912
rect 136732 199724 136784 199776
rect 136640 199656 136692 199708
rect 136548 199588 136600 199640
rect 137192 199588 137244 199640
rect 114928 199520 114980 199572
rect 132960 199520 133012 199572
rect 133696 199520 133748 199572
rect 136824 199520 136876 199572
rect 137284 199520 137336 199572
rect 137790 199860 137842 199912
rect 137882 199860 137934 199912
rect 137974 199860 138026 199912
rect 138066 199860 138118 199912
rect 138250 199860 138302 199912
rect 138526 199860 138578 199912
rect 137514 199792 137566 199844
rect 137606 199792 137658 199844
rect 137928 199724 137980 199776
rect 138020 199724 138072 199776
rect 138434 199792 138486 199844
rect 137560 199588 137612 199640
rect 137652 199588 137704 199640
rect 137744 199588 137796 199640
rect 138112 199588 138164 199640
rect 138480 199588 138532 199640
rect 138710 199860 138762 199912
rect 138802 199860 138854 199912
rect 138894 199860 138946 199912
rect 138756 199724 138808 199776
rect 138848 199656 138900 199708
rect 139170 199860 139222 199912
rect 139354 199860 139406 199912
rect 139032 199588 139084 199640
rect 139308 199588 139360 199640
rect 137836 199520 137888 199572
rect 138388 199520 138440 199572
rect 138664 199520 138716 199572
rect 138756 199520 138808 199572
rect 139538 199860 139590 199912
rect 139722 199860 139774 199912
rect 139814 199860 139866 199912
rect 139906 199860 139958 199912
rect 139998 199860 140050 199912
rect 140182 199860 140234 199912
rect 140366 199860 140418 199912
rect 140458 199860 140510 199912
rect 139676 199724 139728 199776
rect 139860 199724 139912 199776
rect 139952 199724 140004 199776
rect 139584 199656 139636 199708
rect 140044 199588 140096 199640
rect 140228 199520 140280 199572
rect 140412 199724 140464 199776
rect 140734 199860 140786 199912
rect 140826 199860 140878 199912
rect 141010 199860 141062 199912
rect 141286 199860 141338 199912
rect 140734 199724 140786 199776
rect 141470 199860 141522 199912
rect 141746 199860 141798 199912
rect 140872 199656 140924 199708
rect 141424 199656 141476 199708
rect 141608 199588 141660 199640
rect 142022 199860 142074 199912
rect 141930 199792 141982 199844
rect 142206 199860 142258 199912
rect 142160 199656 142212 199708
rect 141884 199588 141936 199640
rect 141976 199588 142028 199640
rect 141148 199520 141200 199572
rect 141516 199520 141568 199572
rect 141792 199520 141844 199572
rect 142574 199860 142626 199912
rect 142666 199860 142718 199912
rect 142758 199860 142810 199912
rect 142482 199724 142534 199776
rect 142528 199588 142580 199640
rect 142942 199860 142994 199912
rect 143126 199860 143178 199912
rect 143218 199792 143270 199844
rect 143310 199792 143362 199844
rect 143402 199792 143454 199844
rect 143080 199656 143132 199708
rect 143172 199656 143224 199708
rect 143678 199860 143730 199912
rect 143770 199860 143822 199912
rect 144046 199860 144098 199912
rect 144138 199860 144190 199912
rect 144414 199860 144466 199912
rect 144506 199860 144558 199912
rect 144598 199860 144650 199912
rect 145058 199860 145110 199912
rect 145150 199860 145202 199912
rect 143816 199724 143868 199776
rect 142712 199588 142764 199640
rect 143264 199588 143316 199640
rect 143448 199588 143500 199640
rect 143540 199588 143592 199640
rect 143724 199588 143776 199640
rect 142620 199520 142672 199572
rect 143356 199520 143408 199572
rect 118332 199452 118384 199504
rect 142436 199452 142488 199504
rect 122472 199384 122524 199436
rect 126612 199384 126664 199436
rect 127900 199384 127952 199436
rect 135168 199384 135220 199436
rect 143356 199384 143408 199436
rect 143908 199520 143960 199572
rect 144460 199656 144512 199708
rect 144782 199792 144834 199844
rect 144552 199588 144604 199640
rect 144184 199520 144236 199572
rect 144644 199520 144696 199572
rect 145104 199656 145156 199708
rect 145012 199588 145064 199640
rect 145334 199860 145386 199912
rect 145610 199860 145662 199912
rect 145794 199860 145846 199912
rect 145886 199860 145938 199912
rect 146070 199860 146122 199912
rect 146162 199860 146214 199912
rect 146530 199860 146582 199912
rect 146622 199860 146674 199912
rect 145472 199588 145524 199640
rect 145840 199656 145892 199708
rect 146208 199724 146260 199776
rect 146116 199656 146168 199708
rect 146806 199860 146858 199912
rect 146898 199860 146950 199912
rect 146990 199860 147042 199912
rect 146852 199724 146904 199776
rect 146944 199656 146996 199708
rect 146760 199588 146812 199640
rect 145288 199520 145340 199572
rect 145748 199520 145800 199572
rect 146024 199520 146076 199572
rect 147818 199860 147870 199912
rect 148370 199860 148422 199912
rect 148462 199860 148514 199912
rect 148646 199860 148698 199912
rect 148738 199860 148790 199912
rect 147680 199588 147732 199640
rect 148416 199724 148468 199776
rect 148508 199724 148560 199776
rect 148600 199724 148652 199776
rect 147404 199452 147456 199504
rect 147588 199452 147640 199504
rect 147312 199384 147364 199436
rect 121368 199316 121420 199368
rect 132132 199248 132184 199300
rect 132776 199248 132828 199300
rect 132960 199248 133012 199300
rect 133696 199248 133748 199300
rect 135812 199316 135864 199368
rect 142160 199316 142212 199368
rect 142528 199316 142580 199368
rect 139492 199248 139544 199300
rect 145104 199248 145156 199300
rect 146392 199316 146444 199368
rect 147404 199316 147456 199368
rect 149014 199860 149066 199912
rect 149290 199860 149342 199912
rect 149474 199860 149526 199912
rect 149566 199860 149618 199912
rect 149658 199860 149710 199912
rect 149336 199588 149388 199640
rect 149520 199588 149572 199640
rect 148968 199520 149020 199572
rect 149152 199520 149204 199572
rect 149612 199452 149664 199504
rect 118424 199180 118476 199232
rect 145656 199180 145708 199232
rect 117136 199112 117188 199164
rect 145380 199112 145432 199164
rect 114376 199044 114428 199096
rect 142344 199044 142396 199096
rect 143356 199044 143408 199096
rect 150118 199860 150170 199912
rect 150946 199860 150998 199912
rect 151222 199860 151274 199912
rect 151774 199860 151826 199912
rect 151958 199860 152010 199912
rect 152234 199860 152286 199912
rect 152326 199860 152378 199912
rect 152418 199860 152470 199912
rect 152694 199860 152746 199912
rect 152786 199860 152838 199912
rect 152878 199860 152930 199912
rect 152004 199724 152056 199776
rect 151912 199656 151964 199708
rect 152280 199724 152332 199776
rect 152372 199724 152424 199776
rect 152740 199724 152792 199776
rect 152832 199724 152884 199776
rect 152188 199588 152240 199640
rect 153062 199860 153114 199912
rect 152740 199452 152792 199504
rect 177764 200608 177816 200660
rect 184204 200676 184256 200728
rect 180064 200608 180116 200660
rect 153338 199860 153390 199912
rect 153430 199860 153482 199912
rect 153384 199724 153436 199776
rect 153614 199860 153666 199912
rect 153706 199860 153758 199912
rect 153798 199860 153850 199912
rect 153890 199860 153942 199912
rect 153982 199860 154034 199912
rect 154258 199860 154310 199912
rect 153660 199724 153712 199776
rect 153936 199724 153988 199776
rect 153752 199656 153804 199708
rect 154442 199860 154494 199912
rect 155178 199860 155230 199912
rect 153568 199588 153620 199640
rect 154304 199588 154356 199640
rect 153844 199520 153896 199572
rect 154120 199520 154172 199572
rect 155362 199860 155414 199912
rect 155454 199860 155506 199912
rect 155730 199860 155782 199912
rect 155822 199860 155874 199912
rect 155914 199860 155966 199912
rect 156374 199860 156426 199912
rect 156466 199860 156518 199912
rect 156558 199860 156610 199912
rect 155408 199724 155460 199776
rect 155224 199656 155276 199708
rect 155776 199724 155828 199776
rect 155868 199724 155920 199776
rect 155684 199588 155736 199640
rect 153200 199452 153252 199504
rect 156236 199452 156288 199504
rect 156604 199588 156656 199640
rect 156926 199860 156978 199912
rect 157018 199860 157070 199912
rect 157110 199860 157162 199912
rect 157478 199860 157530 199912
rect 157064 199656 157116 199708
rect 156972 199588 157024 199640
rect 157524 199724 157576 199776
rect 157846 199860 157898 199912
rect 158030 199860 158082 199912
rect 158306 199860 158358 199912
rect 158398 199860 158450 199912
rect 158582 199860 158634 199912
rect 158674 199860 158726 199912
rect 158766 199860 158818 199912
rect 158628 199724 158680 199776
rect 158720 199724 158772 199776
rect 158352 199656 158404 199708
rect 158536 199656 158588 199708
rect 157984 199588 158036 199640
rect 178040 200540 178092 200592
rect 178132 200540 178184 200592
rect 191932 200540 191984 200592
rect 177948 200472 178000 200524
rect 193220 200472 193272 200524
rect 180340 200404 180392 200456
rect 158950 199860 159002 199912
rect 159042 199860 159094 199912
rect 159134 199860 159186 199912
rect 158996 199656 159048 199708
rect 159088 199656 159140 199708
rect 159594 199860 159646 199912
rect 159778 199860 159830 199912
rect 159870 199860 159922 199912
rect 160054 199860 160106 199912
rect 160146 199860 160198 199912
rect 160238 199860 160290 199912
rect 160330 199860 160382 199912
rect 159640 199724 159692 199776
rect 159272 199588 159324 199640
rect 159456 199588 159508 199640
rect 159732 199588 159784 199640
rect 158628 199520 158680 199572
rect 158812 199520 158864 199572
rect 160192 199724 160244 199776
rect 160284 199724 160336 199776
rect 160698 199860 160750 199912
rect 160882 199860 160934 199912
rect 161066 199860 161118 199912
rect 161158 199860 161210 199912
rect 161618 199860 161670 199912
rect 161710 199860 161762 199912
rect 161802 199860 161854 199912
rect 161894 199860 161946 199912
rect 160652 199724 160704 199776
rect 161112 199656 161164 199708
rect 160836 199588 160888 199640
rect 161020 199588 161072 199640
rect 161480 199520 161532 199572
rect 160468 199452 160520 199504
rect 161664 199724 161716 199776
rect 162078 199792 162130 199844
rect 161848 199656 161900 199708
rect 162032 199520 162084 199572
rect 162630 199860 162682 199912
rect 162722 199860 162774 199912
rect 162538 199792 162590 199844
rect 162308 199588 162360 199640
rect 162906 199860 162958 199912
rect 163090 199860 163142 199912
rect 163182 199860 163234 199912
rect 163274 199860 163326 199912
rect 163366 199860 163418 199912
rect 162768 199588 162820 199640
rect 163136 199724 163188 199776
rect 163228 199724 163280 199776
rect 163458 199792 163510 199844
rect 163826 199860 163878 199912
rect 163918 199860 163970 199912
rect 164378 199860 164430 199912
rect 163642 199792 163694 199844
rect 163412 199656 163464 199708
rect 163044 199588 163096 199640
rect 162400 199520 162452 199572
rect 162492 199520 162544 199572
rect 164470 199792 164522 199844
rect 163596 199656 163648 199708
rect 163780 199656 163832 199708
rect 164240 199656 164292 199708
rect 164332 199588 164384 199640
rect 163872 199452 163924 199504
rect 164240 199520 164292 199572
rect 164424 199520 164476 199572
rect 164148 199452 164200 199504
rect 165206 199860 165258 199912
rect 165298 199860 165350 199912
rect 165390 199860 165442 199912
rect 165482 199860 165534 199912
rect 164746 199792 164798 199844
rect 164930 199724 164982 199776
rect 165252 199724 165304 199776
rect 165160 199656 165212 199708
rect 164884 199588 164936 199640
rect 165850 199860 165902 199912
rect 165942 199860 165994 199912
rect 166034 199860 166086 199912
rect 165574 199724 165626 199776
rect 165804 199656 165856 199708
rect 165988 199656 166040 199708
rect 166494 199860 166546 199912
rect 166862 199860 166914 199912
rect 166678 199792 166730 199844
rect 166310 199724 166362 199776
rect 165436 199588 165488 199640
rect 165896 199588 165948 199640
rect 166080 199588 166132 199640
rect 166632 199588 166684 199640
rect 165528 199520 165580 199572
rect 166356 199520 166408 199572
rect 166448 199520 166500 199572
rect 167598 199860 167650 199912
rect 167690 199860 167742 199912
rect 167782 199860 167834 199912
rect 167874 199860 167926 199912
rect 167230 199792 167282 199844
rect 167414 199792 167466 199844
rect 167138 199724 167190 199776
rect 167000 199588 167052 199640
rect 167552 199656 167604 199708
rect 167644 199656 167696 199708
rect 167736 199656 167788 199708
rect 167184 199588 167236 199640
rect 167368 199588 167420 199640
rect 167828 199588 167880 199640
rect 167092 199520 167144 199572
rect 178408 200336 178460 200388
rect 177764 200268 177816 200320
rect 189264 200268 189316 200320
rect 177856 200200 177908 200252
rect 191840 200200 191892 200252
rect 178040 200132 178092 200184
rect 196348 200132 196400 200184
rect 168058 199860 168110 199912
rect 168150 199860 168202 199912
rect 168518 199860 168570 199912
rect 168794 199860 168846 199912
rect 168886 199860 168938 199912
rect 169070 199860 169122 199912
rect 169162 199860 169214 199912
rect 168426 199792 168478 199844
rect 168104 199724 168156 199776
rect 168472 199656 168524 199708
rect 169024 199724 169076 199776
rect 168840 199656 168892 199708
rect 169116 199656 169168 199708
rect 169530 199860 169582 199912
rect 169714 199860 169766 199912
rect 169806 199860 169858 199912
rect 169898 199860 169950 199912
rect 170174 199860 170226 199912
rect 169484 199724 169536 199776
rect 169852 199724 169904 199776
rect 169668 199656 169720 199708
rect 169760 199656 169812 199708
rect 169300 199588 169352 199640
rect 170450 199792 170502 199844
rect 171002 199860 171054 199912
rect 171186 199860 171238 199912
rect 171370 199860 171422 199912
rect 171462 199860 171514 199912
rect 171554 199860 171606 199912
rect 171646 199860 171698 199912
rect 171922 199860 171974 199912
rect 172198 199860 172250 199912
rect 172290 199860 172342 199912
rect 172658 199860 172710 199912
rect 172842 199860 172894 199912
rect 173578 199860 173630 199912
rect 174038 199860 174090 199912
rect 174590 199860 174642 199912
rect 174682 199860 174734 199912
rect 174866 199860 174918 199912
rect 175234 199860 175286 199912
rect 170726 199792 170778 199844
rect 170818 199792 170870 199844
rect 170910 199792 170962 199844
rect 170312 199588 170364 199640
rect 170496 199588 170548 199640
rect 168564 199520 168616 199572
rect 167920 199452 167972 199504
rect 168288 199452 168340 199504
rect 170772 199588 170824 199640
rect 170956 199588 171008 199640
rect 171140 199588 171192 199640
rect 170680 199520 170732 199572
rect 171416 199656 171468 199708
rect 171508 199656 171560 199708
rect 170864 199452 170916 199504
rect 171324 199452 171376 199504
rect 172336 199724 172388 199776
rect 172244 199656 172296 199708
rect 172704 199656 172756 199708
rect 172060 199588 172112 199640
rect 172612 199588 172664 199640
rect 174084 199724 174136 199776
rect 173808 199520 173860 199572
rect 174636 199656 174688 199708
rect 175188 199724 175240 199776
rect 175096 199588 175148 199640
rect 175418 199860 175470 199912
rect 175510 199860 175562 199912
rect 175878 199860 175930 199912
rect 176062 199860 176114 199912
rect 176246 199860 176298 199912
rect 176338 199860 176390 199912
rect 176798 199860 176850 199912
rect 177074 199860 177126 199912
rect 177166 199860 177218 199912
rect 177258 199860 177310 199912
rect 177350 199860 177402 199912
rect 177856 199860 177908 199912
rect 175464 199656 175516 199708
rect 175740 199588 175792 199640
rect 175924 199588 175976 199640
rect 174912 199520 174964 199572
rect 175280 199452 175332 199504
rect 176292 199724 176344 199776
rect 176844 199520 176896 199572
rect 176660 199452 176712 199504
rect 186688 199860 186740 199912
rect 187608 199792 187660 199844
rect 177120 199588 177172 199640
rect 177212 199588 177264 199640
rect 177396 199588 177448 199640
rect 215668 199588 215720 199640
rect 178592 199520 178644 199572
rect 215392 199520 215444 199572
rect 177304 199452 177356 199504
rect 152924 199384 152976 199436
rect 153108 199384 153160 199436
rect 156420 199384 156472 199436
rect 158352 199384 158404 199436
rect 178684 199384 178736 199436
rect 182824 199384 182876 199436
rect 190460 199384 190512 199436
rect 152556 199316 152608 199368
rect 160100 199316 160152 199368
rect 153568 199248 153620 199300
rect 156788 199248 156840 199300
rect 152004 199180 152056 199232
rect 215484 199316 215536 199368
rect 164424 199248 164476 199300
rect 198740 199248 198792 199300
rect 116952 198976 117004 199028
rect 145932 198976 145984 199028
rect 115664 198908 115716 198960
rect 147036 198908 147088 198960
rect 155132 198908 155184 198960
rect 190000 199180 190052 199232
rect 170128 199112 170180 199164
rect 200304 199112 200356 199164
rect 178408 199044 178460 199096
rect 203156 199044 203208 199096
rect 161940 198976 161992 199028
rect 196164 198976 196216 199028
rect 168380 198908 168432 198960
rect 180156 198908 180208 198960
rect 126428 198840 126480 198892
rect 144920 198840 144972 198892
rect 161480 198840 161532 198892
rect 178868 198840 178920 198892
rect 121184 198772 121236 198824
rect 139492 198772 139544 198824
rect 141148 198772 141200 198824
rect 141700 198772 141752 198824
rect 143908 198772 143960 198824
rect 144092 198772 144144 198824
rect 158076 198772 158128 198824
rect 178776 198772 178828 198824
rect 129096 198704 129148 198756
rect 149152 198704 149204 198756
rect 162584 198704 162636 198756
rect 185584 198772 185636 198824
rect 181076 198704 181128 198756
rect 187700 198704 187752 198756
rect 125876 198636 125928 198688
rect 130752 198636 130804 198688
rect 132500 198636 132552 198688
rect 146208 198636 146260 198688
rect 167460 198636 167512 198688
rect 122196 198568 122248 198620
rect 146852 198568 146904 198620
rect 164976 198568 165028 198620
rect 167920 198568 167972 198620
rect 169944 198568 169996 198620
rect 173900 198636 173952 198688
rect 202512 198636 202564 198688
rect 129280 198500 129332 198552
rect 154672 198500 154724 198552
rect 158996 198500 159048 198552
rect 165620 198500 165672 198552
rect 166448 198500 166500 198552
rect 166816 198500 166868 198552
rect 105820 198432 105872 198484
rect 132408 198432 132460 198484
rect 142436 198432 142488 198484
rect 143908 198432 143960 198484
rect 159732 198432 159784 198484
rect 172520 198500 172572 198552
rect 201592 198568 201644 198620
rect 174360 198500 174412 198552
rect 207112 198500 207164 198552
rect 208584 198432 208636 198484
rect 122288 198364 122340 198416
rect 149428 198364 149480 198416
rect 165528 198364 165580 198416
rect 171600 198364 171652 198416
rect 172060 198364 172112 198416
rect 107108 198296 107160 198348
rect 136088 198296 136140 198348
rect 163136 198296 163188 198348
rect 171048 198296 171100 198348
rect 172428 198296 172480 198348
rect 174820 198296 174872 198348
rect 175648 198364 175700 198416
rect 212816 198364 212868 198416
rect 211344 198296 211396 198348
rect 110328 198228 110380 198280
rect 143356 198228 143408 198280
rect 165712 198228 165764 198280
rect 167460 198228 167512 198280
rect 170588 198228 170640 198280
rect 209964 198228 210016 198280
rect 107200 198160 107252 198212
rect 137008 198160 137060 198212
rect 155592 198160 155644 198212
rect 171140 198160 171192 198212
rect 172796 198160 172848 198212
rect 212908 198160 212960 198212
rect 110236 198092 110288 198144
rect 144736 198092 144788 198144
rect 162768 198092 162820 198144
rect 163320 198092 163372 198144
rect 165620 198092 165672 198144
rect 172060 198092 172112 198144
rect 172336 198092 172388 198144
rect 212724 198092 212776 198144
rect 108672 198024 108724 198076
rect 142068 198024 142120 198076
rect 156604 198024 156656 198076
rect 165712 198024 165764 198076
rect 166080 198024 166132 198076
rect 166448 198024 166500 198076
rect 171324 198024 171376 198076
rect 213000 198024 213052 198076
rect 126520 197956 126572 198008
rect 132500 197956 132552 198008
rect 155316 197956 155368 198008
rect 164976 197956 165028 198008
rect 165620 197956 165672 198008
rect 165988 197956 166040 198008
rect 167460 197956 167512 198008
rect 133880 197888 133932 197940
rect 150716 197888 150768 197940
rect 154856 197888 154908 197940
rect 169300 197956 169352 198008
rect 209780 197956 209832 198008
rect 127716 197820 127768 197872
rect 144184 197820 144236 197872
rect 156512 197820 156564 197872
rect 158076 197820 158128 197872
rect 159180 197820 159232 197872
rect 161296 197820 161348 197872
rect 162952 197820 163004 197872
rect 163228 197820 163280 197872
rect 167092 197820 167144 197872
rect 167460 197820 167512 197872
rect 170772 197888 170824 197940
rect 171140 197888 171192 197940
rect 172336 197888 172388 197940
rect 172612 197888 172664 197940
rect 172888 197888 172940 197940
rect 177120 197888 177172 197940
rect 177764 197888 177816 197940
rect 174636 197820 174688 197872
rect 127808 197752 127860 197804
rect 143540 197752 143592 197804
rect 97632 197684 97684 197736
rect 130660 197684 130712 197736
rect 133880 197684 133932 197736
rect 131856 197616 131908 197668
rect 136732 197616 136784 197668
rect 143540 197616 143592 197668
rect 143724 197616 143776 197668
rect 148048 197616 148100 197668
rect 148324 197616 148376 197668
rect 157524 197616 157576 197668
rect 172152 197752 172204 197804
rect 172520 197752 172572 197804
rect 178132 197752 178184 197804
rect 137652 197548 137704 197600
rect 161848 197548 161900 197600
rect 173072 197684 173124 197736
rect 168288 197616 168340 197668
rect 179420 197616 179472 197668
rect 125140 197480 125192 197532
rect 133328 197480 133380 197532
rect 156236 197480 156288 197532
rect 159180 197480 159232 197532
rect 161296 197480 161348 197532
rect 173808 197480 173860 197532
rect 132868 197412 132920 197464
rect 133512 197412 133564 197464
rect 134248 197412 134300 197464
rect 135168 197412 135220 197464
rect 145196 197412 145248 197464
rect 149428 197412 149480 197464
rect 159548 197412 159600 197464
rect 172428 197412 172480 197464
rect 173992 197412 174044 197464
rect 178960 197412 179012 197464
rect 134156 197344 134208 197396
rect 134616 197344 134668 197396
rect 143908 197344 143960 197396
rect 144552 197344 144604 197396
rect 121000 197276 121052 197328
rect 146760 197276 146812 197328
rect 155868 197276 155920 197328
rect 165344 197276 165396 197328
rect 121092 197208 121144 197260
rect 149888 197208 149940 197260
rect 163872 197208 163924 197260
rect 171324 197208 171376 197260
rect 172060 197208 172112 197260
rect 193404 197208 193456 197260
rect 114284 197140 114336 197192
rect 144368 197140 144420 197192
rect 166908 197140 166960 197192
rect 170404 197140 170456 197192
rect 171048 197140 171100 197192
rect 194876 197140 194928 197192
rect 116860 197072 116912 197124
rect 147588 197072 147640 197124
rect 157248 197072 157300 197124
rect 158720 197072 158772 197124
rect 160836 197072 160888 197124
rect 194600 197072 194652 197124
rect 107016 197004 107068 197056
rect 137468 197004 137520 197056
rect 148508 197004 148560 197056
rect 149796 197004 149848 197056
rect 167920 197004 167972 197056
rect 198832 197004 198884 197056
rect 112720 196936 112772 196988
rect 132960 196936 133012 196988
rect 140872 196936 140924 196988
rect 141148 196936 141200 196988
rect 171600 196936 171652 196988
rect 198924 196936 198976 196988
rect 111708 196868 111760 196920
rect 143816 196868 143868 196920
rect 167184 196868 167236 196920
rect 201684 196868 201736 196920
rect 114192 196800 114244 196852
rect 147312 196800 147364 196852
rect 155960 196800 156012 196852
rect 109868 196732 109920 196784
rect 133236 196732 133288 196784
rect 146300 196732 146352 196784
rect 146484 196732 146536 196784
rect 114468 196664 114520 196716
rect 147680 196664 147732 196716
rect 105912 196596 105964 196648
rect 138756 196596 138808 196648
rect 141884 196596 141936 196648
rect 142252 196596 142304 196648
rect 164148 196800 164200 196852
rect 170588 196800 170640 196852
rect 171232 196800 171284 196852
rect 171600 196800 171652 196852
rect 172520 196800 172572 196852
rect 200488 196800 200540 196852
rect 163596 196732 163648 196784
rect 197636 196732 197688 196784
rect 169852 196664 169904 196716
rect 170220 196664 170272 196716
rect 170588 196664 170640 196716
rect 197728 196664 197780 196716
rect 190644 196596 190696 196648
rect 129464 196528 129516 196580
rect 149980 196528 150032 196580
rect 158628 196528 158680 196580
rect 160284 196528 160336 196580
rect 164700 196528 164752 196580
rect 164884 196528 164936 196580
rect 171324 196528 171376 196580
rect 179052 196528 179104 196580
rect 132776 196460 132828 196512
rect 133788 196460 133840 196512
rect 134156 196460 134208 196512
rect 135076 196460 135128 196512
rect 137284 196460 137336 196512
rect 139400 196460 139452 196512
rect 131764 196392 131816 196444
rect 139676 196392 139728 196444
rect 129372 196324 129424 196376
rect 147864 196324 147916 196376
rect 167736 196324 167788 196376
rect 180524 196324 180576 196376
rect 133236 196256 133288 196308
rect 142804 196256 142856 196308
rect 132960 196188 133012 196240
rect 144092 196188 144144 196240
rect 129740 196120 129792 196172
rect 134708 196120 134760 196172
rect 132132 195984 132184 196036
rect 133144 195984 133196 196036
rect 134524 195984 134576 196036
rect 134984 195984 135036 196036
rect 120632 195916 120684 195968
rect 144828 195916 144880 195968
rect 152188 195916 152240 195968
rect 152832 195916 152884 195968
rect 157800 195916 157852 195968
rect 115204 195848 115256 195900
rect 146116 195848 146168 195900
rect 154488 195848 154540 195900
rect 114100 195780 114152 195832
rect 145472 195780 145524 195832
rect 154764 195780 154816 195832
rect 159456 195848 159508 195900
rect 115756 195712 115808 195764
rect 109960 195644 110012 195696
rect 143172 195644 143224 195696
rect 111616 195576 111668 195628
rect 145840 195576 145892 195628
rect 108856 195508 108908 195560
rect 143448 195508 143500 195560
rect 157616 195712 157668 195764
rect 162124 195916 162176 195968
rect 171876 195916 171928 195968
rect 173808 195916 173860 195968
rect 176936 195984 176988 196036
rect 176200 195848 176252 195900
rect 192208 195916 192260 195968
rect 198188 195848 198240 195900
rect 175004 195780 175056 195832
rect 181352 195780 181404 195832
rect 174360 195712 174412 195764
rect 176292 195712 176344 195764
rect 201040 195712 201092 195764
rect 186596 195644 186648 195696
rect 153936 195576 153988 195628
rect 188712 195576 188764 195628
rect 148968 195508 149020 195560
rect 151912 195508 151964 195560
rect 152280 195508 152332 195560
rect 160468 195508 160520 195560
rect 193312 195508 193364 195560
rect 104624 195440 104676 195492
rect 132592 195440 132644 195492
rect 132684 195440 132736 195492
rect 133420 195440 133472 195492
rect 135812 195440 135864 195492
rect 136272 195440 136324 195492
rect 149336 195440 149388 195492
rect 149980 195440 150032 195492
rect 150716 195440 150768 195492
rect 151084 195440 151136 195492
rect 152004 195440 152056 195492
rect 152464 195440 152516 195492
rect 156696 195440 156748 195492
rect 111156 195372 111208 195424
rect 145288 195372 145340 195424
rect 153476 195372 153528 195424
rect 154212 195372 154264 195424
rect 158076 195440 158128 195492
rect 173256 195440 173308 195492
rect 181352 195440 181404 195492
rect 208676 195440 208728 195492
rect 190552 195372 190604 195424
rect 112812 195304 112864 195356
rect 146300 195304 146352 195356
rect 149336 195304 149388 195356
rect 149704 195304 149756 195356
rect 150624 195304 150676 195356
rect 151084 195304 151136 195356
rect 153568 195304 153620 195356
rect 154304 195304 154356 195356
rect 111340 195236 111392 195288
rect 145012 195236 145064 195288
rect 149060 195236 149112 195288
rect 149520 195236 149572 195288
rect 150532 195236 150584 195288
rect 150900 195236 150952 195288
rect 151268 195236 151320 195288
rect 151636 195236 151688 195288
rect 153476 195236 153528 195288
rect 154028 195236 154080 195288
rect 155960 195236 156012 195288
rect 156880 195236 156932 195288
rect 126704 195168 126756 195220
rect 145748 195168 145800 195220
rect 153292 195168 153344 195220
rect 153844 195168 153896 195220
rect 154120 195168 154172 195220
rect 188436 195304 188488 195356
rect 157616 195236 157668 195288
rect 162124 195236 162176 195288
rect 130384 195100 130436 195152
rect 147220 195100 147272 195152
rect 152372 195100 152424 195152
rect 153108 195100 153160 195152
rect 153384 195100 153436 195152
rect 154396 195100 154448 195152
rect 155408 195100 155460 195152
rect 155684 195100 155736 195152
rect 135536 195032 135588 195084
rect 136088 195032 136140 195084
rect 136732 195032 136784 195084
rect 137468 195032 137520 195084
rect 135720 194964 135772 195016
rect 136456 194964 136508 195016
rect 152832 194964 152884 195016
rect 211528 195236 211580 195288
rect 169576 195100 169628 195152
rect 182916 195100 182968 195152
rect 172612 194964 172664 195016
rect 172980 194964 173032 195016
rect 131948 194828 132000 194880
rect 139308 194896 139360 194948
rect 172336 194896 172388 194948
rect 190092 195168 190144 195220
rect 135444 194828 135496 194880
rect 136364 194828 136416 194880
rect 171876 194828 171928 194880
rect 179144 194828 179196 194880
rect 132592 194760 132644 194812
rect 139124 194760 139176 194812
rect 126244 194692 126296 194744
rect 131120 194692 131172 194744
rect 122104 194488 122156 194540
rect 148048 194488 148100 194540
rect 168656 194488 168708 194540
rect 202880 194488 202932 194540
rect 103336 194420 103388 194472
rect 127900 194420 127952 194472
rect 135352 194420 135404 194472
rect 136180 194420 136232 194472
rect 169116 194420 169168 194472
rect 202972 194420 203024 194472
rect 102968 194352 103020 194404
rect 134892 194352 134944 194404
rect 168472 194352 168524 194404
rect 168656 194352 168708 194404
rect 173532 194352 173584 194404
rect 207204 194352 207256 194404
rect 103244 194284 103296 194336
rect 124772 194284 124824 194336
rect 174544 194284 174596 194336
rect 208492 194284 208544 194336
rect 107384 194216 107436 194268
rect 140044 194216 140096 194268
rect 175464 194216 175516 194268
rect 210148 194216 210200 194268
rect 108948 194148 109000 194200
rect 143080 194148 143132 194200
rect 177856 194148 177908 194200
rect 211620 194148 211672 194200
rect 110144 194080 110196 194132
rect 143540 194080 143592 194132
rect 163964 194080 164016 194132
rect 164148 194080 164200 194132
rect 170680 194080 170732 194132
rect 204720 194080 204772 194132
rect 105728 194012 105780 194064
rect 140412 194012 140464 194064
rect 172796 194012 172848 194064
rect 207480 194012 207532 194064
rect 104256 193944 104308 193996
rect 139032 193944 139084 193996
rect 157432 193944 157484 193996
rect 157892 193944 157944 193996
rect 174268 193944 174320 193996
rect 208860 193944 208912 193996
rect 97908 193876 97960 193928
rect 141332 193876 141384 193928
rect 150716 193876 150768 193928
rect 151176 193876 151228 193928
rect 97816 193808 97868 193860
rect 143908 193808 143960 193860
rect 155500 193808 155552 193860
rect 174544 193876 174596 193928
rect 181352 193876 181404 193928
rect 208952 193876 209004 193928
rect 155040 193740 155092 193792
rect 174544 193740 174596 193792
rect 175280 193740 175332 193792
rect 175740 193740 175792 193792
rect 183192 193808 183244 193860
rect 216772 193808 216824 193860
rect 153200 193672 153252 193724
rect 181536 193672 181588 193724
rect 156052 193604 156104 193656
rect 181628 193604 181680 193656
rect 173992 193536 174044 193588
rect 181352 193536 181404 193588
rect 130568 193128 130620 193180
rect 148692 193128 148744 193180
rect 160468 193128 160520 193180
rect 160652 193128 160704 193180
rect 176660 193128 176712 193180
rect 177028 193128 177080 193180
rect 188344 193128 188396 193180
rect 580172 193128 580224 193180
rect 102784 193060 102836 193112
rect 129740 193060 129792 193112
rect 170312 193060 170364 193112
rect 204444 193060 204496 193112
rect 101680 192992 101732 193044
rect 130936 192992 130988 193044
rect 171600 192992 171652 193044
rect 205916 192992 205968 193044
rect 117044 192924 117096 192976
rect 146944 192924 146996 192976
rect 171508 192924 171560 192976
rect 206008 192924 206060 192976
rect 108764 192856 108816 192908
rect 140596 192856 140648 192908
rect 170220 192856 170272 192908
rect 204628 192856 204680 192908
rect 115112 192788 115164 192840
rect 147496 192788 147548 192840
rect 172704 192788 172756 192840
rect 207572 192788 207624 192840
rect 116216 192720 116268 192772
rect 150072 192720 150124 192772
rect 173164 192720 173216 192772
rect 207664 192720 207716 192772
rect 123944 192652 123996 192704
rect 157156 192652 157208 192704
rect 160836 192652 160888 192704
rect 208768 192652 208820 192704
rect 99104 192584 99156 192636
rect 133328 192584 133380 192636
rect 159180 192584 159232 192636
rect 211252 192584 211304 192636
rect 108304 192516 108356 192568
rect 142896 192516 142948 192568
rect 157984 192516 158036 192568
rect 211160 192516 211212 192568
rect 108396 192448 108448 192500
rect 142620 192448 142672 192500
rect 155776 192448 155828 192500
rect 210700 192448 210752 192500
rect 130844 192380 130896 192432
rect 148508 192380 148560 192432
rect 174820 192380 174872 192432
rect 205640 192380 205692 192432
rect 162584 192312 162636 192364
rect 191104 192312 191156 192364
rect 177948 192244 178000 192296
rect 189172 192244 189224 192296
rect 162676 192176 162728 192228
rect 162952 192176 163004 192228
rect 137008 192108 137060 192160
rect 137928 192108 137980 192160
rect 167368 191768 167420 191820
rect 201500 191768 201552 191820
rect 166080 191700 166132 191752
rect 166908 191700 166960 191752
rect 168564 191700 168616 191752
rect 159272 191632 159324 191684
rect 166632 191632 166684 191684
rect 173900 191632 173952 191684
rect 174912 191632 174964 191684
rect 175096 191700 175148 191752
rect 201776 191700 201828 191752
rect 203248 191632 203300 191684
rect 163780 191564 163832 191616
rect 204352 191564 204404 191616
rect 142436 191496 142488 191548
rect 142988 191496 143040 191548
rect 164700 191496 164752 191548
rect 205732 191496 205784 191548
rect 122472 191428 122524 191480
rect 151452 191428 151504 191480
rect 159916 191428 159968 191480
rect 106096 191360 106148 191412
rect 137744 191360 137796 191412
rect 159364 191360 159416 191412
rect 108580 191292 108632 191344
rect 141240 191292 141292 191344
rect 104164 191224 104216 191276
rect 137560 191224 137612 191276
rect 142528 191224 142580 191276
rect 142988 191224 143040 191276
rect 160284 191224 160336 191276
rect 161296 191224 161348 191276
rect 166540 191428 166592 191480
rect 207388 191428 207440 191480
rect 167184 191360 167236 191412
rect 167552 191360 167604 191412
rect 174176 191360 174228 191412
rect 174728 191360 174780 191412
rect 175004 191360 175056 191412
rect 209044 191360 209096 191412
rect 207296 191292 207348 191344
rect 216864 191224 216916 191276
rect 99196 191156 99248 191208
rect 132868 191156 132920 191208
rect 106924 191088 106976 191140
rect 140872 191156 140924 191208
rect 160192 191156 160244 191208
rect 160468 191156 160520 191208
rect 161572 191156 161624 191208
rect 161756 191156 161808 191208
rect 163136 191156 163188 191208
rect 163504 191156 163556 191208
rect 164240 191156 164292 191208
rect 165252 191156 165304 191208
rect 165712 191156 165764 191208
rect 166356 191156 166408 191208
rect 166632 191156 166684 191208
rect 218152 191156 218204 191208
rect 138296 191088 138348 191140
rect 139216 191088 139268 191140
rect 139952 191088 140004 191140
rect 140688 191088 140740 191140
rect 141332 191088 141384 191140
rect 141976 191088 142028 191140
rect 145380 191088 145432 191140
rect 146024 191088 146076 191140
rect 146668 191088 146720 191140
rect 147404 191088 147456 191140
rect 151728 191088 151780 191140
rect 218244 191088 218296 191140
rect 146392 191020 146444 191072
rect 147036 191020 147088 191072
rect 157524 191020 157576 191072
rect 158444 191020 158496 191072
rect 160192 191020 160244 191072
rect 161204 191020 161256 191072
rect 161572 191020 161624 191072
rect 162032 191020 162084 191072
rect 163412 191020 163464 191072
rect 164056 191020 164108 191072
rect 164608 191020 164660 191072
rect 165068 191020 165120 191072
rect 165896 191020 165948 191072
rect 166724 191020 166776 191072
rect 164332 190952 164384 191004
rect 164792 190952 164844 191004
rect 165620 190952 165672 191004
rect 200120 191020 200172 191072
rect 167000 190952 167052 191004
rect 167828 190952 167880 191004
rect 168564 190952 168616 191004
rect 168932 190952 168984 191004
rect 169852 190952 169904 191004
rect 170588 190952 170640 191004
rect 171140 190952 171192 191004
rect 171968 190952 172020 191004
rect 172704 190952 172756 191004
rect 173624 190952 173676 191004
rect 173992 190952 174044 191004
rect 174452 190952 174504 191004
rect 175556 190952 175608 191004
rect 176108 190952 176160 191004
rect 165804 190884 165856 190936
rect 166172 190884 166224 190936
rect 167092 190884 167144 190936
rect 168288 190884 168340 190936
rect 169760 190884 169812 190936
rect 170864 190884 170916 190936
rect 171232 190884 171284 190936
rect 172244 190884 172296 190936
rect 176936 190884 176988 190936
rect 177672 190884 177724 190936
rect 167460 190816 167512 190868
rect 175096 190816 175148 190868
rect 176844 190816 176896 190868
rect 177396 190816 177448 190868
rect 167644 190748 167696 190800
rect 175004 190748 175056 190800
rect 148140 190544 148192 190596
rect 148784 190544 148836 190596
rect 156144 190544 156196 190596
rect 157064 190544 157116 190596
rect 167920 190408 167972 190460
rect 185768 190408 185820 190460
rect 162400 190340 162452 190392
rect 183100 190340 183152 190392
rect 125324 190272 125376 190324
rect 139860 190272 139912 190324
rect 160008 190272 160060 190324
rect 185676 190272 185728 190324
rect 104716 190204 104768 190256
rect 137468 190204 137520 190256
rect 153660 190204 153712 190256
rect 181720 190204 181772 190256
rect 103428 190136 103480 190188
rect 135444 190136 135496 190188
rect 152372 190136 152424 190188
rect 183008 190136 183060 190188
rect 111524 190068 111576 190120
rect 144460 190068 144512 190120
rect 177120 190068 177172 190120
rect 210240 190068 210292 190120
rect 111064 190000 111116 190052
rect 144092 190000 144144 190052
rect 176476 190000 176528 190052
rect 210332 190000 210384 190052
rect 104072 189932 104124 189984
rect 136916 189932 136968 189984
rect 176016 189932 176068 189984
rect 210424 189932 210476 189984
rect 103060 189864 103112 189916
rect 137192 189864 137244 189916
rect 177212 189864 177264 189916
rect 211896 189864 211948 189916
rect 101588 189796 101640 189848
rect 135352 189796 135404 189848
rect 158536 189796 158588 189848
rect 212540 189796 212592 189848
rect 109684 189728 109736 189780
rect 144276 189728 144328 189780
rect 152280 189728 152332 189780
rect 218336 189728 218388 189780
rect 172520 189592 172572 189644
rect 173348 189592 173400 189644
rect 3424 188980 3476 189032
rect 120540 188980 120592 189032
rect 175372 188572 175424 188624
rect 175648 188572 175700 188624
rect 175372 188436 175424 188488
rect 176384 188436 176436 188488
rect 169944 188368 169996 188420
rect 170312 188368 170364 188420
rect 121828 187484 121880 187536
rect 149244 187484 149296 187536
rect 109776 187416 109828 187468
rect 140504 187416 140556 187468
rect 109592 187348 109644 187400
rect 141884 187348 141936 187400
rect 169024 187348 169076 187400
rect 103152 187280 103204 187332
rect 135904 187280 135956 187332
rect 168472 187280 168524 187332
rect 169668 187280 169720 187332
rect 203340 187280 203392 187332
rect 100484 187212 100536 187264
rect 132776 187212 132828 187264
rect 153568 187212 153620 187264
rect 214012 187212 214064 187264
rect 101496 187144 101548 187196
rect 134524 187144 134576 187196
rect 149796 187144 149848 187196
rect 211436 187144 211488 187196
rect 99012 187076 99064 187128
rect 133144 187076 133196 187128
rect 149336 187076 149388 187128
rect 211712 187076 211764 187128
rect 100300 187008 100352 187060
rect 135076 187008 135128 187060
rect 151084 187008 151136 187060
rect 215852 187008 215904 187060
rect 100392 186940 100444 186992
rect 134248 186940 134300 186992
rect 150992 186940 151044 186992
rect 218428 186940 218480 186992
rect 188344 178032 188396 178084
rect 580172 178032 580224 178084
rect 189908 165588 189960 165640
rect 580172 165588 580224 165640
rect 98920 164840 98972 164892
rect 130660 164840 130712 164892
rect 175740 159740 175792 159792
rect 199200 159740 199252 159792
rect 172796 159672 172848 159724
rect 196624 159672 196676 159724
rect 161848 159604 161900 159656
rect 195152 159604 195204 159656
rect 172612 159536 172664 159588
rect 211988 159536 212040 159588
rect 149980 159468 150032 159520
rect 209136 159468 209188 159520
rect 152096 159400 152148 159452
rect 213920 159400 213972 159452
rect 152188 159332 152240 159384
rect 214196 159332 214248 159384
rect 177856 157292 177908 157344
rect 203432 157292 203484 157344
rect 163596 157224 163648 157276
rect 192392 157224 192444 157276
rect 161940 157156 161992 157208
rect 193772 157156 193824 157208
rect 176936 157088 176988 157140
rect 210608 157088 210660 157140
rect 168564 157020 168616 157072
rect 203800 157020 203852 157072
rect 167276 156952 167328 157004
rect 201960 156952 202012 157004
rect 168656 156884 168708 156936
rect 203432 156884 203484 156936
rect 167184 156816 167236 156868
rect 202144 156816 202196 156868
rect 164884 156748 164936 156800
rect 201868 156748 201920 156800
rect 160744 156680 160796 156732
rect 200580 156680 200632 156732
rect 155868 156612 155920 156664
rect 200948 156612 201000 156664
rect 163504 156544 163556 156596
rect 188252 156544 188304 156596
rect 166264 156476 166316 156528
rect 189724 156476 189776 156528
rect 165896 154504 165948 154556
rect 185860 154504 185912 154556
rect 160652 154436 160704 154488
rect 185952 154436 186004 154488
rect 158904 154368 158956 154420
rect 184296 154368 184348 154420
rect 158996 154300 159048 154352
rect 183744 154300 183796 154352
rect 157524 154232 157576 154284
rect 186136 154232 186188 154284
rect 157616 154164 157668 154216
rect 186044 154164 186096 154216
rect 157248 154096 157300 154148
rect 186228 154096 186280 154148
rect 164792 154028 164844 154080
rect 199200 154028 199252 154080
rect 165988 153960 166040 154012
rect 200580 153960 200632 154012
rect 166908 153892 166960 153944
rect 200672 153892 200724 153944
rect 121920 153824 121972 153876
rect 143632 153824 143684 153876
rect 146208 153824 146260 153876
rect 202052 153824 202104 153876
rect 166172 153756 166224 153808
rect 183284 153756 183336 153808
rect 164700 152736 164752 152788
rect 206192 152736 206244 152788
rect 154856 152668 154908 152720
rect 203064 152668 203116 152720
rect 163412 152600 163464 152652
rect 213092 152600 213144 152652
rect 121644 152532 121696 152584
rect 150900 152532 150952 152584
rect 153568 152532 153620 152584
rect 204536 152532 204588 152584
rect 121552 152464 121604 152516
rect 150808 152464 150860 152516
rect 155684 152464 155736 152516
rect 214288 152464 214340 152516
rect 185492 152396 185544 152448
rect 185676 152396 185728 152448
rect 188252 151784 188304 151836
rect 579988 151784 580040 151836
rect 99840 151716 99892 151768
rect 132684 151716 132736 151768
rect 100116 151648 100168 151700
rect 134340 151648 134392 151700
rect 100208 151580 100260 151632
rect 134432 151580 134484 151632
rect 164608 151580 164660 151632
rect 181812 151580 181864 151632
rect 98828 151512 98880 151564
rect 133052 151512 133104 151564
rect 161756 151512 161808 151564
rect 185400 151512 185452 151564
rect 100024 151444 100076 151496
rect 134616 151444 134668 151496
rect 157432 151444 157484 151496
rect 184388 151444 184440 151496
rect 101404 151376 101456 151428
rect 135628 151376 135680 151428
rect 157340 151376 157392 151428
rect 184848 151376 184900 151428
rect 101312 151308 101364 151360
rect 135536 151308 135588 151360
rect 175556 151308 175608 151360
rect 205088 151308 205140 151360
rect 99932 151240 99984 151292
rect 134156 151240 134208 151292
rect 175648 151240 175700 151292
rect 206376 151240 206428 151292
rect 122012 151172 122064 151224
rect 158720 151172 158772 151224
rect 174176 151172 174228 151224
rect 204996 151172 205048 151224
rect 122380 151104 122432 151156
rect 160100 151104 160152 151156
rect 176752 151104 176804 151156
rect 207756 151104 207808 151156
rect 97448 151036 97500 151088
rect 141148 151036 141200 151088
rect 174084 151036 174136 151088
rect 206284 151036 206336 151088
rect 102600 150968 102652 151020
rect 135996 150968 136048 151020
rect 123668 150900 123720 150952
rect 138388 150900 138440 150952
rect 172244 150356 172296 150408
rect 192760 150356 192812 150408
rect 173256 150288 173308 150340
rect 196716 150288 196768 150340
rect 158904 150220 158956 150272
rect 188160 150220 188212 150272
rect 163136 150152 163188 150204
rect 195152 150152 195204 150204
rect 167000 150084 167052 150136
rect 200856 150084 200908 150136
rect 163228 150016 163280 150068
rect 198280 150016 198332 150068
rect 164424 149948 164476 150000
rect 199752 149948 199804 150000
rect 163320 149880 163372 149932
rect 198464 149880 198516 149932
rect 165804 149812 165856 149864
rect 200764 149812 200816 149864
rect 164516 149744 164568 149796
rect 199476 149744 199528 149796
rect 158628 149676 158680 149728
rect 195520 149676 195572 149728
rect 165528 149608 165580 149660
rect 182088 149608 182140 149660
rect 180892 149540 180944 149592
rect 198096 149540 198148 149592
rect 3148 149132 3200 149184
rect 180892 149132 180944 149184
rect 119344 149064 119396 149116
rect 580540 149064 580592 149116
rect 112536 148996 112588 149048
rect 142528 148996 142580 149048
rect 112076 148928 112128 148980
rect 142436 148928 142488 148980
rect 112168 148860 112220 148912
rect 143908 148860 143960 148912
rect 162676 148860 162728 148912
rect 188620 148860 188672 148912
rect 110788 148792 110840 148844
rect 142620 148792 142672 148844
rect 156144 148792 156196 148844
rect 184572 148792 184624 148844
rect 118976 148724 119028 148776
rect 150624 148724 150676 148776
rect 170036 148724 170088 148776
rect 199292 148724 199344 148776
rect 117688 148656 117740 148708
rect 150716 148656 150768 148708
rect 173808 148656 173860 148708
rect 204536 148656 204588 148708
rect 114836 148588 114888 148640
rect 149520 148588 149572 148640
rect 171232 148588 171284 148640
rect 202236 148588 202288 148640
rect 98736 148520 98788 148572
rect 132960 148520 133012 148572
rect 171416 148520 171468 148572
rect 203524 148520 203576 148572
rect 101220 148452 101272 148504
rect 135720 148452 135772 148504
rect 171324 148452 171376 148504
rect 203708 148452 203760 148504
rect 97540 148384 97592 148436
rect 141056 148384 141108 148436
rect 173992 148384 174044 148436
rect 206468 148384 206520 148436
rect 113640 148316 113692 148368
rect 128636 148316 128688 148368
rect 188252 148316 188304 148368
rect 115572 148248 115624 148300
rect 115848 148248 115900 148300
rect 113456 148112 113508 148164
rect 142988 148248 143040 148300
rect 105452 148044 105504 148096
rect 131856 148044 131908 148096
rect 124036 147636 124088 147688
rect 580448 147636 580500 147688
rect 126796 147568 126848 147620
rect 140136 147568 140188 147620
rect 179052 147568 179104 147620
rect 196992 147568 197044 147620
rect 123484 147500 123536 147552
rect 140320 147500 140372 147552
rect 174728 147500 174780 147552
rect 194140 147500 194192 147552
rect 112444 147432 112496 147484
rect 131764 147432 131816 147484
rect 164148 147432 164200 147484
rect 181904 147432 181956 147484
rect 110972 147364 111024 147416
rect 131948 147364 132000 147416
rect 160376 147364 160428 147416
rect 188160 147364 188212 147416
rect 118884 147296 118936 147348
rect 141332 147296 141384 147348
rect 164056 147296 164108 147348
rect 192852 147296 192904 147348
rect 121920 147228 121972 147280
rect 145564 147228 145616 147280
rect 160008 147228 160060 147280
rect 191380 147228 191432 147280
rect 108120 147160 108172 147212
rect 138572 147160 138624 147212
rect 160560 147160 160612 147212
rect 193864 147160 193916 147212
rect 109500 147092 109552 147144
rect 141700 147092 141752 147144
rect 158812 147092 158864 147144
rect 192392 147092 192444 147144
rect 105360 147024 105412 147076
rect 138664 147024 138716 147076
rect 160468 147024 160520 147076
rect 195244 147024 195296 147076
rect 112628 146956 112680 147008
rect 112904 146956 112956 147008
rect 106740 146888 106792 146940
rect 141884 146956 141936 147008
rect 161664 146956 161716 147008
rect 197176 146956 197228 147008
rect 103980 146820 104032 146872
rect 138848 146888 138900 146940
rect 174912 146888 174964 146940
rect 214472 146888 214524 146940
rect 126612 146820 126664 146872
rect 126888 146820 126940 146872
rect 179144 146820 179196 146872
rect 185768 146820 185820 146872
rect 186044 146820 186096 146872
rect 181720 146752 181772 146804
rect 187240 146752 187292 146804
rect 183192 146684 183244 146736
rect 189724 146684 189776 146736
rect 189172 146616 189224 146668
rect 181628 146548 181680 146600
rect 191472 146752 191524 146804
rect 113916 146208 113968 146260
rect 129832 146208 129884 146260
rect 178224 146208 178276 146260
rect 191012 146208 191064 146260
rect 113824 146140 113876 146192
rect 131672 146140 131724 146192
rect 178040 146140 178092 146192
rect 199108 146140 199160 146192
rect 112352 146072 112404 146124
rect 131120 146072 131172 146124
rect 177212 146072 177264 146124
rect 198004 146072 198056 146124
rect 111248 146004 111300 146056
rect 129924 146004 129976 146056
rect 173992 146004 174044 146056
rect 197912 146004 197964 146056
rect 122564 145936 122616 145988
rect 149152 145936 149204 145988
rect 169852 145936 169904 145988
rect 195060 145936 195112 145988
rect 120448 145868 120500 145920
rect 148600 145868 148652 145920
rect 165712 145868 165764 145920
rect 196440 145868 196492 145920
rect 116308 145800 116360 145852
rect 145380 145800 145432 145852
rect 153292 145800 153344 145852
rect 186780 145800 186832 145852
rect 116492 145732 116544 145784
rect 147036 145732 147088 145784
rect 161572 145732 161624 145784
rect 197084 145732 197136 145784
rect 113548 145664 113600 145716
rect 146760 145664 146812 145716
rect 162768 145664 162820 145716
rect 197912 145664 197964 145716
rect 115020 145596 115072 145648
rect 147956 145596 148008 145648
rect 166816 145596 166868 145648
rect 214564 145596 214616 145648
rect 3516 145528 3568 145580
rect 115388 145460 115440 145512
rect 129740 145460 129792 145512
rect 115296 145392 115348 145444
rect 130660 145392 130712 145444
rect 179420 145528 179472 145580
rect 190920 145528 190972 145580
rect 178316 145460 178368 145512
rect 189632 145460 189684 145512
rect 179512 145392 179564 145444
rect 189540 145392 189592 145444
rect 113824 145324 113876 145376
rect 127808 145324 127860 145376
rect 183744 145324 183796 145376
rect 194232 145324 194284 145376
rect 185676 144916 185728 144968
rect 115848 144848 115900 144900
rect 184020 144848 184072 144900
rect 187792 144848 187844 144900
rect 199568 144848 199620 144900
rect 181536 144780 181588 144832
rect 188068 144780 188120 144832
rect 188252 144780 188304 144832
rect 198188 144780 198240 144832
rect 173808 144712 173860 144764
rect 192116 144712 192168 144764
rect 133880 144644 133932 144696
rect 170588 144644 170640 144696
rect 192300 144644 192352 144696
rect 117780 144576 117832 144628
rect 143632 144576 143684 144628
rect 172428 144576 172480 144628
rect 193680 144576 193732 144628
rect 115572 144508 115624 144560
rect 140872 144508 140924 144560
rect 169116 144508 169168 144560
rect 193588 144508 193640 144560
rect 117780 144440 117832 144492
rect 148232 144440 148284 144492
rect 168012 144440 168064 144492
rect 194968 144440 195020 144492
rect 111248 144372 111300 144424
rect 142528 144372 142580 144424
rect 160284 144372 160336 144424
rect 189816 144372 189868 144424
rect 118792 144304 118844 144356
rect 151912 144304 151964 144356
rect 154672 144304 154724 144356
rect 188804 144304 188856 144356
rect 111432 144236 111484 144288
rect 131212 144236 131264 144288
rect 118148 144168 118200 144220
rect 130200 144168 130252 144220
rect 183284 144236 183336 144288
rect 188252 144236 188304 144288
rect 188344 144168 188396 144220
rect 182088 144100 182140 144152
rect 195060 144100 195112 144152
rect 189908 144032 189960 144084
rect 118148 143692 118200 143744
rect 145288 143692 145340 143744
rect 117228 143624 117280 143676
rect 148600 143624 148652 143676
rect 112904 143556 112956 143608
rect 145840 143556 145892 143608
rect 177120 143488 177172 143540
rect 179420 143488 179472 143540
rect 183008 143488 183060 143540
rect 187424 143488 187476 143540
rect 186044 143420 186096 143472
rect 187516 143420 187568 143472
rect 116676 143352 116728 143404
rect 128544 143352 128596 143404
rect 129832 143352 129884 143404
rect 135444 143352 135496 143404
rect 185492 143352 185544 143404
rect 191288 143352 191340 143404
rect 116768 143284 116820 143336
rect 131488 143284 131540 143336
rect 182732 143284 182784 143336
rect 197820 143284 197872 143336
rect 118056 143216 118108 143268
rect 133144 143216 133196 143268
rect 175648 143216 175700 143268
rect 192024 143216 192076 143268
rect 112260 143148 112312 143200
rect 127716 143148 127768 143200
rect 129740 143148 129792 143200
rect 137008 143148 137060 143200
rect 173532 143148 173584 143200
rect 189356 143148 189408 143200
rect 120816 143080 120868 143132
rect 139768 143080 139820 143132
rect 168288 143080 168340 143132
rect 190828 143080 190880 143132
rect 120908 143012 120960 143064
rect 141424 143012 141476 143064
rect 155960 143012 156012 143064
rect 184204 143012 184256 143064
rect 185676 143012 185728 143064
rect 196532 143012 196584 143064
rect 120724 142944 120776 142996
rect 151452 142944 151504 142996
rect 158628 142944 158680 142996
rect 187976 142944 188028 142996
rect 119804 142876 119856 142928
rect 143080 142876 143132 142928
rect 178868 142876 178920 142928
rect 214656 142876 214708 142928
rect 119528 142808 119580 142860
rect 149704 142808 149756 142860
rect 151268 142808 151320 142860
rect 209228 142808 209280 142860
rect 177948 142536 178000 142588
rect 184480 142536 184532 142588
rect 128268 142468 128320 142520
rect 580724 142468 580776 142520
rect 128544 142400 128596 142452
rect 133512 142400 133564 142452
rect 119528 142332 119580 142384
rect 182732 142400 182784 142452
rect 177856 142332 177908 142384
rect 181996 142332 182048 142384
rect 120172 142264 120224 142316
rect 186044 142264 186096 142316
rect 129924 142196 129976 142248
rect 132592 142196 132644 142248
rect 133512 142196 133564 142248
rect 580908 142196 580960 142248
rect 131120 142128 131172 142180
rect 134248 142128 134300 142180
rect 115848 142060 115900 142112
rect 150532 142128 150584 142180
rect 155776 142128 155828 142180
rect 157432 142128 157484 142180
rect 183652 142128 183704 142180
rect 191012 142128 191064 142180
rect 185952 142060 186004 142112
rect 195336 142060 195388 142112
rect 116400 141992 116452 142044
rect 127808 141992 127860 142044
rect 176476 141992 176528 142044
rect 187332 141992 187384 142044
rect 111248 141924 111300 141976
rect 123484 141924 123536 141976
rect 128912 141924 128964 141976
rect 129280 141924 129332 141976
rect 175188 141924 175240 141976
rect 187884 141924 187936 141976
rect 114008 141856 114060 141908
rect 127348 141856 127400 141908
rect 180340 141856 180392 141908
rect 193496 141856 193548 141908
rect 112628 141788 112680 141840
rect 129280 141788 129332 141840
rect 176200 141788 176252 141840
rect 182916 141788 182968 141840
rect 185584 141788 185636 141840
rect 185952 141788 186004 141840
rect 117964 141720 118016 141772
rect 134800 141720 134852 141772
rect 170220 141720 170272 141772
rect 189448 141720 189500 141772
rect 117872 141652 117924 141704
rect 119620 141584 119672 141636
rect 127808 141652 127860 141704
rect 136640 141652 136692 141704
rect 171876 141652 171928 141704
rect 190736 141652 190788 141704
rect 119344 141516 119396 141568
rect 124864 141516 124916 141568
rect 140320 141584 140372 141636
rect 163964 141584 164016 141636
rect 188528 141584 188580 141636
rect 153660 141516 153712 141568
rect 160192 141516 160244 141568
rect 186964 141516 187016 141568
rect 117228 141448 117280 141500
rect 142252 141448 142304 141500
rect 169300 141448 169352 141500
rect 196256 141448 196308 141500
rect 119436 141380 119488 141432
rect 149428 141380 149480 141432
rect 154212 141380 154264 141432
rect 187148 141380 187200 141432
rect 182916 141312 182968 141364
rect 192300 141312 192352 141364
rect 184112 141108 184164 141160
rect 189632 141108 189684 141160
rect 13084 140836 13136 140888
rect 182824 140836 182876 140888
rect 184204 140836 184256 140888
rect 187332 140836 187384 140888
rect 127348 140768 127400 140820
rect 580816 140768 580868 140820
rect 119712 140700 119764 140752
rect 126244 140700 126296 140752
rect 158720 140700 158772 140752
rect 159640 140700 159692 140752
rect 159548 140632 159600 140684
rect 193496 140700 193548 140752
rect 161848 140632 161900 140684
rect 162400 140632 162452 140684
rect 169852 140632 169904 140684
rect 170680 140632 170732 140684
rect 178040 140632 178092 140684
rect 178960 140632 179012 140684
rect 119252 140564 119304 140616
rect 126704 140564 126756 140616
rect 173900 140564 173952 140616
rect 189080 140564 189132 140616
rect 120908 140496 120960 140548
rect 129188 140496 129240 140548
rect 184848 140496 184900 140548
rect 192484 140496 192536 140548
rect 119344 140428 119396 140480
rect 127624 140428 127676 140480
rect 178776 140428 178828 140480
rect 187976 140428 188028 140480
rect 118148 140360 118200 140412
rect 126428 140360 126480 140412
rect 180064 140360 180116 140412
rect 189356 140360 189408 140412
rect 117964 140292 118016 140344
rect 129372 140292 129424 140344
rect 178684 140292 178736 140344
rect 188344 140292 188396 140344
rect 116676 140224 116728 140276
rect 129096 140224 129148 140276
rect 180248 140224 180300 140276
rect 190736 140224 190788 140276
rect 115296 140156 115348 140208
rect 146668 140156 146720 140208
rect 185860 140156 185912 140208
rect 196808 140156 196860 140208
rect 116400 140088 116452 140140
rect 148140 140088 148192 140140
rect 185952 140088 186004 140140
rect 202328 140088 202380 140140
rect 113640 140020 113692 140072
rect 126520 140020 126572 140072
rect 132500 140020 132552 140072
rect 189908 140020 189960 140072
rect 118056 139952 118108 140004
rect 125048 139952 125100 140004
rect 184572 139952 184624 140004
rect 189448 139952 189500 140004
rect 129464 139680 129516 139732
rect 187700 139680 187752 139732
rect 118700 139612 118752 139664
rect 180064 139612 180116 139664
rect 21364 139544 21416 139596
rect 185032 139544 185084 139596
rect 8944 139476 8996 139528
rect 181168 139476 181220 139528
rect 126060 139408 126112 139460
rect 327724 139408 327776 139460
rect 123024 139340 123076 139392
rect 123668 139340 123720 139392
rect 3424 138660 3476 138712
rect 120172 138660 120224 138712
rect 188620 138660 188672 138712
rect 198004 138660 198056 138712
rect 3240 137912 3292 137964
rect 118700 137912 118752 137964
rect 186872 137776 186924 137828
rect 187424 137776 187476 137828
rect 117780 136416 117832 136468
rect 118148 136416 118200 136468
rect 3056 111392 3108 111444
rect 8944 111392 8996 111444
rect 211804 88952 211856 89004
rect 212080 88952 212132 89004
rect 464344 86912 464396 86964
rect 579620 86912 579672 86964
rect 109592 81064 109644 81116
rect 122012 81064 122064 81116
rect 116308 80928 116360 80980
rect 188436 81064 188488 81116
rect 115204 80860 115256 80912
rect 111064 80792 111116 80844
rect 111156 80724 111208 80776
rect 122288 80724 122340 80776
rect 108304 80656 108356 80708
rect 131028 80588 131080 80640
rect 132224 80588 132276 80640
rect 121920 80520 121972 80572
rect 122288 80452 122340 80504
rect 105268 80248 105320 80300
rect 105636 80248 105688 80300
rect 132224 80248 132276 80300
rect 131120 80180 131172 80232
rect 129096 79976 129148 80028
rect 123484 79908 123536 79960
rect 132914 79908 132966 79960
rect 133558 79908 133610 79960
rect 133650 79908 133702 79960
rect 133742 79908 133794 79960
rect 133926 79908 133978 79960
rect 134294 79908 134346 79960
rect 134386 79908 134438 79960
rect 134570 79908 134622 79960
rect 128176 79840 128228 79892
rect 133282 79840 133334 79892
rect 131396 79772 131448 79824
rect 133604 79704 133656 79756
rect 113640 79636 113692 79688
rect 132500 79636 132552 79688
rect 133236 79636 133288 79688
rect 134018 79840 134070 79892
rect 133880 79636 133932 79688
rect 134156 79636 134208 79688
rect 134662 79840 134714 79892
rect 134524 79772 134576 79824
rect 134432 79704 134484 79756
rect 111340 79568 111392 79620
rect 126336 79568 126388 79620
rect 133972 79568 134024 79620
rect 136318 79908 136370 79960
rect 134938 79840 134990 79892
rect 135582 79840 135634 79892
rect 136042 79840 136094 79892
rect 136594 79840 136646 79892
rect 134800 79636 134852 79688
rect 135260 79636 135312 79688
rect 135444 79636 135496 79688
rect 135674 79772 135726 79824
rect 135536 79568 135588 79620
rect 135628 79568 135680 79620
rect 137330 79908 137382 79960
rect 136870 79840 136922 79892
rect 137054 79840 137106 79892
rect 137974 79908 138026 79960
rect 137514 79840 137566 79892
rect 138250 79840 138302 79892
rect 136272 79636 136324 79688
rect 136640 79636 136692 79688
rect 136732 79636 136784 79688
rect 136916 79636 136968 79688
rect 137100 79636 137152 79688
rect 137376 79636 137428 79688
rect 137468 79636 137520 79688
rect 119436 79500 119488 79552
rect 127900 79500 127952 79552
rect 131948 79500 132000 79552
rect 136456 79568 136508 79620
rect 117780 79432 117832 79484
rect 127808 79432 127860 79484
rect 134340 79432 134392 79484
rect 136732 79432 136784 79484
rect 137836 79636 137888 79688
rect 138204 79636 138256 79688
rect 138802 79908 138854 79960
rect 138434 79840 138486 79892
rect 138756 79772 138808 79824
rect 138664 79636 138716 79688
rect 139354 79908 139406 79960
rect 139446 79908 139498 79960
rect 139630 79908 139682 79960
rect 139906 79908 139958 79960
rect 139078 79840 139130 79892
rect 139170 79772 139222 79824
rect 139032 79568 139084 79620
rect 138940 79432 138992 79484
rect 139814 79840 139866 79892
rect 139676 79772 139728 79824
rect 139492 79636 139544 79688
rect 139584 79636 139636 79688
rect 140366 79840 140418 79892
rect 140550 79908 140602 79960
rect 140734 79908 140786 79960
rect 140826 79908 140878 79960
rect 141010 79908 141062 79960
rect 141654 79908 141706 79960
rect 141838 79908 141890 79960
rect 141930 79908 141982 79960
rect 142022 79908 142074 79960
rect 142206 79908 142258 79960
rect 140412 79704 140464 79756
rect 140228 79636 140280 79688
rect 139952 79500 140004 79552
rect 140412 79500 140464 79552
rect 140596 79636 140648 79688
rect 140504 79432 140556 79484
rect 141470 79840 141522 79892
rect 141608 79704 141660 79756
rect 140872 79636 140924 79688
rect 140964 79636 141016 79688
rect 141148 79636 141200 79688
rect 141700 79568 141752 79620
rect 141332 79500 141384 79552
rect 142068 79772 142120 79824
rect 141976 79500 142028 79552
rect 142160 79704 142212 79756
rect 142390 79908 142442 79960
rect 142482 79908 142534 79960
rect 142574 79908 142626 79960
rect 142850 79908 142902 79960
rect 143954 79908 144006 79960
rect 144046 79908 144098 79960
rect 142390 79772 142442 79824
rect 142252 79636 142304 79688
rect 142528 79636 142580 79688
rect 143034 79840 143086 79892
rect 143402 79840 143454 79892
rect 143218 79772 143270 79824
rect 143080 79636 143132 79688
rect 143172 79636 143224 79688
rect 142344 79500 142396 79552
rect 142620 79500 142672 79552
rect 142712 79500 142764 79552
rect 143770 79772 143822 79824
rect 143540 79568 143592 79620
rect 143816 79500 143868 79552
rect 144230 79908 144282 79960
rect 144414 79840 144466 79892
rect 144506 79840 144558 79892
rect 144690 79840 144742 79892
rect 145150 79908 145202 79960
rect 145334 79908 145386 79960
rect 144322 79772 144374 79824
rect 144276 79636 144328 79688
rect 144368 79636 144420 79688
rect 144644 79704 144696 79756
rect 144460 79568 144512 79620
rect 144874 79772 144926 79824
rect 145196 79772 145248 79824
rect 145518 79908 145570 79960
rect 145702 79840 145754 79892
rect 145104 79704 145156 79756
rect 144920 79568 144972 79620
rect 144736 79500 144788 79552
rect 145472 79432 145524 79484
rect 145840 79636 145892 79688
rect 146254 79908 146306 79960
rect 146070 79840 146122 79892
rect 146162 79840 146214 79892
rect 146438 79840 146490 79892
rect 146622 79840 146674 79892
rect 146300 79704 146352 79756
rect 146484 79636 146536 79688
rect 146116 79568 146168 79620
rect 146392 79500 146444 79552
rect 146806 79908 146858 79960
rect 146898 79840 146950 79892
rect 146852 79704 146904 79756
rect 146852 79568 146904 79620
rect 147174 79840 147226 79892
rect 147542 79840 147594 79892
rect 147358 79772 147410 79824
rect 147128 79704 147180 79756
rect 147220 79704 147272 79756
rect 147312 79636 147364 79688
rect 147726 79908 147778 79960
rect 147818 79908 147870 79960
rect 147910 79908 147962 79960
rect 148462 79908 148514 79960
rect 149014 79908 149066 79960
rect 149198 79908 149250 79960
rect 147772 79704 147824 79756
rect 148278 79840 148330 79892
rect 148002 79772 148054 79824
rect 148094 79772 148146 79824
rect 147680 79500 147732 79552
rect 147956 79636 148008 79688
rect 148738 79840 148790 79892
rect 148830 79840 148882 79892
rect 148508 79772 148560 79824
rect 148600 79636 148652 79688
rect 149290 79840 149342 79892
rect 148968 79636 149020 79688
rect 149474 79908 149526 79960
rect 149750 79908 149802 79960
rect 149934 79908 149986 79960
rect 150026 79908 150078 79960
rect 150118 79908 150170 79960
rect 150210 79908 150262 79960
rect 150670 79908 150722 79960
rect 150762 79908 150814 79960
rect 151314 79908 151366 79960
rect 151406 79908 151458 79960
rect 149382 79772 149434 79824
rect 149336 79636 149388 79688
rect 149428 79636 149480 79688
rect 149612 79636 149664 79688
rect 149888 79636 149940 79688
rect 148140 79500 148192 79552
rect 147864 79432 147916 79484
rect 148048 79432 148100 79484
rect 148600 79500 148652 79552
rect 148876 79500 148928 79552
rect 149060 79568 149112 79620
rect 151038 79840 151090 79892
rect 150716 79772 150768 79824
rect 150946 79772 150998 79824
rect 150256 79636 150308 79688
rect 150164 79568 150216 79620
rect 151130 79772 151182 79824
rect 151084 79636 151136 79688
rect 151360 79704 151412 79756
rect 150900 79568 150952 79620
rect 151176 79568 151228 79620
rect 151452 79568 151504 79620
rect 152326 79908 152378 79960
rect 152418 79908 152470 79960
rect 153154 79908 153206 79960
rect 151958 79840 152010 79892
rect 152234 79840 152286 79892
rect 150072 79500 150124 79552
rect 151728 79500 151780 79552
rect 152970 79840 153022 79892
rect 152372 79772 152424 79824
rect 152280 79704 152332 79756
rect 152924 79568 152976 79620
rect 152832 79500 152884 79552
rect 148416 79432 148468 79484
rect 148784 79432 148836 79484
rect 151820 79432 151872 79484
rect 153430 79908 153482 79960
rect 153522 79908 153574 79960
rect 153706 79908 153758 79960
rect 153890 79908 153942 79960
rect 153476 79772 153528 79824
rect 153844 79772 153896 79824
rect 153660 79704 153712 79756
rect 199476 80928 199528 80980
rect 198188 80860 198240 80912
rect 188436 80792 188488 80844
rect 215668 80792 215720 80844
rect 270500 80792 270552 80844
rect 215852 80724 215904 80776
rect 234620 80724 234672 80776
rect 178684 80588 178736 80640
rect 178776 80588 178828 80640
rect 189908 80520 189960 80572
rect 302240 80656 302292 80708
rect 154442 79908 154494 79960
rect 154810 79908 154862 79960
rect 154994 79908 155046 79960
rect 155362 79908 155414 79960
rect 155546 79908 155598 79960
rect 155914 79908 155966 79960
rect 156190 79908 156242 79960
rect 156282 79908 156334 79960
rect 154074 79840 154126 79892
rect 154120 79704 154172 79756
rect 153752 79500 153804 79552
rect 154856 79704 154908 79756
rect 155316 79772 155368 79824
rect 155730 79840 155782 79892
rect 155822 79840 155874 79892
rect 155592 79772 155644 79824
rect 155040 79636 155092 79688
rect 155408 79568 155460 79620
rect 156282 79772 156334 79824
rect 156144 79704 156196 79756
rect 155868 79568 155920 79620
rect 156926 79908 156978 79960
rect 156650 79840 156702 79892
rect 156834 79840 156886 79892
rect 156328 79500 156380 79552
rect 156788 79704 156840 79756
rect 156880 79704 156932 79756
rect 157110 79908 157162 79960
rect 157386 79908 157438 79960
rect 157754 79908 157806 79960
rect 157846 79908 157898 79960
rect 157938 79908 157990 79960
rect 158214 79908 158266 79960
rect 156972 79636 157024 79688
rect 157662 79840 157714 79892
rect 157478 79772 157530 79824
rect 157340 79704 157392 79756
rect 157156 79636 157208 79688
rect 157708 79704 157760 79756
rect 156788 79568 156840 79620
rect 157524 79568 157576 79620
rect 157616 79568 157668 79620
rect 157800 79568 157852 79620
rect 158398 79908 158450 79960
rect 158490 79908 158542 79960
rect 158260 79704 158312 79756
rect 158444 79772 158496 79824
rect 158352 79636 158404 79688
rect 157984 79568 158036 79620
rect 156696 79500 156748 79552
rect 177764 80112 177816 80164
rect 238760 80112 238812 80164
rect 179236 80044 179288 80096
rect 184480 80044 184532 80096
rect 187240 80044 187292 80096
rect 211988 80044 212040 80096
rect 212356 80044 212408 80096
rect 523132 80044 523184 80096
rect 158766 79908 158818 79960
rect 158950 79908 159002 79960
rect 159226 79908 159278 79960
rect 159962 79908 160014 79960
rect 160054 79908 160106 79960
rect 160146 79908 160198 79960
rect 160330 79908 160382 79960
rect 158858 79840 158910 79892
rect 158904 79704 158956 79756
rect 159594 79840 159646 79892
rect 159778 79840 159830 79892
rect 159502 79772 159554 79824
rect 159180 79568 159232 79620
rect 159548 79636 159600 79688
rect 159456 79568 159508 79620
rect 160054 79772 160106 79824
rect 159364 79500 159416 79552
rect 159824 79500 159876 79552
rect 160192 79636 160244 79688
rect 160008 79568 160060 79620
rect 160698 79908 160750 79960
rect 161158 79908 161210 79960
rect 161618 79908 161670 79960
rect 162170 79908 162222 79960
rect 160514 79772 160566 79824
rect 160560 79636 160612 79688
rect 160836 79500 160888 79552
rect 160928 79500 160980 79552
rect 161710 79840 161762 79892
rect 161894 79840 161946 79892
rect 162262 79772 162314 79824
rect 162722 79772 162774 79824
rect 162492 79636 162544 79688
rect 162584 79636 162636 79688
rect 162676 79636 162728 79688
rect 163090 79908 163142 79960
rect 163366 79908 163418 79960
rect 162906 79840 162958 79892
rect 163550 79908 163602 79960
rect 163320 79772 163372 79824
rect 163412 79772 163464 79824
rect 163826 79840 163878 79892
rect 164102 79840 164154 79892
rect 163596 79636 163648 79688
rect 162032 79568 162084 79620
rect 162768 79568 162820 79620
rect 163136 79568 163188 79620
rect 164286 79772 164338 79824
rect 164240 79636 164292 79688
rect 164746 79908 164798 79960
rect 164838 79908 164890 79960
rect 164930 79840 164982 79892
rect 165390 79840 165442 79892
rect 164608 79568 164660 79620
rect 161664 79500 161716 79552
rect 161756 79500 161808 79552
rect 158720 79432 158772 79484
rect 163228 79500 163280 79552
rect 163780 79500 163832 79552
rect 164056 79500 164108 79552
rect 164700 79500 164752 79552
rect 165206 79772 165258 79824
rect 165160 79636 165212 79688
rect 165252 79636 165304 79688
rect 166678 79908 166730 79960
rect 166770 79908 166822 79960
rect 165666 79840 165718 79892
rect 166034 79840 166086 79892
rect 166218 79840 166270 79892
rect 165528 79568 165580 79620
rect 165896 79568 165948 79620
rect 166586 79772 166638 79824
rect 166678 79772 166730 79824
rect 166862 79840 166914 79892
rect 167782 79908 167834 79960
rect 167874 79908 167926 79960
rect 167966 79908 168018 79960
rect 168334 79908 168386 79960
rect 168518 79908 168570 79960
rect 167414 79840 167466 79892
rect 167598 79840 167650 79892
rect 166954 79772 167006 79824
rect 167322 79772 167374 79824
rect 166724 79636 166776 79688
rect 166816 79636 166868 79688
rect 167276 79636 167328 79688
rect 167460 79636 167512 79688
rect 166172 79568 166224 79620
rect 166908 79568 166960 79620
rect 165620 79500 165672 79552
rect 167368 79500 167420 79552
rect 108212 79364 108264 79416
rect 121920 79364 121972 79416
rect 135628 79364 135680 79416
rect 144552 79364 144604 79416
rect 145288 79364 145340 79416
rect 146300 79364 146352 79416
rect 167460 79432 167512 79484
rect 162860 79364 162912 79416
rect 168196 79568 168248 79620
rect 168426 79840 168478 79892
rect 168978 79908 169030 79960
rect 169254 79908 169306 79960
rect 169530 79908 169582 79960
rect 169898 79908 169950 79960
rect 170082 79908 170134 79960
rect 170174 79908 170226 79960
rect 171002 79908 171054 79960
rect 171462 79908 171514 79960
rect 171554 79908 171606 79960
rect 172474 79908 172526 79960
rect 172566 79908 172618 79960
rect 168702 79840 168754 79892
rect 168794 79840 168846 79892
rect 168472 79636 168524 79688
rect 168564 79636 168616 79688
rect 167920 79500 167972 79552
rect 168012 79500 168064 79552
rect 168564 79500 168616 79552
rect 168840 79704 168892 79756
rect 169070 79840 169122 79892
rect 169162 79840 169214 79892
rect 169208 79704 169260 79756
rect 169484 79636 169536 79688
rect 169024 79568 169076 79620
rect 169116 79568 169168 79620
rect 169806 79772 169858 79824
rect 170036 79772 170088 79824
rect 170634 79840 170686 79892
rect 170450 79772 170502 79824
rect 170128 79704 170180 79756
rect 169852 79568 169904 79620
rect 169944 79568 169996 79620
rect 170496 79568 170548 79620
rect 171094 79840 171146 79892
rect 170956 79636 171008 79688
rect 169300 79500 169352 79552
rect 170680 79500 170732 79552
rect 170956 79500 171008 79552
rect 171370 79772 171422 79824
rect 172014 79772 172066 79824
rect 172474 79772 172526 79824
rect 171968 79636 172020 79688
rect 172612 79568 172664 79620
rect 180524 79976 180576 80028
rect 172842 79908 172894 79960
rect 173302 79840 173354 79892
rect 173854 79908 173906 79960
rect 174222 79908 174274 79960
rect 172980 79568 173032 79620
rect 173164 79568 173216 79620
rect 173394 79772 173446 79824
rect 173946 79772 173998 79824
rect 174038 79772 174090 79824
rect 174130 79772 174182 79824
rect 173348 79636 173400 79688
rect 173440 79636 173492 79688
rect 173624 79568 173676 79620
rect 174084 79568 174136 79620
rect 174498 79908 174550 79960
rect 174590 79908 174642 79960
rect 174774 79840 174826 79892
rect 174866 79840 174918 79892
rect 174544 79704 174596 79756
rect 174912 79704 174964 79756
rect 174360 79636 174412 79688
rect 175142 79908 175194 79960
rect 175234 79908 175286 79960
rect 175602 79908 175654 79960
rect 175418 79840 175470 79892
rect 175510 79840 175562 79892
rect 175188 79704 175240 79756
rect 175280 79704 175332 79756
rect 175464 79704 175516 79756
rect 175694 79772 175746 79824
rect 175970 79908 176022 79960
rect 176706 79908 176758 79960
rect 176798 79908 176850 79960
rect 177856 79908 177908 79960
rect 175878 79840 175930 79892
rect 176430 79840 176482 79892
rect 177074 79840 177126 79892
rect 178040 79840 178092 79892
rect 175924 79704 175976 79756
rect 176016 79704 176068 79756
rect 175740 79636 175792 79688
rect 177580 79772 177632 79824
rect 177672 79772 177724 79824
rect 181628 79772 181680 79824
rect 174728 79568 174780 79620
rect 175004 79568 175056 79620
rect 175556 79568 175608 79620
rect 175648 79568 175700 79620
rect 176292 79568 176344 79620
rect 177764 79568 177816 79620
rect 214656 79568 214708 79620
rect 171324 79500 171376 79552
rect 171416 79500 171468 79552
rect 171508 79500 171560 79552
rect 168656 79432 168708 79484
rect 179420 79500 179472 79552
rect 181352 79500 181404 79552
rect 202328 79500 202380 79552
rect 172244 79432 172296 79484
rect 192668 79432 192720 79484
rect 324320 79432 324372 79484
rect 108672 79296 108724 79348
rect 122656 79296 122708 79348
rect 122748 79296 122800 79348
rect 135076 79296 135128 79348
rect 136180 79296 136232 79348
rect 143632 79296 143684 79348
rect 144368 79296 144420 79348
rect 119252 79228 119304 79280
rect 135812 79228 135864 79280
rect 148324 79296 148376 79348
rect 165988 79296 166040 79348
rect 116492 79160 116544 79212
rect 152096 79228 152148 79280
rect 153016 79228 153068 79280
rect 158628 79228 158680 79280
rect 166264 79228 166316 79280
rect 167828 79364 167880 79416
rect 170588 79364 170640 79416
rect 170864 79364 170916 79416
rect 172520 79364 172572 79416
rect 179144 79364 179196 79416
rect 179236 79364 179288 79416
rect 214564 79364 214616 79416
rect 214656 79364 214708 79416
rect 358820 79364 358872 79416
rect 166540 79296 166592 79348
rect 166908 79296 166960 79348
rect 167092 79296 167144 79348
rect 180156 79296 180208 79348
rect 184388 79296 184440 79348
rect 194048 79296 194100 79348
rect 191104 79228 191156 79280
rect 136180 79160 136232 79212
rect 146116 79160 146168 79212
rect 147496 79160 147548 79212
rect 150900 79160 150952 79212
rect 156972 79160 157024 79212
rect 157892 79160 157944 79212
rect 158352 79160 158404 79212
rect 188344 79160 188396 79212
rect 113824 79092 113876 79144
rect 126244 79092 126296 79144
rect 126336 79092 126388 79144
rect 135628 79092 135680 79144
rect 135812 79092 135864 79144
rect 145748 79092 145800 79144
rect 161572 79092 161624 79144
rect 161756 79092 161808 79144
rect 164332 79092 164384 79144
rect 165068 79092 165120 79144
rect 166816 79092 166868 79144
rect 196808 79092 196860 79144
rect 116400 79024 116452 79076
rect 150072 79024 150124 79076
rect 158996 79024 159048 79076
rect 159732 79024 159784 79076
rect 160008 79024 160060 79076
rect 193864 79024 193916 79076
rect 115112 78956 115164 79008
rect 147220 78956 147272 79008
rect 147404 78956 147456 79008
rect 161848 78956 161900 79008
rect 196348 78956 196400 79008
rect 376760 79296 376812 79348
rect 113548 78888 113600 78940
rect 147128 78888 147180 78940
rect 158996 78888 159048 78940
rect 159640 78888 159692 78940
rect 166264 78888 166316 78940
rect 172244 78888 172296 78940
rect 173072 78888 173124 78940
rect 212356 78888 212408 78940
rect 115020 78820 115072 78872
rect 147772 78820 147824 78872
rect 166448 78820 166500 78872
rect 127900 78752 127952 78804
rect 130936 78752 130988 78804
rect 135536 78752 135588 78804
rect 143724 78752 143776 78804
rect 144552 78752 144604 78804
rect 159640 78752 159692 78804
rect 159916 78752 159968 78804
rect 160376 78752 160428 78804
rect 161204 78752 161256 78804
rect 127808 78684 127860 78736
rect 131028 78684 131080 78736
rect 145012 78684 145064 78736
rect 153200 78684 153252 78736
rect 153936 78684 153988 78736
rect 169944 78684 169996 78736
rect 170588 78684 170640 78736
rect 171048 78684 171100 78736
rect 171692 78684 171744 78736
rect 171968 78684 172020 78736
rect 172244 78684 172296 78736
rect 172428 78684 172480 78736
rect 173348 78684 173400 78736
rect 175372 78820 175424 78872
rect 176016 78820 176068 78872
rect 174544 78752 174596 78804
rect 178776 78684 178828 78736
rect 210424 78752 210476 78804
rect 212448 78752 212500 78804
rect 480260 78752 480312 78804
rect 201040 78684 201092 78736
rect 539692 78684 539744 78736
rect 106832 78616 106884 78668
rect 107568 78616 107620 78668
rect 135628 78616 135680 78668
rect 142436 78616 142488 78668
rect 153476 78616 153528 78668
rect 153660 78616 153712 78668
rect 157432 78616 157484 78668
rect 157616 78616 157668 78668
rect 158812 78616 158864 78668
rect 159088 78616 159140 78668
rect 160836 78616 160888 78668
rect 162216 78616 162268 78668
rect 168656 78616 168708 78668
rect 169208 78616 169260 78668
rect 169668 78616 169720 78668
rect 98920 78548 98972 78600
rect 150624 78548 150676 78600
rect 151176 78548 151228 78600
rect 176844 78616 176896 78668
rect 177580 78616 177632 78668
rect 212080 78548 212132 78600
rect 212448 78548 212500 78600
rect 103980 78480 104032 78532
rect 104348 78480 104400 78532
rect 132500 78480 132552 78532
rect 136180 78480 136232 78532
rect 152188 78480 152240 78532
rect 153476 78480 153528 78532
rect 158904 78480 158956 78532
rect 163412 78480 163464 78532
rect 164884 78480 164936 78532
rect 178684 78480 178736 78532
rect 205824 78480 205876 78532
rect 110420 78412 110472 78464
rect 110880 78412 110932 78464
rect 140964 78412 141016 78464
rect 157156 78412 157208 78464
rect 161296 78412 161348 78464
rect 181444 78412 181496 78464
rect 202144 78412 202196 78464
rect 105636 78344 105688 78396
rect 136640 78344 136692 78396
rect 168748 78344 168800 78396
rect 203156 78344 203208 78396
rect 204168 78344 204220 78396
rect 207480 78344 207532 78396
rect 207940 78344 207992 78396
rect 60740 78276 60792 78328
rect 107200 78276 107252 78328
rect 133696 78276 133748 78328
rect 75920 78208 75972 78260
rect 104440 78208 104492 78260
rect 136916 78276 136968 78328
rect 165712 78276 165764 78328
rect 166448 78276 166500 78328
rect 169024 78276 169076 78328
rect 203340 78276 203392 78328
rect 204076 78276 204128 78328
rect 205916 78276 205968 78328
rect 57980 78072 58032 78124
rect 107292 78072 107344 78124
rect 135076 78208 135128 78260
rect 149612 78208 149664 78260
rect 153016 78208 153068 78260
rect 163228 78208 163280 78260
rect 166632 78208 166684 78260
rect 168012 78208 168064 78260
rect 199016 78208 199068 78260
rect 53840 78004 53892 78056
rect 105636 78004 105688 78056
rect 46940 77936 46992 77988
rect 107108 77936 107160 77988
rect 136272 78140 136324 78192
rect 165804 78140 165856 78192
rect 171876 78140 171928 78192
rect 175464 78140 175516 78192
rect 176384 78140 176436 78192
rect 180708 78140 180760 78192
rect 207848 78140 207900 78192
rect 122104 78072 122156 78124
rect 148692 78072 148744 78124
rect 164056 78072 164108 78124
rect 178776 78072 178828 78124
rect 179144 78072 179196 78124
rect 197912 78072 197964 78124
rect 199016 78072 199068 78124
rect 199568 78072 199620 78124
rect 456800 78072 456852 78124
rect 107016 77868 107068 77920
rect 129832 78004 129884 78056
rect 134340 78004 134392 78056
rect 163596 78004 163648 78056
rect 179328 78004 179380 78056
rect 195152 78004 195204 78056
rect 204168 78004 204220 78056
rect 465172 78004 465224 78056
rect 108396 77936 108448 77988
rect 159732 77936 159784 77988
rect 159916 77936 159968 77988
rect 160192 77936 160244 77988
rect 162308 77936 162360 77988
rect 165804 77936 165856 77988
rect 166540 77936 166592 77988
rect 167552 77936 167604 77988
rect 168104 77936 168156 77988
rect 121920 77868 121972 77920
rect 122104 77868 122156 77920
rect 132316 77868 132368 77920
rect 161664 77868 161716 77920
rect 164056 77868 164108 77920
rect 165160 77868 165212 77920
rect 180524 77936 180576 77988
rect 180708 77936 180760 77988
rect 171876 77868 171928 77920
rect 181904 77868 181956 77920
rect 200948 77936 201000 77988
rect 204076 77936 204128 77988
rect 471980 77936 472032 77988
rect 166356 77800 166408 77852
rect 180708 77800 180760 77852
rect 125600 77732 125652 77784
rect 139676 77732 139728 77784
rect 167644 77732 167696 77784
rect 181628 77732 181680 77784
rect 131304 77664 131356 77716
rect 142528 77664 142580 77716
rect 163044 77664 163096 77716
rect 172520 77664 172572 77716
rect 178040 77664 178092 77716
rect 211896 77664 211948 77716
rect 104440 77596 104492 77648
rect 137836 77596 137888 77648
rect 149336 77596 149388 77648
rect 209136 77596 209188 77648
rect 107568 77528 107620 77580
rect 141240 77528 141292 77580
rect 154672 77528 154724 77580
rect 155040 77528 155092 77580
rect 167644 77528 167696 77580
rect 167828 77528 167880 77580
rect 174728 77528 174780 77580
rect 177580 77528 177632 77580
rect 118884 77460 118936 77512
rect 131672 77460 131724 77512
rect 134524 77460 134576 77512
rect 175464 77460 175516 77512
rect 176660 77460 176712 77512
rect 122012 77392 122064 77444
rect 124864 77392 124916 77444
rect 142988 77392 143040 77444
rect 143264 77392 143316 77444
rect 162124 77392 162176 77444
rect 162860 77392 162912 77444
rect 173992 77392 174044 77444
rect 175004 77392 175056 77444
rect 176292 77392 176344 77444
rect 176568 77392 176620 77444
rect 161112 77324 161164 77376
rect 153200 77256 153252 77308
rect 154028 77256 154080 77308
rect 156696 77256 156748 77308
rect 157156 77256 157208 77308
rect 161848 77256 161900 77308
rect 162676 77256 162728 77308
rect 167368 77324 167420 77376
rect 181444 77324 181496 77376
rect 166448 77256 166500 77308
rect 172888 77256 172940 77308
rect 177488 77256 177540 77308
rect 97632 77188 97684 77240
rect 137652 77188 137704 77240
rect 151728 77188 151780 77240
rect 151912 77188 151964 77240
rect 162124 77188 162176 77240
rect 213920 77188 213972 77240
rect 113732 77120 113784 77172
rect 146668 77120 146720 77172
rect 148508 77120 148560 77172
rect 154856 77120 154908 77172
rect 155224 77120 155276 77172
rect 155500 77120 155552 77172
rect 214288 77120 214340 77172
rect 214564 77120 214616 77172
rect 104164 77052 104216 77104
rect 104440 77052 104492 77104
rect 136732 77052 136784 77104
rect 158076 77052 158128 77104
rect 104072 76984 104124 77036
rect 104348 76984 104400 77036
rect 137008 76984 137060 77036
rect 138296 76984 138348 77036
rect 138572 76984 138624 77036
rect 154672 76984 154724 77036
rect 155500 76984 155552 77036
rect 160836 76984 160888 77036
rect 195336 76984 195388 77036
rect 114192 76916 114244 76968
rect 142896 76916 142948 76968
rect 115664 76848 115716 76900
rect 147036 76916 147088 76968
rect 162492 76916 162544 76968
rect 162860 76916 162912 76968
rect 168196 76916 168248 76968
rect 114100 76780 114152 76832
rect 145656 76848 145708 76900
rect 159640 76848 159692 76900
rect 175648 76916 175700 76968
rect 175832 76916 175884 76968
rect 175924 76916 175976 76968
rect 207664 76916 207716 76968
rect 144000 76780 144052 76832
rect 147036 76780 147088 76832
rect 190828 76848 190880 76900
rect 192392 76780 192444 76832
rect 253940 76848 253992 76900
rect 117964 76712 118016 76764
rect 147956 76712 148008 76764
rect 148692 76712 148744 76764
rect 153476 76712 153528 76764
rect 162124 76712 162176 76764
rect 162308 76712 162360 76764
rect 67640 76644 67692 76696
rect 97632 76644 97684 76696
rect 114008 76644 114060 76696
rect 66260 76576 66312 76628
rect 104440 76576 104492 76628
rect 114284 76576 114336 76628
rect 126244 76576 126296 76628
rect 133880 76644 133932 76696
rect 134156 76644 134208 76696
rect 137560 76644 137612 76696
rect 143540 76644 143592 76696
rect 144092 76644 144144 76696
rect 147220 76644 147272 76696
rect 180064 76644 180116 76696
rect 135352 76576 135404 76628
rect 135536 76576 135588 76628
rect 135904 76576 135956 76628
rect 136364 76576 136416 76628
rect 137008 76576 137060 76628
rect 137744 76576 137796 76628
rect 138112 76576 138164 76628
rect 138296 76576 138348 76628
rect 140044 76576 140096 76628
rect 140412 76576 140464 76628
rect 142896 76576 142948 76628
rect 146760 76576 146812 76628
rect 59360 76508 59412 76560
rect 104348 76508 104400 76560
rect 112720 76508 112772 76560
rect 143816 76508 143868 76560
rect 150072 76576 150124 76628
rect 182824 76576 182876 76628
rect 214472 76780 214524 76832
rect 289820 76780 289872 76832
rect 214564 76712 214616 76764
rect 296720 76712 296772 76764
rect 353300 76644 353352 76696
rect 195244 76576 195296 76628
rect 357532 76576 357584 76628
rect 184940 76508 184992 76560
rect 195336 76508 195388 76560
rect 367100 76508 367152 76560
rect 112444 76440 112496 76492
rect 126980 76440 127032 76492
rect 134340 76440 134392 76492
rect 134892 76440 134944 76492
rect 135720 76440 135772 76492
rect 136548 76440 136600 76492
rect 139400 76440 139452 76492
rect 141884 76440 141936 76492
rect 164332 76440 164384 76492
rect 164884 76440 164936 76492
rect 170588 76440 170640 76492
rect 199292 76440 199344 76492
rect 129648 76372 129700 76424
rect 142160 76372 142212 76424
rect 154580 76372 154632 76424
rect 155132 76372 155184 76424
rect 163964 76372 164016 76424
rect 165068 76372 165120 76424
rect 192852 76372 192904 76424
rect 134248 76304 134300 76356
rect 135168 76304 135220 76356
rect 139768 76304 139820 76356
rect 140228 76304 140280 76356
rect 141700 76304 141752 76356
rect 146024 76304 146076 76356
rect 173348 76304 173400 76356
rect 173808 76304 173860 76356
rect 174084 76304 174136 76356
rect 174636 76304 174688 76356
rect 181628 76304 181680 76356
rect 181904 76304 181956 76356
rect 201500 76304 201552 76356
rect 139676 76236 139728 76288
rect 140596 76236 140648 76288
rect 180432 76236 180484 76288
rect 180708 76236 180760 76288
rect 214380 76236 214432 76288
rect 126244 76168 126296 76220
rect 140320 76168 140372 76220
rect 140964 76168 141016 76220
rect 141424 76168 141476 76220
rect 156052 76168 156104 76220
rect 161020 76168 161072 76220
rect 162124 76168 162176 76220
rect 162952 76168 163004 76220
rect 174360 76168 174412 76220
rect 175004 76168 175056 76220
rect 126980 76100 127032 76152
rect 141976 76100 142028 76152
rect 144184 76100 144236 76152
rect 144920 76100 144972 76152
rect 172796 76100 172848 76152
rect 177212 76100 177264 76152
rect 139492 76032 139544 76084
rect 140228 76032 140280 76084
rect 162584 76032 162636 76084
rect 168012 76032 168064 76084
rect 172704 76032 172756 76084
rect 178408 76032 178460 76084
rect 173532 75964 173584 76016
rect 173716 75964 173768 76016
rect 167828 75896 167880 75948
rect 168196 75896 168248 75948
rect 108580 75828 108632 75880
rect 113180 75828 113232 75880
rect 114284 75828 114336 75880
rect 123944 75828 123996 75880
rect 148232 75828 148284 75880
rect 112812 75760 112864 75812
rect 146208 75760 146260 75812
rect 146484 75760 146536 75812
rect 102876 75692 102928 75744
rect 135168 75692 135220 75744
rect 136732 75692 136784 75744
rect 138020 75692 138072 75744
rect 171508 75828 171560 75880
rect 172060 75828 172112 75880
rect 175832 75828 175884 75880
rect 176660 75828 176712 75880
rect 185032 75828 185084 75880
rect 185124 75828 185176 75880
rect 212908 75828 212960 75880
rect 172336 75760 172388 75812
rect 206376 75760 206428 75812
rect 159548 75692 159600 75744
rect 171232 75692 171284 75744
rect 205824 75692 205876 75744
rect 116860 75624 116912 75676
rect 147312 75624 147364 75676
rect 175832 75624 175884 75676
rect 206008 75624 206060 75676
rect 114192 75556 114244 75608
rect 144276 75556 144328 75608
rect 117136 75488 117188 75540
rect 145564 75488 145616 75540
rect 157064 75488 157116 75540
rect 159088 75488 159140 75540
rect 160376 75488 160428 75540
rect 161388 75488 161440 75540
rect 171784 75556 171836 75608
rect 205916 75556 205968 75608
rect 192208 75488 192260 75540
rect 118424 75420 118476 75472
rect 135260 75420 135312 75472
rect 157340 75420 157392 75472
rect 157616 75420 157668 75472
rect 158812 75420 158864 75472
rect 159732 75420 159784 75472
rect 160192 75420 160244 75472
rect 160744 75420 160796 75472
rect 161572 75420 161624 75472
rect 162400 75420 162452 75472
rect 163044 75420 163096 75472
rect 163780 75420 163832 75472
rect 168472 75420 168524 75472
rect 169024 75420 169076 75472
rect 178408 75420 178460 75472
rect 207480 75420 207532 75472
rect 121000 75352 121052 75404
rect 136180 75352 136232 75404
rect 121184 75284 121236 75336
rect 131120 75284 131172 75336
rect 85580 75216 85632 75268
rect 103888 75216 103940 75268
rect 104440 75216 104492 75268
rect 106924 75216 106976 75268
rect 131488 75216 131540 75268
rect 141792 75352 141844 75404
rect 153016 75352 153068 75404
rect 216680 75352 216732 75404
rect 148508 75284 148560 75336
rect 157064 75284 157116 75336
rect 159088 75284 159140 75336
rect 176660 75284 176712 75336
rect 176752 75284 176804 75336
rect 177028 75284 177080 75336
rect 177212 75284 177264 75336
rect 177764 75284 177816 75336
rect 185124 75284 185176 75336
rect 205824 75284 205876 75336
rect 478144 75284 478196 75336
rect 145472 75216 145524 75268
rect 147220 75216 147272 75268
rect 147404 75216 147456 75268
rect 99196 75148 99248 75200
rect 131396 75148 131448 75200
rect 131580 75148 131632 75200
rect 133144 75148 133196 75200
rect 136180 75148 136232 75200
rect 146576 75148 146628 75200
rect 152096 75148 152148 75200
rect 152924 75148 152976 75200
rect 154028 75148 154080 75200
rect 154396 75148 154448 75200
rect 193864 75216 193916 75268
rect 205916 75216 205968 75268
rect 506480 75216 506532 75268
rect 159548 75148 159600 75200
rect 201500 75148 201552 75200
rect 207480 75148 207532 75200
rect 517520 75148 517572 75200
rect 120632 75080 120684 75132
rect 144184 75080 144236 75132
rect 151820 75080 151872 75132
rect 152464 75080 152516 75132
rect 156052 75080 156104 75132
rect 157248 75080 157300 75132
rect 157432 75080 157484 75132
rect 158168 75080 158220 75132
rect 158812 75080 158864 75132
rect 159824 75080 159876 75132
rect 160376 75080 160428 75132
rect 160560 75080 160612 75132
rect 161664 75080 161716 75132
rect 162032 75080 162084 75132
rect 162952 75080 163004 75132
rect 163320 75080 163372 75132
rect 164332 75080 164384 75132
rect 164516 75080 164568 75132
rect 165988 75080 166040 75132
rect 166172 75080 166224 75132
rect 168932 75080 168984 75132
rect 169484 75080 169536 75132
rect 175004 75080 175056 75132
rect 206284 75080 206336 75132
rect 104440 75012 104492 75064
rect 138848 75012 138900 75064
rect 146208 75012 146260 75064
rect 180800 75012 180852 75064
rect 108488 74944 108540 74996
rect 125600 74944 125652 74996
rect 165620 74944 165672 74996
rect 166172 74944 166224 74996
rect 168748 74944 168800 74996
rect 169116 74944 169168 74996
rect 176660 74944 176712 74996
rect 177304 74944 177356 74996
rect 135260 74876 135312 74928
rect 145472 74876 145524 74928
rect 164608 74876 164660 74928
rect 165252 74876 165304 74928
rect 168472 74876 168524 74928
rect 169300 74876 169352 74928
rect 165620 74808 165672 74860
rect 166908 74808 166960 74860
rect 138480 74672 138532 74724
rect 139308 74672 139360 74724
rect 131120 74536 131172 74588
rect 134800 74536 134852 74588
rect 206376 74536 206428 74588
rect 511264 74536 511316 74588
rect 104256 74468 104308 74520
rect 138664 74468 138716 74520
rect 142160 74468 142212 74520
rect 143264 74468 143316 74520
rect 152280 74468 152332 74520
rect 211528 74468 211580 74520
rect 109684 74400 109736 74452
rect 142344 74400 142396 74452
rect 142804 74400 142856 74452
rect 143448 74400 143500 74452
rect 145380 74400 145432 74452
rect 146024 74400 146076 74452
rect 171324 74400 171376 74452
rect 172244 74400 172296 74452
rect 100392 74332 100444 74384
rect 129096 74332 129148 74384
rect 170864 74332 170916 74384
rect 204720 74400 204772 74452
rect 177396 74332 177448 74384
rect 211620 74332 211672 74384
rect 116676 74264 116728 74316
rect 149704 74264 149756 74316
rect 149980 74264 150032 74316
rect 153384 74264 153436 74316
rect 188068 74264 188120 74316
rect 109868 74196 109920 74248
rect 142804 74196 142856 74248
rect 143448 74196 143500 74248
rect 143816 74196 143868 74248
rect 153660 74196 153712 74248
rect 154212 74196 154264 74248
rect 187148 74196 187200 74248
rect 111708 74128 111760 74180
rect 144092 74128 144144 74180
rect 172244 74128 172296 74180
rect 203708 74128 203760 74180
rect 108764 74060 108816 74112
rect 140504 74060 140556 74112
rect 171692 74060 171744 74112
rect 203616 74060 203668 74112
rect 119896 73992 119948 74044
rect 151728 73992 151780 74044
rect 163412 73992 163464 74044
rect 193772 73992 193824 74044
rect 89720 73924 89772 73976
rect 104256 73924 104308 73976
rect 121276 73924 121328 73976
rect 152188 73924 152240 73976
rect 161388 73924 161440 73976
rect 186964 73924 187016 73976
rect 211528 73924 211580 73976
rect 255320 73924 255372 73976
rect 22744 73856 22796 73908
rect 100392 73856 100444 73908
rect 112996 73856 113048 73908
rect 142160 73856 142212 73908
rect 146392 73856 146444 73908
rect 146944 73856 146996 73908
rect 188068 73856 188120 73908
rect 269120 73856 269172 73908
rect 8944 73788 8996 73840
rect 105820 73788 105872 73840
rect 106832 73788 106884 73840
rect 131120 73788 131172 73840
rect 131212 73788 131264 73840
rect 145104 73788 145156 73840
rect 111800 73720 111852 73772
rect 140688 73720 140740 73772
rect 175096 73788 175148 73840
rect 189080 73788 189132 73840
rect 193772 73788 193824 73840
rect 340880 73788 340932 73840
rect 152464 73720 152516 73772
rect 170772 73720 170824 73772
rect 196900 73720 196952 73772
rect 105820 73584 105872 73636
rect 132408 73584 132460 73636
rect 145012 73584 145064 73636
rect 145748 73584 145800 73636
rect 131304 73516 131356 73568
rect 131672 73516 131724 73568
rect 135628 73516 135680 73568
rect 136088 73516 136140 73568
rect 107660 73176 107712 73228
rect 108764 73176 108816 73228
rect 142344 73176 142396 73228
rect 144736 73176 144788 73228
rect 149704 73176 149756 73228
rect 97724 73108 97776 73160
rect 151268 73108 151320 73160
rect 153752 73108 153804 73160
rect 154396 73108 154448 73160
rect 155684 73108 155736 73160
rect 216772 73108 216824 73160
rect 327724 73108 327776 73160
rect 580172 73108 580224 73160
rect 122472 73040 122524 73092
rect 151084 73040 151136 73092
rect 151452 73040 151504 73092
rect 161480 73040 161532 73092
rect 162676 73040 162728 73092
rect 163228 73040 163280 73092
rect 198004 73040 198056 73092
rect 98828 72972 98880 73024
rect 133788 72972 133840 73024
rect 142344 72972 142396 73024
rect 143172 72972 143224 73024
rect 153108 72972 153160 73024
rect 186872 72972 186924 73024
rect 99012 72904 99064 72956
rect 132960 72904 133012 72956
rect 157156 72904 157208 72956
rect 191196 72904 191248 72956
rect 191748 72904 191800 72956
rect 96620 72836 96672 72888
rect 105912 72836 105964 72888
rect 140044 72836 140096 72888
rect 161480 72836 161532 72888
rect 162124 72836 162176 72888
rect 163228 72836 163280 72888
rect 163872 72836 163924 72888
rect 169852 72836 169904 72888
rect 171048 72836 171100 72888
rect 204628 72836 204680 72888
rect 216772 72836 216824 72888
rect 220084 72836 220136 72888
rect 118608 72768 118660 72820
rect 150992 72768 151044 72820
rect 162676 72768 162728 72820
rect 181352 72768 181404 72820
rect 191748 72768 191800 72820
rect 287704 72768 287756 72820
rect 114928 72700 114980 72752
rect 147680 72700 147732 72752
rect 148876 72700 148928 72752
rect 154396 72700 154448 72752
rect 187332 72700 187384 72752
rect 191656 72700 191708 72752
rect 305000 72700 305052 72752
rect 109960 72632 110012 72684
rect 142344 72632 142396 72684
rect 150992 72632 151044 72684
rect 151636 72632 151688 72684
rect 157524 72632 157576 72684
rect 192760 72632 192812 72684
rect 322940 72632 322992 72684
rect 108304 72564 108356 72616
rect 138388 72564 138440 72616
rect 156788 72564 156840 72616
rect 157064 72564 157116 72616
rect 157708 72564 157760 72616
rect 192300 72564 192352 72616
rect 323584 72564 323636 72616
rect 21456 72496 21508 72548
rect 98828 72496 98880 72548
rect 121092 72496 121144 72548
rect 149796 72496 149848 72548
rect 159180 72496 159232 72548
rect 194140 72496 194192 72548
rect 342904 72496 342956 72548
rect 9680 72428 9732 72480
rect 98736 72428 98788 72480
rect 119068 72428 119120 72480
rect 148140 72428 148192 72480
rect 161020 72428 161072 72480
rect 191656 72428 191708 72480
rect 198004 72428 198056 72480
rect 396724 72428 396776 72480
rect 110972 72360 111024 72412
rect 138112 72360 138164 72412
rect 138940 72360 138992 72412
rect 121368 72292 121420 72344
rect 129924 72292 129976 72344
rect 141516 72292 141568 72344
rect 170312 72292 170364 72344
rect 180524 72360 180576 72412
rect 207112 72360 207164 72412
rect 98736 72224 98788 72276
rect 128636 72224 128688 72276
rect 159916 72224 159968 72276
rect 194232 72224 194284 72276
rect 132868 72020 132920 72072
rect 133512 72020 133564 72072
rect 149796 71952 149848 72004
rect 150256 71952 150308 72004
rect 3516 71680 3568 71732
rect 13084 71680 13136 71732
rect 119712 71680 119764 71732
rect 128452 71680 128504 71732
rect 129648 71680 129700 71732
rect 135352 71680 135404 71732
rect 137468 71680 137520 71732
rect 142436 71680 142488 71732
rect 142988 71680 143040 71732
rect 144092 71680 144144 71732
rect 146300 71680 146352 71732
rect 149336 71680 149388 71732
rect 150164 71680 150216 71732
rect 150716 71680 150768 71732
rect 151452 71680 151504 71732
rect 157984 71680 158036 71732
rect 158536 71680 158588 71732
rect 159364 71680 159416 71732
rect 159548 71680 159600 71732
rect 164240 71680 164292 71732
rect 165068 71680 165120 71732
rect 165528 71680 165580 71732
rect 206192 71680 206244 71732
rect 105728 71612 105780 71664
rect 139768 71612 139820 71664
rect 140780 71612 140832 71664
rect 143356 71612 143408 71664
rect 157340 71612 157392 71664
rect 158260 71612 158312 71664
rect 118056 71544 118108 71596
rect 149336 71544 149388 71596
rect 150440 71544 150492 71596
rect 151544 71544 151596 71596
rect 157616 71544 157668 71596
rect 158444 71544 158496 71596
rect 164240 71544 164292 71596
rect 164884 71544 164936 71596
rect 166816 71612 166868 71664
rect 207388 71612 207440 71664
rect 193956 71544 194008 71596
rect 104256 71476 104308 71528
rect 104532 71476 104584 71528
rect 135352 71476 135404 71528
rect 149152 71476 149204 71528
rect 150164 71476 150216 71528
rect 157340 71476 157392 71528
rect 157892 71476 157944 71528
rect 158352 71476 158404 71528
rect 192576 71476 192628 71528
rect 84844 71068 84896 71120
rect 106004 71408 106056 71460
rect 138204 71408 138256 71460
rect 162492 71408 162544 71460
rect 197084 71408 197136 71460
rect 120908 71340 120960 71392
rect 152004 71340 152056 71392
rect 158444 71340 158496 71392
rect 192484 71340 192536 71392
rect 117596 71272 117648 71324
rect 149428 71272 149480 71324
rect 165068 71272 165120 71324
rect 199200 71272 199252 71324
rect 112536 71204 112588 71256
rect 142436 71204 142488 71256
rect 158260 71204 158312 71256
rect 191012 71204 191064 71256
rect 135260 71136 135312 71188
rect 135720 71136 135772 71188
rect 146576 71136 146628 71188
rect 181444 71136 181496 71188
rect 181812 71136 181864 71188
rect 203248 71136 203300 71188
rect 114376 71068 114428 71120
rect 128360 71068 128412 71120
rect 141240 71068 141292 71120
rect 147128 71068 147180 71120
rect 184296 71068 184348 71120
rect 71780 71000 71832 71052
rect 104256 71000 104308 71052
rect 110788 71000 110840 71052
rect 140780 71000 140832 71052
rect 148876 71000 148928 71052
rect 200856 71000 200908 71052
rect 121552 70932 121604 70984
rect 151452 70932 151504 70984
rect 156328 70932 156380 70984
rect 157248 70932 157300 70984
rect 187700 70932 187752 70984
rect 117228 70864 117280 70916
rect 140964 70864 141016 70916
rect 152004 70864 152056 70916
rect 152924 70864 152976 70916
rect 158536 70864 158588 70916
rect 188252 70864 188304 70916
rect 114836 70796 114888 70848
rect 149152 70796 149204 70848
rect 121644 70728 121696 70780
rect 150440 70796 150492 70848
rect 158628 70796 158680 70848
rect 187056 70796 187108 70848
rect 149428 70728 149480 70780
rect 150072 70728 150124 70780
rect 167368 70728 167420 70780
rect 167736 70728 167788 70780
rect 171232 70728 171284 70780
rect 171968 70728 172020 70780
rect 175004 70728 175056 70780
rect 175188 70728 175240 70780
rect 103520 70388 103572 70440
rect 105728 70388 105780 70440
rect 100116 70320 100168 70372
rect 134340 70320 134392 70372
rect 165344 70320 165396 70372
rect 205732 70320 205784 70372
rect 209136 70320 209188 70372
rect 210424 70320 210476 70372
rect 100760 70252 100812 70304
rect 101312 70252 101364 70304
rect 135996 70252 136048 70304
rect 162400 70252 162452 70304
rect 196624 70252 196676 70304
rect 104624 70184 104676 70236
rect 138756 70184 138808 70236
rect 163872 70184 163924 70236
rect 198280 70184 198332 70236
rect 97908 70116 97960 70168
rect 115940 70116 115992 70168
rect 117228 70116 117280 70168
rect 117688 70116 117740 70168
rect 151360 70116 151412 70168
rect 162584 70116 162636 70168
rect 197176 70116 197228 70168
rect 118792 70048 118844 70100
rect 151820 70048 151872 70100
rect 171232 70048 171284 70100
rect 172152 70048 172204 70100
rect 205640 70048 205692 70100
rect 107384 69980 107436 70032
rect 140136 69980 140188 70032
rect 161756 69980 161808 70032
rect 162400 69980 162452 70032
rect 164700 69980 164752 70032
rect 165344 69980 165396 70032
rect 169024 69980 169076 70032
rect 169484 69980 169536 70032
rect 203432 69980 203484 70032
rect 102140 69912 102192 69964
rect 102968 69912 103020 69964
rect 134892 69912 134944 69964
rect 161940 69912 161992 69964
rect 162584 69912 162636 69964
rect 163136 69912 163188 69964
rect 163872 69912 163924 69964
rect 164792 69912 164844 69964
rect 165528 69912 165580 69964
rect 199752 69912 199804 69964
rect 112168 69844 112220 69896
rect 143540 69844 143592 69896
rect 144460 69844 144512 69896
rect 159088 69844 159140 69896
rect 159916 69844 159968 69896
rect 191380 69844 191432 69896
rect 85672 69776 85724 69828
rect 104624 69776 104676 69828
rect 112076 69776 112128 69828
rect 142528 69776 142580 69828
rect 143080 69776 143132 69828
rect 154488 69776 154540 69828
rect 184480 69776 184532 69828
rect 45560 69708 45612 69760
rect 100760 69708 100812 69760
rect 102784 69708 102836 69760
rect 107384 69708 107436 69760
rect 113088 69708 113140 69760
rect 139400 69708 139452 69760
rect 158996 69708 159048 69760
rect 159640 69708 159692 69760
rect 189632 69708 189684 69760
rect 201684 69708 201736 69760
rect 201868 69708 201920 69760
rect 35164 69640 35216 69692
rect 102140 69640 102192 69692
rect 147588 69640 147640 69692
rect 183560 69640 183612 69692
rect 153568 69572 153620 69624
rect 154488 69572 154540 69624
rect 160468 69572 160520 69624
rect 161112 69572 161164 69624
rect 188160 69572 188212 69624
rect 162308 69504 162360 69556
rect 185400 69504 185452 69556
rect 180156 69436 180208 69488
rect 197268 69436 197320 69488
rect 210516 69640 210568 69692
rect 151820 69028 151872 69080
rect 152556 69028 152608 69080
rect 185400 69028 185452 69080
rect 354680 69028 354732 69080
rect 107568 68960 107620 69012
rect 114560 68960 114612 69012
rect 110328 68892 110380 68944
rect 110144 68824 110196 68876
rect 132040 68892 132092 68944
rect 141516 68960 141568 69012
rect 142160 68960 142212 69012
rect 158904 68960 158956 69012
rect 159732 68960 159784 69012
rect 207296 68960 207348 69012
rect 144000 68892 144052 68944
rect 144460 68892 144512 68944
rect 166080 68892 166132 68944
rect 166816 68892 166868 68944
rect 177580 68892 177632 68944
rect 212816 68892 212868 68944
rect 213828 68892 213880 68944
rect 121736 68824 121788 68876
rect 132224 68824 132276 68876
rect 132408 68824 132460 68876
rect 156052 68824 156104 68876
rect 165988 68824 166040 68876
rect 166908 68824 166960 68876
rect 167000 68824 167052 68876
rect 167920 68824 167972 68876
rect 202052 68824 202104 68876
rect 48320 68416 48372 68468
rect 101588 68756 101640 68808
rect 131948 68756 132000 68808
rect 132040 68756 132092 68808
rect 144276 68756 144328 68808
rect 144552 68756 144604 68808
rect 167092 68756 167144 68808
rect 168012 68756 168064 68808
rect 201960 68756 202012 68808
rect 108856 68688 108908 68740
rect 142712 68688 142764 68740
rect 166908 68688 166960 68740
rect 200764 68688 200816 68740
rect 26240 68348 26292 68400
rect 101680 68348 101732 68400
rect 134432 68620 134484 68672
rect 142160 68620 142212 68672
rect 142344 68620 142396 68672
rect 153292 68620 153344 68672
rect 154304 68620 154356 68672
rect 166816 68620 166868 68672
rect 200672 68620 200724 68672
rect 106924 68552 106976 68604
rect 109776 68552 109828 68604
rect 139676 68552 139728 68604
rect 169852 68552 169904 68604
rect 170956 68552 171008 68604
rect 204444 68552 204496 68604
rect 18604 68280 18656 68332
rect 101772 68280 101824 68332
rect 133604 68484 133656 68536
rect 142436 68484 142488 68536
rect 186320 68484 186372 68536
rect 186688 68484 186740 68536
rect 252560 68484 252612 68536
rect 131948 68416 132000 68468
rect 135628 68416 135680 68468
rect 166172 68416 166224 68468
rect 200580 68416 200632 68468
rect 427820 68416 427872 68468
rect 164608 68348 164660 68400
rect 195060 68348 195112 68400
rect 423680 68348 423732 68400
rect 147312 68280 147364 68332
rect 189724 68280 189776 68332
rect 213828 68280 213880 68332
rect 536840 68280 536892 68332
rect 142436 68212 142488 68264
rect 168840 68212 168892 68264
rect 169576 68212 169628 68264
rect 203800 68212 203852 68264
rect 168932 68144 168984 68196
rect 169668 68144 169720 68196
rect 199384 68144 199436 68196
rect 152740 68076 152792 68128
rect 186320 68076 186372 68128
rect 154304 68008 154356 68060
rect 186780 68008 186832 68060
rect 156052 67600 156104 67652
rect 156788 67600 156840 67652
rect 114468 67532 114520 67584
rect 147956 67532 148008 67584
rect 161296 67532 161348 67584
rect 189080 67532 189132 67584
rect 189448 67532 189500 67584
rect 108948 67464 109000 67516
rect 142620 67464 142672 67516
rect 160284 67464 160336 67516
rect 160928 67464 160980 67516
rect 195520 67464 195572 67516
rect 115388 67396 115440 67448
rect 148508 67396 148560 67448
rect 148784 67396 148836 67448
rect 174360 67396 174412 67448
rect 175004 67396 175056 67448
rect 176292 67396 176344 67448
rect 208860 67396 208912 67448
rect 116216 67328 116268 67380
rect 149060 67328 149112 67380
rect 149888 67328 149940 67380
rect 155040 67328 155092 67380
rect 155868 67328 155920 67380
rect 189172 67328 189224 67380
rect 103244 67260 103296 67312
rect 40040 66920 40092 66972
rect 135812 67260 135864 67312
rect 174268 67260 174320 67312
rect 174912 67260 174964 67312
rect 175004 67260 175056 67312
rect 208676 67260 208728 67312
rect 109040 67192 109092 67244
rect 138572 67192 138624 67244
rect 164056 67192 164108 67244
rect 196992 67192 197044 67244
rect 174176 67124 174228 67176
rect 174820 67124 174872 67176
rect 175556 67124 175608 67176
rect 201684 67124 201736 67176
rect 202788 67124 202840 67176
rect 172888 67056 172940 67108
rect 199200 67056 199252 67108
rect 169760 66988 169812 67040
rect 193404 66988 193456 67040
rect 194508 66988 194560 67040
rect 168104 66920 168156 66972
rect 184388 66920 184440 66972
rect 97448 66852 97500 66904
rect 113180 66852 113232 66904
rect 141056 66852 141108 66904
rect 174912 66852 174964 66904
rect 176292 66852 176344 66904
rect 189080 66852 189132 66904
rect 317420 66852 317472 66904
rect 174820 66784 174872 66836
rect 208952 66784 209004 66836
rect 194508 66376 194560 66428
rect 494060 66376 494112 66428
rect 199200 66308 199252 66360
rect 529940 66308 529992 66360
rect 202788 66240 202840 66292
rect 554044 66240 554096 66292
rect 121828 66172 121880 66224
rect 155960 66172 156012 66224
rect 160192 66172 160244 66224
rect 161296 66172 161348 66224
rect 208768 66172 208820 66224
rect 101404 66104 101456 66156
rect 135536 66104 135588 66156
rect 138112 66104 138164 66156
rect 138664 66104 138716 66156
rect 163044 66104 163096 66156
rect 163780 66104 163832 66156
rect 204352 66104 204404 66156
rect 108304 66036 108356 66088
rect 140228 66036 140280 66088
rect 154856 66036 154908 66088
rect 189080 66036 189132 66088
rect 204168 66036 204220 66088
rect 211436 66036 211488 66088
rect 102140 65968 102192 66020
rect 103336 65968 103388 66020
rect 134248 65968 134300 66020
rect 164516 65968 164568 66020
rect 198924 65968 198976 66020
rect 108120 65900 108172 65952
rect 138112 65900 138164 65952
rect 158812 65900 158864 65952
rect 191932 65900 191984 65952
rect 193036 65900 193088 65952
rect 104624 65832 104676 65884
rect 133052 65832 133104 65884
rect 172796 65832 172848 65884
rect 196164 65832 196216 65884
rect 111248 65764 111300 65816
rect 139952 65764 140004 65816
rect 155960 65764 156012 65816
rect 156788 65764 156840 65816
rect 148140 65696 148192 65748
rect 207664 65696 207716 65748
rect 189080 65628 189132 65680
rect 295340 65628 295392 65680
rect 193036 65560 193088 65612
rect 351920 65560 351972 65612
rect 35992 65492 36044 65544
rect 102140 65492 102192 65544
rect 109500 65492 109552 65544
rect 117320 65492 117372 65544
rect 141148 65492 141200 65544
rect 198924 65492 198976 65544
rect 414664 65492 414716 65544
rect 196164 64880 196216 64932
rect 525800 64880 525852 64932
rect 103060 64812 103112 64864
rect 137284 64812 137336 64864
rect 164424 64812 164476 64864
rect 199660 64812 199712 64864
rect 104716 64744 104768 64796
rect 136824 64744 136876 64796
rect 156144 64744 156196 64796
rect 190644 64744 190696 64796
rect 191748 64744 191800 64796
rect 111248 64676 111300 64728
rect 139860 64676 139912 64728
rect 165896 64676 165948 64728
rect 200120 64676 200172 64728
rect 168748 64608 168800 64660
rect 202972 64608 203024 64660
rect 174084 64540 174136 64592
rect 198924 64540 198976 64592
rect 161572 64472 161624 64524
rect 162308 64472 162360 64524
rect 185676 64472 185728 64524
rect 62120 64200 62172 64252
rect 103060 64200 103112 64252
rect 191748 64200 191800 64252
rect 306380 64200 306432 64252
rect 57244 64132 57296 64184
rect 104716 64132 104768 64184
rect 106740 64132 106792 64184
rect 120080 64132 120132 64184
rect 141240 64132 141292 64184
rect 146392 64132 146444 64184
rect 185584 64132 185636 64184
rect 202972 64132 203024 64184
rect 472624 64132 472676 64184
rect 164424 63860 164476 63912
rect 165252 63860 165304 63912
rect 165896 63860 165948 63912
rect 166632 63860 166684 63912
rect 144460 63520 144512 63572
rect 147220 63520 147272 63572
rect 198924 63520 198976 63572
rect 543740 63520 543792 63572
rect 106096 63452 106148 63504
rect 137008 63452 137060 63504
rect 164332 63452 164384 63504
rect 198740 63452 198792 63504
rect 115112 63384 115164 63436
rect 138480 63384 138532 63436
rect 154764 63384 154816 63436
rect 189080 63384 189132 63436
rect 166448 63316 166500 63368
rect 187240 63316 187292 63368
rect 144368 63180 144420 63232
rect 148324 63180 148376 63232
rect 150808 62908 150860 62960
rect 245660 62908 245712 62960
rect 189080 62840 189132 62892
rect 190000 62840 190052 62892
rect 292580 62840 292632 62892
rect 69020 62772 69072 62824
rect 106096 62772 106148 62824
rect 198740 62772 198792 62824
rect 412640 62772 412692 62824
rect 138664 62568 138716 62620
rect 142436 62568 142488 62620
rect 187240 62092 187292 62144
rect 368480 62092 368532 62144
rect 102140 62024 102192 62076
rect 103152 62024 103204 62076
rect 135444 62024 135496 62076
rect 162952 62024 163004 62076
rect 197728 62024 197780 62076
rect 198188 62024 198240 62076
rect 153200 61956 153252 62008
rect 187884 61956 187936 62008
rect 157064 61888 157116 61940
rect 190552 61888 190604 61940
rect 191748 61888 191800 61940
rect 172704 61820 172756 61872
rect 202144 61820 202196 61872
rect 202788 61820 202840 61872
rect 187884 61480 187936 61532
rect 188712 61480 188764 61532
rect 277400 61480 277452 61532
rect 191748 61412 191800 61464
rect 313280 61412 313332 61464
rect 43444 61344 43496 61396
rect 102140 61344 102192 61396
rect 147772 61344 147824 61396
rect 197452 61344 197504 61396
rect 198188 61344 198240 61396
rect 398840 61344 398892 61396
rect 202788 60732 202840 60784
rect 527824 60732 527876 60784
rect 102140 60664 102192 60716
rect 103428 60664 103480 60716
rect 135904 60664 135956 60716
rect 158720 60664 158772 60716
rect 193496 60664 193548 60716
rect 194508 60664 194560 60716
rect 162860 60596 162912 60648
rect 197728 60596 197780 60648
rect 154672 60528 154724 60580
rect 189080 60528 189132 60580
rect 166540 60460 166592 60512
rect 197820 60460 197872 60512
rect 147956 60324 148008 60376
rect 198740 60324 198792 60376
rect 149612 60256 149664 60308
rect 231860 60256 231912 60308
rect 145288 60188 145340 60240
rect 148416 60188 148468 60240
rect 189080 60188 189132 60240
rect 190092 60188 190144 60240
rect 299480 60188 299532 60240
rect 194508 60120 194560 60172
rect 340972 60120 341024 60172
rect 197728 60052 197780 60104
rect 198372 60052 198424 60104
rect 394700 60052 394752 60104
rect 52552 59984 52604 60036
rect 102140 59984 102192 60036
rect 197820 59984 197872 60036
rect 198464 59984 198516 60036
rect 396080 59984 396132 60036
rect 157524 59304 157576 59356
rect 191932 59304 191984 59356
rect 193036 59304 193088 59356
rect 139400 58760 139452 58812
rect 142160 58760 142212 58812
rect 151728 58692 151780 58744
rect 249800 58692 249852 58744
rect 193036 58624 193088 58676
rect 327080 58624 327132 58676
rect 168656 57876 168708 57928
rect 203248 57876 203300 57928
rect 204076 57876 204128 57928
rect 173992 57808 174044 57860
rect 204996 57808 205048 57860
rect 176936 57740 176988 57792
rect 198004 57740 198056 57792
rect 152372 57264 152424 57316
rect 263600 57264 263652 57316
rect 145656 57196 145708 57248
rect 169760 57196 169812 57248
rect 204996 57196 205048 57248
rect 545120 57196 545172 57248
rect 204076 56652 204128 56704
rect 473452 56652 473504 56704
rect 198004 56584 198056 56636
rect 567844 56584 567896 56636
rect 104440 56516 104492 56568
rect 137100 56516 137152 56568
rect 157432 56516 157484 56568
rect 187976 56516 188028 56568
rect 149428 55904 149480 55956
rect 229100 55904 229152 55956
rect 187976 55836 188028 55888
rect 331220 55836 331272 55888
rect 136640 55224 136692 55276
rect 142344 55224 142396 55276
rect 156972 55156 157024 55208
rect 189356 55156 189408 55208
rect 150440 54544 150492 54596
rect 239404 54544 239456 54596
rect 189356 54476 189408 54528
rect 315304 54476 315356 54528
rect 163504 53728 163556 53780
rect 194324 53728 194376 53780
rect 148692 53184 148744 53236
rect 201592 53184 201644 53236
rect 153016 53116 153068 53168
rect 267740 53116 267792 53168
rect 194324 53048 194376 53100
rect 389180 53048 389232 53100
rect 99472 52368 99524 52420
rect 100484 52368 100536 52420
rect 133144 52368 133196 52420
rect 168380 52368 168432 52420
rect 202880 52368 202932 52420
rect 204076 52368 204128 52420
rect 150256 51756 150308 51808
rect 224960 51756 225012 51808
rect 17960 51688 18012 51740
rect 99472 51688 99524 51740
rect 204076 51688 204128 51740
rect 464344 51688 464396 51740
rect 176844 51008 176896 51060
rect 207112 51008 207164 51060
rect 207756 51008 207808 51060
rect 207112 50328 207164 50380
rect 569960 50328 570012 50380
rect 172612 49648 172664 49700
rect 204904 49648 204956 49700
rect 148600 49104 148652 49156
rect 204260 49104 204312 49156
rect 167644 49036 167696 49088
rect 455420 49036 455472 49088
rect 145196 48968 145248 49020
rect 168656 48968 168708 49020
rect 204904 48968 204956 49020
rect 516140 48968 516192 49020
rect 168564 48220 168616 48272
rect 203064 48220 203116 48272
rect 204076 48220 204128 48272
rect 150164 47608 150216 47660
rect 215300 47608 215352 47660
rect 149520 47540 149572 47592
rect 218152 47540 218204 47592
rect 204076 46928 204128 46980
rect 466460 46928 466512 46980
rect 176752 46860 176804 46912
rect 207112 46860 207164 46912
rect 150072 46248 150124 46300
rect 219440 46248 219492 46300
rect 155316 46180 155368 46232
rect 285680 46180 285732 46232
rect 135352 45568 135404 45620
rect 142252 45568 142304 45620
rect 207848 45568 207900 45620
rect 571984 45568 572036 45620
rect 151636 44888 151688 44940
rect 242900 44888 242952 44940
rect 161480 44820 161532 44872
rect 390560 44820 390612 44872
rect 176660 44072 176712 44124
rect 207020 44072 207072 44124
rect 167460 43392 167512 43444
rect 458180 43392 458232 43444
rect 207020 42780 207072 42832
rect 576860 42780 576912 42832
rect 158260 42236 158312 42288
rect 324412 42236 324464 42288
rect 164240 42168 164292 42220
rect 426440 42168 426492 42220
rect 167736 42100 167788 42152
rect 452660 42100 452712 42152
rect 70400 42032 70452 42084
rect 136732 42032 136784 42084
rect 170496 42032 170548 42084
rect 495440 42032 495492 42084
rect 154580 41352 154632 41404
rect 187792 41352 187844 41404
rect 151544 41012 151596 41064
rect 233240 41012 233292 41064
rect 187792 40944 187844 40996
rect 188804 40944 188856 40996
rect 292672 40944 292724 40996
rect 157340 40876 157392 40928
rect 333980 40876 334032 40928
rect 165804 40808 165856 40860
rect 444380 40808 444432 40860
rect 171968 40740 172020 40792
rect 498292 40740 498344 40792
rect 74540 40672 74592 40724
rect 138296 40672 138348 40724
rect 174820 40672 174872 40724
rect 535460 40672 535512 40724
rect 153108 39516 153160 39568
rect 266360 39516 266412 39568
rect 165068 39448 165120 39500
rect 409880 39448 409932 39500
rect 167828 39380 167880 39432
rect 462320 39380 462372 39432
rect 77392 39312 77444 39364
rect 138112 39312 138164 39364
rect 176292 39312 176344 39364
rect 562324 39312 562376 39364
rect 156880 38088 156932 38140
rect 318800 38088 318852 38140
rect 169484 38020 169536 38072
rect 463700 38020 463752 38072
rect 168472 37952 168524 38004
rect 476120 37952 476172 38004
rect 13820 37884 13872 37936
rect 132868 37884 132920 37936
rect 172520 37884 172572 37936
rect 525064 37884 525116 37936
rect 148508 36796 148560 36848
rect 205640 36796 205692 36848
rect 153660 36728 153712 36780
rect 267832 36728 267884 36780
rect 160928 36660 160980 36712
rect 356704 36660 356756 36712
rect 170680 36592 170732 36644
rect 481640 36592 481692 36644
rect 23480 36524 23532 36576
rect 134064 36524 134116 36576
rect 172060 36524 172112 36576
rect 503720 36524 503772 36576
rect 156788 35368 156840 35420
rect 303620 35368 303672 35420
rect 170588 35300 170640 35352
rect 488540 35300 488592 35352
rect 174912 35232 174964 35284
rect 538864 35232 538916 35284
rect 31760 35164 31812 35216
rect 134156 35164 134208 35216
rect 176384 35164 176436 35216
rect 552020 35164 552072 35216
rect 151452 34076 151504 34128
rect 236000 34076 236052 34128
rect 152924 34008 152976 34060
rect 251180 34008 251232 34060
rect 159548 33940 159600 33992
rect 339500 33940 339552 33992
rect 166632 33872 166684 33924
rect 431960 33872 432012 33924
rect 175648 33804 175700 33856
rect 558920 33804 558972 33856
rect 38660 33736 38712 33788
rect 135536 33736 135588 33788
rect 177672 33736 177724 33788
rect 578240 33736 578292 33788
rect 148968 32648 149020 32700
rect 208400 32648 208452 32700
rect 151360 32580 151412 32632
rect 242992 32580 243044 32632
rect 158352 32512 158404 32564
rect 332692 32512 332744 32564
rect 161020 32444 161072 32496
rect 372620 32444 372672 32496
rect 165712 32376 165764 32428
rect 438860 32376 438912 32428
rect 149980 31288 150032 31340
rect 222200 31288 222252 31340
rect 152280 31220 152332 31272
rect 264980 31220 265032 31272
rect 159640 31152 159692 31204
rect 346400 31152 346452 31204
rect 162216 31084 162268 31136
rect 390652 31084 390704 31136
rect 42800 31016 42852 31068
rect 136548 31016 136600 31068
rect 145564 31016 145616 31068
rect 164884 31016 164936 31068
rect 169576 31016 169628 31068
rect 470600 31016 470652 31068
rect 144276 30268 144328 30320
rect 145104 30268 145156 30320
rect 155224 29860 155276 29912
rect 299572 29860 299624 29912
rect 163964 29792 164016 29844
rect 398932 29792 398984 29844
rect 170772 29724 170824 29776
rect 491300 29724 491352 29776
rect 145932 29656 145984 29708
rect 175924 29656 175976 29708
rect 176476 29656 176528 29708
rect 553400 29656 553452 29708
rect 175464 29588 175516 29640
rect 567936 29588 567988 29640
rect 158444 28432 158496 28484
rect 321560 28432 321612 28484
rect 165160 28364 165212 28416
rect 420920 28364 420972 28416
rect 172244 28296 172296 28348
rect 502340 28296 502392 28348
rect 177764 28228 177816 28280
rect 518900 28228 518952 28280
rect 154212 27140 154264 27192
rect 271880 27140 271932 27192
rect 161112 27072 161164 27124
rect 360200 27072 360252 27124
rect 162308 27004 162360 27056
rect 386420 27004 386472 27056
rect 170864 26936 170916 26988
rect 492680 26936 492732 26988
rect 46204 26868 46256 26920
rect 135720 26868 135772 26920
rect 172336 26868 172388 26920
rect 506572 26868 506624 26920
rect 154028 25712 154080 25764
rect 278780 25712 278832 25764
rect 162400 25644 162452 25696
rect 374092 25644 374144 25696
rect 172428 25576 172480 25628
rect 509240 25576 509292 25628
rect 145012 25508 145064 25560
rect 171784 25508 171836 25560
rect 172152 25508 172204 25560
rect 510620 25508 510672 25560
rect 163872 24216 163924 24268
rect 391940 24216 391992 24268
rect 171140 24148 171192 24200
rect 513380 24148 513432 24200
rect 173624 24080 173676 24132
rect 531412 24080 531464 24132
rect 153844 22992 153896 23044
rect 282920 22992 282972 23044
rect 162492 22924 162544 22976
rect 382280 22924 382332 22976
rect 163780 22856 163832 22908
rect 404360 22856 404412 22908
rect 173716 22788 173768 22840
rect 520280 22788 520332 22840
rect 173808 22720 173860 22772
rect 524420 22720 524472 22772
rect 159732 21428 159784 21480
rect 350540 21428 350592 21480
rect 165344 21360 165396 21412
rect 418160 21360 418212 21412
rect 155868 20068 155920 20120
rect 287060 20068 287112 20120
rect 155776 20000 155828 20052
rect 291200 20000 291252 20052
rect 143632 19932 143684 19984
rect 154580 19932 154632 19984
rect 161204 19932 161256 19984
rect 361580 19932 361632 19984
rect 152832 18844 152884 18896
rect 251272 18844 251324 18896
rect 159824 18776 159876 18828
rect 345020 18776 345072 18828
rect 165252 18708 165304 18760
rect 411260 18708 411312 18760
rect 177856 18640 177908 18692
rect 571340 18640 571392 18692
rect 177948 18572 178000 18624
rect 574100 18572 574152 18624
rect 152648 17416 152700 17468
rect 259552 17416 259604 17468
rect 167920 17348 167972 17400
rect 445760 17348 445812 17400
rect 168012 17280 168064 17332
rect 448612 17280 448664 17332
rect 146024 17212 146076 17264
rect 167000 17212 167052 17264
rect 169668 17212 169720 17264
rect 477500 17212 477552 17264
rect 154396 16124 154448 16176
rect 284392 16124 284444 16176
rect 160100 16056 160152 16108
rect 364616 16056 364668 16108
rect 165436 15988 165488 16040
rect 417424 15988 417476 16040
rect 166724 15920 166776 15972
rect 440332 15920 440384 15972
rect 175004 15852 175056 15904
rect 546500 15852 546552 15904
rect 154304 14696 154356 14748
rect 276020 14696 276072 14748
rect 157248 14628 157300 14680
rect 314660 14628 314712 14680
rect 168104 14560 168156 14612
rect 382372 14560 382424 14612
rect 162676 14492 162728 14544
rect 385960 14492 386012 14544
rect 170956 14424 171008 14476
rect 486424 14424 486476 14476
rect 152556 13336 152608 13388
rect 258264 13336 258316 13388
rect 156696 13268 156748 13320
rect 307944 13268 307996 13320
rect 164056 13200 164108 13252
rect 376024 13200 376076 13252
rect 162584 13132 162636 13184
rect 378416 13132 378468 13184
rect 171048 13064 171100 13116
rect 482192 13064 482244 13116
rect 149796 11976 149848 12028
rect 226340 11976 226392 12028
rect 158536 11908 158588 11960
rect 328736 11908 328788 11960
rect 164148 11840 164200 11892
rect 407212 11840 407264 11892
rect 168196 11772 168248 11824
rect 454040 11772 454092 11824
rect 175372 11704 175424 11756
rect 560392 11704 560444 11756
rect 184940 11636 184992 11688
rect 186136 11636 186188 11688
rect 201500 11636 201552 11688
rect 202696 11636 202748 11688
rect 234620 11636 234672 11688
rect 235816 11636 235868 11688
rect 151176 10548 151228 10600
rect 234620 10548 234672 10600
rect 158628 10480 158680 10532
rect 336280 10480 336332 10532
rect 161296 10412 161348 10464
rect 365812 10412 365864 10464
rect 166816 10344 166868 10396
rect 432052 10344 432104 10396
rect 30104 10276 30156 10328
rect 133972 10276 134024 10328
rect 175096 10276 175148 10328
rect 548616 10276 548668 10328
rect 149888 9188 149940 9240
rect 227536 9188 227588 9240
rect 156604 9120 156656 9172
rect 316224 9120 316276 9172
rect 165528 9052 165580 9104
rect 414296 9052 414348 9104
rect 184204 8984 184256 9036
rect 562048 8984 562100 9036
rect 6460 8916 6512 8968
rect 132592 8916 132644 8968
rect 175280 8916 175332 8968
rect 556160 8916 556212 8968
rect 151268 7828 151320 7880
rect 241704 7828 241756 7880
rect 160008 7760 160060 7812
rect 343364 7760 343416 7812
rect 162768 7692 162820 7744
rect 379980 7692 380032 7744
rect 166908 7624 166960 7676
rect 435548 7624 435600 7676
rect 103336 7556 103388 7608
rect 139584 7556 139636 7608
rect 175188 7556 175240 7608
rect 538404 7556 538456 7608
rect 3424 6808 3476 6860
rect 21364 6808 21416 6860
rect 154488 6740 154540 6792
rect 273628 6740 273680 6792
rect 159916 6672 159968 6724
rect 350448 6672 350500 6724
rect 180708 6604 180760 6656
rect 422576 6604 422628 6656
rect 181996 6536 182048 6588
rect 429660 6536 429712 6588
rect 180616 6468 180668 6520
rect 436744 6468 436796 6520
rect 179144 6400 179196 6452
rect 443828 6400 443880 6452
rect 181904 6332 181956 6384
rect 450912 6332 450964 6384
rect 165620 6264 165672 6316
rect 442632 6264 442684 6316
rect 176568 6196 176620 6248
rect 563244 6196 563296 6248
rect 87972 6128 88024 6180
rect 138204 6128 138256 6180
rect 144184 6128 144236 6180
rect 161296 6128 161348 6180
rect 182088 6128 182140 6180
rect 583392 6128 583444 6180
rect 143540 5652 143592 5704
rect 144736 5652 144788 5704
rect 138848 5516 138900 5568
rect 142528 5516 142580 5568
rect 142804 5516 142856 5568
rect 143540 5516 143592 5568
rect 151084 4972 151136 5024
rect 245200 4972 245252 5024
rect 161388 4904 161440 4956
rect 371700 4904 371752 4956
rect 168288 4836 168340 4888
rect 456892 4836 456944 4888
rect 25320 4768 25372 4820
rect 133880 4768 133932 4820
rect 173900 4768 173952 4820
rect 541992 4768 542044 4820
rect 572 4088 624 4140
rect 7564 4088 7616 4140
rect 73804 4088 73856 4140
rect 75184 4088 75236 4140
rect 83280 4088 83332 4140
rect 84844 4088 84896 4140
rect 112812 4088 112864 4140
rect 113272 4088 113324 4140
rect 148324 4088 148376 4140
rect 154212 4088 154264 4140
rect 181812 4088 181864 4140
rect 187424 4088 187476 4140
rect 188344 4088 188396 4140
rect 196808 4088 196860 4140
rect 197268 4088 197320 4140
rect 203892 4088 203944 4140
rect 207664 4088 207716 4140
rect 210976 4088 211028 4140
rect 211804 4088 211856 4140
rect 223948 4088 224000 4140
rect 242164 4088 242216 4140
rect 260656 4088 260708 4140
rect 315304 4088 315356 4140
rect 317328 4088 317380 4140
rect 323584 4088 323636 4140
rect 326804 4088 326856 4140
rect 450544 4088 450596 4140
rect 452108 4088 452160 4140
rect 180064 4020 180116 4072
rect 189816 4020 189868 4072
rect 193864 4020 193916 4072
rect 195612 4020 195664 4072
rect 195704 4020 195756 4072
rect 247592 4020 247644 4072
rect 284300 4020 284352 4072
rect 285036 4020 285088 4072
rect 287704 4020 287756 4072
rect 312636 4020 312688 4072
rect 566464 4020 566516 4072
rect 568028 4020 568080 4072
rect 146944 3952 146996 4004
rect 148508 3952 148560 4004
rect 149704 3952 149756 4004
rect 153016 3952 153068 4004
rect 182824 3952 182876 4004
rect 212172 3952 212224 4004
rect 220084 3952 220136 4004
rect 298468 3952 298520 4004
rect 299572 3952 299624 4004
rect 300768 3952 300820 4004
rect 147128 3884 147180 3936
rect 149612 3884 149664 3936
rect 179236 3884 179288 3936
rect 394240 3884 394292 3936
rect 44272 3816 44324 3868
rect 46204 3816 46256 3868
rect 148416 3816 148468 3868
rect 163688 3816 163740 3868
rect 179328 3816 179380 3868
rect 401324 3816 401376 3868
rect 122288 3748 122340 3800
rect 127072 3748 127124 3800
rect 130844 3748 130896 3800
rect 151820 3748 151872 3800
rect 152464 3748 152516 3800
rect 164516 3748 164568 3800
rect 178776 3748 178828 3800
rect 408408 3748 408460 3800
rect 119896 3680 119948 3732
rect 131488 3680 131540 3732
rect 147036 3680 147088 3732
rect 149520 3680 149572 3732
rect 149612 3680 149664 3732
rect 171968 3680 172020 3732
rect 178684 3680 178736 3732
rect 415492 3680 415544 3732
rect 454684 3680 454736 3732
rect 497096 3680 497148 3732
rect 51356 3612 51408 3664
rect 54484 3612 54536 3664
rect 65524 3612 65576 3664
rect 17040 3544 17092 3596
rect 18604 3544 18656 3596
rect 19432 3544 19484 3596
rect 21456 3544 21508 3596
rect 27620 3544 27672 3596
rect 28540 3544 28592 3596
rect 52460 3544 52512 3596
rect 53380 3544 53432 3596
rect 56048 3544 56100 3596
rect 57244 3544 57296 3596
rect 60740 3544 60792 3596
rect 61660 3544 61712 3596
rect 69112 3544 69164 3596
rect 71044 3544 71096 3596
rect 93952 3612 94004 3664
rect 125600 3612 125652 3664
rect 129832 3612 129884 3664
rect 131028 3612 131080 3664
rect 162492 3612 162544 3664
rect 179052 3612 179104 3664
rect 461584 3612 461636 3664
rect 125876 3544 125928 3596
rect 129924 3544 129976 3596
rect 130936 3544 130988 3596
rect 166080 3544 166132 3596
rect 170404 3544 170456 3596
rect 174268 3544 174320 3596
rect 185584 3544 185636 3596
rect 187332 3544 187384 3596
rect 187424 3544 187476 3596
rect 468300 3544 468352 3596
rect 468484 3544 468536 3596
rect 469864 3544 469916 3596
rect 15936 3476 15988 3528
rect 1676 3408 1728 3460
rect 8944 3408 8996 3460
rect 11152 3408 11204 3460
rect 91560 3340 91612 3392
rect 93124 3340 93176 3392
rect 101036 3340 101088 3392
rect 102784 3340 102836 3392
rect 105728 3340 105780 3392
rect 106924 3340 106976 3392
rect 110420 3340 110472 3392
rect 111616 3340 111668 3392
rect 109316 3272 109368 3324
rect 112444 3272 112496 3324
rect 123484 3476 123536 3528
rect 124864 3476 124916 3528
rect 126980 3476 127032 3528
rect 128452 3476 128504 3528
rect 136456 3476 136508 3528
rect 141516 3476 141568 3528
rect 147220 3476 147272 3528
rect 148324 3476 148376 3528
rect 148508 3476 148560 3528
rect 124680 3408 124732 3460
rect 131304 3408 131356 3460
rect 141424 3408 141476 3460
rect 131396 3340 131448 3392
rect 143448 3340 143500 3392
rect 150624 3340 150676 3392
rect 157984 3340 158036 3392
rect 158904 3340 158956 3392
rect 131580 3272 131632 3324
rect 171784 3476 171836 3528
rect 173164 3476 173216 3528
rect 178960 3476 179012 3528
rect 472624 3476 472676 3528
rect 473452 3476 473504 3528
rect 478236 3544 478288 3596
rect 500592 3544 500644 3596
rect 525064 3544 525116 3596
rect 527824 3544 527876 3596
rect 560944 3544 560996 3596
rect 564440 3544 564492 3596
rect 574744 3544 574796 3596
rect 576308 3544 576360 3596
rect 479340 3476 479392 3528
rect 506480 3476 506532 3528
rect 507308 3476 507360 3528
rect 514024 3476 514076 3528
rect 515956 3476 516008 3528
rect 538864 3476 538916 3528
rect 539600 3476 539652 3528
rect 549904 3476 549956 3528
rect 551468 3476 551520 3528
rect 554044 3476 554096 3528
rect 554964 3476 555016 3528
rect 563704 3476 563756 3528
rect 565636 3476 565688 3528
rect 567936 3476 567988 3528
rect 569132 3476 569184 3528
rect 180524 3408 180576 3460
rect 487620 3408 487672 3460
rect 511356 3408 511408 3460
rect 514760 3408 514812 3460
rect 527916 3408 527968 3460
rect 533712 3408 533764 3460
rect 567844 3408 567896 3460
rect 572720 3408 572772 3460
rect 176660 3340 176712 3392
rect 184296 3340 184348 3392
rect 189724 3340 189776 3392
rect 189816 3340 189868 3392
rect 190828 3340 190880 3392
rect 193128 3340 193180 3392
rect 195704 3340 195756 3392
rect 204168 3340 204220 3392
rect 207388 3340 207440 3392
rect 239404 3340 239456 3392
rect 240508 3340 240560 3392
rect 261484 3340 261536 3392
rect 262956 3340 263008 3392
rect 275284 3340 275336 3392
rect 277124 3340 277176 3392
rect 279424 3340 279476 3392
rect 280712 3340 280764 3392
rect 307024 3340 307076 3392
rect 309048 3340 309100 3392
rect 324412 3340 324464 3392
rect 325608 3340 325660 3392
rect 329104 3340 329156 3392
rect 330392 3340 330444 3392
rect 340972 3340 341024 3392
rect 342168 3340 342220 3392
rect 342904 3340 342956 3392
rect 344560 3340 344612 3392
rect 356704 3340 356756 3392
rect 358728 3340 358780 3392
rect 364984 3340 365036 3392
rect 367008 3340 367060 3392
rect 374092 3340 374144 3392
rect 375288 3340 375340 3392
rect 382372 3340 382424 3392
rect 383568 3340 383620 3392
rect 390560 3340 390612 3392
rect 391848 3340 391900 3392
rect 398932 3340 398984 3392
rect 400128 3340 400180 3392
rect 400864 3340 400916 3392
rect 402520 3340 402572 3392
rect 414664 3340 414716 3392
rect 416688 3340 416740 3392
rect 418804 3340 418856 3392
rect 420184 3340 420236 3392
rect 423680 3340 423732 3392
rect 424968 3340 425020 3392
rect 432604 3340 432656 3392
rect 434444 3340 434496 3392
rect 440240 3340 440292 3392
rect 441528 3340 441580 3392
rect 446404 3340 446456 3392
rect 447416 3340 447468 3392
rect 448612 3340 448664 3392
rect 449808 3340 449860 3392
rect 456800 3340 456852 3392
rect 458088 3340 458140 3392
rect 482284 3340 482336 3392
rect 484032 3340 484084 3392
rect 534724 3340 534776 3392
rect 550272 3340 550324 3392
rect 175464 3272 175516 3324
rect 189908 3272 189960 3324
rect 193220 3272 193272 3324
rect 210424 3272 210476 3324
rect 218060 3272 218112 3324
rect 224224 3272 224276 3324
rect 231032 3272 231084 3324
rect 260104 3272 260156 3324
rect 261760 3272 261812 3324
rect 396724 3272 396776 3324
rect 397736 3272 397788 3324
rect 431960 3272 432012 3324
rect 433248 3272 433300 3324
rect 520924 3272 520976 3324
rect 524236 3272 524288 3324
rect 562324 3272 562376 3324
rect 566832 3272 566884 3324
rect 571984 3272 572036 3324
rect 573916 3272 573968 3324
rect 134156 3204 134208 3256
rect 138664 3204 138716 3256
rect 33600 3136 33652 3188
rect 35164 3136 35216 3188
rect 38384 3136 38436 3188
rect 39304 3136 39356 3188
rect 41880 3136 41932 3188
rect 43444 3136 43496 3188
rect 118792 3136 118844 3188
rect 122104 3136 122156 3188
rect 164884 3136 164936 3188
rect 168380 3136 168432 3188
rect 12348 3068 12400 3120
rect 17224 3068 17276 3120
rect 382924 3068 382976 3120
rect 384764 3068 384816 3120
rect 20628 3000 20680 3052
rect 22744 3000 22796 3052
rect 175924 3000 175976 3052
rect 177856 3000 177908 3052
rect 464344 3000 464396 3052
rect 466276 3000 466328 3052
rect 132960 2932 133012 2984
rect 139492 2932 139544 2984
rect 23020 2864 23072 2916
rect 25504 2864 25556 2916
rect 128176 2864 128228 2916
rect 129004 2864 129056 2916
rect 181444 2864 181496 2916
rect 182548 2864 182600 2916
rect 332600 1096 332652 1148
rect 333888 1096 333940 1148
<< metal2 >>
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40052 703582 40356 703610
rect 8128 700534 8156 703520
rect 24320 700602 24348 703520
rect 24308 700596 24360 700602
rect 24308 700538 24360 700544
rect 8116 700528 8168 700534
rect 8116 700470 8168 700476
rect 3422 684312 3478 684321
rect 3422 684247 3478 684256
rect 3436 683262 3464 684247
rect 3424 683256 3476 683262
rect 3424 683198 3476 683204
rect 3514 671256 3570 671265
rect 3514 671191 3570 671200
rect 3528 670750 3556 671191
rect 3516 670744 3568 670750
rect 3516 670686 3568 670692
rect 3422 658200 3478 658209
rect 3422 658135 3478 658144
rect 3436 656946 3464 658135
rect 3424 656940 3476 656946
rect 3424 656882 3476 656888
rect 3424 632120 3476 632126
rect 3422 632088 3424 632097
rect 3476 632088 3478 632097
rect 3422 632023 3478 632032
rect 3146 619168 3202 619177
rect 3146 619103 3202 619112
rect 3160 618322 3188 619103
rect 3148 618316 3200 618322
rect 3148 618258 3200 618264
rect 3238 606112 3294 606121
rect 3238 606047 3294 606056
rect 3252 605878 3280 606047
rect 3240 605872 3292 605878
rect 3240 605814 3292 605820
rect 3330 580000 3386 580009
rect 3330 579935 3386 579944
rect 3344 579698 3372 579935
rect 3332 579692 3384 579698
rect 3332 579634 3384 579640
rect 3422 566944 3478 566953
rect 3422 566879 3478 566888
rect 3436 565894 3464 566879
rect 3424 565888 3476 565894
rect 3424 565830 3476 565836
rect 3422 553888 3478 553897
rect 3422 553823 3478 553832
rect 3436 553450 3464 553823
rect 3424 553444 3476 553450
rect 3424 553386 3476 553392
rect 3422 527912 3478 527921
rect 3422 527847 3478 527856
rect 3436 527202 3464 527847
rect 3424 527196 3476 527202
rect 3424 527138 3476 527144
rect 3422 514856 3478 514865
rect 3422 514791 3424 514800
rect 3476 514791 3478 514800
rect 8944 514820 8996 514826
rect 3424 514762 3476 514768
rect 8944 514762 8996 514768
rect 3054 501800 3110 501809
rect 3054 501735 3110 501744
rect 3068 501022 3096 501735
rect 3056 501016 3108 501022
rect 3056 500958 3108 500964
rect 3422 475688 3478 475697
rect 3422 475623 3478 475632
rect 3146 449576 3202 449585
rect 3146 449511 3202 449520
rect 3160 448594 3188 449511
rect 3148 448588 3200 448594
rect 3148 448530 3200 448536
rect 2870 410544 2926 410553
rect 2870 410479 2926 410488
rect 2884 409902 2912 410479
rect 2872 409896 2924 409902
rect 2872 409838 2924 409844
rect 2778 371376 2834 371385
rect 2778 371311 2780 371320
rect 2832 371311 2834 371320
rect 2780 371282 2832 371288
rect 3146 358456 3202 358465
rect 3146 358391 3202 358400
rect 3160 357474 3188 358391
rect 3148 357468 3200 357474
rect 3148 357410 3200 357416
rect 3330 319288 3386 319297
rect 3330 319223 3386 319232
rect 3344 318850 3372 319223
rect 3332 318844 3384 318850
rect 3332 318786 3384 318792
rect 3054 267200 3110 267209
rect 3054 267135 3110 267144
rect 3068 266422 3096 267135
rect 3056 266416 3108 266422
rect 3056 266358 3108 266364
rect 3436 265674 3464 475623
rect 3514 462632 3570 462641
rect 3514 462567 3570 462576
rect 3528 462398 3556 462567
rect 3516 462392 3568 462398
rect 3516 462334 3568 462340
rect 3514 423600 3570 423609
rect 3514 423535 3570 423544
rect 3528 422346 3556 423535
rect 3516 422340 3568 422346
rect 3516 422282 3568 422288
rect 3516 397520 3568 397526
rect 3514 397488 3516 397497
rect 3568 397488 3570 397497
rect 3514 397423 3570 397432
rect 4804 371340 4856 371346
rect 4804 371282 4856 371288
rect 3514 345400 3570 345409
rect 3514 345335 3570 345344
rect 3528 345234 3556 345335
rect 3516 345228 3568 345234
rect 3516 345170 3568 345176
rect 3514 306232 3570 306241
rect 3514 306167 3570 306176
rect 3528 305046 3556 306167
rect 3516 305040 3568 305046
rect 3516 304982 3568 304988
rect 3514 293176 3570 293185
rect 3514 293111 3570 293120
rect 3528 292602 3556 293111
rect 3516 292596 3568 292602
rect 3516 292538 3568 292544
rect 4816 268394 4844 371282
rect 7564 345228 7616 345234
rect 7564 345170 7616 345176
rect 7576 271250 7604 345170
rect 8956 274038 8984 514762
rect 10324 357468 10376 357474
rect 10324 357410 10376 357416
rect 10336 289134 10364 357410
rect 10324 289128 10376 289134
rect 10324 289070 10376 289076
rect 40052 279478 40080 703582
rect 40328 703474 40356 703582
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218072 703582 218836 703610
rect 40512 703474 40540 703520
rect 40328 703446 40540 703474
rect 72988 703050 73016 703520
rect 71780 703044 71832 703050
rect 71780 702986 71832 702992
rect 72976 703044 73028 703050
rect 72976 702986 73028 702992
rect 40040 279472 40092 279478
rect 40040 279414 40092 279420
rect 8944 274032 8996 274038
rect 8944 273974 8996 273980
rect 7564 271244 7616 271250
rect 7564 271186 7616 271192
rect 71792 269822 71820 702986
rect 89180 700738 89208 703520
rect 89168 700732 89220 700738
rect 89168 700674 89220 700680
rect 105464 699718 105492 703520
rect 137848 700874 137876 703520
rect 154132 702434 154160 703520
rect 170324 702434 170352 703520
rect 153212 702406 154160 702434
rect 169772 702406 170352 702434
rect 137836 700868 137888 700874
rect 137836 700810 137888 700816
rect 153108 700392 153160 700398
rect 153108 700334 153160 700340
rect 148324 700324 148376 700330
rect 148324 700266 148376 700272
rect 105452 699712 105504 699718
rect 105452 699654 105504 699660
rect 106924 699712 106976 699718
rect 106924 699654 106976 699660
rect 71780 269816 71832 269822
rect 71780 269758 71832 269764
rect 4804 268388 4856 268394
rect 4804 268330 4856 268336
rect 3424 265668 3476 265674
rect 3424 265610 3476 265616
rect 106936 264246 106964 699654
rect 146300 696992 146352 696998
rect 146300 696934 146352 696940
rect 143632 616888 143684 616894
rect 143632 616830 143684 616836
rect 142160 590708 142212 590714
rect 142160 590650 142212 590656
rect 139400 484424 139452 484430
rect 139400 484366 139452 484372
rect 138664 430636 138716 430642
rect 138664 430578 138716 430584
rect 135260 351960 135312 351966
rect 135260 351902 135312 351908
rect 134524 324352 134576 324358
rect 134524 324294 134576 324300
rect 133144 271924 133196 271930
rect 133144 271866 133196 271872
rect 121460 269816 121512 269822
rect 121460 269758 121512 269764
rect 121472 269142 121500 269758
rect 121460 269136 121512 269142
rect 121460 269078 121512 269084
rect 122380 269136 122432 269142
rect 122380 269078 122432 269084
rect 120816 264308 120868 264314
rect 120816 264250 120868 264256
rect 106924 264240 106976 264246
rect 106924 264182 106976 264188
rect 118240 264172 118292 264178
rect 118240 264114 118292 264120
rect 115572 264104 115624 264110
rect 115572 264046 115624 264052
rect 115388 263968 115440 263974
rect 115388 263910 115440 263916
rect 3424 262948 3476 262954
rect 3424 262890 3476 262896
rect 2780 241256 2832 241262
rect 2780 241198 2832 241204
rect 2792 241097 2820 241198
rect 2778 241088 2834 241097
rect 2778 241023 2834 241032
rect 3436 201929 3464 262890
rect 113824 262880 113876 262886
rect 113824 262822 113876 262828
rect 112904 262608 112956 262614
rect 112904 262550 112956 262556
rect 3516 262472 3568 262478
rect 3516 262414 3568 262420
rect 3528 254153 3556 262414
rect 111248 261112 111300 261118
rect 111248 261054 111300 261060
rect 4804 260976 4856 260982
rect 4804 260918 4856 260924
rect 3514 254144 3570 254153
rect 3514 254079 3570 254088
rect 4816 241262 4844 260918
rect 7564 259548 7616 259554
rect 7564 259490 7616 259496
rect 4804 241256 4856 241262
rect 4804 241198 4856 241204
rect 7576 215150 7604 259490
rect 3516 215144 3568 215150
rect 3516 215086 3568 215092
rect 7564 215144 7616 215150
rect 7564 215086 7616 215092
rect 3528 214985 3556 215086
rect 3514 214976 3570 214985
rect 3514 214911 3570 214920
rect 3422 201920 3478 201929
rect 3422 201855 3478 201864
rect 104440 200592 104492 200598
rect 104440 200534 104492 200540
rect 102876 199708 102928 199714
rect 102876 199650 102928 199656
rect 101770 197976 101826 197985
rect 101770 197911 101826 197920
rect 97632 197736 97684 197742
rect 97632 197678 97684 197684
rect 3424 189032 3476 189038
rect 3424 188974 3476 188980
rect 3436 188873 3464 188974
rect 3422 188864 3478 188873
rect 3422 188799 3478 188808
rect 3514 162888 3570 162897
rect 3514 162823 3570 162832
rect 3146 149832 3202 149841
rect 3146 149767 3202 149776
rect 3160 149190 3188 149767
rect 3148 149184 3200 149190
rect 3148 149126 3200 149132
rect 3528 145586 3556 162823
rect 97448 151088 97500 151094
rect 97448 151030 97500 151036
rect 3516 145580 3568 145586
rect 3516 145522 3568 145528
rect 13084 140888 13136 140894
rect 13084 140830 13136 140836
rect 8944 139528 8996 139534
rect 8944 139470 8996 139476
rect 3424 138712 3476 138718
rect 3424 138654 3476 138660
rect 3240 137964 3292 137970
rect 3240 137906 3292 137912
rect 3252 136785 3280 137906
rect 3238 136776 3294 136785
rect 3238 136711 3294 136720
rect 3056 111444 3108 111450
rect 3056 111386 3108 111392
rect 3068 110673 3096 111386
rect 3054 110664 3110 110673
rect 3054 110599 3110 110608
rect 2778 77888 2834 77897
rect 2778 77823 2834 77832
rect 2792 6914 2820 77823
rect 2870 62792 2926 62801
rect 2870 62727 2926 62736
rect 2884 16574 2912 62727
rect 3436 19417 3464 138654
rect 8956 111450 8984 139470
rect 8944 111444 8996 111450
rect 8944 111386 8996 111392
rect 6918 78024 6974 78033
rect 6918 77959 6974 77968
rect 3516 71732 3568 71738
rect 3516 71674 3568 71680
rect 3528 71641 3556 71674
rect 3514 71632 3570 71641
rect 3514 71567 3570 71576
rect 4158 59936 4214 59945
rect 4158 59871 4214 59880
rect 3422 19408 3478 19417
rect 3422 19343 3478 19352
rect 4172 16574 4200 59871
rect 6932 16574 6960 77959
rect 7562 75168 7618 75177
rect 7562 75103 7618 75112
rect 2884 16546 3648 16574
rect 4172 16546 5304 16574
rect 6932 16546 7512 16574
rect 2792 6886 2912 6914
rect 572 4140 624 4146
rect 572 4082 624 4088
rect 584 480 612 4082
rect 1676 3460 1728 3466
rect 1676 3402 1728 3408
rect 1688 480 1716 3402
rect 2884 480 2912 6886
rect 3424 6860 3476 6866
rect 3424 6802 3476 6808
rect 3436 6497 3464 6802
rect 3422 6488 3478 6497
rect 3422 6423 3478 6432
rect 542 -960 654 480
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 3620 354 3648 16546
rect 5276 480 5304 16546
rect 6460 8968 6512 8974
rect 6460 8910 6512 8916
rect 6472 480 6500 8910
rect 7484 3482 7512 16546
rect 7576 4146 7604 75103
rect 8944 73840 8996 73846
rect 8944 73782 8996 73788
rect 8298 65512 8354 65521
rect 8298 65447 8354 65456
rect 8312 16574 8340 65447
rect 8312 16546 8800 16574
rect 7564 4140 7616 4146
rect 7564 4082 7616 4088
rect 7484 3454 7696 3482
rect 7668 480 7696 3454
rect 8772 480 8800 16546
rect 8956 3466 8984 73782
rect 9680 72480 9732 72486
rect 9680 72422 9732 72428
rect 8944 3460 8996 3466
rect 8944 3402 8996 3408
rect 4038 354 4150 480
rect 3620 326 4150 354
rect 4038 -960 4150 326
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8730 -960 8842 480
rect 9692 354 9720 72422
rect 13096 71738 13124 140830
rect 21364 139596 21416 139602
rect 21364 139538 21416 139544
rect 20718 78160 20774 78169
rect 20718 78095 20774 78104
rect 13084 71732 13136 71738
rect 13084 71674 13136 71680
rect 17222 71088 17278 71097
rect 17222 71023 17278 71032
rect 12438 55856 12494 55865
rect 12438 55791 12494 55800
rect 12452 16574 12480 55791
rect 13820 37936 13872 37942
rect 13820 37878 13872 37884
rect 13832 16574 13860 37878
rect 12452 16546 13584 16574
rect 13832 16546 14320 16574
rect 11152 3460 11204 3466
rect 11152 3402 11204 3408
rect 11164 480 11192 3402
rect 12348 3120 12400 3126
rect 12348 3062 12400 3068
rect 12360 480 12388 3062
rect 13556 480 13584 16546
rect 9926 354 10038 480
rect 9692 326 10038 354
rect 9926 -960 10038 326
rect 11122 -960 11234 480
rect 12318 -960 12430 480
rect 13514 -960 13626 480
rect 14292 354 14320 16546
rect 17040 3596 17092 3602
rect 17040 3538 17092 3544
rect 15936 3528 15988 3534
rect 15936 3470 15988 3476
rect 15948 480 15976 3470
rect 17052 480 17080 3538
rect 17236 3126 17264 71023
rect 18604 68332 18656 68338
rect 18604 68274 18656 68280
rect 17960 51740 18012 51746
rect 17960 51682 18012 51688
rect 17224 3120 17276 3126
rect 17224 3062 17276 3068
rect 14710 354 14822 480
rect 14292 326 14822 354
rect 14710 -960 14822 326
rect 15906 -960 16018 480
rect 17010 -960 17122 480
rect 17972 354 18000 51682
rect 18616 3602 18644 68274
rect 20732 16574 20760 78095
rect 20732 16546 21312 16574
rect 18604 3596 18656 3602
rect 18604 3538 18656 3544
rect 19432 3596 19484 3602
rect 19432 3538 19484 3544
rect 19444 480 19472 3538
rect 21284 3482 21312 16546
rect 21376 6866 21404 139538
rect 60740 78328 60792 78334
rect 60740 78270 60792 78276
rect 57980 78124 58032 78130
rect 57980 78066 58032 78072
rect 53840 78056 53892 78062
rect 53840 77998 53892 78004
rect 46940 77988 46992 77994
rect 46940 77930 46992 77936
rect 34518 76528 34574 76537
rect 34518 76463 34574 76472
rect 22744 73908 22796 73914
rect 22744 73850 22796 73856
rect 21456 72548 21508 72554
rect 21456 72490 21508 72496
rect 21364 6860 21416 6866
rect 21364 6802 21416 6808
rect 21468 3602 21496 72490
rect 21456 3596 21508 3602
rect 21456 3538 21508 3544
rect 21284 3454 21864 3482
rect 20628 3052 20680 3058
rect 20628 2994 20680 3000
rect 20640 480 20668 2994
rect 21836 480 21864 3454
rect 22756 3058 22784 73850
rect 26240 68400 26292 68406
rect 26240 68342 26292 68348
rect 25502 57216 25558 57225
rect 25502 57151 25558 57160
rect 23480 36576 23532 36582
rect 23480 36518 23532 36524
rect 23492 16574 23520 36518
rect 23492 16546 24256 16574
rect 22744 3052 22796 3058
rect 22744 2994 22796 3000
rect 23020 2916 23072 2922
rect 23020 2858 23072 2864
rect 23032 480 23060 2858
rect 24228 480 24256 16546
rect 25320 4820 25372 4826
rect 25320 4762 25372 4768
rect 25332 480 25360 4762
rect 25516 2922 25544 57151
rect 25504 2916 25556 2922
rect 25504 2858 25556 2864
rect 18206 354 18318 480
rect 17972 326 18318 354
rect 18206 -960 18318 326
rect 19402 -960 19514 480
rect 20598 -960 20710 480
rect 21794 -960 21906 480
rect 22990 -960 23102 480
rect 24186 -960 24298 480
rect 25290 -960 25402 480
rect 26252 354 26280 68342
rect 27618 61432 27674 61441
rect 27618 61367 27674 61376
rect 27632 3602 27660 61367
rect 27710 50280 27766 50289
rect 27710 50215 27766 50224
rect 27620 3596 27672 3602
rect 27620 3538 27672 3544
rect 27724 480 27752 50215
rect 30378 48920 30434 48929
rect 30378 48855 30434 48864
rect 30392 16574 30420 48855
rect 31760 35216 31812 35222
rect 31760 35158 31812 35164
rect 31772 16574 31800 35158
rect 30392 16546 30880 16574
rect 31772 16546 31984 16574
rect 30104 10328 30156 10334
rect 30104 10270 30156 10276
rect 28540 3596 28592 3602
rect 28540 3538 28592 3544
rect 26486 354 26598 480
rect 26252 326 26598 354
rect 26486 -960 26598 326
rect 27682 -960 27794 480
rect 28552 354 28580 3538
rect 30116 480 30144 10270
rect 28878 354 28990 480
rect 28552 326 28990 354
rect 28878 -960 28990 326
rect 30074 -960 30186 480
rect 30852 354 30880 16546
rect 31270 354 31382 480
rect 30852 326 31382 354
rect 31956 354 31984 16546
rect 33600 3188 33652 3194
rect 33600 3130 33652 3136
rect 33612 480 33640 3130
rect 32374 354 32486 480
rect 31956 326 32486 354
rect 31270 -960 31382 326
rect 32374 -960 32486 326
rect 33570 -960 33682 480
rect 34532 354 34560 76463
rect 35898 75304 35954 75313
rect 35898 75239 35954 75248
rect 35164 69692 35216 69698
rect 35164 69634 35216 69640
rect 35176 3194 35204 69634
rect 35912 6914 35940 75239
rect 45560 69760 45612 69766
rect 45560 69702 45612 69708
rect 40040 66972 40092 66978
rect 40040 66914 40092 66920
rect 35992 65544 36044 65550
rect 35992 65486 36044 65492
rect 36004 16574 36032 65486
rect 39302 47560 39358 47569
rect 39302 47495 39358 47504
rect 38660 33788 38712 33794
rect 38660 33730 38712 33736
rect 38672 16574 38700 33730
rect 36004 16546 36768 16574
rect 38672 16546 39160 16574
rect 35912 6886 36032 6914
rect 35164 3188 35216 3194
rect 35164 3130 35216 3136
rect 36004 480 36032 6886
rect 34766 354 34878 480
rect 34532 326 34878 354
rect 34766 -960 34878 326
rect 35962 -960 36074 480
rect 36740 354 36768 16546
rect 38384 3188 38436 3194
rect 38384 3130 38436 3136
rect 38396 480 38424 3130
rect 37158 354 37270 480
rect 36740 326 37270 354
rect 37158 -960 37270 326
rect 38354 -960 38466 480
rect 39132 354 39160 16546
rect 39316 3194 39344 47495
rect 40052 16574 40080 66914
rect 43444 61396 43496 61402
rect 43444 61338 43496 61344
rect 42800 31068 42852 31074
rect 42800 31010 42852 31016
rect 40052 16546 40264 16574
rect 39304 3188 39356 3194
rect 39304 3130 39356 3136
rect 39550 354 39662 480
rect 39132 326 39662 354
rect 40236 354 40264 16546
rect 41880 3188 41932 3194
rect 41880 3130 41932 3136
rect 41892 480 41920 3130
rect 40654 354 40766 480
rect 40236 326 40766 354
rect 39550 -960 39662 326
rect 40654 -960 40766 326
rect 41850 -960 41962 480
rect 42812 354 42840 31010
rect 43456 3194 43484 61338
rect 44178 46200 44234 46209
rect 44178 46135 44234 46144
rect 44192 16574 44220 46135
rect 45572 16574 45600 69702
rect 46204 26920 46256 26926
rect 46204 26862 46256 26868
rect 44192 16546 45048 16574
rect 45572 16546 46152 16574
rect 44272 3868 44324 3874
rect 44272 3810 44324 3816
rect 43444 3188 43496 3194
rect 43444 3130 43496 3136
rect 44284 480 44312 3810
rect 43046 354 43158 480
rect 42812 326 43158 354
rect 43046 -960 43158 326
rect 44242 -960 44354 480
rect 45020 354 45048 16546
rect 46124 3482 46152 16546
rect 46216 3874 46244 26862
rect 46952 16574 46980 77930
rect 52458 71224 52514 71233
rect 52458 71159 52514 71168
rect 48320 68468 48372 68474
rect 48320 68410 48372 68416
rect 48332 16574 48360 68410
rect 49698 53136 49754 53145
rect 49698 53071 49754 53080
rect 49712 16574 49740 53071
rect 46952 16546 47440 16574
rect 48332 16546 48544 16574
rect 49712 16546 50200 16574
rect 46204 3868 46256 3874
rect 46204 3810 46256 3816
rect 46124 3454 46704 3482
rect 46676 480 46704 3454
rect 45438 354 45550 480
rect 45020 326 45550 354
rect 45438 -960 45550 326
rect 46634 -960 46746 480
rect 47412 354 47440 16546
rect 47830 354 47942 480
rect 47412 326 47942 354
rect 48516 354 48544 16546
rect 50172 480 50200 16546
rect 51356 3664 51408 3670
rect 51356 3606 51408 3612
rect 51368 480 51396 3606
rect 52472 3602 52500 71159
rect 52552 60036 52604 60042
rect 52552 59978 52604 59984
rect 52460 3596 52512 3602
rect 52460 3538 52512 3544
rect 52564 480 52592 59978
rect 53852 16574 53880 77998
rect 54482 73808 54538 73817
rect 54482 73743 54538 73752
rect 53852 16546 54432 16574
rect 53380 3596 53432 3602
rect 53380 3538 53432 3544
rect 48934 354 49046 480
rect 48516 326 49046 354
rect 47830 -960 47942 326
rect 48934 -960 49046 326
rect 50130 -960 50242 480
rect 51326 -960 51438 480
rect 52522 -960 52634 480
rect 53392 354 53420 3538
rect 54404 3482 54432 16546
rect 54496 3670 54524 73743
rect 57244 64184 57296 64190
rect 57244 64126 57296 64132
rect 56598 54496 56654 54505
rect 56598 54431 56654 54440
rect 56612 16574 56640 54431
rect 56612 16546 56824 16574
rect 54484 3664 54536 3670
rect 54484 3606 54536 3612
rect 56048 3596 56100 3602
rect 56048 3538 56100 3544
rect 54404 3454 54984 3482
rect 54956 480 54984 3454
rect 56060 480 56088 3538
rect 53718 354 53830 480
rect 53392 326 53830 354
rect 53718 -960 53830 326
rect 54914 -960 55026 480
rect 56018 -960 56130 480
rect 56796 354 56824 16546
rect 57256 3602 57284 64126
rect 57992 16574 58020 78066
rect 59360 76560 59412 76566
rect 59360 76502 59412 76508
rect 57992 16546 58480 16574
rect 57244 3596 57296 3602
rect 57244 3538 57296 3544
rect 58452 480 58480 16546
rect 57214 354 57326 480
rect 56796 326 57326 354
rect 57214 -960 57326 326
rect 58410 -960 58522 480
rect 59372 354 59400 76502
rect 60752 3602 60780 78270
rect 75920 78260 75972 78266
rect 75920 78202 75972 78208
rect 67640 76696 67692 76702
rect 67640 76638 67692 76644
rect 66260 76628 66312 76634
rect 66260 76570 66312 76576
rect 62120 64252 62172 64258
rect 62120 64194 62172 64200
rect 60830 55992 60886 56001
rect 60830 55927 60886 55936
rect 60740 3596 60792 3602
rect 60740 3538 60792 3544
rect 60844 480 60872 55927
rect 62132 16574 62160 64194
rect 63498 43480 63554 43489
rect 63498 43415 63554 43424
rect 63512 16574 63540 43415
rect 66272 16574 66300 76570
rect 62132 16546 63264 16574
rect 63512 16546 64368 16574
rect 66272 16546 66760 16574
rect 61660 3596 61712 3602
rect 61660 3538 61712 3544
rect 59606 354 59718 480
rect 59372 326 59718 354
rect 59606 -960 59718 326
rect 60802 -960 60914 480
rect 61672 354 61700 3538
rect 63236 480 63264 16546
rect 64340 480 64368 16546
rect 65524 3664 65576 3670
rect 65524 3606 65576 3612
rect 65536 480 65564 3606
rect 66732 480 66760 16546
rect 61998 354 62110 480
rect 61672 326 62110 354
rect 61998 -960 62110 326
rect 63194 -960 63306 480
rect 64298 -960 64410 480
rect 65494 -960 65606 480
rect 66690 -960 66802 480
rect 67652 354 67680 76638
rect 71042 75440 71098 75449
rect 71042 75375 71098 75384
rect 69020 62824 69072 62830
rect 69020 62766 69072 62772
rect 69032 16574 69060 62766
rect 70400 42084 70452 42090
rect 70400 42026 70452 42032
rect 70412 16574 70440 42026
rect 69032 16546 69888 16574
rect 70412 16546 70992 16574
rect 69112 3596 69164 3602
rect 69112 3538 69164 3544
rect 69124 480 69152 3538
rect 67886 354 67998 480
rect 67652 326 67998 354
rect 67886 -960 67998 326
rect 69082 -960 69194 480
rect 69860 354 69888 16546
rect 70964 3482 70992 16546
rect 71056 3602 71084 75375
rect 71780 71052 71832 71058
rect 71780 70994 71832 71000
rect 71792 16574 71820 70994
rect 75182 61568 75238 61577
rect 75182 61503 75238 61512
rect 74540 40724 74592 40730
rect 74540 40666 74592 40672
rect 74552 16574 74580 40666
rect 71792 16546 72648 16574
rect 74552 16546 75040 16574
rect 71044 3596 71096 3602
rect 71044 3538 71096 3544
rect 70964 3454 71544 3482
rect 71516 480 71544 3454
rect 72620 480 72648 16546
rect 73804 4140 73856 4146
rect 73804 4082 73856 4088
rect 73816 480 73844 4082
rect 75012 480 75040 16546
rect 75196 4146 75224 61503
rect 75184 4140 75236 4146
rect 75184 4082 75236 4088
rect 70278 354 70390 480
rect 69860 326 70390 354
rect 70278 -960 70390 326
rect 71474 -960 71586 480
rect 72578 -960 72690 480
rect 73774 -960 73886 480
rect 74970 -960 75082 480
rect 75932 354 75960 78202
rect 85580 75268 85632 75274
rect 85580 75210 85632 75216
rect 78678 72448 78734 72457
rect 78678 72383 78734 72392
rect 77298 66872 77354 66881
rect 77298 66807 77354 66816
rect 77312 6914 77340 66807
rect 77392 39364 77444 39370
rect 77392 39306 77444 39312
rect 77404 16574 77432 39306
rect 78692 16574 78720 72383
rect 84844 71120 84896 71126
rect 84844 71062 84896 71068
rect 81438 60072 81494 60081
rect 81438 60007 81494 60016
rect 80058 57352 80114 57361
rect 80058 57287 80114 57296
rect 80072 16574 80100 57287
rect 81452 16574 81480 60007
rect 84198 55176 84254 55185
rect 84198 55111 84254 55120
rect 77404 16546 78168 16574
rect 78692 16546 79272 16574
rect 80072 16546 80928 16574
rect 81452 16546 81664 16574
rect 77312 6886 77432 6914
rect 77404 480 77432 6886
rect 76166 354 76278 480
rect 75932 326 76278 354
rect 76166 -960 76278 326
rect 77362 -960 77474 480
rect 78140 354 78168 16546
rect 78558 354 78670 480
rect 78140 326 78670 354
rect 79244 354 79272 16546
rect 80900 480 80928 16546
rect 79662 354 79774 480
rect 79244 326 79774 354
rect 78558 -960 78670 326
rect 79662 -960 79774 326
rect 80858 -960 80970 480
rect 81636 354 81664 16546
rect 83280 4140 83332 4146
rect 83280 4082 83332 4088
rect 83292 480 83320 4082
rect 82054 354 82166 480
rect 81636 326 82166 354
rect 82054 -960 82166 326
rect 83250 -960 83362 480
rect 84212 354 84240 55111
rect 84856 4146 84884 71062
rect 85592 6914 85620 75210
rect 89720 73976 89772 73982
rect 89720 73918 89772 73924
rect 85672 69828 85724 69834
rect 85672 69770 85724 69776
rect 85684 16574 85712 69770
rect 88338 62928 88394 62937
rect 88338 62863 88394 62872
rect 88352 16574 88380 62863
rect 89732 16574 89760 73918
rect 96620 72888 96672 72894
rect 96620 72830 96672 72836
rect 93122 65648 93178 65657
rect 93122 65583 93178 65592
rect 92478 58712 92534 58721
rect 92478 58647 92534 58656
rect 85684 16546 86448 16574
rect 88352 16546 89208 16574
rect 89732 16546 89944 16574
rect 85592 6886 85712 6914
rect 84844 4140 84896 4146
rect 84844 4082 84896 4088
rect 85684 480 85712 6886
rect 84446 354 84558 480
rect 84212 326 84558 354
rect 84446 -960 84558 326
rect 85642 -960 85754 480
rect 86420 354 86448 16546
rect 87972 6180 88024 6186
rect 87972 6122 88024 6128
rect 87984 480 88012 6122
rect 89180 480 89208 16546
rect 86838 354 86950 480
rect 86420 326 86950 354
rect 86838 -960 86950 326
rect 87942 -960 88054 480
rect 89138 -960 89250 480
rect 89916 354 89944 16546
rect 91560 3392 91612 3398
rect 91560 3334 91612 3340
rect 91572 480 91600 3334
rect 90334 354 90446 480
rect 89916 326 90446 354
rect 90334 -960 90446 326
rect 91530 -960 91642 480
rect 92492 354 92520 58647
rect 93136 3398 93164 65583
rect 93858 58848 93914 58857
rect 93858 58783 93914 58792
rect 93872 16574 93900 58783
rect 95238 50416 95294 50425
rect 95238 50351 95294 50360
rect 95252 16574 95280 50351
rect 96632 16574 96660 72830
rect 97460 66910 97488 151030
rect 97540 148436 97592 148442
rect 97540 148378 97592 148384
rect 97448 66904 97500 66910
rect 97448 66846 97500 66852
rect 97552 58585 97580 148378
rect 97644 77246 97672 197678
rect 97722 195392 97778 195401
rect 97722 195327 97778 195336
rect 97632 77240 97684 77246
rect 97632 77182 97684 77188
rect 97644 76702 97672 77182
rect 97632 76696 97684 76702
rect 97632 76638 97684 76644
rect 97736 73166 97764 195327
rect 97908 193928 97960 193934
rect 97908 193870 97960 193876
rect 97816 193860 97868 193866
rect 97816 193802 97868 193808
rect 97724 73160 97776 73166
rect 97724 73102 97776 73108
rect 97828 71777 97856 193802
rect 97814 71768 97870 71777
rect 97814 71703 97870 71712
rect 97920 70174 97948 193870
rect 101680 193044 101732 193050
rect 101680 192986 101732 192992
rect 99104 192636 99156 192642
rect 99104 192578 99156 192584
rect 99012 187128 99064 187134
rect 99012 187070 99064 187076
rect 98920 164892 98972 164898
rect 98920 164834 98972 164840
rect 98828 151564 98880 151570
rect 98828 151506 98880 151512
rect 98736 148572 98788 148578
rect 98736 148514 98788 148520
rect 98748 72486 98776 148514
rect 98840 73030 98868 151506
rect 98932 78606 98960 164834
rect 98920 78600 98972 78606
rect 98920 78542 98972 78548
rect 98828 73024 98880 73030
rect 98828 72966 98880 72972
rect 98840 72554 98868 72966
rect 99024 72962 99052 187070
rect 99116 76673 99144 192578
rect 100666 191584 100722 191593
rect 100666 191519 100722 191528
rect 99196 191208 99248 191214
rect 99196 191150 99248 191156
rect 100574 191176 100630 191185
rect 99102 76664 99158 76673
rect 99102 76599 99158 76608
rect 99208 75206 99236 191150
rect 100574 191111 100630 191120
rect 100484 187264 100536 187270
rect 100484 187206 100536 187212
rect 100300 187060 100352 187066
rect 100300 187002 100352 187008
rect 99286 186960 99342 186969
rect 99286 186895 99342 186904
rect 99196 75200 99248 75206
rect 99196 75142 99248 75148
rect 99012 72956 99064 72962
rect 99012 72898 99064 72904
rect 98828 72548 98880 72554
rect 98828 72490 98880 72496
rect 98736 72480 98788 72486
rect 98736 72422 98788 72428
rect 98748 72282 98776 72422
rect 98736 72276 98788 72282
rect 98736 72218 98788 72224
rect 97908 70168 97960 70174
rect 97908 70110 97960 70116
rect 97998 64152 98054 64161
rect 97998 64087 98054 64096
rect 97538 58576 97594 58585
rect 97538 58511 97594 58520
rect 98012 16574 98040 64087
rect 99300 60625 99328 186895
rect 99840 151768 99892 151774
rect 99840 151710 99892 151716
rect 99852 77217 99880 151710
rect 100116 151700 100168 151706
rect 100116 151642 100168 151648
rect 100024 151496 100076 151502
rect 100024 151438 100076 151444
rect 99932 151292 99984 151298
rect 99932 151234 99984 151240
rect 99838 77208 99894 77217
rect 99838 77143 99894 77152
rect 99378 76800 99434 76809
rect 99378 76735 99434 76744
rect 98826 60616 98882 60625
rect 98826 60551 98882 60560
rect 99286 60616 99342 60625
rect 99286 60551 99342 60560
rect 98840 59945 98868 60551
rect 98826 59936 98882 59945
rect 98826 59871 98882 59880
rect 99392 16574 99420 76735
rect 99944 75857 99972 151234
rect 99470 75848 99526 75857
rect 99470 75783 99526 75792
rect 99930 75848 99986 75857
rect 99930 75783 99986 75792
rect 99484 75313 99512 75783
rect 99470 75304 99526 75313
rect 99470 75239 99526 75248
rect 100036 71369 100064 151438
rect 100022 71360 100078 71369
rect 100022 71295 100078 71304
rect 100128 70378 100156 151642
rect 100208 151632 100260 151638
rect 100208 151574 100260 151580
rect 100116 70372 100168 70378
rect 100116 70314 100168 70320
rect 100220 64874 100248 151574
rect 100312 78849 100340 187002
rect 100392 186992 100444 186998
rect 100392 186934 100444 186940
rect 100298 78840 100354 78849
rect 100298 78775 100354 78784
rect 100404 74390 100432 186934
rect 100392 74384 100444 74390
rect 100392 74326 100444 74332
rect 100404 73914 100432 74326
rect 100392 73908 100444 73914
rect 100392 73850 100444 73856
rect 100128 64846 100248 64874
rect 100128 62121 100156 64846
rect 100114 62112 100170 62121
rect 100114 62047 100170 62056
rect 100128 61441 100156 62047
rect 100114 61432 100170 61441
rect 100114 61367 100170 61376
rect 100496 52426 100524 187206
rect 99472 52420 99524 52426
rect 99472 52362 99524 52368
rect 100484 52420 100536 52426
rect 100484 52362 100536 52368
rect 99484 51746 99512 52362
rect 99472 51740 99524 51746
rect 99472 51682 99524 51688
rect 100588 50969 100616 191111
rect 99470 50960 99526 50969
rect 99470 50895 99526 50904
rect 100574 50960 100630 50969
rect 100574 50895 100630 50904
rect 99484 50289 99512 50895
rect 99470 50280 99526 50289
rect 99470 50215 99526 50224
rect 100680 49609 100708 191519
rect 101588 189848 101640 189854
rect 101588 189790 101640 189796
rect 101496 187196 101548 187202
rect 101496 187138 101548 187144
rect 101404 151428 101456 151434
rect 101404 151370 101456 151376
rect 101312 151360 101364 151366
rect 101312 151302 101364 151308
rect 101220 148504 101272 148510
rect 101220 148446 101272 148452
rect 101232 71641 101260 148446
rect 101218 71632 101274 71641
rect 101218 71567 101274 71576
rect 101324 70310 101352 151302
rect 100760 70304 100812 70310
rect 100760 70246 100812 70252
rect 101312 70304 101364 70310
rect 101312 70246 101364 70252
rect 100772 69766 100800 70246
rect 100760 69760 100812 69766
rect 100760 69702 100812 69708
rect 101416 66162 101444 151370
rect 101508 77081 101536 187138
rect 101494 77072 101550 77081
rect 101494 77007 101550 77016
rect 101600 68814 101628 189790
rect 101588 68808 101640 68814
rect 101588 68750 101640 68756
rect 101692 68406 101720 192986
rect 101680 68400 101732 68406
rect 101680 68342 101732 68348
rect 101784 68338 101812 197911
rect 101862 196752 101918 196761
rect 101862 196687 101918 196696
rect 101772 68332 101824 68338
rect 101772 68274 101824 68280
rect 101404 66156 101456 66162
rect 101404 66098 101456 66104
rect 101876 57905 101904 196687
rect 102784 193112 102836 193118
rect 102784 193054 102836 193060
rect 102046 191312 102102 191321
rect 102046 191247 102102 191256
rect 101954 191040 102010 191049
rect 101954 190975 102010 190984
rect 100758 57896 100814 57905
rect 100758 57831 100814 57840
rect 101862 57896 101918 57905
rect 101862 57831 101918 57840
rect 100772 57225 100800 57831
rect 100758 57216 100814 57225
rect 100758 57151 100814 57160
rect 99470 49600 99526 49609
rect 99470 49535 99526 49544
rect 100666 49600 100722 49609
rect 100666 49535 100722 49544
rect 99484 48929 99512 49535
rect 99470 48920 99526 48929
rect 99470 48855 99526 48864
rect 101968 48249 101996 190975
rect 100758 48240 100814 48249
rect 100758 48175 100814 48184
rect 101954 48240 102010 48249
rect 101954 48175 102010 48184
rect 100772 47569 100800 48175
rect 100758 47560 100814 47569
rect 100758 47495 100814 47504
rect 102060 46889 102088 191247
rect 102600 151020 102652 151026
rect 102600 150962 102652 150968
rect 102612 80753 102640 150962
rect 102690 146976 102746 146985
rect 102690 146911 102746 146920
rect 102598 80744 102654 80753
rect 102598 80679 102654 80688
rect 102140 69964 102192 69970
rect 102140 69906 102192 69912
rect 102152 69698 102180 69906
rect 102140 69692 102192 69698
rect 102140 69634 102192 69640
rect 102140 66020 102192 66026
rect 102140 65962 102192 65968
rect 102152 65550 102180 65962
rect 102140 65544 102192 65550
rect 102140 65486 102192 65492
rect 102140 62076 102192 62082
rect 102140 62018 102192 62024
rect 102152 61402 102180 62018
rect 102140 61396 102192 61402
rect 102140 61338 102192 61344
rect 102140 60716 102192 60722
rect 102140 60658 102192 60664
rect 102152 60042 102180 60658
rect 102140 60036 102192 60042
rect 102140 59978 102192 59984
rect 102138 53272 102194 53281
rect 102138 53207 102194 53216
rect 100758 46880 100814 46889
rect 100758 46815 100814 46824
rect 102046 46880 102102 46889
rect 102046 46815 102102 46824
rect 100772 46209 100800 46815
rect 100758 46200 100814 46209
rect 100758 46135 100814 46144
rect 102152 16574 102180 53207
rect 102704 44169 102732 146911
rect 102796 75585 102824 193054
rect 102888 75750 102916 199650
rect 104346 196616 104402 196625
rect 104346 196551 104402 196560
rect 103336 194472 103388 194478
rect 103336 194414 103388 194420
rect 102968 194404 103020 194410
rect 102968 194346 103020 194352
rect 102876 75744 102928 75750
rect 102876 75686 102928 75692
rect 102782 75576 102838 75585
rect 102782 75511 102838 75520
rect 102980 69970 103008 194346
rect 103244 194336 103296 194342
rect 103244 194278 103296 194284
rect 103060 189916 103112 189922
rect 103060 189858 103112 189864
rect 102968 69964 103020 69970
rect 102968 69906 103020 69912
rect 102784 69760 102836 69766
rect 102784 69702 102836 69708
rect 102230 44160 102286 44169
rect 102230 44095 102286 44104
rect 102690 44160 102746 44169
rect 102690 44095 102746 44104
rect 102244 43489 102272 44095
rect 102230 43480 102286 43489
rect 102230 43415 102286 43424
rect 93872 16546 94728 16574
rect 95252 16546 95832 16574
rect 96632 16546 97488 16574
rect 98012 16546 98224 16574
rect 99392 16546 99880 16574
rect 102152 16546 102272 16574
rect 93952 3664 94004 3670
rect 93952 3606 94004 3612
rect 93124 3392 93176 3398
rect 93124 3334 93176 3340
rect 93964 480 93992 3606
rect 92726 354 92838 480
rect 92492 326 92838 354
rect 92726 -960 92838 326
rect 93922 -960 94034 480
rect 94700 354 94728 16546
rect 95118 354 95230 480
rect 94700 326 95230 354
rect 95804 354 95832 16546
rect 97460 480 97488 16546
rect 96222 354 96334 480
rect 95804 326 96334 354
rect 95118 -960 95230 326
rect 96222 -960 96334 326
rect 97418 -960 97530 480
rect 98196 354 98224 16546
rect 99852 480 99880 16546
rect 101036 3392 101088 3398
rect 101036 3334 101088 3340
rect 101048 480 101076 3334
rect 102244 480 102272 16546
rect 102796 3398 102824 69702
rect 103072 64870 103100 189858
rect 103152 187332 103204 187338
rect 103152 187274 103204 187280
rect 103060 64864 103112 64870
rect 103060 64806 103112 64812
rect 103072 64258 103100 64806
rect 103060 64252 103112 64258
rect 103060 64194 103112 64200
rect 103164 62082 103192 187274
rect 103256 67318 103284 194278
rect 103244 67312 103296 67318
rect 103244 67254 103296 67260
rect 103348 66026 103376 194414
rect 104256 193996 104308 194002
rect 104256 193938 104308 193944
rect 104164 191276 104216 191282
rect 104164 191218 104216 191224
rect 103428 190188 103480 190194
rect 103428 190130 103480 190136
rect 103336 66020 103388 66026
rect 103336 65962 103388 65968
rect 103152 62076 103204 62082
rect 103152 62018 103204 62024
rect 103440 60722 103468 190130
rect 104072 189984 104124 189990
rect 104072 189926 104124 189932
rect 103980 146872 104032 146878
rect 103980 146814 104032 146820
rect 103992 84194 104020 146814
rect 103900 84166 104020 84194
rect 103900 75274 103928 84166
rect 103980 78532 104032 78538
rect 103980 78474 104032 78480
rect 103992 75721 104020 78474
rect 104084 77042 104112 189926
rect 104176 77110 104204 191218
rect 104164 77104 104216 77110
rect 104164 77046 104216 77052
rect 104072 77036 104124 77042
rect 104072 76978 104124 76984
rect 103978 75712 104034 75721
rect 103978 75647 104034 75656
rect 103888 75268 103940 75274
rect 103888 75210 103940 75216
rect 104268 74526 104296 193938
rect 104360 78538 104388 196551
rect 104348 78532 104400 78538
rect 104348 78474 104400 78480
rect 104452 78266 104480 200534
rect 106004 199640 106056 199646
rect 106004 199582 106056 199588
rect 107290 199608 107346 199617
rect 105820 198484 105872 198490
rect 105820 198426 105872 198432
rect 105634 198112 105690 198121
rect 105634 198047 105690 198056
rect 105542 197024 105598 197033
rect 105542 196959 105598 196968
rect 104530 195800 104586 195809
rect 104530 195735 104586 195744
rect 104440 78260 104492 78266
rect 104440 78202 104492 78208
rect 104452 77654 104480 78202
rect 104440 77648 104492 77654
rect 104440 77590 104492 77596
rect 104440 77104 104492 77110
rect 104440 77046 104492 77052
rect 104348 77036 104400 77042
rect 104348 76978 104400 76984
rect 104360 76566 104388 76978
rect 104452 76634 104480 77046
rect 104440 76628 104492 76634
rect 104440 76570 104492 76576
rect 104348 76560 104400 76566
rect 104348 76502 104400 76508
rect 104440 75268 104492 75274
rect 104440 75210 104492 75216
rect 104452 75070 104480 75210
rect 104440 75064 104492 75070
rect 104440 75006 104492 75012
rect 104256 74520 104308 74526
rect 104256 74462 104308 74468
rect 104268 73982 104296 74462
rect 104256 73976 104308 73982
rect 104256 73918 104308 73924
rect 104544 71534 104572 195735
rect 104624 195492 104676 195498
rect 104624 195434 104676 195440
rect 104256 71528 104308 71534
rect 104256 71470 104308 71476
rect 104532 71528 104584 71534
rect 104532 71470 104584 71476
rect 104268 71058 104296 71470
rect 104256 71052 104308 71058
rect 104256 70994 104308 71000
rect 103520 70440 103572 70446
rect 103520 70382 103572 70388
rect 103428 60716 103480 60722
rect 103428 60658 103480 60664
rect 103532 16574 103560 70382
rect 104636 70242 104664 195434
rect 104716 190256 104768 190262
rect 104716 190198 104768 190204
rect 104624 70236 104676 70242
rect 104624 70178 104676 70184
rect 104636 69834 104664 70178
rect 104624 69828 104676 69834
rect 104624 69770 104676 69776
rect 104624 65884 104676 65890
rect 104624 65826 104676 65832
rect 104636 65521 104664 65826
rect 104622 65512 104678 65521
rect 104622 65447 104678 65456
rect 104728 64802 104756 190198
rect 104806 187096 104862 187105
rect 104806 187031 104862 187040
rect 104716 64796 104768 64802
rect 104716 64738 104768 64744
rect 104728 64190 104756 64738
rect 104716 64184 104768 64190
rect 104716 64126 104768 64132
rect 104440 56568 104492 56574
rect 104440 56510 104492 56516
rect 104452 56001 104480 56510
rect 104438 55992 104494 56001
rect 104438 55927 104494 55936
rect 104820 55185 104848 187031
rect 105452 148096 105504 148102
rect 105452 148038 105504 148044
rect 105360 147076 105412 147082
rect 105360 147018 105412 147024
rect 105268 80300 105320 80306
rect 105268 80242 105320 80248
rect 105280 78305 105308 80242
rect 105266 78296 105322 78305
rect 105266 78231 105322 78240
rect 105372 60489 105400 147018
rect 105358 60480 105414 60489
rect 105358 60415 105414 60424
rect 104806 55176 104862 55185
rect 104806 55111 104862 55120
rect 105464 55049 105492 148038
rect 105556 80186 105584 196959
rect 105648 80306 105676 198047
rect 105728 194064 105780 194070
rect 105728 194006 105780 194012
rect 105636 80300 105688 80306
rect 105636 80242 105688 80248
rect 105556 80158 105676 80186
rect 105648 78402 105676 80158
rect 105636 78396 105688 78402
rect 105636 78338 105688 78344
rect 105648 78062 105676 78338
rect 105636 78056 105688 78062
rect 105636 77998 105688 78004
rect 105740 71670 105768 194006
rect 105832 73846 105860 198426
rect 105912 196648 105964 196654
rect 105912 196590 105964 196596
rect 105820 73840 105872 73846
rect 105820 73782 105872 73788
rect 105832 73642 105860 73782
rect 105820 73636 105872 73642
rect 105820 73578 105872 73584
rect 105924 72894 105952 196590
rect 105912 72888 105964 72894
rect 105912 72830 105964 72836
rect 105728 71664 105780 71670
rect 105728 71606 105780 71612
rect 105740 70446 105768 71606
rect 106016 71466 106044 199582
rect 107290 199543 107346 199552
rect 107108 198348 107160 198354
rect 107108 198290 107160 198296
rect 107016 197056 107068 197062
rect 107016 196998 107068 197004
rect 106096 191412 106148 191418
rect 106096 191354 106148 191360
rect 106004 71460 106056 71466
rect 106004 71402 106056 71408
rect 105728 70440 105780 70446
rect 105728 70382 105780 70388
rect 106108 63510 106136 191354
rect 106924 191140 106976 191146
rect 106924 191082 106976 191088
rect 106186 190224 106242 190233
rect 106186 190159 106242 190168
rect 106096 63504 106148 63510
rect 106096 63446 106148 63452
rect 106108 62830 106136 63446
rect 106096 62824 106148 62830
rect 106096 62766 106148 62772
rect 106200 61985 106228 190159
rect 106830 189816 106886 189825
rect 106830 189751 106886 189760
rect 106646 187232 106702 187241
rect 106646 187167 106702 187176
rect 106278 73672 106334 73681
rect 106278 73607 106334 73616
rect 106186 61976 106242 61985
rect 106186 61911 106242 61920
rect 105450 55040 105506 55049
rect 105450 54975 105506 54984
rect 105464 54505 105492 54975
rect 105450 54496 105506 54505
rect 105450 54431 105506 54440
rect 106292 16574 106320 73607
rect 106660 53689 106688 187167
rect 106740 146940 106792 146946
rect 106740 146882 106792 146888
rect 106752 64190 106780 146882
rect 106844 78674 106872 189751
rect 106832 78668 106884 78674
rect 106832 78610 106884 78616
rect 106936 75274 106964 191082
rect 107028 77926 107056 196998
rect 107120 77994 107148 198290
rect 107200 198212 107252 198218
rect 107200 198154 107252 198160
rect 107212 78334 107240 198154
rect 107200 78328 107252 78334
rect 107200 78270 107252 78276
rect 107304 78130 107332 199543
rect 110328 198280 110380 198286
rect 110328 198222 110380 198228
rect 110236 198144 110288 198150
rect 110236 198086 110288 198092
rect 108672 198076 108724 198082
rect 108672 198018 108724 198024
rect 107384 194268 107436 194274
rect 107384 194210 107436 194216
rect 107292 78124 107344 78130
rect 107292 78066 107344 78072
rect 107108 77988 107160 77994
rect 107108 77930 107160 77936
rect 107016 77920 107068 77926
rect 107016 77862 107068 77868
rect 106924 75268 106976 75274
rect 106924 75210 106976 75216
rect 106830 74080 106886 74089
rect 106830 74015 106886 74024
rect 106844 73846 106872 74015
rect 106832 73840 106884 73846
rect 106830 73808 106832 73817
rect 106884 73808 106886 73817
rect 106830 73743 106886 73752
rect 107396 70038 107424 194210
rect 108304 192568 108356 192574
rect 108304 192510 108356 192516
rect 108210 189680 108266 189689
rect 108210 189615 108266 189624
rect 107474 187368 107530 187377
rect 107474 187303 107530 187312
rect 107384 70032 107436 70038
rect 107384 69974 107436 69980
rect 107396 69766 107424 69974
rect 107384 69760 107436 69766
rect 107384 69702 107436 69708
rect 106924 68604 106976 68610
rect 106924 68546 106976 68552
rect 106740 64184 106792 64190
rect 106740 64126 106792 64132
rect 106646 53680 106702 53689
rect 106646 53615 106702 53624
rect 106660 53281 106688 53615
rect 106646 53272 106702 53281
rect 106646 53207 106702 53216
rect 103532 16546 104112 16574
rect 106292 16546 106504 16574
rect 103336 7608 103388 7614
rect 103336 7550 103388 7556
rect 102784 3392 102836 3398
rect 102784 3334 102836 3340
rect 103348 480 103376 7550
rect 98614 354 98726 480
rect 98196 326 98726 354
rect 98614 -960 98726 326
rect 99810 -960 99922 480
rect 101006 -960 101118 480
rect 102202 -960 102314 480
rect 103306 -960 103418 480
rect 104084 354 104112 16546
rect 105728 3392 105780 3398
rect 105728 3334 105780 3340
rect 105740 480 105768 3334
rect 104502 354 104614 480
rect 104084 326 104614 354
rect 104502 -960 104614 326
rect 105698 -960 105810 480
rect 106476 354 106504 16546
rect 106936 3398 106964 68546
rect 107488 57769 107516 187303
rect 108120 147212 108172 147218
rect 108120 147154 108172 147160
rect 107568 78668 107620 78674
rect 107568 78610 107620 78616
rect 107580 77586 107608 78610
rect 107568 77580 107620 77586
rect 107568 77522 107620 77528
rect 107580 69018 107608 77522
rect 107660 73228 107712 73234
rect 107660 73170 107712 73176
rect 107568 69012 107620 69018
rect 107568 68954 107620 68960
rect 107474 57760 107530 57769
rect 107474 57695 107530 57704
rect 107672 16574 107700 73170
rect 108132 65958 108160 147154
rect 108224 79422 108252 189615
rect 108316 80714 108344 192510
rect 108396 192500 108448 192506
rect 108396 192442 108448 192448
rect 108304 80708 108356 80714
rect 108304 80650 108356 80656
rect 108212 79416 108264 79422
rect 108212 79358 108264 79364
rect 108408 77994 108436 192442
rect 108580 191344 108632 191350
rect 108580 191286 108632 191292
rect 108486 190088 108542 190097
rect 108486 190023 108542 190032
rect 108396 77988 108448 77994
rect 108396 77930 108448 77936
rect 108500 75002 108528 190023
rect 108592 75886 108620 191286
rect 108684 79354 108712 198018
rect 109868 196784 109920 196790
rect 109868 196726 109920 196732
rect 108856 195560 108908 195566
rect 108856 195502 108908 195508
rect 108764 192908 108816 192914
rect 108764 192850 108816 192856
rect 108672 79348 108724 79354
rect 108672 79290 108724 79296
rect 108580 75880 108632 75886
rect 108580 75822 108632 75828
rect 108488 74996 108540 75002
rect 108488 74938 108540 74944
rect 108776 74118 108804 192850
rect 108764 74112 108816 74118
rect 108764 74054 108816 74060
rect 108776 73234 108804 74054
rect 108764 73228 108816 73234
rect 108764 73170 108816 73176
rect 108302 73128 108358 73137
rect 108302 73063 108358 73072
rect 108316 72622 108344 73063
rect 108304 72616 108356 72622
rect 108304 72558 108356 72564
rect 108316 72457 108344 72558
rect 108302 72448 108358 72457
rect 108302 72383 108358 72392
rect 108868 68746 108896 195502
rect 108948 194200 109000 194206
rect 108948 194142 109000 194148
rect 108856 68740 108908 68746
rect 108856 68682 108908 68688
rect 108960 67522 108988 194142
rect 109684 189780 109736 189786
rect 109684 189722 109736 189728
rect 109592 187400 109644 187406
rect 109592 187342 109644 187348
rect 109500 147144 109552 147150
rect 109500 147086 109552 147092
rect 108948 67516 109000 67522
rect 108948 67458 109000 67464
rect 109040 67244 109092 67250
rect 109040 67186 109092 67192
rect 109052 66881 109080 67186
rect 109038 66872 109094 66881
rect 109038 66807 109094 66816
rect 108304 66088 108356 66094
rect 108304 66030 108356 66036
rect 108120 65952 108172 65958
rect 108120 65894 108172 65900
rect 108316 65657 108344 66030
rect 108302 65648 108358 65657
rect 108302 65583 108358 65592
rect 109512 65550 109540 147086
rect 109604 81122 109632 187342
rect 109592 81116 109644 81122
rect 109592 81058 109644 81064
rect 109696 74458 109724 189722
rect 109776 187468 109828 187474
rect 109776 187410 109828 187416
rect 109684 74452 109736 74458
rect 109684 74394 109736 74400
rect 109788 68610 109816 187410
rect 109880 74254 109908 196726
rect 109960 195696 110012 195702
rect 109960 195638 110012 195644
rect 109868 74248 109920 74254
rect 109868 74190 109920 74196
rect 109972 72690 110000 195638
rect 110144 194132 110196 194138
rect 110144 194074 110196 194080
rect 110050 189952 110106 189961
rect 110050 189887 110106 189896
rect 109960 72684 110012 72690
rect 109960 72626 110012 72632
rect 109776 68604 109828 68610
rect 109776 68546 109828 68552
rect 110064 67561 110092 189887
rect 110156 68882 110184 194074
rect 110144 68876 110196 68882
rect 110144 68818 110196 68824
rect 110248 68105 110276 198086
rect 110340 68950 110368 198222
rect 111156 195424 111208 195430
rect 111156 195366 111208 195372
rect 111064 190052 111116 190058
rect 111064 189994 111116 190000
rect 110788 148844 110840 148850
rect 110788 148786 110840 148792
rect 110420 78464 110472 78470
rect 110420 78406 110472 78412
rect 110328 68944 110380 68950
rect 110328 68886 110380 68892
rect 110234 68096 110290 68105
rect 110234 68031 110290 68040
rect 110050 67552 110106 67561
rect 110050 67487 110106 67496
rect 109500 65544 109552 65550
rect 109500 65486 109552 65492
rect 107672 16546 108160 16574
rect 106924 3392 106976 3398
rect 106924 3334 106976 3340
rect 108132 480 108160 16546
rect 110432 3398 110460 78406
rect 110800 71058 110828 148786
rect 110972 147416 111024 147422
rect 110972 147358 111024 147364
rect 110878 144120 110934 144129
rect 110878 144055 110934 144064
rect 110892 78470 110920 144055
rect 110880 78464 110932 78470
rect 110880 78406 110932 78412
rect 110984 72418 111012 147358
rect 111076 80850 111104 189994
rect 111064 80844 111116 80850
rect 111064 80786 111116 80792
rect 111168 80782 111196 195366
rect 111260 146062 111288 261054
rect 111432 261044 111484 261050
rect 111432 260986 111484 260992
rect 111340 195288 111392 195294
rect 111340 195230 111392 195236
rect 111248 146056 111300 146062
rect 111248 145998 111300 146004
rect 111246 145888 111302 145897
rect 111246 145823 111302 145832
rect 111260 144430 111288 145823
rect 111248 144424 111300 144430
rect 111248 144366 111300 144372
rect 111248 141976 111300 141982
rect 111248 141918 111300 141924
rect 111156 80776 111208 80782
rect 111156 80718 111208 80724
rect 110972 72412 111024 72418
rect 110972 72354 111024 72360
rect 110788 71052 110840 71058
rect 110788 70994 110840 71000
rect 111260 65822 111288 141918
rect 111352 79626 111380 195230
rect 111444 144294 111472 260986
rect 112628 260908 112680 260914
rect 112628 260850 112680 260856
rect 111708 196920 111760 196926
rect 111708 196862 111760 196868
rect 111616 195628 111668 195634
rect 111616 195570 111668 195576
rect 111524 190120 111576 190126
rect 111524 190062 111576 190068
rect 111432 144288 111484 144294
rect 111432 144230 111484 144236
rect 111340 79620 111392 79626
rect 111340 79562 111392 79568
rect 111536 68513 111564 190062
rect 111628 73001 111656 195570
rect 111720 74186 111748 196862
rect 112640 151814 112668 260850
rect 112720 196988 112772 196994
rect 112720 196930 112772 196936
rect 112364 151786 112668 151814
rect 112076 148980 112128 148986
rect 112076 148922 112128 148928
rect 111708 74180 111760 74186
rect 111708 74122 111760 74128
rect 111800 73772 111852 73778
rect 111800 73714 111852 73720
rect 111812 73681 111840 73714
rect 111798 73672 111854 73681
rect 111798 73607 111854 73616
rect 111614 72992 111670 73001
rect 111614 72927 111670 72936
rect 112088 69834 112116 148922
rect 112168 148912 112220 148918
rect 112168 148854 112220 148860
rect 112180 69902 112208 148854
rect 112364 146130 112392 151786
rect 112536 149048 112588 149054
rect 112536 148990 112588 148996
rect 112444 147484 112496 147490
rect 112444 147426 112496 147432
rect 112352 146124 112404 146130
rect 112352 146066 112404 146072
rect 112260 143200 112312 143206
rect 112260 143142 112312 143148
rect 112272 81297 112300 143142
rect 112350 138816 112406 138825
rect 112350 138751 112406 138760
rect 112258 81288 112314 81297
rect 112258 81223 112314 81232
rect 112364 70281 112392 138751
rect 112456 76498 112484 147426
rect 112444 76492 112496 76498
rect 112444 76434 112496 76440
rect 112548 71262 112576 148990
rect 112628 147008 112680 147014
rect 112628 146950 112680 146956
rect 112640 141846 112668 146950
rect 112628 141840 112680 141846
rect 112628 141782 112680 141788
rect 112732 76566 112760 196930
rect 112812 195356 112864 195362
rect 112812 195298 112864 195304
rect 112720 76560 112772 76566
rect 112720 76502 112772 76508
rect 112824 75818 112852 195298
rect 112916 147014 112944 262550
rect 113640 260024 113692 260030
rect 113640 259966 113692 259972
rect 113088 200456 113140 200462
rect 113088 200398 113140 200404
rect 112996 200388 113048 200394
rect 112996 200330 113048 200336
rect 112904 147008 112956 147014
rect 112904 146950 112956 146956
rect 112902 144800 112958 144809
rect 112902 144735 112958 144744
rect 112916 143614 112944 144735
rect 112904 143608 112956 143614
rect 112904 143550 112956 143556
rect 112812 75812 112864 75818
rect 112812 75754 112864 75760
rect 113008 73914 113036 200330
rect 112996 73908 113048 73914
rect 112996 73850 113048 73856
rect 112536 71256 112588 71262
rect 112536 71198 112588 71204
rect 112350 70272 112406 70281
rect 112350 70207 112406 70216
rect 112168 69896 112220 69902
rect 112168 69838 112220 69844
rect 112076 69828 112128 69834
rect 112076 69770 112128 69776
rect 113100 69766 113128 200398
rect 113652 148374 113680 259966
rect 113730 192672 113786 192681
rect 113730 192607 113786 192616
rect 113640 148368 113692 148374
rect 113640 148310 113692 148316
rect 113456 148164 113508 148170
rect 113456 148106 113508 148112
rect 113180 75880 113232 75886
rect 113180 75822 113232 75828
rect 113192 74534 113220 75822
rect 113468 75313 113496 148106
rect 113548 145716 113600 145722
rect 113548 145658 113600 145664
rect 113560 78946 113588 145658
rect 113640 140072 113692 140078
rect 113640 140014 113692 140020
rect 113652 79694 113680 140014
rect 113640 79688 113692 79694
rect 113640 79630 113692 79636
rect 113548 78940 113600 78946
rect 113548 78882 113600 78888
rect 113744 77178 113772 192607
rect 113836 146198 113864 262822
rect 113916 262812 113968 262818
rect 113916 262754 113968 262760
rect 113928 146266 113956 262754
rect 115296 262676 115348 262682
rect 115296 262618 115348 262624
rect 114008 260092 114060 260098
rect 114008 260034 114060 260040
rect 113916 146260 113968 146266
rect 113916 146202 113968 146208
rect 113824 146192 113876 146198
rect 113824 146134 113876 146140
rect 113824 145376 113876 145382
rect 113824 145318 113876 145324
rect 113836 79150 113864 145318
rect 114020 141914 114048 260034
rect 114928 199572 114980 199578
rect 114928 199514 114980 199520
rect 114376 199096 114428 199102
rect 114376 199038 114428 199044
rect 114284 197192 114336 197198
rect 114284 197134 114336 197140
rect 114192 196852 114244 196858
rect 114192 196794 114244 196800
rect 114100 195832 114152 195838
rect 114100 195774 114152 195780
rect 114008 141908 114060 141914
rect 114008 141850 114060 141856
rect 113824 79144 113876 79150
rect 113824 79086 113876 79092
rect 113732 77172 113784 77178
rect 113732 77114 113784 77120
rect 114112 76838 114140 195774
rect 114204 76974 114232 196794
rect 114192 76968 114244 76974
rect 114192 76910 114244 76916
rect 114100 76832 114152 76838
rect 114006 76800 114062 76809
rect 114296 76786 114324 197134
rect 114100 76774 114152 76780
rect 114006 76735 114062 76744
rect 114204 76758 114324 76786
rect 114020 76702 114048 76735
rect 114008 76696 114060 76702
rect 114008 76638 114060 76644
rect 114204 75614 114232 76758
rect 114284 76628 114336 76634
rect 114284 76570 114336 76576
rect 114296 75886 114324 76570
rect 114284 75880 114336 75886
rect 114284 75822 114336 75828
rect 114192 75608 114244 75614
rect 114192 75550 114244 75556
rect 113454 75304 113510 75313
rect 113454 75239 113510 75248
rect 113192 74506 113312 74534
rect 113088 69760 113140 69766
rect 113088 69702 113140 69708
rect 112442 68912 112498 68921
rect 112442 68847 112498 68856
rect 111522 68504 111578 68513
rect 111522 68439 111578 68448
rect 111248 65816 111300 65822
rect 111248 65758 111300 65764
rect 111248 64728 111300 64734
rect 111248 64670 111300 64676
rect 111260 64161 111288 64670
rect 111246 64152 111302 64161
rect 111246 64087 111302 64096
rect 110510 58576 110566 58585
rect 110510 58511 110566 58520
rect 110420 3392 110472 3398
rect 110420 3334 110472 3340
rect 109316 3324 109368 3330
rect 109316 3266 109368 3272
rect 109328 480 109356 3266
rect 110524 480 110552 58511
rect 111616 3392 111668 3398
rect 111616 3334 111668 3340
rect 111628 480 111656 3334
rect 112456 3330 112484 68847
rect 113180 66904 113232 66910
rect 113180 66846 113232 66852
rect 112812 4140 112864 4146
rect 112812 4082 112864 4088
rect 112444 3324 112496 3330
rect 112444 3266 112496 3272
rect 112824 480 112852 4082
rect 113192 3482 113220 66846
rect 113284 4146 113312 74506
rect 114388 71126 114416 199038
rect 114468 196716 114520 196722
rect 114468 196658 114520 196664
rect 114376 71120 114428 71126
rect 114376 71062 114428 71068
rect 114480 67590 114508 196658
rect 114836 148640 114888 148646
rect 114836 148582 114888 148588
rect 114848 70854 114876 148582
rect 114940 72758 114968 199514
rect 115204 195900 115256 195906
rect 115204 195842 115256 195848
rect 115112 192840 115164 192846
rect 115112 192782 115164 192788
rect 115020 145648 115072 145654
rect 115020 145590 115072 145596
rect 115032 78878 115060 145590
rect 115124 79014 115152 192782
rect 115216 80918 115244 195842
rect 115308 145450 115336 262618
rect 115400 145518 115428 263910
rect 115478 187640 115534 187649
rect 115478 187575 115534 187584
rect 115388 145512 115440 145518
rect 115388 145454 115440 145460
rect 115296 145444 115348 145450
rect 115296 145386 115348 145392
rect 115296 140208 115348 140214
rect 115296 140150 115348 140156
rect 115204 80912 115256 80918
rect 115204 80854 115256 80860
rect 115112 79008 115164 79014
rect 115112 78950 115164 78956
rect 115020 78872 115072 78878
rect 115020 78814 115072 78820
rect 115308 74225 115336 140150
rect 115386 138952 115442 138961
rect 115386 138887 115442 138896
rect 115294 74216 115350 74225
rect 115294 74151 115350 74160
rect 114928 72752 114980 72758
rect 114928 72694 114980 72700
rect 114836 70848 114888 70854
rect 114836 70790 114888 70796
rect 114560 69012 114612 69018
rect 114560 68954 114612 68960
rect 114468 67584 114520 67590
rect 114468 67526 114520 67532
rect 114572 16574 114600 68954
rect 115400 67454 115428 138887
rect 115492 68921 115520 187575
rect 115584 148306 115612 264046
rect 116768 263016 116820 263022
rect 116768 262958 116820 262964
rect 116676 262744 116728 262750
rect 116676 262686 116728 262692
rect 116584 260228 116636 260234
rect 116584 260170 116636 260176
rect 115664 198960 115716 198966
rect 115664 198902 115716 198908
rect 115572 148300 115624 148306
rect 115572 148242 115624 148248
rect 115570 146296 115626 146305
rect 115570 146231 115626 146240
rect 115584 144566 115612 146231
rect 115572 144560 115624 144566
rect 115572 144502 115624 144508
rect 115676 76906 115704 198902
rect 115756 195764 115808 195770
rect 115756 195706 115808 195712
rect 115664 76900 115716 76906
rect 115664 76842 115716 76848
rect 115768 72865 115796 195706
rect 116216 192772 116268 192778
rect 116216 192714 116268 192720
rect 115848 148300 115900 148306
rect 115848 148242 115900 148248
rect 115860 144906 115888 148242
rect 115848 144900 115900 144906
rect 115848 144842 115900 144848
rect 115846 144800 115902 144809
rect 115846 144735 115902 144744
rect 115860 142118 115888 144735
rect 115848 142112 115900 142118
rect 115848 142054 115900 142060
rect 115754 72856 115810 72865
rect 115754 72791 115810 72800
rect 115940 70168 115992 70174
rect 115940 70110 115992 70116
rect 115478 68912 115534 68921
rect 115478 68847 115534 68856
rect 115388 67448 115440 67454
rect 115388 67390 115440 67396
rect 115112 63436 115164 63442
rect 115112 63378 115164 63384
rect 115124 63345 115152 63378
rect 115110 63336 115166 63345
rect 115110 63271 115166 63280
rect 115124 62937 115152 63271
rect 115110 62928 115166 62937
rect 115110 62863 115166 62872
rect 115952 16574 115980 70110
rect 116228 67386 116256 192714
rect 116596 151814 116624 260170
rect 116412 151786 116624 151814
rect 116308 145852 116360 145858
rect 116308 145794 116360 145800
rect 116320 80986 116348 145794
rect 116412 142050 116440 151786
rect 116492 145784 116544 145790
rect 116492 145726 116544 145732
rect 116400 142044 116452 142050
rect 116400 141986 116452 141992
rect 116400 140140 116452 140146
rect 116400 140082 116452 140088
rect 116308 80980 116360 80986
rect 116308 80922 116360 80928
rect 116412 79082 116440 140082
rect 116504 79218 116532 145726
rect 116688 143410 116716 262686
rect 116676 143404 116728 143410
rect 116676 143346 116728 143352
rect 116780 143342 116808 262958
rect 118148 262404 118200 262410
rect 118148 262346 118200 262352
rect 118056 261180 118108 261186
rect 118056 261122 118108 261128
rect 117872 259956 117924 259962
rect 117872 259898 117924 259904
rect 117136 199164 117188 199170
rect 117136 199106 117188 199112
rect 116952 199028 117004 199034
rect 116952 198970 117004 198976
rect 116860 197124 116912 197130
rect 116860 197066 116912 197072
rect 116768 143336 116820 143342
rect 116768 143278 116820 143284
rect 116676 140276 116728 140282
rect 116676 140218 116728 140224
rect 116492 79212 116544 79218
rect 116492 79154 116544 79160
rect 116400 79076 116452 79082
rect 116400 79018 116452 79024
rect 116688 74322 116716 140218
rect 116766 139224 116822 139233
rect 116766 139159 116822 139168
rect 116676 74316 116728 74322
rect 116676 74258 116728 74264
rect 116216 67380 116268 67386
rect 116216 67322 116268 67328
rect 116780 67289 116808 139159
rect 116872 75682 116900 197066
rect 116964 76809 116992 198970
rect 117044 192976 117096 192982
rect 117044 192918 117096 192924
rect 116950 76800 117006 76809
rect 116950 76735 117006 76744
rect 116860 75676 116912 75682
rect 116860 75618 116912 75624
rect 117056 69601 117084 192918
rect 117148 75546 117176 199106
rect 117884 151814 117912 259898
rect 117964 259480 118016 259486
rect 117964 259422 118016 259428
rect 117792 151786 117912 151814
rect 117688 148708 117740 148714
rect 117688 148650 117740 148656
rect 117226 144800 117282 144809
rect 117226 144735 117282 144744
rect 117240 143682 117268 144735
rect 117594 144256 117650 144265
rect 117594 144191 117650 144200
rect 117228 143676 117280 143682
rect 117228 143618 117280 143624
rect 117226 143440 117282 143449
rect 117226 143375 117282 143384
rect 117240 141506 117268 143375
rect 117228 141500 117280 141506
rect 117228 141442 117280 141448
rect 117136 75540 117188 75546
rect 117136 75482 117188 75488
rect 117608 71330 117636 144191
rect 117596 71324 117648 71330
rect 117596 71266 117648 71272
rect 117228 70916 117280 70922
rect 117228 70858 117280 70864
rect 117240 70174 117268 70858
rect 117700 70174 117728 148650
rect 117792 144634 117820 151786
rect 117976 146690 118004 259422
rect 117884 146662 118004 146690
rect 117780 144628 117832 144634
rect 117780 144570 117832 144576
rect 117780 144492 117832 144498
rect 117780 144434 117832 144440
rect 117792 137306 117820 144434
rect 117884 141710 117912 146662
rect 118068 143274 118096 261122
rect 118160 144226 118188 262346
rect 118148 144220 118200 144226
rect 118148 144162 118200 144168
rect 118146 143984 118202 143993
rect 118146 143919 118202 143928
rect 118160 143750 118188 143919
rect 118148 143744 118200 143750
rect 118148 143686 118200 143692
rect 118056 143268 118108 143274
rect 118056 143210 118108 143216
rect 118252 142154 118280 264114
rect 119804 263900 119856 263906
rect 119804 263842 119856 263848
rect 119712 263764 119764 263770
rect 119712 263706 119764 263712
rect 119344 260840 119396 260846
rect 119344 260782 119396 260788
rect 119068 200524 119120 200530
rect 119068 200466 119120 200472
rect 118608 200252 118660 200258
rect 118608 200194 118660 200200
rect 118332 199504 118384 199510
rect 118332 199446 118384 199452
rect 117976 142126 118280 142154
rect 117976 141778 118004 142126
rect 117964 141772 118016 141778
rect 117964 141714 118016 141720
rect 117872 141704 117924 141710
rect 117872 141646 117924 141652
rect 118148 140412 118200 140418
rect 118148 140354 118200 140360
rect 117964 140344 118016 140350
rect 117964 140286 118016 140292
rect 117792 137278 117912 137306
rect 117780 136468 117832 136474
rect 117780 136410 117832 136416
rect 117792 79490 117820 136410
rect 117884 80481 117912 137278
rect 117870 80472 117926 80481
rect 117870 80407 117926 80416
rect 117780 79484 117832 79490
rect 117780 79426 117832 79432
rect 117976 76770 118004 140286
rect 118056 140004 118108 140010
rect 118056 139946 118108 139952
rect 117964 76764 118016 76770
rect 117964 76706 118016 76712
rect 118068 71602 118096 139946
rect 118160 136474 118188 140354
rect 118148 136468 118200 136474
rect 118148 136410 118200 136416
rect 118344 76945 118372 199446
rect 118424 199232 118476 199238
rect 118424 199174 118476 199180
rect 118330 76936 118386 76945
rect 118330 76871 118386 76880
rect 118436 75478 118464 199174
rect 118514 197160 118570 197169
rect 118514 197095 118570 197104
rect 118424 75472 118476 75478
rect 118424 75414 118476 75420
rect 118528 72729 118556 197095
rect 118620 72826 118648 200194
rect 118976 148776 119028 148782
rect 118976 148718 119028 148724
rect 118884 147348 118936 147354
rect 118884 147290 118936 147296
rect 118792 144356 118844 144362
rect 118792 144298 118844 144304
rect 118700 139664 118752 139670
rect 118700 139606 118752 139612
rect 118712 137970 118740 139606
rect 118700 137964 118752 137970
rect 118700 137906 118752 137912
rect 118608 72820 118660 72826
rect 118608 72762 118660 72768
rect 118514 72720 118570 72729
rect 118514 72655 118570 72664
rect 118056 71596 118108 71602
rect 118056 71538 118108 71544
rect 117228 70168 117280 70174
rect 117228 70110 117280 70116
rect 117688 70168 117740 70174
rect 117688 70110 117740 70116
rect 118804 70106 118832 144298
rect 118896 77518 118924 147290
rect 118988 79257 119016 148718
rect 118974 79248 119030 79257
rect 118974 79183 119030 79192
rect 118884 77512 118936 77518
rect 118884 77454 118936 77460
rect 119080 72486 119108 200466
rect 119356 149122 119384 260782
rect 119436 259888 119488 259894
rect 119436 259830 119488 259836
rect 119344 149116 119396 149122
rect 119344 149058 119396 149064
rect 119356 141574 119384 149058
rect 119448 146169 119476 259830
rect 119528 259820 119580 259826
rect 119528 259762 119580 259768
rect 119434 146160 119490 146169
rect 119434 146095 119490 146104
rect 119540 142866 119568 259762
rect 119620 259752 119672 259758
rect 119620 259694 119672 259700
rect 119528 142860 119580 142866
rect 119528 142802 119580 142808
rect 119528 142384 119580 142390
rect 119528 142326 119580 142332
rect 119344 141568 119396 141574
rect 119344 141510 119396 141516
rect 119436 141432 119488 141438
rect 119436 141374 119488 141380
rect 119252 140616 119304 140622
rect 119252 140558 119304 140564
rect 119264 79286 119292 140558
rect 119344 140480 119396 140486
rect 119344 140422 119396 140428
rect 119252 79280 119304 79286
rect 119252 79222 119304 79228
rect 119356 79121 119384 140422
rect 119448 79558 119476 141374
rect 119540 139505 119568 142326
rect 119632 141642 119660 259694
rect 119724 142769 119752 263706
rect 119816 142934 119844 263842
rect 120724 263696 120776 263702
rect 120724 263638 120776 263644
rect 120540 259616 120592 259622
rect 120540 259558 120592 259564
rect 119896 200320 119948 200326
rect 119896 200262 119948 200268
rect 119804 142928 119856 142934
rect 119804 142870 119856 142876
rect 119710 142760 119766 142769
rect 119710 142695 119766 142704
rect 119620 141636 119672 141642
rect 119620 141578 119672 141584
rect 119712 140752 119764 140758
rect 119712 140694 119764 140700
rect 119526 139496 119582 139505
rect 119526 139431 119582 139440
rect 119436 79552 119488 79558
rect 119436 79494 119488 79500
rect 119342 79112 119398 79121
rect 119342 79047 119398 79056
rect 119068 72480 119120 72486
rect 119068 72422 119120 72428
rect 119724 71738 119752 140694
rect 119908 74050 119936 200262
rect 120552 189038 120580 259558
rect 120632 195968 120684 195974
rect 120632 195910 120684 195916
rect 120540 189032 120592 189038
rect 120540 188974 120592 188980
rect 120448 145920 120500 145926
rect 120448 145862 120500 145868
rect 120172 142316 120224 142322
rect 120172 142258 120224 142264
rect 120184 138718 120212 142258
rect 120172 138712 120224 138718
rect 120172 138654 120224 138660
rect 120460 80889 120488 145862
rect 120446 80880 120502 80889
rect 120446 80815 120502 80824
rect 120644 75138 120672 195910
rect 120736 143002 120764 263638
rect 120828 143138 120856 264250
rect 121460 264240 121512 264246
rect 121460 264182 121512 264188
rect 120908 264036 120960 264042
rect 120908 263978 120960 263984
rect 120816 143132 120868 143138
rect 120816 143074 120868 143080
rect 120920 143070 120948 263978
rect 121472 263634 121500 264182
rect 121460 263628 121512 263634
rect 121460 263570 121512 263576
rect 122012 263628 122064 263634
rect 122012 263570 122064 263576
rect 121920 262540 121972 262546
rect 121920 262482 121972 262488
rect 121368 199368 121420 199374
rect 121368 199310 121420 199316
rect 121274 198928 121330 198937
rect 121274 198863 121330 198872
rect 121184 198824 121236 198830
rect 121184 198766 121236 198772
rect 121000 197328 121052 197334
rect 121000 197270 121052 197276
rect 120908 143064 120960 143070
rect 120908 143006 120960 143012
rect 120724 142996 120776 143002
rect 120724 142938 120776 142944
rect 120908 140548 120960 140554
rect 120908 140490 120960 140496
rect 120722 138680 120778 138689
rect 120722 138615 120778 138624
rect 120736 81977 120764 138615
rect 120814 86184 120870 86193
rect 120814 86119 120870 86128
rect 120722 81968 120778 81977
rect 120722 81903 120778 81912
rect 120828 80617 120856 86119
rect 120814 80608 120870 80617
rect 120814 80543 120870 80552
rect 120632 75132 120684 75138
rect 120632 75074 120684 75080
rect 119896 74044 119948 74050
rect 119896 73986 119948 73992
rect 119712 71732 119764 71738
rect 119712 71674 119764 71680
rect 120920 71398 120948 140490
rect 121012 75410 121040 197270
rect 121092 197260 121144 197266
rect 121092 197202 121144 197208
rect 121000 75404 121052 75410
rect 121000 75346 121052 75352
rect 121104 72554 121132 197202
rect 121196 75342 121224 198766
rect 121184 75336 121236 75342
rect 121184 75278 121236 75284
rect 121288 73982 121316 198863
rect 121276 73976 121328 73982
rect 121276 73918 121328 73924
rect 121092 72548 121144 72554
rect 121092 72490 121144 72496
rect 121380 72350 121408 199310
rect 121828 187536 121880 187542
rect 121828 187478 121880 187484
rect 121644 152584 121696 152590
rect 121644 152526 121696 152532
rect 121552 152516 121604 152522
rect 121552 152458 121604 152464
rect 121458 81288 121514 81297
rect 121458 81223 121514 81232
rect 121472 77625 121500 81223
rect 121458 77616 121514 77625
rect 121458 77551 121514 77560
rect 121368 72344 121420 72350
rect 121368 72286 121420 72292
rect 120908 71392 120960 71398
rect 120908 71334 120960 71340
rect 121564 70990 121592 152458
rect 121552 70984 121604 70990
rect 121552 70926 121604 70932
rect 121656 70786 121684 152526
rect 121840 133929 121868 187478
rect 121932 153882 121960 262482
rect 121920 153876 121972 153882
rect 121920 153818 121972 153824
rect 122024 151230 122052 263570
rect 122196 198620 122248 198626
rect 122196 198562 122248 198568
rect 122104 194540 122156 194546
rect 122104 194482 122156 194488
rect 122012 151224 122064 151230
rect 122012 151166 122064 151172
rect 121920 147280 121972 147286
rect 121920 147222 121972 147228
rect 121826 133920 121882 133929
rect 121826 133855 121882 133864
rect 121734 86048 121790 86057
rect 121734 85983 121790 85992
rect 121644 70780 121696 70786
rect 121644 70722 121696 70728
rect 118792 70100 118844 70106
rect 118792 70042 118844 70048
rect 117042 69592 117098 69601
rect 117042 69527 117098 69536
rect 121748 68882 121776 85983
rect 121932 80578 121960 147222
rect 122012 81116 122064 81122
rect 122012 81058 122064 81064
rect 121920 80572 121972 80578
rect 121920 80514 121972 80520
rect 121826 80200 121882 80209
rect 121826 80135 121882 80144
rect 121736 68876 121788 68882
rect 121736 68818 121788 68824
rect 116766 67280 116822 67289
rect 116766 67215 116822 67224
rect 121840 66230 121868 80135
rect 121920 79416 121972 79422
rect 121920 79358 121972 79364
rect 121932 77926 121960 79358
rect 121920 77920 121972 77926
rect 121920 77862 121972 77868
rect 122024 77450 122052 81058
rect 122116 78130 122144 194482
rect 122208 81161 122236 198562
rect 122288 198416 122340 198422
rect 122288 198358 122340 198364
rect 122194 81152 122250 81161
rect 122194 81087 122250 81096
rect 122300 81025 122328 198358
rect 122392 151162 122420 269078
rect 133156 264110 133184 271866
rect 134248 264172 134300 264178
rect 134248 264114 134300 264120
rect 133144 264104 133196 264110
rect 133144 264046 133196 264052
rect 122564 263832 122616 263838
rect 122564 263774 122616 263780
rect 122472 262268 122524 262274
rect 122472 262210 122524 262216
rect 122484 199442 122512 262210
rect 122472 199436 122524 199442
rect 122472 199378 122524 199384
rect 122472 191480 122524 191486
rect 122472 191422 122524 191428
rect 122380 151156 122432 151162
rect 122380 151098 122432 151104
rect 122378 81968 122434 81977
rect 122378 81903 122434 81912
rect 122286 81016 122342 81025
rect 122286 80951 122342 80960
rect 122288 80776 122340 80782
rect 122288 80718 122340 80724
rect 122300 80510 122328 80718
rect 122288 80504 122340 80510
rect 122288 80446 122340 80452
rect 122104 78124 122156 78130
rect 122104 78066 122156 78072
rect 122104 77920 122156 77926
rect 122104 77862 122156 77868
rect 122012 77444 122064 77450
rect 122012 77386 122064 77392
rect 121828 66224 121880 66230
rect 121828 66166 121880 66172
rect 117320 65544 117372 65550
rect 117320 65486 117372 65492
rect 114572 16546 114784 16574
rect 115952 16546 116440 16574
rect 113272 4140 113324 4146
rect 113272 4082 113324 4088
rect 113192 3454 114048 3482
rect 114020 480 114048 3454
rect 106894 354 107006 480
rect 106476 326 107006 354
rect 106894 -960 107006 326
rect 108090 -960 108202 480
rect 109286 -960 109398 480
rect 110482 -960 110594 480
rect 111586 -960 111698 480
rect 112782 -960 112894 480
rect 113978 -960 114090 480
rect 114756 354 114784 16546
rect 116412 480 116440 16546
rect 115174 354 115286 480
rect 114756 326 115286 354
rect 115174 -960 115286 326
rect 116370 -960 116482 480
rect 117332 354 117360 65486
rect 120080 64184 120132 64190
rect 120080 64126 120132 64132
rect 120092 16574 120120 64126
rect 120092 16546 120672 16574
rect 119896 3732 119948 3738
rect 119896 3674 119948 3680
rect 118792 3188 118844 3194
rect 118792 3130 118844 3136
rect 118804 480 118832 3130
rect 119908 480 119936 3674
rect 117566 354 117678 480
rect 117332 326 117678 354
rect 117566 -960 117678 326
rect 118762 -960 118874 480
rect 119866 -960 119978 480
rect 120644 354 120672 16546
rect 122116 3194 122144 77862
rect 122392 74089 122420 81903
rect 122378 74080 122434 74089
rect 122378 74015 122434 74024
rect 122484 73098 122512 191422
rect 122576 145994 122604 263774
rect 127346 263120 127402 263129
rect 127346 263055 127402 263064
rect 125598 262440 125654 262449
rect 125598 262375 125654 262384
rect 124312 260840 124364 260846
rect 123206 260808 123262 260817
rect 124312 260782 124364 260788
rect 123206 260743 123262 260752
rect 123220 259978 123248 260743
rect 124324 259978 124352 260782
rect 125612 259978 125640 262375
rect 125968 262268 126020 262274
rect 125968 262210 126020 262216
rect 125980 259978 126008 262210
rect 127254 260128 127310 260137
rect 126842 260092 126894 260098
rect 127254 260063 127310 260072
rect 126842 260034 126894 260040
rect 123220 259950 123556 259978
rect 124324 259950 124660 259978
rect 125612 259950 125764 259978
rect 125980 259950 126316 259978
rect 126854 259964 126882 260034
rect 127268 259729 127296 260063
rect 127360 259978 127388 263055
rect 131120 263016 131172 263022
rect 131120 262958 131172 262964
rect 132040 263016 132092 263022
rect 132040 262958 132092 262964
rect 127716 262744 127768 262750
rect 127716 262686 127768 262692
rect 127622 260536 127678 260545
rect 127622 260471 127678 260480
rect 127636 260137 127664 260471
rect 127622 260128 127678 260137
rect 127622 260063 127678 260072
rect 127728 259978 127756 262686
rect 129832 262676 129884 262682
rect 129832 262618 129884 262624
rect 128728 262608 128780 262614
rect 128728 262550 128780 262556
rect 128360 260024 128412 260030
rect 127360 259950 127420 259978
rect 127728 259950 127972 259978
rect 128740 259978 128768 262550
rect 129280 262404 129332 262410
rect 129280 262346 129332 262352
rect 129292 259978 129320 262346
rect 129844 261458 129872 262618
rect 129832 261452 129884 261458
rect 129832 261394 129884 261400
rect 129844 259978 129872 261394
rect 131132 261322 131160 262958
rect 131764 262880 131816 262886
rect 131764 262822 131816 262828
rect 131120 261316 131172 261322
rect 131120 261258 131172 261264
rect 130384 261044 130436 261050
rect 130384 260986 130436 260992
rect 130396 259978 130424 260986
rect 131132 259978 131160 261258
rect 131776 259978 131804 262822
rect 132052 261118 132080 262958
rect 132868 261180 132920 261186
rect 132868 261122 132920 261128
rect 132040 261112 132092 261118
rect 132040 261054 132092 261060
rect 132052 259978 132080 261054
rect 132880 260250 132908 261122
rect 132880 260222 132954 260250
rect 132926 260166 132954 260222
rect 132914 260160 132966 260166
rect 132914 260102 132966 260108
rect 128412 259972 128524 259978
rect 128360 259966 128524 259972
rect 128372 259950 128524 259966
rect 128740 259950 129076 259978
rect 129292 259950 129628 259978
rect 129844 259950 130180 259978
rect 130396 259950 130732 259978
rect 131132 259950 131284 259978
rect 131776 259950 131836 259978
rect 132052 259950 132388 259978
rect 132926 259964 132954 260102
rect 133156 259978 133184 264046
rect 133972 260908 134024 260914
rect 133972 260850 134024 260856
rect 133984 259978 134012 260850
rect 134260 259978 134288 264114
rect 134536 262818 134564 324294
rect 134616 298172 134668 298178
rect 134616 298114 134668 298120
rect 134628 264178 134656 298114
rect 134616 264172 134668 264178
rect 134616 264114 134668 264120
rect 134524 262812 134576 262818
rect 134524 262754 134576 262760
rect 134800 262812 134852 262818
rect 134800 262754 134852 262760
rect 134812 259978 134840 262754
rect 135272 260234 135300 351902
rect 135904 311908 135956 311914
rect 135904 311850 135956 311856
rect 135916 265169 135944 311850
rect 137284 286340 137336 286346
rect 137284 286282 137336 286288
rect 137296 267734 137324 286282
rect 137204 267706 137324 267734
rect 135902 265160 135958 265169
rect 135902 265095 135958 265104
rect 135260 260228 135312 260234
rect 135260 260170 135312 260176
rect 135916 259978 135944 265095
rect 137204 263974 137232 267706
rect 137836 267028 137888 267034
rect 137836 266970 137888 266976
rect 137192 263968 137244 263974
rect 137192 263910 137244 263916
rect 136226 260228 136278 260234
rect 136226 260170 136278 260176
rect 133156 259950 133492 259978
rect 133984 259964 134044 259978
rect 133984 259950 134058 259964
rect 134260 259950 134596 259978
rect 134812 259950 135148 259978
rect 135700 259950 135944 259978
rect 136238 259964 136266 260170
rect 137204 259978 137232 263910
rect 137848 263809 137876 266970
rect 137834 263800 137890 263809
rect 137834 263735 137890 263744
rect 137468 263560 137520 263566
rect 137468 263502 137520 263508
rect 137480 261089 137508 263502
rect 137466 261080 137522 261089
rect 137466 261015 137522 261024
rect 136804 259950 137232 259978
rect 124862 259720 124918 259729
rect 127254 259720 127310 259729
rect 124918 259678 125212 259706
rect 124862 259655 124918 259664
rect 134030 259706 134058 259950
rect 137480 259842 137508 261015
rect 137356 259814 137508 259842
rect 137848 259842 137876 263735
rect 138676 262585 138704 430578
rect 138756 418192 138808 418198
rect 138756 418134 138808 418140
rect 138768 265033 138796 418134
rect 138754 265024 138810 265033
rect 138754 264959 138810 264968
rect 138662 262576 138718 262585
rect 138662 262511 138718 262520
rect 138676 259978 138704 262511
rect 138460 259950 138704 259978
rect 138768 259978 138796 264959
rect 138768 259950 139012 259978
rect 137848 259814 137908 259842
rect 134030 259692 134380 259706
rect 134044 259690 134380 259692
rect 134044 259684 134392 259690
rect 134044 259678 134340 259684
rect 127254 259655 127310 259664
rect 134340 259626 134392 259632
rect 123298 259584 123354 259593
rect 123004 259542 123298 259570
rect 123298 259519 123354 259528
rect 123772 259542 124108 259570
rect 123772 259457 123800 259542
rect 139412 259486 139440 484366
rect 140044 470620 140096 470626
rect 140044 470562 140096 470568
rect 140056 267734 140084 470562
rect 140780 280832 140832 280838
rect 140780 280774 140832 280780
rect 140056 267706 140360 267734
rect 139492 264308 139544 264314
rect 139492 264250 139544 264256
rect 139504 259978 139532 264250
rect 140332 262721 140360 267706
rect 140318 262712 140374 262721
rect 140318 262647 140374 262656
rect 140332 259978 140360 262647
rect 140792 260137 140820 280774
rect 141700 265736 141752 265742
rect 141700 265678 141752 265684
rect 141712 264042 141740 265678
rect 141148 264036 141200 264042
rect 141148 263978 141200 263984
rect 141700 264036 141752 264042
rect 141700 263978 141752 263984
rect 140778 260128 140834 260137
rect 140778 260063 140834 260072
rect 141160 259978 141188 263978
rect 141744 260128 141800 260137
rect 141744 260063 141800 260072
rect 139504 259950 139564 259978
rect 140332 259950 140668 259978
rect 141160 259950 141220 259978
rect 141758 259964 141786 260063
rect 142172 259962 142200 590650
rect 142804 563100 142856 563106
rect 142804 563042 142856 563048
rect 142816 267734 142844 563042
rect 142896 524476 142948 524482
rect 142896 524418 142948 524424
rect 142632 267706 142844 267734
rect 142632 263906 142660 267706
rect 142620 263900 142672 263906
rect 142620 263842 142672 263848
rect 142250 262984 142306 262993
rect 142250 262919 142306 262928
rect 142264 259978 142292 262919
rect 142632 259978 142660 263842
rect 142908 262993 142936 524418
rect 142894 262984 142950 262993
rect 142894 262919 142950 262928
rect 143644 260273 143672 616830
rect 144184 576904 144236 576910
rect 144184 576846 144236 576852
rect 144196 262546 144224 576846
rect 145564 287700 145616 287706
rect 145564 287642 145616 287648
rect 145104 282192 145156 282198
rect 145104 282134 145156 282140
rect 144184 262540 144236 262546
rect 144184 262482 144236 262488
rect 143630 260264 143686 260273
rect 143630 260199 143686 260208
rect 144196 259978 144224 262482
rect 144504 260264 144560 260273
rect 145116 260250 145144 282134
rect 145576 263673 145604 287642
rect 146208 268456 146260 268462
rect 146208 268398 146260 268404
rect 146220 263770 146248 268398
rect 146208 263764 146260 263770
rect 146208 263706 146260 263712
rect 145286 263664 145342 263673
rect 145286 263599 145342 263608
rect 145562 263664 145618 263673
rect 145562 263599 145618 263608
rect 144504 260199 144560 260208
rect 145070 260222 145144 260250
rect 142160 259956 142212 259962
rect 142264 259950 142324 259978
rect 142632 259950 142876 259978
rect 143092 259962 143428 259978
rect 143080 259956 143428 259962
rect 142160 259898 142212 259904
rect 143132 259950 143428 259956
rect 143980 259950 144224 259978
rect 144518 259964 144546 260199
rect 143080 259898 143132 259904
rect 144918 259856 144974 259865
rect 145070 259842 145098 260222
rect 145300 259978 145328 263599
rect 146220 260250 146248 263706
rect 146174 260222 146248 260250
rect 145300 259950 145636 259978
rect 146174 259964 146202 260222
rect 146312 259978 146340 696934
rect 146944 683188 146996 683194
rect 146944 683130 146996 683136
rect 146956 262857 146984 683130
rect 147956 283620 148008 283626
rect 147956 283562 148008 283568
rect 147772 269816 147824 269822
rect 147772 269758 147824 269764
rect 146942 262848 146998 262857
rect 146942 262783 146998 262792
rect 146956 259978 146984 262783
rect 147678 259992 147734 260001
rect 146312 259950 146740 259978
rect 146956 259950 147292 259978
rect 146312 259894 146340 259950
rect 147784 259978 147812 269758
rect 147968 259978 147996 283562
rect 148336 267734 148364 700266
rect 149060 660340 149112 660346
rect 149060 660282 149112 660288
rect 148336 267706 148548 267734
rect 148520 263838 148548 267706
rect 148508 263832 148560 263838
rect 148508 263774 148560 263780
rect 148520 259978 148548 263774
rect 149072 260273 149100 660282
rect 150440 284368 150492 284374
rect 150440 284310 150492 284316
rect 149152 271176 149204 271182
rect 149152 271118 149204 271124
rect 149058 260264 149114 260273
rect 149058 260199 149114 260208
rect 149164 259978 149192 271118
rect 150452 263498 150480 284310
rect 151820 274712 151872 274718
rect 151820 274654 151872 274660
rect 151084 273964 151136 273970
rect 151084 273906 151136 273912
rect 151096 263702 151124 273906
rect 151832 267734 151860 274654
rect 151832 267706 152412 267734
rect 152188 264988 152240 264994
rect 152188 264930 152240 264936
rect 151084 263696 151136 263702
rect 151084 263638 151136 263644
rect 150440 263492 150492 263498
rect 150440 263434 150492 263440
rect 150898 262848 150954 262857
rect 150898 262783 150954 262792
rect 150024 260264 150080 260273
rect 150024 260199 150080 260208
rect 147734 259950 147844 259978
rect 147968 259950 148396 259978
rect 148520 259950 148948 259978
rect 149164 259950 149500 259978
rect 150038 259964 150066 260199
rect 150912 259978 150940 262783
rect 150604 259950 150940 259978
rect 151096 259978 151124 263638
rect 151360 263492 151412 263498
rect 151360 263434 151412 263440
rect 151372 259978 151400 263434
rect 152200 259978 152228 264930
rect 152384 259978 152412 267706
rect 153120 264994 153148 700334
rect 153108 264988 153160 264994
rect 153108 264930 153160 264936
rect 153212 262682 153240 702406
rect 157340 700868 157392 700874
rect 157340 700810 157392 700816
rect 155960 700800 156012 700806
rect 155960 700742 156012 700748
rect 154580 700664 154632 700670
rect 154580 700606 154632 700612
rect 153292 700460 153344 700466
rect 153292 700402 153344 700408
rect 153200 262676 153252 262682
rect 153200 262618 153252 262624
rect 153304 259978 153332 700402
rect 153384 276072 153436 276078
rect 153384 276014 153436 276020
rect 153396 267734 153424 276014
rect 153396 267706 154068 267734
rect 153842 262576 153898 262585
rect 153842 262511 153898 262520
rect 153856 259978 153884 262511
rect 154040 259978 154068 267706
rect 154592 259978 154620 700606
rect 155866 262440 155922 262449
rect 155866 262375 155922 262384
rect 155880 259978 155908 262375
rect 155972 260273 156000 700742
rect 156050 277536 156106 277545
rect 156050 277471 156106 277480
rect 155958 260264 156014 260273
rect 155958 260199 156014 260208
rect 151096 259950 151156 259978
rect 151372 259950 151708 259978
rect 152200 259950 152260 259978
rect 152384 259950 152812 259978
rect 153304 259950 153364 259978
rect 153856 259950 153916 259978
rect 154040 259950 154468 259978
rect 154592 259964 155020 259978
rect 154592 259950 155034 259964
rect 155572 259950 155908 259978
rect 156064 259978 156092 277471
rect 157156 262608 157208 262614
rect 157156 262550 157208 262556
rect 156648 260264 156704 260273
rect 156648 260199 156704 260208
rect 156064 259950 156124 259978
rect 147678 259927 147734 259936
rect 144974 259828 145098 259842
rect 146300 259888 146352 259894
rect 146300 259830 146352 259836
rect 144974 259814 145084 259828
rect 144918 259791 144974 259800
rect 148152 259729 148180 259950
rect 149164 259826 149192 259950
rect 153304 259842 153332 259950
rect 149152 259820 149204 259826
rect 149152 259762 149204 259768
rect 153212 259814 153332 259842
rect 153212 259758 153240 259814
rect 153200 259752 153252 259758
rect 148138 259720 148194 259729
rect 153200 259694 153252 259700
rect 155006 259706 155034 259950
rect 156662 259842 156690 260199
rect 157168 259978 157196 262550
rect 157352 260234 157380 700810
rect 160744 700732 160796 700738
rect 160744 700674 160796 700680
rect 157432 447840 157484 447846
rect 157432 447782 157484 447788
rect 157340 260228 157392 260234
rect 157340 260170 157392 260176
rect 157444 259978 157472 447782
rect 160100 279472 160152 279478
rect 160100 279414 160152 279420
rect 158720 269136 158772 269142
rect 158720 269078 158772 269084
rect 158732 267734 158760 269078
rect 158732 267706 159588 267734
rect 159088 263628 159140 263634
rect 159088 263570 159140 263576
rect 158720 262676 158772 262682
rect 158720 262618 158772 262624
rect 158732 260953 158760 262618
rect 158718 260944 158774 260953
rect 158718 260879 158774 260888
rect 158306 260228 158358 260234
rect 158306 260170 158358 260176
rect 158318 259978 158346 260170
rect 158732 259978 158760 260879
rect 159100 259978 159128 263570
rect 159560 259978 159588 267706
rect 160112 260273 160140 279414
rect 160756 262546 160784 700674
rect 162216 700596 162268 700602
rect 162216 700538 162268 700544
rect 162124 700528 162176 700534
rect 162124 700470 162176 700476
rect 162136 267734 162164 700470
rect 162044 267706 162164 267734
rect 162044 262750 162072 267706
rect 162032 262744 162084 262750
rect 162032 262686 162084 262692
rect 160744 262540 160796 262546
rect 160744 262482 160796 262488
rect 160098 260264 160154 260273
rect 160098 260199 160154 260208
rect 160756 259978 160784 262482
rect 161064 260264 161120 260273
rect 161064 260199 161120 260208
rect 157168 259950 157228 259978
rect 157444 259950 158116 259978
rect 158318 259964 158668 259978
rect 158332 259950 158668 259964
rect 158732 259950 158884 259978
rect 159100 259950 159436 259978
rect 159560 259950 159988 259978
rect 160540 259950 160784 259978
rect 161078 259978 161106 260199
rect 161202 259992 161258 260001
rect 161078 259964 161202 259978
rect 161092 259950 161202 259964
rect 156878 259856 156934 259865
rect 156662 259828 156878 259842
rect 156676 259814 156878 259828
rect 158088 259826 158116 259950
rect 156878 259791 156934 259800
rect 158076 259820 158128 259826
rect 158076 259762 158128 259768
rect 158640 259758 158668 259950
rect 162044 259978 162072 262686
rect 162228 262682 162256 700538
rect 162308 683256 162360 683262
rect 162308 683198 162360 683204
rect 162320 265266 162348 683198
rect 163504 670744 163556 670750
rect 163504 670686 163556 670692
rect 162308 265260 162360 265266
rect 162308 265202 162360 265208
rect 162216 262676 162268 262682
rect 162216 262618 162268 262624
rect 162228 260250 162256 262618
rect 161644 259950 162072 259978
rect 162182 260222 162256 260250
rect 162182 259964 162210 260222
rect 162320 259978 162348 265202
rect 163516 265033 163544 670686
rect 163596 656940 163648 656946
rect 163596 656882 163648 656888
rect 163502 265024 163558 265033
rect 163502 264959 163558 264968
rect 163412 263288 163464 263294
rect 163412 263230 163464 263236
rect 163424 262818 163452 263230
rect 163412 262812 163464 262818
rect 163412 262754 163464 262760
rect 163424 259978 163452 262754
rect 162320 259950 162748 259978
rect 163300 259950 163452 259978
rect 163516 259978 163544 264959
rect 163608 263294 163636 656882
rect 164240 632120 164292 632126
rect 164240 632062 164292 632068
rect 163596 263288 163648 263294
rect 163596 263230 163648 263236
rect 164252 259978 164280 632062
rect 164884 618316 164936 618322
rect 164884 618258 164936 618264
rect 164896 265062 164924 618258
rect 164976 605872 165028 605878
rect 164976 605814 165028 605820
rect 164884 265056 164936 265062
rect 164884 264998 164936 265004
rect 164988 262721 165016 605814
rect 165620 579692 165672 579698
rect 165620 579634 165672 579640
rect 165344 265056 165396 265062
rect 165344 264998 165396 265004
rect 164974 262712 165030 262721
rect 164974 262647 165030 262656
rect 164988 260250 165016 262647
rect 164942 260222 165016 260250
rect 163516 259950 163852 259978
rect 164252 259950 164648 259978
rect 164942 259964 164970 260222
rect 165356 259978 165384 264998
rect 165632 259978 165660 579634
rect 167644 565888 167696 565894
rect 167644 565830 167696 565836
rect 166264 553444 166316 553450
rect 166264 553386 166316 553392
rect 166276 265169 166304 553386
rect 167000 527196 167052 527202
rect 167000 527138 167052 527144
rect 166262 265160 166318 265169
rect 166262 265095 166318 265104
rect 166032 260128 166088 260137
rect 166032 260063 166088 260072
rect 166046 259978 166074 260063
rect 165356 259950 165508 259978
rect 165632 259964 166074 259978
rect 166276 259978 166304 265095
rect 167012 260234 167040 527138
rect 167656 267734 167684 565830
rect 167736 501016 167788 501022
rect 167736 500958 167788 500964
rect 167472 267706 167684 267734
rect 167748 267734 167776 500958
rect 169772 447846 169800 702406
rect 202800 700806 202828 703520
rect 202788 700800 202840 700806
rect 202788 700742 202840 700748
rect 185584 670744 185636 670750
rect 185584 670686 185636 670692
rect 184204 643136 184256 643142
rect 184204 643078 184256 643084
rect 178684 536852 178736 536858
rect 178684 536794 178736 536800
rect 170404 462392 170456 462398
rect 170404 462334 170456 462340
rect 169760 447840 169812 447846
rect 169760 447782 169812 447788
rect 169760 422340 169812 422346
rect 169760 422282 169812 422288
rect 169024 274032 169076 274038
rect 169024 273974 169076 273980
rect 169036 267734 169064 273974
rect 167748 267706 167868 267734
rect 169036 267706 169156 267734
rect 167472 265130 167500 267706
rect 167840 265334 167868 267706
rect 167828 265328 167880 265334
rect 167828 265270 167880 265276
rect 167460 265124 167512 265130
rect 167460 265066 167512 265072
rect 167000 260228 167052 260234
rect 167000 260170 167052 260176
rect 167472 259978 167500 265066
rect 167690 260228 167742 260234
rect 167690 260170 167742 260176
rect 165632 259950 166060 259964
rect 166276 259950 166612 259978
rect 167164 259950 167500 259978
rect 167702 259964 167730 260170
rect 167840 259978 167868 265270
rect 169128 265198 169156 267706
rect 169208 265668 169260 265674
rect 169208 265610 169260 265616
rect 169116 265192 169168 265198
rect 169116 265134 169168 265140
rect 169128 259978 169156 265134
rect 167840 259950 168268 259978
rect 168820 259950 169156 259978
rect 169220 259978 169248 265610
rect 169772 260234 169800 422282
rect 170416 265470 170444 462334
rect 170496 448588 170548 448594
rect 170496 448530 170548 448536
rect 170404 265464 170456 265470
rect 170404 265406 170456 265412
rect 170508 263090 170536 448530
rect 171784 409896 171836 409902
rect 171784 409838 171836 409844
rect 171140 397520 171192 397526
rect 171140 397462 171192 397468
rect 170680 265464 170732 265470
rect 170680 265406 170732 265412
rect 170220 263084 170272 263090
rect 170220 263026 170272 263032
rect 170496 263084 170548 263090
rect 170496 263026 170548 263032
rect 169760 260228 169812 260234
rect 169760 260170 169812 260176
rect 170232 259978 170260 263026
rect 170692 259978 170720 265406
rect 171002 260228 171054 260234
rect 171002 260170 171054 260176
rect 171014 260098 171042 260170
rect 171002 260092 171054 260098
rect 171002 260034 171054 260040
rect 169220 259950 169524 259978
rect 169924 259950 170260 259978
rect 170476 259950 170720 259978
rect 171014 259964 171042 260034
rect 171152 259978 171180 397462
rect 171796 265402 171824 409838
rect 173900 318844 173952 318850
rect 173900 318786 173952 318792
rect 173164 289128 173216 289134
rect 173164 289070 173216 289076
rect 172704 268388 172756 268394
rect 172704 268330 172756 268336
rect 171784 265396 171836 265402
rect 171784 265338 171836 265344
rect 171796 259978 171824 265338
rect 172716 263702 172744 268330
rect 172704 263696 172756 263702
rect 172704 263638 172756 263644
rect 172716 260250 172744 263638
rect 173176 263634 173204 289070
rect 173256 271244 173308 271250
rect 173256 271186 173308 271192
rect 173268 265606 173296 271186
rect 173256 265600 173308 265606
rect 173256 265542 173308 265548
rect 173164 263628 173216 263634
rect 173164 263570 173216 263576
rect 173268 260250 173296 265542
rect 173716 263628 173768 263634
rect 173716 263570 173768 263576
rect 172670 260222 172744 260250
rect 173222 260222 173296 260250
rect 171152 259962 171732 259978
rect 171152 259956 171744 259962
rect 171152 259950 171692 259956
rect 161202 259927 161258 259936
rect 158628 259752 158680 259758
rect 155222 259720 155278 259729
rect 155006 259692 155222 259706
rect 155020 259678 155222 259692
rect 148138 259655 148194 259664
rect 158628 259694 158680 259700
rect 155222 259655 155278 259664
rect 164620 259593 164648 259950
rect 169496 259894 169524 259950
rect 171796 259950 172132 259978
rect 172670 259964 172698 260222
rect 173222 259964 173250 260222
rect 173728 259978 173756 263570
rect 173912 260438 173940 318786
rect 175924 305040 175976 305046
rect 175924 304982 175976 304988
rect 174544 292596 174596 292602
rect 174544 292538 174596 292544
rect 174556 265810 174584 292538
rect 175936 267734 175964 304982
rect 178696 280838 178724 536794
rect 181444 510672 181496 510678
rect 181444 510614 181496 510620
rect 180064 456816 180116 456822
rect 180064 456758 180116 456764
rect 178684 280832 178736 280838
rect 178684 280774 178736 280780
rect 175844 267706 175964 267734
rect 174544 265804 174596 265810
rect 174544 265746 174596 265752
rect 173900 260432 173952 260438
rect 173900 260374 173952 260380
rect 173912 259978 173940 260374
rect 174556 259978 174584 265746
rect 175844 265538 175872 267706
rect 175924 266416 175976 266422
rect 175924 266358 175976 266364
rect 175832 265532 175884 265538
rect 175832 265474 175884 265480
rect 175844 259978 175872 265474
rect 175936 260302 175964 266358
rect 180076 264246 180104 456758
rect 181456 265742 181484 510614
rect 182824 378208 182876 378214
rect 182824 378150 182876 378156
rect 182836 286346 182864 378150
rect 182824 286340 182876 286346
rect 182824 286282 182876 286288
rect 184216 282198 184244 643078
rect 184204 282192 184256 282198
rect 184204 282134 184256 282140
rect 185596 268462 185624 670686
rect 203524 630692 203576 630698
rect 203524 630634 203576 630640
rect 199384 404388 199436 404394
rect 199384 404330 199436 404336
rect 186320 284980 186372 284986
rect 186320 284922 186372 284928
rect 187148 284980 187200 284986
rect 187148 284922 187200 284928
rect 186332 284374 186360 284922
rect 186320 284368 186372 284374
rect 186320 284310 186372 284316
rect 185584 268456 185636 268462
rect 185584 268398 185636 268404
rect 181444 265736 181496 265742
rect 181444 265678 181496 265684
rect 180064 264240 180116 264246
rect 180064 264182 180116 264188
rect 178500 262948 178552 262954
rect 178500 262890 178552 262896
rect 179236 262948 179288 262954
rect 179236 262890 179288 262896
rect 176752 262472 176804 262478
rect 176752 262414 176804 262420
rect 176764 261390 176792 262414
rect 176752 261384 176804 261390
rect 176752 261326 176804 261332
rect 176200 260976 176252 260982
rect 176200 260918 176252 260924
rect 175924 260296 175976 260302
rect 175924 260238 175976 260244
rect 173728 259950 173788 259978
rect 173912 259950 174340 259978
rect 174556 259950 174892 259978
rect 175444 259950 175872 259978
rect 175936 259978 175964 260238
rect 176108 260228 176160 260234
rect 176108 260170 176160 260176
rect 175936 259950 175996 259978
rect 171692 259898 171744 259904
rect 176120 259894 176148 260170
rect 176212 259978 176240 260918
rect 176764 259978 176792 261326
rect 178512 261118 178540 262890
rect 178500 261112 178552 261118
rect 178500 261054 178552 261060
rect 177580 260908 177632 260914
rect 177580 260850 177632 260856
rect 176212 259950 176548 259978
rect 176764 259950 177100 259978
rect 169484 259888 169536 259894
rect 169484 259830 169536 259836
rect 176108 259888 176160 259894
rect 176108 259830 176160 259836
rect 164606 259584 164662 259593
rect 139780 259542 140116 259570
rect 139780 259486 139808 259542
rect 177592 259570 177620 260850
rect 178408 260296 178460 260302
rect 178408 260238 178460 260244
rect 178040 259616 178092 259622
rect 177316 259554 177652 259570
rect 178420 259570 178448 260238
rect 178512 259978 178540 261054
rect 179248 259978 179276 262890
rect 180156 262472 180208 262478
rect 180156 262414 180208 262420
rect 180168 259978 180196 262414
rect 182916 262404 182968 262410
rect 182916 262346 182968 262352
rect 181260 262268 181312 262274
rect 181260 262210 181312 262216
rect 180524 261180 180576 261186
rect 180524 261122 180576 261128
rect 180536 259978 180564 261122
rect 181272 259978 181300 262210
rect 181996 261044 182048 261050
rect 181996 260986 182048 260992
rect 178512 259950 178756 259978
rect 179248 259950 179308 259978
rect 179860 259950 180196 259978
rect 180412 259950 180564 259978
rect 180964 259950 181300 259978
rect 182008 259978 182036 260986
rect 182928 259978 182956 262346
rect 184572 262336 184624 262342
rect 184572 262278 184624 262284
rect 184020 261248 184072 261254
rect 184020 261190 184072 261196
rect 184032 259978 184060 261190
rect 184584 259978 184612 262278
rect 185584 260432 185636 260438
rect 185584 260374 185636 260380
rect 185596 260098 185624 260374
rect 185584 260092 185636 260098
rect 185584 260034 185636 260040
rect 185676 260092 185728 260098
rect 185676 260034 185728 260040
rect 182008 259950 182068 259978
rect 182620 259950 182956 259978
rect 183724 259950 184060 259978
rect 184276 259950 184612 259978
rect 185688 259894 185716 260034
rect 185676 259888 185728 259894
rect 185676 259830 185728 259836
rect 181812 259616 181864 259622
rect 178092 259564 178448 259570
rect 178040 259558 178448 259564
rect 164606 259519 164662 259528
rect 177304 259548 177652 259554
rect 177356 259542 177652 259548
rect 178052 259542 178448 259558
rect 181516 259564 181812 259570
rect 181516 259558 181864 259564
rect 181516 259542 181852 259558
rect 183172 259554 183508 259570
rect 183172 259548 183520 259554
rect 183172 259542 183468 259548
rect 177304 259490 177356 259496
rect 185380 259542 185716 259570
rect 183468 259490 183520 259496
rect 139400 259480 139452 259486
rect 123758 259448 123814 259457
rect 139400 259422 139452 259428
rect 139768 259480 139820 259486
rect 184940 259480 184992 259486
rect 139768 259422 139820 259428
rect 184828 259428 184940 259434
rect 185688 259457 185716 259542
rect 184828 259422 184992 259428
rect 185674 259448 185730 259457
rect 184828 259406 184980 259422
rect 123758 259383 123814 259392
rect 185674 259383 185730 259392
rect 130844 200728 130896 200734
rect 129002 200696 129058 200705
rect 130844 200670 130896 200676
rect 132040 200728 132092 200734
rect 132040 200670 132092 200676
rect 132132 200728 132184 200734
rect 132132 200670 132184 200676
rect 132224 200728 132276 200734
rect 184204 200728 184256 200734
rect 132224 200670 132276 200676
rect 178222 200696 178278 200705
rect 129002 200631 129058 200640
rect 124862 200560 124918 200569
rect 124862 200495 124918 200504
rect 124034 200152 124090 200161
rect 124034 200087 124090 200096
rect 123944 192704 123996 192710
rect 123944 192646 123996 192652
rect 123668 150952 123720 150958
rect 123668 150894 123720 150900
rect 122838 150512 122894 150521
rect 122838 150447 122894 150456
rect 122564 145988 122616 145994
rect 122564 145930 122616 145936
rect 122852 140060 122880 150447
rect 123484 147552 123536 147558
rect 123484 147494 123536 147500
rect 123496 141982 123524 147494
rect 123484 141976 123536 141982
rect 123484 141918 123536 141924
rect 122852 140032 123156 140060
rect 123128 139890 123156 140032
rect 123128 139862 123556 139890
rect 123680 139398 123708 150894
rect 123024 139392 123076 139398
rect 123022 139360 123024 139369
rect 123668 139392 123720 139398
rect 123076 139360 123078 139369
rect 123956 139369 123984 192646
rect 124048 147694 124076 200087
rect 124770 197568 124826 197577
rect 124770 197503 124826 197512
rect 124784 194342 124812 197503
rect 124772 194336 124824 194342
rect 124772 194278 124824 194284
rect 124036 147688 124088 147694
rect 124036 147630 124088 147636
rect 124048 139890 124076 147630
rect 124770 144800 124826 144809
rect 124770 144735 124826 144744
rect 124784 143585 124812 144735
rect 124770 143576 124826 143585
rect 124770 143511 124826 143520
rect 124784 139890 124812 143511
rect 124876 141658 124904 200495
rect 126060 199776 126112 199782
rect 126060 199718 126112 199724
rect 125046 198792 125102 198801
rect 125046 198727 125102 198736
rect 124954 197296 125010 197305
rect 124954 197231 125010 197240
rect 124968 142154 124996 197231
rect 125060 144809 125088 198727
rect 125876 198688 125928 198694
rect 125876 198630 125928 198636
rect 125140 197532 125192 197538
rect 125140 197474 125192 197480
rect 125152 193905 125180 197474
rect 125138 193896 125194 193905
rect 125138 193831 125194 193840
rect 125888 192817 125916 198630
rect 126072 198121 126100 199718
rect 126612 199436 126664 199442
rect 126612 199378 126664 199384
rect 127900 199436 127952 199442
rect 127900 199378 127952 199384
rect 126334 199336 126390 199345
rect 126334 199271 126390 199280
rect 126058 198112 126114 198121
rect 126058 198047 126114 198056
rect 126244 194744 126296 194750
rect 126244 194686 126296 194692
rect 125874 192808 125930 192817
rect 125874 192743 125930 192752
rect 125324 190324 125376 190330
rect 125324 190266 125376 190272
rect 125336 151814 125364 190266
rect 125336 151786 125548 151814
rect 125046 144800 125102 144809
rect 125046 144735 125102 144744
rect 124968 142126 125088 142154
rect 124876 141630 124996 141658
rect 124864 141568 124916 141574
rect 124864 141510 124916 141516
rect 124048 139862 124108 139890
rect 124660 139862 124812 139890
rect 124876 139890 124904 141510
rect 124968 140049 124996 141630
rect 124954 140040 125010 140049
rect 125060 140010 125088 142126
rect 124954 139975 125010 139984
rect 125048 140004 125100 140010
rect 125048 139946 125100 139952
rect 124876 139862 125212 139890
rect 125520 139369 125548 151786
rect 125690 143304 125746 143313
rect 125690 143239 125746 143248
rect 125704 139482 125732 143239
rect 126150 142080 126206 142089
rect 126150 142015 126206 142024
rect 126164 140865 126192 142015
rect 126150 140856 126206 140865
rect 126150 140791 126206 140800
rect 126164 139890 126192 140791
rect 126256 140758 126284 194686
rect 126244 140752 126296 140758
rect 126244 140694 126296 140700
rect 126348 140593 126376 199271
rect 126428 198892 126480 198898
rect 126428 198834 126480 198840
rect 126334 140584 126390 140593
rect 126334 140519 126390 140528
rect 126440 140418 126468 198834
rect 126520 198008 126572 198014
rect 126520 197950 126572 197956
rect 126428 140412 126480 140418
rect 126428 140354 126480 140360
rect 126532 140078 126560 197950
rect 126624 146878 126652 199378
rect 127622 198520 127678 198529
rect 127622 198455 127678 198464
rect 126704 195220 126756 195226
rect 126704 195162 126756 195168
rect 126612 146872 126664 146878
rect 126612 146814 126664 146820
rect 126716 140622 126744 195162
rect 126796 147620 126848 147626
rect 126796 147562 126848 147568
rect 126808 141273 126836 147562
rect 126888 146872 126940 146878
rect 126888 146814 126940 146820
rect 126794 141264 126850 141273
rect 126794 141199 126850 141208
rect 126794 140992 126850 141001
rect 126900 140978 126928 146814
rect 127348 141908 127400 141914
rect 127348 141850 127400 141856
rect 126850 140950 126928 140978
rect 126794 140927 126850 140936
rect 126704 140616 126756 140622
rect 126704 140558 126756 140564
rect 126520 140072 126572 140078
rect 126520 140014 126572 140020
rect 126808 139890 126836 140927
rect 127360 140826 127388 141850
rect 127348 140820 127400 140826
rect 127348 140762 127400 140768
rect 127360 139890 127388 140762
rect 127636 140486 127664 198455
rect 127716 197872 127768 197878
rect 127716 197814 127768 197820
rect 127728 143206 127756 197814
rect 127808 197804 127860 197810
rect 127808 197746 127860 197752
rect 127820 145382 127848 197746
rect 127912 194478 127940 199378
rect 127900 194472 127952 194478
rect 127900 194414 127952 194420
rect 128636 148368 128688 148374
rect 128636 148310 128688 148316
rect 127808 145376 127860 145382
rect 127808 145318 127860 145324
rect 128544 143404 128596 143410
rect 128544 143346 128596 143352
rect 127716 143200 127768 143206
rect 127716 143142 127768 143148
rect 128266 143168 128322 143177
rect 128266 143103 128322 143112
rect 128280 142526 128308 143103
rect 128268 142520 128320 142526
rect 128268 142462 128320 142468
rect 127808 142044 127860 142050
rect 127808 141986 127860 141992
rect 127820 141710 127848 141986
rect 127808 141704 127860 141710
rect 127808 141646 127860 141652
rect 127624 140480 127676 140486
rect 127624 140422 127676 140428
rect 128280 139890 128308 142462
rect 128556 142458 128584 143346
rect 128544 142452 128596 142458
rect 128544 142394 128596 142400
rect 128556 140162 128584 142394
rect 126164 139862 126316 139890
rect 126808 139862 126868 139890
rect 127360 139862 127420 139890
rect 127972 139862 128308 139890
rect 128510 140134 128584 140162
rect 128510 139876 128538 140134
rect 128648 139890 128676 148310
rect 128912 141976 128964 141982
rect 128912 141918 128964 141924
rect 128924 140049 128952 141918
rect 129016 140457 129044 200631
rect 130856 200122 130884 200670
rect 131120 200660 131172 200666
rect 131120 200602 131172 200608
rect 130934 200152 130990 200161
rect 130844 200116 130896 200122
rect 130934 200087 130990 200096
rect 130844 200058 130896 200064
rect 130752 199708 130804 199714
rect 130752 199650 130804 199656
rect 130660 199640 130712 199646
rect 130660 199582 130712 199588
rect 129186 199200 129242 199209
rect 129186 199135 129242 199144
rect 129096 198756 129148 198762
rect 129096 198698 129148 198704
rect 129002 140448 129058 140457
rect 129002 140383 129058 140392
rect 129108 140282 129136 198698
rect 129200 140554 129228 199135
rect 129280 198552 129332 198558
rect 129280 198494 129332 198500
rect 129292 141982 129320 198494
rect 130672 198393 130700 199582
rect 130764 198694 130792 199650
rect 130752 198688 130804 198694
rect 130752 198630 130804 198636
rect 130658 198384 130714 198393
rect 130658 198319 130714 198328
rect 130660 197736 130712 197742
rect 130660 197678 130712 197684
rect 129464 196580 129516 196586
rect 129464 196522 129516 196528
rect 129372 196376 129424 196382
rect 129372 196318 129424 196324
rect 129280 141976 129332 141982
rect 129280 141918 129332 141924
rect 129280 141840 129332 141846
rect 129280 141782 129332 141788
rect 129188 140548 129240 140554
rect 129188 140490 129240 140496
rect 129096 140276 129148 140282
rect 129096 140218 129148 140224
rect 128910 140040 128966 140049
rect 128910 139975 128966 139984
rect 129292 139890 129320 141782
rect 129384 140350 129412 196318
rect 129372 140344 129424 140350
rect 129476 140321 129504 196522
rect 129740 196172 129792 196178
rect 129740 196114 129792 196120
rect 129752 193118 129780 196114
rect 130384 195152 130436 195158
rect 130384 195094 130436 195100
rect 129740 193112 129792 193118
rect 129740 193054 129792 193060
rect 129832 146260 129884 146266
rect 129832 146202 129884 146208
rect 129740 145512 129792 145518
rect 129740 145454 129792 145460
rect 129752 143206 129780 145454
rect 129844 143410 129872 146202
rect 129924 146056 129976 146062
rect 129924 145998 129976 146004
rect 129832 143404 129884 143410
rect 129832 143346 129884 143352
rect 129740 143200 129792 143206
rect 129740 143142 129792 143148
rect 129936 142254 129964 145998
rect 130200 144220 130252 144226
rect 130200 144162 130252 144168
rect 129924 142248 129976 142254
rect 129924 142190 129976 142196
rect 129372 140286 129424 140292
rect 129462 140312 129518 140321
rect 129462 140247 129518 140256
rect 130212 140162 130240 144162
rect 130166 140134 130240 140162
rect 128648 139862 129076 139890
rect 129292 139862 129628 139890
rect 130166 139876 130194 140134
rect 130396 140049 130424 195094
rect 130568 193180 130620 193186
rect 130568 193122 130620 193128
rect 130474 193080 130530 193089
rect 130474 193015 130530 193024
rect 130488 141953 130516 193015
rect 130474 141944 130530 141953
rect 130474 141879 130530 141888
rect 130382 140040 130438 140049
rect 130382 139975 130438 139984
rect 129476 139738 129504 139862
rect 129464 139732 129516 139738
rect 129464 139674 129516 139680
rect 125704 139466 126100 139482
rect 125704 139460 126112 139466
rect 125704 139454 126060 139460
rect 126060 139402 126112 139408
rect 130580 139369 130608 193122
rect 130672 164898 130700 197678
rect 130948 193050 130976 200087
rect 131132 194750 131160 200602
rect 132052 200598 132080 200670
rect 132040 200592 132092 200598
rect 132040 200534 132092 200540
rect 132144 200326 132172 200670
rect 132236 200598 132264 200670
rect 177764 200660 177816 200666
rect 184204 200670 184256 200676
rect 178222 200631 178278 200640
rect 180064 200660 180116 200666
rect 177764 200602 177816 200608
rect 132224 200592 132276 200598
rect 132224 200534 132276 200540
rect 177776 200326 177804 200602
rect 178040 200592 178092 200598
rect 178040 200534 178092 200540
rect 178132 200592 178184 200598
rect 178132 200534 178184 200540
rect 177948 200524 178000 200530
rect 177948 200466 178000 200472
rect 132132 200320 132184 200326
rect 132132 200262 132184 200268
rect 177764 200320 177816 200326
rect 177764 200262 177816 200268
rect 177856 200252 177908 200258
rect 177856 200194 177908 200200
rect 132052 200110 132388 200138
rect 131856 197668 131908 197674
rect 131856 197610 131908 197616
rect 131764 196444 131816 196450
rect 131764 196386 131816 196392
rect 131120 194744 131172 194750
rect 131120 194686 131172 194692
rect 130936 193044 130988 193050
rect 130936 192986 130988 192992
rect 130844 192432 130896 192438
rect 130844 192374 130896 192380
rect 130660 164892 130712 164898
rect 130660 164834 130712 164840
rect 130660 145444 130712 145450
rect 130660 145386 130712 145392
rect 130672 139890 130700 145386
rect 130672 139862 130732 139890
rect 130856 139369 130884 192374
rect 131776 147490 131804 196386
rect 131868 148102 131896 197610
rect 132052 195265 132080 200110
rect 132466 199866 132494 200124
rect 132420 199838 132494 199866
rect 132132 199300 132184 199306
rect 132132 199242 132184 199248
rect 132144 196042 132172 199242
rect 132314 198656 132370 198665
rect 132314 198591 132370 198600
rect 132132 196036 132184 196042
rect 132132 195978 132184 195984
rect 132038 195256 132094 195265
rect 132038 195191 132094 195200
rect 131948 194880 132000 194886
rect 131948 194822 132000 194828
rect 131856 148096 131908 148102
rect 131856 148038 131908 148044
rect 131764 147484 131816 147490
rect 131764 147426 131816 147432
rect 131960 147422 131988 194822
rect 132328 190454 132356 198591
rect 132420 198490 132448 199838
rect 132558 199628 132586 200124
rect 132650 199730 132678 200124
rect 132742 199923 132770 200124
rect 132728 199914 132784 199923
rect 132728 199849 132784 199858
rect 132834 199730 132862 200124
rect 132926 199918 132954 200124
rect 133018 199918 133046 200124
rect 132914 199912 132966 199918
rect 132914 199854 132966 199860
rect 133006 199912 133058 199918
rect 133006 199854 133058 199860
rect 133110 199764 133138 200124
rect 132650 199702 132724 199730
rect 132558 199600 132632 199628
rect 132500 198688 132552 198694
rect 132500 198630 132552 198636
rect 132408 198484 132460 198490
rect 132408 198426 132460 198432
rect 132512 198014 132540 198630
rect 132604 198257 132632 199600
rect 132590 198248 132646 198257
rect 132590 198183 132646 198192
rect 132500 198008 132552 198014
rect 132500 197950 132552 197956
rect 132696 195673 132724 199702
rect 132788 199702 132862 199730
rect 133064 199736 133138 199764
rect 132788 199306 132816 199702
rect 132960 199572 133012 199578
rect 132960 199514 133012 199520
rect 132972 199306 133000 199514
rect 132776 199300 132828 199306
rect 132776 199242 132828 199248
rect 132960 199300 133012 199306
rect 132960 199242 133012 199248
rect 132868 197464 132920 197470
rect 132868 197406 132920 197412
rect 132776 196512 132828 196518
rect 132776 196454 132828 196460
rect 132682 195664 132738 195673
rect 132682 195599 132738 195608
rect 132592 195492 132644 195498
rect 132592 195434 132644 195440
rect 132684 195492 132736 195498
rect 132684 195434 132736 195440
rect 132604 194818 132632 195434
rect 132592 194812 132644 194818
rect 132592 194754 132644 194760
rect 132328 190426 132448 190454
rect 131948 147416 132000 147422
rect 131948 147358 132000 147364
rect 131672 146192 131724 146198
rect 131672 146134 131724 146140
rect 131120 146124 131172 146130
rect 131120 146066 131172 146072
rect 131132 142186 131160 146066
rect 131212 144288 131264 144294
rect 131212 144230 131264 144236
rect 131120 142180 131172 142186
rect 131120 142122 131172 142128
rect 131224 139890 131252 144230
rect 131488 143336 131540 143342
rect 131488 143278 131540 143284
rect 131500 139890 131528 143278
rect 131684 140060 131712 146134
rect 132420 140162 132448 190426
rect 132696 151774 132724 195434
rect 132788 187270 132816 196454
rect 132880 191214 132908 197406
rect 132960 196988 133012 196994
rect 132960 196930 133012 196936
rect 132972 196246 133000 196930
rect 132960 196240 133012 196246
rect 132960 196182 133012 196188
rect 133064 195974 133092 199736
rect 133202 199696 133230 200124
rect 133294 199918 133322 200124
rect 133282 199912 133334 199918
rect 133282 199854 133334 199860
rect 133386 199764 133414 200124
rect 133478 199918 133506 200124
rect 133466 199912 133518 199918
rect 133466 199854 133518 199860
rect 133570 199764 133598 200124
rect 133662 199918 133690 200124
rect 133754 199918 133782 200124
rect 133650 199912 133702 199918
rect 133650 199854 133702 199860
rect 133742 199912 133794 199918
rect 133846 199889 133874 200124
rect 133938 199918 133966 200124
rect 133926 199912 133978 199918
rect 133742 199854 133794 199860
rect 133832 199880 133888 199889
rect 133926 199854 133978 199860
rect 134030 199850 134058 200124
rect 134122 199923 134150 200124
rect 134108 199914 134164 199923
rect 134214 199918 134242 200124
rect 133832 199815 133888 199824
rect 134018 199844 134070 199850
rect 134108 199849 134164 199858
rect 134202 199912 134254 199918
rect 134202 199854 134254 199860
rect 133340 199736 133414 199764
rect 133524 199736 133598 199764
rect 133648 199778 133704 199787
rect 134018 199786 134070 199792
rect 133202 199668 133276 199696
rect 133248 197354 133276 199668
rect 133340 197538 133368 199736
rect 133420 199640 133472 199646
rect 133420 199582 133472 199588
rect 133328 197532 133380 197538
rect 133328 197474 133380 197480
rect 133248 197326 133368 197354
rect 133236 196784 133288 196790
rect 133236 196726 133288 196732
rect 133248 196314 133276 196726
rect 133236 196308 133288 196314
rect 133236 196250 133288 196256
rect 133144 196036 133196 196042
rect 133144 195978 133196 195984
rect 132972 195946 133092 195974
rect 132868 191208 132920 191214
rect 132868 191150 132920 191156
rect 132776 187264 132828 187270
rect 132776 187206 132828 187212
rect 132684 151768 132736 151774
rect 132684 151710 132736 151716
rect 132972 148578 133000 195946
rect 133050 195256 133106 195265
rect 133050 195191 133106 195200
rect 133064 151570 133092 195191
rect 133156 187134 133184 195978
rect 133340 192642 133368 197326
rect 133432 195498 133460 199582
rect 133524 197470 133552 199736
rect 133648 199713 133704 199722
rect 133880 199776 133932 199782
rect 134306 199764 134334 200124
rect 134398 199923 134426 200124
rect 134384 199914 134440 199923
rect 134490 199918 134518 200124
rect 134582 199923 134610 200124
rect 134384 199849 134440 199858
rect 134478 199912 134530 199918
rect 134478 199854 134530 199860
rect 134568 199914 134624 199923
rect 134568 199849 134624 199858
rect 133880 199718 133932 199724
rect 134062 199744 134118 199753
rect 133788 199708 133840 199714
rect 133788 199650 133840 199656
rect 133604 199640 133656 199646
rect 133604 199582 133656 199588
rect 133512 197464 133564 197470
rect 133512 197406 133564 197412
rect 133420 195492 133472 195498
rect 133420 195434 133472 195440
rect 133616 192953 133644 199582
rect 133696 199572 133748 199578
rect 133696 199514 133748 199520
rect 133708 199306 133736 199514
rect 133696 199300 133748 199306
rect 133696 199242 133748 199248
rect 133800 196518 133828 199650
rect 133892 198098 133920 199718
rect 134260 199736 134334 199764
rect 134522 199744 134578 199753
rect 134062 199679 134118 199688
rect 134156 199708 134208 199714
rect 133892 198070 134012 198098
rect 133880 197940 133932 197946
rect 133880 197882 133932 197888
rect 133892 197742 133920 197882
rect 133880 197736 133932 197742
rect 133880 197678 133932 197684
rect 133984 196602 134012 198070
rect 134076 196761 134104 199679
rect 134156 199650 134208 199656
rect 134168 197402 134196 199650
rect 134260 197470 134288 199736
rect 134432 199708 134484 199714
rect 134522 199679 134578 199688
rect 134432 199650 134484 199656
rect 134248 197464 134300 197470
rect 134444 197441 134472 199650
rect 134248 197406 134300 197412
rect 134430 197432 134486 197441
rect 134156 197396 134208 197402
rect 134430 197367 134486 197376
rect 134156 197338 134208 197344
rect 134536 196874 134564 199679
rect 134674 199560 134702 200124
rect 134766 199918 134794 200124
rect 134858 199923 134886 200124
rect 134754 199912 134806 199918
rect 134754 199854 134806 199860
rect 134844 199914 134900 199923
rect 134844 199849 134900 199858
rect 134950 199764 134978 200124
rect 135042 199918 135070 200124
rect 135134 199918 135162 200124
rect 135226 199918 135254 200124
rect 135318 199918 135346 200124
rect 135410 199918 135438 200124
rect 135030 199912 135082 199918
rect 135030 199854 135082 199860
rect 135122 199912 135174 199918
rect 135122 199854 135174 199860
rect 135214 199912 135266 199918
rect 135214 199854 135266 199860
rect 135306 199912 135358 199918
rect 135306 199854 135358 199860
rect 135398 199912 135450 199918
rect 135502 199889 135530 200124
rect 135398 199854 135450 199860
rect 135488 199880 135544 199889
rect 135488 199815 135544 199824
rect 134904 199736 134978 199764
rect 135076 199776 135128 199782
rect 134800 199708 134852 199714
rect 134800 199650 134852 199656
rect 134674 199532 134748 199560
rect 134616 197396 134668 197402
rect 134616 197338 134668 197344
rect 134444 196846 134564 196874
rect 134062 196752 134118 196761
rect 134062 196687 134118 196696
rect 133984 196574 134288 196602
rect 133788 196512 133840 196518
rect 133788 196454 133840 196460
rect 134156 196512 134208 196518
rect 134156 196454 134208 196460
rect 133602 192944 133658 192953
rect 133602 192879 133658 192888
rect 133328 192636 133380 192642
rect 133328 192578 133380 192584
rect 133144 187128 133196 187134
rect 133144 187070 133196 187076
rect 133052 151564 133104 151570
rect 133052 151506 133104 151512
rect 134168 151298 134196 196454
rect 134260 186998 134288 196574
rect 134338 195936 134394 195945
rect 134338 195871 134394 195880
rect 134248 186992 134300 186998
rect 134248 186934 134300 186940
rect 134352 151706 134380 195871
rect 134340 151700 134392 151706
rect 134340 151642 134392 151648
rect 134444 151638 134472 196846
rect 134524 196036 134576 196042
rect 134524 195978 134576 195984
rect 134536 187202 134564 195978
rect 134628 193214 134656 197338
rect 134720 196178 134748 199532
rect 134708 196172 134760 196178
rect 134708 196114 134760 196120
rect 134628 193186 134748 193214
rect 134524 187196 134576 187202
rect 134524 187138 134576 187144
rect 134720 180794 134748 193186
rect 134812 192953 134840 199650
rect 134904 194410 134932 199736
rect 135490 199776 135542 199782
rect 135364 199753 135490 199764
rect 135076 199718 135128 199724
rect 135350 199744 135490 199753
rect 134984 199640 135036 199646
rect 134984 199582 135036 199588
rect 134996 196042 135024 199582
rect 135088 196518 135116 199718
rect 135406 199736 135490 199744
rect 135594 199764 135622 200124
rect 135686 199889 135714 200124
rect 135778 199918 135806 200124
rect 135870 199923 135898 200124
rect 135766 199912 135818 199918
rect 135672 199880 135728 199889
rect 135766 199854 135818 199860
rect 135856 199914 135912 199923
rect 135856 199849 135912 199858
rect 135672 199815 135728 199824
rect 135962 199764 135990 200124
rect 136054 199918 136082 200124
rect 136146 199918 136174 200124
rect 136238 199923 136266 200124
rect 136042 199912 136094 199918
rect 136042 199854 136094 199860
rect 136134 199912 136186 199918
rect 136134 199854 136186 199860
rect 136224 199914 136280 199923
rect 136224 199849 136280 199858
rect 136330 199850 136358 200124
rect 136422 199923 136450 200124
rect 136408 199914 136464 199923
rect 136318 199844 136370 199850
rect 136408 199849 136464 199858
rect 136318 199786 136370 199792
rect 136088 199776 136140 199782
rect 135594 199736 135668 199764
rect 135490 199718 135542 199724
rect 135350 199679 135406 199688
rect 135168 199640 135220 199646
rect 135168 199582 135220 199588
rect 135306 199640 135358 199646
rect 135306 199582 135358 199588
rect 135444 199640 135496 199646
rect 135640 199594 135668 199736
rect 135718 199744 135774 199753
rect 135962 199736 136036 199764
rect 135718 199679 135774 199688
rect 135444 199582 135496 199588
rect 135180 199442 135208 199582
rect 135168 199436 135220 199442
rect 135168 199378 135220 199384
rect 135318 199322 135346 199582
rect 135180 199294 135346 199322
rect 135180 197713 135208 199294
rect 135456 198734 135484 199582
rect 135548 199566 135668 199594
rect 135548 198914 135576 199566
rect 135732 199458 135760 199679
rect 135732 199430 135944 199458
rect 135812 199368 135864 199374
rect 135732 199316 135812 199322
rect 135732 199310 135864 199316
rect 135732 199294 135852 199310
rect 135732 199073 135760 199294
rect 135718 199064 135774 199073
rect 135718 198999 135774 199008
rect 135548 198886 135760 198914
rect 135456 198706 135668 198734
rect 135166 197704 135222 197713
rect 135166 197639 135222 197648
rect 135168 197464 135220 197470
rect 135168 197406 135220 197412
rect 135076 196512 135128 196518
rect 135076 196454 135128 196460
rect 134984 196036 135036 196042
rect 134984 195978 135036 195984
rect 135180 194594 135208 197406
rect 135536 195084 135588 195090
rect 135536 195026 135588 195032
rect 135444 194880 135496 194886
rect 135444 194822 135496 194828
rect 135088 194566 135208 194594
rect 134892 194404 134944 194410
rect 134892 194346 134944 194352
rect 134798 192944 134854 192953
rect 134798 192879 134854 192888
rect 135088 187066 135116 194566
rect 135352 194472 135404 194478
rect 135352 194414 135404 194420
rect 135364 189854 135392 194414
rect 135456 190194 135484 194822
rect 135444 190188 135496 190194
rect 135444 190130 135496 190136
rect 135352 189848 135404 189854
rect 135352 189790 135404 189796
rect 135076 187060 135128 187066
rect 135076 187002 135128 187008
rect 134628 180766 134748 180794
rect 134432 151632 134484 151638
rect 134432 151574 134484 151580
rect 134628 151502 134656 180766
rect 134616 151496 134668 151502
rect 134616 151438 134668 151444
rect 135548 151366 135576 195026
rect 135640 151434 135668 198706
rect 135732 195974 135760 198886
rect 135916 196738 135944 199430
rect 136008 196874 136036 199736
rect 136514 199764 136542 200124
rect 136606 199918 136634 200124
rect 136698 199918 136726 200124
rect 136790 199918 136818 200124
rect 136882 199923 136910 200124
rect 136594 199912 136646 199918
rect 136594 199854 136646 199860
rect 136686 199912 136738 199918
rect 136686 199854 136738 199860
rect 136778 199912 136830 199918
rect 136778 199854 136830 199860
rect 136868 199914 136924 199923
rect 136868 199849 136924 199858
rect 136088 199718 136140 199724
rect 136178 199744 136234 199753
rect 136100 198354 136128 199718
rect 136362 199744 136418 199753
rect 136234 199702 136312 199730
rect 136178 199679 136234 199688
rect 136180 199640 136232 199646
rect 136180 199582 136232 199588
rect 136088 198348 136140 198354
rect 136088 198290 136140 198296
rect 136008 196846 136128 196874
rect 135916 196710 136036 196738
rect 135732 195946 135944 195974
rect 135812 195492 135864 195498
rect 135812 195434 135864 195440
rect 135720 195016 135772 195022
rect 135720 194958 135772 194964
rect 135628 151428 135680 151434
rect 135628 151370 135680 151376
rect 135536 151360 135588 151366
rect 135536 151302 135588 151308
rect 134156 151292 134208 151298
rect 134156 151234 134208 151240
rect 132960 148572 133012 148578
rect 132960 148514 133012 148520
rect 135732 148510 135760 194958
rect 135824 148617 135852 195434
rect 135916 187338 135944 195946
rect 135904 187332 135956 187338
rect 135904 187274 135956 187280
rect 136008 151026 136036 196710
rect 136100 195090 136128 196846
rect 136088 195084 136140 195090
rect 136088 195026 136140 195032
rect 136192 194478 136220 199582
rect 136284 195498 136312 199702
rect 136362 199679 136418 199688
rect 136468 199736 136542 199764
rect 136732 199776 136784 199782
rect 136272 195492 136324 195498
rect 136272 195434 136324 195440
rect 136376 194886 136404 199679
rect 136468 195022 136496 199736
rect 136974 199730 137002 200124
rect 136732 199718 136784 199724
rect 136640 199708 136692 199714
rect 136640 199650 136692 199656
rect 136548 199640 136600 199646
rect 136548 199582 136600 199588
rect 136560 197033 136588 199582
rect 136652 197354 136680 199650
rect 136744 197674 136772 199718
rect 136928 199702 137002 199730
rect 136824 199572 136876 199578
rect 136824 199514 136876 199520
rect 136836 198393 136864 199514
rect 136822 198384 136878 198393
rect 136822 198319 136878 198328
rect 136732 197668 136784 197674
rect 136732 197610 136784 197616
rect 136652 197326 136772 197354
rect 136546 197024 136602 197033
rect 136546 196959 136602 196968
rect 136744 195090 136772 197326
rect 136732 195084 136784 195090
rect 136732 195026 136784 195032
rect 136456 195016 136508 195022
rect 136456 194958 136508 194964
rect 136364 194880 136416 194886
rect 136364 194822 136416 194828
rect 136180 194472 136232 194478
rect 136180 194414 136232 194420
rect 136928 189990 136956 199702
rect 137066 199628 137094 200124
rect 137158 199753 137186 200124
rect 137250 199918 137278 200124
rect 137342 199918 137370 200124
rect 137434 199923 137462 200124
rect 137238 199912 137290 199918
rect 137238 199854 137290 199860
rect 137330 199912 137382 199918
rect 137330 199854 137382 199860
rect 137420 199914 137476 199923
rect 137420 199849 137476 199858
rect 137526 199850 137554 200124
rect 137618 199850 137646 200124
rect 137514 199844 137566 199850
rect 137514 199786 137566 199792
rect 137606 199844 137658 199850
rect 137606 199786 137658 199792
rect 137710 199764 137738 200124
rect 137802 199918 137830 200124
rect 137894 199918 137922 200124
rect 137986 199918 138014 200124
rect 138078 199918 138106 200124
rect 137790 199912 137842 199918
rect 137790 199854 137842 199860
rect 137882 199912 137934 199918
rect 137882 199854 137934 199860
rect 137974 199912 138026 199918
rect 137974 199854 138026 199860
rect 138066 199912 138118 199918
rect 138066 199854 138118 199860
rect 137928 199776 137980 199782
rect 137710 199753 137784 199764
rect 137144 199744 137200 199753
rect 137710 199744 137798 199753
rect 137710 199736 137742 199744
rect 137144 199679 137200 199688
rect 137928 199718 137980 199724
rect 138020 199776 138072 199782
rect 138170 199764 138198 200124
rect 138262 199918 138290 200124
rect 138250 199912 138302 199918
rect 138250 199854 138302 199860
rect 138354 199764 138382 200124
rect 138446 199850 138474 200124
rect 138538 199918 138566 200124
rect 138526 199912 138578 199918
rect 138630 199889 138658 200124
rect 138722 199918 138750 200124
rect 138814 199918 138842 200124
rect 138906 199918 138934 200124
rect 138710 199912 138762 199918
rect 138526 199854 138578 199860
rect 138616 199880 138672 199889
rect 138434 199844 138486 199850
rect 138710 199854 138762 199860
rect 138802 199912 138854 199918
rect 138802 199854 138854 199860
rect 138894 199912 138946 199918
rect 138894 199854 138946 199860
rect 138616 199815 138672 199824
rect 138434 199786 138486 199792
rect 138170 199736 138244 199764
rect 138020 199718 138072 199724
rect 137742 199679 137798 199688
rect 137192 199640 137244 199646
rect 137066 199600 137140 199628
rect 137006 199064 137062 199073
rect 137006 198999 137062 199008
rect 137020 198218 137048 198999
rect 137008 198212 137060 198218
rect 137008 198154 137060 198160
rect 137112 198121 137140 199600
rect 137560 199640 137612 199646
rect 137192 199582 137244 199588
rect 137466 199608 137522 199617
rect 137098 198112 137154 198121
rect 137098 198047 137154 198056
rect 137008 192160 137060 192166
rect 137008 192102 137060 192108
rect 136916 189984 136968 189990
rect 136916 189926 136968 189932
rect 135996 151020 136048 151026
rect 135996 150962 136048 150968
rect 135810 148608 135866 148617
rect 135810 148543 135866 148552
rect 135720 148504 135772 148510
rect 135720 148446 135772 148452
rect 137020 147393 137048 192102
rect 137204 189922 137232 199582
rect 137284 199572 137336 199578
rect 137560 199582 137612 199588
rect 137652 199640 137704 199646
rect 137652 199582 137704 199588
rect 137744 199640 137796 199646
rect 137744 199582 137796 199588
rect 137834 199608 137890 199617
rect 137466 199543 137522 199552
rect 137284 199514 137336 199520
rect 137296 196761 137324 199514
rect 137480 197062 137508 199543
rect 137468 197056 137520 197062
rect 137468 196998 137520 197004
rect 137282 196752 137338 196761
rect 137282 196687 137338 196696
rect 137284 196512 137336 196518
rect 137284 196454 137336 196460
rect 137192 189916 137244 189922
rect 137192 189858 137244 189864
rect 137296 187513 137324 196454
rect 137468 195084 137520 195090
rect 137468 195026 137520 195032
rect 137480 190262 137508 195026
rect 137572 191282 137600 199582
rect 137664 197606 137692 199582
rect 137652 197600 137704 197606
rect 137652 197542 137704 197548
rect 137756 191418 137784 199582
rect 137834 199543 137836 199552
rect 137888 199543 137890 199552
rect 137836 199514 137888 199520
rect 137940 192166 137968 199718
rect 138032 195809 138060 199718
rect 138112 199640 138164 199646
rect 138112 199582 138164 199588
rect 138018 195800 138074 195809
rect 138018 195735 138074 195744
rect 138124 195265 138152 199582
rect 138110 195256 138166 195265
rect 138110 195191 138166 195200
rect 138216 194392 138244 199736
rect 138308 199736 138382 199764
rect 138756 199776 138808 199782
rect 138754 199744 138756 199753
rect 138998 199764 139026 200124
rect 138808 199744 138810 199753
rect 138308 198121 138336 199736
rect 138952 199736 139026 199764
rect 139090 199764 139118 200124
rect 139182 199918 139210 200124
rect 139170 199912 139222 199918
rect 139170 199854 139222 199860
rect 139274 199764 139302 200124
rect 139366 199918 139394 200124
rect 139354 199912 139406 199918
rect 139354 199854 139406 199860
rect 139458 199764 139486 200124
rect 139550 199918 139578 200124
rect 139642 199923 139670 200124
rect 139538 199912 139590 199918
rect 139538 199854 139590 199860
rect 139628 199914 139684 199923
rect 139734 199918 139762 200124
rect 139826 199918 139854 200124
rect 139918 199918 139946 200124
rect 140010 199918 140038 200124
rect 139628 199849 139684 199858
rect 139722 199912 139774 199918
rect 139722 199854 139774 199860
rect 139814 199912 139866 199918
rect 139814 199854 139866 199860
rect 139906 199912 139958 199918
rect 139906 199854 139958 199860
rect 139998 199912 140050 199918
rect 139998 199854 140050 199860
rect 139090 199736 139164 199764
rect 138754 199679 138810 199688
rect 138848 199708 138900 199714
rect 138848 199650 138900 199656
rect 138480 199640 138532 199646
rect 138480 199582 138532 199588
rect 138388 199572 138440 199578
rect 138388 199514 138440 199520
rect 138294 198112 138350 198121
rect 138294 198047 138350 198056
rect 138400 195242 138428 199514
rect 138492 196897 138520 199582
rect 138664 199572 138716 199578
rect 138664 199514 138716 199520
rect 138756 199572 138808 199578
rect 138756 199514 138808 199520
rect 138478 196888 138534 196897
rect 138478 196823 138534 196832
rect 138400 195214 138612 195242
rect 138216 194364 138428 194392
rect 137928 192160 137980 192166
rect 137928 192102 137980 192108
rect 137744 191412 137796 191418
rect 137744 191354 137796 191360
rect 137560 191276 137612 191282
rect 137560 191218 137612 191224
rect 138296 191140 138348 191146
rect 138296 191082 138348 191088
rect 137468 190256 137520 190262
rect 137468 190198 137520 190204
rect 137282 187504 137338 187513
rect 137282 187439 137338 187448
rect 137006 147384 137062 147393
rect 137006 147319 137062 147328
rect 138308 147257 138336 191082
rect 138400 150958 138428 194364
rect 138388 150952 138440 150958
rect 138388 150894 138440 150900
rect 138294 147248 138350 147257
rect 138584 147218 138612 195214
rect 138294 147183 138350 147192
rect 138572 147212 138624 147218
rect 138572 147154 138624 147160
rect 138676 147082 138704 199514
rect 138768 196654 138796 199514
rect 138756 196648 138808 196654
rect 138756 196590 138808 196596
rect 138860 195129 138888 199650
rect 138846 195120 138902 195129
rect 138846 195055 138902 195064
rect 138952 180794 138980 199736
rect 139032 199640 139084 199646
rect 139032 199582 139084 199588
rect 139044 194002 139072 199582
rect 139136 194818 139164 199736
rect 139228 199736 139302 199764
rect 139412 199736 139486 199764
rect 139676 199776 139728 199782
rect 139674 199744 139676 199753
rect 139860 199776 139912 199782
rect 139728 199744 139730 199753
rect 139124 194812 139176 194818
rect 139124 194754 139176 194760
rect 139032 193996 139084 194002
rect 139032 193938 139084 193944
rect 139228 191146 139256 199736
rect 139308 199640 139360 199646
rect 139308 199582 139360 199588
rect 139320 194954 139348 199582
rect 139412 196518 139440 199736
rect 139584 199708 139636 199714
rect 139860 199718 139912 199724
rect 139952 199776 140004 199782
rect 140102 199764 140130 200124
rect 140194 199918 140222 200124
rect 140286 199923 140314 200124
rect 140182 199912 140234 199918
rect 140182 199854 140234 199860
rect 140272 199914 140328 199923
rect 140378 199918 140406 200124
rect 140470 199918 140498 200124
rect 140272 199849 140328 199858
rect 140366 199912 140418 199918
rect 140366 199854 140418 199860
rect 140458 199912 140510 199918
rect 140458 199854 140510 199860
rect 140412 199776 140464 199782
rect 140102 199736 140176 199764
rect 139952 199718 140004 199724
rect 139674 199679 139730 199688
rect 139584 199650 139636 199656
rect 139492 199300 139544 199306
rect 139492 199242 139544 199248
rect 139504 198830 139532 199242
rect 139492 198824 139544 198830
rect 139492 198766 139544 198772
rect 139400 196512 139452 196518
rect 139400 196454 139452 196460
rect 139308 194948 139360 194954
rect 139308 194890 139360 194896
rect 139596 193214 139624 199650
rect 139674 199200 139730 199209
rect 139674 199135 139730 199144
rect 139688 196450 139716 199135
rect 139872 196761 139900 199718
rect 139858 196752 139914 196761
rect 139858 196687 139914 196696
rect 139676 196444 139728 196450
rect 139676 196386 139728 196392
rect 139596 193186 139716 193214
rect 139216 191140 139268 191146
rect 139216 191082 139268 191088
rect 138860 180766 138980 180794
rect 138664 147076 138716 147082
rect 138664 147018 138716 147024
rect 138860 146946 138888 180766
rect 139688 151065 139716 193186
rect 139964 191264 139992 199718
rect 140044 199640 140096 199646
rect 140044 199582 140096 199588
rect 140056 194274 140084 199582
rect 140044 194268 140096 194274
rect 140044 194210 140096 194216
rect 139872 191236 139992 191264
rect 139872 190330 139900 191236
rect 139952 191140 140004 191146
rect 139952 191082 140004 191088
rect 139860 190324 139912 190330
rect 139860 190266 139912 190272
rect 139674 151056 139730 151065
rect 139674 150991 139730 151000
rect 138848 146940 138900 146946
rect 138848 146882 138900 146888
rect 133880 144696 133932 144702
rect 133880 144638 133932 144644
rect 135902 144664 135958 144673
rect 133144 143268 133196 143274
rect 133144 143210 133196 143216
rect 132592 142248 132644 142254
rect 132592 142190 132644 142196
rect 132420 140134 132540 140162
rect 132512 140078 132540 140134
rect 132500 140072 132552 140078
rect 131684 140032 131988 140060
rect 131960 139890 131988 140032
rect 132500 140014 132552 140020
rect 132604 139890 132632 142190
rect 133156 139890 133184 143210
rect 133512 142452 133564 142458
rect 133512 142394 133564 142400
rect 133524 142254 133552 142394
rect 133512 142248 133564 142254
rect 133512 142190 133564 142196
rect 133892 139890 133920 144638
rect 135902 144599 135958 144608
rect 135444 143404 135496 143410
rect 135444 143346 135496 143352
rect 134248 142180 134300 142186
rect 134248 142122 134300 142128
rect 134260 139890 134288 142122
rect 134800 141772 134852 141778
rect 134800 141714 134852 141720
rect 134812 139890 134840 141714
rect 135456 139890 135484 143346
rect 135916 139890 135944 144599
rect 138662 144528 138718 144537
rect 138662 144463 138718 144472
rect 137558 144392 137614 144401
rect 137558 144327 137614 144336
rect 137008 143200 137060 143206
rect 137008 143142 137060 143148
rect 136640 141704 136692 141710
rect 136640 141646 136692 141652
rect 136652 139890 136680 141646
rect 137020 139890 137048 143142
rect 137572 139890 137600 144327
rect 138110 143984 138166 143993
rect 138110 143919 138166 143928
rect 138124 139890 138152 143919
rect 138676 139890 138704 144463
rect 139768 143132 139820 143138
rect 139768 143074 139820 143080
rect 139398 141808 139454 141817
rect 139398 141743 139454 141752
rect 139412 139890 139440 141743
rect 139780 139890 139808 143074
rect 139964 140185 139992 191082
rect 140148 147626 140176 199736
rect 140562 199764 140590 200124
rect 140654 199923 140682 200124
rect 140640 199914 140696 199923
rect 140746 199918 140774 200124
rect 140838 199918 140866 200124
rect 140930 199923 140958 200124
rect 140640 199849 140696 199858
rect 140734 199912 140786 199918
rect 140734 199854 140786 199860
rect 140826 199912 140878 199918
rect 140826 199854 140878 199860
rect 140916 199914 140972 199923
rect 141022 199918 141050 200124
rect 141114 199923 141142 200124
rect 140916 199849 140972 199858
rect 141010 199912 141062 199918
rect 141010 199854 141062 199860
rect 141100 199914 141156 199923
rect 141100 199849 141156 199858
rect 140412 199718 140464 199724
rect 140516 199736 140590 199764
rect 140734 199776 140786 199782
rect 140228 199572 140280 199578
rect 140228 199514 140280 199520
rect 140240 193214 140268 199514
rect 140424 194070 140452 199718
rect 140412 194064 140464 194070
rect 140412 194006 140464 194012
rect 140240 193186 140360 193214
rect 140136 147620 140188 147626
rect 140136 147562 140188 147568
rect 140332 147558 140360 193186
rect 140516 187474 140544 199736
rect 140654 199724 140734 199730
rect 141206 199764 141234 200124
rect 141298 199918 141326 200124
rect 141390 199923 141418 200124
rect 141286 199912 141338 199918
rect 141286 199854 141338 199860
rect 141376 199914 141432 199923
rect 141482 199918 141510 200124
rect 141574 199923 141602 200124
rect 141376 199849 141432 199858
rect 141470 199912 141522 199918
rect 141470 199854 141522 199860
rect 141560 199914 141616 199923
rect 141560 199849 141616 199858
rect 141666 199764 141694 200124
rect 141758 199918 141786 200124
rect 141850 199923 141878 200124
rect 141746 199912 141798 199918
rect 141746 199854 141798 199860
rect 141836 199914 141892 199923
rect 141836 199849 141892 199858
rect 141942 199850 141970 200124
rect 142034 199918 142062 200124
rect 142126 199923 142154 200124
rect 142022 199912 142074 199918
rect 142022 199854 142074 199860
rect 142112 199914 142168 199923
rect 142218 199918 142246 200124
rect 142310 199923 142338 200124
rect 141930 199844 141982 199850
rect 142112 199849 142168 199858
rect 142206 199912 142258 199918
rect 142206 199854 142258 199860
rect 142296 199914 142352 199923
rect 142296 199849 142352 199858
rect 141930 199786 141982 199792
rect 142402 199764 142430 200124
rect 142494 199923 142522 200124
rect 142480 199914 142536 199923
rect 142586 199918 142614 200124
rect 142678 199918 142706 200124
rect 142770 199918 142798 200124
rect 142862 199923 142890 200124
rect 142480 199849 142536 199858
rect 142574 199912 142626 199918
rect 142574 199854 142626 199860
rect 142666 199912 142718 199918
rect 142666 199854 142718 199860
rect 142758 199912 142810 199918
rect 142758 199854 142810 199860
rect 142848 199914 142904 199923
rect 142954 199918 142982 200124
rect 143046 199923 143074 200124
rect 142848 199849 142904 199858
rect 142942 199912 142994 199918
rect 142942 199854 142994 199860
rect 143032 199914 143088 199923
rect 143138 199918 143166 200124
rect 143032 199849 143088 199858
rect 143126 199912 143178 199918
rect 143126 199854 143178 199860
rect 143230 199850 143258 200124
rect 143322 199850 143350 200124
rect 143414 199850 143442 200124
rect 143218 199844 143270 199850
rect 143218 199786 143270 199792
rect 143310 199844 143362 199850
rect 143310 199786 143362 199792
rect 143402 199844 143454 199850
rect 143402 199786 143454 199792
rect 140654 199718 140786 199724
rect 140962 199744 141018 199753
rect 140654 199702 140774 199718
rect 140872 199708 140924 199714
rect 140654 199594 140682 199702
rect 141160 199736 141234 199764
rect 141620 199753 141694 199764
rect 141330 199744 141386 199753
rect 141160 199730 141188 199736
rect 140962 199679 141018 199688
rect 141068 199702 141188 199730
rect 140872 199650 140924 199656
rect 140608 199566 140682 199594
rect 140778 199608 140834 199617
rect 140608 192914 140636 199566
rect 140778 199543 140834 199552
rect 140792 194594 140820 199543
rect 140884 197577 140912 199650
rect 140870 197568 140926 197577
rect 140870 197503 140926 197512
rect 140872 196988 140924 196994
rect 140872 196930 140924 196936
rect 140700 194566 140820 194594
rect 140596 192908 140648 192914
rect 140596 192850 140648 192856
rect 140700 191146 140728 194566
rect 140884 191214 140912 196930
rect 140976 194594 141004 199679
rect 141068 196704 141096 199702
rect 141606 199744 141694 199753
rect 141330 199679 141386 199688
rect 141424 199708 141476 199714
rect 141238 199608 141294 199617
rect 141148 199572 141200 199578
rect 141238 199543 141294 199552
rect 141148 199514 141200 199520
rect 141160 199209 141188 199514
rect 141146 199200 141202 199209
rect 141146 199135 141202 199144
rect 141148 198824 141200 198830
rect 141148 198766 141200 198772
rect 141160 196994 141188 198766
rect 141148 196988 141200 196994
rect 141148 196930 141200 196936
rect 141068 196676 141188 196704
rect 140976 194566 141096 194594
rect 140872 191208 140924 191214
rect 140872 191150 140924 191156
rect 140688 191140 140740 191146
rect 140688 191082 140740 191088
rect 140504 187468 140556 187474
rect 140504 187410 140556 187416
rect 141068 148442 141096 194566
rect 141160 151094 141188 196676
rect 141252 191350 141280 199543
rect 141344 193934 141372 199679
rect 141662 199736 141694 199744
rect 141882 199744 141938 199753
rect 141804 199702 141882 199730
rect 141804 199696 141832 199702
rect 141606 199679 141662 199688
rect 141424 199650 141476 199656
rect 141712 199668 141832 199696
rect 141882 199679 141938 199688
rect 142066 199744 142122 199753
rect 142356 199736 142430 199764
rect 142482 199776 142534 199782
rect 142480 199744 142482 199753
rect 142534 199744 142536 199753
rect 142066 199679 142122 199688
rect 142160 199708 142212 199714
rect 141332 193928 141384 193934
rect 141332 193870 141384 193876
rect 141436 193214 141464 199650
rect 141608 199640 141660 199646
rect 141606 199608 141608 199617
rect 141660 199608 141662 199617
rect 141516 199572 141568 199578
rect 141606 199543 141662 199552
rect 141516 199514 141568 199520
rect 141528 199458 141556 199514
rect 141712 199458 141740 199668
rect 141884 199640 141936 199646
rect 141884 199582 141936 199588
rect 141976 199640 142028 199646
rect 141976 199582 142028 199588
rect 141792 199572 141844 199578
rect 141792 199514 141844 199520
rect 141528 199430 141740 199458
rect 141514 199200 141570 199209
rect 141514 199135 141570 199144
rect 141698 199200 141754 199209
rect 141698 199135 141754 199144
rect 141528 196761 141556 199135
rect 141712 198830 141740 199135
rect 141700 198824 141752 198830
rect 141700 198766 141752 198772
rect 141514 196752 141570 196761
rect 141514 196687 141570 196696
rect 141436 193186 141740 193214
rect 141240 191344 141292 191350
rect 141240 191286 141292 191292
rect 141332 191140 141384 191146
rect 141332 191082 141384 191088
rect 141148 151088 141200 151094
rect 141148 151030 141200 151036
rect 141056 148436 141108 148442
rect 141056 148378 141108 148384
rect 140320 147552 140372 147558
rect 140320 147494 140372 147500
rect 141344 147354 141372 191082
rect 141332 147348 141384 147354
rect 141332 147290 141384 147296
rect 141712 147150 141740 193186
rect 141804 186314 141832 199514
rect 141896 198665 141924 199582
rect 141882 198656 141938 198665
rect 141882 198591 141938 198600
rect 141884 196648 141936 196654
rect 141884 196590 141936 196596
rect 141896 187406 141924 196590
rect 141988 191146 142016 199582
rect 142080 198082 142108 199679
rect 142212 199668 142292 199696
rect 142160 199650 142212 199656
rect 142160 199368 142212 199374
rect 142160 199310 142212 199316
rect 142172 199209 142200 199310
rect 142158 199200 142214 199209
rect 142158 199135 142214 199144
rect 142068 198076 142120 198082
rect 142068 198018 142120 198024
rect 142264 196654 142292 199668
rect 142356 199102 142384 199736
rect 142480 199679 142536 199688
rect 142894 199744 142950 199753
rect 143400 199744 143456 199753
rect 142894 199679 142950 199688
rect 143080 199708 143132 199714
rect 142528 199640 142580 199646
rect 142528 199582 142580 199588
rect 142712 199640 142764 199646
rect 142712 199582 142764 199588
rect 142436 199504 142488 199510
rect 142436 199446 142488 199452
rect 142344 199096 142396 199102
rect 142344 199038 142396 199044
rect 142448 198490 142476 199446
rect 142540 199374 142568 199582
rect 142620 199572 142672 199578
rect 142620 199514 142672 199520
rect 142528 199368 142580 199374
rect 142528 199310 142580 199316
rect 142526 198520 142582 198529
rect 142436 198484 142488 198490
rect 142526 198455 142582 198464
rect 142436 198426 142488 198432
rect 142252 196648 142304 196654
rect 142252 196590 142304 196596
rect 142436 191548 142488 191554
rect 142436 191490 142488 191496
rect 141976 191140 142028 191146
rect 141976 191082 142028 191088
rect 141884 187400 141936 187406
rect 141884 187342 141936 187348
rect 141804 186286 141924 186314
rect 141700 147144 141752 147150
rect 141700 147086 141752 147092
rect 141896 147014 141924 186286
rect 142448 148986 142476 191490
rect 142540 191282 142568 198455
rect 142632 192506 142660 199514
rect 142620 192500 142672 192506
rect 142620 192442 142672 192448
rect 142528 191276 142580 191282
rect 142528 191218 142580 191224
rect 142724 191162 142752 199582
rect 142802 198520 142858 198529
rect 142802 198455 142858 198464
rect 142816 196314 142844 198455
rect 142804 196308 142856 196314
rect 142804 196250 142856 196256
rect 142908 192574 142936 199679
rect 143080 199650 143132 199656
rect 143172 199708 143224 199714
rect 143506 199730 143534 200124
rect 143598 199764 143626 200124
rect 143690 199918 143718 200124
rect 143782 199918 143810 200124
rect 143874 199923 143902 200124
rect 143678 199912 143730 199918
rect 143678 199854 143730 199860
rect 143770 199912 143822 199918
rect 143770 199854 143822 199860
rect 143860 199914 143916 199923
rect 143860 199849 143916 199858
rect 143816 199776 143868 199782
rect 143598 199736 143672 199764
rect 143456 199702 143534 199730
rect 143400 199679 143456 199688
rect 143172 199650 143224 199656
rect 142986 199200 143042 199209
rect 142986 199135 143042 199144
rect 142896 192568 142948 192574
rect 142896 192510 142948 192516
rect 143000 191554 143028 199135
rect 143092 194206 143120 199650
rect 143184 195702 143212 199650
rect 143264 199640 143316 199646
rect 143448 199640 143500 199646
rect 143264 199582 143316 199588
rect 143354 199608 143410 199617
rect 143172 195696 143224 195702
rect 143172 195638 143224 195644
rect 143080 194200 143132 194206
rect 143080 194142 143132 194148
rect 142988 191548 143040 191554
rect 142988 191490 143040 191496
rect 143276 191434 143304 199582
rect 143448 199582 143500 199588
rect 143540 199640 143592 199646
rect 143540 199582 143592 199588
rect 143354 199543 143356 199552
rect 143408 199543 143410 199552
rect 143356 199514 143408 199520
rect 143356 199436 143408 199442
rect 143356 199378 143408 199384
rect 143368 199102 143396 199378
rect 143356 199096 143408 199102
rect 143356 199038 143408 199044
rect 143354 198520 143410 198529
rect 143354 198455 143410 198464
rect 143368 198286 143396 198455
rect 143356 198280 143408 198286
rect 143356 198222 143408 198228
rect 143460 195566 143488 199582
rect 143552 197810 143580 199582
rect 143540 197804 143592 197810
rect 143540 197746 143592 197752
rect 143540 197668 143592 197674
rect 143540 197610 143592 197616
rect 143448 195560 143500 195566
rect 143448 195502 143500 195508
rect 143552 194138 143580 197610
rect 143540 194132 143592 194138
rect 143540 194074 143592 194080
rect 142540 191134 142752 191162
rect 142908 191406 143304 191434
rect 142540 149054 142568 191134
rect 142908 186314 142936 191406
rect 142988 191276 143040 191282
rect 142988 191218 143040 191224
rect 142632 186286 142936 186314
rect 142528 149048 142580 149054
rect 142528 148990 142580 148996
rect 142436 148980 142488 148986
rect 142436 148922 142488 148928
rect 142632 148850 142660 186286
rect 142620 148844 142672 148850
rect 142620 148786 142672 148792
rect 143000 148306 143028 191218
rect 143644 186314 143672 199736
rect 143816 199718 143868 199724
rect 143724 199640 143776 199646
rect 143724 199582 143776 199588
rect 143736 197674 143764 199582
rect 143724 197668 143776 197674
rect 143724 197610 143776 197616
rect 143828 196926 143856 199718
rect 143966 199696 143994 200124
rect 144058 199918 144086 200124
rect 144150 199918 144178 200124
rect 144046 199912 144098 199918
rect 144046 199854 144098 199860
rect 144138 199912 144190 199918
rect 144138 199854 144190 199860
rect 144242 199696 144270 200124
rect 144334 199764 144362 200124
rect 144426 199918 144454 200124
rect 144518 199918 144546 200124
rect 144610 199918 144638 200124
rect 144414 199912 144466 199918
rect 144414 199854 144466 199860
rect 144506 199912 144558 199918
rect 144506 199854 144558 199860
rect 144598 199912 144650 199918
rect 144598 199854 144650 199860
rect 144334 199736 144408 199764
rect 143966 199668 144040 199696
rect 144242 199668 144316 199696
rect 143908 199572 143960 199578
rect 143908 199514 143960 199520
rect 143920 198830 143948 199514
rect 143908 198824 143960 198830
rect 143908 198766 143960 198772
rect 143906 198520 143962 198529
rect 143906 198455 143908 198464
rect 143960 198455 143962 198464
rect 143908 198426 143960 198432
rect 143908 197396 143960 197402
rect 143908 197338 143960 197344
rect 143816 196920 143868 196926
rect 143816 196862 143868 196868
rect 143920 193866 143948 197338
rect 144012 194594 144040 199668
rect 144184 199572 144236 199578
rect 144184 199514 144236 199520
rect 144092 198824 144144 198830
rect 144092 198766 144144 198772
rect 144104 196246 144132 198766
rect 144196 197878 144224 199514
rect 144184 197872 144236 197878
rect 144184 197814 144236 197820
rect 144092 196240 144144 196246
rect 144092 196182 144144 196188
rect 144012 194566 144132 194594
rect 143908 193860 143960 193866
rect 143908 193802 143960 193808
rect 144104 190058 144132 194566
rect 144092 190052 144144 190058
rect 144092 189994 144144 190000
rect 144288 189786 144316 199668
rect 144380 197198 144408 199736
rect 144702 199730 144730 200124
rect 144794 199850 144822 200124
rect 144886 199923 144914 200124
rect 144872 199914 144928 199923
rect 144782 199844 144834 199850
rect 144872 199849 144928 199858
rect 144782 199786 144834 199792
rect 144978 199764 145006 200124
rect 145070 199918 145098 200124
rect 145162 199918 145190 200124
rect 145058 199912 145110 199918
rect 145058 199854 145110 199860
rect 145150 199912 145202 199918
rect 145150 199854 145202 199860
rect 145254 199764 145282 200124
rect 145346 199918 145374 200124
rect 145334 199912 145386 199918
rect 145334 199854 145386 199860
rect 145438 199764 145466 200124
rect 144826 199744 144882 199753
rect 144460 199708 144512 199714
rect 144702 199702 144776 199730
rect 144460 199650 144512 199656
rect 144368 197192 144420 197198
rect 144368 197134 144420 197140
rect 144472 190126 144500 199650
rect 144552 199640 144604 199646
rect 144552 199582 144604 199588
rect 144564 197402 144592 199582
rect 144644 199572 144696 199578
rect 144644 199514 144696 199520
rect 144656 197441 144684 199514
rect 144748 198150 144776 199702
rect 144826 199679 144882 199688
rect 144932 199736 145006 199764
rect 145208 199736 145282 199764
rect 145392 199736 145466 199764
rect 145530 199764 145558 200124
rect 145622 199918 145650 200124
rect 145610 199912 145662 199918
rect 145610 199854 145662 199860
rect 145714 199764 145742 200124
rect 145806 199918 145834 200124
rect 145898 199918 145926 200124
rect 145990 199923 146018 200124
rect 145794 199912 145846 199918
rect 145794 199854 145846 199860
rect 145886 199912 145938 199918
rect 145886 199854 145938 199860
rect 145976 199914 146032 199923
rect 146082 199918 146110 200124
rect 146174 199918 146202 200124
rect 146266 199923 146294 200124
rect 145976 199849 146032 199858
rect 146070 199912 146122 199918
rect 146070 199854 146122 199860
rect 146162 199912 146214 199918
rect 146162 199854 146214 199860
rect 146252 199914 146308 199923
rect 146252 199849 146308 199858
rect 145530 199736 145604 199764
rect 144736 198144 144788 198150
rect 144736 198086 144788 198092
rect 144642 197432 144698 197441
rect 144552 197396 144604 197402
rect 144642 197367 144698 197376
rect 144552 197338 144604 197344
rect 144840 195974 144868 199679
rect 144932 198898 144960 199736
rect 145104 199708 145156 199714
rect 145104 199650 145156 199656
rect 145012 199640 145064 199646
rect 145012 199582 145064 199588
rect 144920 198892 144972 198898
rect 144920 198834 144972 198840
rect 144828 195968 144880 195974
rect 144828 195910 144880 195916
rect 145024 195294 145052 199582
rect 145116 199306 145144 199650
rect 145104 199300 145156 199306
rect 145104 199242 145156 199248
rect 145208 197470 145236 199736
rect 145288 199572 145340 199578
rect 145288 199514 145340 199520
rect 145196 197464 145248 197470
rect 145196 197406 145248 197412
rect 145300 195430 145328 199514
rect 145392 199170 145420 199736
rect 145472 199640 145524 199646
rect 145472 199582 145524 199588
rect 145380 199164 145432 199170
rect 145380 199106 145432 199112
rect 145484 195838 145512 199582
rect 145472 195832 145524 195838
rect 145472 195774 145524 195780
rect 145288 195424 145340 195430
rect 145288 195366 145340 195372
rect 145012 195288 145064 195294
rect 145012 195230 145064 195236
rect 145380 191140 145432 191146
rect 145380 191082 145432 191088
rect 144460 190120 144512 190126
rect 144460 190062 144512 190068
rect 144276 189780 144328 189786
rect 144276 189722 144328 189728
rect 143644 186286 143948 186314
rect 143632 153876 143684 153882
rect 143632 153818 143684 153824
rect 143644 151814 143672 153818
rect 143644 151786 143856 151814
rect 142988 148300 143040 148306
rect 142988 148242 143040 148248
rect 141884 147008 141936 147014
rect 141884 146950 141936 146956
rect 143632 144628 143684 144634
rect 143632 144570 143684 144576
rect 140872 144560 140924 144566
rect 140872 144502 140924 144508
rect 140320 141636 140372 141642
rect 140320 141578 140372 141584
rect 139950 140176 140006 140185
rect 139950 140111 140006 140120
rect 140332 139890 140360 141578
rect 140884 139890 140912 144502
rect 142528 144424 142580 144430
rect 142528 144366 142580 144372
rect 141424 143064 141476 143070
rect 141424 143006 141476 143012
rect 141436 139890 141464 143006
rect 142252 141500 142304 141506
rect 142252 141442 142304 141448
rect 142264 139890 142292 141442
rect 142540 139890 142568 144366
rect 143080 142928 143132 142934
rect 143080 142870 143132 142876
rect 143092 139890 143120 142870
rect 143644 139890 143672 144570
rect 143828 142154 143856 151786
rect 143920 148918 143948 186286
rect 143908 148912 143960 148918
rect 143908 148854 143960 148860
rect 145392 145858 145420 191082
rect 145576 147286 145604 199736
rect 145668 199736 145742 199764
rect 146208 199776 146260 199782
rect 145668 199238 145696 199736
rect 146358 199764 146386 200124
rect 146208 199718 146260 199724
rect 146312 199736 146386 199764
rect 145840 199708 145892 199714
rect 145840 199650 145892 199656
rect 146116 199708 146168 199714
rect 146116 199650 146168 199656
rect 145748 199572 145800 199578
rect 145748 199514 145800 199520
rect 145656 199232 145708 199238
rect 145656 199174 145708 199180
rect 145760 195226 145788 199514
rect 145852 195634 145880 199650
rect 145930 199608 145986 199617
rect 145930 199543 145986 199552
rect 146024 199572 146076 199578
rect 145944 199034 145972 199543
rect 146024 199514 146076 199520
rect 145932 199028 145984 199034
rect 145932 198970 145984 198976
rect 145840 195628 145892 195634
rect 145840 195570 145892 195576
rect 145748 195220 145800 195226
rect 145748 195162 145800 195168
rect 146036 191146 146064 199514
rect 146128 195906 146156 199650
rect 146220 198694 146248 199718
rect 146208 198688 146260 198694
rect 146208 198630 146260 198636
rect 146206 197976 146262 197985
rect 146206 197911 146262 197920
rect 146116 195900 146168 195906
rect 146116 195842 146168 195848
rect 146024 191140 146076 191146
rect 146024 191082 146076 191088
rect 146220 153882 146248 197911
rect 146312 197354 146340 199736
rect 146450 199696 146478 200124
rect 146542 199918 146570 200124
rect 146634 199918 146662 200124
rect 146530 199912 146582 199918
rect 146530 199854 146582 199860
rect 146622 199912 146674 199918
rect 146622 199854 146674 199860
rect 146726 199764 146754 200124
rect 146818 199918 146846 200124
rect 146910 199918 146938 200124
rect 147002 199918 147030 200124
rect 146806 199912 146858 199918
rect 146806 199854 146858 199860
rect 146898 199912 146950 199918
rect 146898 199854 146950 199860
rect 146990 199912 147042 199918
rect 146990 199854 147042 199860
rect 146680 199736 146754 199764
rect 146852 199776 146904 199782
rect 146450 199668 146524 199696
rect 146390 199608 146446 199617
rect 146390 199543 146446 199552
rect 146404 199374 146432 199543
rect 146392 199368 146444 199374
rect 146392 199310 146444 199316
rect 146312 197326 146432 197354
rect 146300 196784 146352 196790
rect 146300 196726 146352 196732
rect 146312 195362 146340 196726
rect 146300 195356 146352 195362
rect 146300 195298 146352 195304
rect 146404 191078 146432 197326
rect 146496 196790 146524 199668
rect 146680 198665 146708 199736
rect 147094 199764 147122 200124
rect 146852 199718 146904 199724
rect 147048 199736 147122 199764
rect 146760 199640 146812 199646
rect 146760 199582 146812 199588
rect 146666 198656 146722 198665
rect 146666 198591 146722 198600
rect 146772 197334 146800 199582
rect 146864 198626 146892 199718
rect 146944 199708 146996 199714
rect 146944 199650 146996 199656
rect 146852 198620 146904 198626
rect 146852 198562 146904 198568
rect 146760 197328 146812 197334
rect 146760 197270 146812 197276
rect 146484 196784 146536 196790
rect 146484 196726 146536 196732
rect 146956 192982 146984 199650
rect 147048 198966 147076 199736
rect 147186 199628 147214 200124
rect 147140 199600 147214 199628
rect 147036 198960 147088 198966
rect 147036 198902 147088 198908
rect 147140 195974 147168 199600
rect 147278 199560 147306 200124
rect 147370 199764 147398 200124
rect 147462 199923 147490 200124
rect 147448 199914 147504 199923
rect 147448 199849 147504 199858
rect 147554 199764 147582 200124
rect 147646 199923 147674 200124
rect 147632 199914 147688 199923
rect 147632 199849 147688 199858
rect 147370 199736 147444 199764
rect 147048 195946 147168 195974
rect 147232 199532 147306 199560
rect 146944 192976 146996 192982
rect 146944 192918 146996 192924
rect 147048 191264 147076 195946
rect 147232 195158 147260 199532
rect 147416 199510 147444 199736
rect 147508 199736 147582 199764
rect 147738 199764 147766 200124
rect 147830 199918 147858 200124
rect 147818 199912 147870 199918
rect 147818 199854 147870 199860
rect 147922 199764 147950 200124
rect 148014 199923 148042 200124
rect 148000 199914 148056 199923
rect 148000 199849 148056 199858
rect 147738 199736 147812 199764
rect 147922 199736 147996 199764
rect 147404 199504 147456 199510
rect 147404 199446 147456 199452
rect 147312 199436 147364 199442
rect 147312 199378 147364 199384
rect 147324 196858 147352 199378
rect 147404 199368 147456 199374
rect 147404 199310 147456 199316
rect 147312 196852 147364 196858
rect 147312 196794 147364 196800
rect 147220 195152 147272 195158
rect 147220 195094 147272 195100
rect 146772 191236 147076 191264
rect 146668 191140 146720 191146
rect 146668 191082 146720 191088
rect 146392 191072 146444 191078
rect 146392 191014 146444 191020
rect 146208 153876 146260 153882
rect 146208 153818 146260 153824
rect 145564 147280 145616 147286
rect 145564 147222 145616 147228
rect 145380 145852 145432 145858
rect 145380 145794 145432 145800
rect 145288 143744 145340 143750
rect 145288 143686 145340 143692
rect 145010 143032 145066 143041
rect 145010 142967 145066 142976
rect 143828 142126 144132 142154
rect 144104 139890 144132 142126
rect 145024 139890 145052 142967
rect 145300 139890 145328 143686
rect 145840 143608 145892 143614
rect 145840 143550 145892 143556
rect 145852 139890 145880 143550
rect 146390 142760 146446 142769
rect 146390 142695 146446 142704
rect 146404 139890 146432 142695
rect 146680 140214 146708 191082
rect 146772 145722 146800 191236
rect 147416 191146 147444 199310
rect 147508 192846 147536 199736
rect 147680 199640 147732 199646
rect 147680 199582 147732 199588
rect 147588 199504 147640 199510
rect 147588 199446 147640 199452
rect 147600 197130 147628 199446
rect 147588 197124 147640 197130
rect 147588 197066 147640 197072
rect 147692 196722 147720 199582
rect 147680 196716 147732 196722
rect 147680 196658 147732 196664
rect 147496 192840 147548 192846
rect 147496 192782 147548 192788
rect 147404 191140 147456 191146
rect 147404 191082 147456 191088
rect 147036 191072 147088 191078
rect 147036 191014 147088 191020
rect 146942 146160 146998 146169
rect 146942 146095 146998 146104
rect 146760 145716 146812 145722
rect 146760 145658 146812 145664
rect 146668 140208 146720 140214
rect 146668 140150 146720 140156
rect 146956 139890 146984 146095
rect 147048 145790 147076 191014
rect 147784 190454 147812 199736
rect 147862 199608 147918 199617
rect 147862 199543 147918 199552
rect 147876 196382 147904 199543
rect 147968 198914 147996 199736
rect 148106 199560 148134 200124
rect 148198 199628 148226 200124
rect 148290 199889 148318 200124
rect 148382 199918 148410 200124
rect 148474 199918 148502 200124
rect 148566 199923 148594 200124
rect 148370 199912 148422 199918
rect 148276 199880 148332 199889
rect 148370 199854 148422 199860
rect 148462 199912 148514 199918
rect 148462 199854 148514 199860
rect 148552 199914 148608 199923
rect 148658 199918 148686 200124
rect 148750 199918 148778 200124
rect 148552 199849 148608 199858
rect 148646 199912 148698 199918
rect 148646 199854 148698 199860
rect 148738 199912 148790 199918
rect 148738 199854 148790 199860
rect 148276 199815 148332 199824
rect 148416 199776 148468 199782
rect 148322 199744 148378 199753
rect 148416 199718 148468 199724
rect 148508 199776 148560 199782
rect 148508 199718 148560 199724
rect 148600 199776 148652 199782
rect 148842 199764 148870 200124
rect 148796 199736 148870 199764
rect 148652 199724 148732 199730
rect 148600 199718 148732 199724
rect 148322 199679 148378 199688
rect 148198 199600 148272 199628
rect 148106 199532 148180 199560
rect 147968 198886 148088 198914
rect 148060 198393 148088 198886
rect 148046 198384 148102 198393
rect 148046 198319 148102 198328
rect 148048 197668 148100 197674
rect 148048 197610 148100 197616
rect 147864 196376 147916 196382
rect 147864 196318 147916 196324
rect 148060 194546 148088 197610
rect 148152 197354 148180 199532
rect 148244 198665 148272 199600
rect 148230 198656 148286 198665
rect 148230 198591 148286 198600
rect 148336 197674 148364 199679
rect 148324 197668 148376 197674
rect 148324 197610 148376 197616
rect 148152 197326 148272 197354
rect 148048 194540 148100 194546
rect 148048 194482 148100 194488
rect 148140 190596 148192 190602
rect 148140 190538 148192 190544
rect 147784 190426 147996 190454
rect 147770 145888 147826 145897
rect 147770 145823 147826 145832
rect 147036 145784 147088 145790
rect 147036 145726 147088 145732
rect 147784 139890 147812 145823
rect 147968 145654 147996 190426
rect 147956 145648 148008 145654
rect 147956 145590 148008 145596
rect 148046 142896 148102 142905
rect 148046 142831 148102 142840
rect 148060 139890 148088 142831
rect 148152 140146 148180 190538
rect 148244 144498 148272 197326
rect 148428 195974 148456 199718
rect 148520 197062 148548 199718
rect 148612 199702 148732 199718
rect 148598 199608 148654 199617
rect 148598 199543 148654 199552
rect 148508 197056 148560 197062
rect 148508 196998 148560 197004
rect 148428 195946 148548 195974
rect 148520 192438 148548 195946
rect 148508 192432 148560 192438
rect 148508 192374 148560 192380
rect 148612 145926 148640 199543
rect 148704 193186 148732 199702
rect 148692 193180 148744 193186
rect 148692 193122 148744 193128
rect 148796 190602 148824 199736
rect 148934 199696 148962 200124
rect 149026 199918 149054 200124
rect 149014 199912 149066 199918
rect 149014 199854 149066 199860
rect 149118 199730 149146 200124
rect 148888 199668 148962 199696
rect 149072 199702 149146 199730
rect 149210 199730 149238 200124
rect 149302 199918 149330 200124
rect 149290 199912 149342 199918
rect 149290 199854 149342 199860
rect 149394 199764 149422 200124
rect 149486 199918 149514 200124
rect 149578 199918 149606 200124
rect 149670 199918 149698 200124
rect 149474 199912 149526 199918
rect 149474 199854 149526 199860
rect 149566 199912 149618 199918
rect 149566 199854 149618 199860
rect 149658 199912 149710 199918
rect 149658 199854 149710 199860
rect 149762 199764 149790 200124
rect 149394 199736 149468 199764
rect 149210 199702 149284 199730
rect 148888 197033 148916 199668
rect 148968 199572 149020 199578
rect 148968 199514 149020 199520
rect 148874 197024 148930 197033
rect 148874 196959 148930 196968
rect 148980 195566 149008 199514
rect 148968 195560 149020 195566
rect 148968 195502 149020 195508
rect 149072 195294 149100 199702
rect 149152 199572 149204 199578
rect 149152 199514 149204 199520
rect 149164 198762 149192 199514
rect 149152 198756 149204 198762
rect 149152 198698 149204 198704
rect 149060 195288 149112 195294
rect 149060 195230 149112 195236
rect 148784 190596 148836 190602
rect 148784 190538 148836 190544
rect 149256 187542 149284 199702
rect 149336 199640 149388 199646
rect 149336 199582 149388 199588
rect 149348 195498 149376 199582
rect 149440 198422 149468 199736
rect 149716 199736 149790 199764
rect 149520 199640 149572 199646
rect 149520 199582 149572 199588
rect 149428 198416 149480 198422
rect 149428 198358 149480 198364
rect 149532 197577 149560 199582
rect 149612 199504 149664 199510
rect 149612 199446 149664 199452
rect 149624 198121 149652 199446
rect 149610 198112 149666 198121
rect 149610 198047 149666 198056
rect 149518 197568 149574 197577
rect 149518 197503 149574 197512
rect 149428 197464 149480 197470
rect 149428 197406 149480 197412
rect 149336 195492 149388 195498
rect 149336 195434 149388 195440
rect 149336 195356 149388 195362
rect 149336 195298 149388 195304
rect 149244 187536 149296 187542
rect 149244 187478 149296 187484
rect 149348 187134 149376 195298
rect 149336 187128 149388 187134
rect 149336 187070 149388 187076
rect 149152 145988 149204 145994
rect 149152 145930 149204 145936
rect 148600 145920 148652 145926
rect 148600 145862 148652 145868
rect 148232 144492 148284 144498
rect 148232 144434 148284 144440
rect 148600 143676 148652 143682
rect 148600 143618 148652 143624
rect 148140 140140 148192 140146
rect 148140 140082 148192 140088
rect 148612 139890 148640 143618
rect 149164 139890 149192 145930
rect 149440 141438 149468 197406
rect 149716 195362 149744 199736
rect 149854 199628 149882 200124
rect 149946 199696 149974 200124
rect 150038 199764 150066 200124
rect 150130 199918 150158 200124
rect 150118 199912 150170 199918
rect 150118 199854 150170 199860
rect 150222 199764 150250 200124
rect 150038 199736 150112 199764
rect 149946 199668 150020 199696
rect 149854 199600 149928 199628
rect 149900 197266 149928 199600
rect 149888 197260 149940 197266
rect 149888 197202 149940 197208
rect 149796 197056 149848 197062
rect 149796 196998 149848 197004
rect 149704 195356 149756 195362
rect 149704 195298 149756 195304
rect 149520 195288 149572 195294
rect 149520 195230 149572 195236
rect 149532 148646 149560 195230
rect 149808 187202 149836 196998
rect 149992 196586 150020 199668
rect 149980 196580 150032 196586
rect 149980 196522 150032 196528
rect 149980 195492 150032 195498
rect 149980 195434 150032 195440
rect 149796 187196 149848 187202
rect 149796 187138 149848 187144
rect 149992 159526 150020 195434
rect 150084 192778 150112 199736
rect 150176 199736 150250 199764
rect 150176 197305 150204 199736
rect 150314 199696 150342 200124
rect 150268 199668 150342 199696
rect 150268 198121 150296 199668
rect 150406 199628 150434 200124
rect 150498 199730 150526 200124
rect 150590 199889 150618 200124
rect 150576 199880 150632 199889
rect 150576 199815 150632 199824
rect 150682 199764 150710 200124
rect 150636 199736 150710 199764
rect 150498 199702 150572 199730
rect 150360 199600 150434 199628
rect 150360 198257 150388 199600
rect 150346 198248 150402 198257
rect 150346 198183 150402 198192
rect 150254 198112 150310 198121
rect 150254 198047 150310 198056
rect 150162 197296 150218 197305
rect 150162 197231 150218 197240
rect 150438 195664 150494 195673
rect 150438 195599 150494 195608
rect 150452 195401 150480 195599
rect 150438 195392 150494 195401
rect 150438 195327 150494 195336
rect 150544 195294 150572 199702
rect 150636 195362 150664 199736
rect 150774 199696 150802 200124
rect 150866 199764 150894 200124
rect 150958 199918 150986 200124
rect 150946 199912 150998 199918
rect 150946 199854 150998 199860
rect 151050 199764 151078 200124
rect 151142 199923 151170 200124
rect 151128 199914 151184 199923
rect 151234 199918 151262 200124
rect 151128 199849 151184 199858
rect 151222 199912 151274 199918
rect 151222 199854 151274 199860
rect 151326 199764 151354 200124
rect 150866 199736 150940 199764
rect 151050 199736 151124 199764
rect 150774 199668 150848 199696
rect 150714 199608 150770 199617
rect 150714 199543 150770 199552
rect 150728 197946 150756 199543
rect 150716 197940 150768 197946
rect 150716 197882 150768 197888
rect 150716 195492 150768 195498
rect 150716 195434 150768 195440
rect 150624 195356 150676 195362
rect 150624 195298 150676 195304
rect 150532 195288 150584 195294
rect 150728 195242 150756 195434
rect 150532 195230 150584 195236
rect 150636 195214 150756 195242
rect 150072 192772 150124 192778
rect 150072 192714 150124 192720
rect 149980 159520 150032 159526
rect 149980 159462 150032 159468
rect 150636 148782 150664 195214
rect 150716 193928 150768 193934
rect 150716 193870 150768 193876
rect 150624 148776 150676 148782
rect 150624 148718 150676 148724
rect 150728 148714 150756 193870
rect 150820 152522 150848 199668
rect 150912 195974 150940 199736
rect 150912 195946 151032 195974
rect 150900 195288 150952 195294
rect 150900 195230 150952 195236
rect 150912 152590 150940 195230
rect 151004 186998 151032 195946
rect 151096 195498 151124 199736
rect 151174 199744 151230 199753
rect 151174 199679 151230 199688
rect 151280 199736 151354 199764
rect 151188 195673 151216 199679
rect 151174 195664 151230 195673
rect 151174 195599 151230 195608
rect 151084 195492 151136 195498
rect 151084 195434 151136 195440
rect 151280 195378 151308 199736
rect 151418 199594 151446 200124
rect 151510 199696 151538 200124
rect 151602 199764 151630 200124
rect 151694 199923 151722 200124
rect 151680 199914 151736 199923
rect 151786 199918 151814 200124
rect 151878 199923 151906 200124
rect 151680 199849 151736 199858
rect 151774 199912 151826 199918
rect 151774 199854 151826 199860
rect 151864 199914 151920 199923
rect 151970 199918 151998 200124
rect 151864 199849 151920 199858
rect 151958 199912 152010 199918
rect 152062 199889 152090 200124
rect 151958 199854 152010 199860
rect 152048 199880 152104 199889
rect 152048 199815 152104 199824
rect 152004 199776 152056 199782
rect 151602 199736 151676 199764
rect 151510 199668 151584 199696
rect 151418 199566 151492 199594
rect 151084 195356 151136 195362
rect 151084 195298 151136 195304
rect 151188 195350 151308 195378
rect 151096 187066 151124 195298
rect 151188 193934 151216 195350
rect 151268 195288 151320 195294
rect 151268 195230 151320 195236
rect 151176 193928 151228 193934
rect 151176 193870 151228 193876
rect 151084 187060 151136 187066
rect 151084 187002 151136 187008
rect 150992 186992 151044 186998
rect 150992 186934 151044 186940
rect 150900 152584 150952 152590
rect 150900 152526 150952 152532
rect 150808 152516 150860 152522
rect 150808 152458 150860 152464
rect 150716 148708 150768 148714
rect 150716 148650 150768 148656
rect 149520 148640 149572 148646
rect 149520 148582 149572 148588
rect 151280 142866 151308 195230
rect 151358 193896 151414 193905
rect 151358 193831 151414 193840
rect 149704 142860 149756 142866
rect 149704 142802 149756 142808
rect 151268 142860 151320 142866
rect 151268 142802 151320 142808
rect 149428 141432 149480 141438
rect 149428 141374 149480 141380
rect 149716 139890 149744 142802
rect 150532 142180 150584 142186
rect 150532 142122 150584 142128
rect 150544 139890 150572 142122
rect 151372 139890 151400 193831
rect 151464 191486 151492 199566
rect 151556 199481 151584 199668
rect 151542 199472 151598 199481
rect 151542 199407 151598 199416
rect 151648 195294 151676 199736
rect 151726 199744 151782 199753
rect 152154 199764 152182 200124
rect 152246 199918 152274 200124
rect 152338 199918 152366 200124
rect 152430 199918 152458 200124
rect 152234 199912 152286 199918
rect 152234 199854 152286 199860
rect 152326 199912 152378 199918
rect 152326 199854 152378 199860
rect 152418 199912 152470 199918
rect 152418 199854 152470 199860
rect 152004 199718 152056 199724
rect 152108 199736 152182 199764
rect 152280 199776 152332 199782
rect 151726 199679 151782 199688
rect 151912 199708 151964 199714
rect 151636 195288 151688 195294
rect 151636 195230 151688 195236
rect 151452 191480 151504 191486
rect 151452 191422 151504 191428
rect 151740 191146 151768 199679
rect 151912 199650 151964 199656
rect 151924 195650 151952 199650
rect 152016 199238 152044 199718
rect 152004 199232 152056 199238
rect 152004 199174 152056 199180
rect 151832 195622 151952 195650
rect 151832 191457 151860 195622
rect 151912 195560 151964 195566
rect 151912 195502 151964 195508
rect 151818 191448 151874 191457
rect 151818 191383 151874 191392
rect 151728 191140 151780 191146
rect 151728 191082 151780 191088
rect 151924 144362 151952 195502
rect 152004 195492 152056 195498
rect 152004 195434 152056 195440
rect 152016 145761 152044 195434
rect 152108 159458 152136 199736
rect 152280 199718 152332 199724
rect 152372 199776 152424 199782
rect 152522 199764 152550 200124
rect 152372 199718 152424 199724
rect 152476 199736 152550 199764
rect 152188 199640 152240 199646
rect 152188 199582 152240 199588
rect 152200 195974 152228 199582
rect 152292 198121 152320 199718
rect 152278 198112 152334 198121
rect 152278 198047 152334 198056
rect 152384 195974 152412 199718
rect 152188 195968 152240 195974
rect 152188 195910 152240 195916
rect 152292 195946 152412 195974
rect 152292 195566 152320 195946
rect 152280 195560 152332 195566
rect 152280 195502 152332 195508
rect 152476 195498 152504 199736
rect 152614 199696 152642 200124
rect 152706 199918 152734 200124
rect 152798 199918 152826 200124
rect 152890 199918 152918 200124
rect 152694 199912 152746 199918
rect 152694 199854 152746 199860
rect 152786 199912 152838 199918
rect 152786 199854 152838 199860
rect 152878 199912 152930 199918
rect 152982 199889 153010 200124
rect 153074 199918 153102 200124
rect 153062 199912 153114 199918
rect 152878 199854 152930 199860
rect 152968 199880 153024 199889
rect 153062 199854 153114 199860
rect 152968 199815 153024 199824
rect 152740 199776 152792 199782
rect 152740 199718 152792 199724
rect 152832 199776 152884 199782
rect 153166 199764 153194 200124
rect 152832 199718 152884 199724
rect 153120 199736 153194 199764
rect 152568 199668 152642 199696
rect 152568 199374 152596 199668
rect 152752 199594 152780 199718
rect 152660 199566 152780 199594
rect 152556 199368 152608 199374
rect 152556 199310 152608 199316
rect 152464 195492 152516 195498
rect 152464 195434 152516 195440
rect 152660 195378 152688 199566
rect 152740 199504 152792 199510
rect 152740 199446 152792 199452
rect 152200 195350 152688 195378
rect 152096 159452 152148 159458
rect 152096 159394 152148 159400
rect 152200 159390 152228 195350
rect 152752 195276 152780 199446
rect 152844 198937 152872 199718
rect 153014 199472 153070 199481
rect 152924 199436 152976 199442
rect 153120 199442 153148 199736
rect 153258 199696 153286 200124
rect 153350 199918 153378 200124
rect 153442 199918 153470 200124
rect 153338 199912 153390 199918
rect 153338 199854 153390 199860
rect 153430 199912 153482 199918
rect 153430 199854 153482 199860
rect 153384 199776 153436 199782
rect 153534 199764 153562 200124
rect 153626 199918 153654 200124
rect 153718 199918 153746 200124
rect 153810 199918 153838 200124
rect 153902 199918 153930 200124
rect 153994 199918 154022 200124
rect 153614 199912 153666 199918
rect 153614 199854 153666 199860
rect 153706 199912 153758 199918
rect 153706 199854 153758 199860
rect 153798 199912 153850 199918
rect 153798 199854 153850 199860
rect 153890 199912 153942 199918
rect 153890 199854 153942 199860
rect 153982 199912 154034 199918
rect 153982 199854 154034 199860
rect 153384 199718 153436 199724
rect 153488 199736 153562 199764
rect 153660 199776 153712 199782
rect 153212 199668 153286 199696
rect 153212 199617 153240 199668
rect 153198 199608 153254 199617
rect 153198 199543 153254 199552
rect 153200 199504 153252 199510
rect 153200 199446 153252 199452
rect 153014 199407 153070 199416
rect 153108 199436 153160 199442
rect 152924 199378 152976 199384
rect 152830 198928 152886 198937
rect 152830 198863 152886 198872
rect 152832 195968 152884 195974
rect 152832 195910 152884 195916
rect 152292 195248 152780 195276
rect 152292 189786 152320 195248
rect 152372 195152 152424 195158
rect 152372 195094 152424 195100
rect 152384 190194 152412 195094
rect 152844 195022 152872 195910
rect 152936 195537 152964 199378
rect 152922 195528 152978 195537
rect 152922 195463 152978 195472
rect 152832 195016 152884 195022
rect 152832 194958 152884 194964
rect 152372 190188 152424 190194
rect 152372 190130 152424 190136
rect 152280 189780 152332 189786
rect 152280 189722 152332 189728
rect 152188 159384 152240 159390
rect 152188 159326 152240 159332
rect 152002 145752 152058 145761
rect 152002 145687 152058 145696
rect 151912 144356 151964 144362
rect 151912 144298 151964 144304
rect 152554 144256 152610 144265
rect 152554 144191 152610 144200
rect 151452 142996 151504 143002
rect 151452 142938 151504 142944
rect 131224 139862 131284 139890
rect 131500 139862 131836 139890
rect 131960 139862 132388 139890
rect 132604 139862 132940 139890
rect 133156 139862 133492 139890
rect 133892 139862 134044 139890
rect 134260 139862 134596 139890
rect 134812 139862 135148 139890
rect 135456 139862 135700 139890
rect 135916 139862 136252 139890
rect 136652 139862 136804 139890
rect 137020 139862 137356 139890
rect 137572 139862 137908 139890
rect 138124 139862 138460 139890
rect 138676 139862 139012 139890
rect 139412 139862 139564 139890
rect 139780 139862 140116 139890
rect 140332 139862 140668 139890
rect 140884 139862 141220 139890
rect 141436 139862 141772 139890
rect 142264 139862 142324 139890
rect 142540 139862 142876 139890
rect 143092 139862 143428 139890
rect 143644 139862 143980 139890
rect 144104 139862 144532 139890
rect 145024 139862 145084 139890
rect 145300 139862 145636 139890
rect 145852 139862 146188 139890
rect 146404 139862 146740 139890
rect 146956 139862 147292 139890
rect 147784 139862 147844 139890
rect 148060 139862 148396 139890
rect 148612 139862 148948 139890
rect 149164 139862 149500 139890
rect 149716 139862 150052 139890
rect 150544 139862 150604 139890
rect 151156 139862 151400 139890
rect 151464 139890 151492 142938
rect 152568 139890 152596 144191
rect 153028 141681 153056 199407
rect 153108 199378 153160 199384
rect 153212 198734 153240 199446
rect 153120 198706 153240 198734
rect 153120 195158 153148 198706
rect 153396 197354 153424 199718
rect 153304 197326 153424 197354
rect 153304 195974 153332 197326
rect 153212 195946 153332 195974
rect 153108 195152 153160 195158
rect 153108 195094 153160 195100
rect 153212 193730 153240 195946
rect 153488 195430 153516 199736
rect 153660 199718 153712 199724
rect 153936 199776 153988 199782
rect 154086 199730 154114 200124
rect 153936 199718 153988 199724
rect 153568 199640 153620 199646
rect 153568 199582 153620 199588
rect 153580 199306 153608 199582
rect 153568 199300 153620 199306
rect 153568 199242 153620 199248
rect 153476 195424 153528 195430
rect 153476 195366 153528 195372
rect 153568 195356 153620 195362
rect 153568 195298 153620 195304
rect 153476 195288 153528 195294
rect 153476 195230 153528 195236
rect 153292 195220 153344 195226
rect 153292 195162 153344 195168
rect 153200 193724 153252 193730
rect 153200 193666 153252 193672
rect 153304 145858 153332 195162
rect 153384 195152 153436 195158
rect 153384 195094 153436 195100
rect 153396 146033 153424 195094
rect 153488 148345 153516 195230
rect 153580 187270 153608 195298
rect 153672 190262 153700 199718
rect 153752 199708 153804 199714
rect 153752 199650 153804 199656
rect 153764 199345 153792 199650
rect 153844 199572 153896 199578
rect 153844 199514 153896 199520
rect 153750 199336 153806 199345
rect 153750 199271 153806 199280
rect 153856 195226 153884 199514
rect 153948 195634 153976 199718
rect 154040 199702 154114 199730
rect 154178 199730 154206 200124
rect 154270 199918 154298 200124
rect 154258 199912 154310 199918
rect 154258 199854 154310 199860
rect 154362 199764 154390 200124
rect 154454 199918 154482 200124
rect 154442 199912 154494 199918
rect 154442 199854 154494 199860
rect 154546 199764 154574 200124
rect 154362 199736 154436 199764
rect 154178 199702 154252 199730
rect 153936 195628 153988 195634
rect 153936 195570 153988 195576
rect 154040 195294 154068 199702
rect 154120 199572 154172 199578
rect 154120 199514 154172 199520
rect 154028 195288 154080 195294
rect 154028 195230 154080 195236
rect 154132 195226 154160 199514
rect 154224 198121 154252 199702
rect 154304 199640 154356 199646
rect 154304 199582 154356 199588
rect 154210 198112 154266 198121
rect 154210 198047 154266 198056
rect 154212 195424 154264 195430
rect 154212 195366 154264 195372
rect 153844 195220 153896 195226
rect 153844 195162 153896 195168
rect 154120 195220 154172 195226
rect 154120 195162 154172 195168
rect 153660 190256 153712 190262
rect 153660 190198 153712 190204
rect 153568 187264 153620 187270
rect 153568 187206 153620 187212
rect 153568 152584 153620 152590
rect 153568 152526 153620 152532
rect 153474 148336 153530 148345
rect 153474 148271 153530 148280
rect 153382 146024 153438 146033
rect 153382 145959 153438 145968
rect 153292 145852 153344 145858
rect 153292 145794 153344 145800
rect 153106 144120 153162 144129
rect 153106 144055 153162 144064
rect 153014 141672 153070 141681
rect 153014 141607 153070 141616
rect 153120 139890 153148 144055
rect 153580 139890 153608 152526
rect 153660 141568 153712 141574
rect 153660 141510 153712 141516
rect 151464 139862 151708 139890
rect 152260 139862 152596 139890
rect 152812 139862 153148 139890
rect 153364 139862 153608 139890
rect 153672 139890 153700 141510
rect 154224 141438 154252 195366
rect 154316 195362 154344 199582
rect 154304 195356 154356 195362
rect 154304 195298 154356 195304
rect 154408 195158 154436 199736
rect 154500 199736 154574 199764
rect 154500 195906 154528 199736
rect 154638 199696 154666 200124
rect 154730 199764 154758 200124
rect 154822 199889 154850 200124
rect 154808 199880 154864 199889
rect 154808 199815 154864 199824
rect 154914 199764 154942 200124
rect 154730 199736 154804 199764
rect 154638 199668 154712 199696
rect 154684 198558 154712 199668
rect 154672 198552 154724 198558
rect 154672 198494 154724 198500
rect 154488 195900 154540 195906
rect 154488 195842 154540 195848
rect 154776 195838 154804 199736
rect 154868 199736 154942 199764
rect 154868 197946 154896 199736
rect 155006 199696 155034 200124
rect 155098 199764 155126 200124
rect 155190 199918 155218 200124
rect 155178 199912 155230 199918
rect 155282 199889 155310 200124
rect 155374 199918 155402 200124
rect 155466 199918 155494 200124
rect 155362 199912 155414 199918
rect 155178 199854 155230 199860
rect 155268 199880 155324 199889
rect 155362 199854 155414 199860
rect 155454 199912 155506 199918
rect 155558 199889 155586 200124
rect 155454 199854 155506 199860
rect 155544 199880 155600 199889
rect 155268 199815 155324 199824
rect 155544 199815 155600 199824
rect 155408 199776 155460 199782
rect 155098 199736 155172 199764
rect 155006 199668 155080 199696
rect 154856 197940 154908 197946
rect 154856 197882 154908 197888
rect 154764 195832 154816 195838
rect 154764 195774 154816 195780
rect 154396 195152 154448 195158
rect 154396 195094 154448 195100
rect 155052 193798 155080 199668
rect 155144 198966 155172 199736
rect 155314 199744 155370 199753
rect 155224 199708 155276 199714
rect 155650 199764 155678 200124
rect 155742 199918 155770 200124
rect 155834 199918 155862 200124
rect 155926 199918 155954 200124
rect 155730 199912 155782 199918
rect 155730 199854 155782 199860
rect 155822 199912 155874 199918
rect 155822 199854 155874 199860
rect 155914 199912 155966 199918
rect 155914 199854 155966 199860
rect 155408 199718 155460 199724
rect 155498 199744 155554 199753
rect 155314 199679 155370 199688
rect 155224 199650 155276 199656
rect 155132 198960 155184 198966
rect 155132 198902 155184 198908
rect 155040 193792 155092 193798
rect 155040 193734 155092 193740
rect 155236 180794 155264 199650
rect 155328 198014 155356 199679
rect 155316 198008 155368 198014
rect 155316 197950 155368 197956
rect 155420 195158 155448 199718
rect 155498 199679 155554 199688
rect 155604 199736 155678 199764
rect 155776 199776 155828 199782
rect 155408 195152 155460 195158
rect 155408 195094 155460 195100
rect 155512 193866 155540 199679
rect 155604 198218 155632 199736
rect 155776 199718 155828 199724
rect 155868 199776 155920 199782
rect 156018 199730 156046 200124
rect 155868 199718 155920 199724
rect 155684 199640 155736 199646
rect 155684 199582 155736 199588
rect 155592 198212 155644 198218
rect 155592 198154 155644 198160
rect 155696 195276 155724 199582
rect 155604 195248 155724 195276
rect 155500 193860 155552 193866
rect 155500 193802 155552 193808
rect 154684 180766 155264 180794
rect 154486 144392 154542 144401
rect 154684 144362 154712 180766
rect 154856 152720 154908 152726
rect 154856 152662 154908 152668
rect 154486 144327 154542 144336
rect 154672 144356 154724 144362
rect 154212 141432 154264 141438
rect 154212 141374 154264 141380
rect 154500 140162 154528 144327
rect 154672 144298 154724 144304
rect 154454 140134 154528 140162
rect 153672 139862 153916 139890
rect 154454 139876 154482 140134
rect 154868 139890 154896 152662
rect 155604 141545 155632 195248
rect 155684 195152 155736 195158
rect 155684 195094 155736 195100
rect 155696 152522 155724 195094
rect 155788 192506 155816 199718
rect 155880 198801 155908 199718
rect 155972 199702 156046 199730
rect 155972 199617 156000 199702
rect 156110 199628 156138 200124
rect 156202 199696 156230 200124
rect 156294 199764 156322 200124
rect 156386 199918 156414 200124
rect 156478 199918 156506 200124
rect 156570 199918 156598 200124
rect 156374 199912 156426 199918
rect 156374 199854 156426 199860
rect 156466 199912 156518 199918
rect 156466 199854 156518 199860
rect 156558 199912 156610 199918
rect 156558 199854 156610 199860
rect 156662 199764 156690 200124
rect 156294 199736 156368 199764
rect 156202 199668 156276 199696
rect 155958 199608 156014 199617
rect 155958 199543 156014 199552
rect 156064 199600 156138 199628
rect 156248 199617 156276 199668
rect 156234 199608 156290 199617
rect 155958 199200 156014 199209
rect 155958 199135 156014 199144
rect 155866 198792 155922 198801
rect 155866 198727 155922 198736
rect 155868 197328 155920 197334
rect 155868 197270 155920 197276
rect 155776 192500 155828 192506
rect 155776 192442 155828 192448
rect 155880 156670 155908 197270
rect 155972 196858 156000 199135
rect 155960 196852 156012 196858
rect 155960 196794 156012 196800
rect 155960 195288 156012 195294
rect 155960 195230 156012 195236
rect 155868 156664 155920 156670
rect 155868 156606 155920 156612
rect 155684 152516 155736 152522
rect 155684 152458 155736 152464
rect 155972 143070 156000 195230
rect 156064 193662 156092 199600
rect 156234 199543 156290 199552
rect 156236 199504 156288 199510
rect 156236 199446 156288 199452
rect 156142 199336 156198 199345
rect 156142 199271 156198 199280
rect 156156 197849 156184 199271
rect 156142 197840 156198 197849
rect 156142 197775 156198 197784
rect 156248 197538 156276 199446
rect 156236 197532 156288 197538
rect 156236 197474 156288 197480
rect 156052 193656 156104 193662
rect 156052 193598 156104 193604
rect 156144 190596 156196 190602
rect 156144 190538 156196 190544
rect 156156 148850 156184 190538
rect 156340 190454 156368 199736
rect 156524 199736 156690 199764
rect 156420 199436 156472 199442
rect 156420 199378 156472 199384
rect 156432 198121 156460 199378
rect 156418 198112 156474 198121
rect 156418 198047 156474 198056
rect 156524 197878 156552 199736
rect 156754 199696 156782 200124
rect 156846 199730 156874 200124
rect 156938 199918 156966 200124
rect 157030 199918 157058 200124
rect 157122 199918 157150 200124
rect 157214 199923 157242 200124
rect 156926 199912 156978 199918
rect 156926 199854 156978 199860
rect 157018 199912 157070 199918
rect 157018 199854 157070 199860
rect 157110 199912 157162 199918
rect 157110 199854 157162 199860
rect 157200 199914 157256 199923
rect 157200 199849 157256 199858
rect 157306 199764 157334 200124
rect 157398 199923 157426 200124
rect 157384 199914 157440 199923
rect 157490 199918 157518 200124
rect 157582 199923 157610 200124
rect 157384 199849 157440 199858
rect 157478 199912 157530 199918
rect 157478 199854 157530 199860
rect 157568 199914 157624 199923
rect 157568 199849 157624 199858
rect 157154 199744 157210 199753
rect 156846 199702 156920 199730
rect 156708 199668 156782 199696
rect 156604 199640 156656 199646
rect 156604 199582 156656 199588
rect 156616 198082 156644 199582
rect 156604 198076 156656 198082
rect 156604 198018 156656 198024
rect 156512 197872 156564 197878
rect 156512 197814 156564 197820
rect 156708 195498 156736 199668
rect 156786 199336 156842 199345
rect 156786 199271 156788 199280
rect 156840 199271 156842 199280
rect 156788 199242 156840 199248
rect 156696 195492 156748 195498
rect 156696 195434 156748 195440
rect 156892 195294 156920 199702
rect 157064 199708 157116 199714
rect 157154 199679 157210 199688
rect 157260 199736 157334 199764
rect 157524 199776 157576 199782
rect 157064 199650 157116 199656
rect 156972 199640 157024 199646
rect 156972 199582 157024 199588
rect 156880 195288 156932 195294
rect 156880 195230 156932 195236
rect 156984 192545 157012 199582
rect 156970 192536 157026 192545
rect 156970 192471 157026 192480
rect 157076 190602 157104 199650
rect 157168 192710 157196 199679
rect 157260 198121 157288 199736
rect 157674 199730 157702 200124
rect 157524 199718 157576 199724
rect 157338 198248 157394 198257
rect 157338 198183 157394 198192
rect 157246 198112 157302 198121
rect 157246 198047 157302 198056
rect 157248 197124 157300 197130
rect 157248 197066 157300 197072
rect 157156 192704 157208 192710
rect 157156 192646 157208 192652
rect 157064 190596 157116 190602
rect 157064 190538 157116 190544
rect 156340 190426 156920 190454
rect 156144 148844 156196 148850
rect 156144 148786 156196 148792
rect 156892 145625 156920 190426
rect 157260 154154 157288 197066
rect 157248 154148 157300 154154
rect 157248 154090 157300 154096
rect 157352 151434 157380 198183
rect 157536 197674 157564 199718
rect 157628 199702 157702 199730
rect 157628 198393 157656 199702
rect 157766 199696 157794 200124
rect 157858 199918 157886 200124
rect 157846 199912 157898 199918
rect 157846 199854 157898 199860
rect 157950 199764 157978 200124
rect 158042 199918 158070 200124
rect 158134 199923 158162 200124
rect 158030 199912 158082 199918
rect 158030 199854 158082 199860
rect 158120 199914 158176 199923
rect 158120 199849 158176 199858
rect 158226 199764 158254 200124
rect 158318 199918 158346 200124
rect 158410 199918 158438 200124
rect 158502 199923 158530 200124
rect 158306 199912 158358 199918
rect 158306 199854 158358 199860
rect 158398 199912 158450 199918
rect 158398 199854 158450 199860
rect 158488 199914 158544 199923
rect 158594 199918 158622 200124
rect 158686 199918 158714 200124
rect 158778 199918 158806 200124
rect 158488 199849 158544 199858
rect 158582 199912 158634 199918
rect 158582 199854 158634 199860
rect 158674 199912 158726 199918
rect 158674 199854 158726 199860
rect 158766 199912 158818 199918
rect 158766 199854 158818 199860
rect 157904 199736 157978 199764
rect 158074 199744 158130 199753
rect 157766 199668 157840 199696
rect 157614 198384 157670 198393
rect 157614 198319 157670 198328
rect 157524 197668 157576 197674
rect 157524 197610 157576 197616
rect 157812 195974 157840 199668
rect 157800 195968 157852 195974
rect 157800 195910 157852 195916
rect 157616 195764 157668 195770
rect 157616 195706 157668 195712
rect 157628 195294 157656 195706
rect 157616 195288 157668 195294
rect 157616 195230 157668 195236
rect 157904 194002 157932 199736
rect 158074 199679 158130 199688
rect 158180 199736 158254 199764
rect 158628 199776 158680 199782
rect 158626 199744 158628 199753
rect 158720 199776 158772 199782
rect 158680 199744 158682 199753
rect 157984 199640 158036 199646
rect 157984 199582 158036 199588
rect 157432 193996 157484 194002
rect 157432 193938 157484 193944
rect 157892 193996 157944 194002
rect 157892 193938 157944 193944
rect 157444 151502 157472 193938
rect 157996 192574 158024 199582
rect 158088 198830 158116 199679
rect 158076 198824 158128 198830
rect 158076 198766 158128 198772
rect 158076 197872 158128 197878
rect 158076 197814 158128 197820
rect 158088 195498 158116 197814
rect 158076 195492 158128 195498
rect 158076 195434 158128 195440
rect 157984 192568 158036 192574
rect 157984 192510 158036 192516
rect 157524 191072 157576 191078
rect 157524 191014 157576 191020
rect 157536 154290 157564 191014
rect 158180 186314 158208 199736
rect 158352 199708 158404 199714
rect 158352 199650 158404 199656
rect 158536 199708 158588 199714
rect 158870 199764 158898 200124
rect 158962 199918 158990 200124
rect 159054 199918 159082 200124
rect 159146 199918 159174 200124
rect 158950 199912 159002 199918
rect 158950 199854 159002 199860
rect 159042 199912 159094 199918
rect 159042 199854 159094 199860
rect 159134 199912 159186 199918
rect 159134 199854 159186 199860
rect 159238 199764 159266 200124
rect 159330 199923 159358 200124
rect 159316 199914 159372 199923
rect 159316 199849 159372 199858
rect 159422 199764 159450 200124
rect 158870 199753 158944 199764
rect 158870 199744 158958 199753
rect 158870 199736 158902 199744
rect 158720 199718 158772 199724
rect 158626 199679 158682 199688
rect 158536 199650 158588 199656
rect 158258 199608 158314 199617
rect 158258 199543 158314 199552
rect 158272 199073 158300 199543
rect 158364 199442 158392 199650
rect 158442 199608 158498 199617
rect 158442 199543 158498 199552
rect 158352 199436 158404 199442
rect 158352 199378 158404 199384
rect 158258 199064 158314 199073
rect 158258 198999 158314 199008
rect 158456 191078 158484 199543
rect 158444 191072 158496 191078
rect 158444 191014 158496 191020
rect 158548 189854 158576 199650
rect 158628 199572 158680 199578
rect 158628 199514 158680 199520
rect 158640 198801 158668 199514
rect 158626 198792 158682 198801
rect 158626 198727 158682 198736
rect 158732 197130 158760 199718
rect 159192 199736 159266 199764
rect 159376 199736 159450 199764
rect 159514 199764 159542 200124
rect 159606 199918 159634 200124
rect 159698 199923 159726 200124
rect 159594 199912 159646 199918
rect 159594 199854 159646 199860
rect 159684 199914 159740 199923
rect 159790 199918 159818 200124
rect 159882 199918 159910 200124
rect 159684 199849 159740 199858
rect 159778 199912 159830 199918
rect 159778 199854 159830 199860
rect 159870 199912 159922 199918
rect 159870 199854 159922 199860
rect 159640 199776 159692 199782
rect 159514 199736 159588 199764
rect 158902 199679 158958 199688
rect 158996 199708 159048 199714
rect 158996 199650 159048 199656
rect 159088 199708 159140 199714
rect 159088 199650 159140 199656
rect 158902 199608 158958 199617
rect 158812 199572 158864 199578
rect 158902 199543 158958 199552
rect 158812 199514 158864 199520
rect 158720 197124 158772 197130
rect 158720 197066 158772 197072
rect 158628 196580 158680 196586
rect 158628 196522 158680 196528
rect 158536 189848 158588 189854
rect 158536 189790 158588 189796
rect 157628 186286 158208 186314
rect 157524 154284 157576 154290
rect 157524 154226 157576 154232
rect 157628 154222 157656 186286
rect 157616 154216 157668 154222
rect 157616 154158 157668 154164
rect 157432 151496 157484 151502
rect 157432 151438 157484 151444
rect 157340 151428 157392 151434
rect 157340 151370 157392 151376
rect 158640 149734 158668 196522
rect 158720 151224 158772 151230
rect 158720 151166 158772 151172
rect 158628 149728 158680 149734
rect 158628 149670 158680 149676
rect 156878 145616 156934 145625
rect 156878 145551 156934 145560
rect 157338 145616 157394 145625
rect 157338 145551 157394 145560
rect 156418 144528 156474 144537
rect 156418 144463 156474 144472
rect 155960 143064 156012 143070
rect 155960 143006 156012 143012
rect 155776 142180 155828 142186
rect 155776 142122 155828 142128
rect 155590 141536 155646 141545
rect 155590 141471 155646 141480
rect 155788 139890 155816 142122
rect 156432 139890 156460 144463
rect 156970 142896 157026 142905
rect 156970 142831 157026 142840
rect 156984 139890 157012 142831
rect 157154 141672 157210 141681
rect 157154 141607 157210 141616
rect 154868 139862 155020 139890
rect 155572 139862 155816 139890
rect 156124 139862 156460 139890
rect 156676 139862 157012 139890
rect 157168 139890 157196 141607
rect 157352 139890 157380 145551
rect 158628 142996 158680 143002
rect 158628 142938 158680 142944
rect 157432 142180 157484 142186
rect 157432 142122 157484 142128
rect 157444 142089 157472 142122
rect 157430 142080 157486 142089
rect 157430 142015 157486 142024
rect 158640 139890 158668 142938
rect 158732 140758 158760 151166
rect 158824 147150 158852 199514
rect 158916 195265 158944 199543
rect 159008 198558 159036 199650
rect 158996 198552 159048 198558
rect 158996 198494 159048 198500
rect 158902 195256 158958 195265
rect 158902 195191 158958 195200
rect 158902 194032 158958 194041
rect 158902 193967 158958 193976
rect 158916 154426 158944 193967
rect 159100 186402 159128 199650
rect 159192 197878 159220 199736
rect 159272 199640 159324 199646
rect 159272 199582 159324 199588
rect 159180 197872 159232 197878
rect 159180 197814 159232 197820
rect 159180 197532 159232 197538
rect 159180 197474 159232 197480
rect 159192 192642 159220 197474
rect 159180 192636 159232 192642
rect 159180 192578 159232 192584
rect 159284 191690 159312 199582
rect 159272 191684 159324 191690
rect 159272 191626 159324 191632
rect 159376 191418 159404 199736
rect 159456 199640 159508 199646
rect 159456 199582 159508 199588
rect 159468 195906 159496 199582
rect 159560 197470 159588 199736
rect 159974 199764 160002 200124
rect 160066 199918 160094 200124
rect 160158 199918 160186 200124
rect 160250 199918 160278 200124
rect 160342 199918 160370 200124
rect 160054 199912 160106 199918
rect 160054 199854 160106 199860
rect 160146 199912 160198 199918
rect 160146 199854 160198 199860
rect 160238 199912 160290 199918
rect 160238 199854 160290 199860
rect 160330 199912 160382 199918
rect 160330 199854 160382 199860
rect 160192 199776 160244 199782
rect 159974 199736 160048 199764
rect 159640 199718 159692 199724
rect 159548 197464 159600 197470
rect 159548 197406 159600 197412
rect 159456 195900 159508 195906
rect 159456 195842 159508 195848
rect 159364 191412 159416 191418
rect 159364 191354 159416 191360
rect 159008 186374 159128 186402
rect 158904 154420 158956 154426
rect 158904 154362 158956 154368
rect 159008 154358 159036 186374
rect 159652 186314 159680 199718
rect 159732 199640 159784 199646
rect 159732 199582 159784 199588
rect 159914 199608 159970 199617
rect 159744 198490 159772 199582
rect 159914 199543 159970 199552
rect 159732 198484 159784 198490
rect 159732 198426 159784 198432
rect 159928 191486 159956 199543
rect 159916 191480 159968 191486
rect 159916 191422 159968 191428
rect 160020 190330 160048 199736
rect 160192 199718 160244 199724
rect 160284 199776 160336 199782
rect 160434 199764 160462 200124
rect 160284 199718 160336 199724
rect 160388 199736 160462 199764
rect 160526 199764 160554 200124
rect 160618 199923 160646 200124
rect 160604 199914 160660 199923
rect 160710 199918 160738 200124
rect 160604 199849 160660 199858
rect 160698 199912 160750 199918
rect 160698 199854 160750 199860
rect 160652 199776 160704 199782
rect 160526 199753 160600 199764
rect 160526 199744 160614 199753
rect 160526 199736 160558 199744
rect 160100 199368 160152 199374
rect 160100 199310 160152 199316
rect 160112 199209 160140 199310
rect 160098 199200 160154 199209
rect 160098 199135 160154 199144
rect 160204 191214 160232 199718
rect 160296 196586 160324 199718
rect 160284 196580 160336 196586
rect 160284 196522 160336 196528
rect 160284 191276 160336 191282
rect 160284 191218 160336 191224
rect 160192 191208 160244 191214
rect 160192 191150 160244 191156
rect 160192 191072 160244 191078
rect 160192 191014 160244 191020
rect 160008 190324 160060 190330
rect 160008 190266 160060 190272
rect 159652 186286 160048 186314
rect 158996 154352 159048 154358
rect 158996 154294 159048 154300
rect 158904 150272 158956 150278
rect 158904 150214 158956 150220
rect 158812 147144 158864 147150
rect 158812 147086 158864 147092
rect 158720 140752 158772 140758
rect 158720 140694 158772 140700
rect 158916 140162 158944 150214
rect 160020 147286 160048 186286
rect 160100 151156 160152 151162
rect 160100 151098 160152 151104
rect 160008 147280 160060 147286
rect 160008 147222 160060 147228
rect 159640 140752 159692 140758
rect 159640 140694 159692 140700
rect 159548 140684 159600 140690
rect 159548 140626 159600 140632
rect 157168 139862 157228 139890
rect 157352 139862 157780 139890
rect 158332 139862 158668 139890
rect 158870 140134 158944 140162
rect 158870 139876 158898 140134
rect 159560 139890 159588 140626
rect 159436 139862 159588 139890
rect 159652 139890 159680 140694
rect 160112 139890 160140 151098
rect 160204 141574 160232 191014
rect 160296 144430 160324 191218
rect 160388 147422 160416 199736
rect 160802 199730 160830 200124
rect 160894 199918 160922 200124
rect 160882 199912 160934 199918
rect 160882 199854 160934 199860
rect 160986 199764 161014 200124
rect 161078 199918 161106 200124
rect 161170 199918 161198 200124
rect 161066 199912 161118 199918
rect 161066 199854 161118 199860
rect 161158 199912 161210 199918
rect 161158 199854 161210 199860
rect 161262 199764 161290 200124
rect 160652 199718 160704 199724
rect 160558 199679 160614 199688
rect 160558 199608 160614 199617
rect 160558 199543 160614 199552
rect 160468 199504 160520 199510
rect 160468 199446 160520 199452
rect 160480 195566 160508 199446
rect 160468 195560 160520 195566
rect 160468 195502 160520 195508
rect 160468 193180 160520 193186
rect 160468 193122 160520 193128
rect 160480 191298 160508 193122
rect 160572 192930 160600 199543
rect 160664 193186 160692 199718
rect 160756 199702 160830 199730
rect 160940 199736 161014 199764
rect 161216 199736 161290 199764
rect 161354 199764 161382 200124
rect 161446 199923 161474 200124
rect 161432 199914 161488 199923
rect 161432 199849 161488 199858
rect 161538 199764 161566 200124
rect 161630 199918 161658 200124
rect 161722 199918 161750 200124
rect 161814 199918 161842 200124
rect 161906 199918 161934 200124
rect 161618 199912 161670 199918
rect 161618 199854 161670 199860
rect 161710 199912 161762 199918
rect 161710 199854 161762 199860
rect 161802 199912 161854 199918
rect 161802 199854 161854 199860
rect 161894 199912 161946 199918
rect 161894 199854 161946 199860
rect 161664 199776 161716 199782
rect 161354 199736 161428 199764
rect 161538 199736 161612 199764
rect 160756 194594 160784 199702
rect 160836 199640 160888 199646
rect 160836 199582 160888 199588
rect 160848 197130 160876 199582
rect 160836 197124 160888 197130
rect 160836 197066 160888 197072
rect 160756 194566 160876 194594
rect 160652 193180 160704 193186
rect 160652 193122 160704 193128
rect 160572 192902 160692 192930
rect 160480 191270 160600 191298
rect 160468 191208 160520 191214
rect 160468 191150 160520 191156
rect 160376 147416 160428 147422
rect 160376 147358 160428 147364
rect 160480 147082 160508 191150
rect 160572 147218 160600 191270
rect 160664 190097 160692 192902
rect 160848 192710 160876 194566
rect 160836 192704 160888 192710
rect 160836 192646 160888 192652
rect 160650 190088 160706 190097
rect 160650 190023 160706 190032
rect 160940 186314 160968 199736
rect 161112 199708 161164 199714
rect 161112 199650 161164 199656
rect 161020 199640 161072 199646
rect 161020 199582 161072 199588
rect 161032 194594 161060 199582
rect 161124 195401 161152 199650
rect 161110 195392 161166 195401
rect 161110 195327 161166 195336
rect 161032 194566 161152 194594
rect 160664 186286 160968 186314
rect 161124 186314 161152 194566
rect 161216 191078 161244 199736
rect 161296 197872 161348 197878
rect 161296 197814 161348 197820
rect 161308 197538 161336 197814
rect 161296 197532 161348 197538
rect 161296 197474 161348 197480
rect 161400 197354 161428 199736
rect 161480 199572 161532 199578
rect 161480 199514 161532 199520
rect 161492 198898 161520 199514
rect 161480 198892 161532 198898
rect 161480 198834 161532 198840
rect 161308 197326 161428 197354
rect 161308 191282 161336 197326
rect 161296 191276 161348 191282
rect 161296 191218 161348 191224
rect 161584 191214 161612 199736
rect 161998 199764 162026 200124
rect 162090 199850 162118 200124
rect 162182 199923 162210 200124
rect 162168 199914 162224 199923
rect 162078 199844 162130 199850
rect 162168 199849 162224 199858
rect 162078 199786 162130 199792
rect 162274 199764 162302 200124
rect 161664 199718 161716 199724
rect 161952 199736 162026 199764
rect 162228 199736 162302 199764
rect 162366 199764 162394 200124
rect 162458 199923 162486 200124
rect 162444 199914 162500 199923
rect 162444 199849 162500 199858
rect 162550 199850 162578 200124
rect 162642 199918 162670 200124
rect 162734 199918 162762 200124
rect 162630 199912 162682 199918
rect 162630 199854 162682 199860
rect 162722 199912 162774 199918
rect 162722 199854 162774 199860
rect 162538 199844 162590 199850
rect 162538 199786 162590 199792
rect 162366 199736 162486 199764
rect 161572 191208 161624 191214
rect 161572 191150 161624 191156
rect 161204 191072 161256 191078
rect 161204 191014 161256 191020
rect 161572 191072 161624 191078
rect 161572 191014 161624 191020
rect 161124 186286 161244 186314
rect 160664 154494 160692 186286
rect 160744 156732 160796 156738
rect 160744 156674 160796 156680
rect 160652 154488 160704 154494
rect 160652 154430 160704 154436
rect 160560 147212 160612 147218
rect 160560 147154 160612 147160
rect 160468 147076 160520 147082
rect 160468 147018 160520 147024
rect 160284 144424 160336 144430
rect 160284 144366 160336 144372
rect 160192 141568 160244 141574
rect 160192 141510 160244 141516
rect 160756 139890 160784 156674
rect 161216 140185 161244 186286
rect 161584 145790 161612 191014
rect 161676 147014 161704 199718
rect 161848 199708 161900 199714
rect 161848 199650 161900 199656
rect 161860 197606 161888 199650
rect 161952 199034 161980 199736
rect 162032 199572 162084 199578
rect 162032 199514 162084 199520
rect 161940 199028 161992 199034
rect 161940 198970 161992 198976
rect 161848 197600 161900 197606
rect 161848 197542 161900 197548
rect 161756 191208 161808 191214
rect 161756 191150 161808 191156
rect 161768 151570 161796 191150
rect 162044 191078 162072 199514
rect 162228 197033 162256 199736
rect 162458 199730 162486 199736
rect 162826 199730 162854 200124
rect 162918 199918 162946 200124
rect 162906 199912 162958 199918
rect 162906 199854 162958 199860
rect 163010 199764 163038 200124
rect 163102 199918 163130 200124
rect 163194 199918 163222 200124
rect 163286 199918 163314 200124
rect 163378 199918 163406 200124
rect 163090 199912 163142 199918
rect 163090 199854 163142 199860
rect 163182 199912 163234 199918
rect 163182 199854 163234 199860
rect 163274 199912 163326 199918
rect 163274 199854 163326 199860
rect 163366 199912 163418 199918
rect 163366 199854 163418 199860
rect 163470 199850 163498 200124
rect 163562 199923 163590 200124
rect 163548 199914 163604 199923
rect 163458 199844 163510 199850
rect 163548 199849 163604 199858
rect 163654 199850 163682 200124
rect 163746 199889 163774 200124
rect 163838 199918 163866 200124
rect 163930 199918 163958 200124
rect 164022 199923 164050 200124
rect 163826 199912 163878 199918
rect 163732 199880 163788 199889
rect 163458 199786 163510 199792
rect 163642 199844 163694 199850
rect 163826 199854 163878 199860
rect 163918 199912 163970 199918
rect 163918 199854 163970 199860
rect 164008 199914 164064 199923
rect 164008 199849 164064 199858
rect 163732 199815 163788 199824
rect 163642 199786 163694 199792
rect 162458 199702 162624 199730
rect 162308 199640 162360 199646
rect 162308 199582 162360 199588
rect 162320 198257 162348 199582
rect 162400 199572 162452 199578
rect 162400 199514 162452 199520
rect 162492 199572 162544 199578
rect 162492 199514 162544 199520
rect 162306 198248 162362 198257
rect 162306 198183 162362 198192
rect 162412 198064 162440 199514
rect 162320 198036 162440 198064
rect 162214 197024 162270 197033
rect 162214 196959 162270 196968
rect 162214 196888 162270 196897
rect 162214 196823 162270 196832
rect 162124 195968 162176 195974
rect 162124 195910 162176 195916
rect 162136 195294 162164 195910
rect 162124 195288 162176 195294
rect 162124 195230 162176 195236
rect 162032 191072 162084 191078
rect 162032 191014 162084 191020
rect 162228 186314 162256 196823
rect 162320 191049 162348 198036
rect 162398 197840 162454 197849
rect 162398 197775 162454 197784
rect 162306 191040 162362 191049
rect 162306 190975 162362 190984
rect 162412 190398 162440 197775
rect 162504 196897 162532 199514
rect 162596 198762 162624 199702
rect 162688 199702 162854 199730
rect 162918 199736 163038 199764
rect 163136 199776 163188 199782
rect 163134 199744 163136 199753
rect 163228 199776 163280 199782
rect 163188 199744 163190 199753
rect 162584 198756 162636 198762
rect 162584 198698 162636 198704
rect 162490 196888 162546 196897
rect 162490 196823 162546 196832
rect 162688 195974 162716 199702
rect 162768 199640 162820 199646
rect 162918 199628 162946 199736
rect 163228 199718 163280 199724
rect 163502 199744 163558 199753
rect 163134 199679 163190 199688
rect 162768 199582 162820 199588
rect 162872 199600 162946 199628
rect 163044 199640 163096 199646
rect 162780 198150 162808 199582
rect 162768 198144 162820 198150
rect 162768 198086 162820 198092
rect 162596 195946 162716 195974
rect 162596 192370 162624 195946
rect 162872 193214 162900 199600
rect 163044 199582 163096 199588
rect 163134 199608 163190 199617
rect 162952 197872 163004 197878
rect 162952 197814 163004 197820
rect 162780 193186 162900 193214
rect 162584 192364 162636 192370
rect 162584 192306 162636 192312
rect 162676 192228 162728 192234
rect 162676 192170 162728 192176
rect 162400 190392 162452 190398
rect 162400 190334 162452 190340
rect 162228 186286 162532 186314
rect 161848 159656 161900 159662
rect 161848 159598 161900 159604
rect 161756 151564 161808 151570
rect 161756 151506 161808 151512
rect 161664 147008 161716 147014
rect 161664 146950 161716 146956
rect 161572 145784 161624 145790
rect 161572 145726 161624 145732
rect 161754 143032 161810 143041
rect 161754 142967 161810 142976
rect 161202 140176 161258 140185
rect 161202 140111 161258 140120
rect 161768 139890 161796 142967
rect 161860 140690 161888 159598
rect 161940 157208 161992 157214
rect 161940 157150 161992 157156
rect 161848 140684 161900 140690
rect 161848 140626 161900 140632
rect 159652 139862 159988 139890
rect 160112 139862 160540 139890
rect 160756 139862 161092 139890
rect 161644 139862 161796 139890
rect 161952 139890 161980 157150
rect 162504 142154 162532 186286
rect 162688 148918 162716 192170
rect 162676 148912 162728 148918
rect 162676 148854 162728 148860
rect 162780 145722 162808 193186
rect 162964 192234 162992 197814
rect 163056 193214 163084 199582
rect 163134 199543 163190 199552
rect 163148 198354 163176 199543
rect 163136 198348 163188 198354
rect 163136 198290 163188 198296
rect 163240 197878 163268 199718
rect 163412 199708 163464 199714
rect 163686 199744 163742 199753
rect 163502 199679 163558 199688
rect 163596 199708 163648 199714
rect 163412 199650 163464 199656
rect 163320 198144 163372 198150
rect 163320 198086 163372 198092
rect 163228 197872 163280 197878
rect 163228 197814 163280 197820
rect 163056 193186 163268 193214
rect 162952 192228 163004 192234
rect 162952 192170 163004 192176
rect 163136 191208 163188 191214
rect 163136 191150 163188 191156
rect 163148 150210 163176 191150
rect 163136 150204 163188 150210
rect 163136 150146 163188 150152
rect 163240 150074 163268 193186
rect 163228 150068 163280 150074
rect 163228 150010 163280 150016
rect 163332 149938 163360 198086
rect 163424 191078 163452 199650
rect 163516 191214 163544 199679
rect 163686 199679 163742 199688
rect 163780 199708 163832 199714
rect 163596 199650 163648 199656
rect 163608 196790 163636 199650
rect 163596 196784 163648 196790
rect 163596 196726 163648 196732
rect 163504 191208 163556 191214
rect 163504 191150 163556 191156
rect 163412 191072 163464 191078
rect 163412 191014 163464 191020
rect 163700 180794 163728 199679
rect 164114 199696 164142 200124
rect 164206 199889 164234 200124
rect 164192 199880 164248 199889
rect 164192 199815 164248 199824
rect 164298 199730 164326 200124
rect 164390 199918 164418 200124
rect 164378 199912 164430 199918
rect 164378 199854 164430 199860
rect 164482 199850 164510 200124
rect 164574 199889 164602 200124
rect 164560 199880 164616 199889
rect 164470 199844 164522 199850
rect 164560 199815 164616 199824
rect 164470 199786 164522 199792
rect 164252 199714 164326 199730
rect 163780 199650 163832 199656
rect 164068 199668 164142 199696
rect 164240 199708 164326 199714
rect 163792 191622 163820 199650
rect 163962 199608 164018 199617
rect 163962 199543 164018 199552
rect 163872 199504 163924 199510
rect 163872 199446 163924 199452
rect 163884 197266 163912 199446
rect 163872 197260 163924 197266
rect 163872 197202 163924 197208
rect 163976 194138 164004 199543
rect 163964 194132 164016 194138
rect 163964 194074 164016 194080
rect 164068 193214 164096 199668
rect 164292 199702 164326 199708
rect 164514 199744 164570 199753
rect 164514 199679 164570 199688
rect 164240 199650 164292 199656
rect 164332 199640 164384 199646
rect 164332 199582 164384 199588
rect 164240 199572 164292 199578
rect 164240 199514 164292 199520
rect 164148 199504 164200 199510
rect 164148 199446 164200 199452
rect 164160 196858 164188 199446
rect 164148 196852 164200 196858
rect 164148 196794 164200 196800
rect 164252 196625 164280 199514
rect 164238 196616 164294 196625
rect 164238 196551 164294 196560
rect 164148 194132 164200 194138
rect 164148 194074 164200 194080
rect 163976 193186 164096 193214
rect 163780 191616 163832 191622
rect 163780 191558 163832 191564
rect 163424 180766 163728 180794
rect 163424 152658 163452 180766
rect 163596 157276 163648 157282
rect 163596 157218 163648 157224
rect 163504 156596 163556 156602
rect 163504 156538 163556 156544
rect 163412 152652 163464 152658
rect 163412 152594 163464 152600
rect 163320 149932 163372 149938
rect 163320 149874 163372 149880
rect 162768 145716 162820 145722
rect 162768 145658 162820 145664
rect 162320 142126 162532 142154
rect 161952 139862 162196 139890
rect 162320 139369 162348 142126
rect 162400 140684 162452 140690
rect 162400 140626 162452 140632
rect 162412 139890 162440 140626
rect 163516 139890 163544 156538
rect 162412 139862 162748 139890
rect 163300 139862 163544 139890
rect 163608 139890 163636 157218
rect 163976 141642 164004 193186
rect 164056 191072 164108 191078
rect 164056 191014 164108 191020
rect 164068 147354 164096 191014
rect 164160 147490 164188 194074
rect 164240 191208 164292 191214
rect 164240 191150 164292 191156
rect 164148 147484 164200 147490
rect 164148 147426 164200 147432
rect 164056 147348 164108 147354
rect 164056 147290 164108 147296
rect 164252 147121 164280 191150
rect 164344 191010 164372 199582
rect 164424 199572 164476 199578
rect 164424 199514 164476 199520
rect 164436 199306 164464 199514
rect 164424 199300 164476 199306
rect 164424 199242 164476 199248
rect 164528 193214 164556 199679
rect 164666 199628 164694 200124
rect 164758 199850 164786 200124
rect 164746 199844 164798 199850
rect 164746 199786 164798 199792
rect 164850 199730 164878 200124
rect 164942 199782 164970 200124
rect 164436 193186 164556 193214
rect 164620 199600 164694 199628
rect 164804 199702 164878 199730
rect 164930 199776 164982 199782
rect 164930 199718 164982 199724
rect 164332 191004 164384 191010
rect 164332 190946 164384 190952
rect 164436 150006 164464 193186
rect 164620 191162 164648 199600
rect 164700 196580 164752 196586
rect 164700 196522 164752 196528
rect 164712 191554 164740 196522
rect 164700 191548 164752 191554
rect 164700 191490 164752 191496
rect 164804 191162 164832 199702
rect 164884 199640 164936 199646
rect 165034 199594 165062 200124
rect 165126 199889 165154 200124
rect 165218 199918 165246 200124
rect 165310 199918 165338 200124
rect 165402 199918 165430 200124
rect 165494 199918 165522 200124
rect 165206 199912 165258 199918
rect 165112 199880 165168 199889
rect 165206 199854 165258 199860
rect 165298 199912 165350 199918
rect 165298 199854 165350 199860
rect 165390 199912 165442 199918
rect 165390 199854 165442 199860
rect 165482 199912 165534 199918
rect 165482 199854 165534 199860
rect 165112 199815 165168 199824
rect 165586 199782 165614 200124
rect 165252 199776 165304 199782
rect 165574 199776 165626 199782
rect 165252 199718 165304 199724
rect 165342 199744 165398 199753
rect 165160 199708 165212 199714
rect 165160 199650 165212 199656
rect 164884 199582 164936 199588
rect 164896 196586 164924 199582
rect 164988 199566 165062 199594
rect 164988 198626 165016 199566
rect 165066 199472 165122 199481
rect 165066 199407 165122 199416
rect 164976 198620 165028 198626
rect 164976 198562 165028 198568
rect 164976 198008 165028 198014
rect 164976 197950 165028 197956
rect 164988 197849 165016 197950
rect 164974 197840 165030 197849
rect 164974 197775 165030 197784
rect 164884 196580 164936 196586
rect 164884 196522 164936 196528
rect 164528 191134 164648 191162
rect 164712 191134 164832 191162
rect 164424 150000 164476 150006
rect 164424 149942 164476 149948
rect 164528 149802 164556 191134
rect 164608 191072 164660 191078
rect 164608 191014 164660 191020
rect 164620 151638 164648 191014
rect 164712 152794 164740 191134
rect 165080 191078 165108 199407
rect 165172 195974 165200 199650
rect 165264 197305 165292 199718
rect 165574 199718 165626 199724
rect 165342 199679 165398 199688
rect 165678 199696 165706 200124
rect 165770 199923 165798 200124
rect 165756 199914 165812 199923
rect 165862 199918 165890 200124
rect 165954 199918 165982 200124
rect 166046 199918 166074 200124
rect 165756 199849 165812 199858
rect 165850 199912 165902 199918
rect 165850 199854 165902 199860
rect 165942 199912 165994 199918
rect 165942 199854 165994 199860
rect 166034 199912 166086 199918
rect 166034 199854 166086 199860
rect 166138 199764 166166 200124
rect 166092 199753 166166 199764
rect 166078 199744 166166 199753
rect 165804 199708 165856 199714
rect 165356 197334 165384 199679
rect 165678 199668 165752 199696
rect 165436 199640 165488 199646
rect 165436 199582 165488 199588
rect 165344 197328 165396 197334
rect 165250 197296 165306 197305
rect 165344 197270 165396 197276
rect 165250 197231 165306 197240
rect 165172 195946 165292 195974
rect 165264 191214 165292 195946
rect 165448 193214 165476 199582
rect 165528 199572 165580 199578
rect 165528 199514 165580 199520
rect 165540 198422 165568 199514
rect 165620 198552 165672 198558
rect 165620 198494 165672 198500
rect 165528 198416 165580 198422
rect 165528 198358 165580 198364
rect 165632 198150 165660 198494
rect 165724 198370 165752 199668
rect 165804 199650 165856 199656
rect 165988 199708 166040 199714
rect 166134 199736 166166 199744
rect 166230 199696 166258 200124
rect 166322 199782 166350 200124
rect 166414 199923 166442 200124
rect 166400 199914 166456 199923
rect 166506 199918 166534 200124
rect 166400 199849 166456 199858
rect 166494 199912 166546 199918
rect 166494 199854 166546 199860
rect 166310 199776 166362 199782
rect 166598 199764 166626 200124
rect 166690 199850 166718 200124
rect 166782 199923 166810 200124
rect 166768 199914 166824 199923
rect 166874 199918 166902 200124
rect 166678 199844 166730 199850
rect 166768 199849 166824 199858
rect 166862 199912 166914 199918
rect 166862 199854 166914 199860
rect 166678 199786 166730 199792
rect 166310 199718 166362 199724
rect 166552 199736 166626 199764
rect 166078 199679 166134 199688
rect 165988 199650 166040 199656
rect 166184 199668 166258 199696
rect 165816 198529 165844 199650
rect 165896 199640 165948 199646
rect 165896 199582 165948 199588
rect 165802 198520 165858 198529
rect 165802 198455 165858 198464
rect 165724 198342 165844 198370
rect 165712 198280 165764 198286
rect 165712 198222 165764 198228
rect 165620 198144 165672 198150
rect 165620 198086 165672 198092
rect 165724 198082 165752 198222
rect 165712 198076 165764 198082
rect 165712 198018 165764 198024
rect 165620 198008 165672 198014
rect 165620 197950 165672 197956
rect 165448 193186 165568 193214
rect 165252 191208 165304 191214
rect 165252 191150 165304 191156
rect 165068 191072 165120 191078
rect 165068 191014 165120 191020
rect 164792 191004 164844 191010
rect 164792 190946 164844 190952
rect 164804 154086 164832 190946
rect 164884 156800 164936 156806
rect 164884 156742 164936 156748
rect 164792 154080 164844 154086
rect 164792 154022 164844 154028
rect 164700 152788 164752 152794
rect 164700 152730 164752 152736
rect 164608 151632 164660 151638
rect 164608 151574 164660 151580
rect 164516 149796 164568 149802
rect 164516 149738 164568 149744
rect 164238 147112 164294 147121
rect 164238 147047 164294 147056
rect 164238 145752 164294 145761
rect 164238 145687 164294 145696
rect 163964 141636 164016 141642
rect 163964 141578 164016 141584
rect 164252 139890 164280 145687
rect 164896 139890 164924 156742
rect 165540 149666 165568 193186
rect 165632 191010 165660 197950
rect 165816 193214 165844 198342
rect 165908 195974 165936 199582
rect 166000 198014 166028 199650
rect 166080 199640 166132 199646
rect 166080 199582 166132 199588
rect 166092 198082 166120 199582
rect 166080 198076 166132 198082
rect 166080 198018 166132 198024
rect 165988 198008 166040 198014
rect 165988 197950 166040 197956
rect 165908 195946 166120 195974
rect 165816 193186 166028 193214
rect 166000 191400 166028 193186
rect 166092 191758 166120 195946
rect 166080 191752 166132 191758
rect 166080 191694 166132 191700
rect 166000 191372 166120 191400
rect 165712 191208 165764 191214
rect 165712 191150 165764 191156
rect 165620 191004 165672 191010
rect 165620 190946 165672 190952
rect 165528 149660 165580 149666
rect 165528 149602 165580 149608
rect 165724 146985 165752 191150
rect 165896 191072 165948 191078
rect 165896 191014 165948 191020
rect 165804 190936 165856 190942
rect 165804 190878 165856 190884
rect 165816 149870 165844 190878
rect 165908 154562 165936 191014
rect 166092 186314 166120 191372
rect 166184 190942 166212 199668
rect 166356 199572 166408 199578
rect 166356 199514 166408 199520
rect 166448 199572 166500 199578
rect 166448 199514 166500 199520
rect 166368 191214 166396 199514
rect 166460 198558 166488 199514
rect 166448 198552 166500 198558
rect 166448 198494 166500 198500
rect 166448 198076 166500 198082
rect 166448 198018 166500 198024
rect 166356 191208 166408 191214
rect 166356 191150 166408 191156
rect 166172 190936 166224 190942
rect 166172 190878 166224 190884
rect 166000 186286 166120 186314
rect 165896 154556 165948 154562
rect 165896 154498 165948 154504
rect 166000 154018 166028 186286
rect 166460 180794 166488 198018
rect 166552 191486 166580 199736
rect 166966 199730 166994 200124
rect 167058 199787 167086 200124
rect 166920 199702 166994 199730
rect 167044 199778 167100 199787
rect 167150 199782 167178 200124
rect 167242 199850 167270 200124
rect 167230 199844 167282 199850
rect 167230 199786 167282 199792
rect 167044 199713 167100 199722
rect 167138 199776 167190 199782
rect 167334 199730 167362 200124
rect 167426 199850 167454 200124
rect 167518 199889 167546 200124
rect 167610 199918 167638 200124
rect 167702 199918 167730 200124
rect 167794 199918 167822 200124
rect 167886 199918 167914 200124
rect 167598 199912 167650 199918
rect 167504 199880 167560 199889
rect 167414 199844 167466 199850
rect 167598 199854 167650 199860
rect 167690 199912 167742 199918
rect 167690 199854 167742 199860
rect 167782 199912 167834 199918
rect 167782 199854 167834 199860
rect 167874 199912 167926 199918
rect 167874 199854 167926 199860
rect 167504 199815 167560 199824
rect 167414 199786 167466 199792
rect 167978 199764 168006 200124
rect 168070 199918 168098 200124
rect 168162 199918 168190 200124
rect 168254 199923 168282 200124
rect 168058 199912 168110 199918
rect 168058 199854 168110 199860
rect 168150 199912 168202 199918
rect 168150 199854 168202 199860
rect 168240 199914 168296 199923
rect 168240 199849 168296 199858
rect 168104 199776 168156 199782
rect 167138 199718 167190 199724
rect 167288 199702 167362 199730
rect 167458 199744 167514 199753
rect 166632 199640 166684 199646
rect 166632 199582 166684 199588
rect 166644 196761 166672 199582
rect 166816 198552 166868 198558
rect 166816 198494 166868 198500
rect 166722 198112 166778 198121
rect 166722 198047 166778 198056
rect 166630 196752 166686 196761
rect 166630 196687 166686 196696
rect 166632 191684 166684 191690
rect 166632 191626 166684 191632
rect 166540 191480 166592 191486
rect 166540 191422 166592 191428
rect 166644 191214 166672 191626
rect 166632 191208 166684 191214
rect 166632 191150 166684 191156
rect 166736 191078 166764 198047
rect 166724 191072 166776 191078
rect 166724 191014 166776 191020
rect 166184 180766 166488 180794
rect 165988 154012 166040 154018
rect 165988 153954 166040 153960
rect 166184 153814 166212 180766
rect 166264 156528 166316 156534
rect 166264 156470 166316 156476
rect 166172 153808 166224 153814
rect 166172 153750 166224 153756
rect 165804 149864 165856 149870
rect 165804 149806 165856 149812
rect 165710 146976 165766 146985
rect 165710 146911 165766 146920
rect 165712 145920 165764 145926
rect 165712 145862 165764 145868
rect 165526 144800 165582 144809
rect 165526 144735 165582 144744
rect 165540 140162 165568 144735
rect 165494 140134 165568 140162
rect 163608 139862 163852 139890
rect 164252 139862 164404 139890
rect 164896 139862 164956 139890
rect 165494 139876 165522 140134
rect 165724 139890 165752 145862
rect 166276 139890 166304 156470
rect 166828 145654 166856 198494
rect 166920 197198 166948 199702
rect 167000 199640 167052 199646
rect 167000 199582 167052 199588
rect 167184 199640 167236 199646
rect 167184 199582 167236 199588
rect 167012 197441 167040 199582
rect 167092 199572 167144 199578
rect 167092 199514 167144 199520
rect 167104 197878 167132 199514
rect 167092 197872 167144 197878
rect 167092 197814 167144 197820
rect 166998 197432 167054 197441
rect 166998 197367 167054 197376
rect 166908 197192 166960 197198
rect 166908 197134 166960 197140
rect 167196 196926 167224 199582
rect 167184 196920 167236 196926
rect 167184 196862 167236 196868
rect 166908 191752 166960 191758
rect 166908 191694 166960 191700
rect 166920 153950 166948 191694
rect 167184 191412 167236 191418
rect 167184 191354 167236 191360
rect 167000 191004 167052 191010
rect 167000 190946 167052 190952
rect 166908 153944 166960 153950
rect 166908 153886 166960 153892
rect 167012 150142 167040 190946
rect 167092 190936 167144 190942
rect 167092 190878 167144 190884
rect 167000 150136 167052 150142
rect 167000 150078 167052 150084
rect 167104 149841 167132 190878
rect 167196 156874 167224 191354
rect 167288 190890 167316 199702
rect 167978 199736 168052 199764
rect 167458 199679 167514 199688
rect 167552 199708 167604 199714
rect 167368 199640 167420 199646
rect 167368 199582 167420 199588
rect 167380 191826 167408 199582
rect 167472 198694 167500 199679
rect 167552 199650 167604 199656
rect 167644 199708 167696 199714
rect 167644 199650 167696 199656
rect 167736 199708 167788 199714
rect 167736 199650 167788 199656
rect 167460 198688 167512 198694
rect 167460 198630 167512 198636
rect 167460 198280 167512 198286
rect 167460 198222 167512 198228
rect 167472 198014 167500 198222
rect 167460 198008 167512 198014
rect 167460 197950 167512 197956
rect 167460 197872 167512 197878
rect 167460 197814 167512 197820
rect 167368 191820 167420 191826
rect 167368 191762 167420 191768
rect 167288 190862 167408 190890
rect 167472 190874 167500 197814
rect 167564 191418 167592 199650
rect 167552 191412 167604 191418
rect 167552 191354 167604 191360
rect 167380 186402 167408 190862
rect 167460 190868 167512 190874
rect 167460 190810 167512 190816
rect 167656 190806 167684 199650
rect 167748 196382 167776 199650
rect 167828 199640 167880 199646
rect 167828 199582 167880 199588
rect 167918 199608 167974 199617
rect 167736 196376 167788 196382
rect 167736 196318 167788 196324
rect 167840 191010 167868 199582
rect 167918 199543 167974 199552
rect 167932 199510 167960 199543
rect 167920 199504 167972 199510
rect 167920 199446 167972 199452
rect 167920 198620 167972 198626
rect 167920 198562 167972 198568
rect 167932 197062 167960 198562
rect 167920 197056 167972 197062
rect 167920 196998 167972 197004
rect 168024 194594 168052 199736
rect 168104 199718 168156 199724
rect 168194 199744 168250 199753
rect 167932 194566 168052 194594
rect 167828 191004 167880 191010
rect 167828 190946 167880 190952
rect 167644 190800 167696 190806
rect 167644 190742 167696 190748
rect 167932 190466 167960 194566
rect 168116 193361 168144 199718
rect 168194 199679 168250 199688
rect 168102 193352 168158 193361
rect 168102 193287 168158 193296
rect 168208 191834 168236 199679
rect 168346 199628 168374 200124
rect 168438 199850 168466 200124
rect 168530 199918 168558 200124
rect 168518 199912 168570 199918
rect 168518 199854 168570 199860
rect 168426 199844 168478 199850
rect 168426 199786 168478 199792
rect 168472 199708 168524 199714
rect 168622 199696 168650 200124
rect 168714 199764 168742 200124
rect 168806 199918 168834 200124
rect 168898 199918 168926 200124
rect 168794 199912 168846 199918
rect 168794 199854 168846 199860
rect 168886 199912 168938 199918
rect 168990 199889 169018 200124
rect 169082 199918 169110 200124
rect 169174 199918 169202 200124
rect 169070 199912 169122 199918
rect 168886 199854 168938 199860
rect 168976 199880 169032 199889
rect 169070 199854 169122 199860
rect 169162 199912 169214 199918
rect 169162 199854 169214 199860
rect 168976 199815 169032 199824
rect 169024 199776 169076 199782
rect 168714 199736 168788 199764
rect 168622 199668 168696 199696
rect 168472 199650 168524 199656
rect 168346 199600 168420 199628
rect 168288 199504 168340 199510
rect 168288 199446 168340 199452
rect 168300 197674 168328 199446
rect 168392 198966 168420 199600
rect 168380 198960 168432 198966
rect 168380 198902 168432 198908
rect 168288 197668 168340 197674
rect 168288 197610 168340 197616
rect 168484 194410 168512 199650
rect 168564 199572 168616 199578
rect 168564 199514 168616 199520
rect 168472 194404 168524 194410
rect 168472 194346 168524 194352
rect 168208 191806 168328 191834
rect 168300 190942 168328 191806
rect 168576 191758 168604 199514
rect 168668 194546 168696 199668
rect 168760 195945 168788 199736
rect 168930 199744 168986 199753
rect 168840 199708 168892 199714
rect 169266 199764 169294 200124
rect 169024 199718 169076 199724
rect 169220 199736 169294 199764
rect 169358 199764 169386 200124
rect 169450 199923 169478 200124
rect 169436 199914 169492 199923
rect 169542 199918 169570 200124
rect 169634 199923 169662 200124
rect 169436 199849 169492 199858
rect 169530 199912 169582 199918
rect 169530 199854 169582 199860
rect 169620 199914 169676 199923
rect 169726 199918 169754 200124
rect 169818 199918 169846 200124
rect 169910 199918 169938 200124
rect 169620 199849 169676 199858
rect 169714 199912 169766 199918
rect 169714 199854 169766 199860
rect 169806 199912 169858 199918
rect 169806 199854 169858 199860
rect 169898 199912 169950 199918
rect 169898 199854 169950 199860
rect 169484 199776 169536 199782
rect 169358 199736 169432 199764
rect 168930 199679 168986 199688
rect 168840 199650 168892 199656
rect 168746 195936 168802 195945
rect 168746 195871 168802 195880
rect 168656 194540 168708 194546
rect 168656 194482 168708 194488
rect 168656 194404 168708 194410
rect 168656 194346 168708 194352
rect 168564 191752 168616 191758
rect 168564 191694 168616 191700
rect 168564 191004 168616 191010
rect 168564 190946 168616 190952
rect 168288 190936 168340 190942
rect 168288 190878 168340 190884
rect 167920 190460 167972 190466
rect 167920 190402 167972 190408
rect 168472 187332 168524 187338
rect 168472 187274 168524 187280
rect 167288 186374 167408 186402
rect 167288 157010 167316 186374
rect 167276 157004 167328 157010
rect 167276 156946 167328 156952
rect 167184 156868 167236 156874
rect 167184 156810 167236 156816
rect 168484 149977 168512 187274
rect 168576 157078 168604 190946
rect 168564 157072 168616 157078
rect 168564 157014 168616 157020
rect 168668 156942 168696 194346
rect 168852 194313 168880 199650
rect 168838 194304 168894 194313
rect 168838 194239 168894 194248
rect 168944 191010 168972 199679
rect 168932 191004 168984 191010
rect 168932 190946 168984 190952
rect 169036 187406 169064 199718
rect 169116 199708 169168 199714
rect 169116 199650 169168 199656
rect 169128 194478 169156 199650
rect 169116 194472 169168 194478
rect 169116 194414 169168 194420
rect 169024 187400 169076 187406
rect 169024 187342 169076 187348
rect 169220 186314 169248 199736
rect 169300 199640 169352 199646
rect 169300 199582 169352 199588
rect 169312 199073 169340 199582
rect 169298 199064 169354 199073
rect 169298 198999 169354 199008
rect 169300 198008 169352 198014
rect 169300 197950 169352 197956
rect 169312 197849 169340 197950
rect 169298 197840 169354 197849
rect 169298 197775 169354 197784
rect 169404 196353 169432 199736
rect 169852 199776 169904 199782
rect 169484 199718 169536 199724
rect 169574 199744 169630 199753
rect 169390 196344 169446 196353
rect 169390 196279 169446 196288
rect 168760 186286 169248 186314
rect 168656 156936 168708 156942
rect 168656 156878 168708 156884
rect 168760 156641 168788 186286
rect 168746 156632 168802 156641
rect 168746 156567 168802 156576
rect 168470 149968 168526 149977
rect 168470 149903 168526 149912
rect 167090 149832 167146 149841
rect 167090 149767 167146 149776
rect 166816 145648 166868 145654
rect 166816 145590 166868 145596
rect 169116 144560 169168 144566
rect 169116 144502 169168 144508
rect 168012 144492 168064 144498
rect 168012 144434 168064 144440
rect 167458 141808 167514 141817
rect 167458 141743 167514 141752
rect 167472 139890 167500 141743
rect 168024 139890 168052 144434
rect 168288 143132 168340 143138
rect 168288 143074 168340 143080
rect 168300 140162 168328 143074
rect 165724 139862 166060 139890
rect 166276 139862 166612 139890
rect 167164 139862 167500 139890
rect 167716 139862 168052 139890
rect 168254 140134 168328 140162
rect 168254 139876 168282 140134
rect 169128 139890 169156 144502
rect 169300 141500 169352 141506
rect 169300 141442 169352 141448
rect 168820 139862 169156 139890
rect 169312 139754 169340 141442
rect 169312 139726 169372 139754
rect 169496 139369 169524 199718
rect 170002 199764 170030 200124
rect 170094 199923 170122 200124
rect 170080 199914 170136 199923
rect 170186 199918 170214 200124
rect 170080 199849 170136 199858
rect 170174 199912 170226 199918
rect 170174 199854 170226 199860
rect 170278 199764 170306 200124
rect 169852 199718 169904 199724
rect 169956 199736 170030 199764
rect 170126 199744 170182 199753
rect 169574 199679 169630 199688
rect 169668 199708 169720 199714
rect 169588 195158 169616 199679
rect 169668 199650 169720 199656
rect 169760 199708 169812 199714
rect 169760 199650 169812 199656
rect 169680 197985 169708 199650
rect 169666 197976 169722 197985
rect 169666 197911 169722 197920
rect 169666 196480 169722 196489
rect 169666 196415 169722 196424
rect 169576 195152 169628 195158
rect 169576 195094 169628 195100
rect 169680 187338 169708 196415
rect 169772 193214 169800 199650
rect 169864 196722 169892 199718
rect 169956 198626 169984 199736
rect 170126 199679 170182 199688
rect 170232 199736 170306 199764
rect 170140 199170 170168 199679
rect 170128 199164 170180 199170
rect 170128 199106 170180 199112
rect 170232 198937 170260 199736
rect 170370 199730 170398 200124
rect 170462 199850 170490 200124
rect 170450 199844 170502 199850
rect 170450 199786 170502 199792
rect 170554 199730 170582 200124
rect 170646 199923 170674 200124
rect 170632 199914 170688 199923
rect 170632 199849 170688 199858
rect 170738 199850 170766 200124
rect 170830 199850 170858 200124
rect 170922 199850 170950 200124
rect 171014 199918 171042 200124
rect 171002 199912 171054 199918
rect 171002 199854 171054 199860
rect 170726 199844 170778 199850
rect 170726 199786 170778 199792
rect 170818 199844 170870 199850
rect 170818 199786 170870 199792
rect 170910 199844 170962 199850
rect 170910 199786 170962 199792
rect 171106 199764 171134 200124
rect 171198 199918 171226 200124
rect 171290 199923 171318 200124
rect 171186 199912 171238 199918
rect 171186 199854 171238 199860
rect 171276 199914 171332 199923
rect 171382 199918 171410 200124
rect 171474 199918 171502 200124
rect 171566 199918 171594 200124
rect 171658 199918 171686 200124
rect 171276 199849 171332 199858
rect 171370 199912 171422 199918
rect 171370 199854 171422 199860
rect 171462 199912 171514 199918
rect 171462 199854 171514 199860
rect 171554 199912 171606 199918
rect 171554 199854 171606 199860
rect 171646 199912 171698 199918
rect 171646 199854 171698 199860
rect 171750 199764 171778 200124
rect 171842 199923 171870 200124
rect 171828 199914 171884 199923
rect 171934 199918 171962 200124
rect 171828 199849 171884 199858
rect 171922 199912 171974 199918
rect 171922 199854 171974 199860
rect 172026 199764 172054 200124
rect 172118 199889 172146 200124
rect 172210 199918 172238 200124
rect 172302 199918 172330 200124
rect 172394 199923 172422 200124
rect 172198 199912 172250 199918
rect 172104 199880 172160 199889
rect 172198 199854 172250 199860
rect 172290 199912 172342 199918
rect 172290 199854 172342 199860
rect 172380 199914 172436 199923
rect 172380 199849 172436 199858
rect 172104 199815 172160 199824
rect 171060 199736 171134 199764
rect 171704 199736 171778 199764
rect 171980 199736 172054 199764
rect 172336 199776 172388 199782
rect 170370 199702 170444 199730
rect 170554 199702 170628 199730
rect 170312 199640 170364 199646
rect 170312 199582 170364 199588
rect 170218 198928 170274 198937
rect 170218 198863 170274 198872
rect 169944 198620 169996 198626
rect 169944 198562 169996 198568
rect 169852 196716 169904 196722
rect 169852 196658 169904 196664
rect 170220 196716 170272 196722
rect 170220 196658 170272 196664
rect 169772 193186 170076 193214
rect 169852 191004 169904 191010
rect 170048 190992 170076 193186
rect 170232 192914 170260 196658
rect 170324 193118 170352 199582
rect 170416 198064 170444 199702
rect 170496 199640 170548 199646
rect 170496 199582 170548 199588
rect 170508 198257 170536 199582
rect 170600 198286 170628 199702
rect 170772 199640 170824 199646
rect 170772 199582 170824 199588
rect 170956 199640 171008 199646
rect 170956 199582 171008 199588
rect 170680 199572 170732 199578
rect 170680 199514 170732 199520
rect 170588 198280 170640 198286
rect 170494 198248 170550 198257
rect 170588 198222 170640 198228
rect 170494 198183 170550 198192
rect 170416 198036 170536 198064
rect 170404 197192 170456 197198
rect 170404 197134 170456 197140
rect 170416 193225 170444 197134
rect 170402 193216 170458 193225
rect 170402 193151 170458 193160
rect 170312 193112 170364 193118
rect 170312 193054 170364 193060
rect 170220 192908 170272 192914
rect 170220 192850 170272 192856
rect 170508 191834 170536 198036
rect 170588 196852 170640 196858
rect 170588 196794 170640 196800
rect 170600 196722 170628 196794
rect 170588 196716 170640 196722
rect 170588 196658 170640 196664
rect 170586 196480 170642 196489
rect 170586 196415 170642 196424
rect 170324 191806 170536 191834
rect 170048 190964 170168 190992
rect 169852 190946 169904 190952
rect 169760 190936 169812 190942
rect 169760 190878 169812 190884
rect 169668 187332 169720 187338
rect 169668 187274 169720 187280
rect 169772 140321 169800 190878
rect 169864 147529 169892 190946
rect 169944 188420 169996 188426
rect 169944 188362 169996 188368
rect 169850 147520 169906 147529
rect 169850 147455 169906 147464
rect 169852 145988 169904 145994
rect 169852 145930 169904 145936
rect 169864 140690 169892 145930
rect 169852 140684 169904 140690
rect 169852 140626 169904 140632
rect 169956 140457 169984 188362
rect 170140 183554 170168 190964
rect 170324 188426 170352 191806
rect 170600 191010 170628 196415
rect 170692 194138 170720 199514
rect 170784 198529 170812 199582
rect 170864 199504 170916 199510
rect 170864 199446 170916 199452
rect 170770 198520 170826 198529
rect 170770 198455 170826 198464
rect 170772 197940 170824 197946
rect 170772 197882 170824 197888
rect 170680 194132 170732 194138
rect 170680 194074 170732 194080
rect 170588 191004 170640 191010
rect 170588 190946 170640 190952
rect 170312 188420 170364 188426
rect 170312 188362 170364 188368
rect 170784 186314 170812 197882
rect 170876 190942 170904 199446
rect 170968 198665 170996 199582
rect 170954 198656 171010 198665
rect 170954 198591 171010 198600
rect 171060 198506 171088 199736
rect 171416 199708 171468 199714
rect 171416 199650 171468 199656
rect 171508 199708 171560 199714
rect 171508 199650 171560 199656
rect 171140 199640 171192 199646
rect 171322 199608 171378 199617
rect 171140 199582 171192 199588
rect 170968 198478 171088 198506
rect 170968 198257 170996 198478
rect 171152 198393 171180 199582
rect 171244 199566 171322 199594
rect 171138 198384 171194 198393
rect 171048 198348 171100 198354
rect 171138 198319 171194 198328
rect 171048 198290 171100 198296
rect 170954 198248 171010 198257
rect 170954 198183 171010 198192
rect 171060 197198 171088 198290
rect 171140 198212 171192 198218
rect 171140 198154 171192 198160
rect 171152 197946 171180 198154
rect 171140 197940 171192 197946
rect 171140 197882 171192 197888
rect 171048 197192 171100 197198
rect 171048 197134 171100 197140
rect 171244 196858 171272 199566
rect 171322 199543 171378 199552
rect 171324 199504 171376 199510
rect 171324 199446 171376 199452
rect 171336 198082 171364 199446
rect 171428 198734 171456 199650
rect 171520 199424 171548 199650
rect 171520 199396 171640 199424
rect 171428 198706 171548 198734
rect 171520 198608 171548 198706
rect 171428 198580 171548 198608
rect 171324 198076 171376 198082
rect 171324 198018 171376 198024
rect 171324 197260 171376 197266
rect 171324 197202 171376 197208
rect 171232 196852 171284 196858
rect 171232 196794 171284 196800
rect 171336 196586 171364 197202
rect 171324 196580 171376 196586
rect 171324 196522 171376 196528
rect 171140 191004 171192 191010
rect 171140 190946 171192 190952
rect 170864 190936 170916 190942
rect 170864 190878 170916 190884
rect 170784 186286 170904 186314
rect 170048 183526 170168 183554
rect 170048 148782 170076 183526
rect 170036 148776 170088 148782
rect 170036 148718 170088 148724
rect 170876 147393 170904 186286
rect 170862 147384 170918 147393
rect 170862 147319 170918 147328
rect 170588 144696 170640 144702
rect 170588 144638 170640 144644
rect 170220 141772 170272 141778
rect 170220 141714 170272 141720
rect 169942 140448 169998 140457
rect 169942 140383 169998 140392
rect 169758 140312 169814 140321
rect 169758 140247 169814 140256
rect 170232 139890 170260 141714
rect 170600 139890 170628 144638
rect 170680 140684 170732 140690
rect 170680 140626 170732 140632
rect 169924 139862 170260 139890
rect 170476 139862 170628 139890
rect 170692 139890 170720 140626
rect 171152 140593 171180 190946
rect 171232 190936 171284 190942
rect 171232 190878 171284 190884
rect 171244 148646 171272 190878
rect 171428 186314 171456 198580
rect 171612 198506 171640 199396
rect 171704 198734 171732 199736
rect 171874 199608 171930 199617
rect 171874 199543 171930 199552
rect 171704 198706 171824 198734
rect 171796 198506 171824 198706
rect 171520 198478 171640 198506
rect 171704 198478 171824 198506
rect 171520 192982 171548 198478
rect 171600 198416 171652 198422
rect 171600 198358 171652 198364
rect 171612 196994 171640 198358
rect 171600 196988 171652 196994
rect 171600 196930 171652 196936
rect 171600 196852 171652 196858
rect 171600 196794 171652 196800
rect 171612 193050 171640 196794
rect 171600 193044 171652 193050
rect 171600 192986 171652 192992
rect 171508 192976 171560 192982
rect 171508 192918 171560 192924
rect 171336 186286 171456 186314
rect 171232 148640 171284 148646
rect 171232 148582 171284 148588
rect 171336 148510 171364 186286
rect 171704 180794 171732 198478
rect 171888 198064 171916 199543
rect 171796 198036 171916 198064
rect 171796 192681 171824 198036
rect 171876 195968 171928 195974
rect 171876 195910 171928 195916
rect 171888 194886 171916 195910
rect 171876 194880 171928 194886
rect 171876 194822 171928 194828
rect 171782 192672 171838 192681
rect 171782 192607 171838 192616
rect 171980 191010 172008 199736
rect 172486 199764 172514 200124
rect 172578 199923 172606 200124
rect 172564 199914 172620 199923
rect 172670 199918 172698 200124
rect 172762 199923 172790 200124
rect 172564 199849 172620 199858
rect 172658 199912 172710 199918
rect 172658 199854 172710 199860
rect 172748 199914 172804 199923
rect 172854 199918 172882 200124
rect 172748 199849 172804 199858
rect 172842 199912 172894 199918
rect 172842 199854 172894 199860
rect 172946 199764 172974 200124
rect 172486 199736 172560 199764
rect 172336 199718 172388 199724
rect 172244 199708 172296 199714
rect 172244 199650 172296 199656
rect 172060 199640 172112 199646
rect 172060 199582 172112 199588
rect 172072 198422 172100 199582
rect 172060 198416 172112 198422
rect 172060 198358 172112 198364
rect 172060 198144 172112 198150
rect 172060 198086 172112 198092
rect 172072 197266 172100 198086
rect 172152 197804 172204 197810
rect 172152 197746 172204 197752
rect 172060 197260 172112 197266
rect 172060 197202 172112 197208
rect 171968 191004 172020 191010
rect 171968 190946 172020 190952
rect 172164 186314 172192 197746
rect 172256 190942 172284 199650
rect 172348 198150 172376 199718
rect 172426 199608 172482 199617
rect 172426 199543 172482 199552
rect 172440 198354 172468 199543
rect 172532 198801 172560 199736
rect 172794 199744 172850 199753
rect 172704 199708 172756 199714
rect 172794 199679 172850 199688
rect 172900 199736 172974 199764
rect 172704 199650 172756 199656
rect 172612 199640 172664 199646
rect 172612 199582 172664 199588
rect 172518 198792 172574 198801
rect 172518 198727 172574 198736
rect 172520 198552 172572 198558
rect 172520 198494 172572 198500
rect 172428 198348 172480 198354
rect 172428 198290 172480 198296
rect 172336 198144 172388 198150
rect 172336 198086 172388 198092
rect 172336 197940 172388 197946
rect 172336 197882 172388 197888
rect 172348 194954 172376 197882
rect 172426 197840 172482 197849
rect 172532 197810 172560 198494
rect 172624 197946 172652 199582
rect 172612 197940 172664 197946
rect 172612 197882 172664 197888
rect 172426 197775 172482 197784
rect 172520 197804 172572 197810
rect 172440 197470 172468 197775
rect 172520 197746 172572 197752
rect 172428 197464 172480 197470
rect 172428 197406 172480 197412
rect 172518 197432 172574 197441
rect 172518 197367 172574 197376
rect 172532 196858 172560 197367
rect 172520 196852 172572 196858
rect 172520 196794 172572 196800
rect 172612 195016 172664 195022
rect 172612 194958 172664 194964
rect 172336 194948 172388 194954
rect 172336 194890 172388 194896
rect 172244 190936 172296 190942
rect 172244 190878 172296 190884
rect 172520 189644 172572 189650
rect 172520 189586 172572 189592
rect 172164 186286 172284 186314
rect 171428 180766 171732 180794
rect 171428 148578 171456 180766
rect 172256 150414 172284 186286
rect 172244 150408 172296 150414
rect 172244 150350 172296 150356
rect 172532 149025 172560 189586
rect 172624 159594 172652 194958
rect 172716 192846 172744 199650
rect 172808 198218 172836 199679
rect 172796 198212 172848 198218
rect 172796 198154 172848 198160
rect 172900 198064 172928 199736
rect 173038 199424 173066 200124
rect 173130 199923 173158 200124
rect 173116 199914 173172 199923
rect 173116 199849 173172 199858
rect 173222 199764 173250 200124
rect 173314 199889 173342 200124
rect 173300 199880 173356 199889
rect 173300 199815 173356 199824
rect 173406 199764 173434 200124
rect 172808 198036 172928 198064
rect 172992 199396 173066 199424
rect 173176 199736 173250 199764
rect 173360 199736 173434 199764
rect 172808 194070 172836 198036
rect 172888 197940 172940 197946
rect 172888 197882 172940 197888
rect 172796 194064 172848 194070
rect 172796 194006 172848 194012
rect 172704 192840 172756 192846
rect 172704 192782 172756 192788
rect 172704 191004 172756 191010
rect 172704 190946 172756 190952
rect 172612 159588 172664 159594
rect 172612 159530 172664 159536
rect 172518 149016 172574 149025
rect 172518 148951 172574 148960
rect 171416 148572 171468 148578
rect 171416 148514 171468 148520
rect 171324 148504 171376 148510
rect 172716 148481 172744 190946
rect 172796 159724 172848 159730
rect 172796 159666 172848 159672
rect 171324 148446 171376 148452
rect 172702 148472 172758 148481
rect 172702 148407 172758 148416
rect 172428 144628 172480 144634
rect 172428 144570 172480 144576
rect 171876 141704 171928 141710
rect 171876 141646 171928 141652
rect 171138 140584 171194 140593
rect 171138 140519 171194 140528
rect 171888 139890 171916 141646
rect 172440 139890 172468 144570
rect 172808 139890 172836 159666
rect 172900 148209 172928 197882
rect 172992 195022 173020 199396
rect 173072 197736 173124 197742
rect 173072 197678 173124 197684
rect 172980 195016 173032 195022
rect 172980 194958 173032 194964
rect 173084 186314 173112 197678
rect 173176 192778 173204 199736
rect 173360 199628 173388 199736
rect 173498 199696 173526 200124
rect 173590 199918 173618 200124
rect 173578 199912 173630 199918
rect 173578 199854 173630 199860
rect 173314 199600 173388 199628
rect 173452 199668 173526 199696
rect 173314 199560 173342 199600
rect 173314 199532 173388 199560
rect 173256 195492 173308 195498
rect 173256 195434 173308 195440
rect 173164 192772 173216 192778
rect 173164 192714 173216 192720
rect 173268 189530 173296 195434
rect 173360 189650 173388 199532
rect 173452 194177 173480 199668
rect 173682 199628 173710 200124
rect 173774 199889 173802 200124
rect 173760 199880 173816 199889
rect 173760 199815 173816 199824
rect 173866 199696 173894 200124
rect 173958 199764 173986 200124
rect 174050 199918 174078 200124
rect 174142 199923 174170 200124
rect 174038 199912 174090 199918
rect 174038 199854 174090 199860
rect 174128 199914 174184 199923
rect 174128 199849 174184 199858
rect 174084 199776 174136 199782
rect 173958 199736 174032 199764
rect 173866 199668 173940 199696
rect 173682 199600 173756 199628
rect 173530 199064 173586 199073
rect 173530 198999 173586 199008
rect 173544 194410 173572 198999
rect 173622 198792 173678 198801
rect 173622 198727 173678 198736
rect 173636 197849 173664 198727
rect 173622 197840 173678 197849
rect 173622 197775 173678 197784
rect 173532 194404 173584 194410
rect 173532 194346 173584 194352
rect 173438 194168 173494 194177
rect 173438 194103 173494 194112
rect 173728 193214 173756 199600
rect 173806 199608 173862 199617
rect 173806 199543 173808 199552
rect 173860 199543 173862 199552
rect 173808 199514 173860 199520
rect 173912 198694 173940 199668
rect 173900 198688 173952 198694
rect 173900 198630 173952 198636
rect 173808 197532 173860 197538
rect 173808 197474 173860 197480
rect 173820 195974 173848 197474
rect 174004 197470 174032 199736
rect 174234 199764 174262 200124
rect 174326 199923 174354 200124
rect 174312 199914 174368 199923
rect 174312 199849 174368 199858
rect 174418 199764 174446 200124
rect 174084 199718 174136 199724
rect 174188 199736 174262 199764
rect 174372 199736 174446 199764
rect 173992 197464 174044 197470
rect 173992 197406 174044 197412
rect 173808 195968 173860 195974
rect 173808 195910 173860 195916
rect 173806 195664 173862 195673
rect 173806 195599 173862 195608
rect 173636 193186 173756 193214
rect 173636 191010 173664 193186
rect 173624 191004 173676 191010
rect 173624 190946 173676 190952
rect 173348 189644 173400 189650
rect 173348 189586 173400 189592
rect 173268 189502 173388 189530
rect 173084 186286 173296 186314
rect 173268 150346 173296 186286
rect 173360 151814 173388 189502
rect 173360 151786 173664 151814
rect 173256 150340 173308 150346
rect 173256 150282 173308 150288
rect 172886 148200 172942 148209
rect 172886 148135 172942 148144
rect 173532 143200 173584 143206
rect 173532 143142 173584 143148
rect 173544 139890 173572 143142
rect 170692 139862 171028 139890
rect 171580 139862 171916 139890
rect 172132 139862 172468 139890
rect 172684 139862 172836 139890
rect 173236 139862 173572 139890
rect 173636 139369 173664 151786
rect 173820 148714 173848 195599
rect 174096 194698 174124 199718
rect 174004 194670 174124 194698
rect 174004 193594 174032 194670
rect 174188 194594 174216 199736
rect 174372 199617 174400 199736
rect 174510 199628 174538 200124
rect 174602 199918 174630 200124
rect 174694 199918 174722 200124
rect 174590 199912 174642 199918
rect 174590 199854 174642 199860
rect 174682 199912 174734 199918
rect 174786 199889 174814 200124
rect 174878 199918 174906 200124
rect 174866 199912 174918 199918
rect 174682 199854 174734 199860
rect 174772 199880 174828 199889
rect 174970 199889 174998 200124
rect 174866 199854 174918 199860
rect 174956 199880 175012 199889
rect 174772 199815 174828 199824
rect 174956 199815 175012 199824
rect 175062 199764 175090 200124
rect 175154 199923 175182 200124
rect 175140 199914 175196 199923
rect 175246 199918 175274 200124
rect 175140 199849 175196 199858
rect 175234 199912 175286 199918
rect 175234 199854 175286 199860
rect 174726 199744 174782 199753
rect 174636 199708 174688 199714
rect 174726 199679 174782 199688
rect 175016 199736 175090 199764
rect 175188 199776 175240 199782
rect 174636 199650 174688 199656
rect 174358 199608 174414 199617
rect 174358 199543 174414 199552
rect 174464 199600 174538 199628
rect 174358 199472 174414 199481
rect 174096 194566 174216 194594
rect 174280 199430 174358 199458
rect 173992 193588 174044 193594
rect 173992 193530 174044 193536
rect 173900 191684 173952 191690
rect 173900 191626 173952 191632
rect 173808 148708 173860 148714
rect 173808 148650 173860 148656
rect 173808 144764 173860 144770
rect 173808 144706 173860 144712
rect 173820 140162 173848 144706
rect 173912 140622 173940 191626
rect 173992 191004 174044 191010
rect 173992 190946 174044 190952
rect 174004 148442 174032 190946
rect 174096 151094 174124 194566
rect 174280 194002 174308 199430
rect 174358 199407 174414 199416
rect 174358 198928 174414 198937
rect 174358 198863 174414 198872
rect 174372 198558 174400 198863
rect 174360 198552 174412 198558
rect 174360 198494 174412 198500
rect 174360 195764 174412 195770
rect 174360 195706 174412 195712
rect 174268 193996 174320 194002
rect 174268 193938 174320 193944
rect 174176 191412 174228 191418
rect 174176 191354 174228 191360
rect 174188 151230 174216 191354
rect 174372 186314 174400 195706
rect 174464 191010 174492 199600
rect 174648 199481 174676 199650
rect 174634 199472 174690 199481
rect 174634 199407 174690 199416
rect 174542 198928 174598 198937
rect 174542 198863 174598 198872
rect 174556 194342 174584 198863
rect 174636 197872 174688 197878
rect 174636 197814 174688 197820
rect 174544 194336 174596 194342
rect 174544 194278 174596 194284
rect 174544 193928 174596 193934
rect 174544 193870 174596 193876
rect 174556 193798 174584 193870
rect 174544 193792 174596 193798
rect 174544 193734 174596 193740
rect 174648 191162 174676 197814
rect 174740 191418 174768 199679
rect 174912 199572 174964 199578
rect 174912 199514 174964 199520
rect 174924 198937 174952 199514
rect 174910 198928 174966 198937
rect 174910 198863 174966 198872
rect 175016 198744 175044 199736
rect 175338 199764 175366 200124
rect 175430 199918 175458 200124
rect 175522 199918 175550 200124
rect 175418 199912 175470 199918
rect 175418 199854 175470 199860
rect 175510 199912 175562 199918
rect 175510 199854 175562 199860
rect 175338 199736 175412 199764
rect 175188 199718 175240 199724
rect 175096 199640 175148 199646
rect 175096 199582 175148 199588
rect 174924 198716 175044 198744
rect 174820 198348 174872 198354
rect 174820 198290 174872 198296
rect 174832 192438 174860 198290
rect 174820 192432 174872 192438
rect 174820 192374 174872 192380
rect 174924 191690 174952 198716
rect 175108 197354 175136 199582
rect 175016 197326 175136 197354
rect 175016 195838 175044 197326
rect 175004 195832 175056 195838
rect 175004 195774 175056 195780
rect 175200 195673 175228 199718
rect 175280 199504 175332 199510
rect 175280 199446 175332 199452
rect 175292 198393 175320 199446
rect 175278 198384 175334 198393
rect 175278 198319 175334 198328
rect 175186 195664 175242 195673
rect 175186 195599 175242 195608
rect 175280 193792 175332 193798
rect 175280 193734 175332 193740
rect 175096 191752 175148 191758
rect 175096 191694 175148 191700
rect 174912 191684 174964 191690
rect 174912 191626 174964 191632
rect 174728 191412 174780 191418
rect 174728 191354 174780 191360
rect 175004 191412 175056 191418
rect 175004 191354 175056 191360
rect 174648 191134 174952 191162
rect 174452 191004 174504 191010
rect 174452 190946 174504 190952
rect 174372 186286 174860 186314
rect 174832 180794 174860 186286
rect 174740 180766 174860 180794
rect 174176 151224 174228 151230
rect 174176 151166 174228 151172
rect 174084 151088 174136 151094
rect 174084 151030 174136 151036
rect 173992 148436 174044 148442
rect 173992 148378 174044 148384
rect 174740 147558 174768 180766
rect 174728 147552 174780 147558
rect 174728 147494 174780 147500
rect 174924 146946 174952 191134
rect 175016 190806 175044 191354
rect 175108 190874 175136 191694
rect 175096 190868 175148 190874
rect 175096 190810 175148 190816
rect 175004 190800 175056 190806
rect 175004 190742 175056 190748
rect 174912 146940 174964 146946
rect 174912 146882 174964 146888
rect 173992 146056 174044 146062
rect 173992 145998 174044 146004
rect 173900 140616 173952 140622
rect 173900 140558 173952 140564
rect 173774 140134 173848 140162
rect 173774 139876 173802 140134
rect 174004 139890 174032 145998
rect 175292 145897 175320 193734
rect 175384 188630 175412 199736
rect 175614 199730 175642 200124
rect 175706 199923 175734 200124
rect 175692 199914 175748 199923
rect 175692 199849 175748 199858
rect 175798 199764 175826 200124
rect 175890 199918 175918 200124
rect 175878 199912 175930 199918
rect 175878 199854 175930 199860
rect 175982 199764 176010 200124
rect 176074 199918 176102 200124
rect 176062 199912 176114 199918
rect 176062 199854 176114 199860
rect 176166 199764 176194 200124
rect 176258 199918 176286 200124
rect 176350 199918 176378 200124
rect 176246 199912 176298 199918
rect 176246 199854 176298 199860
rect 176338 199912 176390 199918
rect 176442 199889 176470 200124
rect 176338 199854 176390 199860
rect 176428 199880 176484 199889
rect 176428 199815 176484 199824
rect 175798 199736 175872 199764
rect 175982 199736 176056 199764
rect 175464 199708 175516 199714
rect 175464 199650 175516 199656
rect 175568 199702 175642 199730
rect 175476 194274 175504 199650
rect 175464 194268 175516 194274
rect 175464 194210 175516 194216
rect 175568 191162 175596 199702
rect 175740 199640 175792 199646
rect 175740 199582 175792 199588
rect 175646 198792 175702 198801
rect 175646 198727 175702 198736
rect 175660 198422 175688 198727
rect 175648 198416 175700 198422
rect 175648 198358 175700 198364
rect 175752 193798 175780 199582
rect 175844 199073 175872 199736
rect 175924 199640 175976 199646
rect 175924 199582 175976 199588
rect 175830 199064 175886 199073
rect 175830 198999 175886 199008
rect 175936 198801 175964 199582
rect 175922 198792 175978 198801
rect 175922 198727 175978 198736
rect 175740 193792 175792 193798
rect 175740 193734 175792 193740
rect 175476 191134 175596 191162
rect 175372 188624 175424 188630
rect 175372 188566 175424 188572
rect 175372 188488 175424 188494
rect 175372 188430 175424 188436
rect 175384 148889 175412 188430
rect 175476 151337 175504 191134
rect 175556 191004 175608 191010
rect 175556 190946 175608 190952
rect 175568 151366 175596 190946
rect 176028 189990 176056 199736
rect 176120 199736 176194 199764
rect 176292 199776 176344 199782
rect 176120 191010 176148 199736
rect 176534 199764 176562 200124
rect 176292 199718 176344 199724
rect 176488 199736 176562 199764
rect 176200 195900 176252 195906
rect 176200 195842 176252 195848
rect 176108 191004 176160 191010
rect 176108 190946 176160 190952
rect 176016 189984 176068 189990
rect 176016 189926 176068 189932
rect 175648 188624 175700 188630
rect 175648 188566 175700 188572
rect 175556 151360 175608 151366
rect 175462 151328 175518 151337
rect 175556 151302 175608 151308
rect 175660 151298 175688 188566
rect 175740 159792 175792 159798
rect 175740 159734 175792 159740
rect 175462 151263 175518 151272
rect 175648 151292 175700 151298
rect 175648 151234 175700 151240
rect 175370 148880 175426 148889
rect 175370 148815 175426 148824
rect 175278 145888 175334 145897
rect 175278 145823 175334 145832
rect 175648 143268 175700 143274
rect 175648 143210 175700 143216
rect 175188 141976 175240 141982
rect 175188 141918 175240 141924
rect 175200 139890 175228 141918
rect 175660 139890 175688 143210
rect 174004 139862 174340 139890
rect 174892 139862 175228 139890
rect 175444 139862 175688 139890
rect 175752 139890 175780 159734
rect 176212 141846 176240 195842
rect 176304 195770 176332 199718
rect 176382 198928 176438 198937
rect 176382 198863 176438 198872
rect 176292 195764 176344 195770
rect 176292 195706 176344 195712
rect 176396 188494 176424 198863
rect 176488 190058 176516 199736
rect 176626 199628 176654 200124
rect 176718 199764 176746 200124
rect 176810 199918 176838 200124
rect 176798 199912 176850 199918
rect 176798 199854 176850 199860
rect 176718 199736 176792 199764
rect 176580 199600 176654 199628
rect 176580 195945 176608 199600
rect 176660 199504 176712 199510
rect 176660 199446 176712 199452
rect 176566 195936 176622 195945
rect 176566 195871 176622 195880
rect 176672 194041 176700 199446
rect 176658 194032 176714 194041
rect 176658 193967 176714 193976
rect 176660 193180 176712 193186
rect 176660 193122 176712 193128
rect 176476 190052 176528 190058
rect 176476 189994 176528 190000
rect 176384 188488 176436 188494
rect 176384 188430 176436 188436
rect 176672 151201 176700 193122
rect 176658 151192 176714 151201
rect 176764 151162 176792 199736
rect 176902 199696 176930 200124
rect 176994 199764 177022 200124
rect 177086 199918 177114 200124
rect 177178 199918 177206 200124
rect 177270 199918 177298 200124
rect 177362 199918 177390 200124
rect 177074 199912 177126 199918
rect 177074 199854 177126 199860
rect 177166 199912 177218 199918
rect 177166 199854 177218 199860
rect 177258 199912 177310 199918
rect 177258 199854 177310 199860
rect 177350 199912 177402 199918
rect 177454 199900 177482 200124
rect 177546 199968 177574 200124
rect 177652 200110 177804 200138
rect 177546 199940 177620 199968
rect 177454 199889 177528 199900
rect 177454 199880 177542 199889
rect 177454 199872 177486 199880
rect 177350 199854 177402 199860
rect 177486 199815 177542 199824
rect 176994 199736 177068 199764
rect 176902 199668 176976 199696
rect 176844 199572 176896 199578
rect 176844 199514 176896 199520
rect 176856 193066 176884 199514
rect 176948 196042 176976 199668
rect 176936 196036 176988 196042
rect 176936 195978 176988 195984
rect 177040 193186 177068 199736
rect 177120 199640 177172 199646
rect 177120 199582 177172 199588
rect 177212 199640 177264 199646
rect 177212 199582 177264 199588
rect 177396 199640 177448 199646
rect 177396 199582 177448 199588
rect 177132 197946 177160 199582
rect 177224 198801 177252 199582
rect 177304 199504 177356 199510
rect 177304 199446 177356 199452
rect 177210 198792 177266 198801
rect 177210 198727 177266 198736
rect 177120 197940 177172 197946
rect 177120 197882 177172 197888
rect 177316 197354 177344 199446
rect 177408 199345 177436 199582
rect 177394 199336 177450 199345
rect 177394 199271 177450 199280
rect 177394 198792 177450 198801
rect 177394 198727 177450 198736
rect 177224 197326 177344 197354
rect 177028 193180 177080 193186
rect 177028 193122 177080 193128
rect 176856 193038 177160 193066
rect 176936 190936 176988 190942
rect 176936 190878 176988 190884
rect 176844 190868 176896 190874
rect 176844 190810 176896 190816
rect 176856 153785 176884 190810
rect 176948 157146 176976 190878
rect 177132 190126 177160 193038
rect 177120 190120 177172 190126
rect 177120 190062 177172 190068
rect 177224 189922 177252 197326
rect 177408 190874 177436 198727
rect 177396 190868 177448 190874
rect 177396 190810 177448 190816
rect 177212 189916 177264 189922
rect 177212 189858 177264 189864
rect 177592 186314 177620 199940
rect 177776 199730 177804 200110
rect 177868 200002 177896 200194
rect 177960 200161 177988 200466
rect 178052 200190 178080 200534
rect 178040 200184 178092 200190
rect 177946 200152 178002 200161
rect 178040 200126 178092 200132
rect 177946 200087 178002 200096
rect 177868 199974 177988 200002
rect 177856 199912 177908 199918
rect 177856 199854 177908 199860
rect 177684 199702 177804 199730
rect 177684 190942 177712 199702
rect 177764 197940 177816 197946
rect 177764 197882 177816 197888
rect 177776 195129 177804 197882
rect 177762 195120 177818 195129
rect 177762 195055 177818 195064
rect 177868 194206 177896 199854
rect 177960 198665 177988 199974
rect 177946 198656 178002 198665
rect 177946 198591 178002 198600
rect 178144 197810 178172 200534
rect 178236 198665 178264 200631
rect 180064 200602 180116 200608
rect 178408 200388 178460 200394
rect 178408 200330 178460 200336
rect 178420 199102 178448 200330
rect 178592 199572 178644 199578
rect 178592 199514 178644 199520
rect 178604 199209 178632 199514
rect 178684 199436 178736 199442
rect 178684 199378 178736 199384
rect 178590 199200 178646 199209
rect 178590 199135 178646 199144
rect 178408 199096 178460 199102
rect 178408 199038 178460 199044
rect 178222 198656 178278 198665
rect 178222 198591 178278 198600
rect 178132 197804 178184 197810
rect 178132 197746 178184 197752
rect 177856 194200 177908 194206
rect 177856 194142 177908 194148
rect 177948 192296 178000 192302
rect 177948 192238 178000 192244
rect 177672 190936 177724 190942
rect 177672 190878 177724 190884
rect 177040 186286 177620 186314
rect 176936 157140 176988 157146
rect 176936 157082 176988 157088
rect 177040 153921 177068 186286
rect 177856 157344 177908 157350
rect 177856 157286 177908 157292
rect 177026 153912 177082 153921
rect 177026 153847 177082 153856
rect 176842 153776 176898 153785
rect 176842 153711 176898 153720
rect 176658 151127 176714 151136
rect 176752 151156 176804 151162
rect 176752 151098 176804 151104
rect 177212 146124 177264 146130
rect 177212 146066 177264 146072
rect 177120 143540 177172 143546
rect 177120 143482 177172 143488
rect 176476 142044 176528 142050
rect 176476 141986 176528 141992
rect 176200 141840 176252 141846
rect 176200 141782 176252 141788
rect 176488 139890 176516 141986
rect 177132 140162 177160 143482
rect 177086 140134 177160 140162
rect 175752 139862 175996 139890
rect 176488 139862 176548 139890
rect 177086 139876 177114 140134
rect 177224 139890 177252 146066
rect 177868 142390 177896 157286
rect 177960 142594 177988 192238
rect 178224 146260 178276 146266
rect 178224 146202 178276 146208
rect 178040 146192 178092 146198
rect 178040 146134 178092 146140
rect 177948 142588 178000 142594
rect 177948 142530 178000 142536
rect 177856 142384 177908 142390
rect 177856 142326 177908 142332
rect 177868 141409 177896 142326
rect 177854 141400 177910 141409
rect 177854 141335 177910 141344
rect 177960 140049 177988 142530
rect 178052 140690 178080 146134
rect 178040 140684 178092 140690
rect 178040 140626 178092 140632
rect 178236 140162 178264 146202
rect 178316 145512 178368 145518
rect 178316 145454 178368 145460
rect 178190 140134 178264 140162
rect 177946 140040 178002 140049
rect 177946 139975 178002 139984
rect 177224 139862 177652 139890
rect 178190 139876 178218 140134
rect 178328 139890 178356 145454
rect 178696 140350 178724 199378
rect 178868 198892 178920 198898
rect 178868 198834 178920 198840
rect 178776 198824 178828 198830
rect 178776 198766 178828 198772
rect 178788 140486 178816 198766
rect 178880 142934 178908 198834
rect 179420 197668 179472 197674
rect 179420 197610 179472 197616
rect 178960 197464 179012 197470
rect 178960 197406 179012 197412
rect 178868 142928 178920 142934
rect 178868 142870 178920 142876
rect 178972 142769 179000 197406
rect 179052 196580 179104 196586
rect 179052 196522 179104 196528
rect 179064 147626 179092 196522
rect 179144 194880 179196 194886
rect 179144 194822 179196 194828
rect 179052 147620 179104 147626
rect 179052 147562 179104 147568
rect 179156 146878 179184 194822
rect 179432 192409 179460 197610
rect 179418 192400 179474 192409
rect 179418 192335 179474 192344
rect 179144 146872 179196 146878
rect 179144 146814 179196 146820
rect 179420 145580 179472 145586
rect 179420 145522 179472 145528
rect 179432 143546 179460 145522
rect 179512 145444 179564 145450
rect 179512 145386 179564 145392
rect 179420 143540 179472 143546
rect 179420 143482 179472 143488
rect 178958 142760 179014 142769
rect 178958 142695 179014 142704
rect 179524 142154 179552 145386
rect 179432 142126 179552 142154
rect 178960 140684 179012 140690
rect 178960 140626 179012 140632
rect 178776 140480 178828 140486
rect 178776 140422 178828 140428
rect 178684 140344 178736 140350
rect 178684 140286 178736 140292
rect 178972 139890 179000 140626
rect 179432 139890 179460 142126
rect 180076 140418 180104 200602
rect 180340 200456 180392 200462
rect 180340 200398 180392 200404
rect 181442 200424 181498 200433
rect 180156 198960 180208 198966
rect 180156 198902 180208 198908
rect 180064 140412 180116 140418
rect 180064 140354 180116 140360
rect 180168 140049 180196 198902
rect 180246 195800 180302 195809
rect 180246 195735 180302 195744
rect 180260 140282 180288 195735
rect 180352 146169 180380 200398
rect 181442 200359 181498 200368
rect 181076 198756 181128 198762
rect 181076 198698 181128 198704
rect 180524 196376 180576 196382
rect 180524 196318 180576 196324
rect 180338 146160 180394 146169
rect 180338 146095 180394 146104
rect 180536 146033 180564 196318
rect 181088 157334 181116 198698
rect 181352 195832 181404 195838
rect 181352 195774 181404 195780
rect 181364 195498 181392 195774
rect 181352 195492 181404 195498
rect 181352 195434 181404 195440
rect 181352 193928 181404 193934
rect 181352 193870 181404 193876
rect 181364 193594 181392 193870
rect 181352 193588 181404 193594
rect 181352 193530 181404 193536
rect 181088 157306 181208 157334
rect 180892 149592 180944 149598
rect 180892 149534 180944 149540
rect 180904 149190 180932 149534
rect 180892 149184 180944 149190
rect 180892 149126 180944 149132
rect 180522 146024 180578 146033
rect 180522 145959 180578 145968
rect 180340 141908 180392 141914
rect 180340 141850 180392 141856
rect 180248 140276 180300 140282
rect 180248 140218 180300 140224
rect 180154 140040 180210 140049
rect 180154 139975 180210 139984
rect 178328 139862 178756 139890
rect 178972 139862 179308 139890
rect 179432 139862 179860 139890
rect 180064 139664 180116 139670
rect 180352 139618 180380 141850
rect 180904 139890 180932 149126
rect 181180 139890 181208 157306
rect 181456 147665 181484 200359
rect 182824 199436 182876 199442
rect 182824 199378 182876 199384
rect 181536 193724 181588 193730
rect 181536 193666 181588 193672
rect 181442 147656 181498 147665
rect 181442 147591 181498 147600
rect 181548 144838 181576 193666
rect 181628 193656 181680 193662
rect 181628 193598 181680 193604
rect 181640 146606 181668 193598
rect 181720 190256 181772 190262
rect 181720 190198 181772 190204
rect 181732 146810 181760 190198
rect 181812 151632 181864 151638
rect 181812 151574 181864 151580
rect 181720 146804 181772 146810
rect 181720 146746 181772 146752
rect 181628 146600 181680 146606
rect 181628 146542 181680 146548
rect 181536 144832 181588 144838
rect 181536 144774 181588 144780
rect 180904 139862 180964 139890
rect 181180 139862 181516 139890
rect 180116 139612 180412 139618
rect 180064 139606 180412 139612
rect 180076 139590 180412 139606
rect 181180 139534 181208 139862
rect 181824 139777 181852 151574
rect 182088 149660 182140 149666
rect 182088 149602 182140 149608
rect 181904 147484 181956 147490
rect 181904 147426 181956 147432
rect 181916 141409 181944 147426
rect 182100 144158 182128 149602
rect 182088 144152 182140 144158
rect 182088 144094 182140 144100
rect 182732 143336 182784 143342
rect 182732 143278 182784 143284
rect 182744 142458 182772 143278
rect 182732 142452 182784 142458
rect 182732 142394 182784 142400
rect 181996 142384 182048 142390
rect 181996 142326 182048 142332
rect 181902 141400 181958 141409
rect 181902 141335 181958 141344
rect 182008 139890 182036 142326
rect 182744 139890 182772 142394
rect 182836 140894 182864 199378
rect 182916 195152 182968 195158
rect 182916 195094 182968 195100
rect 182928 142154 182956 195094
rect 183192 193860 183244 193866
rect 183192 193802 183244 193808
rect 183100 190392 183152 190398
rect 183100 190334 183152 190340
rect 183008 190188 183060 190194
rect 183008 190130 183060 190136
rect 183020 143546 183048 190130
rect 183008 143540 183060 143546
rect 183008 143482 183060 143488
rect 183112 143449 183140 190334
rect 183204 146742 183232 193802
rect 183744 154352 183796 154358
rect 183744 154294 183796 154300
rect 183284 153808 183336 153814
rect 183284 153750 183336 153756
rect 183192 146736 183244 146742
rect 183192 146678 183244 146684
rect 183296 144294 183324 153750
rect 183650 151056 183706 151065
rect 183650 150991 183706 151000
rect 183284 144288 183336 144294
rect 183284 144230 183336 144236
rect 183098 143440 183154 143449
rect 183098 143375 183154 143384
rect 183664 142186 183692 150991
rect 183756 145382 183784 154294
rect 184216 147674 184244 200670
rect 186688 199912 186740 199918
rect 186688 199854 186740 199860
rect 185584 198824 185636 198830
rect 185584 198766 185636 198772
rect 184296 154420 184348 154426
rect 184296 154362 184348 154368
rect 184032 147646 184244 147674
rect 183744 145376 183796 145382
rect 183744 145318 183796 145324
rect 184032 144906 184060 147646
rect 184308 146962 184336 154362
rect 185492 152448 185544 152454
rect 185492 152390 185544 152396
rect 185400 151564 185452 151570
rect 185400 151506 185452 151512
rect 184388 151496 184440 151502
rect 184388 151438 184440 151444
rect 184124 146934 184336 146962
rect 184020 144900 184072 144906
rect 184020 144842 184072 144848
rect 183742 143168 183798 143177
rect 183742 143103 183798 143112
rect 183756 142361 183784 143103
rect 183742 142352 183798 142361
rect 183742 142287 183798 142296
rect 183652 142180 183704 142186
rect 182928 142126 183048 142154
rect 182916 141840 182968 141846
rect 182916 141782 182968 141788
rect 182928 141370 182956 141782
rect 182916 141364 182968 141370
rect 182916 141306 182968 141312
rect 182824 140888 182876 140894
rect 182824 140830 182876 140836
rect 182008 139862 182068 139890
rect 182620 139862 182772 139890
rect 182836 139890 182864 140830
rect 183020 140729 183048 142126
rect 183652 142122 183704 142128
rect 183006 140720 183062 140729
rect 183006 140655 183062 140664
rect 183374 140176 183430 140185
rect 183756 140162 183784 142287
rect 184124 141166 184152 146934
rect 184294 143304 184350 143313
rect 184294 143239 184350 143248
rect 184204 143064 184256 143070
rect 184204 143006 184256 143012
rect 184112 141160 184164 141166
rect 184112 141102 184164 141108
rect 184216 140894 184244 143006
rect 184308 142225 184336 143239
rect 184294 142216 184350 142225
rect 184294 142151 184350 142160
rect 184204 140888 184256 140894
rect 184204 140830 184256 140836
rect 184308 140162 184336 142151
rect 183374 140111 183430 140120
rect 183710 140134 183784 140162
rect 184262 140134 184336 140162
rect 183388 139913 183416 140111
rect 183374 139904 183430 139913
rect 182836 139862 183172 139890
rect 183710 139876 183738 140134
rect 184262 139876 184290 140134
rect 183374 139839 183430 139848
rect 181810 139768 181866 139777
rect 181810 139703 181866 139712
rect 181168 139528 181220 139534
rect 184400 139505 184428 151438
rect 184848 151428 184900 151434
rect 184848 151370 184900 151376
rect 184572 148844 184624 148850
rect 184572 148786 184624 148792
rect 184480 142588 184532 142594
rect 184480 142530 184532 142536
rect 184492 139890 184520 142530
rect 184584 140010 184612 148786
rect 184860 140554 184888 151370
rect 184848 140548 184900 140554
rect 184848 140490 184900 140496
rect 185412 140185 185440 151506
rect 185504 143410 185532 152390
rect 185492 143404 185544 143410
rect 185492 143346 185544 143352
rect 185596 141846 185624 198766
rect 186596 195696 186648 195702
rect 186596 195638 186648 195644
rect 185768 190460 185820 190466
rect 185768 190402 185820 190408
rect 185676 190324 185728 190330
rect 185676 190266 185728 190272
rect 185688 152454 185716 190266
rect 185676 152448 185728 152454
rect 185676 152390 185728 152396
rect 185780 147674 185808 190402
rect 185860 154556 185912 154562
rect 185860 154498 185912 154504
rect 185688 147646 185808 147674
rect 185688 144974 185716 147646
rect 185768 146872 185820 146878
rect 185768 146814 185820 146820
rect 185676 144968 185728 144974
rect 185676 144910 185728 144916
rect 185676 143064 185728 143070
rect 185676 143006 185728 143012
rect 185584 141840 185636 141846
rect 185584 141782 185636 141788
rect 185688 141250 185716 143006
rect 185504 141222 185716 141250
rect 185398 140176 185454 140185
rect 185398 140111 185454 140120
rect 184572 140004 184624 140010
rect 184572 139946 184624 139952
rect 184492 139862 184828 139890
rect 185504 139618 185532 141222
rect 185582 140584 185638 140593
rect 185582 140519 185638 140528
rect 185596 140185 185624 140519
rect 185582 140176 185638 140185
rect 185582 140111 185638 140120
rect 185044 139602 185532 139618
rect 185032 139596 185532 139602
rect 185084 139590 185532 139596
rect 185582 139632 185638 139641
rect 185780 139618 185808 146814
rect 185872 140214 185900 154498
rect 185952 154488 186004 154494
rect 185952 154430 186004 154436
rect 185964 142118 185992 154430
rect 186136 154284 186188 154290
rect 186136 154226 186188 154232
rect 186044 154216 186096 154222
rect 186044 154158 186096 154164
rect 186056 146878 186084 154158
rect 186044 146872 186096 146878
rect 186044 146814 186096 146820
rect 186044 143472 186096 143478
rect 186044 143414 186096 143420
rect 186056 142322 186084 143414
rect 186044 142316 186096 142322
rect 186044 142258 186096 142264
rect 185952 142112 186004 142118
rect 185952 142054 186004 142060
rect 185952 141840 186004 141846
rect 185952 141782 186004 141788
rect 185860 140208 185912 140214
rect 185860 140150 185912 140156
rect 185964 140146 185992 141782
rect 185952 140140 186004 140146
rect 185952 140082 186004 140088
rect 186056 139890 186084 142258
rect 185932 139862 186084 139890
rect 185638 139590 185808 139618
rect 185582 139567 185638 139576
rect 185032 139538 185084 139544
rect 181168 139470 181220 139476
rect 184386 139496 184442 139505
rect 184386 139431 184442 139440
rect 123668 139334 123720 139340
rect 123942 139360 123998 139369
rect 123022 139295 123078 139304
rect 123942 139295 123998 139304
rect 125506 139360 125562 139369
rect 125506 139295 125562 139304
rect 130566 139360 130622 139369
rect 130566 139295 130622 139304
rect 130842 139360 130898 139369
rect 130842 139295 130898 139304
rect 162306 139360 162362 139369
rect 162306 139295 162362 139304
rect 169482 139360 169538 139369
rect 169482 139295 169538 139304
rect 173622 139360 173678 139369
rect 186148 139346 186176 154226
rect 186228 154148 186280 154154
rect 186228 154090 186280 154096
rect 186240 139505 186268 154090
rect 186226 139496 186282 139505
rect 186226 139431 186282 139440
rect 186226 139360 186282 139369
rect 186148 139318 186226 139346
rect 173622 139295 173678 139304
rect 186226 139295 186282 139304
rect 131028 80640 131080 80646
rect 122746 80608 122802 80617
rect 132224 80640 132276 80646
rect 131946 80608 132002 80617
rect 131080 80588 131160 80594
rect 131028 80582 131160 80588
rect 131040 80566 131160 80582
rect 122746 80543 122802 80552
rect 122760 79354 122788 80543
rect 123942 80472 123998 80481
rect 123942 80407 123998 80416
rect 123484 79960 123536 79966
rect 123484 79902 123536 79908
rect 122656 79348 122708 79354
rect 122656 79290 122708 79296
rect 122748 79348 122800 79354
rect 122748 79290 122800 79296
rect 122668 78441 122696 79290
rect 122654 78432 122710 78441
rect 122654 78367 122710 78376
rect 123496 78305 123524 79902
rect 123482 78296 123538 78305
rect 123482 78231 123538 78240
rect 123956 75886 123984 80407
rect 131132 80238 131160 80566
rect 132224 80582 132276 80588
rect 178684 80640 178736 80646
rect 178684 80582 178736 80588
rect 178776 80640 178828 80646
rect 178776 80582 178828 80588
rect 180522 80608 180578 80617
rect 131946 80543 132002 80552
rect 131120 80232 131172 80238
rect 131120 80174 131172 80180
rect 131670 80200 131726 80209
rect 131670 80135 131726 80144
rect 128634 80064 128690 80073
rect 128634 79999 128690 80008
rect 129096 80028 129148 80034
rect 126058 79928 126114 79937
rect 126058 79863 126114 79872
rect 128176 79892 128228 79898
rect 124862 78160 124918 78169
rect 124862 78095 124918 78104
rect 124876 77450 124904 78095
rect 125600 77784 125652 77790
rect 125600 77726 125652 77732
rect 124864 77444 124916 77450
rect 124864 77386 124916 77392
rect 123944 75880 123996 75886
rect 123944 75822 123996 75828
rect 122472 73092 122524 73098
rect 122472 73034 122524 73040
rect 122288 3800 122340 3806
rect 122288 3742 122340 3748
rect 122104 3188 122156 3194
rect 122104 3130 122156 3136
rect 122300 480 122328 3742
rect 124876 3534 124904 77386
rect 125612 75002 125640 77726
rect 126072 77489 126100 79863
rect 128176 79834 128228 79840
rect 126336 79620 126388 79626
rect 126336 79562 126388 79568
rect 126242 79384 126298 79393
rect 126242 79319 126298 79328
rect 126256 79150 126284 79319
rect 126348 79150 126376 79562
rect 127900 79552 127952 79558
rect 127900 79494 127952 79500
rect 127808 79484 127860 79490
rect 127808 79426 127860 79432
rect 126244 79144 126296 79150
rect 126244 79086 126296 79092
rect 126336 79144 126388 79150
rect 126336 79086 126388 79092
rect 127820 78742 127848 79426
rect 127912 78810 127940 79494
rect 127900 78804 127952 78810
rect 127900 78746 127952 78752
rect 127808 78736 127860 78742
rect 127808 78678 127860 78684
rect 126058 77480 126114 77489
rect 126058 77415 126114 77424
rect 126244 76628 126296 76634
rect 126244 76570 126296 76576
rect 126256 76226 126284 76570
rect 126980 76492 127032 76498
rect 126980 76434 127032 76440
rect 126244 76220 126296 76226
rect 126244 76162 126296 76168
rect 126992 76158 127020 76434
rect 126980 76152 127032 76158
rect 126980 76094 127032 76100
rect 125600 74996 125652 75002
rect 125600 74938 125652 74944
rect 125612 3670 125640 74938
rect 126992 16574 127020 76094
rect 128188 71233 128216 79834
rect 128648 72282 128676 79999
rect 129096 79970 129148 79976
rect 129002 78432 129058 78441
rect 129002 78367 129058 78376
rect 128636 72276 128688 72282
rect 128636 72218 128688 72224
rect 128452 71732 128504 71738
rect 128452 71674 128504 71680
rect 128174 71224 128230 71233
rect 128174 71159 128230 71168
rect 128360 71120 128412 71126
rect 128360 71062 128412 71068
rect 126992 16546 127112 16574
rect 127084 3806 127112 16546
rect 127072 3800 127124 3806
rect 127072 3742 127124 3748
rect 125600 3664 125652 3670
rect 125600 3606 125652 3612
rect 125876 3596 125928 3602
rect 125876 3538 125928 3544
rect 123484 3528 123536 3534
rect 123484 3470 123536 3476
rect 124864 3528 124916 3534
rect 124864 3470 124916 3476
rect 123496 480 123524 3470
rect 124680 3460 124732 3466
rect 124680 3402 124732 3408
rect 124692 480 124720 3402
rect 125888 480 125916 3538
rect 126980 3528 127032 3534
rect 126980 3470 127032 3476
rect 126992 480 127020 3470
rect 128176 2916 128228 2922
rect 128176 2858 128228 2864
rect 128188 480 128216 2858
rect 128372 490 128400 71062
rect 128464 3534 128492 71674
rect 128452 3528 128504 3534
rect 128452 3470 128504 3476
rect 129016 2922 129044 78367
rect 129108 74390 129136 79970
rect 131396 79824 131448 79830
rect 131396 79766 131448 79772
rect 130936 78804 130988 78810
rect 130936 78746 130988 78752
rect 129832 78056 129884 78062
rect 129832 77998 129884 78004
rect 129648 76424 129700 76430
rect 129648 76366 129700 76372
rect 129096 74384 129148 74390
rect 129096 74326 129148 74332
rect 129660 71738 129688 76366
rect 129738 75304 129794 75313
rect 129738 75239 129794 75248
rect 129648 71732 129700 71738
rect 129648 71674 129700 71680
rect 129752 3482 129780 75239
rect 129844 3670 129872 77998
rect 130842 77616 130898 77625
rect 130842 77551 130898 77560
rect 129924 72344 129976 72350
rect 129924 72286 129976 72292
rect 129832 3664 129884 3670
rect 129832 3606 129884 3612
rect 129936 3602 129964 72286
rect 130856 3806 130884 77551
rect 130844 3800 130896 3806
rect 130844 3742 130896 3748
rect 130948 3602 130976 78746
rect 131028 78736 131080 78742
rect 131028 78678 131080 78684
rect 131040 3670 131068 78678
rect 131304 77716 131356 77722
rect 131304 77658 131356 77664
rect 131120 75336 131172 75342
rect 131172 75284 131252 75290
rect 131120 75278 131252 75284
rect 131132 75262 131252 75278
rect 131120 74588 131172 74594
rect 131120 74530 131172 74536
rect 131132 73846 131160 74530
rect 131224 73846 131252 75262
rect 131120 73840 131172 73846
rect 131120 73782 131172 73788
rect 131212 73840 131264 73846
rect 131212 73782 131264 73788
rect 131316 73658 131344 77658
rect 131408 75206 131436 79766
rect 131684 78441 131712 80135
rect 131960 79558 131988 80543
rect 132236 80306 132264 80582
rect 132224 80300 132276 80306
rect 132224 80242 132276 80248
rect 177764 80164 177816 80170
rect 177764 80106 177816 80112
rect 132052 80022 132388 80050
rect 131948 79552 132000 79558
rect 131948 79494 132000 79500
rect 132052 78577 132080 80022
rect 132466 79778 132494 80036
rect 132558 79937 132586 80036
rect 132544 79928 132600 79937
rect 132544 79863 132600 79872
rect 132650 79778 132678 80036
rect 132742 79801 132770 80036
rect 132420 79750 132494 79778
rect 132604 79750 132678 79778
rect 132728 79792 132784 79801
rect 132038 78568 132094 78577
rect 132038 78503 132094 78512
rect 131670 78432 131726 78441
rect 131670 78367 131726 78376
rect 132314 78432 132370 78441
rect 132314 78367 132370 78376
rect 132328 77926 132356 78367
rect 132316 77920 132368 77926
rect 132316 77862 132368 77868
rect 131672 77512 131724 77518
rect 131672 77454 131724 77460
rect 131578 76664 131634 76673
rect 131578 76599 131634 76608
rect 131488 75268 131540 75274
rect 131488 75210 131540 75216
rect 131396 75200 131448 75206
rect 131396 75142 131448 75148
rect 131132 73630 131344 73658
rect 131132 16574 131160 73630
rect 131304 73568 131356 73574
rect 131304 73510 131356 73516
rect 131132 16546 131252 16574
rect 131028 3664 131080 3670
rect 131028 3606 131080 3612
rect 129924 3596 129976 3602
rect 129924 3538 129976 3544
rect 130936 3596 130988 3602
rect 130936 3538 130988 3544
rect 129752 3454 130608 3482
rect 129004 2916 129056 2922
rect 129004 2858 129056 2864
rect 121062 354 121174 480
rect 120644 326 121174 354
rect 121062 -960 121174 326
rect 122258 -960 122370 480
rect 123454 -960 123566 480
rect 124650 -960 124762 480
rect 125846 -960 125958 480
rect 126950 -960 127062 480
rect 128146 -960 128258 480
rect 128372 462 128952 490
rect 130580 480 130608 3454
rect 128924 354 128952 462
rect 129342 354 129454 480
rect 128924 326 129454 354
rect 129342 -960 129454 326
rect 130538 -960 130650 480
rect 131224 354 131252 16546
rect 131316 3466 131344 73510
rect 131304 3460 131356 3466
rect 131304 3402 131356 3408
rect 131408 3398 131436 75142
rect 131500 3738 131528 75210
rect 131592 75206 131620 76599
rect 131580 75200 131632 75206
rect 131580 75142 131632 75148
rect 131488 3732 131540 3738
rect 131488 3674 131540 3680
rect 131396 3392 131448 3398
rect 131396 3334 131448 3340
rect 131592 3330 131620 75142
rect 131684 73574 131712 77454
rect 132420 73642 132448 79750
rect 132500 79688 132552 79694
rect 132500 79630 132552 79636
rect 132512 78538 132540 79630
rect 132500 78532 132552 78538
rect 132500 78474 132552 78480
rect 132604 76673 132632 79750
rect 132834 79778 132862 80036
rect 132926 79966 132954 80036
rect 132914 79960 132966 79966
rect 132914 79902 132966 79908
rect 132834 79750 132908 79778
rect 132728 79727 132784 79736
rect 132590 76664 132646 76673
rect 132590 76599 132646 76608
rect 132408 73636 132460 73642
rect 132408 73578 132460 73584
rect 131672 73568 131724 73574
rect 131672 73510 131724 73516
rect 132880 73154 132908 79750
rect 133018 79676 133046 80036
rect 133110 79937 133138 80036
rect 133096 79928 133152 79937
rect 133096 79863 133152 79872
rect 133202 79778 133230 80036
rect 133294 79898 133322 80036
rect 133282 79892 133334 79898
rect 133282 79834 133334 79840
rect 133386 79778 133414 80036
rect 133478 79971 133506 80036
rect 133464 79962 133520 79971
rect 133570 79966 133598 80036
rect 133662 79966 133690 80036
rect 133754 79966 133782 80036
rect 133464 79897 133520 79906
rect 133558 79960 133610 79966
rect 133558 79902 133610 79908
rect 133650 79960 133702 79966
rect 133650 79902 133702 79908
rect 133742 79960 133794 79966
rect 133742 79902 133794 79908
rect 133846 79812 133874 80036
rect 133938 79966 133966 80036
rect 133926 79960 133978 79966
rect 133926 79902 133978 79908
rect 134030 79898 134058 80036
rect 134018 79892 134070 79898
rect 134018 79834 134070 79840
rect 133156 79750 133230 79778
rect 133340 79750 133414 79778
rect 133510 79792 133566 79801
rect 133018 79648 133092 79676
rect 132880 73126 133000 73154
rect 132972 72962 133000 73126
rect 132960 72956 133012 72962
rect 132960 72898 133012 72904
rect 132972 72162 133000 72898
rect 132604 72134 133000 72162
rect 132040 68944 132092 68950
rect 132040 68886 132092 68892
rect 132052 68814 132080 68886
rect 132236 68882 132448 68898
rect 132224 68876 132460 68882
rect 132276 68870 132408 68876
rect 132224 68818 132276 68824
rect 132408 68818 132460 68824
rect 131948 68808 132000 68814
rect 131948 68750 132000 68756
rect 132040 68808 132092 68814
rect 132040 68750 132092 68756
rect 131960 68474 131988 68750
rect 131948 68468 132000 68474
rect 131948 68410 132000 68416
rect 132604 8974 132632 72134
rect 132868 72072 132920 72078
rect 132868 72014 132920 72020
rect 132880 37942 132908 72014
rect 133064 65890 133092 79648
rect 133156 75206 133184 79750
rect 133236 79688 133288 79694
rect 133236 79630 133288 79636
rect 133144 75200 133196 75206
rect 133144 75142 133196 75148
rect 133052 65884 133104 65890
rect 133052 65826 133104 65832
rect 133248 60734 133276 79630
rect 133340 74633 133368 79750
rect 133800 79784 133874 79812
rect 133510 79727 133566 79736
rect 133604 79756 133656 79762
rect 133524 77217 133552 79727
rect 133604 79698 133656 79704
rect 133510 77208 133566 77217
rect 133510 77143 133566 77152
rect 133326 74624 133382 74633
rect 133326 74559 133382 74568
rect 133524 72078 133552 77143
rect 133512 72072 133564 72078
rect 133512 72014 133564 72020
rect 133616 68542 133644 79698
rect 133694 79656 133750 79665
rect 133694 79591 133750 79600
rect 133708 78334 133736 79591
rect 133696 78328 133748 78334
rect 133696 78270 133748 78276
rect 133800 73030 133828 79784
rect 134122 79778 134150 80036
rect 134214 79812 134242 80036
rect 134306 79966 134334 80036
rect 134398 79966 134426 80036
rect 134294 79960 134346 79966
rect 134294 79902 134346 79908
rect 134386 79960 134438 79966
rect 134490 79937 134518 80036
rect 134582 79966 134610 80036
rect 134570 79960 134622 79966
rect 134386 79902 134438 79908
rect 134476 79928 134532 79937
rect 134570 79902 134622 79908
rect 134674 79898 134702 80036
rect 134766 79971 134794 80036
rect 134752 79962 134808 79971
rect 134476 79863 134532 79872
rect 134662 79892 134714 79898
rect 134752 79897 134808 79906
rect 134662 79834 134714 79840
rect 134524 79824 134576 79830
rect 134214 79784 134288 79812
rect 134076 79750 134150 79778
rect 133880 79688 133932 79694
rect 133880 79630 133932 79636
rect 133892 77353 133920 79630
rect 133972 79620 134024 79626
rect 133972 79562 134024 79568
rect 133878 77344 133934 77353
rect 133878 77279 133934 77288
rect 133880 76696 133932 76702
rect 133880 76638 133932 76644
rect 133788 73024 133840 73030
rect 133788 72966 133840 72972
rect 133604 68536 133656 68542
rect 133604 68478 133656 68484
rect 133156 60706 133276 60734
rect 133156 52426 133184 60706
rect 133144 52420 133196 52426
rect 133144 52362 133196 52368
rect 132868 37936 132920 37942
rect 132868 37878 132920 37884
rect 132592 8968 132644 8974
rect 132592 8910 132644 8916
rect 133892 4826 133920 76638
rect 133984 75585 134012 79562
rect 134076 76673 134104 79750
rect 134156 79688 134208 79694
rect 134156 79630 134208 79636
rect 134168 78849 134196 79630
rect 134154 78840 134210 78849
rect 134154 78775 134210 78784
rect 134168 76702 134196 78775
rect 134156 76696 134208 76702
rect 134062 76664 134118 76673
rect 134156 76638 134208 76644
rect 134062 76599 134118 76608
rect 134260 76514 134288 79784
rect 134524 79766 134576 79772
rect 134858 79778 134886 80036
rect 134950 79898 134978 80036
rect 134938 79892 134990 79898
rect 134938 79834 134990 79840
rect 134432 79756 134484 79762
rect 134432 79698 134484 79704
rect 134340 79484 134392 79490
rect 134340 79426 134392 79432
rect 134352 78062 134380 79426
rect 134340 78056 134392 78062
rect 134340 77998 134392 78004
rect 134076 76486 134288 76514
rect 134340 76492 134392 76498
rect 133970 75576 134026 75585
rect 133970 75511 134026 75520
rect 133984 10334 134012 75511
rect 134076 71369 134104 76486
rect 134340 76434 134392 76440
rect 134248 76356 134300 76362
rect 134248 76298 134300 76304
rect 134062 71360 134118 71369
rect 134062 71295 134118 71304
rect 134076 36582 134104 71295
rect 134260 66026 134288 76298
rect 134352 70378 134380 76434
rect 134340 70372 134392 70378
rect 134340 70314 134392 70320
rect 134248 66020 134300 66026
rect 134248 65962 134300 65968
rect 134352 60734 134380 70314
rect 134444 68678 134472 79698
rect 134536 78033 134564 79766
rect 134858 79750 134932 79778
rect 134800 79688 134852 79694
rect 134800 79630 134852 79636
rect 134522 78024 134578 78033
rect 134522 77959 134578 77968
rect 134522 77888 134578 77897
rect 134522 77823 134578 77832
rect 134536 77518 134564 77823
rect 134524 77512 134576 77518
rect 134524 77454 134576 77460
rect 134812 74594 134840 79630
rect 134904 76498 134932 79750
rect 135042 79676 135070 80036
rect 135134 79937 135162 80036
rect 135120 79928 135176 79937
rect 135120 79863 135176 79872
rect 135226 79778 135254 80036
rect 135318 79937 135346 80036
rect 135304 79928 135360 79937
rect 135304 79863 135360 79872
rect 135410 79778 135438 80036
rect 134996 79648 135070 79676
rect 135180 79750 135254 79778
rect 135364 79750 135438 79778
rect 135502 79778 135530 80036
rect 135594 79898 135622 80036
rect 135582 79892 135634 79898
rect 135582 79834 135634 79840
rect 135686 79830 135714 80036
rect 135778 79937 135806 80036
rect 135764 79928 135820 79937
rect 135764 79863 135820 79872
rect 135674 79824 135726 79830
rect 135502 79750 135576 79778
rect 135870 79812 135898 80036
rect 135674 79766 135726 79772
rect 135824 79784 135898 79812
rect 134996 77081 135024 79648
rect 135076 79348 135128 79354
rect 135076 79290 135128 79296
rect 135088 78266 135116 79290
rect 135076 78260 135128 78266
rect 135076 78202 135128 78208
rect 134982 77072 135038 77081
rect 134982 77007 135038 77016
rect 134892 76492 134944 76498
rect 134892 76434 134944 76440
rect 135180 76362 135208 79750
rect 135260 79688 135312 79694
rect 135260 79630 135312 79636
rect 135168 76356 135220 76362
rect 135168 76298 135220 76304
rect 135272 76242 135300 79630
rect 135364 76634 135392 79750
rect 135444 79688 135496 79694
rect 135444 79630 135496 79636
rect 135352 76628 135404 76634
rect 135352 76570 135404 76576
rect 134904 76214 135300 76242
rect 134800 74588 134852 74594
rect 134800 74530 134852 74536
rect 134904 69970 134932 76214
rect 135168 75744 135220 75750
rect 135168 75686 135220 75692
rect 135180 74746 135208 75686
rect 135260 75472 135312 75478
rect 135260 75414 135312 75420
rect 135272 74934 135300 75414
rect 135260 74928 135312 74934
rect 135260 74870 135312 74876
rect 135258 74760 135314 74769
rect 135180 74718 135258 74746
rect 135258 74695 135314 74704
rect 135272 71194 135300 74695
rect 135352 71732 135404 71738
rect 135352 71674 135404 71680
rect 135364 71534 135392 71674
rect 135352 71528 135404 71534
rect 135352 71470 135404 71476
rect 135260 71188 135312 71194
rect 135260 71130 135312 71136
rect 134892 69964 134944 69970
rect 134892 69906 134944 69912
rect 134432 68672 134484 68678
rect 134432 68614 134484 68620
rect 135456 62082 135484 79630
rect 135548 79626 135576 79750
rect 135536 79620 135588 79626
rect 135536 79562 135588 79568
rect 135628 79620 135680 79626
rect 135628 79562 135680 79568
rect 135534 79520 135590 79529
rect 135640 79506 135668 79562
rect 135640 79478 135760 79506
rect 135534 79455 135590 79464
rect 135548 78810 135576 79455
rect 135628 79416 135680 79422
rect 135628 79358 135680 79364
rect 135640 79150 135668 79358
rect 135628 79144 135680 79150
rect 135628 79086 135680 79092
rect 135536 78804 135588 78810
rect 135536 78746 135588 78752
rect 135628 78668 135680 78674
rect 135628 78610 135680 78616
rect 135536 76628 135588 76634
rect 135536 76570 135588 76576
rect 135548 66162 135576 76570
rect 135640 75313 135668 78610
rect 135732 76650 135760 79478
rect 135824 79370 135852 79784
rect 135962 79778 135990 80036
rect 136054 79898 136082 80036
rect 136042 79892 136094 79898
rect 136042 79834 136094 79840
rect 136146 79778 136174 80036
rect 136238 79801 136266 80036
rect 136330 79966 136358 80036
rect 136318 79960 136370 79966
rect 136318 79902 136370 79908
rect 135962 79750 136036 79778
rect 135824 79342 135944 79370
rect 135812 79280 135864 79286
rect 135812 79222 135864 79228
rect 135824 79150 135852 79222
rect 135812 79144 135864 79150
rect 135812 79086 135864 79092
rect 135916 77081 135944 79342
rect 135902 77072 135958 77081
rect 135902 77007 135958 77016
rect 135732 76622 135852 76650
rect 135720 76492 135772 76498
rect 135720 76434 135772 76440
rect 135626 75304 135682 75313
rect 135626 75239 135682 75248
rect 135628 73568 135680 73574
rect 135628 73510 135680 73516
rect 135640 68474 135668 73510
rect 135732 71641 135760 76434
rect 135718 71632 135774 71641
rect 135718 71567 135774 71576
rect 135720 71188 135772 71194
rect 135720 71130 135772 71136
rect 135628 68468 135680 68474
rect 135628 68410 135680 68416
rect 135536 66156 135588 66162
rect 135536 66098 135588 66104
rect 135444 62076 135496 62082
rect 135444 62018 135496 62024
rect 134168 60706 134380 60734
rect 134064 36576 134116 36582
rect 134064 36518 134116 36524
rect 134168 35222 134196 60706
rect 135352 45620 135404 45626
rect 135352 45562 135404 45568
rect 134156 35216 134208 35222
rect 134156 35158 134208 35164
rect 133972 10328 134024 10334
rect 133972 10270 134024 10276
rect 135364 6914 135392 45562
rect 135548 33794 135576 66098
rect 135536 33788 135588 33794
rect 135536 33730 135588 33736
rect 135732 26926 135760 71130
rect 135824 67318 135852 76622
rect 135904 76628 135956 76634
rect 135904 76570 135956 76576
rect 135812 67312 135864 67318
rect 135812 67254 135864 67260
rect 135916 60722 135944 76570
rect 136008 70310 136036 79750
rect 136100 79750 136174 79778
rect 136224 79792 136280 79801
rect 136100 73574 136128 79750
rect 136422 79778 136450 80036
rect 136224 79727 136280 79736
rect 136376 79750 136450 79778
rect 136514 79778 136542 80036
rect 136606 79898 136634 80036
rect 136594 79892 136646 79898
rect 136594 79834 136646 79840
rect 136698 79778 136726 80036
rect 136790 79937 136818 80036
rect 136776 79928 136832 79937
rect 136882 79898 136910 80036
rect 136776 79863 136832 79872
rect 136870 79892 136922 79898
rect 136870 79834 136922 79840
rect 136974 79778 137002 80036
rect 137066 79898 137094 80036
rect 137054 79892 137106 79898
rect 137054 79834 137106 79840
rect 137158 79801 137186 80036
rect 137144 79792 137200 79801
rect 136514 79750 136588 79778
rect 136698 79750 136864 79778
rect 136974 79750 137048 79778
rect 136272 79688 136324 79694
rect 136272 79630 136324 79636
rect 136178 79384 136234 79393
rect 136178 79319 136180 79328
rect 136232 79319 136234 79328
rect 136180 79290 136232 79296
rect 136180 79212 136232 79218
rect 136180 79154 136232 79160
rect 136192 78538 136220 79154
rect 136180 78532 136232 78538
rect 136180 78474 136232 78480
rect 136284 78198 136312 79630
rect 136272 78192 136324 78198
rect 136272 78134 136324 78140
rect 136376 76634 136404 79750
rect 136456 79620 136508 79626
rect 136456 79562 136508 79568
rect 136364 76628 136416 76634
rect 136364 76570 136416 76576
rect 136180 75404 136232 75410
rect 136180 75346 136232 75352
rect 136192 75206 136220 75346
rect 136180 75200 136232 75206
rect 136180 75142 136232 75148
rect 136088 73568 136140 73574
rect 136088 73510 136140 73516
rect 136468 73154 136496 79562
rect 136560 76498 136588 79750
rect 136640 79688 136692 79694
rect 136732 79688 136784 79694
rect 136640 79630 136692 79636
rect 136730 79656 136732 79665
rect 136784 79656 136786 79665
rect 136652 78402 136680 79630
rect 136730 79591 136786 79600
rect 136732 79484 136784 79490
rect 136732 79426 136784 79432
rect 136640 78396 136692 78402
rect 136640 78338 136692 78344
rect 136744 77110 136772 79426
rect 136732 77104 136784 77110
rect 136732 77046 136784 77052
rect 136548 76492 136600 76498
rect 136548 76434 136600 76440
rect 136732 75744 136784 75750
rect 136732 75686 136784 75692
rect 136744 73953 136772 75686
rect 136730 73944 136786 73953
rect 136730 73879 136786 73888
rect 136468 73126 136588 73154
rect 135996 70304 136048 70310
rect 135996 70246 136048 70252
rect 135904 60716 135956 60722
rect 135904 60658 135956 60664
rect 136560 31074 136588 73126
rect 136640 55276 136692 55282
rect 136640 55218 136692 55224
rect 136548 31068 136600 31074
rect 136548 31010 136600 31016
rect 135720 26920 135772 26926
rect 135720 26862 135772 26868
rect 136652 16574 136680 55218
rect 136744 42090 136772 73879
rect 136836 64802 136864 79750
rect 136916 79688 136968 79694
rect 136916 79630 136968 79636
rect 136928 78334 136956 79630
rect 136916 78328 136968 78334
rect 136916 78270 136968 78276
rect 137020 77042 137048 79750
rect 137250 79778 137278 80036
rect 137342 79966 137370 80036
rect 137330 79960 137382 79966
rect 137330 79902 137382 79908
rect 137434 79778 137462 80036
rect 137526 79898 137554 80036
rect 137514 79892 137566 79898
rect 137514 79834 137566 79840
rect 137250 79750 137324 79778
rect 137144 79727 137200 79736
rect 137100 79688 137152 79694
rect 137100 79630 137152 79636
rect 137008 77036 137060 77042
rect 137008 76978 137060 76984
rect 137008 76628 137060 76634
rect 137008 76570 137060 76576
rect 136824 64796 136876 64802
rect 136824 64738 136876 64744
rect 137020 63510 137048 76570
rect 137008 63504 137060 63510
rect 137008 63446 137060 63452
rect 137112 56574 137140 79630
rect 137296 64870 137324 79750
rect 137388 79750 137462 79778
rect 137618 79778 137646 80036
rect 137710 79937 137738 80036
rect 137696 79928 137752 79937
rect 137696 79863 137752 79872
rect 137802 79778 137830 80036
rect 137618 79750 137692 79778
rect 137388 79694 137416 79750
rect 137376 79688 137428 79694
rect 137376 79630 137428 79636
rect 137468 79688 137520 79694
rect 137468 79630 137520 79636
rect 137558 79656 137614 79665
rect 137480 71738 137508 79630
rect 137558 79591 137614 79600
rect 137572 76702 137600 79591
rect 137664 77246 137692 79750
rect 137756 79750 137830 79778
rect 137894 79778 137922 80036
rect 137986 79966 138014 80036
rect 137974 79960 138026 79966
rect 138078 79937 138106 80036
rect 137974 79902 138026 79908
rect 138064 79928 138120 79937
rect 138064 79863 138120 79872
rect 138170 79778 138198 80036
rect 138262 79898 138290 80036
rect 138250 79892 138302 79898
rect 138250 79834 138302 79840
rect 138354 79778 138382 80036
rect 138446 79898 138474 80036
rect 138434 79892 138486 79898
rect 138434 79834 138486 79840
rect 137894 79750 138060 79778
rect 137652 77240 137704 77246
rect 137652 77182 137704 77188
rect 137560 76696 137612 76702
rect 137560 76638 137612 76644
rect 137756 76634 137784 79750
rect 137836 79688 137888 79694
rect 137836 79630 137888 79636
rect 137848 77654 137876 79630
rect 137836 77648 137888 77654
rect 137836 77590 137888 77596
rect 137744 76628 137796 76634
rect 137744 76570 137796 76576
rect 138032 75750 138060 79750
rect 138124 79750 138198 79778
rect 138308 79750 138382 79778
rect 138124 76634 138152 79750
rect 138204 79688 138256 79694
rect 138204 79630 138256 79636
rect 138112 76628 138164 76634
rect 138112 76570 138164 76576
rect 138020 75744 138072 75750
rect 138020 75686 138072 75692
rect 138112 72412 138164 72418
rect 138112 72354 138164 72360
rect 137468 71732 137520 71738
rect 137468 71674 137520 71680
rect 138124 70394 138152 72354
rect 138216 71466 138244 79630
rect 138308 77042 138336 79750
rect 138538 79676 138566 80036
rect 138630 79801 138658 80036
rect 138722 79971 138750 80036
rect 138708 79962 138764 79971
rect 138814 79966 138842 80036
rect 138708 79897 138764 79906
rect 138802 79960 138854 79966
rect 138906 79937 138934 80036
rect 138802 79902 138854 79908
rect 138892 79928 138948 79937
rect 138892 79863 138948 79872
rect 138756 79824 138808 79830
rect 138616 79792 138672 79801
rect 138998 79812 139026 80036
rect 139090 79898 139118 80036
rect 139078 79892 139130 79898
rect 139078 79834 139130 79840
rect 139182 79830 139210 80036
rect 138756 79766 138808 79772
rect 138860 79784 139026 79812
rect 139170 79824 139222 79830
rect 138616 79727 138672 79736
rect 138400 79648 138566 79676
rect 138664 79688 138716 79694
rect 138296 77036 138348 77042
rect 138296 76978 138348 76984
rect 138296 76628 138348 76634
rect 138296 76570 138348 76576
rect 138204 71460 138256 71466
rect 138204 71402 138256 71408
rect 138124 70366 138244 70394
rect 138112 66156 138164 66162
rect 138112 66098 138164 66104
rect 138124 65958 138152 66098
rect 138112 65952 138164 65958
rect 138112 65894 138164 65900
rect 137284 64864 137336 64870
rect 137284 64806 137336 64812
rect 137100 56568 137152 56574
rect 137100 56510 137152 56516
rect 136732 42084 136784 42090
rect 136732 42026 136784 42032
rect 138124 39370 138152 65894
rect 138112 39364 138164 39370
rect 138112 39306 138164 39312
rect 136652 16546 137232 16574
rect 135272 6886 135392 6914
rect 133880 4820 133932 4826
rect 133880 4762 133932 4768
rect 131580 3324 131632 3330
rect 131580 3266 131632 3272
rect 134156 3256 134208 3262
rect 134156 3198 134208 3204
rect 132960 2984 133012 2990
rect 132960 2926 133012 2932
rect 132972 480 133000 2926
rect 134168 480 134196 3198
rect 135272 480 135300 6886
rect 136456 3528 136508 3534
rect 136456 3470 136508 3476
rect 136468 480 136496 3470
rect 131734 354 131846 480
rect 131224 326 131846 354
rect 131734 -960 131846 326
rect 132930 -960 133042 480
rect 134126 -960 134238 480
rect 135230 -960 135342 480
rect 136426 -960 136538 480
rect 137204 354 137232 16546
rect 138216 6186 138244 70366
rect 138308 68377 138336 76570
rect 138400 72622 138428 79648
rect 138664 79630 138716 79636
rect 138572 77036 138624 77042
rect 138572 76978 138624 76984
rect 138480 74724 138532 74730
rect 138480 74666 138532 74672
rect 138388 72616 138440 72622
rect 138388 72558 138440 72564
rect 138294 68368 138350 68377
rect 138294 68303 138350 68312
rect 138308 40730 138336 68303
rect 138492 63442 138520 74666
rect 138584 67250 138612 76978
rect 138676 74526 138704 79630
rect 138664 74520 138716 74526
rect 138664 74462 138716 74468
rect 138768 73154 138796 79766
rect 138860 75070 138888 79784
rect 139170 79766 139222 79772
rect 139274 79778 139302 80036
rect 139366 79966 139394 80036
rect 139458 79966 139486 80036
rect 139354 79960 139406 79966
rect 139354 79902 139406 79908
rect 139446 79960 139498 79966
rect 139446 79902 139498 79908
rect 139550 79801 139578 80036
rect 139642 79966 139670 80036
rect 139734 79971 139762 80036
rect 139630 79960 139682 79966
rect 139630 79902 139682 79908
rect 139720 79962 139776 79971
rect 139720 79897 139776 79906
rect 139826 79898 139854 80036
rect 139918 79966 139946 80036
rect 139906 79960 139958 79966
rect 139906 79902 139958 79908
rect 139814 79892 139866 79898
rect 139814 79834 139866 79840
rect 139676 79824 139728 79830
rect 139536 79792 139592 79801
rect 139274 79750 139348 79778
rect 139032 79620 139084 79626
rect 139032 79562 139084 79568
rect 138940 79484 138992 79490
rect 138940 79426 138992 79432
rect 138848 75064 138900 75070
rect 138848 75006 138900 75012
rect 138676 73126 138796 73154
rect 138572 67244 138624 67250
rect 138572 67186 138624 67192
rect 138676 66162 138704 73126
rect 138952 72418 138980 79426
rect 138940 72412 138992 72418
rect 138940 72354 138992 72360
rect 139044 70394 139072 79562
rect 139320 74730 139348 79750
rect 140010 79812 140038 80036
rect 140102 79937 140130 80036
rect 140088 79928 140144 79937
rect 140088 79863 140144 79872
rect 139964 79784 140038 79812
rect 139964 79778 139992 79784
rect 140194 79778 140222 80036
rect 140286 79801 140314 80036
rect 140378 79898 140406 80036
rect 140366 79892 140418 79898
rect 140366 79834 140418 79840
rect 139676 79766 139728 79772
rect 139536 79727 139592 79736
rect 139492 79688 139544 79694
rect 139492 79630 139544 79636
rect 139584 79688 139636 79694
rect 139584 79630 139636 79636
rect 139400 76492 139452 76498
rect 139400 76434 139452 76440
rect 139308 74724 139360 74730
rect 139308 74666 139360 74672
rect 138768 70366 139072 70394
rect 138768 70242 138796 70366
rect 138756 70236 138808 70242
rect 138756 70178 138808 70184
rect 139412 69766 139440 76434
rect 139504 76090 139532 79630
rect 139596 76673 139624 79630
rect 139688 77790 139716 79766
rect 139872 79750 139992 79778
rect 140148 79750 140222 79778
rect 140272 79792 140328 79801
rect 139676 77784 139728 77790
rect 139676 77726 139728 77732
rect 139582 76664 139638 76673
rect 139582 76599 139638 76608
rect 139768 76356 139820 76362
rect 139768 76298 139820 76304
rect 139676 76288 139728 76294
rect 139676 76230 139728 76236
rect 139492 76084 139544 76090
rect 139492 76026 139544 76032
rect 139400 69760 139452 69766
rect 139400 69702 139452 69708
rect 138664 66156 138716 66162
rect 138664 66098 138716 66104
rect 139412 64874 139440 69702
rect 139688 68610 139716 76230
rect 139780 71670 139808 76298
rect 139768 71664 139820 71670
rect 139768 71606 139820 71612
rect 139676 68604 139728 68610
rect 139676 68546 139728 68552
rect 139412 64846 139532 64874
rect 138480 63436 138532 63442
rect 138480 63378 138532 63384
rect 138664 62620 138716 62626
rect 138664 62562 138716 62568
rect 138296 40724 138348 40730
rect 138296 40666 138348 40672
rect 138204 6180 138256 6186
rect 138204 6122 138256 6128
rect 138676 3262 138704 62562
rect 139400 58812 139452 58818
rect 139400 58754 139452 58760
rect 138848 5568 138900 5574
rect 138848 5510 138900 5516
rect 138664 3256 138716 3262
rect 138664 3198 138716 3204
rect 138860 480 138888 5510
rect 139412 490 139440 58754
rect 139504 2990 139532 64846
rect 139872 64734 139900 79750
rect 139952 79552 140004 79558
rect 139952 79494 140004 79500
rect 139964 65822 139992 79494
rect 140044 76628 140096 76634
rect 140044 76570 140096 76576
rect 140056 72894 140084 76570
rect 140044 72888 140096 72894
rect 140044 72830 140096 72836
rect 140148 70038 140176 79750
rect 140470 79778 140498 80036
rect 140562 79966 140590 80036
rect 140550 79960 140602 79966
rect 140550 79902 140602 79908
rect 140654 79812 140682 80036
rect 140746 79966 140774 80036
rect 140838 79966 140866 80036
rect 140734 79960 140786 79966
rect 140734 79902 140786 79908
rect 140826 79960 140878 79966
rect 140826 79902 140878 79908
rect 140930 79812 140958 80036
rect 141022 79966 141050 80036
rect 141114 79971 141142 80036
rect 141010 79960 141062 79966
rect 141010 79902 141062 79908
rect 141100 79962 141156 79971
rect 141100 79897 141156 79906
rect 140654 79784 140728 79812
rect 140884 79801 140958 79812
rect 140424 79762 140498 79778
rect 140272 79727 140328 79736
rect 140412 79756 140498 79762
rect 140464 79750 140498 79756
rect 140412 79698 140464 79704
rect 140228 79688 140280 79694
rect 140596 79688 140648 79694
rect 140228 79630 140280 79636
rect 140318 79656 140374 79665
rect 140240 76362 140268 79630
rect 140596 79630 140648 79636
rect 140318 79591 140374 79600
rect 140228 76356 140280 76362
rect 140228 76298 140280 76304
rect 140332 76226 140360 79591
rect 140412 79552 140464 79558
rect 140412 79494 140464 79500
rect 140424 76634 140452 79494
rect 140504 79484 140556 79490
rect 140504 79426 140556 79432
rect 140412 76628 140464 76634
rect 140412 76570 140464 76576
rect 140320 76220 140372 76226
rect 140320 76162 140372 76168
rect 140228 76084 140280 76090
rect 140228 76026 140280 76032
rect 140136 70032 140188 70038
rect 140136 69974 140188 69980
rect 140240 66094 140268 76026
rect 140516 74118 140544 79426
rect 140608 76294 140636 79630
rect 140596 76288 140648 76294
rect 140596 76230 140648 76236
rect 140504 74112 140556 74118
rect 140504 74054 140556 74060
rect 140700 73778 140728 79784
rect 140870 79792 140958 79801
rect 140926 79784 140958 79792
rect 141206 79778 141234 80036
rect 140870 79727 140926 79736
rect 141068 79750 141234 79778
rect 140872 79688 140924 79694
rect 140870 79656 140872 79665
rect 140964 79688 141016 79694
rect 140924 79656 140926 79665
rect 140964 79630 141016 79636
rect 140870 79591 140926 79600
rect 140976 78470 141004 79630
rect 140964 78464 141016 78470
rect 140964 78406 141016 78412
rect 140964 76220 141016 76226
rect 140964 76162 141016 76168
rect 140688 73772 140740 73778
rect 140688 73714 140740 73720
rect 140780 71664 140832 71670
rect 140780 71606 140832 71612
rect 140792 71058 140820 71606
rect 140780 71052 140832 71058
rect 140780 70994 140832 71000
rect 140228 66088 140280 66094
rect 140228 66030 140280 66036
rect 139952 65816 140004 65822
rect 139952 65758 140004 65764
rect 139860 64728 139912 64734
rect 139860 64670 139912 64676
rect 139964 45554 139992 65758
rect 139596 45526 139992 45554
rect 139596 7614 139624 45526
rect 140792 16574 140820 70994
rect 140976 70922 141004 76162
rect 140964 70916 141016 70922
rect 140964 70858 141016 70864
rect 141068 66910 141096 79750
rect 141148 79688 141200 79694
rect 141298 79676 141326 80036
rect 141390 79744 141418 80036
rect 141482 79898 141510 80036
rect 141574 79937 141602 80036
rect 141666 79966 141694 80036
rect 141654 79960 141706 79966
rect 141560 79928 141616 79937
rect 141470 79892 141522 79898
rect 141654 79902 141706 79908
rect 141560 79863 141616 79872
rect 141470 79834 141522 79840
rect 141514 79792 141570 79801
rect 141390 79716 141464 79744
rect 141514 79727 141570 79736
rect 141608 79756 141660 79762
rect 141148 79630 141200 79636
rect 141252 79648 141326 79676
rect 141056 66904 141108 66910
rect 141056 66846 141108 66852
rect 141160 65550 141188 79630
rect 141252 77586 141280 79648
rect 141332 79552 141384 79558
rect 141332 79494 141384 79500
rect 141240 77580 141292 77586
rect 141240 77522 141292 77528
rect 141238 77480 141294 77489
rect 141238 77415 141294 77424
rect 141252 71126 141280 77415
rect 141240 71120 141292 71126
rect 141240 71062 141292 71068
rect 141344 70394 141372 79494
rect 141436 76226 141464 79716
rect 141424 76220 141476 76226
rect 141424 76162 141476 76168
rect 141528 72350 141556 79727
rect 141758 79744 141786 80036
rect 141850 79966 141878 80036
rect 141942 79966 141970 80036
rect 142034 79966 142062 80036
rect 141838 79960 141890 79966
rect 141838 79902 141890 79908
rect 141930 79960 141982 79966
rect 141930 79902 141982 79908
rect 142022 79960 142074 79966
rect 142126 79937 142154 80036
rect 142218 79966 142246 80036
rect 142310 79971 142338 80036
rect 142206 79960 142258 79966
rect 142022 79902 142074 79908
rect 142112 79928 142168 79937
rect 142206 79902 142258 79908
rect 142296 79962 142352 79971
rect 142402 79966 142430 80036
rect 142494 79966 142522 80036
rect 142586 79966 142614 80036
rect 142296 79897 142352 79906
rect 142390 79960 142442 79966
rect 142390 79902 142442 79908
rect 142482 79960 142534 79966
rect 142482 79902 142534 79908
rect 142574 79960 142626 79966
rect 142574 79902 142626 79908
rect 142112 79863 142168 79872
rect 142068 79824 142120 79830
rect 142068 79766 142120 79772
rect 142388 79826 142444 79835
rect 141608 79698 141660 79704
rect 141712 79716 141786 79744
rect 141620 79472 141648 79698
rect 141712 79626 141740 79716
rect 141882 79656 141938 79665
rect 141700 79620 141752 79626
rect 141882 79591 141938 79600
rect 141700 79562 141752 79568
rect 141620 79444 141740 79472
rect 141712 79370 141740 79444
rect 141712 79342 141832 79370
rect 141698 76800 141754 76809
rect 141698 76735 141754 76744
rect 141712 76362 141740 76735
rect 141700 76356 141752 76362
rect 141700 76298 141752 76304
rect 141516 72344 141568 72350
rect 141516 72286 141568 72292
rect 141712 70394 141740 76298
rect 141804 75410 141832 79342
rect 141896 76498 141924 79591
rect 141976 79552 142028 79558
rect 141976 79494 142028 79500
rect 141884 76492 141936 76498
rect 141884 76434 141936 76440
rect 141988 76158 142016 79494
rect 142080 77897 142108 79766
rect 142160 79756 142212 79762
rect 142388 79761 142444 79770
rect 142678 79744 142706 80036
rect 142770 79778 142798 80036
rect 142862 79966 142890 80036
rect 142850 79960 142902 79966
rect 142850 79902 142902 79908
rect 142770 79750 142844 79778
rect 142160 79698 142212 79704
rect 142632 79716 142706 79744
rect 142066 77888 142122 77897
rect 142066 77823 142122 77832
rect 142172 76430 142200 79698
rect 142252 79688 142304 79694
rect 142252 79630 142304 79636
rect 142528 79688 142580 79694
rect 142632 79665 142660 79716
rect 142528 79630 142580 79636
rect 142618 79656 142674 79665
rect 142160 76424 142212 76430
rect 142160 76366 142212 76372
rect 141976 76152 142028 76158
rect 141976 76094 142028 76100
rect 141792 75404 141844 75410
rect 141792 75346 141844 75352
rect 142160 74520 142212 74526
rect 142160 74462 142212 74468
rect 142172 73914 142200 74462
rect 142160 73908 142212 73914
rect 142160 73850 142212 73856
rect 141252 70366 141372 70394
rect 141436 70366 141740 70394
rect 141148 65544 141200 65550
rect 141148 65486 141200 65492
rect 141252 64190 141280 70366
rect 141240 64184 141292 64190
rect 141240 64126 141292 64132
rect 140792 16546 141280 16574
rect 139584 7608 139636 7614
rect 139584 7550 139636 7556
rect 139492 2984 139544 2990
rect 139492 2926 139544 2932
rect 137622 354 137734 480
rect 137204 326 137734 354
rect 137622 -960 137734 326
rect 138818 -960 138930 480
rect 139412 462 139624 490
rect 141252 480 141280 16546
rect 141436 3466 141464 70366
rect 142172 69018 142200 73850
rect 141516 69012 141568 69018
rect 141516 68954 141568 68960
rect 142160 69012 142212 69018
rect 142160 68954 142212 68960
rect 141528 3534 141556 68954
rect 142160 68672 142212 68678
rect 142160 68614 142212 68620
rect 142172 58818 142200 68614
rect 142160 58812 142212 58818
rect 142160 58754 142212 58760
rect 142264 45626 142292 79630
rect 142344 79552 142396 79558
rect 142344 79494 142396 79500
rect 142356 78169 142384 79494
rect 142540 78962 142568 79630
rect 142618 79591 142674 79600
rect 142620 79552 142672 79558
rect 142620 79494 142672 79500
rect 142712 79552 142764 79558
rect 142712 79494 142764 79500
rect 142448 78934 142568 78962
rect 142448 78674 142476 78934
rect 142632 78792 142660 79494
rect 142540 78764 142660 78792
rect 142436 78668 142488 78674
rect 142436 78610 142488 78616
rect 142342 78160 142398 78169
rect 142342 78095 142398 78104
rect 142540 77722 142568 78764
rect 142618 78704 142674 78713
rect 142618 78639 142674 78648
rect 142528 77716 142580 77722
rect 142528 77658 142580 77664
rect 142344 74452 142396 74458
rect 142344 74394 142396 74400
rect 142356 73234 142384 74394
rect 142344 73228 142396 73234
rect 142344 73170 142396 73176
rect 142344 73024 142396 73030
rect 142344 72966 142396 72972
rect 142356 72690 142384 72966
rect 142344 72684 142396 72690
rect 142344 72626 142396 72632
rect 142356 68678 142384 72626
rect 142436 71732 142488 71738
rect 142436 71674 142488 71680
rect 142448 71262 142476 71674
rect 142436 71256 142488 71262
rect 142436 71198 142488 71204
rect 142344 68672 142396 68678
rect 142344 68614 142396 68620
rect 142448 68542 142476 71198
rect 142528 69828 142580 69834
rect 142528 69770 142580 69776
rect 142436 68536 142488 68542
rect 142436 68478 142488 68484
rect 142540 68354 142568 69770
rect 142356 68326 142568 68354
rect 142356 55282 142384 68326
rect 142436 68264 142488 68270
rect 142436 68206 142488 68212
rect 142448 62626 142476 68206
rect 142632 67522 142660 78639
rect 142724 68746 142752 79494
rect 142816 74534 142844 79750
rect 142954 79744 142982 80036
rect 143046 79898 143074 80036
rect 143138 79937 143166 80036
rect 143124 79928 143180 79937
rect 143034 79892 143086 79898
rect 143124 79863 143180 79872
rect 143034 79834 143086 79840
rect 143230 79830 143258 80036
rect 143322 79971 143350 80036
rect 143308 79962 143364 79971
rect 143308 79897 143364 79906
rect 143414 79898 143442 80036
rect 143402 79892 143454 79898
rect 143402 79834 143454 79840
rect 143218 79824 143270 79830
rect 143218 79766 143270 79772
rect 143506 79744 143534 80036
rect 143598 79801 143626 80036
rect 142954 79716 143028 79744
rect 143000 77450 143028 79716
rect 143460 79716 143534 79744
rect 143584 79792 143640 79801
rect 143584 79727 143640 79736
rect 143080 79688 143132 79694
rect 143080 79630 143132 79636
rect 143172 79688 143224 79694
rect 143172 79630 143224 79636
rect 143262 79656 143318 79665
rect 142988 77444 143040 77450
rect 142988 77386 143040 77392
rect 142896 76968 142948 76974
rect 142896 76910 142948 76916
rect 142908 76634 142936 76910
rect 142896 76628 142948 76634
rect 142896 76570 142948 76576
rect 142816 74506 143028 74534
rect 142804 74452 142856 74458
rect 142804 74394 142856 74400
rect 142816 74254 142844 74394
rect 142804 74248 142856 74254
rect 142804 74190 142856 74196
rect 142712 68740 142764 68746
rect 142712 68682 142764 68688
rect 142620 67516 142672 67522
rect 142620 67458 142672 67464
rect 142632 64874 142660 67458
rect 142540 64846 142660 64874
rect 142436 62620 142488 62626
rect 142436 62562 142488 62568
rect 142344 55276 142396 55282
rect 142344 55218 142396 55224
rect 142252 45620 142304 45626
rect 142252 45562 142304 45568
rect 142540 5574 142568 64846
rect 142724 6914 142752 68682
rect 142632 6886 142752 6914
rect 142528 5568 142580 5574
rect 142528 5510 142580 5516
rect 141516 3528 141568 3534
rect 142632 3482 142660 6886
rect 142816 5574 142844 74190
rect 143000 71738 143028 74506
rect 142988 71732 143040 71738
rect 142988 71674 143040 71680
rect 143092 69834 143120 79630
rect 143184 73030 143212 79630
rect 143262 79591 143318 79600
rect 143276 78792 143304 79591
rect 143276 78764 143396 78792
rect 143264 77444 143316 77450
rect 143264 77386 143316 77392
rect 143276 74526 143304 77386
rect 143264 74520 143316 74526
rect 143264 74462 143316 74468
rect 143172 73024 143224 73030
rect 143172 72966 143224 72972
rect 143368 71670 143396 78764
rect 143460 74458 143488 79716
rect 143540 79620 143592 79626
rect 143690 79608 143718 80036
rect 143782 79830 143810 80036
rect 143770 79824 143822 79830
rect 143770 79766 143822 79772
rect 143874 79642 143902 80036
rect 143966 79966 143994 80036
rect 144058 79966 144086 80036
rect 143954 79960 144006 79966
rect 143954 79902 144006 79908
rect 144046 79960 144098 79966
rect 144046 79902 144098 79908
rect 143966 79744 143994 79902
rect 144150 79778 144178 80036
rect 144242 79966 144270 80036
rect 144230 79960 144282 79966
rect 144230 79902 144282 79908
rect 144334 79830 144362 80036
rect 144426 79898 144454 80036
rect 144518 79898 144546 80036
rect 144610 79937 144638 80036
rect 144596 79928 144652 79937
rect 144414 79892 144466 79898
rect 144414 79834 144466 79840
rect 144506 79892 144558 79898
rect 144702 79898 144730 80036
rect 144596 79863 144652 79872
rect 144690 79892 144742 79898
rect 144506 79834 144558 79840
rect 144690 79834 144742 79840
rect 144322 79824 144374 79830
rect 144150 79750 144224 79778
rect 144322 79766 144374 79772
rect 144550 79792 144606 79801
rect 143966 79716 144040 79744
rect 143874 79614 143948 79642
rect 143690 79580 143764 79608
rect 143540 79562 143592 79568
rect 143552 76702 143580 79562
rect 143632 79348 143684 79354
rect 143632 79290 143684 79296
rect 143540 76696 143592 76702
rect 143540 76638 143592 76644
rect 143448 74452 143500 74458
rect 143448 74394 143500 74400
rect 143448 74248 143500 74254
rect 143448 74190 143500 74196
rect 143356 71664 143408 71670
rect 143356 71606 143408 71612
rect 143080 69828 143132 69834
rect 143080 69770 143132 69776
rect 142804 5568 142856 5574
rect 142804 5510 142856 5516
rect 141516 3470 141568 3476
rect 141424 3460 141476 3466
rect 141424 3402 141476 3408
rect 142448 3454 142660 3482
rect 142448 480 142476 3454
rect 143460 3398 143488 74190
rect 143540 69896 143592 69902
rect 143540 69838 143592 69844
rect 143552 5710 143580 69838
rect 143644 19990 143672 79290
rect 143736 78810 143764 79580
rect 143816 79552 143868 79558
rect 143816 79494 143868 79500
rect 143724 78804 143776 78810
rect 143724 78746 143776 78752
rect 143828 76566 143856 79494
rect 143816 76560 143868 76566
rect 143816 76502 143868 76508
rect 143828 74254 143856 76502
rect 143816 74248 143868 74254
rect 143816 74190 143868 74196
rect 143920 70394 143948 79614
rect 144012 76838 144040 79716
rect 144196 77625 144224 79750
rect 144550 79727 144606 79736
rect 144644 79756 144696 79762
rect 144276 79688 144328 79694
rect 144276 79630 144328 79636
rect 144368 79688 144420 79694
rect 144368 79630 144420 79636
rect 144182 77616 144238 77625
rect 144182 77551 144238 77560
rect 144000 76832 144052 76838
rect 144000 76774 144052 76780
rect 144092 76696 144144 76702
rect 144092 76638 144144 76644
rect 144104 74186 144132 76638
rect 144184 76152 144236 76158
rect 144184 76094 144236 76100
rect 144196 75138 144224 76094
rect 144288 75614 144316 79630
rect 144380 79354 144408 79630
rect 144460 79620 144512 79626
rect 144460 79562 144512 79568
rect 144368 79348 144420 79354
rect 144368 79290 144420 79296
rect 144472 77897 144500 79562
rect 144564 79422 144592 79727
rect 144644 79698 144696 79704
rect 144552 79416 144604 79422
rect 144552 79358 144604 79364
rect 144552 78804 144604 78810
rect 144552 78746 144604 78752
rect 144458 77888 144514 77897
rect 144458 77823 144514 77832
rect 144458 77752 144514 77761
rect 144458 77687 144514 77696
rect 144276 75608 144328 75614
rect 144276 75550 144328 75556
rect 144184 75132 144236 75138
rect 144184 75074 144236 75080
rect 144092 74180 144144 74186
rect 144092 74122 144144 74128
rect 144104 71738 144132 74122
rect 144092 71732 144144 71738
rect 144092 71674 144144 71680
rect 143920 70366 144040 70394
rect 144012 68950 144040 70366
rect 144000 68944 144052 68950
rect 144000 68886 144052 68892
rect 143632 19984 143684 19990
rect 143632 19926 143684 19932
rect 144196 6186 144224 75074
rect 144288 73154 144316 75550
rect 144288 73126 144408 73154
rect 144276 68808 144328 68814
rect 144276 68750 144328 68756
rect 144288 30326 144316 68750
rect 144380 63238 144408 73126
rect 144472 69902 144500 77687
rect 144460 69896 144512 69902
rect 144460 69838 144512 69844
rect 144460 68944 144512 68950
rect 144460 68886 144512 68892
rect 144472 63578 144500 68886
rect 144564 68814 144592 78746
rect 144656 74769 144684 79698
rect 144794 79642 144822 80036
rect 144886 79830 144914 80036
rect 144874 79824 144926 79830
rect 144874 79766 144926 79772
rect 144978 79744 145006 80036
rect 145070 79937 145098 80036
rect 145162 79966 145190 80036
rect 145254 79971 145282 80036
rect 145150 79960 145202 79966
rect 145056 79928 145112 79937
rect 145150 79902 145202 79908
rect 145240 79962 145296 79971
rect 145346 79966 145374 80036
rect 145240 79897 145296 79906
rect 145334 79960 145386 79966
rect 145438 79937 145466 80036
rect 145530 79966 145558 80036
rect 145518 79960 145570 79966
rect 145334 79902 145386 79908
rect 145424 79928 145480 79937
rect 145056 79863 145112 79872
rect 145196 79824 145248 79830
rect 145196 79766 145248 79772
rect 145104 79756 145156 79762
rect 144978 79716 145052 79744
rect 144794 79614 144868 79642
rect 144736 79552 144788 79558
rect 144736 79494 144788 79500
rect 144642 74760 144698 74769
rect 144642 74695 144698 74704
rect 144748 73234 144776 79494
rect 144840 76673 144868 79614
rect 144920 79620 144972 79626
rect 144920 79562 144972 79568
rect 144826 76664 144882 76673
rect 144826 76599 144882 76608
rect 144932 76158 144960 79562
rect 145024 78742 145052 79716
rect 145104 79698 145156 79704
rect 145012 78736 145064 78742
rect 145012 78678 145064 78684
rect 144920 76152 144972 76158
rect 144920 76094 144972 76100
rect 145116 73846 145144 79698
rect 145104 73840 145156 73846
rect 145104 73782 145156 73788
rect 145012 73636 145064 73642
rect 145012 73578 145064 73584
rect 144736 73228 144788 73234
rect 144736 73170 144788 73176
rect 144552 68808 144604 68814
rect 144552 68750 144604 68756
rect 144460 63572 144512 63578
rect 144460 63514 144512 63520
rect 144368 63232 144420 63238
rect 144368 63174 144420 63180
rect 144276 30320 144328 30326
rect 144276 30262 144328 30268
rect 145024 25566 145052 73578
rect 145208 49026 145236 79766
rect 145346 79744 145374 79902
rect 145518 79902 145570 79908
rect 145424 79863 145480 79872
rect 145470 79792 145526 79801
rect 145346 79716 145420 79744
rect 145622 79778 145650 80036
rect 145714 79898 145742 80036
rect 145702 79892 145754 79898
rect 145702 79834 145754 79840
rect 145806 79778 145834 80036
rect 145898 79937 145926 80036
rect 145884 79928 145940 79937
rect 145884 79863 145940 79872
rect 145622 79750 145696 79778
rect 145470 79727 145526 79736
rect 145288 79416 145340 79422
rect 145288 79358 145340 79364
rect 145300 70394 145328 79358
rect 145392 74458 145420 79716
rect 145484 79608 145512 79727
rect 145484 79580 145604 79608
rect 145472 79484 145524 79490
rect 145472 79426 145524 79432
rect 145484 75274 145512 79426
rect 145576 75546 145604 79580
rect 145668 76906 145696 79750
rect 145760 79750 145834 79778
rect 145760 79150 145788 79750
rect 145990 79744 146018 80036
rect 146082 79898 146110 80036
rect 146174 79898 146202 80036
rect 146266 79966 146294 80036
rect 146254 79960 146306 79966
rect 146254 79902 146306 79908
rect 146358 79903 146386 80036
rect 146070 79892 146122 79898
rect 146070 79834 146122 79840
rect 146162 79892 146214 79898
rect 146162 79834 146214 79840
rect 146344 79894 146400 79903
rect 146450 79898 146478 80036
rect 146174 79801 146202 79834
rect 146344 79829 146400 79838
rect 146438 79892 146490 79898
rect 146438 79834 146490 79840
rect 146160 79792 146216 79801
rect 145990 79716 146064 79744
rect 146542 79778 146570 80036
rect 146634 79898 146662 80036
rect 146726 79971 146754 80036
rect 146712 79962 146768 79971
rect 146818 79966 146846 80036
rect 146622 79892 146674 79898
rect 146712 79897 146768 79906
rect 146806 79960 146858 79966
rect 146806 79902 146858 79908
rect 146910 79898 146938 80036
rect 146622 79834 146674 79840
rect 146898 79892 146950 79898
rect 146898 79834 146950 79840
rect 146666 79792 146722 79801
rect 146160 79727 146216 79736
rect 146300 79756 146352 79762
rect 145840 79688 145892 79694
rect 145840 79630 145892 79636
rect 145930 79656 145986 79665
rect 145748 79144 145800 79150
rect 145748 79086 145800 79092
rect 145656 76900 145708 76906
rect 145656 76842 145708 76848
rect 145564 75540 145616 75546
rect 145564 75482 145616 75488
rect 145472 75268 145524 75274
rect 145472 75210 145524 75216
rect 145484 74934 145512 75210
rect 145472 74928 145524 74934
rect 145472 74870 145524 74876
rect 145380 74452 145432 74458
rect 145380 74394 145432 74400
rect 145300 70366 145420 70394
rect 145392 64874 145420 70366
rect 145300 64846 145420 64874
rect 145300 60246 145328 64846
rect 145288 60240 145340 60246
rect 145288 60182 145340 60188
rect 145196 49020 145248 49026
rect 145196 48962 145248 48968
rect 145576 31074 145604 75482
rect 145668 57254 145696 76842
rect 145760 73642 145788 79086
rect 145852 76945 145880 79630
rect 145930 79591 145986 79600
rect 145838 76936 145894 76945
rect 145838 76871 145894 76880
rect 145852 76673 145880 76871
rect 145838 76664 145894 76673
rect 145838 76599 145894 76608
rect 145748 73636 145800 73642
rect 145748 73578 145800 73584
rect 145656 57248 145708 57254
rect 145656 57190 145708 57196
rect 145564 31068 145616 31074
rect 145564 31010 145616 31016
rect 145104 30320 145156 30326
rect 145104 30262 145156 30268
rect 145012 25560 145064 25566
rect 145012 25502 145064 25508
rect 145116 16574 145144 30262
rect 145944 29714 145972 79591
rect 146036 76362 146064 79716
rect 146542 79750 146616 79778
rect 146352 79716 146432 79744
rect 146300 79698 146352 79704
rect 146298 79656 146354 79665
rect 146116 79620 146168 79626
rect 146298 79591 146354 79600
rect 146116 79562 146168 79568
rect 146128 79218 146156 79562
rect 146312 79422 146340 79591
rect 146404 79558 146432 79716
rect 146484 79688 146536 79694
rect 146484 79630 146536 79636
rect 146392 79552 146444 79558
rect 146392 79494 146444 79500
rect 146300 79416 146352 79422
rect 146300 79358 146352 79364
rect 146116 79212 146168 79218
rect 146116 79154 146168 79160
rect 146024 76356 146076 76362
rect 146024 76298 146076 76304
rect 146208 75812 146260 75818
rect 146208 75754 146260 75760
rect 146220 75070 146248 75754
rect 146208 75064 146260 75070
rect 146208 75006 146260 75012
rect 146024 74452 146076 74458
rect 146024 74394 146076 74400
rect 145932 29708 145984 29714
rect 145932 29650 145984 29656
rect 146036 17270 146064 74394
rect 146404 73914 146432 79494
rect 146496 75818 146524 79630
rect 146484 75812 146536 75818
rect 146484 75754 146536 75760
rect 146588 75206 146616 79750
rect 146852 79756 146904 79762
rect 146666 79727 146722 79736
rect 146680 77178 146708 79727
rect 146772 79716 146852 79744
rect 146668 77172 146720 77178
rect 146668 77114 146720 77120
rect 146772 76634 146800 79716
rect 146852 79698 146904 79704
rect 147002 79676 147030 80036
rect 147094 79937 147122 80036
rect 147080 79928 147136 79937
rect 147186 79898 147214 80036
rect 147278 79971 147306 80036
rect 147264 79962 147320 79971
rect 147080 79863 147136 79872
rect 147174 79892 147226 79898
rect 147264 79897 147320 79906
rect 147174 79834 147226 79840
rect 147370 79830 147398 80036
rect 147462 79971 147490 80036
rect 147448 79962 147504 79971
rect 147448 79897 147504 79906
rect 147554 79898 147582 80036
rect 147646 79937 147674 80036
rect 147738 79966 147766 80036
rect 147830 79966 147858 80036
rect 147922 79966 147950 80036
rect 147726 79960 147778 79966
rect 147632 79928 147688 79937
rect 147542 79892 147594 79898
rect 147726 79902 147778 79908
rect 147818 79960 147870 79966
rect 147818 79902 147870 79908
rect 147910 79960 147962 79966
rect 147910 79902 147962 79908
rect 147632 79863 147688 79872
rect 147542 79834 147594 79840
rect 148014 79830 148042 80036
rect 148106 79830 148134 80036
rect 147358 79824 147410 79830
rect 147358 79766 147410 79772
rect 148002 79824 148054 79830
rect 148002 79766 148054 79772
rect 148094 79824 148146 79830
rect 148094 79766 148146 79772
rect 147128 79756 147180 79762
rect 147128 79698 147180 79704
rect 147220 79756 147272 79762
rect 147220 79698 147272 79704
rect 147772 79756 147824 79762
rect 148198 79744 148226 80036
rect 148290 79898 148318 80036
rect 148278 79892 148330 79898
rect 148278 79834 148330 79840
rect 148382 79812 148410 80036
rect 148474 79966 148502 80036
rect 148566 79971 148594 80036
rect 148462 79960 148514 79966
rect 148462 79902 148514 79908
rect 148552 79962 148608 79971
rect 148552 79897 148608 79906
rect 148508 79824 148560 79830
rect 148382 79784 148456 79812
rect 148198 79716 148364 79744
rect 147772 79698 147824 79704
rect 146956 79648 147030 79676
rect 146852 79620 146904 79626
rect 146852 79562 146904 79568
rect 146864 79529 146892 79562
rect 146850 79520 146906 79529
rect 146850 79455 146906 79464
rect 146760 76628 146812 76634
rect 146760 76570 146812 76576
rect 146576 75200 146628 75206
rect 146576 75142 146628 75148
rect 146392 73908 146444 73914
rect 146392 73850 146444 73856
rect 146300 71732 146352 71738
rect 146300 71674 146352 71680
rect 146024 17264 146076 17270
rect 146024 17206 146076 17212
rect 146312 16574 146340 71674
rect 146588 71194 146616 75142
rect 146576 71188 146628 71194
rect 146576 71130 146628 71136
rect 146864 70394 146892 79455
rect 146956 76673 146984 79648
rect 147140 78946 147168 79698
rect 147232 79014 147260 79698
rect 147312 79688 147364 79694
rect 147312 79630 147364 79636
rect 147220 79008 147272 79014
rect 147220 78950 147272 78956
rect 147128 78940 147180 78946
rect 147128 78882 147180 78888
rect 147034 78704 147090 78713
rect 147034 78639 147090 78648
rect 147048 76974 147076 78639
rect 147140 77294 147168 78882
rect 147140 77266 147260 77294
rect 147036 76968 147088 76974
rect 147088 76928 147168 76956
rect 147036 76910 147088 76916
rect 147036 76832 147088 76838
rect 147036 76774 147088 76780
rect 146942 76664 146998 76673
rect 146942 76599 146998 76608
rect 146944 73908 146996 73914
rect 146944 73850 146996 73856
rect 146496 70366 146892 70394
rect 146496 64874 146524 70366
rect 146404 64846 146524 64874
rect 146404 64190 146432 64846
rect 146392 64184 146444 64190
rect 146392 64126 146444 64132
rect 145116 16546 145512 16574
rect 146312 16546 146892 16574
rect 144184 6180 144236 6186
rect 144184 6122 144236 6128
rect 143540 5704 143592 5710
rect 143540 5646 143592 5652
rect 144736 5704 144788 5710
rect 144736 5646 144788 5652
rect 143540 5568 143592 5574
rect 143540 5510 143592 5516
rect 143448 3392 143500 3398
rect 143448 3334 143500 3340
rect 143552 480 143580 5510
rect 144748 480 144776 5646
rect 139596 354 139624 462
rect 140014 354 140126 480
rect 139596 326 140126 354
rect 140014 -960 140126 326
rect 141210 -960 141322 480
rect 142406 -960 142518 480
rect 143510 -960 143622 480
rect 144706 -960 144818 480
rect 145484 354 145512 16546
rect 146864 3482 146892 16546
rect 146956 4010 146984 73850
rect 146944 4004 146996 4010
rect 146944 3946 146996 3952
rect 147048 3738 147076 76774
rect 147140 71126 147168 76928
rect 147232 76702 147260 77266
rect 147220 76696 147272 76702
rect 147220 76638 147272 76644
rect 147324 75682 147352 79630
rect 147680 79552 147732 79558
rect 147680 79494 147732 79500
rect 147496 79212 147548 79218
rect 147496 79154 147548 79160
rect 147404 79008 147456 79014
rect 147404 78950 147456 78956
rect 147312 75676 147364 75682
rect 147312 75618 147364 75624
rect 147220 75268 147272 75274
rect 147220 75210 147272 75216
rect 147128 71120 147180 71126
rect 147128 71062 147180 71068
rect 147232 70394 147260 75210
rect 147140 70366 147260 70394
rect 147140 3942 147168 70366
rect 147324 68338 147352 75618
rect 147416 75274 147444 78950
rect 147404 75268 147456 75274
rect 147404 75210 147456 75216
rect 147508 73154 147536 79154
rect 147416 73126 147536 73154
rect 147416 70394 147444 73126
rect 147692 72758 147720 79494
rect 147784 78878 147812 79698
rect 147956 79688 148008 79694
rect 147956 79630 148008 79636
rect 147864 79484 147916 79490
rect 147864 79426 147916 79432
rect 147772 78872 147824 78878
rect 147772 78814 147824 78820
rect 147680 72752 147732 72758
rect 147680 72694 147732 72700
rect 147416 70366 147628 70394
rect 147600 69698 147628 70366
rect 147588 69692 147640 69698
rect 147588 69634 147640 69640
rect 147312 68332 147364 68338
rect 147312 68274 147364 68280
rect 147220 63572 147272 63578
rect 147220 63514 147272 63520
rect 147128 3936 147180 3942
rect 147128 3878 147180 3884
rect 147036 3732 147088 3738
rect 147036 3674 147088 3680
rect 147232 3534 147260 63514
rect 147784 61402 147812 78814
rect 147876 70394 147904 79426
rect 147968 76770 147996 79630
rect 148140 79552 148192 79558
rect 148140 79494 148192 79500
rect 148048 79484 148100 79490
rect 148048 79426 148100 79432
rect 147956 76764 148008 76770
rect 147956 76706 148008 76712
rect 148060 74534 148088 79426
rect 148152 78674 148180 79494
rect 148336 79354 148364 79716
rect 148428 79490 148456 79784
rect 148658 79801 148686 80036
rect 148750 79898 148778 80036
rect 148842 79898 148870 80036
rect 148738 79892 148790 79898
rect 148738 79834 148790 79840
rect 148830 79892 148882 79898
rect 148830 79834 148882 79840
rect 148508 79766 148560 79772
rect 148644 79792 148700 79801
rect 148416 79484 148468 79490
rect 148416 79426 148468 79432
rect 148520 79370 148548 79766
rect 148934 79778 148962 80036
rect 149026 79966 149054 80036
rect 149014 79960 149066 79966
rect 149014 79902 149066 79908
rect 148644 79727 148700 79736
rect 148842 79750 148962 79778
rect 148600 79688 148652 79694
rect 148842 79676 148870 79750
rect 149118 79744 149146 80036
rect 149210 79966 149238 80036
rect 149198 79960 149250 79966
rect 149198 79902 149250 79908
rect 149302 79898 149330 80036
rect 149394 79971 149422 80036
rect 149380 79962 149436 79971
rect 149486 79966 149514 80036
rect 149290 79892 149342 79898
rect 149380 79897 149436 79906
rect 149474 79960 149526 79966
rect 149578 79937 149606 80036
rect 149474 79902 149526 79908
rect 149564 79928 149620 79937
rect 149564 79863 149620 79872
rect 149290 79834 149342 79840
rect 149382 79824 149434 79830
rect 149670 79812 149698 80036
rect 149762 79966 149790 80036
rect 149750 79960 149802 79966
rect 149750 79902 149802 79908
rect 149854 79812 149882 80036
rect 149946 79966 149974 80036
rect 150038 79966 150066 80036
rect 150130 79966 150158 80036
rect 150222 79966 150250 80036
rect 150314 79971 150342 80036
rect 149934 79960 149986 79966
rect 149934 79902 149986 79908
rect 150026 79960 150078 79966
rect 150026 79902 150078 79908
rect 150118 79960 150170 79966
rect 150118 79902 150170 79908
rect 150210 79960 150262 79966
rect 150210 79902 150262 79908
rect 150300 79962 150356 79971
rect 150300 79897 150356 79906
rect 149434 79784 149560 79812
rect 149670 79784 149744 79812
rect 149382 79766 149434 79772
rect 149118 79716 149192 79744
rect 148968 79688 149020 79694
rect 148652 79648 148732 79676
rect 148842 79648 148916 79676
rect 148600 79630 148652 79636
rect 148600 79552 148652 79558
rect 148600 79494 148652 79500
rect 148324 79348 148376 79354
rect 148324 79290 148376 79296
rect 148428 79342 148548 79370
rect 148152 78646 148272 78674
rect 148244 75886 148272 78646
rect 148428 77489 148456 79342
rect 148414 77480 148470 77489
rect 148414 77415 148470 77424
rect 148612 77353 148640 79494
rect 148704 78130 148732 79648
rect 148888 79558 148916 79648
rect 148968 79630 149020 79636
rect 148876 79552 148928 79558
rect 148876 79494 148928 79500
rect 148784 79484 148836 79490
rect 148784 79426 148836 79432
rect 148692 78124 148744 78130
rect 148692 78066 148744 78072
rect 148598 77344 148654 77353
rect 148598 77279 148654 77288
rect 148704 77228 148732 78066
rect 148612 77200 148732 77228
rect 148508 77172 148560 77178
rect 148508 77114 148560 77120
rect 148232 75880 148284 75886
rect 148232 75822 148284 75828
rect 148520 75342 148548 77114
rect 148508 75336 148560 75342
rect 148508 75278 148560 75284
rect 148060 74506 148180 74534
rect 148152 72486 148180 74506
rect 148140 72480 148192 72486
rect 148140 72422 148192 72428
rect 147876 70366 147996 70394
rect 147968 67590 147996 70366
rect 147956 67584 148008 67590
rect 147956 67526 148008 67532
rect 147772 61396 147824 61402
rect 147772 61338 147824 61344
rect 147968 60382 147996 67526
rect 148152 65754 148180 72422
rect 148508 67448 148560 67454
rect 148508 67390 148560 67396
rect 148140 65748 148192 65754
rect 148140 65690 148192 65696
rect 148324 63232 148376 63238
rect 148324 63174 148376 63180
rect 147956 60376 148008 60382
rect 147956 60318 148008 60324
rect 148336 4146 148364 63174
rect 148416 60240 148468 60246
rect 148416 60182 148468 60188
rect 148324 4140 148376 4146
rect 148324 4082 148376 4088
rect 148428 3874 148456 60182
rect 148520 36854 148548 67390
rect 148612 49162 148640 77200
rect 148692 76764 148744 76770
rect 148692 76706 148744 76712
rect 148704 53242 148732 76706
rect 148796 67454 148824 79426
rect 148874 79384 148930 79393
rect 148874 79319 148930 79328
rect 148888 74534 148916 79319
rect 148980 77217 149008 79630
rect 149060 79620 149112 79626
rect 149060 79562 149112 79568
rect 148966 77208 149022 77217
rect 148966 77143 149022 77152
rect 148888 74506 149008 74534
rect 148876 72752 148928 72758
rect 148876 72694 148928 72700
rect 148888 71058 148916 72694
rect 148876 71052 148928 71058
rect 148876 70994 148928 71000
rect 148784 67448 148836 67454
rect 148784 67390 148836 67396
rect 148692 53236 148744 53242
rect 148692 53178 148744 53184
rect 148600 49156 148652 49162
rect 148600 49098 148652 49104
rect 148508 36848 148560 36854
rect 148508 36790 148560 36796
rect 148980 32706 149008 74506
rect 149072 67386 149100 79562
rect 149164 71534 149192 79716
rect 149336 79688 149388 79694
rect 149336 79630 149388 79636
rect 149428 79688 149480 79694
rect 149428 79630 149480 79636
rect 149348 77654 149376 79630
rect 149336 77648 149388 77654
rect 149336 77590 149388 77596
rect 149336 71732 149388 71738
rect 149336 71674 149388 71680
rect 149348 71602 149376 71674
rect 149336 71596 149388 71602
rect 149336 71538 149388 71544
rect 149152 71528 149204 71534
rect 149152 71470 149204 71476
rect 149164 70854 149192 71470
rect 149152 70848 149204 70854
rect 149152 70790 149204 70796
rect 149348 70394 149376 71538
rect 149440 71330 149468 79630
rect 149532 79268 149560 79784
rect 149612 79688 149664 79694
rect 149612 79630 149664 79636
rect 149624 79393 149652 79630
rect 149610 79384 149666 79393
rect 149610 79319 149666 79328
rect 149532 79240 149652 79268
rect 149518 78568 149574 78577
rect 149518 78503 149574 78512
rect 149428 71324 149480 71330
rect 149428 71266 149480 71272
rect 149440 70786 149468 71266
rect 149428 70780 149480 70786
rect 149428 70722 149480 70728
rect 149348 70366 149468 70394
rect 149060 67380 149112 67386
rect 149060 67322 149112 67328
rect 149440 55962 149468 70366
rect 149428 55956 149480 55962
rect 149428 55898 149480 55904
rect 149532 47598 149560 78503
rect 149624 78266 149652 79240
rect 149612 78260 149664 78266
rect 149612 78202 149664 78208
rect 149716 74322 149744 79784
rect 149808 79784 149882 79812
rect 149704 74316 149756 74322
rect 149704 74258 149756 74264
rect 149610 74080 149666 74089
rect 149610 74015 149666 74024
rect 149624 60314 149652 74015
rect 149704 73228 149756 73234
rect 149704 73170 149756 73176
rect 149612 60308 149664 60314
rect 149612 60250 149664 60256
rect 149520 47592 149572 47598
rect 149520 47534 149572 47540
rect 148968 32700 149020 32706
rect 148968 32642 149020 32648
rect 149716 4010 149744 73170
rect 149808 72554 149836 79784
rect 149888 79688 149940 79694
rect 149888 79630 149940 79636
rect 150256 79688 150308 79694
rect 150406 79676 150434 80036
rect 150256 79630 150308 79636
rect 150360 79648 150434 79676
rect 150498 79676 150526 80036
rect 150590 79744 150618 80036
rect 150682 79966 150710 80036
rect 150774 79966 150802 80036
rect 150670 79960 150722 79966
rect 150670 79902 150722 79908
rect 150762 79960 150814 79966
rect 150762 79902 150814 79908
rect 150716 79824 150768 79830
rect 150866 79812 150894 80036
rect 150958 79830 150986 80036
rect 151050 79898 151078 80036
rect 151038 79892 151090 79898
rect 151038 79834 151090 79840
rect 151142 79830 151170 80036
rect 151234 79937 151262 80036
rect 151326 79966 151354 80036
rect 151418 79966 151446 80036
rect 151314 79960 151366 79966
rect 151220 79928 151276 79937
rect 151314 79902 151366 79908
rect 151406 79960 151458 79966
rect 151406 79902 151458 79908
rect 151220 79863 151276 79872
rect 150716 79766 150768 79772
rect 150820 79784 150894 79812
rect 150946 79824 150998 79830
rect 150590 79716 150664 79744
rect 150498 79648 150572 79676
rect 149796 72548 149848 72554
rect 149796 72490 149848 72496
rect 149808 72010 149836 72490
rect 149796 72004 149848 72010
rect 149796 71946 149848 71952
rect 149900 71505 149928 79630
rect 150164 79620 150216 79626
rect 150164 79562 150216 79568
rect 150072 79552 150124 79558
rect 150072 79494 150124 79500
rect 150084 79082 150112 79494
rect 150072 79076 150124 79082
rect 150072 79018 150124 79024
rect 150084 76634 150112 79018
rect 150072 76628 150124 76634
rect 150072 76570 150124 76576
rect 149980 74316 150032 74322
rect 149980 74258 150032 74264
rect 149886 71496 149942 71505
rect 149886 71431 149942 71440
rect 149900 70394 149928 71431
rect 149808 70366 149928 70394
rect 149808 12034 149836 70366
rect 149888 67380 149940 67386
rect 149888 67322 149940 67328
rect 149796 12028 149848 12034
rect 149796 11970 149848 11976
rect 149900 9246 149928 67322
rect 149992 31346 150020 74258
rect 150176 71738 150204 79562
rect 150268 77353 150296 79630
rect 150254 77344 150310 77353
rect 150254 77279 150310 77288
rect 150360 74089 150388 79648
rect 150544 79370 150572 79648
rect 150452 79342 150572 79370
rect 150346 74080 150402 74089
rect 150346 74015 150402 74024
rect 150256 72004 150308 72010
rect 150256 71946 150308 71952
rect 150164 71732 150216 71738
rect 150164 71674 150216 71680
rect 150164 71528 150216 71534
rect 150164 71470 150216 71476
rect 150072 70780 150124 70786
rect 150072 70722 150124 70728
rect 150084 46306 150112 70722
rect 150176 47666 150204 71470
rect 150268 51814 150296 71946
rect 150452 71602 150480 79342
rect 150530 79248 150586 79257
rect 150530 79183 150586 79192
rect 150440 71596 150492 71602
rect 150440 71538 150492 71544
rect 150452 70854 150480 71538
rect 150440 70848 150492 70854
rect 150440 70790 150492 70796
rect 150544 60734 150572 79183
rect 150636 78606 150664 79716
rect 150624 78600 150676 78606
rect 150624 78542 150676 78548
rect 150728 71738 150756 79766
rect 150820 77353 150848 79784
rect 150946 79766 150998 79772
rect 151130 79824 151182 79830
rect 151130 79766 151182 79772
rect 151360 79756 151412 79762
rect 151510 79744 151538 80036
rect 151602 79812 151630 80036
rect 151694 79937 151722 80036
rect 151680 79928 151736 79937
rect 151680 79863 151736 79872
rect 151602 79784 151676 79812
rect 151510 79716 151584 79744
rect 151360 79698 151412 79704
rect 151084 79688 151136 79694
rect 150990 79656 151046 79665
rect 150900 79620 150952 79626
rect 151084 79630 151136 79636
rect 150990 79591 151046 79600
rect 150900 79562 150952 79568
rect 150912 79218 150940 79562
rect 150900 79212 150952 79218
rect 150900 79154 150952 79160
rect 150912 79121 150940 79154
rect 150898 79112 150954 79121
rect 150898 79047 150954 79056
rect 150806 77344 150862 77353
rect 150806 77279 150862 77288
rect 150806 73128 150862 73137
rect 150806 73063 150862 73072
rect 150716 71732 150768 71738
rect 150716 71674 150768 71680
rect 150820 62966 150848 73063
rect 151004 72826 151032 79591
rect 151096 79257 151124 79630
rect 151176 79620 151228 79626
rect 151176 79562 151228 79568
rect 151082 79248 151138 79257
rect 151082 79183 151138 79192
rect 151188 78674 151216 79562
rect 151188 78646 151308 78674
rect 151176 78600 151228 78606
rect 151176 78542 151228 78548
rect 151084 73092 151136 73098
rect 151084 73034 151136 73040
rect 150992 72820 151044 72826
rect 150992 72762 151044 72768
rect 151004 72690 151032 72762
rect 150992 72684 151044 72690
rect 150992 72626 151044 72632
rect 150808 62960 150860 62966
rect 150808 62902 150860 62908
rect 150452 60706 150572 60734
rect 150452 54602 150480 60706
rect 150440 54596 150492 54602
rect 150440 54538 150492 54544
rect 150256 51808 150308 51814
rect 150256 51750 150308 51756
rect 150164 47660 150216 47666
rect 150164 47602 150216 47608
rect 150072 46300 150124 46306
rect 150072 46242 150124 46248
rect 149980 31340 150032 31346
rect 149980 31282 150032 31288
rect 149888 9240 149940 9246
rect 149888 9182 149940 9188
rect 151096 5030 151124 73034
rect 151188 10606 151216 78542
rect 151280 73166 151308 78646
rect 151268 73160 151320 73166
rect 151268 73102 151320 73108
rect 151176 10600 151228 10606
rect 151176 10542 151228 10548
rect 151280 7886 151308 73102
rect 151372 70174 151400 79698
rect 151452 79620 151504 79626
rect 151452 79562 151504 79568
rect 151464 73098 151492 79562
rect 151556 73137 151584 79716
rect 151648 76537 151676 79784
rect 151786 79676 151814 80036
rect 151878 79744 151906 80036
rect 151970 79898 151998 80036
rect 152062 79903 152090 80036
rect 151958 79892 152010 79898
rect 151958 79834 152010 79840
rect 152048 79894 152104 79903
rect 152048 79829 152104 79838
rect 152154 79744 152182 80036
rect 152246 79898 152274 80036
rect 152338 79966 152366 80036
rect 152430 79966 152458 80036
rect 152326 79960 152378 79966
rect 152326 79902 152378 79908
rect 152418 79960 152470 79966
rect 152418 79902 152470 79908
rect 152234 79892 152286 79898
rect 152234 79834 152286 79840
rect 152372 79824 152424 79830
rect 152522 79812 152550 80036
rect 152372 79766 152424 79772
rect 152476 79784 152550 79812
rect 152280 79756 152332 79762
rect 151878 79716 152044 79744
rect 152154 79716 152228 79744
rect 151786 79648 151952 79676
rect 151728 79552 151780 79558
rect 151728 79494 151780 79500
rect 151740 78713 151768 79494
rect 151820 79484 151872 79490
rect 151820 79426 151872 79432
rect 151726 78704 151782 78713
rect 151726 78639 151782 78648
rect 151728 77240 151780 77246
rect 151728 77182 151780 77188
rect 151634 76528 151690 76537
rect 151634 76463 151690 76472
rect 151740 74050 151768 77182
rect 151832 75256 151860 79426
rect 151924 77246 151952 79648
rect 151912 77240 151964 77246
rect 151912 77182 151964 77188
rect 151832 75228 151952 75256
rect 151820 75132 151872 75138
rect 151820 75074 151872 75080
rect 151728 74044 151780 74050
rect 151728 73986 151780 73992
rect 151542 73128 151598 73137
rect 151452 73092 151504 73098
rect 151542 73063 151598 73072
rect 151452 73034 151504 73040
rect 151636 72684 151688 72690
rect 151636 72626 151688 72632
rect 151452 71732 151504 71738
rect 151452 71674 151504 71680
rect 151464 70990 151492 71674
rect 151544 71596 151596 71602
rect 151544 71538 151596 71544
rect 151452 70984 151504 70990
rect 151452 70926 151504 70932
rect 151360 70168 151412 70174
rect 151360 70110 151412 70116
rect 151372 32638 151400 70110
rect 151464 34134 151492 70926
rect 151556 41070 151584 71538
rect 151648 44946 151676 72626
rect 151740 58750 151768 73986
rect 151832 70106 151860 75074
rect 151924 74497 151952 75228
rect 151910 74488 151966 74497
rect 151910 74423 151966 74432
rect 152016 71398 152044 79716
rect 152096 79280 152148 79286
rect 152096 79222 152148 79228
rect 152108 75290 152136 79222
rect 152200 78538 152228 79716
rect 152280 79698 152332 79704
rect 152188 78532 152240 78538
rect 152188 78474 152240 78480
rect 152108 75262 152228 75290
rect 152096 75200 152148 75206
rect 152096 75142 152148 75148
rect 152004 71392 152056 71398
rect 152004 71334 152056 71340
rect 152016 70922 152044 71334
rect 152004 70916 152056 70922
rect 152004 70858 152056 70864
rect 151820 70100 151872 70106
rect 151820 70042 151872 70048
rect 151832 69086 151860 70042
rect 152108 69873 152136 75142
rect 152200 73982 152228 75262
rect 152292 74526 152320 79698
rect 152384 77294 152412 79766
rect 152476 78656 152504 79784
rect 152614 79744 152642 80036
rect 152706 79778 152734 80036
rect 152798 79937 152826 80036
rect 152784 79928 152840 79937
rect 152784 79863 152840 79872
rect 152706 79750 152780 79778
rect 152568 79716 152642 79744
rect 152568 79257 152596 79716
rect 152752 79665 152780 79750
rect 152890 79744 152918 80036
rect 152982 79898 153010 80036
rect 152970 79892 153022 79898
rect 152970 79834 153022 79840
rect 153074 79812 153102 80036
rect 153166 79966 153194 80036
rect 153154 79960 153206 79966
rect 153154 79902 153206 79908
rect 153258 79812 153286 80036
rect 153074 79784 153148 79812
rect 152890 79716 153056 79744
rect 152738 79656 152794 79665
rect 152738 79591 152794 79600
rect 152924 79620 152976 79626
rect 152924 79562 152976 79568
rect 152832 79552 152884 79558
rect 152738 79520 152794 79529
rect 152832 79494 152884 79500
rect 152738 79455 152794 79464
rect 152554 79248 152610 79257
rect 152554 79183 152610 79192
rect 152476 78628 152596 78656
rect 152384 77266 152504 77294
rect 152476 75138 152504 77266
rect 152464 75132 152516 75138
rect 152464 75074 152516 75080
rect 152280 74520 152332 74526
rect 152280 74462 152332 74468
rect 152188 73976 152240 73982
rect 152188 73918 152240 73924
rect 152200 70394 152228 73918
rect 152464 73772 152516 73778
rect 152464 73714 152516 73720
rect 152200 70366 152412 70394
rect 152094 69864 152150 69873
rect 152094 69799 152150 69808
rect 151820 69080 151872 69086
rect 151820 69022 151872 69028
rect 152108 60734 152136 69799
rect 152108 60706 152320 60734
rect 151728 58744 151780 58750
rect 151728 58686 151780 58692
rect 151636 44940 151688 44946
rect 151636 44882 151688 44888
rect 151544 41064 151596 41070
rect 151544 41006 151596 41012
rect 151452 34128 151504 34134
rect 151452 34070 151504 34076
rect 151360 32632 151412 32638
rect 151360 32574 151412 32580
rect 152292 31278 152320 60706
rect 152384 57322 152412 70366
rect 152372 57316 152424 57322
rect 152372 57258 152424 57264
rect 152280 31272 152332 31278
rect 152280 31214 152332 31220
rect 151268 7880 151320 7886
rect 151268 7822 151320 7828
rect 151084 5024 151136 5030
rect 151084 4966 151136 4972
rect 148508 4004 148560 4010
rect 148508 3946 148560 3952
rect 149704 4004 149756 4010
rect 149704 3946 149756 3952
rect 148416 3868 148468 3874
rect 148416 3810 148468 3816
rect 148520 3534 148548 3946
rect 149612 3936 149664 3942
rect 149612 3878 149664 3884
rect 149624 3738 149652 3878
rect 152476 3806 152504 73714
rect 152568 70394 152596 78628
rect 152568 70366 152688 70394
rect 152556 69080 152608 69086
rect 152556 69022 152608 69028
rect 152568 13394 152596 69022
rect 152660 65929 152688 70366
rect 152752 68134 152780 79455
rect 152740 68128 152792 68134
rect 152740 68070 152792 68076
rect 152844 66065 152872 79494
rect 152936 75206 152964 79562
rect 153028 79286 153056 79716
rect 153016 79280 153068 79286
rect 153016 79222 153068 79228
rect 153016 78260 153068 78266
rect 153016 78202 153068 78208
rect 153028 75410 153056 78202
rect 153016 75404 153068 75410
rect 153016 75346 153068 75352
rect 152924 75200 152976 75206
rect 152924 75142 152976 75148
rect 153014 74488 153070 74497
rect 153014 74423 153070 74432
rect 152924 70916 152976 70922
rect 152924 70858 152976 70864
rect 152830 66056 152886 66065
rect 152830 65991 152886 66000
rect 152646 65920 152702 65929
rect 152646 65855 152702 65864
rect 152660 17474 152688 65855
rect 152844 18902 152872 65991
rect 152936 34066 152964 70858
rect 153028 53174 153056 74423
rect 153120 73030 153148 79784
rect 153212 79784 153286 79812
rect 153212 78742 153240 79784
rect 153350 79778 153378 80036
rect 153442 79966 153470 80036
rect 153534 79966 153562 80036
rect 153626 79971 153654 80036
rect 153430 79960 153482 79966
rect 153430 79902 153482 79908
rect 153522 79960 153574 79966
rect 153522 79902 153574 79908
rect 153612 79962 153668 79971
rect 153718 79966 153746 80036
rect 153810 79971 153838 80036
rect 153612 79897 153668 79906
rect 153706 79960 153758 79966
rect 153706 79902 153758 79908
rect 153796 79962 153852 79971
rect 153902 79966 153930 80036
rect 153994 79971 154022 80036
rect 153796 79897 153852 79906
rect 153890 79960 153942 79966
rect 153890 79902 153942 79908
rect 153980 79962 154036 79971
rect 153980 79897 154036 79906
rect 154086 79898 154114 80036
rect 154178 79937 154206 80036
rect 154164 79928 154220 79937
rect 154074 79892 154126 79898
rect 154164 79863 154220 79872
rect 154074 79834 154126 79840
rect 153476 79824 153528 79830
rect 153350 79750 153424 79778
rect 153476 79766 153528 79772
rect 153844 79824 153896 79830
rect 154270 79812 154298 80036
rect 154224 79801 154298 79812
rect 153844 79766 153896 79772
rect 153934 79792 153990 79801
rect 153290 79656 153346 79665
rect 153290 79591 153346 79600
rect 153200 78736 153252 78742
rect 153200 78678 153252 78684
rect 153200 77308 153252 77314
rect 153200 77250 153252 77256
rect 153108 73024 153160 73030
rect 153108 72966 153160 72972
rect 153016 53168 153068 53174
rect 153016 53110 153068 53116
rect 153120 39574 153148 72966
rect 153212 62014 153240 77250
rect 153304 68678 153332 79591
rect 153396 74322 153424 79750
rect 153488 78674 153516 79766
rect 153660 79756 153712 79762
rect 153660 79698 153712 79704
rect 153566 79520 153622 79529
rect 153566 79455 153622 79464
rect 153476 78668 153528 78674
rect 153476 78610 153528 78616
rect 153476 78532 153528 78538
rect 153476 78474 153528 78480
rect 153488 76770 153516 78474
rect 153476 76764 153528 76770
rect 153476 76706 153528 76712
rect 153384 74316 153436 74322
rect 153384 74258 153436 74264
rect 153580 69630 153608 79455
rect 153672 78849 153700 79698
rect 153752 79552 153804 79558
rect 153752 79494 153804 79500
rect 153658 78840 153714 78849
rect 153658 78775 153714 78784
rect 153660 78668 153712 78674
rect 153660 78610 153712 78616
rect 153672 74254 153700 78610
rect 153660 74248 153712 74254
rect 153660 74190 153712 74196
rect 153764 73166 153792 79494
rect 153856 77489 153884 79766
rect 154210 79792 154298 79801
rect 153934 79727 153990 79736
rect 154120 79756 154172 79762
rect 153948 78826 153976 79727
rect 154266 79784 154298 79792
rect 154210 79727 154266 79736
rect 154362 79744 154390 80036
rect 154454 79966 154482 80036
rect 154442 79960 154494 79966
rect 154442 79902 154494 79908
rect 154546 79812 154574 80036
rect 154500 79784 154574 79812
rect 154362 79716 154436 79744
rect 154120 79698 154172 79704
rect 153948 78798 154068 78826
rect 153936 78736 153988 78742
rect 153936 78678 153988 78684
rect 153842 77480 153898 77489
rect 153842 77415 153898 77424
rect 153752 73160 153804 73166
rect 153752 73102 153804 73108
rect 153948 70394 153976 78678
rect 154040 77314 154068 78798
rect 154028 77308 154080 77314
rect 154028 77250 154080 77256
rect 154028 75200 154080 75206
rect 154028 75142 154080 75148
rect 153672 70366 153976 70394
rect 153672 69737 153700 70366
rect 154040 70009 154068 75142
rect 154132 70145 154160 79698
rect 154408 75206 154436 79716
rect 154500 77353 154528 79784
rect 154638 79744 154666 80036
rect 154592 79716 154666 79744
rect 154592 77466 154620 79716
rect 154730 79642 154758 80036
rect 154822 79966 154850 80036
rect 154914 79971 154942 80036
rect 154810 79960 154862 79966
rect 154810 79902 154862 79908
rect 154900 79962 154956 79971
rect 155006 79966 155034 80036
rect 154900 79897 154956 79906
rect 154994 79960 155046 79966
rect 154994 79902 155046 79908
rect 155098 79778 155126 80036
rect 154856 79756 154908 79762
rect 154856 79698 154908 79704
rect 154960 79750 155126 79778
rect 154684 79614 154758 79642
rect 154684 77586 154712 79614
rect 154868 79529 154896 79698
rect 154854 79520 154910 79529
rect 154854 79455 154910 79464
rect 154868 78985 154896 79455
rect 154854 78976 154910 78985
rect 154854 78911 154910 78920
rect 154960 77874 154988 79750
rect 155040 79688 155092 79694
rect 155190 79642 155218 80036
rect 155282 79971 155310 80036
rect 155268 79962 155324 79971
rect 155374 79966 155402 80036
rect 155268 79897 155324 79906
rect 155362 79960 155414 79966
rect 155362 79902 155414 79908
rect 155316 79824 155368 79830
rect 155316 79766 155368 79772
rect 155040 79630 155092 79636
rect 154776 77846 154988 77874
rect 154672 77580 154724 77586
rect 154672 77522 154724 77528
rect 154592 77438 154712 77466
rect 154486 77344 154542 77353
rect 154486 77279 154542 77288
rect 154684 77042 154712 77438
rect 154672 77036 154724 77042
rect 154672 76978 154724 76984
rect 154670 76936 154726 76945
rect 154670 76871 154726 76880
rect 154580 76424 154632 76430
rect 154580 76366 154632 76372
rect 154396 75200 154448 75206
rect 154396 75142 154448 75148
rect 154212 74248 154264 74254
rect 154212 74190 154264 74196
rect 154118 70136 154174 70145
rect 154118 70071 154174 70080
rect 154026 70000 154082 70009
rect 154026 69935 154082 69944
rect 153658 69728 153714 69737
rect 153658 69663 153714 69672
rect 153568 69624 153620 69630
rect 153568 69566 153620 69572
rect 153292 68672 153344 68678
rect 153292 68614 153344 68620
rect 153200 62008 153252 62014
rect 153200 61950 153252 61956
rect 153108 39568 153160 39574
rect 153108 39510 153160 39516
rect 153672 36786 153700 69663
rect 154040 66994 154068 69935
rect 153948 66966 154068 66994
rect 153948 60734 153976 66966
rect 154132 60734 154160 70071
rect 153856 60706 153976 60734
rect 154040 60706 154160 60734
rect 153660 36780 153712 36786
rect 153660 36722 153712 36728
rect 152924 34060 152976 34066
rect 152924 34002 152976 34008
rect 153856 23050 153884 60706
rect 154040 25770 154068 60706
rect 154224 27198 154252 74190
rect 154396 73160 154448 73166
rect 154396 73102 154448 73108
rect 154408 72758 154436 73102
rect 154396 72752 154448 72758
rect 154396 72694 154448 72700
rect 154304 68672 154356 68678
rect 154304 68614 154356 68620
rect 154316 68066 154344 68614
rect 154304 68060 154356 68066
rect 154304 68002 154356 68008
rect 154212 27192 154264 27198
rect 154212 27134 154264 27140
rect 154028 25764 154080 25770
rect 154028 25706 154080 25712
rect 153844 23044 153896 23050
rect 153844 22986 153896 22992
rect 152832 18896 152884 18902
rect 152832 18838 152884 18844
rect 152648 17468 152700 17474
rect 152648 17410 152700 17416
rect 154316 14754 154344 68002
rect 154408 16182 154436 72694
rect 154488 69828 154540 69834
rect 154488 69770 154540 69776
rect 154500 69630 154528 69770
rect 154488 69624 154540 69630
rect 154488 69566 154540 69572
rect 154396 16176 154448 16182
rect 154396 16118 154448 16124
rect 154304 14748 154356 14754
rect 154304 14690 154356 14696
rect 152556 13388 152608 13394
rect 152556 13330 152608 13336
rect 154500 6798 154528 69566
rect 154592 41410 154620 76366
rect 154684 60586 154712 76871
rect 154776 63442 154804 77846
rect 155052 77704 155080 79630
rect 154960 77676 155080 77704
rect 155144 79614 155218 79642
rect 154856 77172 154908 77178
rect 154856 77114 154908 77120
rect 154868 66094 154896 77114
rect 154960 67561 154988 77676
rect 155040 77580 155092 77586
rect 155040 77522 155092 77528
rect 154946 67552 155002 67561
rect 154946 67487 155002 67496
rect 155052 67386 155080 77522
rect 155144 76430 155172 79614
rect 155328 79370 155356 79766
rect 155466 79744 155494 80036
rect 155558 79966 155586 80036
rect 155546 79960 155598 79966
rect 155650 79937 155678 80036
rect 155546 79902 155598 79908
rect 155636 79928 155692 79937
rect 155742 79898 155770 80036
rect 155834 79898 155862 80036
rect 155926 79966 155954 80036
rect 155914 79960 155966 79966
rect 155914 79902 155966 79908
rect 155636 79863 155692 79872
rect 155730 79892 155782 79898
rect 155730 79834 155782 79840
rect 155822 79892 155874 79898
rect 155822 79834 155874 79840
rect 155592 79824 155644 79830
rect 156018 79778 156046 80036
rect 156110 79903 156138 80036
rect 156202 79966 156230 80036
rect 156294 79966 156322 80036
rect 156190 79960 156242 79966
rect 156096 79894 156152 79903
rect 156190 79902 156242 79908
rect 156282 79960 156334 79966
rect 156282 79902 156334 79908
rect 156096 79829 156152 79838
rect 155592 79766 155644 79772
rect 155466 79716 155540 79744
rect 155408 79620 155460 79626
rect 155408 79562 155460 79568
rect 155236 79342 155356 79370
rect 155236 77178 155264 79342
rect 155224 77172 155276 77178
rect 155224 77114 155276 77120
rect 155132 76424 155184 76430
rect 155132 76366 155184 76372
rect 155420 74534 155448 79562
rect 155512 77178 155540 79716
rect 155500 77172 155552 77178
rect 155500 77114 155552 77120
rect 155500 77036 155552 77042
rect 155500 76978 155552 76984
rect 155328 74506 155448 74534
rect 155328 70394 155356 74506
rect 155512 74361 155540 76978
rect 155604 74534 155632 79766
rect 155972 79750 156046 79778
rect 156282 79824 156334 79830
rect 156282 79766 156334 79772
rect 156144 79756 156196 79762
rect 155868 79620 155920 79626
rect 155868 79562 155920 79568
rect 155880 77353 155908 79562
rect 155866 77344 155922 77353
rect 155866 77279 155922 77288
rect 155604 74506 155724 74534
rect 155498 74352 155554 74361
rect 155498 74287 155554 74296
rect 155236 70366 155356 70394
rect 155236 68785 155264 70366
rect 155222 68776 155278 68785
rect 155222 68711 155278 68720
rect 155040 67380 155092 67386
rect 155040 67322 155092 67328
rect 154856 66088 154908 66094
rect 154856 66030 154908 66036
rect 154764 63436 154816 63442
rect 154764 63378 154816 63384
rect 154672 60580 154724 60586
rect 154672 60522 154724 60528
rect 154580 41404 154632 41410
rect 154580 41346 154632 41352
rect 155236 29918 155264 68711
rect 155512 60734 155540 74287
rect 155696 73166 155724 74506
rect 155684 73160 155736 73166
rect 155684 73102 155736 73108
rect 155774 67552 155830 67561
rect 155774 67487 155830 67496
rect 155328 60706 155540 60734
rect 155328 46238 155356 60706
rect 155316 46232 155368 46238
rect 155316 46174 155368 46180
rect 155224 29912 155276 29918
rect 155224 29854 155276 29860
rect 155788 20058 155816 67487
rect 155868 67380 155920 67386
rect 155868 67322 155920 67328
rect 155880 20126 155908 67322
rect 155972 66230 156000 79750
rect 156144 79698 156196 79704
rect 156050 79656 156106 79665
rect 156050 79591 156106 79600
rect 156064 76226 156092 79591
rect 156052 76220 156104 76226
rect 156052 76162 156104 76168
rect 156052 75132 156104 75138
rect 156052 75074 156104 75080
rect 156064 68882 156092 75074
rect 156052 68876 156104 68882
rect 156052 68818 156104 68824
rect 156064 67658 156092 68818
rect 156052 67652 156104 67658
rect 156052 67594 156104 67600
rect 155960 66224 156012 66230
rect 155960 66166 156012 66172
rect 155972 65822 156000 66166
rect 155960 65816 156012 65822
rect 155960 65758 156012 65764
rect 156156 64802 156184 79698
rect 156294 79676 156322 79766
rect 156386 79744 156414 80036
rect 156478 79971 156506 80036
rect 156464 79962 156520 79971
rect 156464 79897 156520 79906
rect 156570 79744 156598 80036
rect 156662 79898 156690 80036
rect 156650 79892 156702 79898
rect 156650 79834 156702 79840
rect 156754 79778 156782 80036
rect 156846 79898 156874 80036
rect 156938 79966 156966 80036
rect 156926 79960 156978 79966
rect 156926 79902 156978 79908
rect 156834 79892 156886 79898
rect 156834 79834 156886 79840
rect 157030 79778 157058 80036
rect 157122 79966 157150 80036
rect 157110 79960 157162 79966
rect 157110 79902 157162 79908
rect 157214 79812 157242 80036
rect 157306 79937 157334 80036
rect 157398 79966 157426 80036
rect 157386 79960 157438 79966
rect 157292 79928 157348 79937
rect 157386 79902 157438 79908
rect 157292 79863 157348 79872
rect 157490 79830 157518 80036
rect 157582 79971 157610 80036
rect 157568 79962 157624 79971
rect 157568 79897 157624 79906
rect 157674 79898 157702 80036
rect 157766 79966 157794 80036
rect 157858 79966 157886 80036
rect 157950 79966 157978 80036
rect 158042 79971 158070 80036
rect 157754 79960 157806 79966
rect 157754 79902 157806 79908
rect 157846 79960 157898 79966
rect 157846 79902 157898 79908
rect 157938 79960 157990 79966
rect 157938 79902 157990 79908
rect 158028 79962 158084 79971
rect 157662 79892 157714 79898
rect 158028 79897 158084 79906
rect 157662 79834 157714 79840
rect 157478 79824 157530 79830
rect 157214 79784 157288 79812
rect 156754 79762 156828 79778
rect 156754 79756 156840 79762
rect 156754 79750 156788 79756
rect 156386 79716 156460 79744
rect 156570 79716 156644 79744
rect 156248 79648 156322 79676
rect 156248 70394 156276 79648
rect 156328 79552 156380 79558
rect 156328 79494 156380 79500
rect 156340 70990 156368 79494
rect 156432 78674 156460 79716
rect 156616 79665 156644 79716
rect 156788 79698 156840 79704
rect 156880 79756 156932 79762
rect 157030 79750 157104 79778
rect 156880 79698 156932 79704
rect 156602 79656 156658 79665
rect 156602 79591 156658 79600
rect 156788 79620 156840 79626
rect 156788 79562 156840 79568
rect 156696 79552 156748 79558
rect 156696 79494 156748 79500
rect 156432 78646 156552 78674
rect 156524 78577 156552 78646
rect 156510 78568 156566 78577
rect 156510 78503 156566 78512
rect 156708 77314 156736 79494
rect 156696 77308 156748 77314
rect 156696 77250 156748 77256
rect 156800 72622 156828 79562
rect 156788 72616 156840 72622
rect 156788 72558 156840 72564
rect 156328 70984 156380 70990
rect 156328 70926 156380 70932
rect 156248 70366 156736 70394
rect 156602 67688 156658 67697
rect 156602 67623 156658 67632
rect 156144 64796 156196 64802
rect 156144 64738 156196 64744
rect 155958 37904 156014 37913
rect 155958 37839 156014 37848
rect 155868 20120 155920 20126
rect 155868 20062 155920 20068
rect 155776 20052 155828 20058
rect 155776 19994 155828 20000
rect 154580 19984 154632 19990
rect 154580 19926 154632 19932
rect 154592 16574 154620 19926
rect 155972 16574 156000 37839
rect 154592 16546 155448 16574
rect 155972 16546 156184 16574
rect 154488 6792 154540 6798
rect 154488 6734 154540 6740
rect 154212 4140 154264 4146
rect 154212 4082 154264 4088
rect 153016 4004 153068 4010
rect 153016 3946 153068 3952
rect 151820 3800 151872 3806
rect 151820 3742 151872 3748
rect 152464 3800 152516 3806
rect 152464 3742 152516 3748
rect 149520 3732 149572 3738
rect 149520 3674 149572 3680
rect 149612 3732 149664 3738
rect 149612 3674 149664 3680
rect 147220 3528 147272 3534
rect 146864 3454 147168 3482
rect 147220 3470 147272 3476
rect 148324 3528 148376 3534
rect 148324 3470 148376 3476
rect 148508 3528 148560 3534
rect 148508 3470 148560 3476
rect 147140 480 147168 3454
rect 148336 480 148364 3470
rect 149532 480 149560 3674
rect 150624 3392 150676 3398
rect 150624 3334 150676 3340
rect 150636 480 150664 3334
rect 151832 480 151860 3742
rect 153028 480 153056 3946
rect 154224 480 154252 4082
rect 155420 480 155448 16546
rect 145902 354 146014 480
rect 145484 326 146014 354
rect 145902 -960 146014 326
rect 147098 -960 147210 480
rect 148294 -960 148406 480
rect 149490 -960 149602 480
rect 150594 -960 150706 480
rect 151790 -960 151902 480
rect 152986 -960 153098 480
rect 154182 -960 154294 480
rect 155378 -960 155490 480
rect 156156 354 156184 16546
rect 156616 9178 156644 67623
rect 156708 66201 156736 70366
rect 156892 68649 156920 79698
rect 156972 79688 157024 79694
rect 156972 79630 157024 79636
rect 156984 79218 157012 79630
rect 156972 79212 157024 79218
rect 156972 79154 157024 79160
rect 157076 78674 157104 79750
rect 157156 79688 157208 79694
rect 157156 79630 157208 79636
rect 156984 78646 157104 78674
rect 156878 68640 156934 68649
rect 156878 68575 156934 68584
rect 156892 67697 156920 68575
rect 156878 67688 156934 67697
rect 156788 67652 156840 67658
rect 156878 67623 156934 67632
rect 156788 67594 156840 67600
rect 156800 67538 156828 67594
rect 156800 67510 156920 67538
rect 156694 66192 156750 66201
rect 156694 66127 156750 66136
rect 156708 13326 156736 66127
rect 156788 65816 156840 65822
rect 156788 65758 156840 65764
rect 156800 35426 156828 65758
rect 156892 38146 156920 67510
rect 156984 55214 157012 78646
rect 157168 78470 157196 79630
rect 157156 78464 157208 78470
rect 157156 78406 157208 78412
rect 157156 77308 157208 77314
rect 157156 77250 157208 77256
rect 157064 75540 157116 75546
rect 157064 75482 157116 75488
rect 157076 75342 157104 75482
rect 157064 75336 157116 75342
rect 157064 75278 157116 75284
rect 157168 72962 157196 77250
rect 157260 75138 157288 79784
rect 157478 79766 157530 79772
rect 158134 79778 158162 80036
rect 158226 79966 158254 80036
rect 158318 79971 158346 80036
rect 158214 79960 158266 79966
rect 158214 79902 158266 79908
rect 158304 79962 158360 79971
rect 158410 79966 158438 80036
rect 158502 79966 158530 80036
rect 158594 79971 158622 80036
rect 158304 79897 158360 79906
rect 158398 79960 158450 79966
rect 158398 79902 158450 79908
rect 158490 79960 158542 79966
rect 158490 79902 158542 79908
rect 158580 79962 158636 79971
rect 158580 79897 158636 79906
rect 158444 79824 158496 79830
rect 157340 79756 157392 79762
rect 157340 79698 157392 79704
rect 157708 79756 157760 79762
rect 158134 79750 158208 79778
rect 158686 79812 158714 80036
rect 158778 79966 158806 80036
rect 158766 79960 158818 79966
rect 158766 79902 158818 79908
rect 158870 79898 158898 80036
rect 158962 79966 158990 80036
rect 158950 79960 159002 79966
rect 158950 79902 159002 79908
rect 158858 79892 158910 79898
rect 158858 79834 158910 79840
rect 158686 79784 158760 79812
rect 158444 79766 158496 79772
rect 157708 79698 157760 79704
rect 157352 75478 157380 79698
rect 157524 79620 157576 79626
rect 157524 79562 157576 79568
rect 157616 79620 157668 79626
rect 157616 79562 157668 79568
rect 157432 78668 157484 78674
rect 157432 78610 157484 78616
rect 157340 75472 157392 75478
rect 157340 75414 157392 75420
rect 157444 75290 157472 78610
rect 157352 75262 157472 75290
rect 157248 75132 157300 75138
rect 157248 75074 157300 75080
rect 157156 72956 157208 72962
rect 157156 72898 157208 72904
rect 157064 72616 157116 72622
rect 157064 72558 157116 72564
rect 157076 61946 157104 72558
rect 157352 71670 157380 75262
rect 157432 75132 157484 75138
rect 157432 75074 157484 75080
rect 157340 71664 157392 71670
rect 157340 71606 157392 71612
rect 157340 71528 157392 71534
rect 157340 71470 157392 71476
rect 157248 70984 157300 70990
rect 157248 70926 157300 70932
rect 157064 61940 157116 61946
rect 157064 61882 157116 61888
rect 156972 55208 157024 55214
rect 156972 55150 157024 55156
rect 156880 38140 156932 38146
rect 156880 38082 156932 38088
rect 156788 35420 156840 35426
rect 156788 35362 156840 35368
rect 157260 14686 157288 70926
rect 157352 40934 157380 71470
rect 157444 56574 157472 75074
rect 157536 72690 157564 79562
rect 157628 78674 157656 79562
rect 157616 78668 157668 78674
rect 157616 78610 157668 78616
rect 157616 75472 157668 75478
rect 157616 75414 157668 75420
rect 157524 72684 157576 72690
rect 157524 72626 157576 72632
rect 157628 71602 157656 75414
rect 157720 72622 157748 79698
rect 157800 79620 157852 79626
rect 157800 79562 157852 79568
rect 157984 79620 158036 79626
rect 157984 79562 158036 79568
rect 157708 72616 157760 72622
rect 157708 72558 157760 72564
rect 157616 71596 157668 71602
rect 157616 71538 157668 71544
rect 157812 70394 157840 79562
rect 157892 79212 157944 79218
rect 157892 79154 157944 79160
rect 157904 71534 157932 79154
rect 157996 71738 158024 79562
rect 158074 78160 158130 78169
rect 158074 78095 158130 78104
rect 158088 77110 158116 78095
rect 158076 77104 158128 77110
rect 158076 77046 158128 77052
rect 158180 75138 158208 79750
rect 158260 79756 158312 79762
rect 158260 79698 158312 79704
rect 158168 75132 158220 75138
rect 158168 75074 158220 75080
rect 158272 73930 158300 79698
rect 158352 79688 158404 79694
rect 158352 79630 158404 79636
rect 158364 79218 158392 79630
rect 158352 79212 158404 79218
rect 158352 79154 158404 79160
rect 158272 73902 158392 73930
rect 157984 71732 158036 71738
rect 157984 71674 158036 71680
rect 158260 71664 158312 71670
rect 158260 71606 158312 71612
rect 157892 71528 157944 71534
rect 157892 71470 157944 71476
rect 158272 71262 158300 71606
rect 158364 71534 158392 73902
rect 158456 73794 158484 79766
rect 158732 79744 158760 79784
rect 158904 79756 158956 79762
rect 158732 79716 158852 79744
rect 158626 79656 158682 79665
rect 158626 79591 158682 79600
rect 158640 79286 158668 79591
rect 158720 79484 158772 79490
rect 158720 79426 158772 79432
rect 158628 79280 158680 79286
rect 158628 79222 158680 79228
rect 158456 73766 158668 73794
rect 158536 71732 158588 71738
rect 158536 71674 158588 71680
rect 158444 71596 158496 71602
rect 158444 71538 158496 71544
rect 158352 71528 158404 71534
rect 158352 71470 158404 71476
rect 158260 71256 158312 71262
rect 158260 71198 158312 71204
rect 157536 70366 157840 70394
rect 157536 59362 157564 70366
rect 157524 59356 157576 59362
rect 157524 59298 157576 59304
rect 157432 56568 157484 56574
rect 157432 56510 157484 56516
rect 158272 42294 158300 71198
rect 158260 42288 158312 42294
rect 158260 42230 158312 42236
rect 157340 40928 157392 40934
rect 157340 40870 157392 40876
rect 158364 32570 158392 71470
rect 158456 71398 158484 71538
rect 158444 71392 158496 71398
rect 158444 71334 158496 71340
rect 158352 32564 158404 32570
rect 158352 32506 158404 32512
rect 158456 28490 158484 71334
rect 158548 70922 158576 71674
rect 158536 70916 158588 70922
rect 158536 70858 158588 70864
rect 158444 28484 158496 28490
rect 158444 28426 158496 28432
rect 157982 28248 158038 28257
rect 157982 28183 158038 28192
rect 157248 14680 157300 14686
rect 157248 14622 157300 14628
rect 156696 13320 156748 13326
rect 156696 13262 156748 13268
rect 157798 10296 157854 10305
rect 157798 10231 157854 10240
rect 156604 9172 156656 9178
rect 156604 9114 156656 9120
rect 157812 480 157840 10231
rect 157996 3398 158024 28183
rect 158548 11966 158576 70858
rect 158640 70854 158668 73766
rect 158628 70848 158680 70854
rect 158628 70790 158680 70796
rect 158536 11960 158588 11966
rect 158536 11902 158588 11908
rect 158640 10538 158668 70790
rect 158732 60722 158760 79426
rect 158824 78985 158852 79716
rect 158904 79698 158956 79704
rect 158810 78976 158866 78985
rect 158810 78911 158866 78920
rect 158812 78668 158864 78674
rect 158812 78610 158864 78616
rect 158824 75478 158852 78610
rect 158916 78538 158944 79698
rect 159054 79676 159082 80036
rect 159146 79937 159174 80036
rect 159238 79966 159266 80036
rect 159226 79960 159278 79966
rect 159132 79928 159188 79937
rect 159226 79902 159278 79908
rect 159132 79863 159188 79872
rect 159330 79676 159358 80036
rect 159422 79801 159450 80036
rect 159514 79830 159542 80036
rect 159606 79898 159634 80036
rect 159594 79892 159646 79898
rect 159594 79834 159646 79840
rect 159502 79824 159554 79830
rect 159408 79792 159464 79801
rect 159502 79766 159554 79772
rect 159408 79727 159464 79736
rect 159008 79648 159082 79676
rect 159284 79648 159358 79676
rect 159548 79688 159600 79694
rect 159008 79082 159036 79648
rect 159180 79620 159232 79626
rect 159180 79562 159232 79568
rect 158996 79076 159048 79082
rect 158996 79018 159048 79024
rect 159192 78962 159220 79562
rect 158996 78940 159048 78946
rect 158996 78882 159048 78888
rect 159100 78934 159220 78962
rect 158904 78532 158956 78538
rect 158904 78474 158956 78480
rect 158812 75472 158864 75478
rect 159008 75426 159036 78882
rect 159100 78674 159128 78934
rect 159178 78704 159234 78713
rect 159088 78668 159140 78674
rect 159178 78639 159234 78648
rect 159088 78610 159140 78616
rect 159088 75540 159140 75546
rect 159088 75482 159140 75488
rect 158812 75414 158864 75420
rect 158916 75398 159036 75426
rect 158812 75132 158864 75138
rect 158812 75074 158864 75080
rect 158824 65958 158852 75074
rect 158916 69018 158944 75398
rect 159100 75342 159128 75482
rect 159088 75336 159140 75342
rect 159088 75278 159140 75284
rect 159192 72554 159220 78639
rect 159180 72548 159232 72554
rect 159180 72490 159232 72496
rect 159284 72434 159312 79648
rect 159698 79676 159726 80036
rect 159790 79898 159818 80036
rect 159778 79892 159830 79898
rect 159778 79834 159830 79840
rect 159882 79812 159910 80036
rect 159974 79966 160002 80036
rect 160066 79966 160094 80036
rect 160158 79966 160186 80036
rect 159962 79960 160014 79966
rect 159962 79902 160014 79908
rect 160054 79960 160106 79966
rect 160054 79902 160106 79908
rect 160146 79960 160198 79966
rect 160146 79902 160198 79908
rect 160052 79826 160108 79835
rect 159882 79784 159956 79812
rect 159548 79630 159600 79636
rect 159652 79648 159726 79676
rect 159456 79620 159508 79626
rect 159456 79562 159508 79568
rect 159364 79552 159416 79558
rect 159364 79494 159416 79500
rect 159008 72406 159312 72434
rect 159008 69766 159036 72406
rect 159376 71738 159404 79494
rect 159364 71732 159416 71738
rect 159364 71674 159416 71680
rect 159468 70394 159496 79562
rect 159560 78577 159588 79630
rect 159652 78946 159680 79648
rect 159824 79552 159876 79558
rect 159824 79494 159876 79500
rect 159732 79076 159784 79082
rect 159732 79018 159784 79024
rect 159640 78940 159692 78946
rect 159640 78882 159692 78888
rect 159640 78804 159692 78810
rect 159640 78746 159692 78752
rect 159546 78568 159602 78577
rect 159546 78503 159602 78512
rect 159652 76906 159680 78746
rect 159744 77994 159772 79018
rect 159732 77988 159784 77994
rect 159732 77930 159784 77936
rect 159640 76900 159692 76906
rect 159640 76842 159692 76848
rect 159548 75744 159600 75750
rect 159548 75686 159600 75692
rect 159560 75206 159588 75686
rect 159732 75472 159784 75478
rect 159732 75414 159784 75420
rect 159548 75200 159600 75206
rect 159548 75142 159600 75148
rect 159548 71732 159600 71738
rect 159548 71674 159600 71680
rect 159100 70366 159496 70394
rect 159100 69902 159128 70366
rect 159088 69896 159140 69902
rect 159088 69838 159140 69844
rect 158996 69760 159048 69766
rect 158996 69702 159048 69708
rect 158904 69012 158956 69018
rect 158904 68954 158956 68960
rect 158812 65952 158864 65958
rect 158812 65894 158864 65900
rect 158720 60716 158772 60722
rect 158720 60658 158772 60664
rect 159560 33998 159588 71674
rect 159744 70394 159772 75414
rect 159836 75138 159864 79494
rect 159928 78810 159956 79784
rect 160052 79761 160108 79770
rect 160250 79778 160278 80036
rect 160342 79966 160370 80036
rect 160330 79960 160382 79966
rect 160330 79902 160382 79908
rect 160250 79750 160324 79778
rect 160192 79688 160244 79694
rect 160192 79630 160244 79636
rect 160008 79620 160060 79626
rect 160008 79562 160060 79568
rect 160020 79082 160048 79562
rect 160008 79076 160060 79082
rect 160008 79018 160060 79024
rect 159916 78804 159968 78810
rect 159916 78746 159968 78752
rect 159916 77988 159968 77994
rect 159916 77930 159968 77936
rect 159824 75132 159876 75138
rect 159824 75074 159876 75080
rect 159928 72282 159956 77930
rect 160020 77294 160048 79018
rect 160204 77994 160232 79630
rect 160192 77988 160244 77994
rect 160192 77930 160244 77936
rect 160020 77266 160140 77294
rect 159916 72276 159968 72282
rect 159916 72218 159968 72224
rect 159928 70394 159956 72218
rect 159744 70366 159864 70394
rect 159928 70366 160048 70394
rect 159640 69760 159692 69766
rect 159640 69702 159692 69708
rect 159548 33992 159600 33998
rect 159548 33934 159600 33940
rect 159652 31210 159680 69702
rect 159732 69012 159784 69018
rect 159732 68954 159784 68960
rect 159640 31204 159692 31210
rect 159640 31146 159692 31152
rect 159744 21486 159772 68954
rect 159732 21480 159784 21486
rect 159732 21422 159784 21428
rect 159836 18834 159864 70366
rect 159916 69896 159968 69902
rect 159916 69838 159968 69844
rect 159824 18828 159876 18834
rect 159824 18770 159876 18776
rect 158628 10532 158680 10538
rect 158628 10474 158680 10480
rect 159928 6730 159956 69838
rect 160020 7818 160048 70366
rect 160112 16114 160140 77266
rect 160192 75472 160244 75478
rect 160192 75414 160244 75420
rect 160204 66230 160232 75414
rect 160296 67522 160324 79750
rect 160434 79744 160462 80036
rect 160526 79830 160554 80036
rect 160514 79824 160566 79830
rect 160618 79812 160646 80036
rect 160710 79966 160738 80036
rect 160698 79960 160750 79966
rect 160698 79902 160750 79908
rect 160618 79784 160692 79812
rect 160514 79766 160566 79772
rect 160388 79716 160462 79744
rect 160388 78962 160416 79716
rect 160560 79688 160612 79694
rect 160560 79630 160612 79636
rect 160388 78934 160508 78962
rect 160376 78804 160428 78810
rect 160376 78746 160428 78752
rect 160388 75546 160416 78746
rect 160376 75540 160428 75546
rect 160376 75482 160428 75488
rect 160376 75132 160428 75138
rect 160376 75074 160428 75080
rect 160284 67516 160336 67522
rect 160284 67458 160336 67464
rect 160388 67289 160416 75074
rect 160480 69630 160508 78934
rect 160572 75138 160600 79630
rect 160664 78713 160692 79784
rect 160802 79778 160830 80036
rect 160894 79937 160922 80036
rect 160880 79928 160936 79937
rect 160880 79863 160936 79872
rect 160802 79750 160922 79778
rect 160894 79676 160922 79750
rect 160756 79648 160922 79676
rect 160986 79676 161014 80036
rect 161078 79744 161106 80036
rect 161170 79966 161198 80036
rect 161158 79960 161210 79966
rect 161158 79902 161210 79908
rect 161262 79744 161290 80036
rect 161078 79716 161152 79744
rect 160986 79648 161060 79676
rect 160650 78704 160706 78713
rect 160650 78639 160706 78648
rect 160756 75478 160784 79648
rect 160836 79552 160888 79558
rect 160836 79494 160888 79500
rect 160928 79552 160980 79558
rect 160928 79494 160980 79500
rect 160848 78674 160876 79494
rect 160940 78713 160968 79494
rect 160926 78704 160982 78713
rect 160836 78668 160888 78674
rect 160926 78639 160982 78648
rect 160836 78610 160888 78616
rect 161032 78554 161060 79648
rect 160848 78526 161060 78554
rect 160848 77042 160876 78526
rect 161124 77382 161152 79716
rect 161216 79716 161290 79744
rect 161216 78810 161244 79716
rect 161354 79642 161382 80036
rect 161446 79937 161474 80036
rect 161432 79928 161488 79937
rect 161432 79863 161488 79872
rect 161538 79778 161566 80036
rect 161630 79966 161658 80036
rect 161618 79960 161670 79966
rect 161618 79902 161670 79908
rect 161722 79898 161750 80036
rect 161710 79892 161762 79898
rect 161710 79834 161762 79840
rect 161538 79750 161704 79778
rect 161676 79642 161704 79750
rect 161814 79676 161842 80036
rect 161906 79898 161934 80036
rect 161998 79937 162026 80036
rect 161984 79928 162040 79937
rect 161894 79892 161946 79898
rect 161984 79863 162040 79872
rect 161894 79834 161946 79840
rect 162090 79744 162118 80036
rect 162182 79966 162210 80036
rect 162170 79960 162222 79966
rect 162170 79902 162222 79908
rect 162274 79830 162302 80036
rect 162366 79971 162394 80036
rect 162352 79962 162408 79971
rect 162352 79897 162408 79906
rect 162262 79824 162314 79830
rect 162458 79812 162486 80036
rect 162262 79766 162314 79772
rect 162412 79784 162486 79812
rect 162550 79801 162578 80036
rect 162642 79971 162670 80036
rect 162628 79962 162684 79971
rect 162628 79897 162684 79906
rect 162734 79830 162762 80036
rect 162722 79824 162774 79830
rect 162536 79792 162592 79801
rect 162090 79716 162164 79744
rect 161814 79648 161888 79676
rect 161308 79614 161382 79642
rect 161584 79614 161704 79642
rect 161204 78804 161256 78810
rect 161204 78746 161256 78752
rect 161308 78656 161336 79614
rect 161584 79150 161612 79614
rect 161664 79552 161716 79558
rect 161664 79494 161716 79500
rect 161756 79552 161808 79558
rect 161756 79494 161808 79500
rect 161572 79144 161624 79150
rect 161572 79086 161624 79092
rect 161216 78628 161336 78656
rect 161112 77376 161164 77382
rect 161112 77318 161164 77324
rect 160836 77036 160888 77042
rect 160836 76978 160888 76984
rect 161020 76220 161072 76226
rect 161020 76162 161072 76168
rect 160744 75472 160796 75478
rect 160744 75414 160796 75420
rect 160560 75132 160612 75138
rect 160560 75074 160612 75080
rect 161032 72486 161060 76162
rect 161020 72480 161072 72486
rect 161020 72422 161072 72428
rect 161216 70394 161244 78628
rect 161296 78464 161348 78470
rect 161296 78406 161348 78412
rect 160572 70366 161244 70394
rect 160468 69624 160520 69630
rect 160468 69566 160520 69572
rect 160374 67280 160430 67289
rect 160374 67215 160430 67224
rect 160572 67153 160600 70366
rect 161112 69624 161164 69630
rect 161112 69566 161164 69572
rect 160928 67516 160980 67522
rect 160928 67458 160980 67464
rect 160558 67144 160614 67153
rect 160558 67079 160614 67088
rect 160192 66224 160244 66230
rect 160192 66166 160244 66172
rect 160190 51776 160246 51785
rect 160190 51711 160246 51720
rect 160100 16108 160152 16114
rect 160100 16050 160152 16056
rect 160008 7812 160060 7818
rect 160008 7754 160060 7760
rect 160204 6914 160232 51711
rect 160940 36718 160968 67458
rect 161018 67144 161074 67153
rect 161018 67079 161074 67088
rect 160928 36712 160980 36718
rect 160928 36654 160980 36660
rect 161032 32502 161060 67079
rect 161020 32496 161072 32502
rect 161020 32438 161072 32444
rect 161124 27130 161152 69566
rect 161308 67590 161336 78406
rect 161478 78296 161534 78305
rect 161478 78231 161534 78240
rect 161388 75540 161440 75546
rect 161388 75482 161440 75488
rect 161400 73982 161428 75482
rect 161388 73976 161440 73982
rect 161388 73918 161440 73924
rect 161296 67584 161348 67590
rect 161296 67526 161348 67532
rect 161202 67280 161258 67289
rect 161202 67215 161258 67224
rect 161112 27124 161164 27130
rect 161112 27066 161164 27072
rect 161216 19990 161244 67215
rect 161296 66224 161348 66230
rect 161296 66166 161348 66172
rect 161204 19984 161256 19990
rect 161204 19926 161256 19932
rect 161308 10470 161336 66166
rect 161296 10464 161348 10470
rect 161296 10406 161348 10412
rect 160112 6886 160232 6914
rect 159916 6724 159968 6730
rect 159916 6666 159968 6672
rect 157984 3392 158036 3398
rect 157984 3334 158036 3340
rect 158904 3392 158956 3398
rect 158904 3334 158956 3340
rect 158916 480 158944 3334
rect 160112 480 160140 6886
rect 161296 6180 161348 6186
rect 161296 6122 161348 6128
rect 161308 480 161336 6122
rect 161400 4962 161428 73918
rect 161492 73098 161520 78231
rect 161676 77926 161704 79494
rect 161768 79234 161796 79494
rect 161860 79370 161888 79648
rect 162032 79620 162084 79626
rect 162032 79562 162084 79568
rect 161860 79342 161980 79370
rect 161768 79206 161888 79234
rect 161756 79144 161808 79150
rect 161756 79086 161808 79092
rect 161664 77920 161716 77926
rect 161664 77862 161716 77868
rect 161572 75472 161624 75478
rect 161572 75414 161624 75420
rect 161480 73092 161532 73098
rect 161480 73034 161532 73040
rect 161480 72888 161532 72894
rect 161480 72830 161532 72836
rect 161492 44878 161520 72830
rect 161584 64530 161612 75414
rect 161664 75132 161716 75138
rect 161664 75074 161716 75080
rect 161676 68649 161704 75074
rect 161768 70038 161796 79086
rect 161860 79014 161888 79206
rect 161848 79008 161900 79014
rect 161848 78950 161900 78956
rect 161848 77308 161900 77314
rect 161848 77250 161900 77256
rect 161756 70032 161808 70038
rect 161756 69974 161808 69980
rect 161860 68785 161888 77250
rect 161952 69970 161980 79342
rect 162044 75138 162072 79562
rect 162136 77450 162164 79716
rect 162216 78668 162268 78674
rect 162216 78610 162268 78616
rect 162124 77444 162176 77450
rect 162124 77386 162176 77392
rect 162124 77240 162176 77246
rect 162124 77182 162176 77188
rect 162136 76770 162164 77182
rect 162124 76764 162176 76770
rect 162124 76706 162176 76712
rect 162124 76220 162176 76226
rect 162124 76162 162176 76168
rect 162032 75132 162084 75138
rect 162032 75074 162084 75080
rect 162136 72894 162164 76162
rect 162124 72888 162176 72894
rect 162124 72830 162176 72836
rect 162228 70394 162256 78610
rect 162308 77988 162360 77994
rect 162308 77930 162360 77936
rect 162320 76770 162348 77930
rect 162308 76764 162360 76770
rect 162308 76706 162360 76712
rect 162412 75478 162440 79784
rect 162722 79766 162774 79772
rect 162826 79778 162854 80036
rect 162918 79898 162946 80036
rect 162906 79892 162958 79898
rect 162906 79834 162958 79840
rect 163010 79778 163038 80036
rect 163102 79966 163130 80036
rect 163090 79960 163142 79966
rect 163090 79902 163142 79908
rect 162826 79750 162900 79778
rect 163010 79750 163084 79778
rect 162536 79727 162592 79736
rect 162492 79688 162544 79694
rect 162492 79630 162544 79636
rect 162584 79688 162636 79694
rect 162584 79630 162636 79636
rect 162676 79688 162728 79694
rect 162676 79630 162728 79636
rect 162504 77353 162532 79630
rect 162490 77344 162546 77353
rect 162490 77279 162546 77288
rect 162492 76968 162544 76974
rect 162492 76910 162544 76916
rect 162400 75472 162452 75478
rect 162400 75414 162452 75420
rect 162504 71466 162532 76910
rect 162596 76090 162624 79630
rect 162688 77314 162716 79630
rect 162768 79620 162820 79626
rect 162768 79562 162820 79568
rect 162676 77308 162728 77314
rect 162676 77250 162728 77256
rect 162584 76084 162636 76090
rect 162584 76026 162636 76032
rect 162780 74534 162808 79562
rect 162872 79422 162900 79750
rect 162860 79416 162912 79422
rect 162860 79358 162912 79364
rect 162872 79234 162900 79358
rect 162872 79206 162992 79234
rect 162860 77444 162912 77450
rect 162860 77386 162912 77392
rect 162872 76974 162900 77386
rect 162860 76968 162912 76974
rect 162860 76910 162912 76916
rect 162964 76226 162992 79206
rect 163056 77722 163084 79750
rect 163194 79744 163222 80036
rect 163286 79937 163314 80036
rect 163378 79966 163406 80036
rect 163470 79971 163498 80036
rect 163366 79960 163418 79966
rect 163272 79928 163328 79937
rect 163366 79902 163418 79908
rect 163456 79962 163512 79971
rect 163562 79966 163590 80036
rect 163456 79897 163512 79906
rect 163550 79960 163602 79966
rect 163550 79902 163602 79908
rect 163272 79863 163328 79872
rect 163320 79824 163372 79830
rect 163412 79824 163464 79830
rect 163320 79766 163372 79772
rect 163410 79792 163412 79801
rect 163654 79801 163682 80036
rect 163464 79792 163466 79801
rect 163148 79716 163222 79744
rect 163148 79626 163176 79716
rect 163136 79620 163188 79626
rect 163136 79562 163188 79568
rect 163228 79552 163280 79558
rect 163228 79494 163280 79500
rect 163240 78266 163268 79494
rect 163228 78260 163280 78266
rect 163228 78202 163280 78208
rect 163332 78112 163360 79766
rect 163410 79727 163466 79736
rect 163640 79792 163696 79801
rect 163640 79727 163696 79736
rect 163596 79688 163648 79694
rect 163746 79676 163774 80036
rect 163838 79898 163866 80036
rect 163826 79892 163878 79898
rect 163826 79834 163878 79840
rect 163930 79744 163958 80036
rect 163596 79630 163648 79636
rect 163700 79648 163774 79676
rect 163884 79716 163958 79744
rect 163412 78532 163464 78538
rect 163412 78474 163464 78480
rect 163148 78084 163360 78112
rect 163044 77716 163096 77722
rect 163044 77658 163096 77664
rect 162952 76220 163004 76226
rect 162952 76162 163004 76168
rect 163044 75472 163096 75478
rect 163044 75414 163096 75420
rect 162952 75132 163004 75138
rect 162952 75074 163004 75080
rect 162780 74506 162900 74534
rect 162676 73092 162728 73098
rect 162676 73034 162728 73040
rect 162688 72826 162716 73034
rect 162676 72820 162728 72826
rect 162676 72762 162728 72768
rect 162492 71460 162544 71466
rect 162492 71402 162544 71408
rect 162228 70366 162348 70394
rect 161940 69964 161992 69970
rect 161940 69906 161992 69912
rect 162320 69562 162348 70366
rect 162400 70304 162452 70310
rect 162400 70246 162452 70252
rect 162412 70038 162440 70246
rect 162400 70032 162452 70038
rect 162400 69974 162452 69980
rect 162308 69556 162360 69562
rect 162308 69498 162360 69504
rect 161846 68776 161902 68785
rect 161846 68711 161902 68720
rect 161662 68640 161718 68649
rect 161662 68575 161718 68584
rect 161860 64874 161888 68711
rect 161860 64846 162256 64874
rect 161572 64524 161624 64530
rect 161572 64466 161624 64472
rect 161480 44872 161532 44878
rect 161480 44814 161532 44820
rect 162228 31142 162256 64846
rect 162308 64524 162360 64530
rect 162308 64466 162360 64472
rect 162216 31136 162268 31142
rect 162216 31078 162268 31084
rect 162320 27062 162348 64466
rect 162308 27056 162360 27062
rect 162308 26998 162360 27004
rect 162412 25702 162440 69974
rect 162400 25696 162452 25702
rect 162400 25638 162452 25644
rect 162504 22982 162532 71402
rect 162584 70168 162636 70174
rect 162584 70110 162636 70116
rect 162596 69970 162624 70110
rect 162584 69964 162636 69970
rect 162584 69906 162636 69912
rect 162492 22976 162544 22982
rect 162492 22918 162544 22924
rect 162596 13190 162624 69906
rect 162688 14550 162716 72762
rect 162766 68640 162822 68649
rect 162766 68575 162822 68584
rect 162676 14544 162728 14550
rect 162676 14486 162728 14492
rect 162584 13184 162636 13190
rect 162584 13126 162636 13132
rect 162780 7750 162808 68575
rect 162872 60654 162900 74506
rect 162964 62082 162992 75074
rect 163056 66162 163084 75414
rect 163148 69970 163176 78084
rect 163226 78024 163282 78033
rect 163226 77959 163282 77968
rect 163240 73098 163268 77959
rect 163318 77888 163374 77897
rect 163318 77823 163374 77832
rect 163332 75138 163360 77823
rect 163320 75132 163372 75138
rect 163320 75074 163372 75080
rect 163424 74050 163452 78474
rect 163608 78062 163636 79630
rect 163596 78056 163648 78062
rect 163596 77998 163648 78004
rect 163700 77353 163728 79648
rect 163780 79552 163832 79558
rect 163780 79494 163832 79500
rect 163502 77344 163558 77353
rect 163502 77279 163558 77288
rect 163686 77344 163742 77353
rect 163686 77279 163742 77288
rect 163412 74044 163464 74050
rect 163412 73986 163464 73992
rect 163228 73092 163280 73098
rect 163228 73034 163280 73040
rect 163228 72888 163280 72894
rect 163228 72830 163280 72836
rect 163136 69964 163188 69970
rect 163136 69906 163188 69912
rect 163240 69873 163268 72830
rect 163226 69864 163282 69873
rect 163226 69799 163282 69808
rect 163044 66156 163096 66162
rect 163044 66098 163096 66104
rect 162952 62076 163004 62082
rect 162952 62018 163004 62024
rect 162860 60648 162912 60654
rect 162860 60590 162912 60596
rect 163516 53786 163544 77279
rect 163792 75478 163820 79494
rect 163884 77761 163912 79716
rect 164022 79676 164050 80036
rect 164114 79898 164142 80036
rect 164102 79892 164154 79898
rect 164102 79834 164154 79840
rect 164206 79778 164234 80036
rect 164298 79830 164326 80036
rect 163976 79648 164050 79676
rect 164160 79750 164234 79778
rect 164286 79824 164338 79830
rect 164286 79766 164338 79772
rect 163870 77752 163926 77761
rect 163870 77687 163926 77696
rect 163976 77294 164004 79648
rect 164056 79552 164108 79558
rect 164056 79494 164108 79500
rect 164068 78130 164096 79494
rect 164056 78124 164108 78130
rect 164056 78066 164108 78072
rect 164056 77920 164108 77926
rect 164160 77897 164188 79750
rect 164390 79744 164418 80036
rect 164482 79812 164510 80036
rect 164574 79937 164602 80036
rect 164560 79928 164616 79937
rect 164560 79863 164616 79872
rect 164666 79812 164694 80036
rect 164758 79966 164786 80036
rect 164850 79966 164878 80036
rect 164746 79960 164798 79966
rect 164746 79902 164798 79908
rect 164838 79960 164890 79966
rect 164838 79902 164890 79908
rect 164942 79898 164970 80036
rect 165034 79937 165062 80036
rect 165020 79928 165076 79937
rect 164930 79892 164982 79898
rect 165020 79863 165076 79872
rect 164930 79834 164982 79840
rect 164482 79784 164556 79812
rect 164666 79784 164786 79812
rect 164390 79716 164464 79744
rect 164240 79688 164292 79694
rect 164240 79630 164292 79636
rect 164330 79656 164386 79665
rect 164056 77862 164108 77868
rect 164146 77888 164202 77897
rect 163884 77266 164004 77294
rect 163780 75472 163832 75478
rect 163780 75414 163832 75420
rect 163884 72894 163912 77266
rect 163964 76424 164016 76430
rect 163964 76366 164016 76372
rect 163872 72888 163924 72894
rect 163872 72830 163924 72836
rect 163872 70236 163924 70242
rect 163872 70178 163924 70184
rect 163884 69970 163912 70178
rect 163872 69964 163924 69970
rect 163872 69906 163924 69912
rect 163780 66156 163832 66162
rect 163780 66098 163832 66104
rect 163504 53780 163556 53786
rect 163504 53722 163556 53728
rect 163792 22914 163820 66098
rect 163884 24274 163912 69906
rect 163976 29850 164004 76366
rect 164068 67250 164096 77862
rect 164146 77823 164202 77832
rect 164252 71738 164280 79630
rect 164330 79591 164386 79600
rect 164344 79150 164372 79591
rect 164332 79144 164384 79150
rect 164332 79086 164384 79092
rect 164330 78976 164386 78985
rect 164330 78911 164386 78920
rect 164344 76498 164372 78911
rect 164332 76492 164384 76498
rect 164332 76434 164384 76440
rect 164332 75132 164384 75138
rect 164332 75074 164384 75080
rect 164240 71732 164292 71738
rect 164240 71674 164292 71680
rect 164240 71596 164292 71602
rect 164240 71538 164292 71544
rect 164146 69864 164202 69873
rect 164146 69799 164202 69808
rect 164056 67244 164108 67250
rect 164056 67186 164108 67192
rect 163964 29844 164016 29850
rect 163964 29786 164016 29792
rect 163872 24268 163924 24274
rect 163872 24210 163924 24216
rect 163780 22908 163832 22914
rect 163780 22850 163832 22856
rect 164068 13258 164096 67186
rect 164056 13252 164108 13258
rect 164056 13194 164108 13200
rect 164160 11898 164188 69799
rect 164252 42226 164280 71538
rect 164344 63510 164372 75074
rect 164436 64870 164464 79716
rect 164528 75138 164556 79784
rect 164758 79778 164786 79784
rect 165126 79778 165154 80036
rect 165218 79830 165246 80036
rect 164758 79750 164924 79778
rect 164790 79656 164846 79665
rect 164608 79620 164660 79626
rect 164790 79591 164846 79600
rect 164608 79562 164660 79568
rect 164516 75132 164568 75138
rect 164516 75074 164568 75080
rect 164620 75018 164648 79562
rect 164700 79552 164752 79558
rect 164700 79494 164752 79500
rect 164528 74990 164648 75018
rect 164528 66026 164556 74990
rect 164608 74928 164660 74934
rect 164608 74870 164660 74876
rect 164620 68406 164648 74870
rect 164712 70038 164740 79494
rect 164700 70032 164752 70038
rect 164700 69974 164752 69980
rect 164804 69970 164832 79591
rect 164896 78538 164924 79750
rect 164988 79750 165154 79778
rect 165206 79824 165258 79830
rect 165310 79801 165338 80036
rect 165402 79898 165430 80036
rect 165390 79892 165442 79898
rect 165390 79834 165442 79840
rect 165494 79801 165522 80036
rect 165206 79766 165258 79772
rect 165296 79792 165352 79801
rect 164884 78532 164936 78538
rect 164884 78474 164936 78480
rect 164884 76492 164936 76498
rect 164884 76434 164936 76440
rect 164896 71602 164924 76434
rect 164988 74338 165016 79750
rect 165296 79727 165352 79736
rect 165480 79792 165536 79801
rect 165480 79727 165536 79736
rect 165586 79744 165614 80036
rect 165678 79898 165706 80036
rect 165666 79892 165718 79898
rect 165666 79834 165718 79840
rect 165770 79744 165798 80036
rect 165862 79937 165890 80036
rect 165848 79928 165904 79937
rect 165848 79863 165904 79872
rect 165954 79744 165982 80036
rect 166046 79898 166074 80036
rect 166034 79892 166086 79898
rect 166034 79834 166086 79840
rect 166138 79778 166166 80036
rect 166230 79898 166258 80036
rect 166218 79892 166270 79898
rect 166218 79834 166270 79840
rect 166092 79750 166166 79778
rect 165586 79716 165660 79744
rect 165770 79716 165844 79744
rect 165954 79716 166028 79744
rect 165160 79688 165212 79694
rect 165160 79630 165212 79636
rect 165252 79688 165304 79694
rect 165632 79676 165660 79716
rect 165632 79648 165752 79676
rect 165252 79630 165304 79636
rect 165068 79144 165120 79150
rect 165068 79086 165120 79092
rect 165080 76430 165108 79086
rect 165172 77926 165200 79630
rect 165160 77920 165212 77926
rect 165160 77862 165212 77868
rect 165068 76424 165120 76430
rect 165068 76366 165120 76372
rect 165264 74934 165292 79630
rect 165528 79620 165580 79626
rect 165528 79562 165580 79568
rect 165252 74928 165304 74934
rect 165252 74870 165304 74876
rect 164988 74310 165200 74338
rect 165172 72593 165200 74310
rect 165158 72584 165214 72593
rect 165158 72519 165214 72528
rect 165068 71732 165120 71738
rect 165068 71674 165120 71680
rect 164884 71596 164936 71602
rect 164884 71538 164936 71544
rect 165080 71330 165108 71674
rect 165068 71324 165120 71330
rect 165068 71266 165120 71272
rect 164792 69964 164844 69970
rect 164792 69906 164844 69912
rect 164608 68400 164660 68406
rect 164608 68342 164660 68348
rect 164516 66020 164568 66026
rect 164516 65962 164568 65968
rect 164424 64864 164476 64870
rect 164424 64806 164476 64812
rect 164436 63918 164464 64806
rect 164424 63912 164476 63918
rect 164424 63854 164476 63860
rect 164332 63504 164384 63510
rect 164332 63446 164384 63452
rect 164240 42220 164292 42226
rect 164240 42162 164292 42168
rect 165080 39506 165108 71266
rect 165068 39500 165120 39506
rect 165068 39442 165120 39448
rect 164884 31068 164936 31074
rect 164884 31010 164936 31016
rect 164148 11892 164200 11898
rect 164148 11834 164200 11840
rect 162768 7744 162820 7750
rect 162768 7686 162820 7692
rect 161388 4956 161440 4962
rect 161388 4898 161440 4904
rect 163688 3868 163740 3874
rect 163688 3810 163740 3816
rect 162492 3664 162544 3670
rect 162492 3606 162544 3612
rect 162504 480 162532 3606
rect 163700 480 163728 3810
rect 164516 3800 164568 3806
rect 164516 3742 164568 3748
rect 156574 354 156686 480
rect 156156 326 156686 354
rect 156574 -960 156686 326
rect 157770 -960 157882 480
rect 158874 -960 158986 480
rect 160070 -960 160182 480
rect 161266 -960 161378 480
rect 162462 -960 162574 480
rect 163658 -960 163770 480
rect 164528 218 164556 3742
rect 164896 3194 164924 31010
rect 165172 28422 165200 72519
rect 165540 71738 165568 79562
rect 165620 79552 165672 79558
rect 165620 79494 165672 79500
rect 165632 75002 165660 79494
rect 165724 79393 165752 79648
rect 165710 79384 165766 79393
rect 165710 79319 165766 79328
rect 165712 78328 165764 78334
rect 165712 78270 165764 78276
rect 165620 74996 165672 75002
rect 165620 74938 165672 74944
rect 165620 74860 165672 74866
rect 165620 74802 165672 74808
rect 165528 71732 165580 71738
rect 165528 71674 165580 71680
rect 165540 70394 165568 71674
rect 165344 70372 165396 70378
rect 165344 70314 165396 70320
rect 165448 70366 165568 70394
rect 165356 70038 165384 70314
rect 165344 70032 165396 70038
rect 165344 69974 165396 69980
rect 165252 63912 165304 63918
rect 165252 63854 165304 63860
rect 165160 28416 165212 28422
rect 165160 28358 165212 28364
rect 165264 18766 165292 63854
rect 165356 21418 165384 69974
rect 165344 21412 165396 21418
rect 165344 21354 165396 21360
rect 165252 18760 165304 18766
rect 165252 18702 165304 18708
rect 165448 16046 165476 70366
rect 165528 69964 165580 69970
rect 165528 69906 165580 69912
rect 165436 16040 165488 16046
rect 165436 15982 165488 15988
rect 165540 9110 165568 69906
rect 165528 9104 165580 9110
rect 165528 9046 165580 9052
rect 165632 6322 165660 74802
rect 165724 32434 165752 78270
rect 165816 78198 165844 79716
rect 165896 79620 165948 79626
rect 165896 79562 165948 79568
rect 165804 78192 165856 78198
rect 165804 78134 165856 78140
rect 165804 77988 165856 77994
rect 165804 77930 165856 77936
rect 165816 40866 165844 77930
rect 165908 64734 165936 79562
rect 166000 79506 166028 79716
rect 166092 79665 166120 79750
rect 166322 79744 166350 80036
rect 166414 79971 166442 80036
rect 166400 79962 166456 79971
rect 166400 79897 166456 79906
rect 166506 79778 166534 80036
rect 166598 79830 166626 80036
rect 166690 79966 166718 80036
rect 166782 79966 166810 80036
rect 166678 79960 166730 79966
rect 166678 79902 166730 79908
rect 166770 79960 166822 79966
rect 166770 79902 166822 79908
rect 166874 79898 166902 80036
rect 166862 79892 166914 79898
rect 166862 79834 166914 79840
rect 166966 79830 166994 80036
rect 167058 79903 167086 80036
rect 167044 79894 167100 79903
rect 166460 79750 166534 79778
rect 166586 79824 166638 79830
rect 166678 79824 166730 79830
rect 166586 79766 166638 79772
rect 166676 79792 166678 79801
rect 166954 79824 167006 79830
rect 167044 79829 167100 79838
rect 166730 79792 166732 79801
rect 166322 79716 166396 79744
rect 166078 79656 166134 79665
rect 166078 79591 166134 79600
rect 166172 79620 166224 79626
rect 166172 79562 166224 79568
rect 166000 79478 166120 79506
rect 165986 79384 166042 79393
rect 165986 79319 165988 79328
rect 166040 79319 166042 79328
rect 165988 79290 166040 79296
rect 165988 75132 166040 75138
rect 165988 75074 166040 75080
rect 166000 68882 166028 75074
rect 166092 68950 166120 79478
rect 166184 75138 166212 79562
rect 166264 79280 166316 79286
rect 166264 79222 166316 79228
rect 166276 78946 166304 79222
rect 166264 78940 166316 78946
rect 166264 78882 166316 78888
rect 166368 77858 166396 79716
rect 166460 78878 166488 79750
rect 166954 79766 167006 79772
rect 166676 79727 166732 79736
rect 167150 79744 167178 80036
rect 167242 79971 167270 80036
rect 167228 79962 167284 79971
rect 167228 79897 167284 79906
rect 167334 79830 167362 80036
rect 167426 79898 167454 80036
rect 167414 79892 167466 79898
rect 167414 79834 167466 79840
rect 167322 79824 167374 79830
rect 167518 79801 167546 80036
rect 167610 79898 167638 80036
rect 167598 79892 167650 79898
rect 167598 79834 167650 79840
rect 167322 79766 167374 79772
rect 167504 79792 167560 79801
rect 167150 79716 167224 79744
rect 167702 79744 167730 80036
rect 167794 79966 167822 80036
rect 167886 79966 167914 80036
rect 167978 79966 168006 80036
rect 168070 79971 168098 80036
rect 167782 79960 167834 79966
rect 167782 79902 167834 79908
rect 167874 79960 167926 79966
rect 167874 79902 167926 79908
rect 167966 79960 168018 79966
rect 167966 79902 168018 79908
rect 168056 79962 168112 79971
rect 168056 79897 168112 79906
rect 168162 79744 168190 80036
rect 168254 79937 168282 80036
rect 168346 79966 168374 80036
rect 168334 79960 168386 79966
rect 168240 79928 168296 79937
rect 168334 79902 168386 79908
rect 168438 79898 168466 80036
rect 168530 79966 168558 80036
rect 168622 79971 168650 80036
rect 168518 79960 168570 79966
rect 168518 79902 168570 79908
rect 168608 79962 168664 79971
rect 168240 79863 168296 79872
rect 168426 79892 168478 79898
rect 168608 79897 168664 79906
rect 168714 79898 168742 80036
rect 168806 79898 168834 80036
rect 168898 79971 168926 80036
rect 168884 79962 168940 79971
rect 168990 79966 169018 80036
rect 168426 79834 168478 79840
rect 168702 79892 168754 79898
rect 168702 79834 168754 79840
rect 168794 79892 168846 79898
rect 168884 79897 168940 79906
rect 168978 79960 169030 79966
rect 168978 79902 169030 79908
rect 169082 79898 169110 80036
rect 169174 79898 169202 80036
rect 169266 79966 169294 80036
rect 169254 79960 169306 79966
rect 169358 79937 169386 80036
rect 169254 79902 169306 79908
rect 169344 79928 169400 79937
rect 168794 79834 168846 79840
rect 169070 79892 169122 79898
rect 169070 79834 169122 79840
rect 169162 79892 169214 79898
rect 169344 79863 169400 79872
rect 169162 79834 169214 79840
rect 169450 79812 169478 80036
rect 169542 79966 169570 80036
rect 169530 79960 169582 79966
rect 169530 79902 169582 79908
rect 169634 79812 169662 80036
rect 167504 79727 167560 79736
rect 166724 79688 166776 79694
rect 166724 79630 166776 79636
rect 166816 79688 166868 79694
rect 166816 79630 166868 79636
rect 166998 79656 167054 79665
rect 166540 79348 166592 79354
rect 166540 79290 166592 79296
rect 166448 78872 166500 78878
rect 166448 78814 166500 78820
rect 166460 78334 166488 78814
rect 166448 78328 166500 78334
rect 166448 78270 166500 78276
rect 166552 77994 166580 79290
rect 166632 78260 166684 78266
rect 166632 78202 166684 78208
rect 166540 77988 166592 77994
rect 166540 77930 166592 77936
rect 166356 77852 166408 77858
rect 166356 77794 166408 77800
rect 166448 77308 166500 77314
rect 166448 77250 166500 77256
rect 166172 75132 166224 75138
rect 166172 75074 166224 75080
rect 166172 74996 166224 75002
rect 166172 74938 166224 74944
rect 166080 68944 166132 68950
rect 166080 68886 166132 68892
rect 165988 68876 166040 68882
rect 165988 68818 166040 68824
rect 166184 68474 166212 74938
rect 166172 68468 166224 68474
rect 166172 68410 166224 68416
rect 165896 64728 165948 64734
rect 165896 64670 165948 64676
rect 165908 63918 165936 64670
rect 165896 63912 165948 63918
rect 165896 63854 165948 63860
rect 166460 63374 166488 77250
rect 166644 70394 166672 78202
rect 166736 75914 166764 79630
rect 166828 79150 166856 79630
rect 166908 79620 166960 79626
rect 166998 79591 167054 79600
rect 166908 79562 166960 79568
rect 166920 79354 166948 79562
rect 166908 79348 166960 79354
rect 166908 79290 166960 79296
rect 166920 79257 166948 79290
rect 166906 79248 166962 79257
rect 166906 79183 166962 79192
rect 166816 79144 166868 79150
rect 166868 79104 166948 79132
rect 166816 79086 166868 79092
rect 166736 75886 166856 75914
rect 166828 71670 166856 75886
rect 166920 74866 166948 79104
rect 166908 74860 166960 74866
rect 166908 74802 166960 74808
rect 166816 71664 166868 71670
rect 166816 71606 166868 71612
rect 166828 70394 166856 71606
rect 166552 70366 166672 70394
rect 166736 70366 166856 70394
rect 166448 63368 166500 63374
rect 166448 63310 166500 63316
rect 166552 60518 166580 70366
rect 166632 63912 166684 63918
rect 166632 63854 166684 63860
rect 166540 60512 166592 60518
rect 166540 60454 166592 60460
rect 165804 40860 165856 40866
rect 165804 40802 165856 40808
rect 166644 33930 166672 63854
rect 166632 33924 166684 33930
rect 166632 33866 166684 33872
rect 165712 32428 165764 32434
rect 165712 32370 165764 32376
rect 166736 15978 166764 70366
rect 166816 68944 166868 68950
rect 166816 68886 166868 68892
rect 166828 68678 166856 68886
rect 167012 68882 167040 79591
rect 167090 79384 167146 79393
rect 167090 79319 167092 79328
rect 167144 79319 167146 79328
rect 167092 79290 167144 79296
rect 167196 77353 167224 79716
rect 167656 79716 167730 79744
rect 168024 79716 168190 79744
rect 168286 79792 168342 79801
rect 169404 79784 169478 79812
rect 169588 79784 169662 79812
rect 168286 79727 168342 79736
rect 168840 79756 168892 79762
rect 167276 79688 167328 79694
rect 167276 79630 167328 79636
rect 167460 79688 167512 79694
rect 167512 79648 167592 79676
rect 167460 79630 167512 79636
rect 167182 77344 167238 77353
rect 167182 77279 167238 77288
rect 167288 70394 167316 79630
rect 167368 79552 167420 79558
rect 167368 79494 167420 79500
rect 167380 77382 167408 79494
rect 167460 79484 167512 79490
rect 167460 79426 167512 79432
rect 167472 79393 167500 79426
rect 167458 79384 167514 79393
rect 167458 79319 167514 79328
rect 167564 78112 167592 79648
rect 167656 78928 167684 79716
rect 167918 79656 167974 79665
rect 168024 79642 168052 79716
rect 167974 79614 168052 79642
rect 168102 79656 168158 79665
rect 167918 79591 167974 79600
rect 168102 79591 168158 79600
rect 168196 79620 168248 79626
rect 167920 79552 167972 79558
rect 167920 79494 167972 79500
rect 168012 79552 168064 79558
rect 168012 79494 168064 79500
rect 167828 79416 167880 79422
rect 167828 79358 167880 79364
rect 167656 78900 167776 78928
rect 167564 78084 167684 78112
rect 167552 77988 167604 77994
rect 167552 77930 167604 77936
rect 167368 77376 167420 77382
rect 167368 77318 167420 77324
rect 167380 70786 167408 77318
rect 167564 75449 167592 77930
rect 167656 77790 167684 78084
rect 167644 77784 167696 77790
rect 167644 77726 167696 77732
rect 167644 77580 167696 77586
rect 167644 77522 167696 77528
rect 167656 75585 167684 77522
rect 167642 75576 167698 75585
rect 167642 75511 167698 75520
rect 167550 75440 167606 75449
rect 167550 75375 167606 75384
rect 167368 70780 167420 70786
rect 167368 70722 167420 70728
rect 167564 70394 167592 75375
rect 167104 70366 167316 70394
rect 167472 70366 167592 70394
rect 166908 68876 166960 68882
rect 166908 68818 166960 68824
rect 167000 68876 167052 68882
rect 167000 68818 167052 68824
rect 166920 68746 166948 68818
rect 167104 68814 167132 70366
rect 167092 68808 167144 68814
rect 167092 68750 167144 68756
rect 166908 68740 166960 68746
rect 166908 68682 166960 68688
rect 166816 68672 166868 68678
rect 166816 68614 166868 68620
rect 166724 15972 166776 15978
rect 166724 15914 166776 15920
rect 166828 10402 166856 68614
rect 166816 10396 166868 10402
rect 166816 10338 166868 10344
rect 166920 7682 166948 68682
rect 167472 43450 167500 70366
rect 167656 49094 167684 75511
rect 167748 71641 167776 78900
rect 167840 77586 167868 79358
rect 167828 77580 167880 77586
rect 167828 77522 167880 77528
rect 167828 75948 167880 75954
rect 167828 75890 167880 75896
rect 167734 71632 167790 71641
rect 167734 71567 167790 71576
rect 167736 70780 167788 70786
rect 167736 70722 167788 70728
rect 167644 49088 167696 49094
rect 167644 49030 167696 49036
rect 167460 43444 167512 43450
rect 167460 43386 167512 43392
rect 167748 42158 167776 70722
rect 167736 42152 167788 42158
rect 167736 42094 167788 42100
rect 167840 39438 167868 75890
rect 167932 71777 167960 79494
rect 168024 78266 168052 79494
rect 168012 78260 168064 78266
rect 168012 78202 168064 78208
rect 168116 77994 168144 79591
rect 168196 79562 168248 79568
rect 168104 77988 168156 77994
rect 168104 77930 168156 77936
rect 168208 76974 168236 79562
rect 168196 76968 168248 76974
rect 168196 76910 168248 76916
rect 168012 76084 168064 76090
rect 168012 76026 168064 76032
rect 167918 71768 167974 71777
rect 167918 71703 167974 71712
rect 168024 70394 168052 76026
rect 168208 75954 168236 76910
rect 168196 75948 168248 75954
rect 168196 75890 168248 75896
rect 168300 75177 168328 79727
rect 168840 79698 168892 79704
rect 169208 79756 169260 79762
rect 169208 79698 169260 79704
rect 168472 79688 168524 79694
rect 168378 79656 168434 79665
rect 168472 79630 168524 79636
rect 168564 79688 168616 79694
rect 168616 79648 168788 79676
rect 168564 79630 168616 79636
rect 168378 79591 168434 79600
rect 168286 75168 168342 75177
rect 168286 75103 168342 75112
rect 168286 71768 168342 71777
rect 168286 71703 168342 71712
rect 168194 71632 168250 71641
rect 168194 71567 168250 71576
rect 168024 70366 168144 70394
rect 167920 68876 167972 68882
rect 167920 68818 167972 68824
rect 167828 39432 167880 39438
rect 167828 39374 167880 39380
rect 167932 17406 167960 68818
rect 168012 68808 168064 68814
rect 168012 68750 168064 68756
rect 167920 17400 167972 17406
rect 167920 17342 167972 17348
rect 168024 17338 168052 68750
rect 168116 66978 168144 70366
rect 168104 66972 168156 66978
rect 168104 66914 168156 66920
rect 168012 17332 168064 17338
rect 168012 17274 168064 17280
rect 167000 17264 167052 17270
rect 167000 17206 167052 17212
rect 167012 16574 167040 17206
rect 167012 16546 167224 16574
rect 166908 7676 166960 7682
rect 166908 7618 166960 7624
rect 165620 6316 165672 6322
rect 165620 6258 165672 6264
rect 166080 3596 166132 3602
rect 166080 3538 166132 3544
rect 164884 3188 164936 3194
rect 164884 3130 164936 3136
rect 166092 480 166120 3538
rect 167196 480 167224 16546
rect 168116 14618 168144 66914
rect 168104 14612 168156 14618
rect 168104 14554 168156 14560
rect 168208 11830 168236 71567
rect 168196 11824 168248 11830
rect 168196 11766 168248 11772
rect 168300 4894 168328 71703
rect 168392 52426 168420 79591
rect 168484 75478 168512 79630
rect 168564 79552 168616 79558
rect 168564 79494 168616 79500
rect 168472 75472 168524 75478
rect 168472 75414 168524 75420
rect 168472 74928 168524 74934
rect 168472 74870 168524 74876
rect 168380 52420 168432 52426
rect 168380 52362 168432 52368
rect 168484 38010 168512 74870
rect 168576 48278 168604 79494
rect 168656 79484 168708 79490
rect 168656 79426 168708 79432
rect 168668 79393 168696 79426
rect 168654 79384 168710 79393
rect 168654 79319 168710 79328
rect 168656 78668 168708 78674
rect 168656 78610 168708 78616
rect 168668 57934 168696 78610
rect 168760 78402 168788 79648
rect 168748 78396 168800 78402
rect 168748 78338 168800 78344
rect 168748 74996 168800 75002
rect 168748 74938 168800 74944
rect 168760 64666 168788 74938
rect 168852 68270 168880 79698
rect 169024 79620 169076 79626
rect 169024 79562 169076 79568
rect 169116 79620 169168 79626
rect 169116 79562 169168 79568
rect 169036 78334 169064 79562
rect 169024 78328 169076 78334
rect 169024 78270 169076 78276
rect 169024 75472 169076 75478
rect 169024 75414 169076 75420
rect 168932 75132 168984 75138
rect 168932 75074 168984 75080
rect 168840 68264 168892 68270
rect 168840 68206 168892 68212
rect 168944 68202 168972 75074
rect 169036 70038 169064 75414
rect 169128 75002 169156 79562
rect 169220 78674 169248 79698
rect 169300 79552 169352 79558
rect 169300 79494 169352 79500
rect 169208 78668 169260 78674
rect 169208 78610 169260 78616
rect 169312 77294 169340 79494
rect 169404 79121 169432 79784
rect 169484 79688 169536 79694
rect 169484 79630 169536 79636
rect 169390 79112 169446 79121
rect 169390 79047 169446 79056
rect 169220 77266 169340 77294
rect 169116 74996 169168 75002
rect 169116 74938 169168 74944
rect 169220 71097 169248 77266
rect 169404 75914 169432 79047
rect 169312 75886 169432 75914
rect 169312 74934 169340 75886
rect 169496 75138 169524 79630
rect 169588 75313 169616 79784
rect 169726 79744 169754 80036
rect 169818 79830 169846 80036
rect 169910 79966 169938 80036
rect 170002 79971 170030 80036
rect 169898 79960 169950 79966
rect 169898 79902 169950 79908
rect 169988 79962 170044 79971
rect 170094 79966 170122 80036
rect 170186 79966 170214 80036
rect 169988 79897 170044 79906
rect 170082 79960 170134 79966
rect 170082 79902 170134 79908
rect 170174 79960 170226 79966
rect 170278 79937 170306 80036
rect 170174 79902 170226 79908
rect 170264 79928 170320 79937
rect 170264 79863 170320 79872
rect 169806 79824 169858 79830
rect 170036 79824 170088 79830
rect 169806 79766 169858 79772
rect 170034 79792 170036 79801
rect 170088 79792 170090 79801
rect 169680 79716 169754 79744
rect 170034 79727 170090 79736
rect 170128 79756 170180 79762
rect 169680 78674 169708 79716
rect 170370 79744 170398 80036
rect 170462 79830 170490 80036
rect 170554 79971 170582 80036
rect 170540 79962 170596 79971
rect 170540 79897 170596 79906
rect 170646 79898 170674 80036
rect 170634 79892 170686 79898
rect 170634 79834 170686 79840
rect 170450 79824 170502 79830
rect 170450 79766 170502 79772
rect 170128 79698 170180 79704
rect 170232 79716 170398 79744
rect 170738 79744 170766 80036
rect 170830 79971 170858 80036
rect 170816 79962 170872 79971
rect 170816 79897 170872 79906
rect 170922 79778 170950 80036
rect 171014 79966 171042 80036
rect 171002 79960 171054 79966
rect 171002 79902 171054 79908
rect 171106 79898 171134 80036
rect 171094 79892 171146 79898
rect 171094 79834 171146 79840
rect 170876 79750 170950 79778
rect 170738 79716 170812 79744
rect 170034 79656 170090 79665
rect 169852 79620 169904 79626
rect 169852 79562 169904 79568
rect 169944 79620 169996 79626
rect 170034 79591 170090 79600
rect 169944 79562 169996 79568
rect 169758 79384 169814 79393
rect 169758 79319 169814 79328
rect 169668 78668 169720 78674
rect 169668 78610 169720 78616
rect 169574 75304 169630 75313
rect 169574 75239 169630 75248
rect 169484 75132 169536 75138
rect 169484 75074 169536 75080
rect 169300 74928 169352 74934
rect 169300 74870 169352 74876
rect 169206 71088 169262 71097
rect 169206 71023 169262 71032
rect 169024 70032 169076 70038
rect 169024 69974 169076 69980
rect 169484 70032 169536 70038
rect 169484 69974 169536 69980
rect 168932 68196 168984 68202
rect 168932 68138 168984 68144
rect 168748 64660 168800 64666
rect 168748 64602 168800 64608
rect 168656 57928 168708 57934
rect 168656 57870 168708 57876
rect 168656 49020 168708 49026
rect 168656 48962 168708 48968
rect 168564 48272 168616 48278
rect 168564 48214 168616 48220
rect 168472 38004 168524 38010
rect 168472 37946 168524 37952
rect 168668 16574 168696 48962
rect 169496 38078 169524 69974
rect 169576 68264 169628 68270
rect 169576 68206 169628 68212
rect 169484 38072 169536 38078
rect 169484 38014 169536 38020
rect 169588 31074 169616 68206
rect 169668 68196 169720 68202
rect 169668 68138 169720 68144
rect 169576 31068 169628 31074
rect 169576 31010 169628 31016
rect 169680 17270 169708 68138
rect 169772 67046 169800 79319
rect 169864 72894 169892 79562
rect 169956 78742 169984 79562
rect 169944 78736 169996 78742
rect 169944 78678 169996 78684
rect 170048 78577 170076 79591
rect 170034 78568 170090 78577
rect 170034 78503 170090 78512
rect 169852 72888 169904 72894
rect 169852 72830 169904 72836
rect 170140 70394 170168 79698
rect 170232 74497 170260 79716
rect 170310 79656 170366 79665
rect 170310 79591 170366 79600
rect 170496 79620 170548 79626
rect 170218 74488 170274 74497
rect 170218 74423 170274 74432
rect 170324 72350 170352 79591
rect 170496 79562 170548 79568
rect 170508 78713 170536 79562
rect 170680 79552 170732 79558
rect 170680 79494 170732 79500
rect 170588 79416 170640 79422
rect 170588 79358 170640 79364
rect 170600 78826 170628 79358
rect 170692 78928 170720 79494
rect 170784 78996 170812 79716
rect 170876 79422 170904 79750
rect 171198 79744 171226 80036
rect 171060 79716 171226 79744
rect 170956 79688 171008 79694
rect 170954 79656 170956 79665
rect 171008 79656 171010 79665
rect 170954 79591 171010 79600
rect 170956 79552 171008 79558
rect 170956 79494 171008 79500
rect 170864 79416 170916 79422
rect 170864 79358 170916 79364
rect 170784 78968 170904 78996
rect 170692 78900 170812 78928
rect 170600 78798 170720 78826
rect 170588 78736 170640 78742
rect 170494 78704 170550 78713
rect 170588 78678 170640 78684
rect 170494 78639 170550 78648
rect 170600 76498 170628 78678
rect 170692 76809 170720 78798
rect 170678 76800 170734 76809
rect 170678 76735 170734 76744
rect 170588 76492 170640 76498
rect 170588 76434 170640 76440
rect 170494 75984 170550 75993
rect 170494 75919 170550 75928
rect 170312 72344 170364 72350
rect 170312 72286 170364 72292
rect 169864 70366 170168 70394
rect 169864 68610 169892 70366
rect 169852 68604 169904 68610
rect 169852 68546 169904 68552
rect 169760 67040 169812 67046
rect 169760 66982 169812 66988
rect 169760 57248 169812 57254
rect 169760 57190 169812 57196
rect 169668 17264 169720 17270
rect 169668 17206 169720 17212
rect 169772 16574 169800 57190
rect 170508 42090 170536 75919
rect 170600 75698 170628 76434
rect 170692 75993 170720 76735
rect 170678 75984 170734 75993
rect 170678 75919 170734 75928
rect 170600 75670 170720 75698
rect 170586 74488 170642 74497
rect 170586 74423 170642 74432
rect 170600 73681 170628 74423
rect 170586 73672 170642 73681
rect 170586 73607 170642 73616
rect 170496 42084 170548 42090
rect 170496 42026 170548 42032
rect 170600 35358 170628 73607
rect 170692 36650 170720 75670
rect 170784 73778 170812 78900
rect 170876 74390 170904 78968
rect 170864 74384 170916 74390
rect 170864 74326 170916 74332
rect 170772 73772 170824 73778
rect 170772 73714 170824 73720
rect 170680 36644 170732 36650
rect 170680 36586 170732 36592
rect 170588 35352 170640 35358
rect 170588 35294 170640 35300
rect 170402 35184 170458 35193
rect 170402 35119 170458 35128
rect 168668 16546 169616 16574
rect 169772 16546 170352 16574
rect 168288 4888 168340 4894
rect 168288 4830 168340 4836
rect 168380 3188 168432 3194
rect 168380 3130 168432 3136
rect 168392 480 168420 3130
rect 169588 480 169616 16546
rect 164854 218 164966 480
rect 164528 190 164966 218
rect 164854 -960 164966 190
rect 166050 -960 166162 480
rect 167154 -960 167266 480
rect 168350 -960 168462 480
rect 169546 -960 169658 480
rect 170324 354 170352 16546
rect 170416 3602 170444 35119
rect 170784 29782 170812 73714
rect 170772 29776 170824 29782
rect 170772 29718 170824 29724
rect 170876 26994 170904 74326
rect 170968 71369 170996 79494
rect 171060 78742 171088 79716
rect 171290 79676 171318 80036
rect 171382 79830 171410 80036
rect 171474 79966 171502 80036
rect 171566 79966 171594 80036
rect 171658 79971 171686 80036
rect 171462 79960 171514 79966
rect 171462 79902 171514 79908
rect 171554 79960 171606 79966
rect 171554 79902 171606 79908
rect 171644 79962 171700 79971
rect 171644 79897 171700 79906
rect 171370 79824 171422 79830
rect 171370 79766 171422 79772
rect 171750 79744 171778 80036
rect 171244 79648 171318 79676
rect 171612 79716 171778 79744
rect 171138 79384 171194 79393
rect 171138 79319 171194 79328
rect 171048 78736 171100 78742
rect 171048 78678 171100 78684
rect 171048 72888 171100 72894
rect 171048 72830 171100 72836
rect 170954 71360 171010 71369
rect 170954 71295 171010 71304
rect 170956 68604 171008 68610
rect 170956 68546 171008 68552
rect 170864 26988 170916 26994
rect 170864 26930 170916 26936
rect 170968 14482 170996 68546
rect 170956 14476 171008 14482
rect 170956 14418 171008 14424
rect 171060 13122 171088 72830
rect 171152 24206 171180 79319
rect 171244 75750 171272 79648
rect 171324 79552 171376 79558
rect 171324 79494 171376 79500
rect 171416 79552 171468 79558
rect 171416 79494 171468 79500
rect 171508 79552 171560 79558
rect 171508 79494 171560 79500
rect 171232 75744 171284 75750
rect 171232 75686 171284 75692
rect 171336 74458 171364 79494
rect 171428 78033 171456 79494
rect 171414 78024 171470 78033
rect 171414 77959 171470 77968
rect 171520 75886 171548 79494
rect 171508 75880 171560 75886
rect 171508 75822 171560 75828
rect 171324 74452 171376 74458
rect 171324 74394 171376 74400
rect 171612 73001 171640 79716
rect 171842 79676 171870 80036
rect 171934 79971 171962 80036
rect 171920 79962 171976 79971
rect 171920 79897 171976 79906
rect 172026 79830 172054 80036
rect 172014 79824 172066 79830
rect 172014 79766 172066 79772
rect 171796 79648 171870 79676
rect 171968 79688 172020 79694
rect 171692 78736 171744 78742
rect 171692 78678 171744 78684
rect 171704 74118 171732 78678
rect 171796 75614 171824 79648
rect 172118 79676 172146 80036
rect 171968 79630 172020 79636
rect 172072 79648 172146 79676
rect 171980 78742 172008 79630
rect 171968 78736 172020 78742
rect 171968 78678 172020 78684
rect 171876 78192 171928 78198
rect 171876 78134 171928 78140
rect 171888 77926 171916 78134
rect 171876 77920 171928 77926
rect 171876 77862 171928 77868
rect 172072 77294 172100 79648
rect 172210 79608 172238 80036
rect 172302 79971 172330 80036
rect 172288 79962 172344 79971
rect 172288 79897 172344 79906
rect 172394 79744 172422 80036
rect 172486 79966 172514 80036
rect 172578 79966 172606 80036
rect 172474 79960 172526 79966
rect 172474 79902 172526 79908
rect 172566 79960 172618 79966
rect 172566 79902 172618 79908
rect 172474 79824 172526 79830
rect 172670 79801 172698 80036
rect 172762 79971 172790 80036
rect 172748 79962 172804 79971
rect 172854 79966 172882 80036
rect 172748 79897 172804 79906
rect 172842 79960 172894 79966
rect 172842 79902 172894 79908
rect 172474 79766 172526 79772
rect 172656 79792 172712 79801
rect 172164 79580 172238 79608
rect 172348 79716 172422 79744
rect 172164 78713 172192 79580
rect 172244 79484 172296 79490
rect 172244 79426 172296 79432
rect 172256 78946 172284 79426
rect 172244 78940 172296 78946
rect 172244 78882 172296 78888
rect 172244 78736 172296 78742
rect 172150 78704 172206 78713
rect 172244 78678 172296 78684
rect 172150 78639 172206 78648
rect 171980 77266 172100 77294
rect 171784 75608 171836 75614
rect 171784 75550 171836 75556
rect 171692 74112 171744 74118
rect 171692 74054 171744 74060
rect 171598 72992 171654 73001
rect 171598 72927 171654 72936
rect 171230 71768 171286 71777
rect 171230 71703 171286 71712
rect 171244 71505 171272 71703
rect 171230 71496 171286 71505
rect 171230 71431 171286 71440
rect 171232 70780 171284 70786
rect 171232 70722 171284 70728
rect 171244 70106 171272 70722
rect 171704 70394 171732 74054
rect 171980 70786 172008 77266
rect 172060 75880 172112 75886
rect 172060 75822 172112 75828
rect 171968 70780 172020 70786
rect 171968 70722 172020 70728
rect 171612 70366 171732 70394
rect 171232 70100 171284 70106
rect 171232 70042 171284 70048
rect 171612 64874 171640 70366
rect 171612 64846 172008 64874
rect 171980 40798 172008 64846
rect 171968 40792 172020 40798
rect 171968 40734 172020 40740
rect 172072 36582 172100 75822
rect 172256 74610 172284 78678
rect 172348 75818 172376 79716
rect 172486 79676 172514 79766
rect 172656 79727 172712 79736
rect 172794 79792 172850 79801
rect 172946 79744 172974 80036
rect 173038 79801 173066 80036
rect 172794 79727 172850 79736
rect 172440 79665 172514 79676
rect 172426 79656 172514 79665
rect 172482 79648 172514 79656
rect 172702 79656 172758 79665
rect 172426 79591 172482 79600
rect 172612 79620 172664 79626
rect 172702 79591 172758 79600
rect 172612 79562 172664 79568
rect 172520 79416 172572 79422
rect 172520 79358 172572 79364
rect 172428 78736 172480 78742
rect 172428 78678 172480 78684
rect 172440 77602 172468 78678
rect 172532 77722 172560 79358
rect 172520 77716 172572 77722
rect 172520 77658 172572 77664
rect 172440 77574 172560 77602
rect 172336 75812 172388 75818
rect 172336 75754 172388 75760
rect 172256 74582 172468 74610
rect 172244 74452 172296 74458
rect 172244 74394 172296 74400
rect 172256 74186 172284 74394
rect 172244 74180 172296 74186
rect 172244 74122 172296 74128
rect 172152 70100 172204 70106
rect 172152 70042 172204 70048
rect 172060 36576 172112 36582
rect 172060 36518 172112 36524
rect 172164 25566 172192 70042
rect 172256 28354 172284 74122
rect 172334 72992 172390 73001
rect 172334 72927 172390 72936
rect 172244 28348 172296 28354
rect 172244 28290 172296 28296
rect 172348 26926 172376 72927
rect 172440 72457 172468 74582
rect 172426 72448 172482 72457
rect 172426 72383 172482 72392
rect 172336 26920 172388 26926
rect 172336 26862 172388 26868
rect 172440 25634 172468 72383
rect 172532 37942 172560 77574
rect 172624 49706 172652 79562
rect 172716 76090 172744 79591
rect 172808 76158 172836 79727
rect 172900 79716 172974 79744
rect 173024 79792 173080 79801
rect 173024 79727 173080 79736
rect 173130 79744 173158 80036
rect 173222 79937 173250 80036
rect 173208 79928 173264 79937
rect 173314 79898 173342 80036
rect 173208 79863 173264 79872
rect 173302 79892 173354 79898
rect 173302 79834 173354 79840
rect 173406 79830 173434 80036
rect 173498 79937 173526 80036
rect 173484 79928 173540 79937
rect 173484 79863 173540 79872
rect 173394 79824 173446 79830
rect 173254 79792 173310 79801
rect 173130 79736 173254 79744
rect 173590 79778 173618 80036
rect 173394 79766 173446 79772
rect 173130 79727 173310 79736
rect 173544 79750 173618 79778
rect 173130 79716 173296 79727
rect 172900 77314 172928 79716
rect 173348 79688 173400 79694
rect 173070 79656 173126 79665
rect 172980 79620 173032 79626
rect 173254 79656 173310 79665
rect 173070 79591 173126 79600
rect 173164 79620 173216 79626
rect 172980 79562 173032 79568
rect 172888 77308 172940 77314
rect 172888 77250 172940 77256
rect 172796 76152 172848 76158
rect 172796 76094 172848 76100
rect 172704 76084 172756 76090
rect 172704 76026 172756 76032
rect 172992 75970 173020 79562
rect 173084 78946 173112 79591
rect 173348 79630 173400 79636
rect 173440 79688 173492 79694
rect 173544 79665 173572 79750
rect 173682 79744 173710 80036
rect 173774 79971 173802 80036
rect 173760 79962 173816 79971
rect 173866 79966 173894 80036
rect 173760 79897 173816 79906
rect 173854 79960 173906 79966
rect 173854 79902 173906 79908
rect 173958 79830 173986 80036
rect 174050 79830 174078 80036
rect 174142 79830 174170 80036
rect 174234 79966 174262 80036
rect 174222 79960 174274 79966
rect 174222 79902 174274 79908
rect 173946 79824 173998 79830
rect 173946 79766 173998 79772
rect 174038 79824 174090 79830
rect 174038 79766 174090 79772
rect 174130 79824 174182 79830
rect 174326 79812 174354 80036
rect 174130 79766 174182 79772
rect 174234 79784 174354 79812
rect 173682 79716 173756 79744
rect 173440 79630 173492 79636
rect 173530 79656 173586 79665
rect 173254 79591 173310 79600
rect 173164 79562 173216 79568
rect 173072 78940 173124 78946
rect 173072 78882 173124 78888
rect 172716 75942 173020 75970
rect 172716 61878 172744 75942
rect 173176 73154 173204 79562
rect 173268 78554 173296 79591
rect 173360 79393 173388 79630
rect 173346 79384 173402 79393
rect 173346 79319 173402 79328
rect 173360 78742 173388 79319
rect 173348 78736 173400 78742
rect 173348 78678 173400 78684
rect 173452 78656 173480 79630
rect 173530 79591 173586 79600
rect 173624 79620 173676 79626
rect 173624 79562 173676 79568
rect 173636 78792 173664 79562
rect 173728 79540 173756 79716
rect 174234 79676 174262 79784
rect 174418 79778 174446 80036
rect 174510 79966 174538 80036
rect 174602 79966 174630 80036
rect 174694 79971 174722 80036
rect 174498 79960 174550 79966
rect 174496 79928 174498 79937
rect 174590 79960 174642 79966
rect 174550 79928 174552 79937
rect 174590 79902 174642 79908
rect 174680 79962 174736 79971
rect 174680 79897 174736 79906
rect 174786 79898 174814 80036
rect 174878 79898 174906 80036
rect 174970 79971 174998 80036
rect 174956 79962 175012 79971
rect 174496 79863 174552 79872
rect 174774 79892 174826 79898
rect 174774 79834 174826 79840
rect 174866 79892 174918 79898
rect 174956 79897 175012 79906
rect 174866 79834 174918 79840
rect 175062 79812 175090 80036
rect 175154 79966 175182 80036
rect 175246 79966 175274 80036
rect 175142 79960 175194 79966
rect 175142 79902 175194 79908
rect 175234 79960 175286 79966
rect 175338 79937 175366 80036
rect 175234 79902 175286 79908
rect 175324 79928 175380 79937
rect 175430 79898 175458 80036
rect 175522 79898 175550 80036
rect 175614 79966 175642 80036
rect 175602 79960 175654 79966
rect 175602 79902 175654 79908
rect 175324 79863 175380 79872
rect 175418 79892 175470 79898
rect 175418 79834 175470 79840
rect 175510 79892 175562 79898
rect 175510 79834 175562 79840
rect 175706 79830 175734 80036
rect 175798 79971 175826 80036
rect 175784 79962 175840 79971
rect 175784 79897 175840 79906
rect 175890 79898 175918 80036
rect 175982 79966 176010 80036
rect 176074 79971 176102 80036
rect 175970 79960 176022 79966
rect 175970 79902 176022 79908
rect 176060 79962 176116 79971
rect 175878 79892 175930 79898
rect 176060 79897 176116 79906
rect 175878 79834 175930 79840
rect 175694 79824 175746 79830
rect 174542 79792 174598 79801
rect 174418 79750 174492 79778
rect 174360 79688 174412 79694
rect 173990 79656 174046 79665
rect 174234 79648 174308 79676
rect 173990 79591 174046 79600
rect 174084 79620 174136 79626
rect 173728 79512 173848 79540
rect 173636 78764 173756 78792
rect 173452 78628 173572 78656
rect 173268 78526 173480 78554
rect 173348 76356 173400 76362
rect 173348 76298 173400 76304
rect 172808 73126 173204 73154
rect 172808 65890 172836 73126
rect 173360 71505 173388 76298
rect 173346 71496 173402 71505
rect 173346 71431 173402 71440
rect 173452 71346 173480 78526
rect 173544 76673 173572 78628
rect 173728 78305 173756 78764
rect 173714 78296 173770 78305
rect 173714 78231 173770 78240
rect 173714 78160 173770 78169
rect 173714 78095 173770 78104
rect 173728 76945 173756 78095
rect 173714 76936 173770 76945
rect 173714 76871 173770 76880
rect 173530 76664 173586 76673
rect 173530 76599 173586 76608
rect 173544 76022 173572 76599
rect 173622 76392 173678 76401
rect 173622 76327 173678 76336
rect 173532 76016 173584 76022
rect 173532 75958 173584 75964
rect 172900 71318 173480 71346
rect 172900 67114 172928 71318
rect 173636 70394 173664 76327
rect 173728 76106 173756 76871
rect 173820 76362 173848 79512
rect 174004 78452 174032 79591
rect 174084 79562 174136 79568
rect 173912 78424 174032 78452
rect 173808 76356 173860 76362
rect 173808 76298 173860 76304
rect 173728 76078 173848 76106
rect 173716 76016 173768 76022
rect 173716 75958 173768 75964
rect 172992 70366 173664 70394
rect 172992 69601 173020 70366
rect 172978 69592 173034 69601
rect 172978 69527 173034 69536
rect 173622 69592 173678 69601
rect 173622 69527 173678 69536
rect 172888 67108 172940 67114
rect 172888 67050 172940 67056
rect 172796 65884 172848 65890
rect 172796 65826 172848 65832
rect 172704 61872 172756 61878
rect 172704 61814 172756 61820
rect 172612 49700 172664 49706
rect 172612 49642 172664 49648
rect 172520 37936 172572 37942
rect 172520 37878 172572 37884
rect 172428 25628 172480 25634
rect 172428 25570 172480 25576
rect 171784 25560 171836 25566
rect 171784 25502 171836 25508
rect 172152 25560 172204 25566
rect 172152 25502 172204 25508
rect 171140 24200 171192 24206
rect 171140 24142 171192 24148
rect 171048 13116 171100 13122
rect 171048 13058 171100 13064
rect 170404 3596 170456 3602
rect 170404 3538 170456 3544
rect 171796 3534 171824 25502
rect 173636 24138 173664 69527
rect 173624 24132 173676 24138
rect 173624 24074 173676 24080
rect 173728 22846 173756 75958
rect 173716 22840 173768 22846
rect 173716 22782 173768 22788
rect 173820 22778 173848 76078
rect 173808 22772 173860 22778
rect 173808 22714 173860 22720
rect 173912 4826 173940 78424
rect 173992 77444 174044 77450
rect 173992 77386 174044 77392
rect 174004 57866 174032 77386
rect 174096 76650 174124 79562
rect 174096 76622 174216 76650
rect 174084 76356 174136 76362
rect 174084 76298 174136 76304
rect 174096 64598 174124 76298
rect 174188 67182 174216 76622
rect 174280 67318 174308 79648
rect 174360 79630 174412 79636
rect 174464 79642 174492 79750
rect 175062 79784 175136 79812
rect 174542 79727 174544 79736
rect 174596 79727 174598 79736
rect 174912 79756 174964 79762
rect 174544 79698 174596 79704
rect 174912 79698 174964 79704
rect 174634 79656 174690 79665
rect 174372 76226 174400 79630
rect 174464 79614 174584 79642
rect 174556 78810 174584 79614
rect 174634 79591 174690 79600
rect 174728 79620 174780 79626
rect 174544 78804 174596 78810
rect 174544 78746 174596 78752
rect 174648 76362 174676 79591
rect 174728 79562 174780 79568
rect 174740 77586 174768 79562
rect 174728 77580 174780 77586
rect 174728 77522 174780 77528
rect 174636 76356 174688 76362
rect 174636 76298 174688 76304
rect 174360 76220 174412 76226
rect 174360 76162 174412 76168
rect 174924 74534 174952 79698
rect 175004 79620 175056 79626
rect 175004 79562 175056 79568
rect 175016 77450 175044 79562
rect 175004 77444 175056 77450
rect 175004 77386 175056 77392
rect 175004 76220 175056 76226
rect 175004 76162 175056 76168
rect 175016 75138 175044 76162
rect 175004 75132 175056 75138
rect 175004 75074 175056 75080
rect 174832 74506 174952 74534
rect 174832 70394 174860 74506
rect 175016 70786 175044 75074
rect 175108 73846 175136 79784
rect 175694 79766 175746 79772
rect 175188 79756 175240 79762
rect 175188 79698 175240 79704
rect 175280 79756 175332 79762
rect 175280 79698 175332 79704
rect 175464 79756 175516 79762
rect 175464 79698 175516 79704
rect 175924 79756 175976 79762
rect 175924 79698 175976 79704
rect 176016 79756 176068 79762
rect 176166 79744 176194 80036
rect 176258 79971 176286 80036
rect 176244 79962 176300 79971
rect 176244 79897 176300 79906
rect 176350 79744 176378 80036
rect 176442 79898 176470 80036
rect 176430 79892 176482 79898
rect 176430 79834 176482 79840
rect 176166 79716 176240 79744
rect 176350 79716 176424 79744
rect 176016 79698 176068 79704
rect 175200 79665 175228 79698
rect 175186 79656 175242 79665
rect 175186 79591 175242 79600
rect 175292 78554 175320 79698
rect 175372 78872 175424 78878
rect 175372 78814 175424 78820
rect 175200 78526 175320 78554
rect 175096 73840 175148 73846
rect 175096 73782 175148 73788
rect 175004 70780 175056 70786
rect 175004 70722 175056 70728
rect 174372 70366 174860 70394
rect 174372 67454 174400 70366
rect 174360 67448 174412 67454
rect 174360 67390 174412 67396
rect 175004 67448 175056 67454
rect 175004 67390 175056 67396
rect 175016 67318 175044 67390
rect 174268 67312 174320 67318
rect 174268 67254 174320 67260
rect 174912 67312 174964 67318
rect 174912 67254 174964 67260
rect 175004 67312 175056 67318
rect 175004 67254 175056 67260
rect 174176 67176 174228 67182
rect 174176 67118 174228 67124
rect 174820 67176 174872 67182
rect 174820 67118 174872 67124
rect 174832 66842 174860 67118
rect 174924 66910 174952 67254
rect 174912 66904 174964 66910
rect 174912 66846 174964 66852
rect 174820 66836 174872 66842
rect 174820 66778 174872 66784
rect 174084 64592 174136 64598
rect 174084 64534 174136 64540
rect 173992 57860 174044 57866
rect 173992 57802 174044 57808
rect 174832 40730 174860 66778
rect 174820 40724 174872 40730
rect 174820 40666 174872 40672
rect 174924 35290 174952 66846
rect 174912 35284 174964 35290
rect 174912 35226 174964 35232
rect 175016 15910 175044 67254
rect 175004 15904 175056 15910
rect 175004 15846 175056 15852
rect 175108 10334 175136 73782
rect 175200 71233 175228 78526
rect 175278 78432 175334 78441
rect 175278 78367 175334 78376
rect 175186 71224 175242 71233
rect 175186 71159 175242 71168
rect 175188 70780 175240 70786
rect 175188 70722 175240 70728
rect 175096 10328 175148 10334
rect 175096 10270 175148 10276
rect 175200 7614 175228 70722
rect 175292 8974 175320 78367
rect 175384 11762 175412 78814
rect 175476 78198 175504 79698
rect 175740 79688 175792 79694
rect 175738 79656 175740 79665
rect 175792 79656 175794 79665
rect 175556 79620 175608 79626
rect 175556 79562 175608 79568
rect 175648 79620 175700 79626
rect 175738 79591 175794 79600
rect 175648 79562 175700 79568
rect 175464 78192 175516 78198
rect 175464 78134 175516 78140
rect 175464 77512 175516 77518
rect 175464 77454 175516 77460
rect 175476 29646 175504 77454
rect 175568 67182 175596 79562
rect 175660 77353 175688 79562
rect 175936 78713 175964 79698
rect 176028 78878 176056 79698
rect 176016 78872 176068 78878
rect 176016 78814 176068 78820
rect 175922 78704 175978 78713
rect 175844 78662 175922 78690
rect 175738 77480 175794 77489
rect 175738 77415 175794 77424
rect 175646 77344 175702 77353
rect 175646 77279 175702 77288
rect 175648 76968 175700 76974
rect 175648 76910 175700 76916
rect 175556 67176 175608 67182
rect 175556 67118 175608 67124
rect 175660 33862 175688 76910
rect 175752 69873 175780 77415
rect 175844 76974 175872 78662
rect 175922 78639 175978 78648
rect 176106 77616 176162 77625
rect 176106 77551 176162 77560
rect 175832 76968 175884 76974
rect 175924 76968 175976 76974
rect 175832 76910 175884 76916
rect 175922 76936 175924 76945
rect 175976 76936 175978 76945
rect 175922 76871 175978 76880
rect 175832 75880 175884 75886
rect 175832 75822 175884 75828
rect 175844 75682 175872 75822
rect 175832 75676 175884 75682
rect 175832 75618 175884 75624
rect 175830 72856 175886 72865
rect 175830 72791 175886 72800
rect 175738 69864 175794 69873
rect 175738 69799 175794 69808
rect 175844 64874 175872 72791
rect 176120 70394 176148 77551
rect 176212 72729 176240 79716
rect 176292 79620 176344 79626
rect 176292 79562 176344 79568
rect 176304 77450 176332 79562
rect 176396 78305 176424 79716
rect 176534 79540 176562 80036
rect 176626 79778 176654 80036
rect 176718 79966 176746 80036
rect 176810 79966 176838 80036
rect 176706 79960 176758 79966
rect 176706 79902 176758 79908
rect 176798 79960 176850 79966
rect 176798 79902 176850 79908
rect 176902 79812 176930 80036
rect 176994 79937 177022 80036
rect 176980 79928 177036 79937
rect 177086 79898 177114 80036
rect 176980 79863 177036 79872
rect 177074 79892 177126 79898
rect 177074 79834 177126 79840
rect 176810 79784 176930 79812
rect 177026 79792 177082 79801
rect 176810 79778 176838 79784
rect 176626 79750 176700 79778
rect 176488 79512 176562 79540
rect 176382 78296 176438 78305
rect 176382 78231 176438 78240
rect 176384 78192 176436 78198
rect 176384 78134 176436 78140
rect 176396 77489 176424 78134
rect 176382 77480 176438 77489
rect 176292 77444 176344 77450
rect 176382 77415 176438 77424
rect 176292 77386 176344 77392
rect 176396 73154 176424 77415
rect 176488 77081 176516 79512
rect 176672 79393 176700 79750
rect 176764 79750 176838 79778
rect 176658 79384 176714 79393
rect 176658 79319 176714 79328
rect 176672 77518 176700 79319
rect 176764 78792 176792 79750
rect 177178 79744 177206 80036
rect 177026 79727 177082 79736
rect 176764 78764 176976 78792
rect 176844 78668 176896 78674
rect 176844 78610 176896 78616
rect 176660 77512 176712 77518
rect 176660 77454 176712 77460
rect 176568 77444 176620 77450
rect 176568 77386 176620 77392
rect 176474 77072 176530 77081
rect 176474 77007 176530 77016
rect 176396 73126 176516 73154
rect 176198 72720 176254 72729
rect 176198 72655 176254 72664
rect 176120 70366 176424 70394
rect 176292 67448 176344 67454
rect 176292 67390 176344 67396
rect 176304 66910 176332 67390
rect 176292 66904 176344 66910
rect 176292 66846 176344 66852
rect 175844 64846 176332 64874
rect 176304 39370 176332 64846
rect 176292 39364 176344 39370
rect 176292 39306 176344 39312
rect 176396 35222 176424 70366
rect 176384 35216 176436 35222
rect 176384 35158 176436 35164
rect 175648 33856 175700 33862
rect 175648 33798 175700 33804
rect 176488 29714 176516 73126
rect 176580 72865 176608 77386
rect 176660 75880 176712 75886
rect 176660 75822 176712 75828
rect 176672 75342 176700 75822
rect 176660 75336 176712 75342
rect 176660 75278 176712 75284
rect 176752 75336 176804 75342
rect 176752 75278 176804 75284
rect 176660 74996 176712 75002
rect 176660 74938 176712 74944
rect 176566 72856 176622 72865
rect 176566 72791 176622 72800
rect 176566 72720 176622 72729
rect 176566 72655 176622 72664
rect 175924 29708 175976 29714
rect 175924 29650 175976 29656
rect 176476 29708 176528 29714
rect 176476 29650 176528 29656
rect 175464 29640 175516 29646
rect 175464 29582 175516 29588
rect 175372 11756 175424 11762
rect 175372 11698 175424 11704
rect 175280 8968 175332 8974
rect 175280 8910 175332 8916
rect 175188 7608 175240 7614
rect 175188 7550 175240 7556
rect 173900 4820 173952 4826
rect 173900 4762 173952 4768
rect 171968 3732 172020 3738
rect 171968 3674 172020 3680
rect 171784 3528 171836 3534
rect 171784 3470 171836 3476
rect 171980 480 172008 3674
rect 174268 3596 174320 3602
rect 174268 3538 174320 3544
rect 173164 3528 173216 3534
rect 173164 3470 173216 3476
rect 173176 480 173204 3470
rect 174280 480 174308 3538
rect 175464 3324 175516 3330
rect 175464 3266 175516 3272
rect 175476 480 175504 3266
rect 175936 3058 175964 29650
rect 176580 6254 176608 72655
rect 176672 44130 176700 74938
rect 176764 46918 176792 75278
rect 176856 51066 176884 78610
rect 176948 57798 176976 78764
rect 177040 75342 177068 79727
rect 177132 79716 177206 79744
rect 177028 75336 177080 75342
rect 177028 75278 177080 75284
rect 177132 70394 177160 79716
rect 177270 79676 177298 80036
rect 177362 79744 177390 80036
rect 177454 79812 177482 80036
rect 177546 79971 177574 80036
rect 177532 79962 177588 79971
rect 177532 79897 177588 79906
rect 177638 79914 177666 80036
rect 177638 79886 177712 79914
rect 177684 79830 177712 79886
rect 177580 79824 177632 79830
rect 177454 79784 177528 79812
rect 177362 79716 177436 79744
rect 177270 79648 177344 79676
rect 177212 76152 177264 76158
rect 177212 76094 177264 76100
rect 177224 75342 177252 76094
rect 177212 75336 177264 75342
rect 177212 75278 177264 75284
rect 177316 75002 177344 79648
rect 177304 74996 177356 75002
rect 177304 74938 177356 74944
rect 177408 74390 177436 79716
rect 177500 78305 177528 79784
rect 177580 79766 177632 79772
rect 177672 79824 177724 79830
rect 177672 79766 177724 79772
rect 177592 78674 177620 79766
rect 177776 79626 177804 80106
rect 177856 79960 177908 79966
rect 177856 79902 177908 79908
rect 177764 79620 177816 79626
rect 177764 79562 177816 79568
rect 177580 78668 177632 78674
rect 177580 78610 177632 78616
rect 177486 78296 177542 78305
rect 177486 78231 177542 78240
rect 177580 77580 177632 77586
rect 177580 77522 177632 77528
rect 177488 77308 177540 77314
rect 177488 77250 177540 77256
rect 177500 75041 177528 77250
rect 177486 75032 177542 75041
rect 177486 74967 177542 74976
rect 177396 74384 177448 74390
rect 177396 74326 177448 74332
rect 177408 70394 177436 74326
rect 177040 70366 177160 70394
rect 177316 70366 177436 70394
rect 177040 68513 177068 70366
rect 177026 68504 177082 68513
rect 177026 68439 177082 68448
rect 177316 64874 177344 70366
rect 177592 68950 177620 77522
rect 177868 76945 177896 79902
rect 178040 79892 178092 79898
rect 178040 79834 178092 79840
rect 178052 77722 178080 79834
rect 178696 78538 178724 80582
rect 178788 78742 178816 80582
rect 180522 80543 180578 80552
rect 179236 80096 179288 80102
rect 179236 80038 179288 80044
rect 179248 79506 179276 80038
rect 180536 80034 180564 80543
rect 185766 80472 185822 80481
rect 185766 80407 185822 80416
rect 184202 80200 184258 80209
rect 184202 80135 184258 80144
rect 180524 80028 180576 80034
rect 180524 79970 180576 79976
rect 180522 79928 180578 79937
rect 180522 79863 180578 79872
rect 179510 79656 179566 79665
rect 179510 79591 179566 79600
rect 179064 79478 179276 79506
rect 179420 79552 179472 79558
rect 179420 79494 179472 79500
rect 178776 78736 178828 78742
rect 178776 78678 178828 78684
rect 178684 78532 178736 78538
rect 178684 78474 178736 78480
rect 178040 77716 178092 77722
rect 178040 77658 178092 77664
rect 178052 77294 178080 77658
rect 177960 77266 178080 77294
rect 177854 76936 177910 76945
rect 177854 76871 177910 76880
rect 177764 75336 177816 75342
rect 177764 75278 177816 75284
rect 177580 68944 177632 68950
rect 177580 68886 177632 68892
rect 177316 64846 177712 64874
rect 176936 57792 176988 57798
rect 176936 57734 176988 57740
rect 176844 51060 176896 51066
rect 176844 51002 176896 51008
rect 176752 46912 176804 46918
rect 176752 46854 176804 46860
rect 176660 44124 176712 44130
rect 176660 44066 176712 44072
rect 177684 33794 177712 64846
rect 177672 33788 177724 33794
rect 177672 33730 177724 33736
rect 177776 28286 177804 75278
rect 177764 28280 177816 28286
rect 177764 28222 177816 28228
rect 177868 18698 177896 76871
rect 177856 18692 177908 18698
rect 177856 18634 177908 18640
rect 177960 18630 177988 77266
rect 178408 76084 178460 76090
rect 178408 76026 178460 76032
rect 178420 75478 178448 76026
rect 178408 75472 178460 75478
rect 178408 75414 178460 75420
rect 178038 68232 178094 68241
rect 178038 68167 178094 68176
rect 177948 18624 178000 18630
rect 177948 18566 178000 18572
rect 178052 16574 178080 68167
rect 178052 16546 178632 16574
rect 176568 6248 176620 6254
rect 176568 6190 176620 6196
rect 176660 3392 176712 3398
rect 176660 3334 176712 3340
rect 175924 3052 175976 3058
rect 175924 2994 175976 3000
rect 176672 480 176700 3334
rect 177856 3052 177908 3058
rect 177856 2994 177908 3000
rect 177868 480 177896 2994
rect 170742 354 170854 480
rect 170324 326 170854 354
rect 170742 -960 170854 326
rect 171938 -960 172050 480
rect 173134 -960 173246 480
rect 174238 -960 174350 480
rect 175434 -960 175546 480
rect 176630 -960 176742 480
rect 177826 -960 177938 480
rect 178604 354 178632 16546
rect 178696 3738 178724 78474
rect 178776 78124 178828 78130
rect 178776 78066 178828 78072
rect 178788 78033 178816 78066
rect 178774 78024 178830 78033
rect 178774 77959 178830 77968
rect 178788 3806 178816 77959
rect 179064 75914 179092 79478
rect 179248 79422 179276 79478
rect 179144 79416 179196 79422
rect 179144 79358 179196 79364
rect 179236 79416 179288 79422
rect 179236 79358 179288 79364
rect 179156 78130 179184 79358
rect 179144 78124 179196 78130
rect 179144 78066 179196 78072
rect 179156 75970 179184 78066
rect 179328 78056 179380 78062
rect 179328 77998 179380 78004
rect 179156 75942 179276 75970
rect 179064 75886 179184 75914
rect 178958 75304 179014 75313
rect 178958 75239 179014 75248
rect 178776 3800 178828 3806
rect 178776 3742 178828 3748
rect 178684 3732 178736 3738
rect 178684 3674 178736 3680
rect 178972 3534 179000 75239
rect 179050 75168 179106 75177
rect 179050 75103 179106 75112
rect 179064 3670 179092 75103
rect 179156 6458 179184 75886
rect 179144 6452 179196 6458
rect 179144 6394 179196 6400
rect 179248 3942 179276 75942
rect 179236 3936 179288 3942
rect 179236 3878 179288 3884
rect 179340 3874 179368 77998
rect 179432 16574 179460 79494
rect 179524 78033 179552 79591
rect 180156 79348 180208 79354
rect 180156 79290 180208 79296
rect 179510 78024 179566 78033
rect 179510 77959 179566 77968
rect 180064 76696 180116 76702
rect 180064 76638 180116 76644
rect 179432 16546 180012 16574
rect 179328 3868 179380 3874
rect 179328 3810 179380 3816
rect 179052 3664 179104 3670
rect 179052 3606 179104 3612
rect 178960 3528 179012 3534
rect 178960 3470 179012 3476
rect 179984 3482 180012 16546
rect 180076 4078 180104 76638
rect 180168 69494 180196 79290
rect 180536 78441 180564 79863
rect 181628 79824 181680 79830
rect 181628 79766 181680 79772
rect 181352 79552 181404 79558
rect 181352 79494 181404 79500
rect 180522 78432 180578 78441
rect 180522 78367 180578 78376
rect 180708 78192 180760 78198
rect 180708 78134 180760 78140
rect 180720 77994 180748 78134
rect 180524 77988 180576 77994
rect 180524 77930 180576 77936
rect 180708 77988 180760 77994
rect 180708 77930 180760 77936
rect 180432 76288 180484 76294
rect 180432 76230 180484 76236
rect 180444 74610 180472 76230
rect 180536 74746 180564 77930
rect 180708 77852 180760 77858
rect 180708 77794 180760 77800
rect 180720 76294 180748 77794
rect 180708 76288 180760 76294
rect 180708 76230 180760 76236
rect 180800 75064 180852 75070
rect 180800 75006 180852 75012
rect 180536 74718 180748 74746
rect 180444 74582 180656 74610
rect 180524 72412 180576 72418
rect 180524 72354 180576 72360
rect 180156 69488 180208 69494
rect 180156 69430 180208 69436
rect 180064 4072 180116 4078
rect 180064 4014 180116 4020
rect 179984 3454 180288 3482
rect 180536 3466 180564 72354
rect 180628 6526 180656 74582
rect 180720 6662 180748 74718
rect 180812 16574 180840 75006
rect 181364 72826 181392 79494
rect 181444 78464 181496 78470
rect 181444 78406 181496 78412
rect 181456 77382 181484 78406
rect 181640 77897 181668 79766
rect 181904 77920 181956 77926
rect 181626 77888 181682 77897
rect 181904 77862 181956 77868
rect 182086 77888 182142 77897
rect 181626 77823 181682 77832
rect 181628 77784 181680 77790
rect 181628 77726 181680 77732
rect 181444 77376 181496 77382
rect 181444 77318 181496 77324
rect 181640 76362 181668 77726
rect 181916 76514 181944 77862
rect 182086 77823 182142 77832
rect 181916 76486 182036 76514
rect 181628 76356 181680 76362
rect 181628 76298 181680 76304
rect 181904 76356 181956 76362
rect 181904 76298 181956 76304
rect 181626 72856 181682 72865
rect 181352 72820 181404 72826
rect 181626 72791 181682 72800
rect 181352 72762 181404 72768
rect 181640 72593 181668 72791
rect 181442 72584 181498 72593
rect 181442 72519 181498 72528
rect 181626 72584 181682 72593
rect 181626 72519 181682 72528
rect 181456 72321 181484 72519
rect 181442 72312 181498 72321
rect 181442 72247 181498 72256
rect 181444 71188 181496 71194
rect 181444 71130 181496 71136
rect 181812 71188 181864 71194
rect 181812 71130 181864 71136
rect 180812 16546 181024 16574
rect 180708 6656 180760 6662
rect 180708 6598 180760 6604
rect 180616 6520 180668 6526
rect 180616 6462 180668 6468
rect 180260 480 180288 3454
rect 180524 3460 180576 3466
rect 180524 3402 180576 3408
rect 179022 354 179134 480
rect 178604 326 179134 354
rect 179022 -960 179134 326
rect 180218 -960 180330 480
rect 180996 354 181024 16546
rect 181456 2922 181484 71130
rect 181824 71097 181852 71130
rect 181810 71088 181866 71097
rect 181810 71023 181866 71032
rect 181824 4146 181852 71023
rect 181916 6390 181944 76298
rect 182008 6594 182036 76486
rect 181996 6588 182048 6594
rect 181996 6530 182048 6536
rect 181904 6384 181956 6390
rect 181904 6326 181956 6332
rect 182100 6186 182128 77823
rect 182824 76628 182876 76634
rect 182824 76570 182876 76576
rect 182088 6180 182140 6186
rect 182088 6122 182140 6128
rect 181812 4140 181864 4146
rect 181812 4082 181864 4088
rect 182836 4010 182864 76570
rect 183560 69692 183612 69698
rect 183560 69634 183612 69640
rect 183572 16574 183600 69634
rect 183572 16546 183784 16574
rect 182824 4004 182876 4010
rect 182824 3946 182876 3952
rect 181444 2916 181496 2922
rect 181444 2858 181496 2864
rect 182548 2916 182600 2922
rect 182548 2858 182600 2864
rect 182560 480 182588 2858
rect 183756 480 183784 16546
rect 184216 9042 184244 80135
rect 184480 80096 184532 80102
rect 184480 80038 184532 80044
rect 184388 79348 184440 79354
rect 184388 79290 184440 79296
rect 184296 71120 184348 71126
rect 184296 71062 184348 71068
rect 184204 9036 184256 9042
rect 184204 8978 184256 8984
rect 184308 3398 184336 71062
rect 184400 66978 184428 79290
rect 184492 69834 184520 80038
rect 184940 76560 184992 76566
rect 184940 76502 184992 76508
rect 184480 69828 184532 69834
rect 184480 69770 184532 69776
rect 184388 66972 184440 66978
rect 184388 66914 184440 66920
rect 184952 11694 184980 76502
rect 185032 75880 185084 75886
rect 185032 75822 185084 75828
rect 185124 75880 185176 75886
rect 185124 75822 185176 75828
rect 184940 11688 184992 11694
rect 184940 11630 184992 11636
rect 185044 6914 185072 75822
rect 185136 75342 185164 75822
rect 185124 75336 185176 75342
rect 185124 75278 185176 75284
rect 185398 70408 185454 70417
rect 185398 70343 185454 70352
rect 185412 69562 185440 70343
rect 185400 69556 185452 69562
rect 185400 69498 185452 69504
rect 185412 69086 185440 69498
rect 185400 69080 185452 69086
rect 185400 69022 185452 69028
rect 185780 64874 185808 80407
rect 186320 68536 186372 68542
rect 186320 68478 186372 68484
rect 186332 68134 186360 68478
rect 186320 68128 186372 68134
rect 186320 68070 186372 68076
rect 185688 64846 185808 64874
rect 185688 64530 185716 64846
rect 185676 64524 185728 64530
rect 185676 64466 185728 64472
rect 185584 64184 185636 64190
rect 185584 64126 185636 64132
rect 184952 6886 185072 6914
rect 184296 3392 184348 3398
rect 184296 3334 184348 3340
rect 184952 480 184980 6886
rect 185596 3602 185624 64126
rect 186608 56273 186636 195638
rect 186700 68542 186728 199854
rect 186780 145852 186832 145858
rect 186780 145794 186832 145800
rect 186688 68536 186740 68542
rect 186688 68478 186740 68484
rect 186792 68066 186820 145794
rect 187160 144265 187188 284922
rect 199396 267034 199424 404330
rect 203536 287706 203564 630634
rect 203524 287700 203576 287706
rect 203524 287642 203576 287648
rect 204168 276684 204220 276690
rect 204168 276626 204220 276632
rect 204180 276078 204208 276626
rect 203064 276072 203116 276078
rect 203064 276014 203116 276020
rect 204168 276072 204220 276078
rect 204168 276014 204220 276020
rect 199384 267028 199436 267034
rect 199384 266970 199436 266976
rect 192024 265668 192076 265674
rect 192024 265610 192076 265616
rect 188252 265260 188304 265266
rect 188252 265202 188304 265208
rect 187516 264988 187568 264994
rect 187516 264930 187568 264936
rect 187332 260228 187384 260234
rect 187332 260170 187384 260176
rect 187240 146804 187292 146810
rect 187240 146746 187292 146752
rect 187146 144256 187202 144265
rect 187146 144191 187202 144200
rect 186964 141568 187016 141574
rect 186964 141510 187016 141516
rect 186872 137828 186924 137834
rect 186872 137770 186924 137776
rect 186884 73030 186912 137770
rect 186976 73982 187004 141510
rect 187148 141432 187200 141438
rect 187148 141374 187200 141380
rect 187054 139360 187110 139369
rect 187054 139295 187110 139304
rect 186964 73976 187016 73982
rect 186964 73918 187016 73924
rect 186872 73024 186924 73030
rect 186872 72966 186924 72972
rect 187068 70854 187096 139295
rect 187160 74254 187188 141374
rect 187252 80102 187280 146746
rect 187344 142050 187372 260170
rect 187422 213888 187478 213897
rect 187422 213823 187478 213832
rect 187436 143698 187464 213823
rect 187528 144129 187556 264930
rect 188066 262576 188122 262585
rect 188066 262511 188122 262520
rect 187792 262268 187844 262274
rect 187792 262210 187844 262216
rect 187700 259684 187752 259690
rect 187700 259626 187752 259632
rect 187712 259418 187740 259626
rect 187700 259412 187752 259418
rect 187700 259354 187752 259360
rect 187804 258618 187832 262210
rect 187884 260364 187936 260370
rect 187884 260306 187936 260312
rect 187712 258590 187832 258618
rect 187608 199844 187660 199850
rect 187608 199786 187660 199792
rect 187514 144120 187570 144129
rect 187514 144055 187570 144064
rect 187436 143670 187556 143698
rect 187424 143540 187476 143546
rect 187424 143482 187476 143488
rect 187332 142044 187384 142050
rect 187332 141986 187384 141992
rect 187332 140888 187384 140894
rect 187332 140830 187384 140836
rect 187344 132494 187372 140830
rect 187436 137834 187464 143482
rect 187528 143478 187556 143670
rect 187516 143472 187568 143478
rect 187516 143414 187568 143420
rect 187620 138145 187648 199786
rect 187712 198762 187740 258590
rect 187792 258528 187844 258534
rect 187792 258470 187844 258476
rect 187700 198756 187752 198762
rect 187700 198698 187752 198704
rect 187804 151814 187832 258470
rect 187712 151786 187832 151814
rect 187712 144401 187740 151786
rect 187792 144900 187844 144906
rect 187792 144842 187844 144848
rect 187698 144392 187754 144401
rect 187698 144327 187754 144336
rect 187700 139732 187752 139738
rect 187700 139674 187752 139680
rect 187712 139641 187740 139674
rect 187698 139632 187754 139641
rect 187698 139567 187754 139576
rect 187606 138136 187662 138145
rect 187606 138071 187662 138080
rect 187424 137828 187476 137834
rect 187424 137770 187476 137776
rect 187344 132466 187464 132494
rect 187436 89842 187464 132466
rect 187436 89814 187740 89842
rect 187240 80096 187292 80102
rect 187240 80038 187292 80044
rect 187330 79928 187386 79937
rect 187330 79863 187386 79872
rect 187148 74248 187200 74254
rect 187148 74190 187200 74196
rect 187344 72758 187372 79863
rect 187332 72752 187384 72758
rect 187332 72694 187384 72700
rect 187712 70990 187740 89814
rect 187700 70984 187752 70990
rect 187700 70926 187752 70932
rect 187056 70848 187108 70854
rect 187056 70790 187108 70796
rect 186780 68060 186832 68066
rect 186780 68002 186832 68008
rect 187238 63472 187294 63481
rect 187238 63407 187294 63416
rect 187252 63374 187280 63407
rect 187240 63368 187292 63374
rect 187240 63310 187292 63316
rect 187252 62150 187280 63310
rect 187240 62144 187292 62150
rect 187240 62086 187292 62092
rect 187698 57216 187754 57225
rect 187698 57151 187754 57160
rect 186594 56264 186650 56273
rect 186594 56199 186650 56208
rect 187712 16574 187740 57151
rect 187804 55214 187832 144842
rect 187896 141982 187924 260306
rect 187976 259820 188028 259826
rect 187976 259762 188028 259768
rect 187988 143002 188016 259762
rect 188080 258534 188108 262511
rect 188160 259752 188212 259758
rect 188160 259694 188212 259700
rect 188068 258528 188120 258534
rect 188068 258470 188120 258476
rect 188172 150278 188200 259694
rect 188264 156602 188292 265202
rect 189356 263696 189408 263702
rect 189356 263638 189408 263644
rect 188526 262984 188582 262993
rect 188526 262919 188582 262928
rect 188540 262585 188568 262919
rect 188526 262576 188582 262585
rect 188526 262511 188582 262520
rect 189172 262336 189224 262342
rect 189172 262278 189224 262284
rect 188344 261452 188396 261458
rect 188344 261394 188396 261400
rect 188356 193186 188384 261394
rect 188894 259992 188950 260001
rect 188894 259927 188950 259936
rect 188712 195628 188764 195634
rect 188712 195570 188764 195576
rect 188436 195356 188488 195362
rect 188436 195298 188488 195304
rect 188344 193180 188396 193186
rect 188344 193122 188396 193128
rect 188344 178084 188396 178090
rect 188344 178026 188396 178032
rect 188252 156596 188304 156602
rect 188252 156538 188304 156544
rect 188252 151836 188304 151842
rect 188252 151778 188304 151784
rect 188160 150272 188212 150278
rect 188160 150214 188212 150220
rect 188264 148374 188292 151778
rect 188252 148368 188304 148374
rect 188252 148310 188304 148316
rect 188160 147416 188212 147422
rect 188160 147358 188212 147364
rect 188068 144832 188120 144838
rect 188068 144774 188120 144780
rect 187976 142996 188028 143002
rect 187976 142938 188028 142944
rect 187884 141976 187936 141982
rect 187884 141918 187936 141924
rect 187976 140480 188028 140486
rect 187976 140422 188028 140428
rect 187884 62008 187936 62014
rect 187884 61950 187936 61956
rect 187896 61538 187924 61950
rect 187884 61532 187936 61538
rect 187884 61474 187936 61480
rect 187988 56574 188016 140422
rect 188080 74322 188108 144774
rect 188068 74316 188120 74322
rect 188068 74258 188120 74264
rect 188080 73914 188108 74258
rect 188068 73908 188120 73914
rect 188068 73850 188120 73856
rect 188172 69630 188200 147358
rect 188252 144832 188304 144838
rect 188252 144774 188304 144780
rect 188264 144294 188292 144774
rect 188252 144288 188304 144294
rect 188252 144230 188304 144236
rect 188356 144226 188384 178026
rect 188344 144220 188396 144226
rect 188344 144162 188396 144168
rect 188344 140344 188396 140350
rect 188344 140286 188396 140292
rect 188250 139224 188306 139233
rect 188250 139159 188306 139168
rect 188264 70922 188292 139159
rect 188356 79218 188384 140286
rect 188448 118017 188476 195298
rect 188620 148912 188672 148918
rect 188620 148854 188672 148860
rect 188528 141636 188580 141642
rect 188528 141578 188580 141584
rect 188434 118008 188490 118017
rect 188434 117943 188490 117952
rect 188540 81433 188568 141578
rect 188632 138718 188660 148854
rect 188620 138712 188672 138718
rect 188620 138654 188672 138660
rect 188526 81424 188582 81433
rect 188526 81359 188582 81368
rect 188436 81116 188488 81122
rect 188436 81058 188488 81064
rect 188448 80850 188476 81058
rect 188436 80844 188488 80850
rect 188436 80786 188488 80792
rect 188344 79212 188396 79218
rect 188344 79154 188396 79160
rect 188252 70916 188304 70922
rect 188252 70858 188304 70864
rect 188160 69624 188212 69630
rect 188160 69566 188212 69572
rect 188342 64152 188398 64161
rect 188342 64087 188398 64096
rect 187976 56568 188028 56574
rect 187976 56510 188028 56516
rect 187988 55894 188016 56510
rect 187976 55888 188028 55894
rect 187976 55830 188028 55836
rect 187804 55186 187924 55214
rect 187792 41404 187844 41410
rect 187792 41346 187844 41352
rect 187804 41002 187832 41346
rect 187792 40996 187844 41002
rect 187792 40938 187844 40944
rect 187790 38584 187846 38593
rect 187896 38570 187924 55186
rect 187846 38542 187924 38570
rect 187790 38519 187846 38528
rect 187804 37913 187832 38519
rect 187790 37904 187846 37913
rect 187790 37839 187846 37848
rect 187712 16546 188292 16574
rect 186136 11688 186188 11694
rect 186136 11630 186188 11636
rect 185584 3596 185636 3602
rect 185584 3538 185636 3544
rect 186148 480 186176 11630
rect 187424 4140 187476 4146
rect 187424 4082 187476 4088
rect 187436 3602 187464 4082
rect 187332 3596 187384 3602
rect 187332 3538 187384 3544
rect 187424 3596 187476 3602
rect 187424 3538 187476 3544
rect 187344 480 187372 3538
rect 188264 3482 188292 16546
rect 188356 4146 188384 64087
rect 188724 61538 188752 195570
rect 188804 144356 188856 144362
rect 188804 144298 188856 144304
rect 188712 61532 188764 61538
rect 188712 61474 188764 61480
rect 188816 41002 188844 144298
rect 188908 143041 188936 259927
rect 189184 192302 189212 262278
rect 189264 200320 189316 200326
rect 189264 200262 189316 200268
rect 189172 192296 189224 192302
rect 189172 192238 189224 192244
rect 189172 146668 189224 146674
rect 189172 146610 189224 146616
rect 188894 143032 188950 143041
rect 188894 142967 188950 142976
rect 189080 140616 189132 140622
rect 189078 140584 189080 140593
rect 189132 140584 189134 140593
rect 189078 140519 189134 140528
rect 189078 81560 189134 81569
rect 189078 81495 189134 81504
rect 189092 73846 189120 81495
rect 189080 73840 189132 73846
rect 189080 73782 189132 73788
rect 189080 67584 189132 67590
rect 189080 67526 189132 67532
rect 189092 66910 189120 67526
rect 189184 67386 189212 146610
rect 189172 67380 189224 67386
rect 189172 67322 189224 67328
rect 189080 66904 189132 66910
rect 189080 66846 189132 66852
rect 189276 66722 189304 200262
rect 189368 143206 189396 263638
rect 189540 262948 189592 262954
rect 189540 262890 189592 262896
rect 189448 260024 189500 260030
rect 189448 259966 189500 259972
rect 189356 143200 189408 143206
rect 189356 143142 189408 143148
rect 189460 141778 189488 259966
rect 189552 145450 189580 262890
rect 190460 262336 190512 262342
rect 190460 262278 190512 262284
rect 189632 260296 189684 260302
rect 189632 260238 189684 260244
rect 189644 145518 189672 260238
rect 189722 260128 189778 260137
rect 189722 260063 189778 260072
rect 189736 156534 189764 260063
rect 190472 199442 190500 262278
rect 190920 260976 190972 260982
rect 190920 260918 190972 260924
rect 190736 260432 190788 260438
rect 190736 260374 190788 260380
rect 190460 199436 190512 199442
rect 190460 199378 190512 199384
rect 190000 199232 190052 199238
rect 190000 199174 190052 199180
rect 189908 165640 189960 165646
rect 189908 165582 189960 165588
rect 189724 156528 189776 156534
rect 189724 156470 189776 156476
rect 189724 146736 189776 146742
rect 189724 146678 189776 146684
rect 189632 145512 189684 145518
rect 189632 145454 189684 145460
rect 189540 145444 189592 145450
rect 189540 145386 189592 145392
rect 189448 141772 189500 141778
rect 189448 141714 189500 141720
rect 189632 141160 189684 141166
rect 189632 141102 189684 141108
rect 189356 140412 189408 140418
rect 189356 140354 189408 140360
rect 189092 66694 189304 66722
rect 189092 66094 189120 66694
rect 189080 66088 189132 66094
rect 189080 66030 189132 66036
rect 189092 65686 189120 66030
rect 189080 65680 189132 65686
rect 189080 65622 189132 65628
rect 189080 63436 189132 63442
rect 189080 63378 189132 63384
rect 189092 62898 189120 63378
rect 189080 62892 189132 62898
rect 189080 62834 189132 62840
rect 189080 60580 189132 60586
rect 189080 60522 189132 60528
rect 189092 60246 189120 60522
rect 189080 60240 189132 60246
rect 189080 60182 189132 60188
rect 189368 55214 189396 140354
rect 189448 140004 189500 140010
rect 189448 139946 189500 139952
rect 189460 67590 189488 139946
rect 189538 81832 189594 81841
rect 189538 81767 189594 81776
rect 189552 79665 189580 81767
rect 189538 79656 189594 79665
rect 189538 79591 189594 79600
rect 189644 69766 189672 141102
rect 189736 80345 189764 146678
rect 189816 144424 189868 144430
rect 189816 144366 189868 144372
rect 189828 81977 189856 144366
rect 189920 144090 189948 165582
rect 189908 144084 189960 144090
rect 189908 144026 189960 144032
rect 189908 140072 189960 140078
rect 189908 140014 189960 140020
rect 189814 81968 189870 81977
rect 189814 81903 189870 81912
rect 189920 80578 189948 140014
rect 189908 80572 189960 80578
rect 189908 80514 189960 80520
rect 189722 80336 189778 80345
rect 189722 80271 189778 80280
rect 189632 69760 189684 69766
rect 189632 69702 189684 69708
rect 189724 68332 189776 68338
rect 189724 68274 189776 68280
rect 189448 67584 189500 67590
rect 189448 67526 189500 67532
rect 189356 55208 189408 55214
rect 189356 55150 189408 55156
rect 189368 54534 189396 55150
rect 189356 54528 189408 54534
rect 189356 54470 189408 54476
rect 188804 40996 188856 41002
rect 188804 40938 188856 40944
rect 189736 16574 189764 68274
rect 190012 62898 190040 199174
rect 190644 196648 190696 196654
rect 190644 196590 190696 196596
rect 190458 195528 190514 195537
rect 190458 195463 190514 195472
rect 190092 195220 190144 195226
rect 190092 195162 190144 195168
rect 190000 62892 190052 62898
rect 190000 62834 190052 62840
rect 190104 60246 190132 195162
rect 190092 60240 190144 60246
rect 190092 60182 190144 60188
rect 190472 44033 190500 195463
rect 190552 195424 190604 195430
rect 190552 195366 190604 195372
rect 190564 61946 190592 195366
rect 190656 64802 190684 196590
rect 190748 141710 190776 260374
rect 190828 260092 190880 260098
rect 190828 260034 190880 260040
rect 190840 143138 190868 260034
rect 190932 145586 190960 260918
rect 191012 260908 191064 260914
rect 191012 260850 191064 260856
rect 191024 146266 191052 260850
rect 191932 200592 191984 200598
rect 191932 200534 191984 200540
rect 191840 200252 191892 200258
rect 191840 200194 191892 200200
rect 191104 192364 191156 192370
rect 191104 192306 191156 192312
rect 191012 146260 191064 146266
rect 191012 146202 191064 146208
rect 190920 145580 190972 145586
rect 190920 145522 190972 145528
rect 190828 143132 190880 143138
rect 190828 143074 190880 143080
rect 191012 142180 191064 142186
rect 191012 142122 191064 142128
rect 190736 141704 190788 141710
rect 190736 141646 190788 141652
rect 190736 140276 190788 140282
rect 190736 140218 190788 140224
rect 190644 64796 190696 64802
rect 190644 64738 190696 64744
rect 190552 61940 190604 61946
rect 190552 61882 190604 61888
rect 190748 52193 190776 140218
rect 190826 78296 190882 78305
rect 190826 78231 190882 78240
rect 190840 76906 190868 78231
rect 190828 76900 190880 76906
rect 190828 76842 190880 76848
rect 191024 71262 191052 142122
rect 191116 79286 191144 192306
rect 191380 147280 191432 147286
rect 191380 147222 191432 147228
rect 191288 143404 191340 143410
rect 191288 143346 191340 143352
rect 191194 136640 191250 136649
rect 191194 136575 191250 136584
rect 191104 79280 191156 79286
rect 191104 79222 191156 79228
rect 191208 72962 191236 136575
rect 191300 82113 191328 143346
rect 191286 82104 191342 82113
rect 191286 82039 191342 82048
rect 191196 72956 191248 72962
rect 191196 72898 191248 72904
rect 191012 71256 191064 71262
rect 191012 71198 191064 71204
rect 191392 69902 191420 147222
rect 191472 146804 191524 146810
rect 191472 146746 191524 146752
rect 191484 74534 191512 146746
rect 191484 74506 191696 74534
rect 191668 72758 191696 74506
rect 191748 72956 191800 72962
rect 191748 72898 191800 72904
rect 191760 72826 191788 72898
rect 191748 72820 191800 72826
rect 191748 72762 191800 72768
rect 191656 72752 191708 72758
rect 191656 72694 191708 72700
rect 191668 72486 191696 72694
rect 191656 72480 191708 72486
rect 191656 72422 191708 72428
rect 191380 69896 191432 69902
rect 191380 69838 191432 69844
rect 191852 64874 191880 200194
rect 191944 65958 191972 200534
rect 192036 143274 192064 265610
rect 192116 265600 192168 265606
rect 192116 265542 192168 265548
rect 192128 144770 192156 265542
rect 199200 265532 199252 265538
rect 199200 265474 199252 265480
rect 195060 265464 195112 265470
rect 195060 265406 195112 265412
rect 193588 265328 193640 265334
rect 193588 265270 193640 265276
rect 193128 263492 193180 263498
rect 193128 263434 193180 263440
rect 192300 263084 192352 263090
rect 192300 263026 192352 263032
rect 192208 195968 192260 195974
rect 192208 195910 192260 195916
rect 192116 144764 192168 144770
rect 192116 144706 192168 144712
rect 192024 143268 192076 143274
rect 192024 143210 192076 143216
rect 192220 75546 192248 195910
rect 192312 144702 192340 263026
rect 192666 262848 192722 262857
rect 192392 262812 192444 262818
rect 192666 262783 192722 262792
rect 192392 262754 192444 262760
rect 192404 157282 192432 262754
rect 192484 262608 192536 262614
rect 192484 262550 192536 262556
rect 192496 262313 192524 262550
rect 192482 262304 192538 262313
rect 192482 262239 192538 262248
rect 192680 193905 192708 262783
rect 193140 262614 193168 263434
rect 193128 262608 193180 262614
rect 193128 262550 193180 262556
rect 193496 262472 193548 262478
rect 193496 262414 193548 262420
rect 193220 200524 193272 200530
rect 193220 200466 193272 200472
rect 192666 193896 192722 193905
rect 192666 193831 192722 193840
rect 192392 157276 192444 157282
rect 192392 157218 192444 157224
rect 192760 150408 192812 150414
rect 192760 150350 192812 150356
rect 192666 147248 192722 147257
rect 192666 147183 192722 147192
rect 192392 147144 192444 147150
rect 192392 147086 192444 147092
rect 192300 144696 192352 144702
rect 192300 144638 192352 144644
rect 192300 141364 192352 141370
rect 192300 141306 192352 141312
rect 192208 75540 192260 75546
rect 192208 75482 192260 75488
rect 192312 72622 192340 141306
rect 192404 76838 192432 147086
rect 192484 140548 192536 140554
rect 192484 140490 192536 140496
rect 192392 76832 192444 76838
rect 192392 76774 192444 76780
rect 192300 72616 192352 72622
rect 192300 72558 192352 72564
rect 192496 71398 192524 140490
rect 192574 139360 192630 139369
rect 192574 139295 192630 139304
rect 192588 71534 192616 139295
rect 192680 79490 192708 147183
rect 192668 79484 192720 79490
rect 192668 79426 192720 79432
rect 192772 72690 192800 150350
rect 192852 147348 192904 147354
rect 192852 147290 192904 147296
rect 192864 76430 192892 147290
rect 193126 76528 193182 76537
rect 193126 76463 193182 76472
rect 192852 76424 192904 76430
rect 192852 76366 192904 76372
rect 192760 72684 192812 72690
rect 192760 72626 192812 72632
rect 192576 71528 192628 71534
rect 192576 71470 192628 71476
rect 192484 71392 192536 71398
rect 192484 71334 192536 71340
rect 191932 65952 191984 65958
rect 191932 65894 191984 65900
rect 193036 65952 193088 65958
rect 193036 65894 193088 65900
rect 193048 65618 193076 65894
rect 193036 65612 193088 65618
rect 193036 65554 193088 65560
rect 191852 64846 191972 64874
rect 191748 64796 191800 64802
rect 191748 64738 191800 64744
rect 191760 64258 191788 64738
rect 191748 64252 191800 64258
rect 191748 64194 191800 64200
rect 191748 61940 191800 61946
rect 191748 61882 191800 61888
rect 191760 61470 191788 61882
rect 191748 61464 191800 61470
rect 191748 61406 191800 61412
rect 191944 59362 191972 64846
rect 191932 59356 191984 59362
rect 191932 59298 191984 59304
rect 193036 59356 193088 59362
rect 193036 59298 193088 59304
rect 193048 58682 193076 59298
rect 193036 58676 193088 58682
rect 193036 58618 193088 58624
rect 190734 52184 190790 52193
rect 190734 52119 190790 52128
rect 191838 46200 191894 46209
rect 191838 46135 191894 46144
rect 190458 44024 190514 44033
rect 190458 43959 190514 43968
rect 191746 44024 191802 44033
rect 191746 43959 191802 43968
rect 191760 43761 191788 43959
rect 191746 43752 191802 43761
rect 191746 43687 191802 43696
rect 191852 16574 191880 46135
rect 189736 16546 189948 16574
rect 191852 16546 192064 16574
rect 188344 4140 188396 4146
rect 188344 4082 188396 4088
rect 189816 4072 189868 4078
rect 189816 4014 189868 4020
rect 188264 3454 188568 3482
rect 188540 480 188568 3454
rect 189828 3398 189856 4014
rect 189724 3392 189776 3398
rect 189724 3334 189776 3340
rect 189816 3392 189868 3398
rect 189816 3334 189868 3340
rect 189736 480 189764 3334
rect 189920 3330 189948 16546
rect 190828 3392 190880 3398
rect 190828 3334 190880 3340
rect 189908 3324 189960 3330
rect 189908 3266 189960 3272
rect 190840 480 190868 3334
rect 192036 480 192064 16546
rect 193140 3398 193168 76463
rect 193232 57905 193260 200466
rect 193404 197260 193456 197266
rect 193404 197202 193456 197208
rect 193312 195560 193364 195566
rect 193312 195502 193364 195508
rect 193218 57896 193274 57905
rect 193218 57831 193274 57840
rect 193324 52329 193352 195502
rect 193416 74534 193444 197202
rect 193508 141914 193536 262414
rect 193600 144566 193628 265270
rect 194968 265124 195020 265130
rect 194968 265066 195020 265072
rect 193772 262744 193824 262750
rect 193772 262686 193824 262692
rect 193680 259956 193732 259962
rect 193680 259898 193732 259904
rect 193692 144634 193720 259898
rect 193784 157214 193812 262686
rect 194876 197192 194928 197198
rect 194876 197134 194928 197140
rect 194600 197124 194652 197130
rect 194600 197066 194652 197072
rect 193772 157208 193824 157214
rect 193772 157150 193824 157156
rect 193770 149696 193826 149705
rect 193770 149631 193826 149640
rect 193680 144628 193732 144634
rect 193680 144570 193732 144576
rect 193588 144560 193640 144566
rect 193588 144502 193640 144508
rect 193496 141908 193548 141914
rect 193496 141850 193548 141856
rect 193496 140752 193548 140758
rect 193494 140720 193496 140729
rect 193548 140720 193550 140729
rect 193494 140655 193550 140664
rect 193416 74506 193536 74534
rect 193402 67552 193458 67561
rect 193402 67487 193458 67496
rect 193416 67046 193444 67487
rect 193404 67040 193456 67046
rect 193404 66982 193456 66988
rect 193508 60722 193536 74506
rect 193784 74050 193812 149631
rect 194140 147552 194192 147558
rect 194140 147494 194192 147500
rect 193864 147212 193916 147218
rect 193864 147154 193916 147160
rect 193876 79082 193904 147154
rect 193954 139088 194010 139097
rect 193954 139023 194010 139032
rect 193864 79076 193916 79082
rect 193864 79018 193916 79024
rect 193864 75268 193916 75274
rect 193864 75210 193916 75216
rect 193772 74044 193824 74050
rect 193772 73986 193824 73992
rect 193784 73846 193812 73986
rect 193772 73840 193824 73846
rect 193772 73782 193824 73788
rect 193496 60716 193548 60722
rect 193496 60658 193548 60664
rect 193310 52320 193366 52329
rect 193310 52255 193366 52264
rect 193310 50280 193366 50289
rect 193310 50215 193366 50224
rect 193324 16574 193352 50215
rect 193324 16546 193812 16574
rect 193784 3482 193812 16546
rect 193876 4078 193904 75210
rect 193968 71602 193996 139023
rect 194046 135960 194102 135969
rect 194046 135895 194102 135904
rect 194060 79354 194088 135895
rect 194048 79348 194100 79354
rect 194048 79290 194100 79296
rect 194152 72554 194180 147494
rect 194232 145376 194284 145382
rect 194232 145318 194284 145324
rect 194140 72548 194192 72554
rect 194140 72490 194192 72496
rect 194244 72282 194272 145318
rect 194322 144664 194378 144673
rect 194322 144599 194378 144608
rect 194232 72276 194284 72282
rect 194232 72218 194284 72224
rect 193956 71596 194008 71602
rect 193956 71538 194008 71544
rect 194336 53786 194364 144599
rect 194508 67040 194560 67046
rect 194508 66982 194560 66988
rect 194520 66434 194548 66982
rect 194508 66428 194560 66434
rect 194508 66370 194560 66376
rect 194508 60716 194560 60722
rect 194508 60658 194560 60664
rect 194520 60178 194548 60658
rect 194508 60172 194560 60178
rect 194508 60114 194560 60120
rect 194324 53780 194376 53786
rect 194324 53722 194376 53728
rect 194336 53106 194364 53722
rect 194612 53689 194640 197066
rect 194782 195392 194838 195401
rect 194782 195327 194838 195336
rect 194690 192944 194746 192953
rect 194690 192879 194746 192888
rect 194598 53680 194654 53689
rect 194598 53615 194654 53624
rect 194324 53100 194376 53106
rect 194324 53042 194376 53048
rect 194506 52320 194562 52329
rect 194506 52255 194562 52264
rect 194520 52057 194548 52255
rect 194506 52048 194562 52057
rect 194506 51983 194562 51992
rect 194704 50425 194732 192879
rect 194796 54913 194824 195327
rect 194888 64569 194916 197134
rect 194980 144498 195008 265066
rect 195072 145994 195100 265406
rect 196624 265396 196676 265402
rect 196624 265338 196676 265344
rect 196256 265192 196308 265198
rect 196256 265134 196308 265140
rect 195152 262676 195204 262682
rect 195152 262618 195204 262624
rect 195164 159662 195192 262618
rect 196164 199028 196216 199034
rect 196164 198970 196216 198976
rect 196070 197024 196126 197033
rect 196070 196959 196126 196968
rect 195978 196888 196034 196897
rect 195978 196823 196034 196832
rect 195152 159656 195204 159662
rect 195152 159598 195204 159604
rect 195152 150204 195204 150210
rect 195152 150146 195204 150152
rect 195060 145988 195112 145994
rect 195060 145930 195112 145936
rect 194968 144492 195020 144498
rect 194968 144434 195020 144440
rect 195060 144152 195112 144158
rect 195060 144094 195112 144100
rect 195072 68406 195100 144094
rect 195164 78062 195192 150146
rect 195520 149728 195572 149734
rect 195520 149670 195572 149676
rect 195244 147076 195296 147082
rect 195244 147018 195296 147024
rect 195152 78056 195204 78062
rect 195152 77998 195204 78004
rect 195256 76634 195284 147018
rect 195336 142112 195388 142118
rect 195336 142054 195388 142060
rect 195348 77042 195376 142054
rect 195426 137864 195482 137873
rect 195426 137799 195482 137808
rect 195440 82249 195468 137799
rect 195426 82240 195482 82249
rect 195426 82175 195482 82184
rect 195336 77036 195388 77042
rect 195336 76978 195388 76984
rect 195244 76628 195296 76634
rect 195244 76570 195296 76576
rect 195348 76566 195376 76978
rect 195336 76560 195388 76566
rect 195336 76502 195388 76508
rect 195060 68400 195112 68406
rect 195060 68342 195112 68348
rect 195532 67522 195560 149670
rect 195520 67516 195572 67522
rect 195520 67458 195572 67464
rect 194874 64560 194930 64569
rect 194874 64495 194930 64504
rect 194888 64297 194916 64495
rect 194874 64288 194930 64297
rect 194874 64223 194930 64232
rect 194782 54904 194838 54913
rect 194782 54839 194838 54848
rect 194690 50416 194746 50425
rect 194690 50351 194746 50360
rect 195992 49473 196020 196823
rect 196084 56409 196112 196959
rect 196176 74534 196204 198970
rect 196268 141506 196296 265134
rect 196440 265056 196492 265062
rect 196440 264998 196492 265004
rect 196348 200184 196400 200190
rect 196348 200126 196400 200132
rect 196256 141500 196308 141506
rect 196256 141442 196308 141448
rect 196360 79014 196388 200126
rect 196452 145926 196480 264998
rect 196532 259480 196584 259486
rect 196532 259422 196584 259428
rect 196440 145920 196492 145926
rect 196440 145862 196492 145868
rect 196544 143070 196572 259422
rect 196636 159730 196664 265338
rect 197912 263628 197964 263634
rect 197912 263570 197964 263576
rect 197820 261044 197872 261050
rect 197820 260986 197872 260992
rect 197358 197160 197414 197169
rect 197358 197095 197414 197104
rect 196624 159724 196676 159730
rect 196624 159666 196676 159672
rect 196716 150340 196768 150346
rect 196716 150282 196768 150288
rect 196532 143064 196584 143070
rect 196532 143006 196584 143012
rect 196622 138952 196678 138961
rect 196622 138887 196678 138896
rect 196348 79008 196400 79014
rect 196348 78950 196400 78956
rect 196176 74506 196296 74534
rect 196162 66192 196218 66201
rect 196162 66127 196218 66136
rect 196176 65890 196204 66127
rect 196164 65884 196216 65890
rect 196164 65826 196216 65832
rect 196176 64938 196204 65826
rect 196164 64932 196216 64938
rect 196164 64874 196216 64880
rect 196268 59129 196296 74506
rect 196636 70310 196664 138887
rect 196728 81841 196756 150282
rect 196992 147620 197044 147626
rect 196992 147562 197044 147568
rect 196808 140208 196860 140214
rect 196808 140150 196860 140156
rect 196714 81832 196770 81841
rect 196714 81767 196770 81776
rect 196820 79150 196848 140150
rect 196898 81560 196954 81569
rect 196898 81495 196954 81504
rect 196808 79144 196860 79150
rect 196808 79086 196860 79092
rect 196912 73778 196940 81495
rect 196900 73772 196952 73778
rect 196900 73714 196952 73720
rect 196624 70304 196676 70310
rect 196624 70246 196676 70252
rect 197004 67250 197032 147562
rect 197176 147008 197228 147014
rect 197176 146950 197228 146956
rect 197084 145784 197136 145790
rect 197084 145726 197136 145732
rect 197096 71466 197124 145726
rect 197084 71460 197136 71466
rect 197084 71402 197136 71408
rect 197188 70174 197216 146950
rect 197176 70168 197228 70174
rect 197176 70110 197228 70116
rect 197268 69488 197320 69494
rect 197268 69430 197320 69436
rect 196992 67244 197044 67250
rect 196992 67186 197044 67192
rect 196254 59120 196310 59129
rect 196254 59055 196310 59064
rect 196070 56400 196126 56409
rect 196070 56335 196126 56344
rect 196084 56137 196112 56335
rect 196070 56128 196126 56137
rect 196070 56063 196126 56072
rect 195978 49464 196034 49473
rect 195978 49399 196034 49408
rect 196438 49464 196494 49473
rect 196438 49399 196494 49408
rect 196452 49201 196480 49399
rect 196438 49192 196494 49201
rect 196438 49127 196494 49136
rect 197280 4146 197308 69430
rect 197372 44169 197400 197095
rect 197636 196784 197688 196790
rect 197636 196726 197688 196732
rect 197542 196616 197598 196625
rect 197542 196551 197598 196560
rect 197452 61396 197504 61402
rect 197452 61338 197504 61344
rect 197358 44160 197414 44169
rect 197358 44095 197414 44104
rect 197372 43625 197400 44095
rect 197358 43616 197414 43625
rect 197358 43551 197414 43560
rect 197464 16574 197492 61338
rect 197556 48113 197584 196551
rect 197648 52465 197676 196726
rect 197728 196716 197780 196722
rect 197728 196658 197780 196664
rect 197740 62082 197768 196658
rect 197832 143342 197860 260986
rect 197924 146062 197952 263570
rect 198004 261384 198056 261390
rect 198004 261326 198056 261332
rect 198016 146130 198044 261326
rect 199016 261248 199068 261254
rect 199016 261190 199068 261196
rect 198096 261180 198148 261186
rect 198096 261122 198148 261128
rect 198108 149598 198136 261122
rect 198370 200560 198426 200569
rect 198370 200495 198426 200504
rect 198188 195900 198240 195906
rect 198188 195842 198240 195848
rect 198096 149592 198148 149598
rect 198096 149534 198148 149540
rect 198200 149161 198228 195842
rect 198280 150068 198332 150074
rect 198280 150010 198332 150016
rect 198186 149152 198242 149161
rect 198186 149087 198242 149096
rect 198004 146124 198056 146130
rect 198004 146066 198056 146072
rect 197912 146056 197964 146062
rect 197912 145998 197964 146004
rect 197912 145716 197964 145722
rect 197912 145658 197964 145664
rect 197820 143336 197872 143342
rect 197820 143278 197872 143284
rect 197924 78130 197952 145658
rect 198188 144832 198240 144838
rect 198188 144774 198240 144780
rect 198004 138712 198056 138718
rect 198004 138654 198056 138660
rect 197912 78124 197964 78130
rect 197912 78066 197964 78072
rect 198016 73098 198044 138654
rect 198200 80918 198228 144774
rect 198188 80912 198240 80918
rect 198188 80854 198240 80860
rect 198004 73092 198056 73098
rect 198004 73034 198056 73040
rect 198016 72486 198044 73034
rect 198004 72480 198056 72486
rect 198004 72422 198056 72428
rect 198292 70242 198320 150010
rect 198280 70236 198332 70242
rect 198280 70178 198332 70184
rect 197728 62076 197780 62082
rect 197728 62018 197780 62024
rect 198188 62076 198240 62082
rect 198188 62018 198240 62024
rect 198200 61402 198228 62018
rect 198188 61396 198240 61402
rect 198188 61338 198240 61344
rect 197728 60648 197780 60654
rect 197728 60590 197780 60596
rect 197740 60110 197768 60590
rect 197820 60512 197872 60518
rect 197820 60454 197872 60460
rect 197728 60104 197780 60110
rect 197728 60046 197780 60052
rect 197832 60042 197860 60454
rect 198384 60110 198412 200495
rect 198740 199300 198792 199306
rect 198740 199242 198792 199248
rect 198464 149932 198516 149938
rect 198464 149874 198516 149880
rect 198372 60104 198424 60110
rect 198372 60046 198424 60052
rect 198476 60042 198504 149874
rect 198752 63510 198780 199242
rect 198832 197056 198884 197062
rect 198832 196998 198884 197004
rect 198740 63504 198792 63510
rect 198740 63446 198792 63452
rect 198752 62830 198780 63446
rect 198740 62824 198792 62830
rect 198740 62766 198792 62772
rect 198740 60376 198792 60382
rect 198740 60318 198792 60324
rect 197820 60036 197872 60042
rect 197820 59978 197872 59984
rect 198464 60036 198516 60042
rect 198464 59978 198516 59984
rect 198004 57792 198056 57798
rect 198004 57734 198056 57740
rect 198016 57633 198044 57734
rect 198002 57624 198058 57633
rect 198002 57559 198058 57568
rect 198016 56642 198044 57559
rect 198004 56636 198056 56642
rect 198004 56578 198056 56584
rect 197634 52456 197690 52465
rect 197634 52391 197690 52400
rect 198278 52456 198334 52465
rect 198278 52391 198334 52400
rect 198292 51921 198320 52391
rect 198278 51912 198334 51921
rect 198278 51847 198334 51856
rect 197542 48104 197598 48113
rect 197542 48039 197598 48048
rect 197556 47841 197584 48039
rect 197542 47832 197598 47841
rect 197542 47767 197598 47776
rect 197464 16546 197952 16574
rect 196808 4140 196860 4146
rect 196808 4082 196860 4088
rect 197268 4140 197320 4146
rect 197268 4082 197320 4088
rect 193864 4072 193916 4078
rect 193864 4014 193916 4020
rect 195612 4072 195664 4078
rect 195612 4014 195664 4020
rect 195704 4072 195756 4078
rect 195704 4014 195756 4020
rect 193784 3454 194456 3482
rect 193128 3392 193180 3398
rect 193128 3334 193180 3340
rect 193220 3324 193272 3330
rect 193220 3266 193272 3272
rect 193232 480 193260 3266
rect 194428 480 194456 3454
rect 195624 480 195652 4014
rect 195716 3398 195744 4014
rect 195704 3392 195756 3398
rect 195704 3334 195756 3340
rect 196820 480 196848 4082
rect 197924 480 197952 16546
rect 181414 354 181526 480
rect 180996 326 181526 354
rect 181414 -960 181526 326
rect 182518 -960 182630 480
rect 183714 -960 183826 480
rect 184910 -960 185022 480
rect 186106 -960 186218 480
rect 187302 -960 187414 480
rect 188498 -960 188610 480
rect 189694 -960 189806 480
rect 190798 -960 190910 480
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195582 -960 195694 480
rect 196778 -960 196890 480
rect 197882 -960 197994 480
rect 198752 354 198780 60318
rect 198844 57769 198872 196998
rect 198924 196988 198976 196994
rect 198924 196930 198976 196936
rect 198936 66026 198964 196930
rect 199028 143313 199056 261190
rect 199108 261112 199160 261118
rect 199108 261054 199160 261060
rect 199120 146198 199148 261054
rect 199212 159798 199240 265474
rect 200580 262540 200632 262546
rect 200580 262482 200632 262488
rect 200394 200288 200450 200297
rect 200394 200223 200450 200232
rect 200304 199164 200356 199170
rect 200304 199106 200356 199112
rect 200210 196752 200266 196761
rect 200210 196687 200266 196696
rect 200120 191072 200172 191078
rect 200120 191014 200172 191020
rect 199200 159792 199252 159798
rect 199200 159734 199252 159740
rect 199200 154080 199252 154086
rect 199200 154022 199252 154028
rect 199108 146192 199160 146198
rect 199108 146134 199160 146140
rect 199014 143304 199070 143313
rect 199014 143239 199070 143248
rect 199016 78260 199068 78266
rect 199016 78202 199068 78208
rect 199028 78130 199056 78202
rect 199016 78124 199068 78130
rect 199016 78066 199068 78072
rect 199212 71330 199240 154022
rect 199752 150000 199804 150006
rect 199752 149942 199804 149948
rect 199476 149796 199528 149802
rect 199476 149738 199528 149744
rect 199292 148776 199344 148782
rect 199292 148718 199344 148724
rect 199304 76498 199332 148718
rect 199382 138816 199438 138825
rect 199382 138751 199438 138760
rect 199292 76492 199344 76498
rect 199292 76434 199344 76440
rect 199200 71324 199252 71330
rect 199200 71266 199252 71272
rect 199396 68202 199424 138751
rect 199488 80986 199516 149738
rect 199658 147656 199714 147665
rect 199658 147591 199714 147600
rect 199568 144900 199620 144906
rect 199568 144842 199620 144848
rect 199476 80980 199528 80986
rect 199476 80922 199528 80928
rect 199580 78130 199608 144842
rect 199568 78124 199620 78130
rect 199568 78066 199620 78072
rect 199384 68196 199436 68202
rect 199384 68138 199436 68144
rect 199200 67108 199252 67114
rect 199200 67050 199252 67056
rect 199212 66473 199240 67050
rect 199198 66464 199254 66473
rect 199198 66399 199254 66408
rect 199212 66366 199240 66399
rect 199200 66360 199252 66366
rect 199200 66302 199252 66308
rect 198924 66020 198976 66026
rect 198924 65962 198976 65968
rect 198936 65550 198964 65962
rect 198924 65544 198976 65550
rect 198924 65486 198976 65492
rect 199672 64870 199700 147591
rect 199764 69970 199792 149942
rect 199752 69964 199804 69970
rect 199752 69906 199804 69912
rect 199660 64864 199712 64870
rect 198922 64832 198978 64841
rect 199660 64806 199712 64812
rect 198922 64767 198978 64776
rect 198936 64598 198964 64767
rect 200132 64734 200160 191014
rect 200120 64728 200172 64734
rect 200120 64670 200172 64676
rect 198924 64592 198976 64598
rect 198924 64534 198976 64540
rect 198936 63578 198964 64534
rect 198924 63572 198976 63578
rect 198924 63514 198976 63520
rect 198830 57760 198886 57769
rect 198830 57695 198886 57704
rect 200224 45393 200252 196687
rect 200316 53825 200344 199106
rect 200408 55049 200436 200223
rect 200488 196852 200540 196858
rect 200488 196794 200540 196800
rect 200500 69737 200528 196794
rect 200592 156738 200620 262482
rect 201866 259584 201922 259593
rect 201866 259519 201922 259528
rect 201592 198620 201644 198626
rect 201592 198562 201644 198568
rect 201040 195764 201092 195770
rect 201040 195706 201092 195712
rect 200580 156732 200632 156738
rect 200580 156674 200632 156680
rect 200948 156664 201000 156670
rect 200948 156606 201000 156612
rect 200580 154012 200632 154018
rect 200580 153954 200632 153960
rect 200486 69728 200542 69737
rect 200486 69663 200542 69672
rect 200592 68474 200620 153954
rect 200672 153944 200724 153950
rect 200672 153886 200724 153892
rect 200684 68678 200712 153886
rect 200856 150136 200908 150142
rect 200856 150078 200908 150084
rect 200764 149864 200816 149870
rect 200764 149806 200816 149812
rect 200776 68746 200804 149806
rect 200868 71641 200896 150078
rect 200960 77994 200988 156606
rect 201052 149161 201080 195706
rect 201500 191820 201552 191826
rect 201500 191762 201552 191768
rect 201038 149152 201094 149161
rect 201038 149087 201094 149096
rect 201038 80064 201094 80073
rect 201038 79999 201094 80008
rect 201052 78742 201080 79999
rect 201040 78736 201092 78742
rect 201040 78678 201092 78684
rect 200948 77988 201000 77994
rect 200948 77930 201000 77936
rect 201512 76362 201540 191762
rect 201500 76356 201552 76362
rect 201500 76298 201552 76304
rect 201500 75200 201552 75206
rect 201500 75142 201552 75148
rect 200854 71632 200910 71641
rect 200854 71567 200910 71576
rect 200856 71052 200908 71058
rect 200856 70994 200908 71000
rect 200764 68740 200816 68746
rect 200764 68682 200816 68688
rect 200672 68672 200724 68678
rect 200672 68614 200724 68620
rect 200580 68468 200632 68474
rect 200580 68410 200632 68416
rect 200394 55040 200450 55049
rect 200394 54975 200450 54984
rect 200302 53816 200358 53825
rect 200302 53751 200358 53760
rect 200210 45384 200266 45393
rect 200210 45319 200266 45328
rect 200868 6914 200896 70994
rect 201406 55040 201462 55049
rect 201406 54975 201462 54984
rect 201420 54777 201448 54975
rect 201406 54768 201462 54777
rect 201406 54703 201462 54712
rect 201406 53816 201462 53825
rect 201406 53751 201462 53760
rect 201420 53281 201448 53751
rect 201406 53272 201462 53281
rect 201406 53207 201462 53216
rect 201512 11694 201540 75142
rect 201604 56001 201632 198562
rect 201684 196920 201736 196926
rect 201684 196862 201736 196868
rect 201696 69766 201724 196862
rect 201776 191752 201828 191758
rect 201776 191694 201828 191700
rect 201684 69760 201736 69766
rect 201684 69702 201736 69708
rect 201682 67552 201738 67561
rect 201682 67487 201738 67496
rect 201696 67182 201724 67487
rect 201684 67176 201736 67182
rect 201684 67118 201736 67124
rect 201788 63345 201816 191694
rect 201880 156806 201908 259519
rect 202512 198688 202564 198694
rect 202512 198630 202564 198636
rect 201960 157004 202012 157010
rect 201960 156946 202012 156952
rect 201868 156800 201920 156806
rect 201868 156742 201920 156748
rect 201868 69760 201920 69766
rect 201868 69702 201920 69708
rect 201774 63336 201830 63345
rect 201774 63271 201830 63280
rect 201880 58721 201908 69702
rect 201972 68814 202000 156946
rect 202418 156904 202474 156913
rect 202144 156868 202196 156874
rect 202418 156839 202474 156848
rect 202144 156810 202196 156816
rect 202052 153876 202104 153882
rect 202052 153818 202104 153824
rect 202064 68882 202092 153818
rect 202156 78470 202184 156810
rect 202236 148640 202288 148646
rect 202236 148582 202288 148588
rect 202248 81025 202276 148582
rect 202328 140140 202380 140146
rect 202328 140082 202380 140088
rect 202234 81016 202290 81025
rect 202234 80951 202290 80960
rect 202340 79558 202368 140082
rect 202328 79552 202380 79558
rect 202328 79494 202380 79500
rect 202144 78464 202196 78470
rect 202144 78406 202196 78412
rect 202052 68876 202104 68882
rect 202052 68818 202104 68824
rect 201960 68808 202012 68814
rect 201960 68750 202012 68756
rect 202142 62112 202198 62121
rect 202142 62047 202198 62056
rect 202156 61878 202184 62047
rect 202144 61872 202196 61878
rect 202144 61814 202196 61820
rect 202432 61577 202460 156839
rect 202524 139505 202552 198630
rect 202880 194540 202932 194546
rect 202880 194482 202932 194488
rect 202510 139496 202566 139505
rect 202510 139431 202566 139440
rect 202788 67176 202840 67182
rect 202788 67118 202840 67124
rect 202800 66298 202828 67118
rect 202788 66292 202840 66298
rect 202788 66234 202840 66240
rect 202786 63336 202842 63345
rect 202786 63271 202842 63280
rect 202800 62801 202828 63271
rect 202786 62792 202842 62801
rect 202786 62727 202842 62736
rect 202788 61872 202840 61878
rect 202788 61814 202840 61820
rect 202418 61568 202474 61577
rect 202418 61503 202474 61512
rect 202800 60790 202828 61814
rect 202788 60784 202840 60790
rect 202788 60726 202840 60732
rect 201866 58712 201922 58721
rect 201866 58647 201922 58656
rect 201590 55992 201646 56001
rect 201590 55927 201646 55936
rect 201592 53236 201644 53242
rect 201592 53178 201644 53184
rect 201500 11688 201552 11694
rect 201500 11630 201552 11636
rect 201604 6914 201632 53178
rect 202892 52426 202920 194482
rect 202972 194472 203024 194478
rect 202972 194414 203024 194420
rect 202984 64666 203012 194414
rect 203076 152726 203104 276014
rect 204812 275324 204864 275330
rect 204812 275266 204864 275272
rect 204824 274718 204852 275266
rect 204536 274712 204588 274718
rect 204536 274654 204588 274660
rect 204812 274712 204864 274718
rect 204812 274654 204864 274660
rect 203432 259616 203484 259622
rect 203432 259558 203484 259564
rect 203156 199096 203208 199102
rect 203156 199038 203208 199044
rect 203064 152720 203116 152726
rect 203064 152662 203116 152668
rect 203168 78402 203196 199038
rect 203248 191684 203300 191690
rect 203248 191626 203300 191632
rect 203156 78396 203208 78402
rect 203156 78338 203208 78344
rect 203260 71194 203288 191626
rect 203340 187332 203392 187338
rect 203340 187274 203392 187280
rect 203352 78334 203380 187274
rect 203444 157350 203472 259558
rect 204444 193112 204496 193118
rect 204444 193054 204496 193060
rect 204352 191616 204404 191622
rect 204352 191558 204404 191564
rect 203432 157344 203484 157350
rect 203432 157286 203484 157292
rect 203800 157072 203852 157078
rect 203800 157014 203852 157020
rect 203432 156936 203484 156942
rect 203432 156878 203484 156884
rect 203340 78328 203392 78334
rect 203340 78270 203392 78276
rect 203248 71188 203300 71194
rect 203248 71130 203300 71136
rect 203444 70038 203472 156878
rect 203524 148572 203576 148578
rect 203524 148514 203576 148520
rect 203536 73001 203564 148514
rect 203708 148504 203760 148510
rect 203708 148446 203760 148452
rect 203614 148336 203670 148345
rect 203614 148271 203670 148280
rect 203628 74118 203656 148271
rect 203720 74186 203748 148446
rect 203708 74180 203760 74186
rect 203708 74122 203760 74128
rect 203616 74112 203668 74118
rect 203616 74054 203668 74060
rect 203522 72992 203578 73001
rect 203522 72927 203578 72936
rect 203432 70032 203484 70038
rect 203432 69974 203484 69980
rect 203812 68270 203840 157014
rect 204168 78396 204220 78402
rect 204168 78338 204220 78344
rect 204076 78328 204128 78334
rect 204076 78270 204128 78276
rect 204088 77994 204116 78270
rect 204180 78062 204208 78338
rect 204168 78056 204220 78062
rect 204168 77998 204220 78004
rect 204076 77988 204128 77994
rect 204076 77930 204128 77936
rect 203800 68264 203852 68270
rect 203800 68206 203852 68212
rect 204166 66872 204222 66881
rect 204166 66807 204222 66816
rect 204180 66094 204208 66807
rect 204364 66162 204392 191558
rect 204456 68610 204484 193054
rect 204548 152590 204576 274654
rect 218072 263498 218100 703582
rect 218808 703474 218836 703582
rect 218950 703520 219062 704960
rect 234632 703582 235028 703610
rect 218992 703474 219020 703520
rect 218808 703446 219020 703474
rect 234632 278089 234660 703582
rect 235000 703474 235028 703582
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 299492 703582 299980 703610
rect 235184 703474 235212 703520
rect 235000 703446 235212 703474
rect 267660 700670 267688 703520
rect 283852 702434 283880 703520
rect 282932 702406 283880 702434
rect 267648 700664 267700 700670
rect 267648 700606 267700 700612
rect 234618 278080 234674 278089
rect 234618 278015 234674 278024
rect 218060 263492 218112 263498
rect 218060 263434 218112 263440
rect 282932 263129 282960 702406
rect 299492 276690 299520 703582
rect 299952 703474 299980 703582
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 413622 703520 413734 704960
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494072 703582 494652 703610
rect 300136 703474 300164 703520
rect 299952 703446 300164 703474
rect 332520 700466 332548 703520
rect 348804 702434 348832 703520
rect 364996 702434 365024 703520
rect 347792 702406 348832 702434
rect 364352 702406 365024 702434
rect 332508 700460 332560 700466
rect 332508 700402 332560 700408
rect 299480 276684 299532 276690
rect 299480 276626 299532 276632
rect 282918 263120 282974 263129
rect 282918 263055 282974 263064
rect 347792 262993 347820 702406
rect 364352 275330 364380 702406
rect 397472 699718 397500 703520
rect 413664 700398 413692 703520
rect 413652 700392 413704 700398
rect 413652 700334 413704 700340
rect 429856 699718 429884 703520
rect 396724 699712 396776 699718
rect 396724 699654 396776 699660
rect 397460 699712 397512 699718
rect 397460 699654 397512 699660
rect 428464 699712 428516 699718
rect 428464 699654 428516 699660
rect 429844 699712 429896 699718
rect 429844 699654 429896 699660
rect 396736 284986 396764 699654
rect 396724 284980 396776 284986
rect 396724 284922 396776 284928
rect 364340 275324 364392 275330
rect 364340 275266 364392 275272
rect 428476 273970 428504 699654
rect 462332 660346 462360 703520
rect 478524 702434 478552 703520
rect 477512 702406 478552 702434
rect 462320 660340 462372 660346
rect 462320 660282 462372 660288
rect 428464 273964 428516 273970
rect 428464 273906 428516 273912
rect 347778 262984 347834 262993
rect 347778 262919 347834 262928
rect 477512 262857 477540 702406
rect 494072 271182 494100 703582
rect 494624 703474 494652 703582
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 494808 703474 494836 703520
rect 494624 703446 494836 703474
rect 527192 283626 527220 703520
rect 543476 700330 543504 703520
rect 559668 700330 559696 703520
rect 543464 700324 543516 700330
rect 543464 700266 543516 700272
rect 559656 700324 559708 700330
rect 559656 700266 559708 700272
rect 543004 700256 543056 700262
rect 543004 700198 543056 700204
rect 527180 283620 527232 283626
rect 527180 283562 527232 283568
rect 494060 271176 494112 271182
rect 494060 271118 494112 271124
rect 543016 269822 543044 700198
rect 580170 697232 580226 697241
rect 580170 697167 580226 697176
rect 580184 696998 580212 697167
rect 580172 696992 580224 696998
rect 580172 696934 580224 696940
rect 580170 683904 580226 683913
rect 580170 683839 580226 683848
rect 580184 683194 580212 683839
rect 580172 683188 580224 683194
rect 580172 683130 580224 683136
rect 580172 670744 580224 670750
rect 580170 670712 580172 670721
rect 580224 670712 580226 670721
rect 580170 670647 580226 670656
rect 580170 644056 580226 644065
rect 580170 643991 580226 644000
rect 580184 643142 580212 643991
rect 580172 643136 580224 643142
rect 580172 643078 580224 643084
rect 580170 630864 580226 630873
rect 580170 630799 580226 630808
rect 580184 630698 580212 630799
rect 580172 630692 580224 630698
rect 580172 630634 580224 630640
rect 580170 617536 580226 617545
rect 580170 617471 580226 617480
rect 580184 616894 580212 617471
rect 580172 616888 580224 616894
rect 580172 616830 580224 616836
rect 579802 591016 579858 591025
rect 579802 590951 579858 590960
rect 579816 590714 579844 590951
rect 579804 590708 579856 590714
rect 579804 590650 579856 590656
rect 580170 577688 580226 577697
rect 580170 577623 580226 577632
rect 580184 576910 580212 577623
rect 580172 576904 580224 576910
rect 580172 576846 580224 576852
rect 579802 564360 579858 564369
rect 579802 564295 579858 564304
rect 579816 563106 579844 564295
rect 579804 563100 579856 563106
rect 579804 563042 579856 563048
rect 580170 537840 580226 537849
rect 580170 537775 580226 537784
rect 580184 536858 580212 537775
rect 580172 536852 580224 536858
rect 580172 536794 580224 536800
rect 580170 524512 580226 524521
rect 580170 524447 580172 524456
rect 580224 524447 580226 524456
rect 580172 524418 580224 524424
rect 580170 511320 580226 511329
rect 580170 511255 580226 511264
rect 580184 510678 580212 511255
rect 580172 510672 580224 510678
rect 580172 510614 580224 510620
rect 580170 484664 580226 484673
rect 580170 484599 580226 484608
rect 580184 484430 580212 484599
rect 580172 484424 580224 484430
rect 580172 484366 580224 484372
rect 579986 471472 580042 471481
rect 579986 471407 580042 471416
rect 580000 470626 580028 471407
rect 579988 470620 580040 470626
rect 579988 470562 580040 470568
rect 580170 458144 580226 458153
rect 580170 458079 580226 458088
rect 580184 456822 580212 458079
rect 580172 456816 580224 456822
rect 580172 456758 580224 456764
rect 580170 431624 580226 431633
rect 580170 431559 580226 431568
rect 580184 430642 580212 431559
rect 580172 430636 580224 430642
rect 580172 430578 580224 430584
rect 580170 418296 580226 418305
rect 580170 418231 580226 418240
rect 580184 418198 580212 418231
rect 580172 418192 580224 418198
rect 580172 418134 580224 418140
rect 580170 404968 580226 404977
rect 580170 404903 580226 404912
rect 580184 404394 580212 404903
rect 580172 404388 580224 404394
rect 580172 404330 580224 404336
rect 580170 378448 580226 378457
rect 580170 378383 580226 378392
rect 580184 378214 580212 378383
rect 580172 378208 580224 378214
rect 580172 378150 580224 378156
rect 580262 365120 580318 365129
rect 580262 365055 580318 365064
rect 580172 351960 580224 351966
rect 580170 351928 580172 351937
rect 580224 351928 580226 351937
rect 580170 351863 580226 351872
rect 580170 325272 580226 325281
rect 580170 325207 580226 325216
rect 580184 324358 580212 325207
rect 580172 324352 580224 324358
rect 580172 324294 580224 324300
rect 579986 312080 580042 312089
rect 579986 312015 580042 312024
rect 580000 311914 580028 312015
rect 579988 311908 580040 311914
rect 579988 311850 580040 311856
rect 580170 298752 580226 298761
rect 580170 298687 580226 298696
rect 580184 298178 580212 298687
rect 580172 298172 580224 298178
rect 580172 298114 580224 298120
rect 580170 272232 580226 272241
rect 580170 272167 580226 272176
rect 580184 271930 580212 272167
rect 580172 271924 580224 271930
rect 580172 271866 580224 271872
rect 543004 269816 543056 269822
rect 543004 269758 543056 269764
rect 580276 263566 580304 365055
rect 580264 263560 580316 263566
rect 580264 263502 580316 263508
rect 580356 263016 580408 263022
rect 580356 262958 580408 262964
rect 477498 262848 477554 262857
rect 477498 262783 477554 262792
rect 471244 261316 471296 261322
rect 471244 261258 471296 261264
rect 206100 259548 206152 259554
rect 206100 259490 206152 259496
rect 204720 194132 204772 194138
rect 204720 194074 204772 194080
rect 204628 192908 204680 192914
rect 204628 192850 204680 192856
rect 204536 152584 204588 152590
rect 204536 152526 204588 152532
rect 204536 148708 204588 148714
rect 204536 148650 204588 148656
rect 204444 68604 204496 68610
rect 204444 68546 204496 68552
rect 204352 66156 204404 66162
rect 204352 66098 204404 66104
rect 204168 66088 204220 66094
rect 204168 66030 204220 66036
rect 202972 64660 203024 64666
rect 202972 64602 203024 64608
rect 202984 64190 203012 64602
rect 202972 64184 203024 64190
rect 202972 64126 203024 64132
rect 203248 57928 203300 57934
rect 203248 57870 203300 57876
rect 204076 57928 204128 57934
rect 204076 57870 204128 57876
rect 203260 57769 203288 57870
rect 203246 57760 203302 57769
rect 203246 57695 203302 57704
rect 204088 56710 204116 57870
rect 204076 56704 204128 56710
rect 204076 56646 204128 56652
rect 202880 52420 202932 52426
rect 202880 52362 202932 52368
rect 204076 52420 204128 52426
rect 204076 52362 204128 52368
rect 204088 51746 204116 52362
rect 204076 51740 204128 51746
rect 204076 51682 204128 51688
rect 203064 48272 203116 48278
rect 203062 48240 203064 48249
rect 204076 48272 204128 48278
rect 203116 48240 203118 48249
rect 204076 48214 204128 48220
rect 203062 48175 203118 48184
rect 204088 46986 204116 48214
rect 204076 46980 204128 46986
rect 204076 46922 204128 46928
rect 202696 11688 202748 11694
rect 202696 11630 202748 11636
rect 200776 6886 200896 6914
rect 201512 6886 201632 6914
rect 199078 354 199190 480
rect 198752 326 199190 354
rect 199078 -960 199190 326
rect 200274 354 200386 480
rect 200776 354 200804 6886
rect 201512 480 201540 6886
rect 202708 480 202736 11630
rect 203892 4140 203944 4146
rect 203892 4082 203944 4088
rect 203904 480 203932 4082
rect 204180 3398 204208 66030
rect 204260 49156 204312 49162
rect 204260 49098 204312 49104
rect 204272 16574 204300 49098
rect 204548 44985 204576 148650
rect 204640 72894 204668 192850
rect 204732 74458 204760 194074
rect 205916 193044 205968 193050
rect 205916 192986 205968 192992
rect 205178 192808 205234 192817
rect 205178 192743 205234 192752
rect 204810 192536 204866 192545
rect 204810 192471 204866 192480
rect 204824 75313 204852 192471
rect 205088 151360 205140 151366
rect 205088 151302 205140 151308
rect 204996 151224 205048 151230
rect 204996 151166 205048 151172
rect 204902 148744 204958 148753
rect 204902 148679 204958 148688
rect 204810 75304 204866 75313
rect 204810 75239 204866 75248
rect 204720 74452 204772 74458
rect 204720 74394 204772 74400
rect 204628 72888 204680 72894
rect 204628 72830 204680 72836
rect 204916 49706 204944 148679
rect 205008 57866 205036 151166
rect 205100 72865 205128 151302
rect 205086 72856 205142 72865
rect 205086 72791 205142 72800
rect 204996 57860 205048 57866
rect 204996 57802 205048 57808
rect 205008 57254 205036 57802
rect 204996 57248 205048 57254
rect 204996 57190 205048 57196
rect 205192 55214 205220 192743
rect 205822 192672 205878 192681
rect 205822 192607 205878 192616
rect 205640 192432 205692 192438
rect 205640 192374 205692 192380
rect 205652 70106 205680 192374
rect 205732 191548 205784 191554
rect 205732 191490 205784 191496
rect 205744 70378 205772 191490
rect 205836 78538 205864 192607
rect 205824 78532 205876 78538
rect 205824 78474 205876 78480
rect 205928 78418 205956 192986
rect 206008 192976 206060 192982
rect 206008 192918 206060 192924
rect 205836 78390 205956 78418
rect 205836 75750 205864 78390
rect 205916 78328 205968 78334
rect 205916 78270 205968 78276
rect 205824 75744 205876 75750
rect 205824 75686 205876 75692
rect 205836 75342 205864 75686
rect 205928 75614 205956 78270
rect 206020 75682 206048 192918
rect 206112 143177 206140 259490
rect 471256 206990 471284 261258
rect 485044 260160 485096 260166
rect 485044 260102 485096 260108
rect 485056 245614 485084 260102
rect 580172 259412 580224 259418
rect 580172 259354 580224 259360
rect 580184 258913 580212 259354
rect 580170 258904 580226 258913
rect 580170 258839 580226 258848
rect 485044 245608 485096 245614
rect 580172 245608 580224 245614
rect 485044 245550 485096 245556
rect 580170 245576 580172 245585
rect 580224 245576 580226 245585
rect 580170 245511 580226 245520
rect 580368 219065 580396 262958
rect 580448 262880 580500 262886
rect 580448 262822 580500 262828
rect 580460 232393 580488 262822
rect 580446 232384 580502 232393
rect 580446 232319 580502 232328
rect 580354 219056 580410 219065
rect 580354 218991 580410 219000
rect 471244 206984 471296 206990
rect 471244 206926 471296 206932
rect 579804 206984 579856 206990
rect 579804 206926 579856 206932
rect 579816 205737 579844 206926
rect 579802 205728 579858 205737
rect 579802 205663 579858 205672
rect 215668 199640 215720 199646
rect 215668 199582 215720 199588
rect 215392 199572 215444 199578
rect 215392 199514 215444 199520
rect 207112 198552 207164 198558
rect 207112 198494 207164 198500
rect 207018 194168 207074 194177
rect 207018 194103 207074 194112
rect 206192 152788 206244 152794
rect 206192 152730 206244 152736
rect 206098 143168 206154 143177
rect 206098 143103 206154 143112
rect 206098 141536 206154 141545
rect 206098 141471 206154 141480
rect 206008 75676 206060 75682
rect 206008 75618 206060 75624
rect 205916 75608 205968 75614
rect 205916 75550 205968 75556
rect 205824 75336 205876 75342
rect 205824 75278 205876 75284
rect 205928 75274 205956 75550
rect 205916 75268 205968 75274
rect 205916 75210 205968 75216
rect 205732 70372 205784 70378
rect 205732 70314 205784 70320
rect 205640 70100 205692 70106
rect 205640 70042 205692 70048
rect 205008 55186 205220 55214
rect 204904 49700 204956 49706
rect 204904 49642 204956 49648
rect 204916 49026 204944 49642
rect 205008 49337 205036 55186
rect 204994 49328 205050 49337
rect 204994 49263 205050 49272
rect 205008 49065 205036 49263
rect 204994 49056 205050 49065
rect 204904 49020 204956 49026
rect 204994 48991 205050 49000
rect 204904 48962 204956 48968
rect 204534 44976 204590 44985
rect 204534 44911 204590 44920
rect 205640 36848 205692 36854
rect 205640 36790 205692 36796
rect 205652 16574 205680 36790
rect 206112 35873 206140 141471
rect 206204 71738 206232 152730
rect 206376 151292 206428 151298
rect 206376 151234 206428 151240
rect 206284 151088 206336 151094
rect 206284 151030 206336 151036
rect 206296 75138 206324 151030
rect 206388 78033 206416 151234
rect 206468 148436 206520 148442
rect 206468 148378 206520 148384
rect 206480 80889 206508 148378
rect 206466 80880 206522 80889
rect 206466 80815 206522 80824
rect 206374 78024 206430 78033
rect 206374 77959 206430 77968
rect 206374 75848 206430 75857
rect 206374 75783 206376 75792
rect 206428 75783 206430 75792
rect 206376 75754 206428 75760
rect 206284 75132 206336 75138
rect 206284 75074 206336 75080
rect 206388 74594 206416 75754
rect 206376 74588 206428 74594
rect 206376 74530 206428 74536
rect 206192 71732 206244 71738
rect 206192 71674 206244 71680
rect 207032 45257 207060 194103
rect 207124 72418 207152 198494
rect 208584 198484 208636 198490
rect 208584 198426 208636 198432
rect 207204 194404 207256 194410
rect 207204 194346 207256 194352
rect 207112 72412 207164 72418
rect 207112 72354 207164 72360
rect 207216 69465 207244 194346
rect 208492 194336 208544 194342
rect 208492 194278 208544 194284
rect 207480 194064 207532 194070
rect 207480 194006 207532 194012
rect 207388 191480 207440 191486
rect 207388 191422 207440 191428
rect 207296 191344 207348 191350
rect 207296 191286 207348 191292
rect 207202 69456 207258 69465
rect 207202 69391 207258 69400
rect 207308 69018 207336 191286
rect 207400 71670 207428 191422
rect 207492 78402 207520 194006
rect 207572 192840 207624 192846
rect 207572 192782 207624 192788
rect 207480 78396 207532 78402
rect 207480 78338 207532 78344
rect 207584 78282 207612 192782
rect 207664 192772 207716 192778
rect 207664 192714 207716 192720
rect 207492 78254 207612 78282
rect 207492 75478 207520 78254
rect 207676 76974 207704 192714
rect 208398 189816 208454 189825
rect 208398 189751 208454 189760
rect 207756 151156 207808 151162
rect 207756 151098 207808 151104
rect 207664 76968 207716 76974
rect 207664 76910 207716 76916
rect 207480 75472 207532 75478
rect 207480 75414 207532 75420
rect 207492 75206 207520 75414
rect 207480 75200 207532 75206
rect 207480 75142 207532 75148
rect 207388 71664 207440 71670
rect 207388 71606 207440 71612
rect 207296 69012 207348 69018
rect 207296 68954 207348 68960
rect 207664 65748 207716 65754
rect 207664 65690 207716 65696
rect 207112 51060 207164 51066
rect 207112 51002 207164 51008
rect 207124 50386 207152 51002
rect 207112 50380 207164 50386
rect 207112 50322 207164 50328
rect 207112 46912 207164 46918
rect 207112 46854 207164 46860
rect 207124 46617 207152 46854
rect 207110 46608 207166 46617
rect 207110 46543 207166 46552
rect 207018 45248 207074 45257
rect 207018 45183 207074 45192
rect 207032 44849 207060 45183
rect 207018 44840 207074 44849
rect 207018 44775 207074 44784
rect 207018 44160 207074 44169
rect 207018 44095 207020 44104
rect 207072 44095 207074 44104
rect 207020 44066 207072 44072
rect 207032 42838 207060 44066
rect 207020 42832 207072 42838
rect 207020 42774 207072 42780
rect 206098 35864 206154 35873
rect 206098 35799 206154 35808
rect 206112 35193 206140 35799
rect 206098 35184 206154 35193
rect 206098 35119 206154 35128
rect 204272 16546 205128 16574
rect 205652 16546 206232 16574
rect 204168 3392 204220 3398
rect 204168 3334 204220 3340
rect 205100 480 205128 16546
rect 206204 480 206232 16546
rect 207676 4146 207704 65690
rect 207768 51066 207796 151098
rect 207846 147112 207902 147121
rect 207846 147047 207902 147056
rect 207860 78198 207888 147047
rect 207940 78396 207992 78402
rect 207940 78338 207992 78344
rect 207848 78192 207900 78198
rect 207848 78134 207900 78140
rect 207952 75041 207980 78338
rect 207938 75032 207994 75041
rect 207938 74967 207994 74976
rect 207756 51060 207808 51066
rect 207756 51002 207808 51008
rect 207846 46608 207902 46617
rect 207846 46543 207902 46552
rect 207860 45626 207888 46543
rect 207848 45620 207900 45626
rect 207848 45562 207900 45568
rect 208412 43489 208440 189751
rect 208504 51785 208532 194278
rect 208596 56545 208624 198426
rect 212816 198416 212868 198422
rect 212816 198358 212868 198364
rect 211344 198348 211396 198354
rect 211344 198290 211396 198296
rect 209964 198280 210016 198286
rect 209964 198222 210016 198228
rect 209780 198008 209832 198014
rect 209780 197950 209832 197956
rect 208676 195492 208728 195498
rect 208676 195434 208728 195440
rect 208688 67318 208716 195434
rect 208860 193996 208912 194002
rect 208860 193938 208912 193944
rect 208768 192704 208820 192710
rect 208768 192646 208820 192652
rect 208676 67312 208728 67318
rect 208676 67254 208728 67260
rect 208780 66230 208808 192646
rect 208872 67454 208900 193938
rect 208952 193928 209004 193934
rect 208952 193870 209004 193876
rect 208860 67448 208912 67454
rect 208860 67390 208912 67396
rect 208964 66842 208992 193870
rect 209044 191412 209096 191418
rect 209044 191354 209096 191360
rect 209056 71777 209084 191354
rect 209136 159520 209188 159526
rect 209136 159462 209188 159468
rect 209148 77654 209176 159462
rect 209228 142860 209280 142866
rect 209228 142802 209280 142808
rect 209136 77648 209188 77654
rect 209136 77590 209188 77596
rect 209042 71768 209098 71777
rect 209042 71703 209098 71712
rect 209148 70378 209176 77590
rect 209240 76537 209268 142802
rect 209226 76528 209282 76537
rect 209226 76463 209282 76472
rect 209136 70372 209188 70378
rect 209136 70314 209188 70320
rect 208952 66836 209004 66842
rect 208952 66778 209004 66784
rect 208768 66224 208820 66230
rect 208768 66166 208820 66172
rect 208582 56536 208638 56545
rect 208582 56471 208638 56480
rect 208950 56536 209006 56545
rect 208950 56471 209006 56480
rect 208964 55865 208992 56471
rect 208950 55856 209006 55865
rect 208950 55791 209006 55800
rect 208490 51776 208546 51785
rect 208490 51711 208546 51720
rect 208398 43480 208454 43489
rect 208398 43415 208454 43424
rect 208400 32700 208452 32706
rect 208400 32642 208452 32648
rect 208412 16574 208440 32642
rect 209792 20641 209820 197950
rect 209976 47569 210004 198222
rect 210148 194268 210200 194274
rect 210148 194210 210200 194216
rect 210054 147384 210110 147393
rect 210054 147319 210110 147328
rect 209962 47560 210018 47569
rect 209962 47495 210018 47504
rect 209870 43888 209926 43897
rect 209870 43823 209926 43832
rect 209778 20632 209834 20641
rect 209778 20567 209834 20576
rect 208412 16546 208624 16574
rect 207664 4140 207716 4146
rect 207664 4082 207716 4088
rect 207388 3392 207440 3398
rect 207388 3334 207440 3340
rect 207400 480 207428 3334
rect 208596 480 208624 16546
rect 209884 6914 209912 43823
rect 210068 24857 210096 147319
rect 210160 77489 210188 194210
rect 211252 192636 211304 192642
rect 211252 192578 211304 192584
rect 211160 192568 211212 192574
rect 211160 192510 211212 192516
rect 210700 192500 210752 192506
rect 210700 192442 210752 192448
rect 210240 190120 210292 190126
rect 210240 190062 210292 190068
rect 210146 77480 210202 77489
rect 210146 77415 210202 77424
rect 210252 76945 210280 190062
rect 210332 190052 210384 190058
rect 210332 189994 210384 190000
rect 210344 77081 210372 189994
rect 210424 189984 210476 189990
rect 210424 189926 210476 189932
rect 210436 78810 210464 189926
rect 210514 159352 210570 159361
rect 210514 159287 210570 159296
rect 210424 78804 210476 78810
rect 210424 78746 210476 78752
rect 210330 77072 210386 77081
rect 210330 77007 210386 77016
rect 210238 76936 210294 76945
rect 210238 76871 210294 76880
rect 210424 70372 210476 70378
rect 210424 70314 210476 70320
rect 210054 24848 210110 24857
rect 210054 24783 210110 24792
rect 209792 6886 209912 6914
rect 209792 480 209820 6886
rect 210436 3330 210464 70314
rect 210528 69698 210556 159287
rect 210608 157140 210660 157146
rect 210608 157082 210660 157088
rect 210620 77897 210648 157082
rect 210606 77888 210662 77897
rect 210606 77823 210662 77832
rect 210516 69692 210568 69698
rect 210516 69634 210568 69640
rect 210712 42809 210740 192442
rect 210698 42800 210754 42809
rect 210698 42735 210754 42744
rect 211066 42800 211122 42809
rect 211066 42735 211122 42744
rect 211080 42129 211108 42735
rect 211066 42120 211122 42129
rect 211066 42055 211122 42064
rect 211066 24848 211122 24857
rect 211066 24783 211122 24792
rect 211080 24177 211108 24783
rect 211066 24168 211122 24177
rect 211066 24103 211122 24112
rect 211172 21457 211200 192510
rect 211264 28937 211292 192578
rect 211356 55185 211384 198290
rect 212724 198144 212776 198150
rect 212724 198086 212776 198092
rect 211802 197976 211858 197985
rect 211802 197911 211858 197920
rect 211528 195288 211580 195294
rect 211528 195230 211580 195236
rect 211436 187196 211488 187202
rect 211436 187138 211488 187144
rect 211448 66094 211476 187138
rect 211540 74526 211568 195230
rect 211620 194200 211672 194206
rect 211620 194142 211672 194148
rect 211528 74520 211580 74526
rect 211528 74462 211580 74468
rect 211540 73982 211568 74462
rect 211632 74390 211660 194142
rect 211712 187128 211764 187134
rect 211712 187070 211764 187076
rect 211724 84194 211752 187070
rect 211816 89010 211844 197911
rect 211896 189916 211948 189922
rect 211896 189858 211948 189864
rect 211804 89004 211856 89010
rect 211804 88946 211856 88952
rect 211724 84166 211844 84194
rect 211620 74384 211672 74390
rect 211620 74326 211672 74332
rect 211528 73976 211580 73982
rect 211816 73953 211844 84166
rect 211908 77722 211936 189858
rect 212540 189848 212592 189854
rect 212540 189790 212592 189796
rect 211988 159588 212040 159594
rect 211988 159530 212040 159536
rect 212000 80102 212028 159530
rect 212080 89004 212132 89010
rect 212080 88946 212132 88952
rect 211988 80096 212040 80102
rect 211988 80038 212040 80044
rect 212092 78606 212120 88946
rect 212356 80096 212408 80102
rect 212356 80038 212408 80044
rect 212368 78946 212396 80038
rect 212356 78940 212408 78946
rect 212356 78882 212408 78888
rect 212448 78804 212500 78810
rect 212448 78746 212500 78752
rect 212460 78606 212488 78746
rect 212080 78600 212132 78606
rect 212080 78542 212132 78548
rect 212448 78600 212500 78606
rect 212448 78542 212500 78548
rect 211896 77716 211948 77722
rect 211896 77658 211948 77664
rect 211528 73918 211580 73924
rect 211802 73944 211858 73953
rect 211802 73879 211858 73888
rect 211436 66088 211488 66094
rect 211436 66030 211488 66036
rect 211342 55176 211398 55185
rect 211342 55111 211398 55120
rect 211356 54641 211384 55111
rect 211342 54632 211398 54641
rect 211342 54567 211398 54576
rect 211250 28928 211306 28937
rect 211250 28863 211306 28872
rect 211158 21448 211214 21457
rect 211158 21383 211214 21392
rect 211066 20632 211122 20641
rect 211066 20567 211122 20576
rect 211080 19961 211108 20567
rect 211066 19952 211122 19961
rect 211066 19887 211122 19896
rect 211816 4146 211844 73879
rect 212446 28928 212502 28937
rect 212446 28863 212502 28872
rect 212460 28257 212488 28863
rect 212446 28248 212502 28257
rect 212446 28183 212502 28192
rect 212552 22001 212580 189790
rect 212630 187368 212686 187377
rect 212630 187303 212686 187312
rect 212644 49609 212672 187303
rect 212736 64705 212764 198086
rect 212828 68950 212856 198358
rect 212908 198212 212960 198218
rect 212908 198154 212960 198160
rect 212920 75886 212948 198154
rect 213000 198076 213052 198082
rect 213000 198018 213052 198024
rect 213012 77625 213040 198018
rect 214012 187264 214064 187270
rect 214012 187206 214064 187212
rect 215298 187232 215354 187241
rect 213920 159452 213972 159458
rect 213920 159394 213972 159400
rect 213092 152652 213144 152658
rect 213092 152594 213144 152600
rect 212998 77616 213054 77625
rect 212998 77551 213054 77560
rect 212908 75880 212960 75886
rect 212908 75822 212960 75828
rect 212816 68944 212868 68950
rect 212816 68886 212868 68892
rect 213104 65521 213132 152594
rect 213826 78160 213882 78169
rect 213826 78095 213882 78104
rect 213840 77625 213868 78095
rect 213826 77616 213882 77625
rect 213826 77551 213882 77560
rect 213932 77246 213960 159394
rect 213920 77240 213972 77246
rect 213920 77182 213972 77188
rect 213828 68944 213880 68950
rect 213828 68886 213880 68892
rect 213840 68338 213868 68886
rect 213828 68332 213880 68338
rect 213828 68274 213880 68280
rect 213090 65512 213146 65521
rect 213090 65447 213146 65456
rect 212722 64696 212778 64705
rect 212722 64631 212778 64640
rect 212736 64161 212764 64631
rect 212722 64152 212778 64161
rect 212722 64087 212778 64096
rect 213918 62928 213974 62937
rect 213918 62863 213974 62872
rect 212630 49600 212686 49609
rect 212630 49535 212686 49544
rect 213826 49600 213882 49609
rect 213826 49535 213882 49544
rect 213840 48929 213868 49535
rect 213826 48920 213882 48929
rect 213826 48855 213882 48864
rect 212538 21992 212594 22001
rect 212538 21927 212594 21936
rect 213826 21992 213882 22001
rect 213826 21927 213882 21936
rect 213840 21321 213868 21927
rect 213826 21312 213882 21321
rect 213826 21247 213882 21256
rect 213932 16574 213960 62863
rect 214024 58993 214052 187206
rect 215298 187167 215354 187176
rect 214196 159384 214248 159390
rect 214196 159326 214248 159332
rect 214102 142760 214158 142769
rect 214102 142695 214158 142704
rect 214010 58984 214066 58993
rect 214010 58919 214066 58928
rect 214116 37233 214144 142695
rect 214208 77217 214236 159326
rect 214288 152516 214340 152522
rect 214288 152458 214340 152464
rect 214194 77208 214250 77217
rect 214300 77178 214328 152458
rect 214378 146976 214434 146985
rect 214378 146911 214434 146920
rect 214472 146940 214524 146946
rect 214194 77143 214250 77152
rect 214288 77172 214340 77178
rect 214288 77114 214340 77120
rect 214392 76294 214420 146911
rect 214472 146882 214524 146888
rect 214484 76838 214512 146882
rect 214564 145648 214616 145654
rect 214564 145590 214616 145596
rect 214576 79422 214604 145590
rect 214656 142928 214708 142934
rect 214656 142870 214708 142876
rect 214668 79626 214696 142870
rect 214656 79620 214708 79626
rect 214656 79562 214708 79568
rect 214668 79422 214696 79562
rect 214564 79416 214616 79422
rect 214564 79358 214616 79364
rect 214656 79416 214708 79422
rect 214656 79358 214708 79364
rect 214564 77172 214616 77178
rect 214564 77114 214616 77120
rect 214472 76832 214524 76838
rect 214472 76774 214524 76780
rect 214576 76770 214604 77114
rect 214564 76764 214616 76770
rect 214564 76706 214616 76712
rect 214380 76288 214432 76294
rect 214380 76230 214432 76236
rect 215312 50969 215340 187167
rect 215404 64433 215432 199514
rect 215484 199368 215536 199374
rect 215484 199310 215536 199316
rect 215496 67017 215524 199310
rect 215574 186960 215630 186969
rect 215574 186895 215630 186904
rect 215588 68921 215616 186895
rect 215680 80850 215708 199582
rect 216772 193860 216824 193866
rect 216772 193802 216824 193808
rect 215758 187096 215814 187105
rect 215758 187031 215814 187040
rect 215852 187060 215904 187066
rect 215668 80844 215720 80850
rect 215668 80786 215720 80792
rect 215772 74225 215800 187031
rect 215852 187002 215904 187008
rect 215864 80782 215892 187002
rect 215852 80776 215904 80782
rect 215852 80718 215904 80724
rect 216680 75404 216732 75410
rect 216680 75346 216732 75352
rect 215758 74216 215814 74225
rect 215758 74151 215814 74160
rect 215772 73681 215800 74151
rect 215758 73672 215814 73681
rect 215758 73607 215814 73616
rect 215574 68912 215630 68921
rect 215574 68847 215630 68856
rect 215482 67008 215538 67017
rect 215482 66943 215538 66952
rect 215390 64424 215446 64433
rect 215390 64359 215446 64368
rect 215298 50960 215354 50969
rect 215298 50895 215354 50904
rect 215300 47660 215352 47666
rect 215300 47602 215352 47608
rect 214102 37224 214158 37233
rect 214102 37159 214158 37168
rect 214378 37224 214434 37233
rect 214378 37159 214434 37168
rect 214392 36553 214420 37159
rect 214378 36544 214434 36553
rect 214378 36479 214434 36488
rect 213932 16546 214512 16574
rect 213366 8936 213422 8945
rect 213366 8871 213422 8880
rect 210976 4140 211028 4146
rect 210976 4082 211028 4088
rect 211804 4140 211856 4146
rect 211804 4082 211856 4088
rect 210424 3324 210476 3330
rect 210424 3266 210476 3272
rect 210988 480 211016 4082
rect 212172 4004 212224 4010
rect 212172 3946 212224 3952
rect 212184 480 212212 3946
rect 213380 480 213408 8871
rect 214484 480 214512 16546
rect 200274 326 200804 354
rect 200274 -960 200386 326
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203862 -960 203974 480
rect 205058 -960 205170 480
rect 206162 -960 206274 480
rect 207358 -960 207470 480
rect 208554 -960 208666 480
rect 209750 -960 209862 480
rect 210946 -960 211058 480
rect 212142 -960 212254 480
rect 213338 -960 213450 480
rect 214442 -960 214554 480
rect 215312 354 215340 47602
rect 216692 16574 216720 75346
rect 216784 73166 216812 193802
rect 580172 193180 580224 193186
rect 580172 193122 580224 193128
rect 580184 192545 580212 193122
rect 580170 192536 580226 192545
rect 580170 192471 580226 192480
rect 216864 191276 216916 191282
rect 216864 191218 216916 191224
rect 216876 73817 216904 191218
rect 218152 191208 218204 191214
rect 218152 191150 218204 191156
rect 218058 189680 218114 189689
rect 218058 189615 218114 189624
rect 216862 73808 216918 73817
rect 216862 73743 216918 73752
rect 216772 73160 216824 73166
rect 216772 73102 216824 73108
rect 216784 72894 216812 73102
rect 216772 72888 216824 72894
rect 216772 72830 216824 72836
rect 218072 45529 218100 189615
rect 218164 73137 218192 191150
rect 218244 191140 218296 191146
rect 218244 191082 218296 191088
rect 218256 74225 218284 191082
rect 218336 189780 218388 189786
rect 218336 189722 218388 189728
rect 218242 74216 218298 74225
rect 218242 74151 218298 74160
rect 218256 73409 218284 74151
rect 218348 74089 218376 189722
rect 218428 186992 218480 186998
rect 218428 186934 218480 186940
rect 218440 74361 218468 186934
rect 580170 179208 580226 179217
rect 580170 179143 580226 179152
rect 580184 178090 580212 179143
rect 580172 178084 580224 178090
rect 580172 178026 580224 178032
rect 580170 165880 580226 165889
rect 580170 165815 580226 165824
rect 580184 165646 580212 165815
rect 580172 165640 580224 165646
rect 580172 165582 580224 165588
rect 579986 152688 580042 152697
rect 579986 152623 580042 152632
rect 580000 151842 580028 152623
rect 579988 151836 580040 151842
rect 579988 151778 580040 151784
rect 580262 150512 580318 150521
rect 580262 150447 580318 150456
rect 464342 140992 464398 141001
rect 464342 140927 464398 140936
rect 327724 139460 327776 139466
rect 327724 139402 327776 139408
rect 270500 80844 270552 80850
rect 270500 80786 270552 80792
rect 234620 80776 234672 80782
rect 234620 80718 234672 80724
rect 218426 74352 218482 74361
rect 218426 74287 218482 74296
rect 218334 74080 218390 74089
rect 218334 74015 218390 74024
rect 218440 73545 218468 74287
rect 224222 73672 224278 73681
rect 224222 73607 224278 73616
rect 218426 73536 218482 73545
rect 218426 73471 218482 73480
rect 218242 73400 218298 73409
rect 218242 73335 218298 73344
rect 218150 73128 218206 73137
rect 218150 73063 218206 73072
rect 218164 72457 218192 73063
rect 220084 72888 220136 72894
rect 220084 72830 220136 72836
rect 218150 72448 218206 72457
rect 218150 72383 218206 72392
rect 218152 47592 218204 47598
rect 218152 47534 218204 47540
rect 218058 45520 218114 45529
rect 218058 45455 218114 45464
rect 218164 16574 218192 47534
rect 219440 46300 219492 46306
rect 219440 46242 219492 46248
rect 219452 16574 219480 46242
rect 216692 16546 216904 16574
rect 218164 16546 219296 16574
rect 219452 16546 220032 16574
rect 216876 480 216904 16546
rect 218060 3324 218112 3330
rect 218060 3266 218112 3272
rect 218072 480 218100 3266
rect 219268 480 219296 16546
rect 215638 354 215750 480
rect 215312 326 215750 354
rect 215638 -960 215750 326
rect 216834 -960 216946 480
rect 218030 -960 218142 480
rect 219226 -960 219338 480
rect 220004 354 220032 16546
rect 220096 4010 220124 72830
rect 220818 68912 220874 68921
rect 220818 68847 220874 68856
rect 220832 16574 220860 68847
rect 222200 31340 222252 31346
rect 222200 31282 222252 31288
rect 222212 16574 222240 31282
rect 220832 16546 221136 16574
rect 222212 16546 222792 16574
rect 220084 4004 220136 4010
rect 220084 3946 220136 3952
rect 220422 354 220534 480
rect 220004 326 220534 354
rect 221108 354 221136 16546
rect 222764 480 222792 16546
rect 223948 4140 224000 4146
rect 223948 4082 224000 4088
rect 223960 480 223988 4082
rect 224236 3330 224264 73607
rect 227718 67008 227774 67017
rect 227718 66943 227774 66952
rect 224960 51808 225012 51814
rect 224960 51750 225012 51756
rect 224972 16574 225000 51750
rect 227732 16574 227760 66943
rect 231860 60308 231912 60314
rect 231860 60250 231912 60256
rect 229100 55956 229152 55962
rect 229100 55898 229152 55904
rect 229112 16574 229140 55898
rect 224972 16546 225184 16574
rect 227732 16546 228312 16574
rect 229112 16546 229416 16574
rect 224224 3324 224276 3330
rect 224224 3266 224276 3272
rect 225156 480 225184 16546
rect 226340 12028 226392 12034
rect 226340 11970 226392 11976
rect 226352 480 226380 11970
rect 227536 9240 227588 9246
rect 227536 9182 227588 9188
rect 227548 480 227576 9182
rect 221526 354 221638 480
rect 221108 326 221638 354
rect 220422 -960 220534 326
rect 221526 -960 221638 326
rect 222722 -960 222834 480
rect 223918 -960 224030 480
rect 225114 -960 225226 480
rect 226310 -960 226422 480
rect 227506 -960 227618 480
rect 228284 354 228312 16546
rect 228702 354 228814 480
rect 228284 326 228814 354
rect 229388 354 229416 16546
rect 231032 3324 231084 3330
rect 231032 3266 231084 3272
rect 231044 480 231072 3266
rect 229806 354 229918 480
rect 229388 326 229918 354
rect 228702 -960 228814 326
rect 229806 -960 229918 326
rect 231002 -960 231114 480
rect 231872 354 231900 60250
rect 233240 41064 233292 41070
rect 233240 41006 233292 41012
rect 233252 16574 233280 41006
rect 233252 16546 233464 16574
rect 233436 480 233464 16546
rect 234632 11694 234660 80718
rect 238760 80164 238812 80170
rect 238760 80106 238812 80112
rect 237378 74352 237434 74361
rect 237378 74287 237434 74296
rect 236000 34128 236052 34134
rect 236000 34070 236052 34076
rect 236012 16574 236040 34070
rect 237392 16574 237420 74287
rect 238772 16574 238800 80106
rect 253940 76900 253992 76906
rect 253940 76842 253992 76848
rect 248418 74216 248474 74225
rect 248418 74151 248474 74160
rect 242162 64424 242218 64433
rect 242162 64359 242218 64368
rect 239404 54596 239456 54602
rect 239404 54538 239456 54544
rect 236012 16546 236592 16574
rect 237392 16546 237696 16574
rect 238772 16546 239352 16574
rect 234620 11688 234672 11694
rect 234620 11630 234672 11636
rect 235816 11688 235868 11694
rect 235816 11630 235868 11636
rect 234620 10600 234672 10606
rect 234620 10542 234672 10548
rect 234632 480 234660 10542
rect 235828 480 235856 11630
rect 232198 354 232310 480
rect 231872 326 232310 354
rect 232198 -960 232310 326
rect 233394 -960 233506 480
rect 234590 -960 234702 480
rect 235786 -960 235898 480
rect 236564 354 236592 16546
rect 236982 354 237094 480
rect 236564 326 237094 354
rect 237668 354 237696 16546
rect 239324 480 239352 16546
rect 239416 3398 239444 54538
rect 241704 7880 241756 7886
rect 241704 7822 241756 7828
rect 239404 3392 239456 3398
rect 239404 3334 239456 3340
rect 240508 3392 240560 3398
rect 240508 3334 240560 3340
rect 240520 480 240548 3334
rect 241716 480 241744 7822
rect 242176 4146 242204 64359
rect 245660 62960 245712 62966
rect 245660 62902 245712 62908
rect 242900 44940 242952 44946
rect 242900 44882 242952 44888
rect 242164 4140 242216 4146
rect 242164 4082 242216 4088
rect 242912 480 242940 44882
rect 242992 32632 243044 32638
rect 242992 32574 243044 32580
rect 243004 16574 243032 32574
rect 245672 16574 245700 62902
rect 243004 16546 244136 16574
rect 245672 16546 245976 16574
rect 244108 480 244136 16546
rect 245200 5024 245252 5030
rect 245200 4966 245252 4972
rect 245212 480 245240 4966
rect 238086 354 238198 480
rect 237668 326 238198 354
rect 236982 -960 237094 326
rect 238086 -960 238198 326
rect 239282 -960 239394 480
rect 240478 -960 240590 480
rect 241674 -960 241786 480
rect 242870 -960 242982 480
rect 244066 -960 244178 480
rect 245170 -960 245282 480
rect 245948 354 245976 16546
rect 247592 4072 247644 4078
rect 247592 4014 247644 4020
rect 247604 480 247632 4014
rect 246366 354 246478 480
rect 245948 326 246478 354
rect 246366 -960 246478 326
rect 247562 -960 247674 480
rect 248432 354 248460 74151
rect 252560 68536 252612 68542
rect 252560 68478 252612 68484
rect 249800 58744 249852 58750
rect 249800 58686 249852 58692
rect 249812 16574 249840 58686
rect 251180 34060 251232 34066
rect 251180 34002 251232 34008
rect 249812 16546 250024 16574
rect 249996 480 250024 16546
rect 251192 480 251220 34002
rect 251272 18896 251324 18902
rect 251272 18838 251324 18844
rect 251284 16574 251312 18838
rect 252572 16574 252600 68478
rect 253952 16574 253980 76842
rect 260102 76664 260158 76673
rect 260102 76599 260158 76608
rect 255320 73976 255372 73982
rect 255320 73918 255372 73924
rect 255332 16574 255360 73918
rect 256698 50688 256754 50697
rect 256698 50623 256754 50632
rect 251284 16546 252416 16574
rect 252572 16546 253520 16574
rect 253952 16546 254256 16574
rect 255332 16546 255912 16574
rect 252388 480 252416 16546
rect 253492 480 253520 16546
rect 248758 354 248870 480
rect 248432 326 248870 354
rect 248758 -960 248870 326
rect 249954 -960 250066 480
rect 251150 -960 251262 480
rect 252346 -960 252458 480
rect 253450 -960 253562 480
rect 254228 354 254256 16546
rect 255884 480 255912 16546
rect 254646 354 254758 480
rect 254228 326 254758 354
rect 254646 -960 254758 326
rect 255842 -960 255954 480
rect 256712 354 256740 50623
rect 259552 17468 259604 17474
rect 259552 17410 259604 17416
rect 258264 13388 258316 13394
rect 258264 13330 258316 13336
rect 258276 480 258304 13330
rect 259564 6914 259592 17410
rect 259472 6886 259592 6914
rect 259472 480 259500 6886
rect 260116 3330 260144 76599
rect 261482 73944 261538 73953
rect 261482 73879 261538 73888
rect 269120 73908 269172 73914
rect 260656 4140 260708 4146
rect 260656 4082 260708 4088
rect 260104 3324 260156 3330
rect 260104 3266 260156 3272
rect 260668 480 260696 4082
rect 261496 3398 261524 73879
rect 269120 73850 269172 73856
rect 263600 57316 263652 57322
rect 263600 57258 263652 57264
rect 263612 16574 263640 57258
rect 267740 53168 267792 53174
rect 267740 53110 267792 53116
rect 266360 39568 266412 39574
rect 266360 39510 266412 39516
rect 264980 31272 265032 31278
rect 264980 31214 265032 31220
rect 263612 16546 264192 16574
rect 261484 3392 261536 3398
rect 261484 3334 261536 3340
rect 262956 3392 263008 3398
rect 262956 3334 263008 3340
rect 261760 3324 261812 3330
rect 261760 3266 261812 3272
rect 261772 480 261800 3266
rect 262968 480 262996 3334
rect 264164 480 264192 16546
rect 257038 354 257150 480
rect 256712 326 257150 354
rect 257038 -960 257150 326
rect 258234 -960 258346 480
rect 259430 -960 259542 480
rect 260626 -960 260738 480
rect 261730 -960 261842 480
rect 262926 -960 263038 480
rect 264122 -960 264234 480
rect 264992 354 265020 31214
rect 266372 16574 266400 39510
rect 266372 16546 266584 16574
rect 266556 480 266584 16546
rect 267752 480 267780 53110
rect 267832 36780 267884 36786
rect 267832 36722 267884 36728
rect 267844 16574 267872 36722
rect 269132 16574 269160 73850
rect 270512 16574 270540 80786
rect 302240 80708 302292 80714
rect 302240 80650 302292 80656
rect 288438 79520 288494 79529
rect 288438 79455 288494 79464
rect 274638 78840 274694 78849
rect 274638 78775 274694 78784
rect 271880 27192 271932 27198
rect 271880 27134 271932 27140
rect 271892 16574 271920 27134
rect 274652 16574 274680 78775
rect 287704 72820 287756 72826
rect 287704 72762 287756 72768
rect 277400 61532 277452 61538
rect 277400 61474 277452 61480
rect 275282 37904 275338 37913
rect 275282 37839 275338 37848
rect 267844 16546 268424 16574
rect 269132 16546 270080 16574
rect 270512 16546 270816 16574
rect 271892 16546 272472 16574
rect 274652 16546 274864 16574
rect 265318 354 265430 480
rect 264992 326 265430 354
rect 265318 -960 265430 326
rect 266514 -960 266626 480
rect 267710 -960 267822 480
rect 268396 354 268424 16546
rect 270052 480 270080 16546
rect 268814 354 268926 480
rect 268396 326 268926 354
rect 268814 -960 268926 326
rect 270010 -960 270122 480
rect 270788 354 270816 16546
rect 272444 480 272472 16546
rect 273628 6792 273680 6798
rect 273628 6734 273680 6740
rect 273640 480 273668 6734
rect 274836 480 274864 16546
rect 275296 3398 275324 37839
rect 277412 16574 277440 61474
rect 281538 58984 281594 58993
rect 281538 58919 281594 58928
rect 279422 45248 279478 45257
rect 279422 45183 279478 45192
rect 278780 25764 278832 25770
rect 278780 25706 278832 25712
rect 278792 16574 278820 25706
rect 277412 16546 278360 16574
rect 278792 16546 279096 16574
rect 276020 14748 276072 14754
rect 276020 14690 276072 14696
rect 275284 3392 275336 3398
rect 275284 3334 275336 3340
rect 276032 480 276060 14690
rect 277124 3392 277176 3398
rect 277124 3334 277176 3340
rect 277136 480 277164 3334
rect 278332 480 278360 16546
rect 271206 354 271318 480
rect 270788 326 271318 354
rect 271206 -960 271318 326
rect 272402 -960 272514 480
rect 273598 -960 273710 480
rect 274794 -960 274906 480
rect 275990 -960 276102 480
rect 277094 -960 277206 480
rect 278290 -960 278402 480
rect 279068 354 279096 16546
rect 279436 3398 279464 45183
rect 279424 3392 279476 3398
rect 279424 3334 279476 3340
rect 280712 3392 280764 3398
rect 280712 3334 280764 3340
rect 280724 480 280752 3334
rect 279486 354 279598 480
rect 279068 326 279598 354
rect 279486 -960 279598 326
rect 280682 -960 280794 480
rect 281552 354 281580 58919
rect 284298 56264 284354 56273
rect 284298 56199 284354 56208
rect 282920 23044 282972 23050
rect 282920 22986 282972 22992
rect 282932 16574 282960 22986
rect 282932 16546 283144 16574
rect 283116 480 283144 16546
rect 284312 4078 284340 56199
rect 285680 46232 285732 46238
rect 285680 46174 285732 46180
rect 285692 16574 285720 46174
rect 287060 20120 287112 20126
rect 287060 20062 287112 20068
rect 287072 16574 287100 20062
rect 285692 16546 286640 16574
rect 287072 16546 287376 16574
rect 284392 16176 284444 16182
rect 284392 16118 284444 16124
rect 284300 4072 284352 4078
rect 284300 4014 284352 4020
rect 284404 3482 284432 16118
rect 285036 4072 285088 4078
rect 285036 4014 285088 4020
rect 284312 3454 284432 3482
rect 284312 480 284340 3454
rect 281878 354 281990 480
rect 281552 326 281990 354
rect 281878 -960 281990 326
rect 283074 -960 283186 480
rect 284270 -960 284382 480
rect 285048 354 285076 4014
rect 286612 480 286640 16546
rect 285374 354 285486 480
rect 285048 326 285486 354
rect 285374 -960 285486 326
rect 286570 -960 286682 480
rect 287348 354 287376 16546
rect 287716 4078 287744 72762
rect 288452 16574 288480 79455
rect 289820 76832 289872 76838
rect 289820 76774 289872 76780
rect 288452 16546 289032 16574
rect 287704 4072 287756 4078
rect 287704 4014 287756 4020
rect 289004 480 289032 16546
rect 287766 354 287878 480
rect 287348 326 287878 354
rect 287766 -960 287878 326
rect 288962 -960 289074 480
rect 289832 354 289860 76774
rect 296720 76764 296772 76770
rect 296720 76706 296772 76712
rect 295340 65680 295392 65686
rect 295340 65622 295392 65628
rect 292580 62892 292632 62898
rect 292580 62834 292632 62840
rect 291200 20052 291252 20058
rect 291200 19994 291252 20000
rect 291212 16574 291240 19994
rect 291212 16546 291424 16574
rect 291396 480 291424 16546
rect 292592 480 292620 62834
rect 292672 40996 292724 41002
rect 292672 40938 292724 40944
rect 292684 16574 292712 40938
rect 293958 19952 294014 19961
rect 293958 19887 294014 19896
rect 293972 16574 294000 19887
rect 295352 16574 295380 65622
rect 296732 16574 296760 76706
rect 299480 60240 299532 60246
rect 299480 60182 299532 60188
rect 292684 16546 293264 16574
rect 293972 16546 294920 16574
rect 295352 16546 295656 16574
rect 296732 16546 297312 16574
rect 290158 354 290270 480
rect 289832 326 290270 354
rect 290158 -960 290270 326
rect 291354 -960 291466 480
rect 292550 -960 292662 480
rect 293236 354 293264 16546
rect 294892 480 294920 16546
rect 293654 354 293766 480
rect 293236 326 293766 354
rect 293654 -960 293766 326
rect 294850 -960 294962 480
rect 295628 354 295656 16546
rect 297284 480 297312 16546
rect 298468 4004 298520 4010
rect 298468 3946 298520 3952
rect 298480 480 298508 3946
rect 299492 3482 299520 60182
rect 300858 42120 300914 42129
rect 300858 42055 300914 42064
rect 299572 29912 299624 29918
rect 299572 29854 299624 29860
rect 299584 4010 299612 29854
rect 300872 16574 300900 42055
rect 302252 16574 302280 80650
rect 324320 79484 324372 79490
rect 324320 79426 324372 79432
rect 305000 72752 305052 72758
rect 305000 72694 305052 72700
rect 303620 35420 303672 35426
rect 303620 35362 303672 35368
rect 303632 16574 303660 35362
rect 305012 16574 305040 72694
rect 322940 72684 322992 72690
rect 322940 72626 322992 72632
rect 317420 66904 317472 66910
rect 317420 66846 317472 66852
rect 306380 64252 306432 64258
rect 306380 64194 306432 64200
rect 300872 16546 301544 16574
rect 302252 16546 303200 16574
rect 303632 16546 303936 16574
rect 305012 16546 305592 16574
rect 299572 4004 299624 4010
rect 299572 3946 299624 3952
rect 300768 4004 300820 4010
rect 300768 3946 300820 3952
rect 299492 3454 299704 3482
rect 299676 480 299704 3454
rect 300780 480 300808 3946
rect 296046 354 296158 480
rect 295628 326 296158 354
rect 296046 -960 296158 326
rect 297242 -960 297354 480
rect 298438 -960 298550 480
rect 299634 -960 299746 480
rect 300738 -960 300850 480
rect 301516 354 301544 16546
rect 303172 480 303200 16546
rect 301934 354 302046 480
rect 301516 326 302046 354
rect 301934 -960 302046 326
rect 303130 -960 303242 480
rect 303908 354 303936 16546
rect 305564 480 305592 16546
rect 304326 354 304438 480
rect 303908 326 304438 354
rect 304326 -960 304438 326
rect 305522 -960 305634 480
rect 306392 354 306420 64194
rect 313280 61464 313332 61470
rect 313280 61406 313332 61412
rect 309138 43752 309194 43761
rect 309138 43687 309194 43696
rect 307022 28248 307078 28257
rect 307022 28183 307078 28192
rect 307036 3398 307064 28183
rect 309152 16574 309180 43687
rect 310518 24168 310574 24177
rect 310518 24103 310574 24112
rect 310532 16574 310560 24103
rect 313292 16574 313320 61406
rect 315304 54528 315356 54534
rect 315304 54470 315356 54476
rect 309152 16546 309824 16574
rect 310532 16546 311480 16574
rect 313292 16546 313872 16574
rect 307944 13320 307996 13326
rect 307944 13262 307996 13268
rect 307024 3392 307076 3398
rect 307024 3334 307076 3340
rect 307956 480 307984 13262
rect 309048 3392 309100 3398
rect 309048 3334 309100 3340
rect 309060 480 309088 3334
rect 306718 354 306830 480
rect 306392 326 306830 354
rect 306718 -960 306830 326
rect 307914 -960 308026 480
rect 309018 -960 309130 480
rect 309796 354 309824 16546
rect 311452 480 311480 16546
rect 312636 4072 312688 4078
rect 312636 4014 312688 4020
rect 312648 480 312676 4014
rect 313844 480 313872 16546
rect 314660 14680 314712 14686
rect 314660 14622 314712 14628
rect 310214 354 310326 480
rect 309796 326 310326 354
rect 310214 -960 310326 326
rect 311410 -960 311522 480
rect 312606 -960 312718 480
rect 313802 -960 313914 480
rect 314672 354 314700 14622
rect 315316 4146 315344 54470
rect 317432 16574 317460 66846
rect 320178 52184 320234 52193
rect 320178 52119 320234 52128
rect 318800 38140 318852 38146
rect 318800 38082 318852 38088
rect 318812 16574 318840 38082
rect 320192 16574 320220 52119
rect 321560 28484 321612 28490
rect 321560 28426 321612 28432
rect 321572 16574 321600 28426
rect 317432 16546 318104 16574
rect 318812 16546 319760 16574
rect 320192 16546 320496 16574
rect 321572 16546 322152 16574
rect 316224 9172 316276 9178
rect 316224 9114 316276 9120
rect 315304 4140 315356 4146
rect 315304 4082 315356 4088
rect 316236 480 316264 9114
rect 317328 4140 317380 4146
rect 317328 4082 317380 4088
rect 317340 480 317368 4082
rect 314998 354 315110 480
rect 314672 326 315110 354
rect 314998 -960 315110 326
rect 316194 -960 316306 480
rect 317298 -960 317410 480
rect 318076 354 318104 16546
rect 319732 480 319760 16546
rect 318494 354 318606 480
rect 318076 326 318606 354
rect 318494 -960 318606 326
rect 319690 -960 319802 480
rect 320468 354 320496 16546
rect 322124 480 322152 16546
rect 320886 354 320998 480
rect 320468 326 320998 354
rect 320886 -960 320998 326
rect 322082 -960 322194 480
rect 322952 354 322980 72626
rect 323584 72616 323636 72622
rect 323584 72558 323636 72564
rect 323596 4146 323624 72558
rect 323584 4140 323636 4146
rect 323584 4082 323636 4088
rect 324332 3210 324360 79426
rect 327736 73166 327764 139402
rect 464356 86970 464384 140927
rect 464344 86964 464396 86970
rect 464344 86906 464396 86912
rect 579620 86964 579672 86970
rect 579620 86906 579672 86912
rect 579632 86193 579660 86906
rect 579618 86184 579674 86193
rect 579618 86119 579674 86128
rect 505098 80744 505154 80753
rect 505098 80679 505154 80688
rect 358820 79416 358872 79422
rect 358820 79358 358872 79364
rect 353300 76696 353352 76702
rect 353300 76638 353352 76644
rect 340880 73840 340932 73846
rect 340880 73782 340932 73788
rect 347778 73808 347834 73817
rect 327724 73160 327776 73166
rect 327724 73102 327776 73108
rect 332598 72448 332654 72457
rect 332598 72383 332654 72392
rect 327080 58676 327132 58682
rect 327080 58618 327132 58624
rect 324412 42288 324464 42294
rect 324412 42230 324464 42236
rect 324424 3398 324452 42230
rect 327092 16574 327120 58618
rect 331220 55888 331272 55894
rect 331220 55830 331272 55836
rect 329102 21448 329158 21457
rect 329102 21383 329158 21392
rect 327092 16546 328040 16574
rect 326804 4140 326856 4146
rect 326804 4082 326856 4088
rect 324412 3392 324464 3398
rect 324412 3334 324464 3340
rect 325608 3392 325660 3398
rect 325608 3334 325660 3340
rect 324332 3182 324452 3210
rect 324424 480 324452 3182
rect 325620 480 325648 3334
rect 326816 480 326844 4082
rect 328012 480 328040 16546
rect 328736 11960 328788 11966
rect 328736 11902 328788 11908
rect 323278 354 323390 480
rect 322952 326 323390 354
rect 323278 -960 323390 326
rect 324382 -960 324494 480
rect 325578 -960 325690 480
rect 326774 -960 326886 480
rect 327970 -960 328082 480
rect 328748 354 328776 11902
rect 329116 3398 329144 21383
rect 329104 3392 329156 3398
rect 329104 3334 329156 3340
rect 330392 3392 330444 3398
rect 330392 3334 330444 3340
rect 330404 480 330432 3334
rect 329166 354 329278 480
rect 328748 326 329278 354
rect 329166 -960 329278 326
rect 330362 -960 330474 480
rect 331232 354 331260 55830
rect 332612 1154 332640 72383
rect 338118 50552 338174 50561
rect 338118 50487 338174 50496
rect 333980 40928 334032 40934
rect 333980 40870 334032 40876
rect 332692 32564 332744 32570
rect 332692 32506 332744 32512
rect 332600 1148 332652 1154
rect 332600 1090 332652 1096
rect 332704 480 332732 32506
rect 333992 16574 334020 40870
rect 336738 21312 336794 21321
rect 336738 21247 336794 21256
rect 336752 16574 336780 21247
rect 338132 16574 338160 50487
rect 339500 33992 339552 33998
rect 339500 33934 339552 33940
rect 333992 16546 334664 16574
rect 336752 16546 337056 16574
rect 338132 16546 338712 16574
rect 333888 1148 333940 1154
rect 333888 1090 333940 1096
rect 333900 480 333928 1090
rect 331558 354 331670 480
rect 331232 326 331670 354
rect 331558 -960 331670 326
rect 332662 -960 332774 480
rect 333858 -960 333970 480
rect 334636 354 334664 16546
rect 336280 10532 336332 10538
rect 336280 10474 336332 10480
rect 336292 480 336320 10474
rect 335054 354 335166 480
rect 334636 326 335166 354
rect 335054 -960 335166 326
rect 336250 -960 336362 480
rect 337028 354 337056 16546
rect 338684 480 338712 16546
rect 337446 354 337558 480
rect 337028 326 337558 354
rect 337446 -960 337558 326
rect 338642 -960 338754 480
rect 339512 354 339540 33934
rect 340892 3210 340920 73782
rect 347778 73743 347834 73752
rect 342904 72548 342956 72554
rect 342904 72490 342956 72496
rect 340972 60172 341024 60178
rect 340972 60114 341024 60120
rect 340984 3398 341012 60114
rect 342916 3398 342944 72490
rect 346400 31204 346452 31210
rect 346400 31146 346452 31152
rect 345020 18828 345072 18834
rect 345020 18770 345072 18776
rect 345032 16574 345060 18770
rect 346412 16574 346440 31146
rect 347792 16574 347820 73743
rect 351920 65612 351972 65618
rect 351920 65554 351972 65560
rect 349158 57352 349214 57361
rect 349158 57287 349214 57296
rect 349172 16574 349200 57287
rect 350540 21480 350592 21486
rect 350540 21422 350592 21428
rect 350552 16574 350580 21422
rect 351932 16574 351960 65554
rect 353312 16574 353340 76638
rect 357532 76628 357584 76634
rect 357532 76570 357584 76576
rect 354680 69080 354732 69086
rect 354680 69022 354732 69028
rect 354692 16574 354720 69022
rect 356058 52048 356114 52057
rect 356058 51983 356114 51992
rect 356072 16574 356100 51983
rect 356704 36712 356756 36718
rect 356704 36654 356756 36660
rect 345032 16546 345336 16574
rect 346412 16546 346992 16574
rect 347792 16546 348096 16574
rect 349172 16546 349292 16574
rect 350552 16546 351224 16574
rect 351932 16546 352880 16574
rect 353312 16546 353616 16574
rect 354692 16546 355272 16574
rect 356072 16546 356376 16574
rect 343364 7812 343416 7818
rect 343364 7754 343416 7760
rect 340972 3392 341024 3398
rect 340972 3334 341024 3340
rect 342168 3392 342220 3398
rect 342168 3334 342220 3340
rect 342904 3392 342956 3398
rect 342904 3334 342956 3340
rect 340892 3182 341012 3210
rect 340984 480 341012 3182
rect 342180 480 342208 3334
rect 343376 480 343404 7754
rect 344560 3392 344612 3398
rect 344560 3334 344612 3340
rect 344572 480 344600 3334
rect 339838 354 339950 480
rect 339512 326 339950 354
rect 339838 -960 339950 326
rect 340942 -960 341054 480
rect 342138 -960 342250 480
rect 343334 -960 343446 480
rect 344530 -960 344642 480
rect 345308 354 345336 16546
rect 346964 480 346992 16546
rect 348068 480 348096 16546
rect 349264 480 349292 16546
rect 350448 6724 350500 6730
rect 350448 6666 350500 6672
rect 350460 480 350488 6666
rect 345726 354 345838 480
rect 345308 326 345838 354
rect 345726 -960 345838 326
rect 346922 -960 347034 480
rect 348026 -960 348138 480
rect 349222 -960 349334 480
rect 350418 -960 350530 480
rect 351196 354 351224 16546
rect 352852 480 352880 16546
rect 351614 354 351726 480
rect 351196 326 351726 354
rect 351614 -960 351726 326
rect 352810 -960 352922 480
rect 353588 354 353616 16546
rect 355244 480 355272 16546
rect 356348 480 356376 16546
rect 356716 3398 356744 36654
rect 356704 3392 356756 3398
rect 356704 3334 356756 3340
rect 357544 480 357572 76570
rect 358832 16574 358860 79358
rect 376760 79348 376812 79354
rect 376760 79290 376812 79296
rect 367100 76560 367152 76566
rect 367100 76502 367152 76508
rect 362958 64288 363014 64297
rect 362958 64223 363014 64232
rect 360200 27124 360252 27130
rect 360200 27066 360252 27072
rect 360212 16574 360240 27066
rect 361580 19984 361632 19990
rect 361580 19926 361632 19932
rect 361592 16574 361620 19926
rect 362972 16574 363000 64223
rect 364982 53408 365038 53417
rect 364982 53343 365038 53352
rect 358832 16546 359504 16574
rect 360212 16546 361160 16574
rect 361592 16546 361896 16574
rect 362972 16546 363552 16574
rect 358728 3392 358780 3398
rect 358728 3334 358780 3340
rect 358740 480 358768 3334
rect 354006 354 354118 480
rect 353588 326 354118 354
rect 354006 -960 354118 326
rect 355202 -960 355314 480
rect 356306 -960 356418 480
rect 357502 -960 357614 480
rect 358698 -960 358810 480
rect 359476 354 359504 16546
rect 361132 480 361160 16546
rect 359894 354 360006 480
rect 359476 326 360006 354
rect 359894 -960 360006 326
rect 361090 -960 361202 480
rect 361868 354 361896 16546
rect 363524 480 363552 16546
rect 364616 16108 364668 16114
rect 364616 16050 364668 16056
rect 364628 480 364656 16050
rect 364996 3398 365024 53343
rect 367112 16574 367140 76502
rect 368480 62144 368532 62150
rect 368480 62086 368532 62092
rect 368492 16574 368520 62086
rect 369858 54904 369914 54913
rect 369858 54839 369914 54848
rect 369872 16574 369900 54839
rect 373998 50416 374054 50425
rect 373998 50351 374054 50360
rect 372620 32496 372672 32502
rect 372620 32438 372672 32444
rect 372632 16574 372660 32438
rect 367112 16546 367784 16574
rect 368492 16546 369440 16574
rect 369872 16546 370176 16574
rect 372632 16546 372936 16574
rect 365812 10464 365864 10470
rect 365812 10406 365864 10412
rect 364984 3392 365036 3398
rect 364984 3334 365036 3340
rect 365824 480 365852 10406
rect 367008 3392 367060 3398
rect 367008 3334 367060 3340
rect 367020 480 367048 3334
rect 362286 354 362398 480
rect 361868 326 362398 354
rect 362286 -960 362398 326
rect 363482 -960 363594 480
rect 364586 -960 364698 480
rect 365782 -960 365894 480
rect 366978 -960 367090 480
rect 367756 354 367784 16546
rect 369412 480 369440 16546
rect 368174 354 368286 480
rect 367756 326 368286 354
rect 368174 -960 368286 326
rect 369370 -960 369482 480
rect 370148 354 370176 16546
rect 371700 4956 371752 4962
rect 371700 4898 371752 4904
rect 371712 480 371740 4898
rect 372908 480 372936 16546
rect 374012 1170 374040 50351
rect 374092 25696 374144 25702
rect 374092 25638 374144 25644
rect 374104 3398 374132 25638
rect 376772 16574 376800 79290
rect 480260 78804 480312 78810
rect 480260 78746 480312 78752
rect 456800 78124 456852 78130
rect 456800 78066 456852 78072
rect 454682 75304 454738 75313
rect 454682 75239 454738 75248
rect 396724 72480 396776 72486
rect 396724 72422 396776 72428
rect 394700 60104 394752 60110
rect 394700 60046 394752 60052
rect 380898 58848 380954 58857
rect 380898 58783 380954 58792
rect 380912 16574 380940 58783
rect 382922 56128 382978 56137
rect 382922 56063 382978 56072
rect 382280 22976 382332 22982
rect 382280 22918 382332 22924
rect 376772 16546 377720 16574
rect 380912 16546 381216 16574
rect 376024 13252 376076 13258
rect 376024 13194 376076 13200
rect 374092 3392 374144 3398
rect 374092 3334 374144 3340
rect 375288 3392 375340 3398
rect 375288 3334 375340 3340
rect 374012 1142 374132 1170
rect 374104 480 374132 1142
rect 375300 480 375328 3334
rect 370566 354 370678 480
rect 370148 326 370678 354
rect 370566 -960 370678 326
rect 371670 -960 371782 480
rect 372866 -960 372978 480
rect 374062 -960 374174 480
rect 375258 -960 375370 480
rect 376036 354 376064 13194
rect 377692 480 377720 16546
rect 378416 13184 378468 13190
rect 378416 13126 378468 13132
rect 376454 354 376566 480
rect 376036 326 376566 354
rect 376454 -960 376566 326
rect 377650 -960 377762 480
rect 378428 354 378456 13126
rect 379980 7744 380032 7750
rect 379980 7686 380032 7692
rect 379992 480 380020 7686
rect 381188 480 381216 16546
rect 382292 3210 382320 22918
rect 382372 14612 382424 14618
rect 382372 14554 382424 14560
rect 382384 3398 382412 14554
rect 382372 3392 382424 3398
rect 382372 3334 382424 3340
rect 382292 3182 382412 3210
rect 382384 480 382412 3182
rect 382936 3126 382964 56063
rect 389180 53100 389232 53106
rect 389180 53042 389232 53048
rect 387798 49192 387854 49201
rect 387798 49127 387854 49136
rect 386420 27056 386472 27062
rect 386420 26998 386472 27004
rect 386432 16574 386460 26998
rect 386432 16546 386736 16574
rect 385960 14544 386012 14550
rect 385960 14486 386012 14492
rect 383568 3392 383620 3398
rect 383568 3334 383620 3340
rect 382924 3120 382976 3126
rect 382924 3062 382976 3068
rect 383580 480 383608 3334
rect 384764 3120 384816 3126
rect 384764 3062 384816 3068
rect 384776 480 384804 3062
rect 385972 480 386000 14486
rect 378846 354 378958 480
rect 378428 326 378958 354
rect 378846 -960 378958 326
rect 379950 -960 380062 480
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384734 -960 384846 480
rect 385930 -960 386042 480
rect 386708 354 386736 16546
rect 387126 354 387238 480
rect 386708 326 387238 354
rect 387812 354 387840 49127
rect 389192 16574 389220 53042
rect 390560 44872 390612 44878
rect 390560 44814 390612 44820
rect 389192 16546 389496 16574
rect 389468 480 389496 16546
rect 390572 3398 390600 44814
rect 390652 31136 390704 31142
rect 390652 31078 390704 31084
rect 390560 3392 390612 3398
rect 390560 3334 390612 3340
rect 390664 480 390692 31078
rect 391940 24268 391992 24274
rect 391940 24210 391992 24216
rect 391952 16574 391980 24210
rect 394712 16574 394740 60046
rect 396080 60036 396132 60042
rect 396080 59978 396132 59984
rect 391952 16546 392624 16574
rect 394712 16546 395384 16574
rect 391848 3392 391900 3398
rect 391848 3334 391900 3340
rect 391860 480 391888 3334
rect 388230 354 388342 480
rect 387812 326 388342 354
rect 387126 -960 387238 326
rect 388230 -960 388342 326
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 392596 354 392624 16546
rect 394240 3936 394292 3942
rect 394240 3878 394292 3884
rect 394252 480 394280 3878
rect 395356 480 395384 16546
rect 393014 354 393126 480
rect 392596 326 393126 354
rect 393014 -960 393126 326
rect 394210 -960 394322 480
rect 395314 -960 395426 480
rect 396092 354 396120 59978
rect 396736 3330 396764 72422
rect 430578 69728 430634 69737
rect 430578 69663 430634 69672
rect 427820 68468 427872 68474
rect 427820 68410 427872 68416
rect 423680 68400 423732 68406
rect 423680 68342 423732 68348
rect 414664 65544 414716 65550
rect 402978 65512 403034 65521
rect 414664 65486 414716 65492
rect 402978 65447 403034 65456
rect 398840 61396 398892 61402
rect 398840 61338 398892 61344
rect 396724 3324 396776 3330
rect 396724 3266 396776 3272
rect 397736 3324 397788 3330
rect 397736 3266 397788 3272
rect 397748 480 397776 3266
rect 398852 3210 398880 61338
rect 400862 51912 400918 51921
rect 400862 51847 400918 51856
rect 398932 29844 398984 29850
rect 398932 29786 398984 29792
rect 398944 3398 398972 29786
rect 400876 3398 400904 51847
rect 402992 16574 403020 65447
rect 412640 62824 412692 62830
rect 412640 62766 412692 62772
rect 405738 47832 405794 47841
rect 405738 47767 405794 47776
rect 404360 22908 404412 22914
rect 404360 22850 404412 22856
rect 402992 16546 403664 16574
rect 401324 3868 401376 3874
rect 401324 3810 401376 3816
rect 398932 3392 398984 3398
rect 398932 3334 398984 3340
rect 400128 3392 400180 3398
rect 400128 3334 400180 3340
rect 400864 3392 400916 3398
rect 400864 3334 400916 3340
rect 398852 3182 398972 3210
rect 398944 480 398972 3182
rect 400140 480 400168 3334
rect 401336 480 401364 3810
rect 402520 3392 402572 3398
rect 402520 3334 402572 3340
rect 402532 480 402560 3334
rect 403636 480 403664 16546
rect 396510 354 396622 480
rect 396092 326 396622 354
rect 396510 -960 396622 326
rect 397706 -960 397818 480
rect 398902 -960 399014 480
rect 400098 -960 400210 480
rect 401294 -960 401406 480
rect 402490 -960 402602 480
rect 403594 -960 403706 480
rect 404372 354 404400 22850
rect 405752 16574 405780 47767
rect 408498 43616 408554 43625
rect 408498 43551 408554 43560
rect 408512 16574 408540 43551
rect 409880 39500 409932 39506
rect 409880 39442 409932 39448
rect 409892 16574 409920 39442
rect 411260 18760 411312 18766
rect 411260 18702 411312 18708
rect 411272 16574 411300 18702
rect 405752 16546 406056 16574
rect 408512 16546 409184 16574
rect 409892 16546 410840 16574
rect 411272 16546 411944 16574
rect 406028 480 406056 16546
rect 407212 11892 407264 11898
rect 407212 11834 407264 11840
rect 407224 480 407252 11834
rect 408408 3800 408460 3806
rect 408408 3742 408460 3748
rect 408420 480 408448 3742
rect 404790 354 404902 480
rect 404372 326 404902 354
rect 404790 -960 404902 326
rect 405986 -960 406098 480
rect 407182 -960 407294 480
rect 408378 -960 408490 480
rect 409156 354 409184 16546
rect 410812 480 410840 16546
rect 411916 480 411944 16546
rect 409574 354 409686 480
rect 409156 326 409686 354
rect 409574 -960 409686 326
rect 410770 -960 410882 480
rect 411874 -960 411986 480
rect 412652 354 412680 62766
rect 414296 9104 414348 9110
rect 414296 9046 414348 9052
rect 414308 480 414336 9046
rect 414676 3398 414704 65486
rect 418802 57216 418858 57225
rect 418802 57151 418858 57160
rect 418160 21412 418212 21418
rect 418160 21354 418212 21360
rect 418172 16574 418200 21354
rect 418172 16546 418568 16574
rect 417424 16040 417476 16046
rect 417424 15982 417476 15988
rect 415492 3732 415544 3738
rect 415492 3674 415544 3680
rect 414664 3392 414716 3398
rect 414664 3334 414716 3340
rect 415504 480 415532 3674
rect 416688 3392 416740 3398
rect 416688 3334 416740 3340
rect 416700 480 416728 3334
rect 413070 354 413182 480
rect 412652 326 413182 354
rect 413070 -960 413182 326
rect 414266 -960 414378 480
rect 415462 -960 415574 480
rect 416658 -960 416770 480
rect 417436 354 417464 15982
rect 417854 354 417966 480
rect 417436 326 417966 354
rect 418540 354 418568 16546
rect 418816 3398 418844 57151
rect 420920 28416 420972 28422
rect 420920 28358 420972 28364
rect 418804 3392 418856 3398
rect 418804 3334 418856 3340
rect 420184 3392 420236 3398
rect 420184 3334 420236 3340
rect 420196 480 420224 3334
rect 418958 354 419070 480
rect 418540 326 419070 354
rect 417854 -960 417966 326
rect 418958 -960 419070 326
rect 420154 -960 420266 480
rect 420932 354 420960 28358
rect 422576 6656 422628 6662
rect 422576 6598 422628 6604
rect 422588 480 422616 6598
rect 423692 3398 423720 68342
rect 423770 46200 423826 46209
rect 423770 46135 423826 46144
rect 423680 3392 423732 3398
rect 423680 3334 423732 3340
rect 423784 480 423812 46135
rect 426440 42220 426492 42226
rect 426440 42162 426492 42168
rect 425058 35184 425114 35193
rect 425058 35119 425114 35128
rect 425072 16574 425100 35119
rect 426452 16574 426480 42162
rect 427832 16574 427860 68410
rect 430592 16574 430620 69663
rect 446402 62792 446458 62801
rect 446402 62727 446458 62736
rect 432602 54768 432658 54777
rect 432602 54703 432658 54712
rect 431960 33924 432012 33930
rect 431960 33866 432012 33872
rect 425072 16546 425744 16574
rect 426452 16546 426848 16574
rect 427832 16546 428504 16574
rect 430592 16546 430896 16574
rect 424968 3392 425020 3398
rect 424968 3334 425020 3340
rect 424980 480 425008 3334
rect 421350 354 421462 480
rect 420932 326 421462 354
rect 421350 -960 421462 326
rect 422546 -960 422658 480
rect 423742 -960 423854 480
rect 424938 -960 425050 480
rect 425716 354 425744 16546
rect 426134 354 426246 480
rect 425716 326 426246 354
rect 426820 354 426848 16546
rect 428476 480 428504 16546
rect 429660 6588 429712 6594
rect 429660 6530 429712 6536
rect 429672 480 429700 6530
rect 430868 480 430896 16546
rect 431972 3330 432000 33866
rect 432052 10396 432104 10402
rect 432052 10338 432104 10344
rect 431960 3324 432012 3330
rect 431960 3266 432012 3272
rect 432064 480 432092 10338
rect 432616 3398 432644 54703
rect 437478 53272 437534 53281
rect 437478 53207 437534 53216
rect 435548 7676 435600 7682
rect 435548 7618 435600 7624
rect 432604 3392 432656 3398
rect 432604 3334 432656 3340
rect 434444 3392 434496 3398
rect 434444 3334 434496 3340
rect 433248 3324 433300 3330
rect 433248 3266 433300 3272
rect 433260 480 433288 3266
rect 434456 480 434484 3334
rect 435560 480 435588 7618
rect 436744 6520 436796 6526
rect 436744 6462 436796 6468
rect 436756 480 436784 6462
rect 427238 354 427350 480
rect 426820 326 427350 354
rect 426134 -960 426246 326
rect 427238 -960 427350 326
rect 428434 -960 428546 480
rect 429630 -960 429742 480
rect 430826 -960 430938 480
rect 432022 -960 432134 480
rect 433218 -960 433330 480
rect 434414 -960 434526 480
rect 435518 -960 435630 480
rect 436714 -960 436826 480
rect 437492 354 437520 53207
rect 440238 45112 440294 45121
rect 440238 45047 440294 45056
rect 438860 32428 438912 32434
rect 438860 32370 438912 32376
rect 438872 16574 438900 32370
rect 438872 16546 439176 16574
rect 439148 480 439176 16546
rect 440252 3398 440280 45047
rect 444380 40860 444432 40866
rect 444380 40802 444432 40808
rect 444392 16574 444420 40802
rect 445760 17400 445812 17406
rect 445760 17342 445812 17348
rect 444392 16546 445064 16574
rect 440332 15972 440384 15978
rect 440332 15914 440384 15920
rect 440240 3392 440292 3398
rect 440240 3334 440292 3340
rect 440344 480 440372 15914
rect 443828 6452 443880 6458
rect 443828 6394 443880 6400
rect 442632 6316 442684 6322
rect 442632 6258 442684 6264
rect 441528 3392 441580 3398
rect 441528 3334 441580 3340
rect 441540 480 441568 3334
rect 442644 480 442672 6258
rect 443840 480 443868 6394
rect 445036 480 445064 16546
rect 437910 354 438022 480
rect 437492 326 438022 354
rect 437910 -960 438022 326
rect 439106 -960 439218 480
rect 440302 -960 440414 480
rect 441498 -960 441610 480
rect 442602 -960 442714 480
rect 443798 -960 443910 480
rect 444994 -960 445106 480
rect 445772 354 445800 17342
rect 446416 3398 446444 62727
rect 448518 58712 448574 58721
rect 448518 58647 448574 58656
rect 446404 3392 446456 3398
rect 446404 3334 446456 3340
rect 447416 3392 447468 3398
rect 447416 3334 447468 3340
rect 447428 480 447456 3334
rect 448532 3210 448560 58647
rect 450542 55992 450598 56001
rect 450542 55927 450598 55936
rect 448612 17332 448664 17338
rect 448612 17274 448664 17280
rect 448624 3398 448652 17274
rect 450556 4146 450584 55927
rect 452660 42152 452712 42158
rect 452660 42094 452712 42100
rect 452672 16574 452700 42094
rect 452672 16546 453344 16574
rect 450912 6384 450964 6390
rect 450912 6326 450964 6332
rect 450544 4140 450596 4146
rect 450544 4082 450596 4088
rect 448612 3392 448664 3398
rect 448612 3334 448664 3340
rect 449808 3392 449860 3398
rect 449808 3334 449860 3340
rect 448532 3182 448652 3210
rect 448624 480 448652 3182
rect 449820 480 449848 3334
rect 450924 480 450952 6326
rect 452108 4140 452160 4146
rect 452108 4082 452160 4088
rect 452120 480 452148 4082
rect 453316 480 453344 16546
rect 454040 11824 454092 11830
rect 454040 11766 454092 11772
rect 446190 354 446302 480
rect 445772 326 446302 354
rect 446190 -960 446302 326
rect 447386 -960 447498 480
rect 448582 -960 448694 480
rect 449778 -960 449890 480
rect 450882 -960 450994 480
rect 452078 -960 452190 480
rect 453274 -960 453386 480
rect 454052 354 454080 11766
rect 454696 3738 454724 75239
rect 455420 49088 455472 49094
rect 455420 49030 455472 49036
rect 455432 16574 455460 49030
rect 455432 16546 455736 16574
rect 454684 3732 454736 3738
rect 454684 3674 454736 3680
rect 455708 480 455736 16546
rect 456812 3398 456840 78066
rect 465172 78056 465224 78062
rect 465172 77998 465224 78004
rect 459558 61568 459614 61577
rect 459558 61503 459614 61512
rect 458180 43444 458232 43450
rect 458180 43386 458232 43392
rect 458192 16574 458220 43386
rect 459572 16574 459600 61503
rect 464344 51740 464396 51746
rect 464344 51682 464396 51688
rect 462320 39432 462372 39438
rect 462320 39374 462372 39380
rect 458192 16546 459232 16574
rect 459572 16546 459968 16574
rect 456892 4888 456944 4894
rect 456892 4830 456944 4836
rect 456800 3392 456852 3398
rect 456800 3334 456852 3340
rect 456904 480 456932 4830
rect 458088 3392 458140 3398
rect 458088 3334 458140 3340
rect 458100 480 458128 3334
rect 459204 480 459232 16546
rect 454470 354 454582 480
rect 454052 326 454582 354
rect 454470 -960 454582 326
rect 455666 -960 455778 480
rect 456862 -960 456974 480
rect 458058 -960 458170 480
rect 459162 -960 459274 480
rect 459940 354 459968 16546
rect 461584 3664 461636 3670
rect 461584 3606 461636 3612
rect 461596 480 461624 3606
rect 460358 354 460470 480
rect 459940 326 460470 354
rect 460358 -960 460470 326
rect 461554 -960 461666 480
rect 462332 354 462360 39374
rect 463700 38072 463752 38078
rect 463700 38014 463752 38020
rect 463712 16574 463740 38014
rect 463712 16546 464016 16574
rect 463988 480 464016 16546
rect 464356 3058 464384 51682
rect 464344 3052 464396 3058
rect 464344 2994 464396 3000
rect 465184 480 465212 77998
rect 471980 77988 472032 77994
rect 471980 77930 472032 77936
rect 468482 47696 468538 47705
rect 468482 47631 468538 47640
rect 466460 46980 466512 46986
rect 466460 46922 466512 46928
rect 466472 16574 466500 46922
rect 466472 16546 467512 16574
rect 466276 3052 466328 3058
rect 466276 2994 466328 3000
rect 466288 480 466316 2994
rect 467484 480 467512 16546
rect 468496 3602 468524 47631
rect 470600 31068 470652 31074
rect 470600 31010 470652 31016
rect 468300 3596 468352 3602
rect 468300 3538 468352 3544
rect 468484 3596 468536 3602
rect 468484 3538 468536 3544
rect 469864 3596 469916 3602
rect 469864 3538 469916 3544
rect 462750 354 462862 480
rect 462332 326 462862 354
rect 462750 -960 462862 326
rect 463946 -960 464058 480
rect 465142 -960 465254 480
rect 466246 -960 466358 480
rect 467442 -960 467554 480
rect 468312 354 468340 3538
rect 469876 480 469904 3538
rect 468638 354 468750 480
rect 468312 326 468750 354
rect 468638 -960 468750 326
rect 469834 -960 469946 480
rect 470612 354 470640 31010
rect 471992 16574 472020 77930
rect 478144 75336 478196 75342
rect 478144 75278 478196 75284
rect 472624 64184 472676 64190
rect 472624 64126 472676 64132
rect 471992 16546 472296 16574
rect 472268 480 472296 16546
rect 472636 3534 472664 64126
rect 473452 56704 473504 56710
rect 473452 56646 473504 56652
rect 473464 16574 473492 56646
rect 474738 53136 474794 53145
rect 474738 53071 474794 53080
rect 474752 16574 474780 53071
rect 476120 38004 476172 38010
rect 476120 37946 476172 37952
rect 476132 16574 476160 37946
rect 477500 17264 477552 17270
rect 477500 17206 477552 17212
rect 473464 16546 474136 16574
rect 474752 16546 475792 16574
rect 476132 16546 476528 16574
rect 472624 3528 472676 3534
rect 472624 3470 472676 3476
rect 473452 3528 473504 3534
rect 473452 3470 473504 3476
rect 473464 480 473492 3470
rect 471030 354 471142 480
rect 470612 326 471142 354
rect 471030 -960 471142 326
rect 472226 -960 472338 480
rect 473422 -960 473534 480
rect 474108 354 474136 16546
rect 475764 480 475792 16546
rect 474526 354 474638 480
rect 474108 326 474638 354
rect 474526 -960 474638 326
rect 475722 -960 475834 480
rect 476500 354 476528 16546
rect 477512 6914 477540 17206
rect 478156 16574 478184 75278
rect 480272 16574 480300 78746
rect 500958 78160 501014 78169
rect 500958 78095 501014 78104
rect 498198 71360 498254 71369
rect 498198 71295 498254 71304
rect 494060 66428 494112 66434
rect 494060 66370 494112 66376
rect 484398 59936 484454 59945
rect 484398 59871 484454 59880
rect 482282 55856 482338 55865
rect 482282 55791 482338 55800
rect 481640 36644 481692 36650
rect 481640 36586 481692 36592
rect 481652 16574 481680 36586
rect 478156 16546 478276 16574
rect 480272 16546 480576 16574
rect 481652 16546 481772 16574
rect 477512 6886 478184 6914
rect 478156 480 478184 6886
rect 478248 3602 478276 16546
rect 478236 3596 478288 3602
rect 478236 3538 478288 3544
rect 479340 3528 479392 3534
rect 479340 3470 479392 3476
rect 479352 480 479380 3470
rect 480548 480 480576 16546
rect 481744 480 481772 16546
rect 482192 13116 482244 13122
rect 482192 13058 482244 13064
rect 482204 490 482232 13058
rect 482296 3398 482324 55791
rect 484412 16574 484440 59871
rect 489918 49056 489974 49065
rect 489918 48991 489974 49000
rect 488540 35352 488592 35358
rect 488540 35294 488592 35300
rect 488552 16574 488580 35294
rect 484412 16546 484808 16574
rect 488552 16546 488856 16574
rect 482284 3392 482336 3398
rect 482284 3334 482336 3340
rect 484032 3392 484084 3398
rect 484032 3334 484084 3340
rect 476918 354 477030 480
rect 476500 326 477030 354
rect 476918 -960 477030 326
rect 478114 -960 478226 480
rect 479310 -960 479422 480
rect 480506 -960 480618 480
rect 481702 -960 481814 480
rect 482204 462 482416 490
rect 484044 480 484072 3334
rect 482388 354 482416 462
rect 482806 354 482918 480
rect 482388 326 482918 354
rect 482806 -960 482918 326
rect 484002 -960 484114 480
rect 484780 354 484808 16546
rect 486424 14476 486476 14482
rect 486424 14418 486476 14424
rect 486436 480 486464 14418
rect 487620 3460 487672 3466
rect 487620 3402 487672 3408
rect 487632 480 487660 3402
rect 488828 480 488856 16546
rect 489932 480 489960 48991
rect 490010 47560 490066 47569
rect 490010 47495 490066 47504
rect 490024 16574 490052 47495
rect 491300 29776 491352 29782
rect 491300 29718 491352 29724
rect 491312 16574 491340 29718
rect 492680 26988 492732 26994
rect 492680 26930 492732 26936
rect 492692 16574 492720 26930
rect 494072 16574 494100 66370
rect 495440 42084 495492 42090
rect 495440 42026 495492 42032
rect 490024 16546 490696 16574
rect 491312 16546 492352 16574
rect 492692 16546 493088 16574
rect 494072 16546 494744 16574
rect 485198 354 485310 480
rect 484780 326 485310 354
rect 485198 -960 485310 326
rect 486394 -960 486506 480
rect 487590 -960 487702 480
rect 488786 -960 488898 480
rect 489890 -960 490002 480
rect 490668 354 490696 16546
rect 492324 480 492352 16546
rect 491086 354 491198 480
rect 490668 326 491198 354
rect 491086 -960 491198 326
rect 492282 -960 492394 480
rect 493060 354 493088 16546
rect 494716 480 494744 16546
rect 493478 354 493590 480
rect 493060 326 493590 354
rect 493478 -960 493590 326
rect 494674 -960 494786 480
rect 495452 354 495480 42026
rect 497096 3732 497148 3738
rect 497096 3674 497148 3680
rect 497108 480 497136 3674
rect 498212 480 498240 71295
rect 498292 40792 498344 40798
rect 498292 40734 498344 40740
rect 498304 16574 498332 40734
rect 500972 16574 501000 78095
rect 503720 36576 503772 36582
rect 503720 36518 503772 36524
rect 502340 28348 502392 28354
rect 502340 28290 502392 28296
rect 502352 16574 502380 28290
rect 498304 16546 498976 16574
rect 500972 16546 501368 16574
rect 502352 16546 503024 16574
rect 495870 354 495982 480
rect 495452 326 495982 354
rect 495870 -960 495982 326
rect 497066 -960 497178 480
rect 498170 -960 498282 480
rect 498948 354 498976 16546
rect 500592 3596 500644 3602
rect 500592 3538 500644 3544
rect 500604 480 500632 3538
rect 499366 354 499478 480
rect 498948 326 499478 354
rect 499366 -960 499478 326
rect 500562 -960 500674 480
rect 501340 354 501368 16546
rect 502996 480 503024 16546
rect 501758 354 501870 480
rect 501340 326 501870 354
rect 501758 -960 501870 326
rect 502954 -960 503066 480
rect 503732 354 503760 36518
rect 505112 16574 505140 80679
rect 523132 80096 523184 80102
rect 523132 80038 523184 80044
rect 506480 75268 506532 75274
rect 506480 75210 506532 75216
rect 505112 16546 505416 16574
rect 505388 480 505416 16546
rect 506492 3534 506520 75210
rect 517520 75200 517572 75206
rect 517520 75142 517572 75148
rect 521658 75168 521714 75177
rect 511264 74588 511316 74594
rect 511264 74530 511316 74536
rect 507858 54632 507914 54641
rect 507858 54567 507914 54576
rect 506572 26920 506624 26926
rect 506572 26862 506624 26868
rect 506480 3528 506532 3534
rect 506480 3470 506532 3476
rect 506584 3346 506612 26862
rect 507872 16574 507900 54567
rect 509240 25628 509292 25634
rect 509240 25570 509292 25576
rect 509252 16574 509280 25570
rect 510620 25560 510672 25566
rect 510620 25502 510672 25508
rect 507872 16546 508912 16574
rect 509252 16546 509648 16574
rect 507308 3528 507360 3534
rect 507308 3470 507360 3476
rect 506492 3318 506612 3346
rect 506492 480 506520 3318
rect 504150 354 504262 480
rect 503732 326 504262 354
rect 504150 -960 504262 326
rect 505346 -960 505458 480
rect 506450 -960 506562 480
rect 507320 354 507348 3470
rect 508884 480 508912 16546
rect 507646 354 507758 480
rect 507320 326 507758 354
rect 507646 -960 507758 326
rect 508842 -960 508954 480
rect 509620 354 509648 16546
rect 510632 6914 510660 25502
rect 511276 16574 511304 74530
rect 511998 64152 512054 64161
rect 511998 64087 512054 64096
rect 511276 16546 511396 16574
rect 510632 6886 511304 6914
rect 511276 480 511304 6886
rect 511368 3466 511396 16546
rect 511356 3460 511408 3466
rect 511356 3402 511408 3408
rect 510038 354 510150 480
rect 509620 326 510150 354
rect 510038 -960 510150 326
rect 511234 -960 511346 480
rect 512012 354 512040 64087
rect 514022 58576 514078 58585
rect 514022 58511 514078 58520
rect 513380 24200 513432 24206
rect 513380 24142 513432 24148
rect 512430 354 512542 480
rect 512012 326 512542 354
rect 513392 354 513420 24142
rect 514036 3534 514064 58511
rect 516140 49020 516192 49026
rect 516140 48962 516192 48968
rect 516152 16574 516180 48962
rect 517532 16574 517560 75142
rect 521658 75103 521714 75112
rect 520922 44976 520978 44985
rect 520922 44911 520978 44920
rect 518900 28280 518952 28286
rect 518900 28222 518952 28228
rect 518912 16574 518940 28222
rect 520280 22840 520332 22846
rect 520280 22782 520332 22788
rect 516152 16546 517192 16574
rect 517532 16546 517928 16574
rect 518912 16546 519584 16574
rect 514024 3528 514076 3534
rect 514024 3470 514076 3476
rect 515956 3528 516008 3534
rect 515956 3470 516008 3476
rect 514760 3460 514812 3466
rect 514760 3402 514812 3408
rect 514772 480 514800 3402
rect 515968 480 515996 3470
rect 517164 480 517192 16546
rect 513534 354 513646 480
rect 513392 326 513646 354
rect 512430 -960 512542 326
rect 513534 -960 513646 326
rect 514730 -960 514842 480
rect 515926 -960 516038 480
rect 517122 -960 517234 480
rect 517900 354 517928 16546
rect 519556 480 519584 16546
rect 518318 354 518430 480
rect 517900 326 518430 354
rect 518318 -960 518430 326
rect 519514 -960 519626 480
rect 520292 354 520320 22782
rect 520936 3330 520964 44911
rect 520924 3324 520976 3330
rect 520924 3266 520976 3272
rect 520710 354 520822 480
rect 520292 326 520822 354
rect 521672 354 521700 75103
rect 523144 6914 523172 80038
rect 539692 78736 539744 78742
rect 539692 78678 539744 78684
rect 531318 71224 531374 71233
rect 531318 71159 531374 71168
rect 529940 66360 529992 66366
rect 529940 66302 529992 66308
rect 525800 64932 525852 64938
rect 525800 64874 525852 64880
rect 525064 37936 525116 37942
rect 525064 37878 525116 37884
rect 524420 22772 524472 22778
rect 524420 22714 524472 22720
rect 524432 16574 524460 22714
rect 524432 16546 525012 16574
rect 523052 6886 523172 6914
rect 523052 480 523080 6886
rect 524984 3482 525012 16546
rect 525076 3602 525104 37878
rect 525812 16574 525840 64874
rect 527824 60784 527876 60790
rect 527824 60726 527876 60732
rect 527836 16574 527864 60726
rect 528558 44840 528614 44849
rect 528558 44775 528614 44784
rect 525812 16546 526208 16574
rect 527836 16546 527956 16574
rect 525064 3596 525116 3602
rect 525064 3538 525116 3544
rect 524984 3454 525472 3482
rect 524236 3324 524288 3330
rect 524236 3266 524288 3272
rect 524248 480 524276 3266
rect 525444 480 525472 3454
rect 521814 354 521926 480
rect 521672 326 521926 354
rect 520710 -960 520822 326
rect 521814 -960 521926 326
rect 523010 -960 523122 480
rect 524206 -960 524318 480
rect 525402 -960 525514 480
rect 526180 354 526208 16546
rect 527824 3596 527876 3602
rect 527824 3538 527876 3544
rect 527836 480 527864 3538
rect 527928 3466 527956 16546
rect 527916 3460 527968 3466
rect 527916 3402 527968 3408
rect 526598 354 526710 480
rect 526180 326 526710 354
rect 526598 -960 526710 326
rect 527794 -960 527906 480
rect 528572 354 528600 44775
rect 528990 354 529102 480
rect 528572 326 529102 354
rect 529952 354 529980 66302
rect 531332 480 531360 71159
rect 536840 68332 536892 68338
rect 536840 68274 536892 68280
rect 534722 43480 534778 43489
rect 534722 43415 534778 43424
rect 534078 36544 534134 36553
rect 534078 36479 534134 36488
rect 531412 24132 531464 24138
rect 531412 24074 531464 24080
rect 531424 16574 531452 24074
rect 534092 16574 534120 36479
rect 531424 16546 532096 16574
rect 534092 16546 534488 16574
rect 530094 354 530206 480
rect 529952 326 530206 354
rect 528990 -960 529102 326
rect 530094 -960 530206 326
rect 531290 -960 531402 480
rect 532068 354 532096 16546
rect 533712 3460 533764 3466
rect 533712 3402 533764 3408
rect 533724 480 533752 3402
rect 532486 354 532598 480
rect 532068 326 532598 354
rect 532486 -960 532598 326
rect 533682 -960 533794 480
rect 534460 354 534488 16546
rect 534736 3398 534764 43415
rect 535460 40724 535512 40730
rect 535460 40666 535512 40672
rect 535472 16574 535500 40666
rect 536852 16574 536880 68274
rect 538864 35284 538916 35290
rect 538864 35226 538916 35232
rect 535472 16546 536144 16574
rect 536852 16546 537248 16574
rect 534724 3392 534776 3398
rect 534724 3334 534776 3340
rect 536116 480 536144 16546
rect 537220 480 537248 16546
rect 538404 7608 538456 7614
rect 538404 7550 538456 7556
rect 538416 480 538444 7550
rect 538876 3534 538904 35226
rect 539704 16574 539732 78678
rect 566462 76528 566518 76537
rect 566462 76463 566518 76472
rect 549902 71088 549958 71097
rect 549902 71023 549958 71032
rect 543740 63572 543792 63578
rect 543740 63514 543792 63520
rect 542358 51776 542414 51785
rect 542358 51711 542414 51720
rect 542372 16574 542400 51711
rect 543752 16574 543780 63514
rect 545120 57248 545172 57254
rect 545120 57190 545172 57196
rect 545132 16574 545160 57190
rect 547878 48920 547934 48929
rect 547878 48855 547934 48864
rect 539704 16546 540376 16574
rect 542372 16546 542768 16574
rect 543752 16546 544424 16574
rect 545132 16546 545528 16574
rect 538864 3528 538916 3534
rect 538864 3470 538916 3476
rect 539600 3528 539652 3534
rect 539600 3470 539652 3476
rect 539612 480 539640 3470
rect 534878 354 534990 480
rect 534460 326 534990 354
rect 534878 -960 534990 326
rect 536074 -960 536186 480
rect 537178 -960 537290 480
rect 538374 -960 538486 480
rect 539570 -960 539682 480
rect 540348 354 540376 16546
rect 541992 4820 542044 4826
rect 541992 4762 542044 4768
rect 542004 480 542032 4762
rect 540766 354 540878 480
rect 540348 326 540878 354
rect 540766 -960 540878 326
rect 541962 -960 542074 480
rect 542740 354 542768 16546
rect 544396 480 544424 16546
rect 545500 480 545528 16546
rect 546500 15904 546552 15910
rect 546500 15846 546552 15852
rect 543158 354 543270 480
rect 542740 326 543270 354
rect 543158 -960 543270 326
rect 544354 -960 544466 480
rect 545458 -960 545570 480
rect 546512 354 546540 15846
rect 547892 480 547920 48855
rect 548616 10328 548668 10334
rect 548616 10270 548668 10276
rect 546654 354 546766 480
rect 546512 326 546766 354
rect 546654 -960 546766 326
rect 547850 -960 547962 480
rect 548628 354 548656 10270
rect 549916 3534 549944 71023
rect 557538 69592 557594 69601
rect 557538 69527 557594 69536
rect 554044 66292 554096 66298
rect 554044 66234 554096 66240
rect 552020 35216 552072 35222
rect 552020 35158 552072 35164
rect 552032 16574 552060 35158
rect 553400 29708 553452 29714
rect 553400 29650 553452 29656
rect 553412 16574 553440 29650
rect 552032 16546 552704 16574
rect 553412 16546 553808 16574
rect 549904 3528 549956 3534
rect 549904 3470 549956 3476
rect 551468 3528 551520 3534
rect 551468 3470 551520 3476
rect 550272 3392 550324 3398
rect 550272 3334 550324 3340
rect 550284 480 550312 3334
rect 551480 480 551508 3470
rect 552676 480 552704 16546
rect 553780 480 553808 16546
rect 554056 3534 554084 66234
rect 556158 50280 556214 50289
rect 556158 50215 556214 50224
rect 556172 16574 556200 50215
rect 557552 16574 557580 69527
rect 563702 61432 563758 61441
rect 563702 61367 563758 61376
rect 560942 54496 560998 54505
rect 560942 54431 560998 54440
rect 558920 33856 558972 33862
rect 558920 33798 558972 33804
rect 558932 16574 558960 33798
rect 556172 16546 556936 16574
rect 557552 16546 558592 16574
rect 558932 16546 559328 16574
rect 556160 8968 556212 8974
rect 556160 8910 556212 8916
rect 554044 3528 554096 3534
rect 554044 3470 554096 3476
rect 554964 3528 555016 3534
rect 554964 3470 555016 3476
rect 554976 480 555004 3470
rect 556172 480 556200 8910
rect 549046 354 549158 480
rect 548628 326 549158 354
rect 549046 -960 549158 326
rect 550242 -960 550354 480
rect 551438 -960 551550 480
rect 552634 -960 552746 480
rect 553738 -960 553850 480
rect 554934 -960 555046 480
rect 556130 -960 556242 480
rect 556908 354 556936 16546
rect 558564 480 558592 16546
rect 557326 354 557438 480
rect 556908 326 557438 354
rect 557326 -960 557438 326
rect 558522 -960 558634 480
rect 559300 354 559328 16546
rect 560392 11756 560444 11762
rect 560392 11698 560444 11704
rect 559718 354 559830 480
rect 559300 326 559830 354
rect 560404 354 560432 11698
rect 560956 3602 560984 54431
rect 562324 39364 562376 39370
rect 562324 39306 562376 39312
rect 562048 9036 562100 9042
rect 562048 8978 562100 8984
rect 560944 3596 560996 3602
rect 560944 3538 560996 3544
rect 562060 480 562088 8978
rect 562336 3330 562364 39306
rect 563244 6248 563296 6254
rect 563244 6190 563296 6196
rect 562324 3324 562376 3330
rect 562324 3266 562376 3272
rect 563256 480 563284 6190
rect 563716 3534 563744 61367
rect 566476 4078 566504 76463
rect 580172 73160 580224 73166
rect 580172 73102 580224 73108
rect 580184 73001 580212 73102
rect 580170 72992 580226 73001
rect 580170 72927 580226 72936
rect 574742 68232 574798 68241
rect 574742 68167 574798 68176
rect 567844 56636 567896 56642
rect 567844 56578 567896 56584
rect 566464 4072 566516 4078
rect 566464 4014 566516 4020
rect 564440 3596 564492 3602
rect 564440 3538 564492 3544
rect 563704 3528 563756 3534
rect 563704 3470 563756 3476
rect 564452 480 564480 3538
rect 565636 3528 565688 3534
rect 565636 3470 565688 3476
rect 565648 480 565676 3470
rect 567856 3466 567884 56578
rect 569960 50380 570012 50386
rect 569960 50322 570012 50328
rect 567936 29640 567988 29646
rect 567936 29582 567988 29588
rect 567948 3534 567976 29582
rect 569972 16574 570000 50322
rect 571984 45620 572036 45626
rect 571984 45562 572036 45568
rect 571340 18692 571392 18698
rect 571340 18634 571392 18640
rect 569972 16546 570368 16574
rect 568028 4072 568080 4078
rect 568028 4014 568080 4020
rect 567936 3528 567988 3534
rect 567936 3470 567988 3476
rect 567844 3460 567896 3466
rect 567844 3402 567896 3408
rect 566832 3324 566884 3330
rect 566832 3266 566884 3272
rect 566844 480 566872 3266
rect 568040 480 568068 4014
rect 569132 3528 569184 3534
rect 569132 3470 569184 3476
rect 569144 480 569172 3470
rect 570340 480 570368 16546
rect 560822 354 560934 480
rect 560404 326 560934 354
rect 559718 -960 559830 326
rect 560822 -960 560934 326
rect 562018 -960 562130 480
rect 563214 -960 563326 480
rect 564410 -960 564522 480
rect 565606 -960 565718 480
rect 566802 -960 566914 480
rect 567998 -960 568110 480
rect 569102 -960 569214 480
rect 570298 -960 570410 480
rect 571352 354 571380 18634
rect 571996 3330 572024 45562
rect 574100 18624 574152 18630
rect 574100 18566 574152 18572
rect 574112 16574 574140 18566
rect 574112 16546 574692 16574
rect 574664 3482 574692 16546
rect 574756 3602 574784 68167
rect 576860 42832 576912 42838
rect 576860 42774 576912 42780
rect 576872 16574 576900 42774
rect 578240 33788 578292 33794
rect 578240 33730 578292 33736
rect 578252 16574 578280 33730
rect 576872 16546 576992 16574
rect 578252 16546 578648 16574
rect 574744 3596 574796 3602
rect 574744 3538 574796 3544
rect 576308 3596 576360 3602
rect 576308 3538 576360 3544
rect 572720 3460 572772 3466
rect 574664 3454 575152 3482
rect 572720 3402 572772 3408
rect 571984 3324 572036 3330
rect 571984 3266 572036 3272
rect 572732 480 572760 3402
rect 573916 3324 573968 3330
rect 573916 3266 573968 3272
rect 573928 480 573956 3266
rect 575124 480 575152 3454
rect 576320 480 576348 3538
rect 571494 354 571606 480
rect 571352 326 571606 354
rect 571494 -960 571606 326
rect 572690 -960 572802 480
rect 573886 -960 573998 480
rect 575082 -960 575194 480
rect 576278 -960 576390 480
rect 576964 354 576992 16546
rect 578620 480 578648 16546
rect 580276 6633 580304 150447
rect 580540 149116 580592 149122
rect 580540 149058 580592 149064
rect 580448 147688 580500 147694
rect 580448 147630 580500 147636
rect 580354 143576 580410 143585
rect 580354 143511 580410 143520
rect 580368 19825 580396 143511
rect 580460 33153 580488 147630
rect 580552 46345 580580 149058
rect 580724 142520 580776 142526
rect 580724 142462 580776 142468
rect 580630 140856 580686 140865
rect 580630 140791 580686 140800
rect 580644 59673 580672 140791
rect 580736 99521 580764 142462
rect 580908 142248 580960 142254
rect 580908 142190 580960 142196
rect 580816 140820 580868 140826
rect 580816 140762 580868 140768
rect 580828 112849 580856 140762
rect 580920 126041 580948 142190
rect 580906 126032 580962 126041
rect 580906 125967 580962 125976
rect 580814 112840 580870 112849
rect 580814 112775 580870 112784
rect 580722 99512 580778 99521
rect 580722 99447 580778 99456
rect 581090 78024 581146 78033
rect 581090 77959 581146 77968
rect 580998 77888 581054 77897
rect 580998 77823 581054 77832
rect 580630 59664 580686 59673
rect 580630 59599 580686 59608
rect 580538 46336 580594 46345
rect 580538 46271 580594 46280
rect 580446 33144 580502 33153
rect 580446 33079 580502 33088
rect 580354 19816 580410 19825
rect 580354 19751 580410 19760
rect 580262 6624 580318 6633
rect 580262 6559 580318 6568
rect 581012 480 581040 77823
rect 581104 16574 581132 77959
rect 581104 16546 581776 16574
rect 577382 354 577494 480
rect 576964 326 577494 354
rect 577382 -960 577494 326
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 581748 354 581776 16546
rect 583392 6180 583444 6186
rect 583392 6122 583444 6128
rect 583404 480 583432 6122
rect 582166 354 582278 480
rect 581748 326 582278 354
rect 582166 -960 582278 326
rect 583362 -960 583474 480
<< via2 >>
rect 3422 684256 3478 684312
rect 3514 671200 3570 671256
rect 3422 658144 3478 658200
rect 3422 632068 3424 632088
rect 3424 632068 3476 632088
rect 3476 632068 3478 632088
rect 3422 632032 3478 632068
rect 3146 619112 3202 619168
rect 3238 606056 3294 606112
rect 3330 579944 3386 580000
rect 3422 566888 3478 566944
rect 3422 553832 3478 553888
rect 3422 527856 3478 527912
rect 3422 514820 3478 514856
rect 3422 514800 3424 514820
rect 3424 514800 3476 514820
rect 3476 514800 3478 514820
rect 3054 501744 3110 501800
rect 3422 475632 3478 475688
rect 3146 449520 3202 449576
rect 2870 410488 2926 410544
rect 2778 371340 2834 371376
rect 2778 371320 2780 371340
rect 2780 371320 2832 371340
rect 2832 371320 2834 371340
rect 3146 358400 3202 358456
rect 3330 319232 3386 319288
rect 3054 267144 3110 267200
rect 3514 462576 3570 462632
rect 3514 423544 3570 423600
rect 3514 397468 3516 397488
rect 3516 397468 3568 397488
rect 3568 397468 3570 397488
rect 3514 397432 3570 397468
rect 3514 345344 3570 345400
rect 3514 306176 3570 306232
rect 3514 293120 3570 293176
rect 2778 241032 2834 241088
rect 3514 254088 3570 254144
rect 3514 214920 3570 214976
rect 3422 201864 3478 201920
rect 101770 197920 101826 197976
rect 3422 188808 3478 188864
rect 3514 162832 3570 162888
rect 3146 149776 3202 149832
rect 3238 136720 3294 136776
rect 3054 110608 3110 110664
rect 2778 77832 2834 77888
rect 2870 62736 2926 62792
rect 6918 77968 6974 78024
rect 3514 71576 3570 71632
rect 4158 59880 4214 59936
rect 3422 19352 3478 19408
rect 7562 75112 7618 75168
rect 3422 6432 3478 6488
rect 8298 65456 8354 65512
rect 20718 78104 20774 78160
rect 17222 71032 17278 71088
rect 12438 55800 12494 55856
rect 34518 76472 34574 76528
rect 25502 57160 25558 57216
rect 27618 61376 27674 61432
rect 27710 50224 27766 50280
rect 30378 48864 30434 48920
rect 35898 75248 35954 75304
rect 39302 47504 39358 47560
rect 44178 46144 44234 46200
rect 52458 71168 52514 71224
rect 49698 53080 49754 53136
rect 54482 73752 54538 73808
rect 56598 54440 56654 54496
rect 60830 55936 60886 55992
rect 63498 43424 63554 43480
rect 71042 75384 71098 75440
rect 75182 61512 75238 61568
rect 78678 72392 78734 72448
rect 77298 66816 77354 66872
rect 81438 60016 81494 60072
rect 80058 57296 80114 57352
rect 84198 55120 84254 55176
rect 88338 62872 88394 62928
rect 93122 65592 93178 65648
rect 92478 58656 92534 58712
rect 93858 58792 93914 58848
rect 95238 50360 95294 50416
rect 97722 195336 97778 195392
rect 97814 71712 97870 71768
rect 100666 191528 100722 191584
rect 99102 76608 99158 76664
rect 100574 191120 100630 191176
rect 99286 186904 99342 186960
rect 97998 64096 98054 64152
rect 97538 58520 97594 58576
rect 99838 77152 99894 77208
rect 99378 76744 99434 76800
rect 98826 60560 98882 60616
rect 99286 60560 99342 60616
rect 98826 59880 98882 59936
rect 99470 75792 99526 75848
rect 99930 75792 99986 75848
rect 99470 75248 99526 75304
rect 100022 71304 100078 71360
rect 100298 78784 100354 78840
rect 100114 62056 100170 62112
rect 100114 61376 100170 61432
rect 99470 50904 99526 50960
rect 100574 50904 100630 50960
rect 99470 50224 99526 50280
rect 101218 71576 101274 71632
rect 101494 77016 101550 77072
rect 101862 196696 101918 196752
rect 102046 191256 102102 191312
rect 101954 190984 102010 191040
rect 100758 57840 100814 57896
rect 101862 57840 101918 57896
rect 100758 57160 100814 57216
rect 99470 49544 99526 49600
rect 100666 49544 100722 49600
rect 99470 48864 99526 48920
rect 100758 48184 100814 48240
rect 101954 48184 102010 48240
rect 100758 47504 100814 47560
rect 102690 146920 102746 146976
rect 102598 80688 102654 80744
rect 102138 53216 102194 53272
rect 100758 46824 100814 46880
rect 102046 46824 102102 46880
rect 100758 46144 100814 46200
rect 104346 196560 104402 196616
rect 102782 75520 102838 75576
rect 102230 44104 102286 44160
rect 102690 44104 102746 44160
rect 102230 43424 102286 43480
rect 103978 75656 104034 75712
rect 105634 198056 105690 198112
rect 105542 196968 105598 197024
rect 104530 195744 104586 195800
rect 104622 65456 104678 65512
rect 104806 187040 104862 187096
rect 104438 55936 104494 55992
rect 105266 78240 105322 78296
rect 105358 60424 105414 60480
rect 104806 55120 104862 55176
rect 107290 199552 107346 199608
rect 106186 190168 106242 190224
rect 106830 189760 106886 189816
rect 106646 187176 106702 187232
rect 106278 73616 106334 73672
rect 106186 61920 106242 61976
rect 105450 54984 105506 55040
rect 105450 54440 105506 54496
rect 106830 74024 106886 74080
rect 106830 73788 106832 73808
rect 106832 73788 106884 73808
rect 106884 73788 106886 73808
rect 106830 73752 106886 73788
rect 108210 189624 108266 189680
rect 107474 187312 107530 187368
rect 106646 53624 106702 53680
rect 106646 53216 106702 53272
rect 107474 57704 107530 57760
rect 108486 190032 108542 190088
rect 108302 73072 108358 73128
rect 108302 72392 108358 72448
rect 109038 66816 109094 66872
rect 108302 65592 108358 65648
rect 110050 189896 110106 189952
rect 110234 68040 110290 68096
rect 110050 67496 110106 67552
rect 110878 144064 110934 144120
rect 111246 145832 111302 145888
rect 111798 73616 111854 73672
rect 111614 72936 111670 72992
rect 112350 138760 112406 138816
rect 112258 81232 112314 81288
rect 112902 144744 112958 144800
rect 112350 70216 112406 70272
rect 113730 192616 113786 192672
rect 114006 76744 114062 76800
rect 113454 75248 113510 75304
rect 112442 68856 112498 68912
rect 111522 68448 111578 68504
rect 111246 64096 111302 64152
rect 110510 58520 110566 58576
rect 115478 187584 115534 187640
rect 115386 138896 115442 138952
rect 115294 74160 115350 74216
rect 115570 146240 115626 146296
rect 115846 144744 115902 144800
rect 115754 72800 115810 72856
rect 115478 68856 115534 68912
rect 115110 63280 115166 63336
rect 115110 62872 115166 62928
rect 116766 139168 116822 139224
rect 116950 76744 117006 76800
rect 117226 144744 117282 144800
rect 117594 144200 117650 144256
rect 117226 143384 117282 143440
rect 118146 143928 118202 143984
rect 117870 80416 117926 80472
rect 118330 76880 118386 76936
rect 118514 197104 118570 197160
rect 118514 72664 118570 72720
rect 118974 79192 119030 79248
rect 119434 146104 119490 146160
rect 119710 142704 119766 142760
rect 119526 139440 119582 139496
rect 119342 79056 119398 79112
rect 120446 80824 120502 80880
rect 121274 198872 121330 198928
rect 120722 138624 120778 138680
rect 120814 86128 120870 86184
rect 120722 81912 120778 81968
rect 120814 80552 120870 80608
rect 121458 81232 121514 81288
rect 121458 77560 121514 77616
rect 121826 133864 121882 133920
rect 121734 85992 121790 86048
rect 117042 69536 117098 69592
rect 121826 80144 121882 80200
rect 116766 67224 116822 67280
rect 122194 81096 122250 81152
rect 122378 81912 122434 81968
rect 122286 80960 122342 81016
rect 122378 74024 122434 74080
rect 127346 263064 127402 263120
rect 125598 262384 125654 262440
rect 123206 260752 123262 260808
rect 127254 260072 127310 260128
rect 127622 260480 127678 260536
rect 127622 260072 127678 260128
rect 135902 265104 135958 265160
rect 137834 263744 137890 263800
rect 137466 261024 137522 261080
rect 124862 259664 124918 259720
rect 127254 259664 127310 259720
rect 138754 264968 138810 265024
rect 138662 262520 138718 262576
rect 123298 259528 123354 259584
rect 140318 262656 140374 262712
rect 140778 260072 140834 260128
rect 141744 260072 141800 260128
rect 142250 262928 142306 262984
rect 142894 262928 142950 262984
rect 143630 260208 143686 260264
rect 144504 260208 144560 260264
rect 145286 263608 145342 263664
rect 145562 263608 145618 263664
rect 144918 259800 144974 259856
rect 146942 262792 146998 262848
rect 147678 259936 147734 259992
rect 149058 260208 149114 260264
rect 150898 262792 150954 262848
rect 150024 260208 150080 260264
rect 153842 262520 153898 262576
rect 155866 262384 155922 262440
rect 156050 277480 156106 277536
rect 155958 260208 156014 260264
rect 156648 260208 156704 260264
rect 148138 259664 148194 259720
rect 158718 260888 158774 260944
rect 160098 260208 160154 260264
rect 161064 260208 161120 260264
rect 156878 259800 156934 259856
rect 161202 259936 161258 259992
rect 163502 264968 163558 265024
rect 164974 262656 165030 262712
rect 166262 265104 166318 265160
rect 166032 260072 166088 260128
rect 155222 259664 155278 259720
rect 164606 259528 164662 259584
rect 123758 259392 123814 259448
rect 185674 259392 185730 259448
rect 129002 200640 129058 200696
rect 124862 200504 124918 200560
rect 124034 200096 124090 200152
rect 122838 150456 122894 150512
rect 123022 139340 123024 139360
rect 123024 139340 123076 139360
rect 123076 139340 123078 139360
rect 123022 139304 123078 139340
rect 124770 197512 124826 197568
rect 124770 144744 124826 144800
rect 124770 143520 124826 143576
rect 125046 198736 125102 198792
rect 124954 197240 125010 197296
rect 125138 193840 125194 193896
rect 126334 199280 126390 199336
rect 126058 198056 126114 198112
rect 125874 192752 125930 192808
rect 125046 144744 125102 144800
rect 124954 139984 125010 140040
rect 125690 143248 125746 143304
rect 126150 142024 126206 142080
rect 126150 140800 126206 140856
rect 126334 140528 126390 140584
rect 127622 198464 127678 198520
rect 126794 141208 126850 141264
rect 126794 140936 126850 140992
rect 128266 143112 128322 143168
rect 130934 200096 130990 200152
rect 129186 199144 129242 199200
rect 129002 140392 129058 140448
rect 130658 198328 130714 198384
rect 128910 139984 128966 140040
rect 129462 140256 129518 140312
rect 130474 193024 130530 193080
rect 130474 141888 130530 141944
rect 130382 139984 130438 140040
rect 178222 200640 178278 200696
rect 132314 198600 132370 198656
rect 132038 195200 132094 195256
rect 132728 199858 132784 199914
rect 132590 198192 132646 198248
rect 132682 195608 132738 195664
rect 133832 199824 133888 199880
rect 134108 199858 134164 199914
rect 133648 199776 133704 199778
rect 133050 195200 133106 195256
rect 133648 199724 133650 199776
rect 133650 199724 133702 199776
rect 133702 199724 133704 199776
rect 133648 199722 133704 199724
rect 134384 199858 134440 199914
rect 134568 199858 134624 199914
rect 134062 199688 134118 199744
rect 134522 199688 134578 199744
rect 134430 197376 134486 197432
rect 134844 199858 134900 199914
rect 135488 199824 135544 199880
rect 134062 196696 134118 196752
rect 133602 192888 133658 192944
rect 134338 195880 134394 195936
rect 135350 199688 135406 199744
rect 135672 199824 135728 199880
rect 135856 199858 135912 199914
rect 136224 199858 136280 199914
rect 136408 199858 136464 199914
rect 135718 199688 135774 199744
rect 135718 199008 135774 199064
rect 135166 197648 135222 197704
rect 134798 192888 134854 192944
rect 136868 199858 136924 199914
rect 136178 199688 136234 199744
rect 136362 199688 136418 199744
rect 136822 198328 136878 198384
rect 136546 196968 136602 197024
rect 137420 199858 137476 199914
rect 137144 199688 137200 199744
rect 137742 199688 137798 199744
rect 138616 199824 138672 199880
rect 137006 199008 137062 199064
rect 137098 198056 137154 198112
rect 135810 148552 135866 148608
rect 137466 199552 137522 199608
rect 137282 196696 137338 196752
rect 137834 199572 137890 199608
rect 137834 199552 137836 199572
rect 137836 199552 137888 199572
rect 137888 199552 137890 199572
rect 138018 195744 138074 195800
rect 138110 195200 138166 195256
rect 138754 199724 138756 199744
rect 138756 199724 138808 199744
rect 138808 199724 138810 199744
rect 138754 199688 138810 199724
rect 139628 199858 139684 199914
rect 138294 198056 138350 198112
rect 138478 196832 138534 196888
rect 137282 187448 137338 187504
rect 137006 147328 137062 147384
rect 138294 147192 138350 147248
rect 138846 195064 138902 195120
rect 139674 199724 139676 199744
rect 139676 199724 139728 199744
rect 139728 199724 139730 199744
rect 139674 199688 139730 199724
rect 140272 199858 140328 199914
rect 139674 199144 139730 199200
rect 139858 196696 139914 196752
rect 139674 151000 139730 151056
rect 135902 144608 135958 144664
rect 138662 144472 138718 144528
rect 137558 144336 137614 144392
rect 138110 143928 138166 143984
rect 139398 141752 139454 141808
rect 140640 199858 140696 199914
rect 140916 199858 140972 199914
rect 141100 199858 141156 199914
rect 141376 199858 141432 199914
rect 141560 199858 141616 199914
rect 141836 199858 141892 199914
rect 142112 199858 142168 199914
rect 142296 199858 142352 199914
rect 142480 199858 142536 199914
rect 142848 199858 142904 199914
rect 143032 199858 143088 199914
rect 140962 199688 141018 199744
rect 140778 199552 140834 199608
rect 140870 197512 140926 197568
rect 141330 199688 141386 199744
rect 141238 199552 141294 199608
rect 141146 199144 141202 199200
rect 141606 199688 141662 199744
rect 141882 199688 141938 199744
rect 142066 199688 142122 199744
rect 141606 199588 141608 199608
rect 141608 199588 141660 199608
rect 141660 199588 141662 199608
rect 141606 199552 141662 199588
rect 141514 199144 141570 199200
rect 141698 199144 141754 199200
rect 141514 196696 141570 196752
rect 141882 198600 141938 198656
rect 142158 199144 142214 199200
rect 142480 199724 142482 199744
rect 142482 199724 142534 199744
rect 142534 199724 142536 199744
rect 142480 199688 142536 199724
rect 142894 199688 142950 199744
rect 142526 198464 142582 198520
rect 142802 198464 142858 198520
rect 143400 199688 143456 199744
rect 143860 199858 143916 199914
rect 142986 199144 143042 199200
rect 143354 199572 143410 199608
rect 143354 199552 143356 199572
rect 143356 199552 143408 199572
rect 143408 199552 143410 199572
rect 143354 198464 143410 198520
rect 143906 198484 143962 198520
rect 143906 198464 143908 198484
rect 143908 198464 143960 198484
rect 143960 198464 143962 198484
rect 144872 199858 144928 199914
rect 144826 199688 144882 199744
rect 145976 199858 146032 199914
rect 146252 199858 146308 199914
rect 144642 197376 144698 197432
rect 139950 140120 140006 140176
rect 145930 199552 145986 199608
rect 146206 197920 146262 197976
rect 146390 199552 146446 199608
rect 146666 198600 146722 198656
rect 147448 199858 147504 199914
rect 147632 199858 147688 199914
rect 148000 199858 148056 199914
rect 145010 142976 145066 143032
rect 146390 142704 146446 142760
rect 146942 146104 146998 146160
rect 147862 199552 147918 199608
rect 148276 199824 148332 199880
rect 148552 199858 148608 199914
rect 148322 199688 148378 199744
rect 148046 198328 148102 198384
rect 148230 198600 148286 198656
rect 147770 145832 147826 145888
rect 148046 142840 148102 142896
rect 148598 199552 148654 199608
rect 148874 196968 148930 197024
rect 149610 198056 149666 198112
rect 149518 197512 149574 197568
rect 150576 199824 150632 199880
rect 150346 198192 150402 198248
rect 150254 198056 150310 198112
rect 150162 197240 150218 197296
rect 150438 195608 150494 195664
rect 150438 195336 150494 195392
rect 151128 199858 151184 199914
rect 150714 199552 150770 199608
rect 151174 199688 151230 199744
rect 151174 195608 151230 195664
rect 151680 199858 151736 199914
rect 151864 199858 151920 199914
rect 152048 199824 152104 199880
rect 151358 193840 151414 193896
rect 151542 199416 151598 199472
rect 151726 199688 151782 199744
rect 151818 191392 151874 191448
rect 152278 198056 152334 198112
rect 152968 199824 153024 199880
rect 153014 199416 153070 199472
rect 153198 199552 153254 199608
rect 152830 198872 152886 198928
rect 152922 195472 152978 195528
rect 152002 145696 152058 145752
rect 152554 144200 152610 144256
rect 153750 199280 153806 199336
rect 154210 198056 154266 198112
rect 153474 148280 153530 148336
rect 153382 145968 153438 146024
rect 153106 144064 153162 144120
rect 153014 141616 153070 141672
rect 154808 199824 154864 199880
rect 155268 199824 155324 199880
rect 155544 199824 155600 199880
rect 155314 199688 155370 199744
rect 155498 199688 155554 199744
rect 154486 144336 154542 144392
rect 155958 199552 156014 199608
rect 155958 199144 156014 199200
rect 155866 198736 155922 198792
rect 156234 199552 156290 199608
rect 156142 199280 156198 199336
rect 156142 197784 156198 197840
rect 156418 198056 156474 198112
rect 157200 199858 157256 199914
rect 157384 199858 157440 199914
rect 157568 199858 157624 199914
rect 156786 199300 156842 199336
rect 156786 199280 156788 199300
rect 156788 199280 156840 199300
rect 156840 199280 156842 199300
rect 157154 199688 157210 199744
rect 156970 192480 157026 192536
rect 157338 198192 157394 198248
rect 157246 198056 157302 198112
rect 158120 199858 158176 199914
rect 158488 199858 158544 199914
rect 157614 198328 157670 198384
rect 158074 199688 158130 199744
rect 158626 199724 158628 199744
rect 158628 199724 158680 199744
rect 158680 199724 158682 199744
rect 158626 199688 158682 199724
rect 159316 199858 159372 199914
rect 158258 199552 158314 199608
rect 158442 199552 158498 199608
rect 158258 199008 158314 199064
rect 158626 198736 158682 198792
rect 158902 199688 158958 199744
rect 159684 199858 159740 199914
rect 158902 199552 158958 199608
rect 156878 145560 156934 145616
rect 157338 145560 157394 145616
rect 156418 144472 156474 144528
rect 155590 141480 155646 141536
rect 156970 142840 157026 142896
rect 157154 141616 157210 141672
rect 157430 142024 157486 142080
rect 158902 195200 158958 195256
rect 158902 193976 158958 194032
rect 159914 199552 159970 199608
rect 160604 199858 160660 199914
rect 160098 199144 160154 199200
rect 160558 199688 160614 199744
rect 160558 199552 160614 199608
rect 161432 199858 161488 199914
rect 160650 190032 160706 190088
rect 161110 195336 161166 195392
rect 162168 199858 162224 199914
rect 162444 199858 162500 199914
rect 163548 199858 163604 199914
rect 163732 199824 163788 199880
rect 164008 199858 164064 199914
rect 162306 198192 162362 198248
rect 162214 196968 162270 197024
rect 162214 196832 162270 196888
rect 162398 197784 162454 197840
rect 162306 190984 162362 191040
rect 162490 196832 162546 196888
rect 163134 199724 163136 199744
rect 163136 199724 163188 199744
rect 163188 199724 163190 199744
rect 163134 199688 163190 199724
rect 161754 142976 161810 143032
rect 161202 140120 161258 140176
rect 163134 199552 163190 199608
rect 163502 199688 163558 199744
rect 163686 199688 163742 199744
rect 164192 199824 164248 199880
rect 164560 199824 164616 199880
rect 163962 199552 164018 199608
rect 164514 199688 164570 199744
rect 164238 196560 164294 196616
rect 165112 199824 165168 199880
rect 165066 199416 165122 199472
rect 164974 197784 165030 197840
rect 165342 199688 165398 199744
rect 165756 199858 165812 199914
rect 165250 197240 165306 197296
rect 166078 199688 166134 199744
rect 166400 199858 166456 199914
rect 166768 199858 166824 199914
rect 165802 198464 165858 198520
rect 164238 147056 164294 147112
rect 164238 145696 164294 145752
rect 167044 199722 167100 199778
rect 167504 199824 167560 199880
rect 168240 199858 168296 199914
rect 166722 198056 166778 198112
rect 166630 196696 166686 196752
rect 165710 146920 165766 146976
rect 165526 144744 165582 144800
rect 166998 197376 167054 197432
rect 167458 199688 167514 199744
rect 167918 199552 167974 199608
rect 168194 199688 168250 199744
rect 168102 193296 168158 193352
rect 168976 199824 169032 199880
rect 168930 199688 168986 199744
rect 169436 199858 169492 199914
rect 169620 199858 169676 199914
rect 168746 195880 168802 195936
rect 168838 194248 168894 194304
rect 169298 199008 169354 199064
rect 169298 197784 169354 197840
rect 169390 196288 169446 196344
rect 168746 156576 168802 156632
rect 168470 149912 168526 149968
rect 167090 149776 167146 149832
rect 167458 141752 167514 141808
rect 169574 199688 169630 199744
rect 170080 199858 170136 199914
rect 169666 197920 169722 197976
rect 169666 196424 169722 196480
rect 170126 199688 170182 199744
rect 170632 199858 170688 199914
rect 171276 199858 171332 199914
rect 171828 199858 171884 199914
rect 172104 199824 172160 199880
rect 172380 199858 172436 199914
rect 170218 198872 170274 198928
rect 170494 198192 170550 198248
rect 170402 193160 170458 193216
rect 170586 196424 170642 196480
rect 169850 147464 169906 147520
rect 170770 198464 170826 198520
rect 170954 198600 171010 198656
rect 171138 198328 171194 198384
rect 170954 198192 171010 198248
rect 171322 199552 171378 199608
rect 170862 147328 170918 147384
rect 169942 140392 169998 140448
rect 169758 140256 169814 140312
rect 171874 199552 171930 199608
rect 171782 192616 171838 192672
rect 172564 199858 172620 199914
rect 172748 199858 172804 199914
rect 172426 199552 172482 199608
rect 172794 199688 172850 199744
rect 172518 198736 172574 198792
rect 172426 197784 172482 197840
rect 172518 197376 172574 197432
rect 173116 199858 173172 199914
rect 173300 199824 173356 199880
rect 172518 148960 172574 149016
rect 172702 148416 172758 148472
rect 171138 140528 171194 140584
rect 173760 199824 173816 199880
rect 174128 199858 174184 199914
rect 173530 199008 173586 199064
rect 173622 198736 173678 198792
rect 173622 197784 173678 197840
rect 173438 194112 173494 194168
rect 173806 199572 173862 199608
rect 173806 199552 173808 199572
rect 173808 199552 173860 199572
rect 173860 199552 173862 199572
rect 174312 199858 174368 199914
rect 173806 195608 173862 195664
rect 172886 148144 172942 148200
rect 174772 199824 174828 199880
rect 174956 199824 175012 199880
rect 175140 199858 175196 199914
rect 174726 199688 174782 199744
rect 174358 199552 174414 199608
rect 174358 199416 174414 199472
rect 174358 198872 174414 198928
rect 174634 199416 174690 199472
rect 174542 198872 174598 198928
rect 174910 198872 174966 198928
rect 175278 198328 175334 198384
rect 175186 195608 175242 195664
rect 175692 199858 175748 199914
rect 176428 199824 176484 199880
rect 175646 198736 175702 198792
rect 175830 199008 175886 199064
rect 175922 198736 175978 198792
rect 175462 151272 175518 151328
rect 175370 148824 175426 148880
rect 175278 145832 175334 145888
rect 176382 198872 176438 198928
rect 176566 195880 176622 195936
rect 176658 193976 176714 194032
rect 176658 151136 176714 151192
rect 177486 199824 177542 199880
rect 177210 198736 177266 198792
rect 177394 199280 177450 199336
rect 177394 198736 177450 198792
rect 177946 200096 178002 200152
rect 177762 195064 177818 195120
rect 177946 198600 178002 198656
rect 178590 199144 178646 199200
rect 178222 198600 178278 198656
rect 177026 153856 177082 153912
rect 176842 153720 176898 153776
rect 177854 141344 177910 141400
rect 177946 139984 178002 140040
rect 179418 192344 179474 192400
rect 178958 142704 179014 142760
rect 180246 195744 180302 195800
rect 181442 200368 181498 200424
rect 180338 146104 180394 146160
rect 180522 145968 180578 146024
rect 180154 139984 180210 140040
rect 181442 147600 181498 147656
rect 181902 141344 181958 141400
rect 183650 151000 183706 151056
rect 183098 143384 183154 143440
rect 183742 143112 183798 143168
rect 183742 142296 183798 142352
rect 183006 140664 183062 140720
rect 183374 140120 183430 140176
rect 184294 143248 184350 143304
rect 184294 142160 184350 142216
rect 183374 139848 183430 139904
rect 181810 139712 181866 139768
rect 185398 140120 185454 140176
rect 185582 140528 185638 140584
rect 185582 140120 185638 140176
rect 185582 139576 185638 139632
rect 184386 139440 184442 139496
rect 123942 139304 123998 139360
rect 125506 139304 125562 139360
rect 130566 139304 130622 139360
rect 130842 139304 130898 139360
rect 162306 139304 162362 139360
rect 169482 139304 169538 139360
rect 173622 139304 173678 139360
rect 186226 139440 186282 139496
rect 186226 139304 186282 139360
rect 122746 80552 122802 80608
rect 123942 80416 123998 80472
rect 122654 78376 122710 78432
rect 123482 78240 123538 78296
rect 131946 80552 132002 80608
rect 131670 80144 131726 80200
rect 128634 80008 128690 80064
rect 126058 79872 126114 79928
rect 124862 78104 124918 78160
rect 126242 79328 126298 79384
rect 126058 77424 126114 77480
rect 129002 78376 129058 78432
rect 128174 71168 128230 71224
rect 129738 75248 129794 75304
rect 130842 77560 130898 77616
rect 132544 79872 132600 79928
rect 132038 78512 132094 78568
rect 131670 78376 131726 78432
rect 132314 78376 132370 78432
rect 131578 76608 131634 76664
rect 132728 79736 132784 79792
rect 132590 76608 132646 76664
rect 133096 79872 133152 79928
rect 133464 79906 133520 79962
rect 133510 79736 133566 79792
rect 133510 77152 133566 77208
rect 133326 74568 133382 74624
rect 133694 79600 133750 79656
rect 134476 79872 134532 79928
rect 134752 79906 134808 79962
rect 133878 77288 133934 77344
rect 134154 78784 134210 78840
rect 134062 76608 134118 76664
rect 133970 75520 134026 75576
rect 134062 71304 134118 71360
rect 134522 77968 134578 78024
rect 134522 77832 134578 77888
rect 135120 79872 135176 79928
rect 135304 79872 135360 79928
rect 135764 79872 135820 79928
rect 134982 77016 135038 77072
rect 135258 74704 135314 74760
rect 135534 79464 135590 79520
rect 135902 77016 135958 77072
rect 135626 75248 135682 75304
rect 135718 71576 135774 71632
rect 136224 79736 136280 79792
rect 136776 79872 136832 79928
rect 136178 79348 136234 79384
rect 136178 79328 136180 79348
rect 136180 79328 136232 79348
rect 136232 79328 136234 79348
rect 136730 79636 136732 79656
rect 136732 79636 136784 79656
rect 136784 79636 136786 79656
rect 136730 79600 136786 79636
rect 136730 73888 136786 73944
rect 137144 79736 137200 79792
rect 137696 79872 137752 79928
rect 137558 79600 137614 79656
rect 138064 79872 138120 79928
rect 138708 79906 138764 79962
rect 138892 79872 138948 79928
rect 138616 79736 138672 79792
rect 138294 68312 138350 68368
rect 139720 79906 139776 79962
rect 139536 79736 139592 79792
rect 140088 79872 140144 79928
rect 139582 76608 139638 76664
rect 140272 79736 140328 79792
rect 141100 79906 141156 79962
rect 140318 79600 140374 79656
rect 140870 79736 140926 79792
rect 140870 79636 140872 79656
rect 140872 79636 140924 79656
rect 140924 79636 140926 79656
rect 140870 79600 140926 79636
rect 141560 79872 141616 79928
rect 141514 79736 141570 79792
rect 141238 77424 141294 77480
rect 142112 79872 142168 79928
rect 142296 79906 142352 79962
rect 142388 79824 142444 79826
rect 142388 79772 142390 79824
rect 142390 79772 142442 79824
rect 142442 79772 142444 79824
rect 142388 79770 142444 79772
rect 141882 79600 141938 79656
rect 141698 76744 141754 76800
rect 142066 77832 142122 77888
rect 142618 79600 142674 79656
rect 142342 78104 142398 78160
rect 142618 78648 142674 78704
rect 143124 79872 143180 79928
rect 143308 79906 143364 79962
rect 143584 79736 143640 79792
rect 143262 79600 143318 79656
rect 144596 79872 144652 79928
rect 144550 79736 144606 79792
rect 144182 77560 144238 77616
rect 144458 77832 144514 77888
rect 144458 77696 144514 77752
rect 145056 79872 145112 79928
rect 145240 79906 145296 79962
rect 144642 74704 144698 74760
rect 144826 76608 144882 76664
rect 145424 79872 145480 79928
rect 145470 79736 145526 79792
rect 145884 79872 145940 79928
rect 146344 79838 146400 79894
rect 146160 79736 146216 79792
rect 146712 79906 146768 79962
rect 145930 79600 145986 79656
rect 145838 76880 145894 76936
rect 145838 76608 145894 76664
rect 146298 79600 146354 79656
rect 146666 79736 146722 79792
rect 147080 79872 147136 79928
rect 147264 79906 147320 79962
rect 147448 79906 147504 79962
rect 147632 79872 147688 79928
rect 148552 79906 148608 79962
rect 146850 79464 146906 79520
rect 147034 78648 147090 78704
rect 146942 76608 146998 76664
rect 148644 79736 148700 79792
rect 149380 79906 149436 79962
rect 149564 79872 149620 79928
rect 150300 79906 150356 79962
rect 148414 77424 148470 77480
rect 148598 77288 148654 77344
rect 148874 79328 148930 79384
rect 148966 77152 149022 77208
rect 149610 79328 149666 79384
rect 149518 78512 149574 78568
rect 149610 74024 149666 74080
rect 151220 79872 151276 79928
rect 149886 71440 149942 71496
rect 150254 77288 150310 77344
rect 150346 74024 150402 74080
rect 150530 79192 150586 79248
rect 151680 79872 151736 79928
rect 150990 79600 151046 79656
rect 150898 79056 150954 79112
rect 150806 77288 150862 77344
rect 150806 73072 150862 73128
rect 151082 79192 151138 79248
rect 152048 79838 152104 79894
rect 151726 78648 151782 78704
rect 151634 76472 151690 76528
rect 151542 73072 151598 73128
rect 151910 74432 151966 74488
rect 152784 79872 152840 79928
rect 152738 79600 152794 79656
rect 152738 79464 152794 79520
rect 152554 79192 152610 79248
rect 152094 69808 152150 69864
rect 153014 74432 153070 74488
rect 152830 66000 152886 66056
rect 152646 65864 152702 65920
rect 153612 79906 153668 79962
rect 153796 79906 153852 79962
rect 153980 79906 154036 79962
rect 154164 79872 154220 79928
rect 153290 79600 153346 79656
rect 153566 79464 153622 79520
rect 153658 78784 153714 78840
rect 153934 79736 153990 79792
rect 154210 79736 154266 79792
rect 153842 77424 153898 77480
rect 154900 79906 154956 79962
rect 154854 79464 154910 79520
rect 154854 78920 154910 78976
rect 155268 79906 155324 79962
rect 154486 77288 154542 77344
rect 154670 76880 154726 76936
rect 154118 70080 154174 70136
rect 154026 69944 154082 70000
rect 153658 69672 153714 69728
rect 154946 67496 155002 67552
rect 155636 79872 155692 79928
rect 156096 79838 156152 79894
rect 155866 77288 155922 77344
rect 155498 74296 155554 74352
rect 155222 68720 155278 68776
rect 155774 67496 155830 67552
rect 156050 79600 156106 79656
rect 156464 79906 156520 79962
rect 157292 79872 157348 79928
rect 157568 79906 157624 79962
rect 158028 79906 158084 79962
rect 156602 79600 156658 79656
rect 156510 78512 156566 78568
rect 156602 67632 156658 67688
rect 155958 37848 156014 37904
rect 156878 68584 156934 68640
rect 156878 67632 156934 67688
rect 156694 66136 156750 66192
rect 158304 79906 158360 79962
rect 158580 79906 158636 79962
rect 158074 78104 158130 78160
rect 158626 79600 158682 79656
rect 157982 28192 158038 28248
rect 157798 10240 157854 10296
rect 158810 78920 158866 78976
rect 159132 79872 159188 79928
rect 159408 79736 159464 79792
rect 159178 78648 159234 78704
rect 160052 79824 160108 79826
rect 159546 78512 159602 78568
rect 160052 79772 160054 79824
rect 160054 79772 160106 79824
rect 160106 79772 160108 79824
rect 160052 79770 160108 79772
rect 160880 79872 160936 79928
rect 160650 78648 160706 78704
rect 160926 78648 160982 78704
rect 161432 79872 161488 79928
rect 161984 79872 162040 79928
rect 162352 79906 162408 79962
rect 162628 79906 162684 79962
rect 160374 67224 160430 67280
rect 160558 67088 160614 67144
rect 160190 51720 160246 51776
rect 161018 67088 161074 67144
rect 161478 78240 161534 78296
rect 161202 67224 161258 67280
rect 162536 79736 162592 79792
rect 162490 77288 162546 77344
rect 163272 79872 163328 79928
rect 163456 79906 163512 79962
rect 163410 79772 163412 79792
rect 163412 79772 163464 79792
rect 163464 79772 163466 79792
rect 163410 79736 163466 79772
rect 163640 79736 163696 79792
rect 161846 68720 161902 68776
rect 161662 68584 161718 68640
rect 162766 68584 162822 68640
rect 163226 77968 163282 78024
rect 163318 77832 163374 77888
rect 163502 77288 163558 77344
rect 163686 77288 163742 77344
rect 163226 69808 163282 69864
rect 163870 77696 163926 77752
rect 164560 79872 164616 79928
rect 165020 79872 165076 79928
rect 164146 77832 164202 77888
rect 164330 79600 164386 79656
rect 164330 78920 164386 78976
rect 164146 69808 164202 69864
rect 164790 79600 164846 79656
rect 165296 79736 165352 79792
rect 165480 79736 165536 79792
rect 165848 79872 165904 79928
rect 165158 72528 165214 72584
rect 165710 79328 165766 79384
rect 166400 79906 166456 79962
rect 167044 79838 167100 79894
rect 166676 79772 166678 79792
rect 166678 79772 166730 79792
rect 166730 79772 166732 79792
rect 166078 79600 166134 79656
rect 165986 79348 166042 79384
rect 165986 79328 165988 79348
rect 165988 79328 166040 79348
rect 166040 79328 166042 79348
rect 166676 79736 166732 79772
rect 167228 79906 167284 79962
rect 167504 79736 167560 79792
rect 168056 79906 168112 79962
rect 168240 79872 168296 79928
rect 168608 79906 168664 79962
rect 168884 79906 168940 79962
rect 169344 79872 169400 79928
rect 166998 79600 167054 79656
rect 166906 79192 166962 79248
rect 167090 79348 167146 79384
rect 167090 79328 167092 79348
rect 167092 79328 167144 79348
rect 167144 79328 167146 79348
rect 168286 79736 168342 79792
rect 167182 77288 167238 77344
rect 167458 79328 167514 79384
rect 167918 79600 167974 79656
rect 168102 79600 168158 79656
rect 167642 75520 167698 75576
rect 167550 75384 167606 75440
rect 167734 71576 167790 71632
rect 167918 71712 167974 71768
rect 168378 79600 168434 79656
rect 168286 75112 168342 75168
rect 168286 71712 168342 71768
rect 168194 71576 168250 71632
rect 168654 79328 168710 79384
rect 169390 79056 169446 79112
rect 169988 79906 170044 79962
rect 170264 79872 170320 79928
rect 170034 79772 170036 79792
rect 170036 79772 170088 79792
rect 170088 79772 170090 79792
rect 170034 79736 170090 79772
rect 170540 79906 170596 79962
rect 170816 79906 170872 79962
rect 170034 79600 170090 79656
rect 169758 79328 169814 79384
rect 169574 75248 169630 75304
rect 169206 71032 169262 71088
rect 170034 78512 170090 78568
rect 170310 79600 170366 79656
rect 170218 74432 170274 74488
rect 170954 79636 170956 79656
rect 170956 79636 171008 79656
rect 171008 79636 171010 79656
rect 170954 79600 171010 79636
rect 170494 78648 170550 78704
rect 170678 76744 170734 76800
rect 170494 75928 170550 75984
rect 170678 75928 170734 75984
rect 170586 74432 170642 74488
rect 170586 73616 170642 73672
rect 170402 35128 170458 35184
rect 171644 79906 171700 79962
rect 171138 79328 171194 79384
rect 170954 71304 171010 71360
rect 171414 77968 171470 78024
rect 171920 79906 171976 79962
rect 172288 79906 172344 79962
rect 172748 79906 172804 79962
rect 172150 78648 172206 78704
rect 171598 72936 171654 72992
rect 171230 71712 171286 71768
rect 171230 71440 171286 71496
rect 172656 79736 172712 79792
rect 172794 79736 172850 79792
rect 172426 79600 172482 79656
rect 172702 79600 172758 79656
rect 172334 72936 172390 72992
rect 172426 72392 172482 72448
rect 173024 79736 173080 79792
rect 173208 79872 173264 79928
rect 173484 79872 173540 79928
rect 173254 79736 173310 79792
rect 173070 79600 173126 79656
rect 173254 79600 173310 79656
rect 173760 79906 173816 79962
rect 173346 79328 173402 79384
rect 173530 79600 173586 79656
rect 174496 79908 174498 79928
rect 174498 79908 174550 79928
rect 174550 79908 174552 79928
rect 174496 79872 174552 79908
rect 174680 79906 174736 79962
rect 174956 79906 175012 79962
rect 175324 79872 175380 79928
rect 175784 79906 175840 79962
rect 176060 79906 176116 79962
rect 173990 79600 174046 79656
rect 173346 71440 173402 71496
rect 173714 78240 173770 78296
rect 173714 78104 173770 78160
rect 173714 76880 173770 76936
rect 173530 76608 173586 76664
rect 173622 76336 173678 76392
rect 172978 69536 173034 69592
rect 173622 69536 173678 69592
rect 174542 79756 174598 79792
rect 174542 79736 174544 79756
rect 174544 79736 174596 79756
rect 174596 79736 174598 79756
rect 174634 79600 174690 79656
rect 176244 79906 176300 79962
rect 175186 79600 175242 79656
rect 175278 78376 175334 78432
rect 175186 71168 175242 71224
rect 175738 79636 175740 79656
rect 175740 79636 175792 79656
rect 175792 79636 175794 79656
rect 175738 79600 175794 79636
rect 175738 77424 175794 77480
rect 175646 77288 175702 77344
rect 175922 78648 175978 78704
rect 176106 77560 176162 77616
rect 175922 76916 175924 76936
rect 175924 76916 175976 76936
rect 175976 76916 175978 76936
rect 175922 76880 175978 76916
rect 175830 72800 175886 72856
rect 175738 69808 175794 69864
rect 176980 79872 177036 79928
rect 176382 78240 176438 78296
rect 176382 77424 176438 77480
rect 176658 79328 176714 79384
rect 177026 79736 177082 79792
rect 176474 77016 176530 77072
rect 176198 72664 176254 72720
rect 176566 72800 176622 72856
rect 176566 72664 176622 72720
rect 177532 79906 177588 79962
rect 177486 78240 177542 78296
rect 177486 74976 177542 75032
rect 177026 68448 177082 68504
rect 180522 80552 180578 80608
rect 185766 80416 185822 80472
rect 184202 80144 184258 80200
rect 180522 79872 180578 79928
rect 179510 79600 179566 79656
rect 177854 76880 177910 76936
rect 178038 68176 178094 68232
rect 178774 77968 178830 78024
rect 178958 75248 179014 75304
rect 179050 75112 179106 75168
rect 179510 77968 179566 78024
rect 180522 78376 180578 78432
rect 181626 77832 181682 77888
rect 182086 77832 182142 77888
rect 181626 72800 181682 72856
rect 181442 72528 181498 72584
rect 181626 72528 181682 72584
rect 181442 72256 181498 72312
rect 181810 71032 181866 71088
rect 185398 70352 185454 70408
rect 187146 144200 187202 144256
rect 187054 139304 187110 139360
rect 187422 213832 187478 213888
rect 188066 262520 188122 262576
rect 187514 144064 187570 144120
rect 187698 144336 187754 144392
rect 187698 139576 187754 139632
rect 187606 138080 187662 138136
rect 187330 79872 187386 79928
rect 187238 63416 187294 63472
rect 187698 57160 187754 57216
rect 186594 56208 186650 56264
rect 188526 262928 188582 262984
rect 188526 262520 188582 262576
rect 188894 259936 188950 259992
rect 188250 139168 188306 139224
rect 188434 117952 188490 118008
rect 188526 81368 188582 81424
rect 188342 64096 188398 64152
rect 187790 38528 187846 38584
rect 187790 37848 187846 37904
rect 188894 142976 188950 143032
rect 189078 140564 189080 140584
rect 189080 140564 189132 140584
rect 189132 140564 189134 140584
rect 189078 140528 189134 140564
rect 189078 81504 189134 81560
rect 189722 260072 189778 260128
rect 189538 81776 189594 81832
rect 189538 79600 189594 79656
rect 189814 81912 189870 81968
rect 189722 80280 189778 80336
rect 190458 195472 190514 195528
rect 190826 78240 190882 78296
rect 191194 136584 191250 136640
rect 191286 82048 191342 82104
rect 192666 262792 192722 262848
rect 192482 262248 192538 262304
rect 192666 193840 192722 193896
rect 192666 147192 192722 147248
rect 192574 139304 192630 139360
rect 193126 76472 193182 76528
rect 190734 52128 190790 52184
rect 191838 46144 191894 46200
rect 190458 43968 190514 44024
rect 191746 43968 191802 44024
rect 191746 43696 191802 43752
rect 193218 57840 193274 57896
rect 193770 149640 193826 149696
rect 193494 140700 193496 140720
rect 193496 140700 193548 140720
rect 193548 140700 193550 140720
rect 193494 140664 193550 140700
rect 193402 67496 193458 67552
rect 193954 139032 194010 139088
rect 193310 52264 193366 52320
rect 193310 50224 193366 50280
rect 194046 135904 194102 135960
rect 194322 144608 194378 144664
rect 194782 195336 194838 195392
rect 194690 192888 194746 192944
rect 194598 53624 194654 53680
rect 194506 52264 194562 52320
rect 194506 51992 194562 52048
rect 196070 196968 196126 197024
rect 195978 196832 196034 196888
rect 195426 137808 195482 137864
rect 195426 82184 195482 82240
rect 194874 64504 194930 64560
rect 194874 64232 194930 64288
rect 194782 54848 194838 54904
rect 194690 50360 194746 50416
rect 197358 197104 197414 197160
rect 196622 138896 196678 138952
rect 196162 66136 196218 66192
rect 196714 81776 196770 81832
rect 196898 81504 196954 81560
rect 196254 59064 196310 59120
rect 196070 56344 196126 56400
rect 196070 56072 196126 56128
rect 195978 49408 196034 49464
rect 196438 49408 196494 49464
rect 196438 49136 196494 49192
rect 197542 196560 197598 196616
rect 197358 44104 197414 44160
rect 197358 43560 197414 43616
rect 198370 200504 198426 200560
rect 198186 149096 198242 149152
rect 198002 57568 198058 57624
rect 197634 52400 197690 52456
rect 198278 52400 198334 52456
rect 198278 51856 198334 51912
rect 197542 48048 197598 48104
rect 197542 47776 197598 47832
rect 200394 200232 200450 200288
rect 200210 196696 200266 196752
rect 199014 143248 199070 143304
rect 199382 138760 199438 138816
rect 199658 147600 199714 147656
rect 199198 66408 199254 66464
rect 198922 64776 198978 64832
rect 198830 57704 198886 57760
rect 201866 259528 201922 259584
rect 200486 69672 200542 69728
rect 201038 149096 201094 149152
rect 201038 80008 201094 80064
rect 200854 71576 200910 71632
rect 200394 54984 200450 55040
rect 200302 53760 200358 53816
rect 200210 45328 200266 45384
rect 201406 54984 201462 55040
rect 201406 54712 201462 54768
rect 201406 53760 201462 53816
rect 201406 53216 201462 53272
rect 201682 67496 201738 67552
rect 201774 63280 201830 63336
rect 202418 156848 202474 156904
rect 202234 80960 202290 81016
rect 202142 62056 202198 62112
rect 202510 139440 202566 139496
rect 202786 63280 202842 63336
rect 202786 62736 202842 62792
rect 202418 61512 202474 61568
rect 201866 58656 201922 58712
rect 201590 55936 201646 55992
rect 203614 148280 203670 148336
rect 203522 72936 203578 72992
rect 204166 66816 204222 66872
rect 234618 278024 234674 278080
rect 282918 263064 282974 263120
rect 347778 262928 347834 262984
rect 580170 697176 580226 697232
rect 580170 683848 580226 683904
rect 580170 670692 580172 670712
rect 580172 670692 580224 670712
rect 580224 670692 580226 670712
rect 580170 670656 580226 670692
rect 580170 644000 580226 644056
rect 580170 630808 580226 630864
rect 580170 617480 580226 617536
rect 579802 590960 579858 591016
rect 580170 577632 580226 577688
rect 579802 564304 579858 564360
rect 580170 537784 580226 537840
rect 580170 524476 580226 524512
rect 580170 524456 580172 524476
rect 580172 524456 580224 524476
rect 580224 524456 580226 524476
rect 580170 511264 580226 511320
rect 580170 484608 580226 484664
rect 579986 471416 580042 471472
rect 580170 458088 580226 458144
rect 580170 431568 580226 431624
rect 580170 418240 580226 418296
rect 580170 404912 580226 404968
rect 580170 378392 580226 378448
rect 580262 365064 580318 365120
rect 580170 351908 580172 351928
rect 580172 351908 580224 351928
rect 580224 351908 580226 351928
rect 580170 351872 580226 351908
rect 580170 325216 580226 325272
rect 579986 312024 580042 312080
rect 580170 298696 580226 298752
rect 580170 272176 580226 272232
rect 477498 262792 477554 262848
rect 203246 57704 203302 57760
rect 203062 48220 203064 48240
rect 203064 48220 203116 48240
rect 203116 48220 203118 48240
rect 203062 48184 203118 48220
rect 205178 192752 205234 192808
rect 204810 192480 204866 192536
rect 204902 148688 204958 148744
rect 204810 75248 204866 75304
rect 205086 72800 205142 72856
rect 205822 192616 205878 192672
rect 580170 258848 580226 258904
rect 580170 245556 580172 245576
rect 580172 245556 580224 245576
rect 580224 245556 580226 245576
rect 580170 245520 580226 245556
rect 580446 232328 580502 232384
rect 580354 219000 580410 219056
rect 579802 205672 579858 205728
rect 207018 194112 207074 194168
rect 206098 143112 206154 143168
rect 206098 141480 206154 141536
rect 204994 49272 205050 49328
rect 204994 49000 205050 49056
rect 204534 44920 204590 44976
rect 206466 80824 206522 80880
rect 206374 77968 206430 78024
rect 206374 75812 206430 75848
rect 206374 75792 206376 75812
rect 206376 75792 206428 75812
rect 206428 75792 206430 75812
rect 207202 69400 207258 69456
rect 208398 189760 208454 189816
rect 207110 46552 207166 46608
rect 207018 45192 207074 45248
rect 207018 44784 207074 44840
rect 207018 44124 207074 44160
rect 207018 44104 207020 44124
rect 207020 44104 207072 44124
rect 207072 44104 207074 44124
rect 206098 35808 206154 35864
rect 206098 35128 206154 35184
rect 207846 147056 207902 147112
rect 207938 74976 207994 75032
rect 207846 46552 207902 46608
rect 209042 71712 209098 71768
rect 209226 76472 209282 76528
rect 208582 56480 208638 56536
rect 208950 56480 209006 56536
rect 208950 55800 209006 55856
rect 208490 51720 208546 51776
rect 208398 43424 208454 43480
rect 210054 147328 210110 147384
rect 209962 47504 210018 47560
rect 209870 43832 209926 43888
rect 209778 20576 209834 20632
rect 210146 77424 210202 77480
rect 210514 159296 210570 159352
rect 210330 77016 210386 77072
rect 210238 76880 210294 76936
rect 210054 24792 210110 24848
rect 210606 77832 210662 77888
rect 210698 42744 210754 42800
rect 211066 42744 211122 42800
rect 211066 42064 211122 42120
rect 211066 24792 211122 24848
rect 211066 24112 211122 24168
rect 211802 197920 211858 197976
rect 211802 73888 211858 73944
rect 211342 55120 211398 55176
rect 211342 54576 211398 54632
rect 211250 28872 211306 28928
rect 211158 21392 211214 21448
rect 211066 20576 211122 20632
rect 211066 19896 211122 19952
rect 212446 28872 212502 28928
rect 212446 28192 212502 28248
rect 212630 187312 212686 187368
rect 212998 77560 213054 77616
rect 213826 78104 213882 78160
rect 213826 77560 213882 77616
rect 213090 65456 213146 65512
rect 212722 64640 212778 64696
rect 212722 64096 212778 64152
rect 213918 62872 213974 62928
rect 212630 49544 212686 49600
rect 213826 49544 213882 49600
rect 213826 48864 213882 48920
rect 212538 21936 212594 21992
rect 213826 21936 213882 21992
rect 213826 21256 213882 21312
rect 215298 187176 215354 187232
rect 214102 142704 214158 142760
rect 214010 58928 214066 58984
rect 214194 77152 214250 77208
rect 214378 146920 214434 146976
rect 215574 186904 215630 186960
rect 215758 187040 215814 187096
rect 215758 74160 215814 74216
rect 215758 73616 215814 73672
rect 215574 68856 215630 68912
rect 215482 66952 215538 67008
rect 215390 64368 215446 64424
rect 215298 50904 215354 50960
rect 214102 37168 214158 37224
rect 214378 37168 214434 37224
rect 214378 36488 214434 36544
rect 213366 8880 213422 8936
rect 580170 192480 580226 192536
rect 218058 189624 218114 189680
rect 216862 73752 216918 73808
rect 218242 74160 218298 74216
rect 580170 179152 580226 179208
rect 580170 165824 580226 165880
rect 579986 152632 580042 152688
rect 580262 150456 580318 150512
rect 464342 140936 464398 140992
rect 218426 74296 218482 74352
rect 218334 74024 218390 74080
rect 224222 73616 224278 73672
rect 218426 73480 218482 73536
rect 218242 73344 218298 73400
rect 218150 73072 218206 73128
rect 218150 72392 218206 72448
rect 218058 45464 218114 45520
rect 220818 68856 220874 68912
rect 227718 66952 227774 67008
rect 237378 74296 237434 74352
rect 248418 74160 248474 74216
rect 242162 64368 242218 64424
rect 260102 76608 260158 76664
rect 256698 50632 256754 50688
rect 261482 73888 261538 73944
rect 288438 79464 288494 79520
rect 274638 78784 274694 78840
rect 275282 37848 275338 37904
rect 281538 58928 281594 58984
rect 279422 45192 279478 45248
rect 284298 56208 284354 56264
rect 293958 19896 294014 19952
rect 300858 42064 300914 42120
rect 309138 43696 309194 43752
rect 307022 28192 307078 28248
rect 310518 24112 310574 24168
rect 320178 52128 320234 52184
rect 579618 86128 579674 86184
rect 505098 80688 505154 80744
rect 332598 72392 332654 72448
rect 329102 21392 329158 21448
rect 338118 50496 338174 50552
rect 336738 21256 336794 21312
rect 347778 73752 347834 73808
rect 349158 57296 349214 57352
rect 356058 51992 356114 52048
rect 362958 64232 363014 64288
rect 364982 53352 365038 53408
rect 369858 54848 369914 54904
rect 373998 50360 374054 50416
rect 454682 75248 454738 75304
rect 380898 58792 380954 58848
rect 382922 56072 382978 56128
rect 387798 49136 387854 49192
rect 430578 69672 430634 69728
rect 402978 65456 403034 65512
rect 400862 51856 400918 51912
rect 405738 47776 405794 47832
rect 408498 43560 408554 43616
rect 418802 57160 418858 57216
rect 423770 46144 423826 46200
rect 425058 35128 425114 35184
rect 446402 62736 446458 62792
rect 432602 54712 432658 54768
rect 437478 53216 437534 53272
rect 440238 45056 440294 45112
rect 448518 58656 448574 58712
rect 450542 55936 450598 55992
rect 459558 61512 459614 61568
rect 468482 47640 468538 47696
rect 474738 53080 474794 53136
rect 500958 78104 501014 78160
rect 498198 71304 498254 71360
rect 484398 59880 484454 59936
rect 482282 55800 482338 55856
rect 489918 49000 489974 49056
rect 490010 47504 490066 47560
rect 507858 54576 507914 54632
rect 511998 64096 512054 64152
rect 514022 58520 514078 58576
rect 521658 75112 521714 75168
rect 520922 44920 520978 44976
rect 531318 71168 531374 71224
rect 528558 44784 528614 44840
rect 534722 43424 534778 43480
rect 534078 36488 534134 36544
rect 566462 76472 566518 76528
rect 549902 71032 549958 71088
rect 542358 51720 542414 51776
rect 547878 48864 547934 48920
rect 557538 69536 557594 69592
rect 556158 50224 556214 50280
rect 563702 61376 563758 61432
rect 560942 54440 560998 54496
rect 580170 72936 580226 72992
rect 574742 68176 574798 68232
rect 580354 143520 580410 143576
rect 580630 140800 580686 140856
rect 580906 125976 580962 126032
rect 580814 112784 580870 112840
rect 580722 99456 580778 99512
rect 581090 77968 581146 78024
rect 580998 77832 581054 77888
rect 580630 59608 580686 59664
rect 580538 46280 580594 46336
rect 580446 33088 580502 33144
rect 580354 19760 580410 19816
rect 580262 6568 580318 6624
<< metal3 >>
rect -960 697220 480 697460
rect 580165 697234 580231 697237
rect 583520 697234 584960 697324
rect 580165 697232 584960 697234
rect 580165 697176 580170 697232
rect 580226 697176 584960 697232
rect 580165 697174 584960 697176
rect 580165 697171 580231 697174
rect 583520 697084 584960 697174
rect -960 684314 480 684404
rect 3417 684314 3483 684317
rect -960 684312 3483 684314
rect -960 684256 3422 684312
rect 3478 684256 3483 684312
rect -960 684254 3483 684256
rect -960 684164 480 684254
rect 3417 684251 3483 684254
rect 580165 683906 580231 683909
rect 583520 683906 584960 683996
rect 580165 683904 584960 683906
rect 580165 683848 580170 683904
rect 580226 683848 584960 683904
rect 580165 683846 584960 683848
rect 580165 683843 580231 683846
rect 583520 683756 584960 683846
rect -960 671258 480 671348
rect 3509 671258 3575 671261
rect -960 671256 3575 671258
rect -960 671200 3514 671256
rect 3570 671200 3575 671256
rect -960 671198 3575 671200
rect -960 671108 480 671198
rect 3509 671195 3575 671198
rect 580165 670714 580231 670717
rect 583520 670714 584960 670804
rect 580165 670712 584960 670714
rect 580165 670656 580170 670712
rect 580226 670656 584960 670712
rect 580165 670654 584960 670656
rect 580165 670651 580231 670654
rect 583520 670564 584960 670654
rect -960 658202 480 658292
rect 3417 658202 3483 658205
rect -960 658200 3483 658202
rect -960 658144 3422 658200
rect 3478 658144 3483 658200
rect -960 658142 3483 658144
rect -960 658052 480 658142
rect 3417 658139 3483 658142
rect 583520 657236 584960 657476
rect -960 644996 480 645236
rect 580165 644058 580231 644061
rect 583520 644058 584960 644148
rect 580165 644056 584960 644058
rect 580165 644000 580170 644056
rect 580226 644000 584960 644056
rect 580165 643998 584960 644000
rect 580165 643995 580231 643998
rect 583520 643908 584960 643998
rect -960 632090 480 632180
rect 3417 632090 3483 632093
rect -960 632088 3483 632090
rect -960 632032 3422 632088
rect 3478 632032 3483 632088
rect -960 632030 3483 632032
rect -960 631940 480 632030
rect 3417 632027 3483 632030
rect 580165 630866 580231 630869
rect 583520 630866 584960 630956
rect 580165 630864 584960 630866
rect 580165 630808 580170 630864
rect 580226 630808 584960 630864
rect 580165 630806 584960 630808
rect 580165 630803 580231 630806
rect 583520 630716 584960 630806
rect -960 619170 480 619260
rect 3141 619170 3207 619173
rect -960 619168 3207 619170
rect -960 619112 3146 619168
rect 3202 619112 3207 619168
rect -960 619110 3207 619112
rect -960 619020 480 619110
rect 3141 619107 3207 619110
rect 580165 617538 580231 617541
rect 583520 617538 584960 617628
rect 580165 617536 584960 617538
rect 580165 617480 580170 617536
rect 580226 617480 584960 617536
rect 580165 617478 584960 617480
rect 580165 617475 580231 617478
rect 583520 617388 584960 617478
rect -960 606114 480 606204
rect 3233 606114 3299 606117
rect -960 606112 3299 606114
rect -960 606056 3238 606112
rect 3294 606056 3299 606112
rect -960 606054 3299 606056
rect -960 605964 480 606054
rect 3233 606051 3299 606054
rect 583520 604060 584960 604300
rect -960 592908 480 593148
rect 579797 591018 579863 591021
rect 583520 591018 584960 591108
rect 579797 591016 584960 591018
rect 579797 590960 579802 591016
rect 579858 590960 584960 591016
rect 579797 590958 584960 590960
rect 579797 590955 579863 590958
rect 583520 590868 584960 590958
rect -960 580002 480 580092
rect 3325 580002 3391 580005
rect -960 580000 3391 580002
rect -960 579944 3330 580000
rect 3386 579944 3391 580000
rect -960 579942 3391 579944
rect -960 579852 480 579942
rect 3325 579939 3391 579942
rect 580165 577690 580231 577693
rect 583520 577690 584960 577780
rect 580165 577688 584960 577690
rect 580165 577632 580170 577688
rect 580226 577632 584960 577688
rect 580165 577630 584960 577632
rect 580165 577627 580231 577630
rect 583520 577540 584960 577630
rect -960 566946 480 567036
rect 3417 566946 3483 566949
rect -960 566944 3483 566946
rect -960 566888 3422 566944
rect 3478 566888 3483 566944
rect -960 566886 3483 566888
rect -960 566796 480 566886
rect 3417 566883 3483 566886
rect 579797 564362 579863 564365
rect 583520 564362 584960 564452
rect 579797 564360 584960 564362
rect 579797 564304 579802 564360
rect 579858 564304 584960 564360
rect 579797 564302 584960 564304
rect 579797 564299 579863 564302
rect 583520 564212 584960 564302
rect -960 553890 480 553980
rect 3417 553890 3483 553893
rect -960 553888 3483 553890
rect -960 553832 3422 553888
rect 3478 553832 3483 553888
rect -960 553830 3483 553832
rect -960 553740 480 553830
rect 3417 553827 3483 553830
rect 583520 551020 584960 551260
rect -960 540684 480 540924
rect 580165 537842 580231 537845
rect 583520 537842 584960 537932
rect 580165 537840 584960 537842
rect 580165 537784 580170 537840
rect 580226 537784 584960 537840
rect 580165 537782 584960 537784
rect 580165 537779 580231 537782
rect 583520 537692 584960 537782
rect -960 527914 480 528004
rect 3417 527914 3483 527917
rect -960 527912 3483 527914
rect -960 527856 3422 527912
rect 3478 527856 3483 527912
rect -960 527854 3483 527856
rect -960 527764 480 527854
rect 3417 527851 3483 527854
rect 580165 524514 580231 524517
rect 583520 524514 584960 524604
rect 580165 524512 584960 524514
rect 580165 524456 580170 524512
rect 580226 524456 584960 524512
rect 580165 524454 584960 524456
rect 580165 524451 580231 524454
rect 583520 524364 584960 524454
rect -960 514858 480 514948
rect 3417 514858 3483 514861
rect -960 514856 3483 514858
rect -960 514800 3422 514856
rect 3478 514800 3483 514856
rect -960 514798 3483 514800
rect -960 514708 480 514798
rect 3417 514795 3483 514798
rect 580165 511322 580231 511325
rect 583520 511322 584960 511412
rect 580165 511320 584960 511322
rect 580165 511264 580170 511320
rect 580226 511264 584960 511320
rect 580165 511262 584960 511264
rect 580165 511259 580231 511262
rect 583520 511172 584960 511262
rect -960 501802 480 501892
rect 3049 501802 3115 501805
rect -960 501800 3115 501802
rect -960 501744 3054 501800
rect 3110 501744 3115 501800
rect -960 501742 3115 501744
rect -960 501652 480 501742
rect 3049 501739 3115 501742
rect 583520 497844 584960 498084
rect -960 488596 480 488836
rect 580165 484666 580231 484669
rect 583520 484666 584960 484756
rect 580165 484664 584960 484666
rect 580165 484608 580170 484664
rect 580226 484608 584960 484664
rect 580165 484606 584960 484608
rect 580165 484603 580231 484606
rect 583520 484516 584960 484606
rect -960 475690 480 475780
rect 3417 475690 3483 475693
rect -960 475688 3483 475690
rect -960 475632 3422 475688
rect 3478 475632 3483 475688
rect -960 475630 3483 475632
rect -960 475540 480 475630
rect 3417 475627 3483 475630
rect 579981 471474 580047 471477
rect 583520 471474 584960 471564
rect 579981 471472 584960 471474
rect 579981 471416 579986 471472
rect 580042 471416 584960 471472
rect 579981 471414 584960 471416
rect 579981 471411 580047 471414
rect 583520 471324 584960 471414
rect -960 462634 480 462724
rect 3509 462634 3575 462637
rect -960 462632 3575 462634
rect -960 462576 3514 462632
rect 3570 462576 3575 462632
rect -960 462574 3575 462576
rect -960 462484 480 462574
rect 3509 462571 3575 462574
rect 580165 458146 580231 458149
rect 583520 458146 584960 458236
rect 580165 458144 584960 458146
rect 580165 458088 580170 458144
rect 580226 458088 584960 458144
rect 580165 458086 584960 458088
rect 580165 458083 580231 458086
rect 583520 457996 584960 458086
rect -960 449578 480 449668
rect 3141 449578 3207 449581
rect -960 449576 3207 449578
rect -960 449520 3146 449576
rect 3202 449520 3207 449576
rect -960 449518 3207 449520
rect -960 449428 480 449518
rect 3141 449515 3207 449518
rect 583520 444668 584960 444908
rect -960 436508 480 436748
rect 580165 431626 580231 431629
rect 583520 431626 584960 431716
rect 580165 431624 584960 431626
rect 580165 431568 580170 431624
rect 580226 431568 584960 431624
rect 580165 431566 584960 431568
rect 580165 431563 580231 431566
rect 583520 431476 584960 431566
rect -960 423602 480 423692
rect 3509 423602 3575 423605
rect -960 423600 3575 423602
rect -960 423544 3514 423600
rect 3570 423544 3575 423600
rect -960 423542 3575 423544
rect -960 423452 480 423542
rect 3509 423539 3575 423542
rect 580165 418298 580231 418301
rect 583520 418298 584960 418388
rect 580165 418296 584960 418298
rect 580165 418240 580170 418296
rect 580226 418240 584960 418296
rect 580165 418238 584960 418240
rect 580165 418235 580231 418238
rect 583520 418148 584960 418238
rect -960 410546 480 410636
rect 2865 410546 2931 410549
rect -960 410544 2931 410546
rect -960 410488 2870 410544
rect 2926 410488 2931 410544
rect -960 410486 2931 410488
rect -960 410396 480 410486
rect 2865 410483 2931 410486
rect 580165 404970 580231 404973
rect 583520 404970 584960 405060
rect 580165 404968 584960 404970
rect 580165 404912 580170 404968
rect 580226 404912 584960 404968
rect 580165 404910 584960 404912
rect 580165 404907 580231 404910
rect 583520 404820 584960 404910
rect -960 397490 480 397580
rect 3509 397490 3575 397493
rect -960 397488 3575 397490
rect -960 397432 3514 397488
rect 3570 397432 3575 397488
rect -960 397430 3575 397432
rect -960 397340 480 397430
rect 3509 397427 3575 397430
rect 583520 391628 584960 391868
rect -960 384284 480 384524
rect 580165 378450 580231 378453
rect 583520 378450 584960 378540
rect 580165 378448 584960 378450
rect 580165 378392 580170 378448
rect 580226 378392 584960 378448
rect 580165 378390 584960 378392
rect 580165 378387 580231 378390
rect 583520 378300 584960 378390
rect -960 371378 480 371468
rect 2773 371378 2839 371381
rect -960 371376 2839 371378
rect -960 371320 2778 371376
rect 2834 371320 2839 371376
rect -960 371318 2839 371320
rect -960 371228 480 371318
rect 2773 371315 2839 371318
rect 580257 365122 580323 365125
rect 583520 365122 584960 365212
rect 580257 365120 584960 365122
rect 580257 365064 580262 365120
rect 580318 365064 584960 365120
rect 580257 365062 584960 365064
rect 580257 365059 580323 365062
rect 583520 364972 584960 365062
rect -960 358458 480 358548
rect 3141 358458 3207 358461
rect -960 358456 3207 358458
rect -960 358400 3146 358456
rect 3202 358400 3207 358456
rect -960 358398 3207 358400
rect -960 358308 480 358398
rect 3141 358395 3207 358398
rect 580165 351930 580231 351933
rect 583520 351930 584960 352020
rect 580165 351928 584960 351930
rect 580165 351872 580170 351928
rect 580226 351872 584960 351928
rect 580165 351870 584960 351872
rect 580165 351867 580231 351870
rect 583520 351780 584960 351870
rect -960 345402 480 345492
rect 3509 345402 3575 345405
rect -960 345400 3575 345402
rect -960 345344 3514 345400
rect 3570 345344 3575 345400
rect -960 345342 3575 345344
rect -960 345252 480 345342
rect 3509 345339 3575 345342
rect 583520 338452 584960 338692
rect -960 332196 480 332436
rect 580165 325274 580231 325277
rect 583520 325274 584960 325364
rect 580165 325272 584960 325274
rect 580165 325216 580170 325272
rect 580226 325216 584960 325272
rect 580165 325214 584960 325216
rect 580165 325211 580231 325214
rect 583520 325124 584960 325214
rect -960 319290 480 319380
rect 3325 319290 3391 319293
rect -960 319288 3391 319290
rect -960 319232 3330 319288
rect 3386 319232 3391 319288
rect -960 319230 3391 319232
rect -960 319140 480 319230
rect 3325 319227 3391 319230
rect 579981 312082 580047 312085
rect 583520 312082 584960 312172
rect 579981 312080 584960 312082
rect 579981 312024 579986 312080
rect 580042 312024 584960 312080
rect 579981 312022 584960 312024
rect 579981 312019 580047 312022
rect 583520 311932 584960 312022
rect -960 306234 480 306324
rect 3509 306234 3575 306237
rect -960 306232 3575 306234
rect -960 306176 3514 306232
rect 3570 306176 3575 306232
rect -960 306174 3575 306176
rect -960 306084 480 306174
rect 3509 306171 3575 306174
rect 580165 298754 580231 298757
rect 583520 298754 584960 298844
rect 580165 298752 584960 298754
rect 580165 298696 580170 298752
rect 580226 298696 584960 298752
rect 580165 298694 584960 298696
rect 580165 298691 580231 298694
rect 583520 298604 584960 298694
rect -960 293178 480 293268
rect 3509 293178 3575 293181
rect -960 293176 3575 293178
rect -960 293120 3514 293176
rect 3570 293120 3575 293176
rect -960 293118 3575 293120
rect -960 293028 480 293118
rect 3509 293115 3575 293118
rect 583520 285276 584960 285516
rect -960 279972 480 280212
rect 187734 278020 187740 278084
rect 187804 278082 187810 278084
rect 234613 278082 234679 278085
rect 187804 278080 234679 278082
rect 187804 278024 234618 278080
rect 234674 278024 234679 278080
rect 187804 278022 234679 278024
rect 187804 278020 187810 278022
rect 234613 278019 234679 278022
rect 156045 277538 156111 277541
rect 187734 277538 187740 277540
rect 156045 277536 187740 277538
rect 156045 277480 156050 277536
rect 156106 277480 187740 277536
rect 156045 277478 187740 277480
rect 156045 277475 156111 277478
rect 187734 277476 187740 277478
rect 187804 277476 187810 277540
rect 580165 272234 580231 272237
rect 583520 272234 584960 272324
rect 580165 272232 584960 272234
rect 580165 272176 580170 272232
rect 580226 272176 584960 272232
rect 580165 272174 584960 272176
rect 580165 272171 580231 272174
rect 583520 272084 584960 272174
rect -960 267202 480 267292
rect 3049 267202 3115 267205
rect -960 267200 3115 267202
rect -960 267144 3054 267200
rect 3110 267144 3115 267200
rect -960 267142 3115 267144
rect -960 267052 480 267142
rect 3049 267139 3115 267142
rect 111558 265100 111564 265164
rect 111628 265162 111634 265164
rect 135897 265162 135963 265165
rect 111628 265160 135963 265162
rect 111628 265104 135902 265160
rect 135958 265104 135963 265160
rect 111628 265102 135963 265104
rect 111628 265100 111634 265102
rect 135897 265099 135963 265102
rect 166257 265162 166323 265165
rect 192150 265162 192156 265164
rect 166257 265160 192156 265162
rect 166257 265104 166262 265160
rect 166318 265104 192156 265160
rect 166257 265102 192156 265104
rect 166257 265099 166323 265102
rect 192150 265100 192156 265102
rect 192220 265100 192226 265164
rect 108798 264964 108804 265028
rect 108868 265026 108874 265028
rect 138749 265026 138815 265029
rect 108868 265024 138815 265026
rect 108868 264968 138754 265024
rect 138810 264968 138815 265024
rect 108868 264966 138815 264968
rect 108868 264964 108874 264966
rect 138749 264963 138815 264966
rect 163497 265026 163563 265029
rect 196382 265026 196388 265028
rect 163497 265024 196388 265026
rect 163497 264968 163502 265024
rect 163558 264968 196388 265024
rect 163497 264966 196388 264968
rect 163497 264963 163563 264966
rect 196382 264964 196388 264966
rect 196452 264964 196458 265028
rect 116894 263740 116900 263804
rect 116964 263802 116970 263804
rect 137829 263802 137895 263805
rect 116964 263800 137895 263802
rect 116964 263744 137834 263800
rect 137890 263744 137895 263800
rect 116964 263742 137895 263744
rect 116964 263740 116970 263742
rect 137829 263739 137895 263742
rect 113030 263604 113036 263668
rect 113100 263666 113106 263668
rect 145281 263666 145347 263669
rect 145557 263666 145623 263669
rect 113100 263664 145623 263666
rect 113100 263608 145286 263664
rect 145342 263608 145562 263664
rect 145618 263608 145623 263664
rect 113100 263606 145623 263608
rect 113100 263604 113106 263606
rect 145281 263603 145347 263606
rect 145557 263603 145623 263606
rect 111190 263060 111196 263124
rect 111260 263122 111266 263124
rect 127341 263122 127407 263125
rect 111260 263120 127407 263122
rect 111260 263064 127346 263120
rect 127402 263064 127407 263120
rect 111260 263062 127407 263064
rect 111260 263060 111266 263062
rect 127341 263059 127407 263062
rect 191782 263060 191788 263124
rect 191852 263122 191858 263124
rect 282913 263122 282979 263125
rect 191852 263120 282979 263122
rect 191852 263064 282918 263120
rect 282974 263064 282979 263120
rect 191852 263062 282979 263064
rect 191852 263060 191858 263062
rect 282913 263059 282979 263062
rect 111006 262924 111012 262988
rect 111076 262986 111082 262988
rect 142245 262986 142311 262989
rect 142889 262986 142955 262989
rect 111076 262984 142955 262986
rect 111076 262928 142250 262984
rect 142306 262928 142894 262984
rect 142950 262928 142955 262984
rect 111076 262926 142955 262928
rect 111076 262924 111082 262926
rect 142245 262923 142311 262926
rect 142889 262923 142955 262926
rect 188521 262986 188587 262989
rect 347773 262986 347839 262989
rect 188521 262984 347839 262986
rect 188521 262928 188526 262984
rect 188582 262928 347778 262984
rect 347834 262928 347839 262984
rect 188521 262926 347839 262928
rect 188521 262923 188587 262926
rect 347773 262923 347839 262926
rect 112846 262788 112852 262852
rect 112916 262850 112922 262852
rect 146937 262850 147003 262853
rect 112916 262848 147003 262850
rect 112916 262792 146942 262848
rect 146998 262792 147003 262848
rect 112916 262790 147003 262792
rect 112916 262788 112922 262790
rect 146937 262787 147003 262790
rect 150893 262850 150959 262853
rect 192661 262850 192727 262853
rect 477493 262850 477559 262853
rect 150893 262848 477559 262850
rect 150893 262792 150898 262848
rect 150954 262792 192666 262848
rect 192722 262792 477498 262848
rect 477554 262792 477559 262848
rect 150893 262790 477559 262792
rect 150893 262787 150959 262790
rect 192661 262787 192727 262790
rect 477493 262787 477559 262790
rect 115790 262652 115796 262716
rect 115860 262714 115866 262716
rect 140313 262714 140379 262717
rect 115860 262712 140379 262714
rect 115860 262656 140318 262712
rect 140374 262656 140379 262712
rect 115860 262654 140379 262656
rect 115860 262652 115866 262654
rect 140313 262651 140379 262654
rect 164969 262714 165035 262717
rect 193622 262714 193628 262716
rect 164969 262712 193628 262714
rect 164969 262656 164974 262712
rect 165030 262656 193628 262712
rect 164969 262654 193628 262656
rect 164969 262651 165035 262654
rect 193622 262652 193628 262654
rect 193692 262652 193698 262716
rect 114134 262516 114140 262580
rect 114204 262578 114210 262580
rect 138657 262578 138723 262581
rect 114204 262576 138723 262578
rect 114204 262520 138662 262576
rect 138718 262520 138723 262576
rect 114204 262518 138723 262520
rect 114204 262516 114210 262518
rect 138657 262515 138723 262518
rect 153837 262578 153903 262581
rect 188061 262578 188127 262581
rect 188521 262578 188587 262581
rect 153837 262576 188587 262578
rect 153837 262520 153842 262576
rect 153898 262520 188066 262576
rect 188122 262520 188526 262576
rect 188582 262520 188587 262576
rect 153837 262518 188587 262520
rect 153837 262515 153903 262518
rect 188061 262515 188127 262518
rect 188521 262515 188587 262518
rect 111374 262380 111380 262444
rect 111444 262442 111450 262444
rect 125593 262442 125659 262445
rect 111444 262440 125659 262442
rect 111444 262384 125598 262440
rect 125654 262384 125659 262440
rect 111444 262382 125659 262384
rect 111444 262380 111450 262382
rect 125593 262379 125659 262382
rect 155861 262442 155927 262445
rect 190494 262442 190500 262444
rect 155861 262440 190500 262442
rect 155861 262384 155866 262440
rect 155922 262384 190500 262440
rect 155861 262382 190500 262384
rect 155861 262379 155927 262382
rect 190494 262380 190500 262382
rect 190564 262442 190570 262444
rect 191782 262442 191788 262444
rect 190564 262382 191788 262442
rect 190564 262380 190570 262382
rect 191782 262380 191788 262382
rect 191852 262380 191858 262444
rect 192334 262244 192340 262308
rect 192404 262306 192410 262308
rect 192477 262306 192543 262309
rect 192404 262304 192543 262306
rect 192404 262248 192482 262304
rect 192538 262248 192543 262304
rect 192404 262246 192543 262248
rect 192404 262244 192410 262246
rect 192477 262243 192543 262246
rect 112662 261020 112668 261084
rect 112732 261082 112738 261084
rect 137461 261082 137527 261085
rect 112732 261080 137527 261082
rect 112732 261024 137466 261080
rect 137522 261024 137527 261080
rect 112732 261022 137527 261024
rect 112732 261020 112738 261022
rect 137461 261019 137527 261022
rect 158713 260946 158779 260949
rect 193438 260946 193444 260948
rect 158713 260944 193444 260946
rect 158713 260888 158718 260944
rect 158774 260888 193444 260944
rect 158713 260886 193444 260888
rect 158713 260883 158779 260886
rect 193438 260884 193444 260886
rect 193508 260884 193514 260948
rect 122782 260748 122788 260812
rect 122852 260810 122858 260812
rect 123201 260810 123267 260813
rect 122852 260808 123267 260810
rect 122852 260752 123206 260808
rect 123262 260752 123267 260808
rect 122852 260750 123267 260752
rect 122852 260748 122858 260750
rect 123201 260747 123267 260750
rect 116710 260476 116716 260540
rect 116780 260538 116786 260540
rect 127617 260538 127683 260541
rect 116780 260536 127683 260538
rect 116780 260480 127622 260536
rect 127678 260480 127683 260536
rect 116780 260478 127683 260480
rect 116780 260476 116786 260478
rect 127617 260475 127683 260478
rect 115606 260340 115612 260404
rect 115676 260402 115682 260404
rect 115676 260342 147138 260402
rect 115676 260340 115682 260342
rect 121126 260204 121132 260268
rect 121196 260266 121202 260268
rect 143625 260266 143691 260269
rect 144499 260266 144565 260269
rect 121196 260264 144565 260266
rect 121196 260208 143630 260264
rect 143686 260208 144504 260264
rect 144560 260208 144565 260264
rect 121196 260206 144565 260208
rect 147078 260266 147138 260342
rect 149053 260266 149119 260269
rect 150019 260266 150085 260269
rect 147078 260264 150085 260266
rect 147078 260208 149058 260264
rect 149114 260208 150024 260264
rect 150080 260208 150085 260264
rect 147078 260206 150085 260208
rect 121196 260204 121202 260206
rect 143625 260203 143691 260206
rect 144499 260203 144565 260206
rect 149053 260203 149119 260206
rect 150019 260203 150085 260206
rect 155953 260266 156019 260269
rect 156643 260266 156709 260269
rect 155953 260264 156709 260266
rect 155953 260208 155958 260264
rect 156014 260208 156648 260264
rect 156704 260208 156709 260264
rect 155953 260206 156709 260208
rect 155953 260203 156019 260206
rect 156643 260203 156709 260206
rect 160093 260266 160159 260269
rect 161059 260266 161125 260269
rect 160093 260264 161125 260266
rect 160093 260208 160098 260264
rect 160154 260208 161064 260264
rect 161120 260208 161125 260264
rect 160093 260206 161125 260208
rect 160093 260203 160159 260206
rect 161059 260203 161125 260206
rect 116526 260068 116532 260132
rect 116596 260130 116602 260132
rect 127249 260130 127315 260133
rect 116596 260128 127315 260130
rect 116596 260072 127254 260128
rect 127310 260072 127315 260128
rect 116596 260070 127315 260072
rect 116596 260068 116602 260070
rect 127249 260067 127315 260070
rect 127617 260130 127683 260133
rect 140773 260130 140839 260133
rect 141739 260130 141805 260133
rect 127617 260128 141805 260130
rect 127617 260072 127622 260128
rect 127678 260072 140778 260128
rect 140834 260072 141744 260128
rect 141800 260072 141805 260128
rect 127617 260070 141805 260072
rect 127617 260067 127683 260070
rect 140773 260067 140839 260070
rect 141739 260067 141805 260070
rect 166027 260130 166093 260133
rect 189717 260130 189783 260133
rect 166027 260128 189783 260130
rect 166027 260072 166032 260128
rect 166088 260072 189722 260128
rect 189778 260072 189783 260128
rect 166027 260070 189783 260072
rect 166027 260067 166093 260070
rect 189717 260067 189783 260070
rect 121310 259932 121316 259996
rect 121380 259994 121386 259996
rect 147673 259994 147739 259997
rect 121380 259992 147739 259994
rect 121380 259936 147678 259992
rect 147734 259936 147739 259992
rect 121380 259934 147739 259936
rect 121380 259932 121386 259934
rect 147673 259931 147739 259934
rect 161197 259994 161263 259997
rect 188889 259994 188955 259997
rect 161197 259992 188955 259994
rect 161197 259936 161202 259992
rect 161258 259936 188894 259992
rect 188950 259936 188955 259992
rect 161197 259934 188955 259936
rect 161197 259931 161263 259934
rect 188889 259931 188955 259934
rect 118182 259796 118188 259860
rect 118252 259858 118258 259860
rect 144913 259858 144979 259861
rect 118252 259856 144979 259858
rect 118252 259800 144918 259856
rect 144974 259800 144979 259856
rect 118252 259798 144979 259800
rect 118252 259796 118258 259798
rect 144913 259795 144979 259798
rect 156873 259858 156939 259861
rect 189022 259858 189028 259860
rect 156873 259856 189028 259858
rect 156873 259800 156878 259856
rect 156934 259800 189028 259856
rect 156873 259798 189028 259800
rect 156873 259795 156939 259798
rect 189022 259796 189028 259798
rect 189092 259796 189098 259860
rect 124857 259722 124923 259725
rect 122790 259720 124923 259722
rect 122790 259664 124862 259720
rect 124918 259664 124923 259720
rect 122790 259662 124923 259664
rect 113950 259524 113956 259588
rect 114020 259586 114026 259588
rect 122790 259586 122850 259662
rect 124857 259659 124923 259662
rect 127249 259722 127315 259725
rect 148133 259722 148199 259725
rect 127249 259720 148199 259722
rect 127249 259664 127254 259720
rect 127310 259664 148138 259720
rect 148194 259664 148199 259720
rect 127249 259662 148199 259664
rect 127249 259659 127315 259662
rect 148133 259659 148199 259662
rect 155217 259722 155283 259725
rect 189206 259722 189212 259724
rect 155217 259720 189212 259722
rect 155217 259664 155222 259720
rect 155278 259664 189212 259720
rect 155217 259662 189212 259664
rect 155217 259659 155283 259662
rect 189206 259660 189212 259662
rect 189276 259660 189282 259724
rect 114020 259526 122850 259586
rect 123293 259586 123359 259589
rect 124070 259586 124076 259588
rect 123293 259584 124076 259586
rect 123293 259528 123298 259584
rect 123354 259528 124076 259584
rect 123293 259526 124076 259528
rect 114020 259524 114026 259526
rect 123293 259523 123359 259526
rect 124070 259524 124076 259526
rect 124140 259524 124146 259588
rect 164601 259586 164667 259589
rect 201861 259586 201927 259589
rect 164601 259584 201927 259586
rect 164601 259528 164606 259584
rect 164662 259528 201866 259584
rect 201922 259528 201927 259584
rect 164601 259526 201927 259528
rect 164601 259523 164667 259526
rect 201861 259523 201927 259526
rect 122966 259388 122972 259452
rect 123036 259450 123042 259452
rect 123753 259450 123819 259453
rect 123036 259448 123819 259450
rect 123036 259392 123758 259448
rect 123814 259392 123819 259448
rect 123036 259390 123819 259392
rect 123036 259388 123042 259390
rect 123753 259387 123819 259390
rect 185669 259450 185735 259453
rect 186078 259450 186084 259452
rect 185669 259448 186084 259450
rect 185669 259392 185674 259448
rect 185730 259392 186084 259448
rect 185669 259390 186084 259392
rect 185669 259387 185735 259390
rect 186078 259388 186084 259390
rect 186148 259388 186154 259452
rect 580165 258906 580231 258909
rect 583520 258906 584960 258996
rect 580165 258904 584960 258906
rect 580165 258848 580170 258904
rect 580226 258848 584960 258904
rect 580165 258846 584960 258848
rect 580165 258843 580231 258846
rect 583520 258756 584960 258846
rect -960 254146 480 254236
rect 3509 254146 3575 254149
rect -960 254144 3575 254146
rect -960 254088 3514 254144
rect 3570 254088 3575 254144
rect -960 254086 3575 254088
rect -960 253996 480 254086
rect 3509 254083 3575 254086
rect 580165 245578 580231 245581
rect 583520 245578 584960 245668
rect 580165 245576 584960 245578
rect 580165 245520 580170 245576
rect 580226 245520 584960 245576
rect 580165 245518 584960 245520
rect 580165 245515 580231 245518
rect 583520 245428 584960 245518
rect -960 241090 480 241180
rect 2773 241090 2839 241093
rect -960 241088 2839 241090
rect -960 241032 2778 241088
rect 2834 241032 2839 241088
rect -960 241030 2839 241032
rect -960 240940 480 241030
rect 2773 241027 2839 241030
rect 580441 232386 580507 232389
rect 583520 232386 584960 232476
rect 580441 232384 584960 232386
rect 580441 232328 580446 232384
rect 580502 232328 584960 232384
rect 580441 232326 584960 232328
rect 580441 232323 580507 232326
rect 583520 232236 584960 232326
rect -960 227884 480 228124
rect 580349 219058 580415 219061
rect 583520 219058 584960 219148
rect 580349 219056 584960 219058
rect 580349 219000 580354 219056
rect 580410 219000 584960 219056
rect 580349 218998 584960 219000
rect 580349 218995 580415 218998
rect 583520 218908 584960 218998
rect -960 214978 480 215068
rect 3509 214978 3575 214981
rect -960 214976 3575 214978
rect -960 214920 3514 214976
rect 3570 214920 3575 214976
rect -960 214918 3575 214920
rect -960 214828 480 214918
rect 3509 214915 3575 214918
rect 186078 213828 186084 213892
rect 186148 213890 186154 213892
rect 187417 213890 187483 213893
rect 186148 213888 187483 213890
rect 186148 213832 187422 213888
rect 187478 213832 187483 213888
rect 186148 213830 187483 213832
rect 186148 213828 186154 213830
rect 187417 213827 187483 213830
rect 579797 205730 579863 205733
rect 583520 205730 584960 205820
rect 579797 205728 584960 205730
rect 579797 205672 579802 205728
rect 579858 205672 584960 205728
rect 579797 205670 584960 205672
rect 579797 205667 579863 205670
rect 583520 205580 584960 205670
rect -960 201922 480 202012
rect 3417 201922 3483 201925
rect -960 201920 3483 201922
rect -960 201864 3422 201920
rect 3478 201864 3483 201920
rect -960 201862 3483 201864
rect -960 201772 480 201862
rect 3417 201859 3483 201862
rect 131614 201452 131620 201516
rect 131684 201514 131690 201516
rect 139526 201514 139532 201516
rect 131684 201454 139532 201514
rect 131684 201452 131690 201454
rect 139526 201452 139532 201454
rect 139596 201452 139602 201516
rect 128997 200698 129063 200701
rect 154614 200698 154620 200700
rect 128997 200696 154620 200698
rect 128997 200640 129002 200696
rect 129058 200640 154620 200696
rect 128997 200638 154620 200640
rect 128997 200635 129063 200638
rect 154614 200636 154620 200638
rect 154684 200636 154690 200700
rect 173566 200636 173572 200700
rect 173636 200698 173642 200700
rect 178217 200698 178283 200701
rect 173636 200696 178283 200698
rect 173636 200640 178222 200696
rect 178278 200640 178283 200696
rect 173636 200638 178283 200640
rect 173636 200636 173642 200638
rect 178217 200635 178283 200638
rect 124857 200562 124923 200565
rect 150934 200562 150940 200564
rect 124857 200560 150940 200562
rect 124857 200504 124862 200560
rect 124918 200504 150940 200560
rect 124857 200502 150940 200504
rect 124857 200499 124923 200502
rect 150934 200500 150940 200502
rect 151004 200500 151010 200564
rect 163078 200500 163084 200564
rect 163148 200562 163154 200564
rect 198365 200562 198431 200565
rect 163148 200560 198431 200562
rect 163148 200504 198370 200560
rect 198426 200504 198431 200560
rect 163148 200502 198431 200504
rect 163148 200500 163154 200502
rect 198365 200499 198431 200502
rect 106774 200364 106780 200428
rect 106844 200426 106850 200428
rect 106844 200366 135178 200426
rect 106844 200364 106850 200366
rect 122782 200092 122788 200156
rect 122852 200154 122858 200156
rect 124029 200154 124095 200157
rect 122852 200152 124095 200154
rect 122852 200096 124034 200152
rect 124090 200096 124095 200152
rect 122852 200094 124095 200096
rect 122852 200092 122858 200094
rect 124029 200091 124095 200094
rect 130929 200154 130995 200157
rect 130929 200152 134442 200154
rect 130929 200096 130934 200152
rect 130990 200096 134442 200152
rect 130929 200094 134442 200096
rect 130929 200091 130995 200094
rect 134382 199919 134442 200094
rect 132723 199914 132789 199919
rect 134103 199916 134169 199919
rect 132723 199884 132728 199914
rect 132784 199884 132789 199914
rect 134060 199914 134169 199916
rect 133827 199884 133893 199885
rect 132718 199820 132724 199884
rect 132788 199882 132794 199884
rect 132788 199822 132846 199882
rect 132788 199820 132794 199822
rect 133822 199820 133828 199884
rect 133892 199882 133898 199884
rect 133892 199822 133984 199882
rect 134060 199858 134108 199914
rect 134164 199858 134169 199914
rect 134060 199853 134169 199858
rect 134379 199914 134445 199919
rect 134379 199858 134384 199914
rect 134440 199858 134445 199914
rect 134379 199853 134445 199858
rect 134563 199914 134629 199919
rect 134839 199916 134905 199919
rect 134563 199858 134568 199914
rect 134624 199858 134629 199914
rect 134796 199914 134905 199916
rect 134796 199884 134844 199914
rect 134563 199853 134629 199858
rect 133892 199820 133898 199822
rect 133827 199819 133893 199820
rect 133643 199778 133709 199783
rect 133643 199748 133648 199778
rect 133704 199748 133709 199778
rect 134060 199749 134120 199853
rect 134566 199749 134626 199853
rect 134742 199820 134748 199884
rect 134812 199858 134844 199884
rect 134900 199858 134905 199914
rect 134812 199853 134905 199858
rect 134812 199822 134856 199853
rect 134812 199820 134818 199822
rect 133638 199684 133644 199748
rect 133708 199746 133714 199748
rect 133708 199686 133766 199746
rect 134057 199744 134123 199749
rect 134057 199688 134062 199744
rect 134118 199688 134123 199744
rect 133708 199684 133714 199686
rect 134057 199683 134123 199688
rect 134517 199744 134626 199749
rect 134517 199688 134522 199744
rect 134578 199688 134626 199744
rect 134517 199686 134626 199688
rect 135118 199746 135178 200366
rect 171174 200364 171180 200428
rect 171244 200426 171250 200428
rect 181437 200426 181503 200429
rect 171244 200424 181503 200426
rect 171244 200368 181442 200424
rect 181498 200368 181503 200424
rect 171244 200366 181503 200368
rect 171244 200364 171250 200366
rect 181437 200363 181503 200366
rect 200389 200290 200455 200293
rect 166076 200288 200455 200290
rect 166076 200232 200394 200288
rect 200450 200232 200455 200288
rect 166076 200230 200455 200232
rect 142286 200154 142292 200156
rect 139764 200094 142292 200154
rect 135851 199914 135917 199919
rect 135483 199884 135549 199885
rect 135478 199882 135484 199884
rect 135392 199822 135484 199882
rect 135478 199820 135484 199822
rect 135548 199820 135554 199884
rect 135667 199880 135733 199885
rect 135851 199884 135856 199914
rect 135912 199884 135917 199914
rect 136219 199914 136285 199919
rect 135667 199824 135672 199880
rect 135728 199824 135733 199880
rect 135483 199819 135549 199820
rect 135667 199819 135733 199824
rect 135846 199820 135852 199884
rect 135916 199882 135922 199884
rect 135916 199822 135974 199882
rect 136219 199858 136224 199914
rect 136280 199858 136285 199914
rect 136219 199853 136285 199858
rect 136403 199914 136469 199919
rect 136863 199916 136929 199919
rect 136403 199858 136408 199914
rect 136464 199858 136469 199914
rect 136403 199853 136469 199858
rect 136820 199914 136929 199916
rect 136820 199858 136868 199914
rect 136924 199858 136929 199914
rect 136820 199853 136929 199858
rect 137415 199916 137481 199919
rect 139623 199916 139689 199919
rect 139764 199916 139824 200094
rect 142286 200092 142292 200094
rect 142356 200092 142362 200156
rect 150014 200092 150020 200156
rect 150084 200154 150090 200156
rect 150084 200094 157626 200154
rect 150084 200092 150090 200094
rect 152046 199958 157074 200018
rect 137415 199914 137662 199916
rect 137415 199858 137420 199914
rect 137476 199858 137662 199914
rect 139623 199914 139824 199916
rect 137415 199856 137662 199858
rect 137415 199853 137481 199856
rect 135916 199820 135922 199822
rect 135670 199749 135730 199819
rect 136222 199749 136282 199853
rect 136406 199749 136466 199853
rect 135345 199746 135411 199749
rect 135118 199744 135411 199746
rect 135118 199688 135350 199744
rect 135406 199688 135411 199744
rect 135118 199686 135411 199688
rect 135670 199744 135779 199749
rect 135670 199688 135718 199744
rect 135774 199688 135779 199744
rect 135670 199686 135779 199688
rect 134517 199683 134583 199686
rect 135345 199683 135411 199686
rect 135713 199683 135779 199686
rect 136173 199744 136282 199749
rect 136173 199688 136178 199744
rect 136234 199688 136282 199744
rect 136173 199686 136282 199688
rect 136357 199744 136466 199749
rect 136357 199688 136362 199744
rect 136418 199688 136466 199744
rect 136357 199686 136466 199688
rect 136173 199683 136239 199686
rect 136357 199683 136423 199686
rect 107285 199610 107351 199613
rect 136820 199610 136880 199853
rect 137139 199748 137205 199749
rect 137134 199746 137140 199748
rect 137048 199686 137140 199746
rect 137134 199684 137140 199686
rect 137204 199684 137210 199748
rect 137139 199683 137205 199684
rect 107285 199608 136880 199610
rect 107285 199552 107290 199608
rect 107346 199552 136880 199608
rect 107285 199550 136880 199552
rect 137461 199610 137527 199613
rect 137602 199610 137662 199856
rect 138238 199820 138244 199884
rect 138308 199882 138314 199884
rect 138611 199882 138677 199885
rect 138308 199880 138677 199882
rect 138308 199824 138616 199880
rect 138672 199824 138677 199880
rect 139623 199858 139628 199914
rect 139684 199858 139824 199914
rect 139623 199856 139824 199858
rect 140267 199914 140333 199919
rect 140267 199858 140272 199914
rect 140328 199858 140333 199914
rect 139623 199853 139689 199856
rect 140267 199853 140333 199858
rect 140635 199914 140701 199919
rect 140911 199916 140977 199919
rect 141095 199916 141161 199919
rect 140635 199858 140640 199914
rect 140696 199858 140701 199914
rect 140635 199853 140701 199858
rect 140776 199914 140977 199916
rect 140776 199858 140916 199914
rect 140972 199858 140977 199914
rect 140776 199856 140977 199858
rect 138308 199822 138677 199824
rect 138308 199820 138314 199822
rect 138611 199819 138677 199822
rect 137737 199746 137803 199749
rect 137870 199746 137876 199748
rect 137737 199744 137876 199746
rect 137737 199688 137742 199744
rect 137798 199688 137876 199744
rect 137737 199686 137876 199688
rect 137737 199683 137803 199686
rect 137870 199684 137876 199686
rect 137940 199684 137946 199748
rect 138749 199746 138815 199749
rect 138749 199744 138858 199746
rect 138749 199688 138754 199744
rect 138810 199688 138858 199744
rect 138749 199683 138858 199688
rect 139526 199684 139532 199748
rect 139596 199746 139602 199748
rect 139669 199746 139735 199749
rect 139596 199744 139735 199746
rect 139596 199688 139674 199744
rect 139730 199688 139735 199744
rect 139596 199686 139735 199688
rect 139596 199684 139602 199686
rect 139669 199683 139735 199686
rect 137461 199608 137662 199610
rect 137461 199552 137466 199608
rect 137522 199552 137662 199608
rect 137461 199550 137662 199552
rect 137829 199610 137895 199613
rect 138798 199610 138858 199683
rect 137829 199608 138858 199610
rect 137829 199552 137834 199608
rect 137890 199552 138858 199608
rect 137829 199550 138858 199552
rect 107285 199547 107351 199550
rect 137461 199547 137527 199550
rect 137829 199547 137895 199550
rect 139526 199548 139532 199612
rect 139596 199610 139602 199612
rect 140270 199610 140330 199853
rect 139596 199550 140330 199610
rect 140638 199610 140698 199853
rect 140776 199746 140836 199856
rect 140911 199853 140977 199856
rect 141052 199914 141161 199916
rect 141052 199858 141100 199914
rect 141156 199882 141161 199914
rect 141371 199914 141437 199919
rect 141156 199858 141250 199882
rect 141052 199822 141250 199858
rect 141371 199858 141376 199914
rect 141432 199858 141437 199914
rect 141555 199914 141621 199919
rect 141555 199884 141560 199914
rect 141616 199884 141621 199914
rect 141831 199916 141897 199919
rect 141831 199914 141940 199916
rect 141371 199853 141437 199858
rect 140957 199746 141023 199749
rect 140776 199744 141023 199746
rect 140776 199688 140962 199744
rect 141018 199688 141023 199744
rect 140776 199686 141023 199688
rect 140957 199683 141023 199686
rect 141190 199613 141250 199822
rect 141374 199749 141434 199853
rect 141550 199820 141556 199884
rect 141620 199882 141626 199884
rect 141620 199822 141678 199882
rect 141831 199858 141836 199914
rect 141892 199858 141940 199914
rect 142107 199914 142173 199919
rect 142107 199884 142112 199914
rect 142168 199884 142173 199914
rect 142291 199914 142357 199919
rect 141831 199853 141940 199858
rect 141620 199820 141626 199822
rect 141880 199749 141940 199853
rect 142102 199820 142108 199884
rect 142172 199882 142178 199884
rect 142172 199822 142230 199882
rect 142291 199858 142296 199914
rect 142352 199858 142357 199914
rect 142291 199853 142357 199858
rect 142475 199914 142541 199919
rect 142475 199858 142480 199914
rect 142536 199882 142541 199914
rect 142843 199914 142909 199919
rect 142654 199882 142660 199884
rect 142536 199858 142660 199882
rect 142475 199853 142660 199858
rect 142172 199820 142178 199822
rect 141325 199744 141434 199749
rect 141325 199688 141330 199744
rect 141386 199688 141434 199744
rect 141325 199686 141434 199688
rect 141601 199746 141667 199749
rect 141734 199746 141740 199748
rect 141601 199744 141740 199746
rect 141601 199688 141606 199744
rect 141662 199688 141740 199744
rect 141601 199686 141740 199688
rect 141325 199683 141391 199686
rect 141601 199683 141667 199686
rect 141734 199684 141740 199686
rect 141804 199684 141810 199748
rect 141877 199744 141943 199749
rect 141877 199688 141882 199744
rect 141938 199688 141943 199744
rect 141877 199683 141943 199688
rect 142061 199746 142127 199749
rect 142294 199746 142354 199853
rect 142478 199822 142660 199853
rect 142654 199820 142660 199822
rect 142724 199820 142730 199884
rect 142843 199858 142848 199914
rect 142904 199858 142909 199914
rect 142843 199853 142909 199858
rect 143027 199914 143093 199919
rect 143855 199916 143921 199919
rect 143027 199858 143032 199914
rect 143088 199882 143093 199914
rect 143628 199914 143921 199916
rect 143206 199882 143212 199884
rect 143088 199858 143212 199882
rect 143027 199853 143212 199858
rect 142846 199749 142906 199853
rect 143030 199822 143212 199853
rect 143206 199820 143212 199822
rect 143276 199820 143282 199884
rect 143390 199820 143396 199884
rect 143460 199882 143466 199884
rect 143628 199882 143860 199914
rect 143460 199858 143860 199882
rect 143916 199858 143921 199914
rect 143460 199856 143921 199858
rect 143460 199822 143688 199856
rect 143855 199853 143921 199856
rect 144867 199914 144933 199919
rect 144867 199858 144872 199914
rect 144928 199858 144933 199914
rect 144867 199853 144933 199858
rect 145971 199914 146037 199919
rect 146247 199916 146313 199919
rect 145971 199858 145976 199914
rect 146032 199858 146037 199914
rect 146204 199914 146313 199916
rect 146204 199884 146252 199914
rect 145971 199853 146037 199858
rect 143460 199820 143466 199822
rect 144870 199749 144930 199853
rect 142061 199744 142354 199746
rect 142061 199688 142066 199744
rect 142122 199688 142354 199744
rect 142061 199686 142354 199688
rect 142475 199746 142541 199749
rect 142475 199744 142676 199746
rect 142475 199688 142480 199744
rect 142536 199688 142676 199744
rect 142475 199686 142676 199688
rect 142846 199744 142955 199749
rect 142846 199688 142894 199744
rect 142950 199688 142955 199744
rect 142846 199686 142955 199688
rect 142061 199683 142127 199686
rect 142475 199683 142541 199686
rect 140773 199610 140839 199613
rect 140638 199608 140839 199610
rect 140638 199552 140778 199608
rect 140834 199552 140839 199608
rect 140638 199550 140839 199552
rect 141190 199608 141299 199613
rect 141190 199552 141238 199608
rect 141294 199552 141299 199608
rect 141190 199550 141299 199552
rect 139596 199548 139602 199550
rect 140773 199547 140839 199550
rect 141233 199547 141299 199550
rect 141601 199610 141667 199613
rect 142470 199610 142476 199612
rect 141601 199608 142476 199610
rect 141601 199552 141606 199608
rect 141662 199552 142476 199608
rect 141601 199550 142476 199552
rect 141601 199547 141667 199550
rect 142470 199548 142476 199550
rect 142540 199548 142546 199612
rect 142616 199610 142676 199686
rect 142889 199683 142955 199686
rect 143022 199684 143028 199748
rect 143092 199746 143098 199748
rect 143395 199746 143461 199749
rect 143092 199744 143461 199746
rect 143092 199688 143400 199744
rect 143456 199688 143461 199744
rect 143092 199686 143461 199688
rect 143092 199684 143098 199686
rect 143395 199683 143461 199686
rect 144821 199744 144930 199749
rect 144821 199688 144826 199744
rect 144882 199688 144930 199744
rect 144821 199686 144930 199688
rect 144821 199683 144887 199686
rect 145974 199613 146034 199853
rect 146150 199820 146156 199884
rect 146220 199858 146252 199884
rect 146308 199858 146313 199914
rect 147443 199914 147509 199919
rect 147443 199882 147448 199914
rect 146220 199853 146313 199858
rect 146526 199858 147448 199882
rect 147504 199858 147509 199914
rect 146526 199853 147509 199858
rect 147627 199914 147693 199919
rect 147627 199858 147632 199914
rect 147688 199858 147693 199914
rect 147627 199853 147693 199858
rect 147995 199914 148061 199919
rect 147995 199858 148000 199914
rect 148056 199858 148061 199914
rect 148547 199914 148613 199919
rect 147995 199853 148061 199858
rect 148271 199882 148337 199885
rect 148271 199880 148380 199882
rect 146220 199822 146264 199853
rect 146526 199822 147506 199853
rect 146220 199820 146226 199822
rect 143349 199610 143415 199613
rect 142616 199608 143415 199610
rect 142616 199552 143354 199608
rect 143410 199552 143415 199608
rect 142616 199550 143415 199552
rect 143349 199547 143415 199550
rect 145925 199608 146034 199613
rect 145925 199552 145930 199608
rect 145986 199552 146034 199608
rect 145925 199550 146034 199552
rect 146385 199610 146451 199613
rect 146526 199610 146586 199822
rect 146385 199608 146586 199610
rect 146385 199552 146390 199608
rect 146446 199552 146586 199608
rect 146385 199550 146586 199552
rect 145925 199547 145991 199550
rect 146385 199547 146451 199550
rect 147438 199548 147444 199612
rect 147508 199610 147514 199612
rect 147630 199610 147690 199853
rect 147508 199550 147690 199610
rect 147857 199610 147923 199613
rect 147998 199610 148058 199853
rect 148271 199824 148276 199880
rect 148332 199824 148380 199880
rect 148547 199858 148552 199914
rect 148608 199858 148613 199914
rect 151123 199914 151189 199919
rect 148547 199853 148613 199858
rect 150571 199880 150637 199885
rect 148271 199819 148380 199824
rect 148320 199749 148380 199819
rect 148317 199744 148383 199749
rect 148317 199688 148322 199744
rect 148378 199688 148383 199744
rect 148317 199683 148383 199688
rect 147857 199608 148058 199610
rect 147857 199552 147862 199608
rect 147918 199552 148058 199608
rect 147857 199550 148058 199552
rect 148550 199613 148610 199853
rect 150571 199824 150576 199880
rect 150632 199824 150637 199880
rect 151123 199858 151128 199914
rect 151184 199858 151189 199914
rect 151123 199853 151189 199858
rect 151675 199914 151741 199919
rect 151675 199858 151680 199914
rect 151736 199858 151741 199914
rect 151859 199914 151925 199919
rect 151859 199884 151864 199914
rect 151920 199884 151925 199914
rect 152046 199885 152106 199958
rect 151675 199853 151741 199858
rect 150571 199819 150637 199824
rect 148550 199608 148659 199613
rect 148550 199552 148598 199608
rect 148654 199552 148659 199608
rect 148550 199550 148659 199552
rect 150574 199610 150634 199819
rect 151126 199749 151186 199853
rect 151678 199749 151738 199853
rect 151854 199820 151860 199884
rect 151924 199882 151930 199884
rect 151924 199822 151982 199882
rect 152043 199880 152109 199885
rect 152043 199824 152048 199880
rect 152104 199824 152109 199880
rect 151924 199820 151930 199822
rect 152043 199819 152109 199824
rect 152963 199882 153029 199885
rect 152963 199880 153394 199882
rect 152963 199824 152968 199880
rect 153024 199824 153394 199880
rect 152963 199822 153394 199824
rect 152963 199819 153029 199822
rect 151126 199744 151235 199749
rect 151126 199688 151174 199744
rect 151230 199688 151235 199744
rect 151126 199686 151235 199688
rect 151678 199744 151787 199749
rect 151678 199688 151726 199744
rect 151782 199688 151787 199744
rect 151678 199686 151787 199688
rect 151169 199683 151235 199686
rect 151721 199683 151787 199686
rect 150709 199610 150775 199613
rect 150574 199608 150775 199610
rect 150574 199552 150714 199608
rect 150770 199552 150775 199608
rect 150574 199550 150775 199552
rect 147508 199548 147514 199550
rect 147857 199547 147923 199550
rect 148593 199547 148659 199550
rect 150709 199547 150775 199550
rect 150934 199548 150940 199612
rect 151004 199610 151010 199612
rect 153193 199610 153259 199613
rect 151004 199608 153259 199610
rect 151004 199552 153198 199608
rect 153254 199552 153259 199608
rect 151004 199550 153259 199552
rect 151004 199548 151010 199550
rect 153193 199547 153259 199550
rect 117078 199412 117084 199476
rect 117148 199474 117154 199476
rect 151537 199474 151603 199477
rect 117148 199472 151603 199474
rect 117148 199416 151542 199472
rect 151598 199416 151603 199472
rect 117148 199414 151603 199416
rect 117148 199412 117154 199414
rect 151537 199411 151603 199414
rect 153009 199474 153075 199477
rect 153334 199474 153394 199822
rect 154614 199820 154620 199884
rect 154684 199882 154690 199884
rect 154803 199882 154869 199885
rect 155263 199882 155329 199885
rect 154684 199880 154869 199882
rect 154684 199824 154808 199880
rect 154864 199824 154869 199880
rect 154684 199822 154869 199824
rect 154684 199820 154690 199822
rect 154803 199819 154869 199822
rect 154990 199880 155329 199882
rect 154990 199824 155268 199880
rect 155324 199824 155329 199880
rect 154990 199822 155329 199824
rect 154990 199746 155050 199822
rect 155263 199819 155329 199822
rect 155539 199880 155605 199885
rect 155539 199824 155544 199880
rect 155600 199824 155605 199880
rect 155539 199819 155605 199824
rect 155542 199749 155602 199819
rect 155309 199746 155375 199749
rect 154990 199744 155375 199746
rect 154990 199688 155314 199744
rect 155370 199688 155375 199744
rect 154990 199686 155375 199688
rect 155309 199683 155375 199686
rect 155493 199744 155602 199749
rect 155493 199688 155498 199744
rect 155554 199688 155602 199744
rect 155493 199686 155602 199688
rect 155493 199683 155559 199686
rect 155953 199610 156019 199613
rect 156229 199610 156295 199613
rect 157014 199610 157074 199958
rect 157566 199919 157626 200094
rect 157195 199914 157261 199919
rect 157195 199858 157200 199914
rect 157256 199858 157261 199914
rect 157379 199914 157445 199919
rect 157379 199884 157384 199914
rect 157440 199884 157445 199914
rect 157563 199914 157629 199919
rect 157195 199853 157261 199858
rect 157198 199749 157258 199853
rect 157374 199820 157380 199884
rect 157444 199882 157450 199884
rect 157444 199822 157502 199882
rect 157563 199858 157568 199914
rect 157624 199858 157629 199914
rect 157563 199853 157629 199858
rect 158115 199914 158181 199919
rect 158115 199858 158120 199914
rect 158176 199858 158181 199914
rect 158115 199853 158181 199858
rect 158483 199914 158549 199919
rect 159311 199916 159377 199919
rect 158483 199858 158488 199914
rect 158544 199858 158549 199914
rect 159038 199914 159377 199916
rect 159038 199884 159316 199914
rect 158483 199853 158549 199858
rect 157444 199820 157450 199822
rect 158118 199749 158178 199853
rect 157149 199744 157258 199749
rect 157149 199688 157154 199744
rect 157210 199688 157258 199744
rect 157149 199686 157258 199688
rect 158069 199744 158178 199749
rect 158069 199688 158074 199744
rect 158130 199688 158178 199744
rect 158069 199686 158178 199688
rect 157149 199683 157215 199686
rect 158069 199683 158135 199686
rect 158486 199613 158546 199853
rect 159030 199820 159036 199884
rect 159100 199858 159316 199884
rect 159372 199858 159377 199914
rect 159100 199856 159377 199858
rect 159100 199820 159106 199856
rect 159311 199853 159377 199856
rect 159679 199916 159745 199919
rect 160599 199916 160665 199919
rect 159679 199914 159788 199916
rect 159679 199858 159684 199914
rect 159740 199858 159788 199914
rect 159679 199853 159788 199858
rect 160599 199914 160938 199916
rect 160599 199858 160604 199914
rect 160660 199858 160938 199914
rect 161427 199914 161493 199919
rect 160599 199856 160938 199858
rect 160599 199853 160665 199856
rect 158621 199744 158687 199749
rect 158621 199688 158626 199744
rect 158682 199688 158687 199744
rect 158621 199683 158687 199688
rect 158897 199746 158963 199749
rect 158897 199744 159098 199746
rect 158897 199688 158902 199744
rect 158958 199688 159098 199744
rect 158897 199686 159098 199688
rect 158897 199683 158963 199686
rect 158253 199610 158319 199613
rect 155953 199608 156154 199610
rect 155953 199552 155958 199608
rect 156014 199552 156154 199608
rect 155953 199550 156154 199552
rect 155953 199547 156019 199550
rect 153009 199472 153394 199474
rect 153009 199416 153014 199472
rect 153070 199416 153394 199472
rect 153009 199414 153394 199416
rect 153009 199411 153075 199414
rect 156094 199341 156154 199550
rect 156229 199608 156338 199610
rect 156229 199552 156234 199608
rect 156290 199552 156338 199608
rect 156229 199547 156338 199552
rect 157014 199608 158319 199610
rect 157014 199552 158258 199608
rect 158314 199552 158319 199608
rect 157014 199550 158319 199552
rect 158253 199547 158319 199550
rect 158437 199608 158546 199613
rect 158437 199552 158442 199608
rect 158498 199552 158546 199608
rect 158437 199550 158546 199552
rect 158624 199610 158684 199683
rect 158897 199610 158963 199613
rect 158624 199608 158963 199610
rect 158624 199552 158902 199608
rect 158958 199552 158963 199608
rect 158624 199550 158963 199552
rect 158437 199547 158503 199550
rect 158897 199547 158963 199550
rect 126329 199338 126395 199341
rect 153745 199338 153811 199341
rect 126329 199336 153811 199338
rect 126329 199280 126334 199336
rect 126390 199280 153750 199336
rect 153806 199280 153811 199336
rect 126329 199278 153811 199280
rect 156094 199336 156203 199341
rect 156094 199280 156142 199336
rect 156198 199280 156203 199336
rect 156094 199278 156203 199280
rect 126329 199275 126395 199278
rect 153745 199275 153811 199278
rect 156137 199275 156203 199278
rect 129181 199202 129247 199205
rect 139669 199202 139735 199205
rect 141141 199202 141207 199205
rect 141509 199204 141575 199205
rect 141693 199204 141759 199205
rect 142153 199204 142219 199205
rect 141509 199202 141556 199204
rect 129181 199200 138030 199202
rect 129181 199144 129186 199200
rect 129242 199144 138030 199200
rect 129181 199142 138030 199144
rect 129181 199139 129247 199142
rect 135156 199004 135162 199068
rect 135226 199066 135232 199068
rect 135713 199066 135779 199069
rect 135226 199064 135779 199066
rect 135226 199008 135718 199064
rect 135774 199008 135779 199064
rect 135226 199006 135779 199008
rect 135226 199004 135232 199006
rect 135713 199003 135779 199006
rect 137001 199066 137067 199069
rect 137134 199066 137140 199068
rect 137001 199064 137140 199066
rect 137001 199008 137006 199064
rect 137062 199008 137140 199064
rect 137001 199006 137140 199008
rect 137001 199003 137067 199006
rect 137134 199004 137140 199006
rect 137204 199004 137210 199068
rect 137970 199066 138030 199142
rect 139669 199200 141207 199202
rect 139669 199144 139674 199200
rect 139730 199144 141146 199200
rect 141202 199144 141207 199200
rect 139669 199142 141207 199144
rect 141464 199200 141556 199202
rect 141464 199144 141514 199200
rect 141464 199142 141556 199144
rect 139669 199139 139735 199142
rect 141141 199139 141207 199142
rect 141509 199140 141556 199142
rect 141620 199140 141626 199204
rect 141693 199200 141740 199204
rect 141804 199202 141810 199204
rect 141693 199144 141698 199200
rect 141693 199140 141740 199144
rect 141804 199142 141850 199202
rect 141804 199140 141810 199142
rect 142102 199140 142108 199204
rect 142172 199202 142219 199204
rect 142981 199202 143047 199205
rect 143206 199202 143212 199204
rect 142172 199200 142264 199202
rect 142214 199144 142264 199200
rect 142172 199142 142264 199144
rect 142981 199200 143212 199202
rect 142981 199144 142986 199200
rect 143042 199144 143212 199200
rect 142981 199142 143212 199144
rect 142172 199140 142219 199142
rect 141509 199139 141575 199140
rect 141693 199139 141759 199140
rect 142153 199139 142219 199140
rect 142981 199139 143047 199142
rect 143206 199140 143212 199142
rect 143276 199140 143282 199204
rect 155953 199202 156019 199205
rect 156278 199202 156338 199547
rect 156822 199412 156828 199476
rect 156892 199474 156898 199476
rect 159038 199474 159098 199686
rect 159728 199610 159788 199853
rect 160553 199746 160619 199749
rect 160510 199744 160619 199746
rect 160510 199688 160558 199744
rect 160614 199688 160619 199744
rect 160510 199683 160619 199688
rect 160510 199613 160570 199683
rect 159909 199610 159975 199613
rect 159728 199608 159975 199610
rect 159728 199552 159914 199608
rect 159970 199552 159975 199608
rect 159728 199550 159975 199552
rect 160510 199608 160619 199613
rect 160510 199552 160558 199608
rect 160614 199552 160619 199608
rect 160510 199550 160619 199552
rect 160878 199610 160938 199856
rect 161054 199820 161060 199884
rect 161124 199882 161130 199884
rect 161427 199882 161432 199914
rect 161124 199858 161432 199882
rect 161488 199858 161493 199914
rect 162163 199914 162229 199919
rect 162163 199884 162168 199914
rect 162224 199884 162229 199914
rect 162439 199916 162505 199919
rect 163543 199916 163609 199919
rect 162439 199914 162548 199916
rect 161124 199853 161493 199858
rect 161124 199822 161490 199853
rect 161124 199820 161130 199822
rect 162158 199820 162164 199884
rect 162228 199882 162234 199884
rect 162228 199822 162286 199882
rect 162439 199858 162444 199914
rect 162500 199884 162548 199914
rect 163270 199914 163609 199916
rect 162500 199858 162532 199884
rect 162439 199853 162532 199858
rect 162488 199822 162532 199853
rect 162228 199820 162234 199822
rect 162526 199820 162532 199822
rect 162596 199820 162602 199884
rect 163270 199858 163548 199914
rect 163604 199858 163609 199914
rect 164003 199914 164069 199919
rect 165751 199916 165817 199919
rect 163727 199882 163793 199885
rect 163270 199856 163609 199858
rect 163129 199748 163195 199749
rect 163078 199746 163084 199748
rect 163038 199686 163084 199746
rect 163148 199744 163195 199748
rect 163190 199688 163195 199744
rect 163078 199684 163084 199686
rect 163148 199684 163195 199688
rect 163270 199746 163330 199856
rect 163543 199853 163609 199856
rect 163684 199880 163793 199882
rect 163684 199824 163732 199880
rect 163788 199824 163793 199880
rect 164003 199858 164008 199914
rect 164064 199858 164069 199914
rect 165616 199914 165817 199916
rect 164187 199884 164253 199885
rect 164003 199853 164069 199858
rect 163684 199819 163793 199824
rect 163684 199749 163744 199819
rect 163497 199746 163563 199749
rect 163270 199744 163563 199746
rect 163270 199688 163502 199744
rect 163558 199688 163563 199744
rect 163270 199686 163563 199688
rect 163129 199683 163195 199684
rect 163497 199683 163563 199686
rect 163681 199744 163747 199749
rect 163681 199688 163686 199744
rect 163742 199688 163747 199744
rect 163681 199683 163747 199688
rect 164006 199613 164066 199853
rect 164182 199820 164188 199884
rect 164252 199882 164258 199884
rect 164252 199822 164344 199882
rect 164555 199880 164621 199885
rect 164555 199824 164560 199880
rect 164616 199824 164621 199880
rect 164252 199820 164258 199822
rect 164187 199819 164253 199820
rect 164555 199819 164621 199824
rect 165107 199880 165173 199885
rect 165616 199882 165756 199914
rect 165107 199824 165112 199880
rect 165168 199824 165173 199880
rect 165107 199819 165173 199824
rect 165340 199858 165756 199882
rect 165812 199858 165817 199914
rect 165340 199856 165817 199858
rect 165340 199822 165676 199856
rect 165751 199853 165817 199856
rect 164558 199749 164618 199819
rect 164509 199744 164618 199749
rect 164509 199688 164514 199744
rect 164570 199688 164618 199744
rect 164509 199686 164618 199688
rect 164509 199683 164575 199686
rect 163129 199610 163195 199613
rect 160878 199608 163195 199610
rect 160878 199552 163134 199608
rect 163190 199552 163195 199608
rect 160878 199550 163195 199552
rect 159909 199547 159975 199550
rect 160553 199547 160619 199550
rect 163129 199547 163195 199550
rect 163957 199608 164066 199613
rect 163957 199552 163962 199608
rect 164018 199552 164066 199608
rect 163957 199550 164066 199552
rect 163957 199547 164023 199550
rect 165110 199477 165170 199819
rect 165340 199749 165400 199822
rect 166076 199749 166136 200230
rect 200389 200227 200455 200230
rect 166398 200094 170000 200154
rect 166398 199919 166458 200094
rect 166395 199914 166461 199919
rect 166395 199858 166400 199914
rect 166456 199858 166461 199914
rect 166763 199914 166829 199919
rect 166763 199884 166768 199914
rect 166824 199884 166829 199914
rect 168235 199914 168301 199919
rect 169431 199916 169497 199919
rect 166395 199853 166461 199858
rect 166758 199820 166764 199884
rect 166828 199882 166834 199884
rect 167499 199882 167565 199885
rect 166828 199822 166886 199882
rect 167456 199880 167565 199882
rect 167456 199824 167504 199880
rect 167560 199824 167565 199880
rect 168235 199858 168240 199914
rect 168296 199858 168301 199914
rect 169296 199914 169497 199916
rect 168235 199853 168301 199858
rect 168971 199880 169037 199885
rect 166828 199820 166834 199822
rect 167456 199819 167565 199824
rect 167039 199780 167105 199783
rect 166996 199778 167105 199780
rect 165337 199744 165403 199749
rect 165337 199688 165342 199744
rect 165398 199688 165403 199744
rect 165337 199683 165403 199688
rect 166073 199744 166139 199749
rect 166073 199688 166078 199744
rect 166134 199688 166139 199744
rect 166073 199683 166139 199688
rect 166206 199684 166212 199748
rect 166276 199746 166282 199748
rect 166996 199746 167044 199778
rect 166276 199722 167044 199746
rect 167100 199722 167105 199778
rect 167456 199749 167516 199819
rect 168238 199749 168298 199853
rect 168971 199824 168976 199880
rect 169032 199824 169037 199880
rect 168971 199819 169037 199824
rect 169296 199858 169436 199914
rect 169492 199858 169497 199914
rect 169296 199856 169497 199858
rect 168974 199749 169034 199819
rect 166276 199717 167105 199722
rect 167453 199744 167519 199749
rect 166276 199686 167056 199717
rect 167453 199688 167458 199744
rect 167514 199688 167519 199744
rect 166276 199684 166282 199686
rect 167453 199683 167519 199688
rect 168189 199744 168298 199749
rect 168189 199688 168194 199744
rect 168250 199688 168298 199744
rect 168189 199686 168298 199688
rect 168925 199744 169034 199749
rect 168925 199688 168930 199744
rect 168986 199688 169034 199744
rect 168925 199686 169034 199688
rect 169296 199746 169356 199856
rect 169431 199853 169497 199856
rect 169615 199916 169681 199919
rect 169615 199914 169816 199916
rect 169615 199858 169620 199914
rect 169676 199858 169816 199914
rect 169615 199856 169816 199858
rect 169615 199853 169681 199856
rect 169569 199746 169635 199749
rect 169756 199748 169816 199856
rect 169296 199744 169635 199746
rect 169296 199688 169574 199744
rect 169630 199688 169635 199744
rect 169296 199686 169635 199688
rect 168189 199683 168255 199686
rect 168925 199683 168991 199686
rect 169569 199683 169635 199686
rect 169702 199684 169708 199748
rect 169772 199686 169816 199748
rect 169940 199746 170000 200094
rect 172278 200092 172284 200156
rect 172348 200154 172354 200156
rect 172348 200094 172622 200154
rect 172348 200092 172354 200094
rect 172562 199919 172622 200094
rect 172830 200092 172836 200156
rect 172900 200154 172906 200156
rect 177941 200154 178007 200157
rect 172900 200152 178007 200154
rect 172900 200096 177946 200152
rect 178002 200096 178007 200152
rect 172900 200094 178007 200096
rect 172900 200092 172906 200094
rect 177941 200091 178007 200094
rect 176694 200018 176700 200020
rect 175966 199958 176700 200018
rect 170075 199914 170141 199919
rect 170075 199858 170080 199914
rect 170136 199882 170141 199914
rect 170627 199914 170693 199919
rect 171271 199916 171337 199919
rect 171823 199916 171889 199919
rect 170438 199882 170444 199884
rect 170136 199858 170444 199882
rect 170075 199853 170444 199858
rect 170078 199822 170444 199853
rect 170438 199820 170444 199822
rect 170508 199820 170514 199884
rect 170627 199858 170632 199914
rect 170688 199882 170693 199914
rect 171136 199914 171337 199916
rect 170806 199882 170812 199884
rect 170688 199858 170812 199882
rect 170627 199853 170812 199858
rect 170630 199822 170812 199853
rect 170806 199820 170812 199822
rect 170876 199820 170882 199884
rect 171136 199858 171276 199914
rect 171332 199858 171337 199914
rect 171136 199856 171337 199858
rect 170121 199746 170187 199749
rect 169940 199744 170187 199746
rect 169940 199688 170126 199744
rect 170182 199688 170187 199744
rect 169940 199686 170187 199688
rect 171136 199746 171196 199856
rect 171271 199853 171337 199856
rect 171550 199914 171889 199916
rect 171550 199858 171828 199914
rect 171884 199858 171889 199914
rect 172375 199914 172441 199919
rect 171550 199856 171889 199858
rect 171136 199686 171426 199746
rect 169772 199684 169778 199686
rect 170121 199683 170187 199686
rect 171366 199613 171426 199686
rect 167913 199610 167979 199613
rect 171174 199610 171180 199612
rect 167913 199608 171180 199610
rect 167913 199552 167918 199608
rect 167974 199552 171180 199608
rect 167913 199550 171180 199552
rect 167913 199547 167979 199550
rect 171174 199548 171180 199550
rect 171244 199548 171250 199612
rect 171317 199608 171426 199613
rect 171317 199552 171322 199608
rect 171378 199552 171426 199608
rect 171317 199550 171426 199552
rect 171550 199610 171610 199856
rect 171823 199853 171889 199856
rect 172099 199880 172165 199885
rect 172099 199824 172104 199880
rect 172160 199824 172165 199880
rect 172375 199858 172380 199914
rect 172436 199858 172441 199914
rect 172375 199853 172441 199858
rect 172559 199914 172625 199919
rect 172559 199858 172564 199914
rect 172620 199858 172625 199914
rect 172559 199853 172625 199858
rect 172743 199916 172809 199919
rect 172743 199914 172852 199916
rect 172743 199858 172748 199914
rect 172804 199858 172852 199914
rect 172743 199853 172852 199858
rect 173111 199914 173177 199919
rect 173111 199858 173116 199914
rect 173172 199858 173177 199914
rect 174123 199914 174189 199919
rect 173111 199853 173177 199858
rect 173295 199882 173361 199885
rect 173755 199884 173821 199885
rect 174123 199884 174128 199914
rect 174184 199884 174189 199914
rect 174307 199914 174373 199919
rect 173566 199882 173572 199884
rect 173295 199880 173572 199882
rect 172099 199819 172165 199824
rect 171869 199610 171935 199613
rect 171550 199608 171935 199610
rect 171550 199552 171874 199608
rect 171930 199552 171935 199608
rect 171550 199550 171935 199552
rect 172102 199610 172162 199819
rect 172378 199746 172438 199853
rect 172792 199749 172852 199853
rect 172646 199746 172652 199748
rect 172378 199686 172652 199746
rect 172646 199684 172652 199686
rect 172716 199684 172722 199748
rect 172789 199744 172855 199749
rect 172789 199688 172794 199744
rect 172850 199688 172855 199744
rect 172789 199683 172855 199688
rect 173114 199746 173174 199853
rect 173295 199824 173300 199880
rect 173356 199824 173572 199880
rect 173295 199822 173572 199824
rect 173295 199819 173361 199822
rect 173566 199820 173572 199822
rect 173636 199820 173642 199884
rect 173750 199820 173756 199884
rect 173820 199882 173826 199884
rect 173820 199822 173912 199882
rect 173820 199820 173826 199822
rect 174118 199820 174124 199884
rect 174188 199882 174194 199884
rect 174188 199822 174246 199882
rect 174307 199858 174312 199914
rect 174368 199858 174373 199914
rect 175135 199916 175201 199919
rect 175687 199916 175753 199919
rect 175135 199914 175244 199916
rect 174767 199882 174833 199885
rect 174307 199853 174373 199858
rect 174494 199880 174833 199882
rect 174188 199820 174194 199822
rect 173755 199819 173821 199820
rect 173382 199746 173388 199748
rect 173114 199686 173388 199746
rect 173382 199684 173388 199686
rect 173452 199684 173458 199748
rect 174310 199746 174370 199853
rect 174172 199686 174370 199746
rect 174494 199824 174772 199880
rect 174828 199824 174833 199880
rect 174494 199822 174833 199824
rect 174494 199746 174554 199822
rect 174767 199819 174833 199822
rect 174951 199882 175017 199885
rect 174951 199880 175060 199882
rect 174951 199824 174956 199880
rect 175012 199824 175060 199880
rect 175135 199858 175140 199914
rect 175196 199884 175244 199914
rect 175687 199914 175796 199916
rect 175196 199858 175228 199884
rect 175135 199853 175228 199858
rect 174951 199819 175060 199824
rect 175184 199822 175228 199853
rect 175222 199820 175228 199822
rect 175292 199820 175298 199884
rect 175687 199858 175692 199914
rect 175748 199882 175796 199914
rect 175966 199882 176026 199958
rect 176694 199956 176700 199958
rect 176764 199956 176770 200020
rect 175748 199858 176026 199882
rect 175687 199853 176026 199858
rect 175736 199822 176026 199853
rect 176142 199820 176148 199884
rect 176212 199882 176218 199884
rect 176423 199882 176489 199885
rect 177481 199884 177547 199885
rect 176212 199880 176489 199882
rect 176212 199824 176428 199880
rect 176484 199824 176489 199880
rect 176212 199822 176489 199824
rect 176212 199820 176218 199822
rect 176423 199819 176489 199822
rect 177430 199820 177436 199884
rect 177500 199882 177547 199884
rect 177500 199880 177592 199882
rect 177542 199824 177592 199880
rect 177500 199822 177592 199824
rect 177500 199820 177547 199822
rect 177481 199819 177547 199820
rect 174721 199746 174787 199749
rect 174494 199744 174787 199746
rect 174494 199688 174726 199744
rect 174782 199688 174787 199744
rect 174494 199686 174787 199688
rect 175000 199748 175060 199819
rect 175000 199686 175044 199748
rect 172421 199610 172487 199613
rect 172102 199608 172487 199610
rect 172102 199552 172426 199608
rect 172482 199552 172487 199608
rect 172102 199550 172487 199552
rect 171317 199547 171383 199550
rect 171869 199547 171935 199550
rect 172421 199547 172487 199550
rect 173566 199548 173572 199612
rect 173636 199610 173642 199612
rect 173801 199610 173867 199613
rect 173636 199608 173867 199610
rect 173636 199552 173806 199608
rect 173862 199552 173867 199608
rect 173636 199550 173867 199552
rect 173636 199548 173642 199550
rect 173801 199547 173867 199550
rect 156892 199414 159098 199474
rect 165061 199472 165170 199477
rect 165061 199416 165066 199472
rect 165122 199416 165170 199472
rect 165061 199414 165170 199416
rect 174172 199474 174232 199686
rect 174721 199683 174787 199686
rect 175038 199684 175044 199686
rect 175108 199684 175114 199748
rect 174353 199610 174419 199613
rect 174353 199608 186330 199610
rect 174353 199552 174358 199608
rect 174414 199552 186330 199608
rect 174353 199550 186330 199552
rect 174353 199547 174419 199550
rect 174353 199474 174419 199477
rect 174172 199472 174419 199474
rect 174172 199416 174358 199472
rect 174414 199416 174419 199472
rect 174172 199414 174419 199416
rect 156892 199412 156898 199414
rect 165061 199411 165127 199414
rect 174353 199411 174419 199414
rect 174629 199474 174695 199477
rect 174629 199472 184950 199474
rect 174629 199416 174634 199472
rect 174690 199416 184950 199472
rect 174629 199414 184950 199416
rect 174629 199411 174695 199414
rect 156781 199338 156847 199341
rect 177389 199338 177455 199341
rect 156781 199336 177455 199338
rect 156781 199280 156786 199336
rect 156842 199280 177394 199336
rect 177450 199280 177455 199336
rect 156781 199278 177455 199280
rect 156781 199275 156847 199278
rect 177389 199275 177455 199278
rect 155953 199200 156338 199202
rect 155953 199144 155958 199200
rect 156014 199144 156338 199200
rect 155953 199142 156338 199144
rect 160093 199202 160159 199205
rect 178585 199202 178651 199205
rect 160093 199200 178651 199202
rect 160093 199144 160098 199200
rect 160154 199144 178590 199200
rect 178646 199144 178651 199200
rect 160093 199142 178651 199144
rect 184890 199202 184950 199414
rect 186270 199338 186330 199550
rect 200798 199338 200804 199340
rect 186270 199278 200804 199338
rect 200798 199276 200804 199278
rect 200868 199276 200874 199340
rect 198958 199202 198964 199204
rect 184890 199142 198964 199202
rect 155953 199139 156019 199142
rect 160093 199139 160159 199142
rect 178585 199139 178651 199142
rect 198958 199140 198964 199142
rect 199028 199140 199034 199204
rect 151854 199066 151860 199068
rect 137970 199006 151860 199066
rect 151854 199004 151860 199006
rect 151924 199004 151930 199068
rect 158253 199066 158319 199069
rect 169293 199066 169359 199069
rect 158253 199064 169359 199066
rect 158253 199008 158258 199064
rect 158314 199008 169298 199064
rect 169354 199008 169359 199064
rect 158253 199006 169359 199008
rect 158253 199003 158319 199006
rect 169293 199003 169359 199006
rect 173525 199066 173591 199069
rect 173750 199066 173756 199068
rect 173525 199064 173756 199066
rect 173525 199008 173530 199064
rect 173586 199008 173756 199064
rect 173525 199006 173756 199008
rect 173525 199003 173591 199006
rect 173750 199004 173756 199006
rect 173820 199004 173826 199068
rect 175825 199066 175891 199069
rect 200614 199066 200620 199068
rect 175825 199064 200620 199066
rect 175825 199008 175830 199064
rect 175886 199008 200620 199064
rect 175825 199006 200620 199008
rect 175825 199003 175891 199006
rect 200614 199004 200620 199006
rect 200684 199004 200690 199068
rect 121269 198930 121335 198933
rect 152825 198930 152891 198933
rect 121269 198928 152891 198930
rect 121269 198872 121274 198928
rect 121330 198872 152830 198928
rect 152886 198872 152891 198928
rect 121269 198870 152891 198872
rect 121269 198867 121335 198870
rect 152825 198867 152891 198870
rect 170213 198930 170279 198933
rect 174353 198930 174419 198933
rect 170213 198928 174419 198930
rect 170213 198872 170218 198928
rect 170274 198872 174358 198928
rect 174414 198872 174419 198928
rect 170213 198870 174419 198872
rect 170213 198867 170279 198870
rect 174353 198867 174419 198870
rect 174537 198930 174603 198933
rect 174905 198930 174971 198933
rect 174537 198928 174971 198930
rect 174537 198872 174542 198928
rect 174598 198872 174910 198928
rect 174966 198872 174971 198928
rect 174537 198870 174971 198872
rect 174537 198867 174603 198870
rect 174905 198867 174971 198870
rect 176142 198868 176148 198932
rect 176212 198930 176218 198932
rect 176377 198930 176443 198933
rect 201534 198930 201540 198932
rect 176212 198928 176443 198930
rect 176212 198872 176382 198928
rect 176438 198872 176443 198928
rect 176212 198870 176443 198872
rect 176212 198868 176218 198870
rect 176377 198867 176443 198870
rect 176886 198870 201540 198930
rect 122966 198732 122972 198796
rect 123036 198794 123042 198796
rect 125041 198794 125107 198797
rect 155861 198794 155927 198797
rect 123036 198792 125107 198794
rect 123036 198736 125046 198792
rect 125102 198736 125107 198792
rect 123036 198734 125107 198736
rect 123036 198732 123042 198734
rect 125041 198731 125107 198734
rect 132358 198792 155927 198794
rect 132358 198736 155866 198792
rect 155922 198736 155927 198792
rect 132358 198734 155927 198736
rect 132358 198661 132418 198734
rect 155861 198731 155927 198734
rect 158621 198794 158687 198797
rect 172513 198794 172579 198797
rect 173617 198794 173683 198797
rect 158621 198792 171242 198794
rect 158621 198736 158626 198792
rect 158682 198736 171242 198792
rect 158621 198734 171242 198736
rect 158621 198731 158687 198734
rect 132309 198656 132418 198661
rect 132309 198600 132314 198656
rect 132370 198600 132418 198656
rect 132309 198598 132418 198600
rect 141877 198658 141943 198661
rect 143574 198658 143580 198660
rect 141877 198656 143580 198658
rect 141877 198600 141882 198656
rect 141938 198600 143580 198656
rect 141877 198598 143580 198600
rect 132309 198595 132375 198598
rect 141877 198595 141943 198598
rect 143574 198596 143580 198598
rect 143644 198596 143650 198660
rect 144310 198596 144316 198660
rect 144380 198658 144386 198660
rect 146661 198658 146727 198661
rect 144380 198656 146727 198658
rect 144380 198600 146666 198656
rect 146722 198600 146727 198656
rect 144380 198598 146727 198600
rect 144380 198596 144386 198598
rect 146661 198595 146727 198598
rect 148225 198658 148291 198661
rect 170949 198660 171015 198661
rect 148726 198658 148732 198660
rect 148225 198656 148732 198658
rect 148225 198600 148230 198656
rect 148286 198600 148732 198656
rect 148225 198598 148732 198600
rect 148225 198595 148291 198598
rect 148726 198596 148732 198598
rect 148796 198596 148802 198660
rect 170949 198656 170996 198660
rect 171060 198658 171066 198660
rect 171182 198658 171242 198734
rect 172513 198792 173683 198794
rect 172513 198736 172518 198792
rect 172574 198736 173622 198792
rect 173678 198736 173683 198792
rect 172513 198734 173683 198736
rect 172513 198731 172579 198734
rect 173617 198731 173683 198734
rect 174118 198732 174124 198796
rect 174188 198794 174194 198796
rect 175641 198794 175707 198797
rect 174188 198792 175707 198794
rect 174188 198736 175646 198792
rect 175702 198736 175707 198792
rect 174188 198734 175707 198736
rect 174188 198732 174194 198734
rect 175641 198731 175707 198734
rect 175917 198794 175983 198797
rect 176886 198794 176946 198870
rect 201534 198868 201540 198870
rect 201604 198868 201610 198932
rect 175917 198792 176946 198794
rect 175917 198736 175922 198792
rect 175978 198736 176946 198792
rect 175917 198734 176946 198736
rect 175917 198731 175983 198734
rect 177062 198732 177068 198796
rect 177132 198794 177138 198796
rect 177205 198794 177271 198797
rect 177132 198792 177271 198794
rect 177132 198736 177210 198792
rect 177266 198736 177271 198792
rect 177132 198734 177271 198736
rect 177132 198732 177138 198734
rect 177205 198731 177271 198734
rect 177389 198796 177455 198797
rect 177389 198792 177436 198796
rect 177500 198794 177506 198796
rect 177389 198736 177394 198792
rect 177389 198732 177436 198736
rect 177500 198734 177546 198794
rect 177500 198732 177506 198734
rect 177389 198731 177455 198732
rect 177941 198658 178007 198661
rect 170949 198600 170954 198656
rect 170949 198596 170996 198600
rect 171060 198598 171106 198658
rect 171182 198656 178007 198658
rect 171182 198600 177946 198656
rect 178002 198600 178007 198656
rect 171182 198598 178007 198600
rect 171060 198596 171066 198598
rect 170949 198595 171015 198596
rect 177941 198595 178007 198598
rect 178217 198658 178283 198661
rect 196014 198658 196020 198660
rect 178217 198656 196020 198658
rect 178217 198600 178222 198656
rect 178278 198600 196020 198656
rect 178217 198598 196020 198600
rect 178217 198595 178283 198598
rect 196014 198596 196020 198598
rect 196084 198596 196090 198660
rect 127617 198522 127683 198525
rect 135110 198522 135116 198524
rect 127617 198520 135116 198522
rect 127617 198464 127622 198520
rect 127678 198464 135116 198520
rect 127617 198462 135116 198464
rect 127617 198459 127683 198462
rect 135110 198460 135116 198462
rect 135180 198460 135186 198524
rect 142521 198522 142587 198525
rect 142654 198522 142660 198524
rect 142521 198520 142660 198522
rect 142521 198464 142526 198520
rect 142582 198464 142660 198520
rect 142521 198462 142660 198464
rect 142521 198459 142587 198462
rect 142654 198460 142660 198462
rect 142724 198460 142730 198524
rect 142797 198522 142863 198525
rect 143349 198524 143415 198525
rect 143022 198522 143028 198524
rect 142797 198520 143028 198522
rect 142797 198464 142802 198520
rect 142858 198464 143028 198520
rect 142797 198462 143028 198464
rect 142797 198459 142863 198462
rect 143022 198460 143028 198462
rect 143092 198460 143098 198524
rect 143349 198520 143396 198524
rect 143460 198522 143466 198524
rect 143901 198522 143967 198525
rect 146150 198522 146156 198524
rect 143349 198464 143354 198520
rect 143349 198460 143396 198464
rect 143460 198462 143506 198522
rect 143901 198520 146156 198522
rect 143901 198464 143906 198520
rect 143962 198464 146156 198520
rect 143901 198462 146156 198464
rect 143460 198460 143466 198462
rect 143349 198459 143415 198460
rect 143901 198459 143967 198462
rect 146150 198460 146156 198462
rect 146220 198460 146226 198524
rect 165470 198460 165476 198524
rect 165540 198522 165546 198524
rect 165797 198522 165863 198525
rect 165540 198520 165863 198522
rect 165540 198464 165802 198520
rect 165858 198464 165863 198520
rect 165540 198462 165863 198464
rect 165540 198460 165546 198462
rect 165797 198459 165863 198462
rect 170765 198522 170831 198525
rect 193254 198522 193260 198524
rect 170765 198520 193260 198522
rect 170765 198464 170770 198520
rect 170826 198464 193260 198520
rect 170765 198462 193260 198464
rect 170765 198459 170831 198462
rect 193254 198460 193260 198462
rect 193324 198460 193330 198524
rect 107510 198324 107516 198388
rect 107580 198386 107586 198388
rect 130653 198386 130719 198389
rect 107580 198384 130719 198386
rect 107580 198328 130658 198384
rect 130714 198328 130719 198384
rect 107580 198326 130719 198328
rect 107580 198324 107586 198326
rect 130653 198323 130719 198326
rect 136817 198386 136883 198389
rect 148041 198386 148107 198389
rect 136817 198384 148107 198386
rect 136817 198328 136822 198384
rect 136878 198328 148046 198384
rect 148102 198328 148107 198384
rect 136817 198326 148107 198328
rect 136817 198323 136883 198326
rect 148041 198323 148107 198326
rect 148910 198324 148916 198388
rect 148980 198386 148986 198388
rect 157609 198386 157675 198389
rect 148980 198384 157675 198386
rect 148980 198328 157614 198384
rect 157670 198328 157675 198384
rect 148980 198326 157675 198328
rect 148980 198324 148986 198326
rect 157609 198323 157675 198326
rect 158478 198324 158484 198388
rect 158548 198386 158554 198388
rect 171133 198386 171199 198389
rect 158548 198384 171199 198386
rect 158548 198328 171138 198384
rect 171194 198328 171199 198384
rect 158548 198326 171199 198328
rect 158548 198324 158554 198326
rect 171133 198323 171199 198326
rect 173566 198324 173572 198388
rect 173636 198386 173642 198388
rect 175273 198386 175339 198389
rect 197302 198386 197308 198388
rect 173636 198326 175106 198386
rect 173636 198324 173642 198326
rect 107326 198188 107332 198252
rect 107396 198250 107402 198252
rect 132585 198250 132651 198253
rect 107396 198248 132651 198250
rect 107396 198192 132590 198248
rect 132646 198192 132651 198248
rect 107396 198190 132651 198192
rect 107396 198188 107402 198190
rect 132585 198187 132651 198190
rect 146886 198188 146892 198252
rect 146956 198250 146962 198252
rect 150341 198250 150407 198253
rect 157333 198252 157399 198253
rect 162301 198252 162367 198253
rect 170489 198252 170555 198253
rect 157333 198250 157380 198252
rect 146956 198248 150407 198250
rect 146956 198192 150346 198248
rect 150402 198192 150407 198248
rect 146956 198190 150407 198192
rect 157288 198248 157380 198250
rect 157288 198192 157338 198248
rect 157288 198190 157380 198192
rect 146956 198188 146962 198190
rect 150341 198187 150407 198190
rect 157333 198188 157380 198190
rect 157444 198188 157450 198252
rect 162301 198248 162348 198252
rect 162412 198250 162418 198252
rect 170438 198250 170444 198252
rect 162301 198192 162306 198248
rect 162301 198188 162348 198192
rect 162412 198190 162458 198250
rect 170398 198190 170444 198250
rect 170508 198248 170555 198252
rect 170550 198192 170555 198248
rect 162412 198188 162418 198190
rect 170438 198188 170444 198190
rect 170508 198188 170555 198192
rect 157333 198187 157399 198188
rect 162301 198187 162367 198188
rect 170489 198187 170555 198188
rect 170949 198250 171015 198253
rect 175046 198250 175106 198326
rect 175273 198384 197308 198386
rect 175273 198328 175278 198384
rect 175334 198328 197308 198384
rect 175273 198326 197308 198328
rect 175273 198323 175339 198326
rect 197302 198324 197308 198326
rect 197372 198324 197378 198388
rect 199142 198250 199148 198252
rect 170949 198248 174600 198250
rect 170949 198192 170954 198248
rect 171010 198192 174600 198248
rect 170949 198190 174600 198192
rect 175046 198190 199148 198250
rect 170949 198187 171015 198190
rect 105629 198114 105695 198117
rect 126053 198114 126119 198117
rect 105629 198112 126119 198114
rect 105629 198056 105634 198112
rect 105690 198056 126058 198112
rect 126114 198056 126119 198112
rect 105629 198054 126119 198056
rect 105629 198051 105695 198054
rect 126053 198051 126119 198054
rect 136766 198052 136772 198116
rect 136836 198114 136842 198116
rect 137093 198114 137159 198117
rect 136836 198112 137159 198114
rect 136836 198056 137098 198112
rect 137154 198056 137159 198112
rect 136836 198054 137159 198056
rect 136836 198052 136842 198054
rect 137093 198051 137159 198054
rect 138289 198114 138355 198117
rect 149605 198116 149671 198117
rect 138790 198114 138796 198116
rect 138289 198112 138796 198114
rect 138289 198056 138294 198112
rect 138350 198056 138796 198112
rect 138289 198054 138796 198056
rect 138289 198051 138355 198054
rect 138790 198052 138796 198054
rect 138860 198052 138866 198116
rect 149605 198112 149652 198116
rect 149716 198114 149722 198116
rect 149605 198056 149610 198112
rect 149605 198052 149652 198056
rect 149716 198054 149762 198114
rect 149716 198052 149722 198054
rect 149830 198052 149836 198116
rect 149900 198114 149906 198116
rect 150249 198114 150315 198117
rect 149900 198112 150315 198114
rect 149900 198056 150254 198112
rect 150310 198056 150315 198112
rect 149900 198054 150315 198056
rect 149900 198052 149906 198054
rect 149605 198051 149671 198052
rect 150249 198051 150315 198054
rect 152273 198114 152339 198117
rect 152958 198114 152964 198116
rect 152273 198112 152964 198114
rect 152273 198056 152278 198112
rect 152334 198056 152964 198112
rect 152273 198054 152964 198056
rect 152273 198051 152339 198054
rect 152958 198052 152964 198054
rect 153028 198052 153034 198116
rect 154205 198114 154271 198117
rect 154430 198114 154436 198116
rect 154205 198112 154436 198114
rect 154205 198056 154210 198112
rect 154266 198056 154436 198112
rect 154205 198054 154436 198056
rect 154205 198051 154271 198054
rect 154430 198052 154436 198054
rect 154500 198052 154506 198116
rect 156413 198114 156479 198117
rect 157241 198116 157307 198117
rect 156638 198114 156644 198116
rect 156413 198112 156644 198114
rect 156413 198056 156418 198112
rect 156474 198056 156644 198112
rect 156413 198054 156644 198056
rect 156413 198051 156479 198054
rect 156638 198052 156644 198054
rect 156708 198052 156714 198116
rect 157190 198114 157196 198116
rect 157150 198054 157196 198114
rect 157260 198112 157307 198116
rect 166717 198116 166783 198117
rect 166717 198114 166764 198116
rect 157302 198056 157307 198112
rect 157190 198052 157196 198054
rect 157260 198052 157307 198056
rect 166672 198112 166764 198114
rect 166672 198056 166722 198112
rect 166672 198054 166764 198056
rect 157241 198051 157307 198052
rect 166717 198052 166764 198054
rect 166828 198052 166834 198116
rect 174540 198114 174600 198190
rect 199142 198188 199148 198190
rect 199212 198188 199218 198252
rect 196198 198114 196204 198116
rect 174540 198054 196204 198114
rect 196198 198052 196204 198054
rect 196268 198052 196274 198116
rect 166717 198051 166783 198052
rect 101765 197978 101831 197981
rect 133638 197978 133644 197980
rect 101765 197976 133644 197978
rect 101765 197920 101770 197976
rect 101826 197920 133644 197976
rect 101765 197918 133644 197920
rect 101765 197915 101831 197918
rect 133638 197916 133644 197918
rect 133708 197916 133714 197980
rect 146201 197978 146267 197981
rect 166206 197978 166212 197980
rect 146201 197976 166212 197978
rect 146201 197920 146206 197976
rect 146262 197920 166212 197976
rect 146201 197918 166212 197920
rect 146201 197915 146267 197918
rect 166206 197916 166212 197918
rect 166276 197916 166282 197980
rect 169661 197978 169727 197981
rect 211797 197978 211863 197981
rect 169661 197976 211863 197978
rect 169661 197920 169666 197976
rect 169722 197920 211802 197976
rect 211858 197920 211863 197976
rect 169661 197918 211863 197920
rect 169661 197915 169727 197918
rect 211797 197915 211863 197918
rect 156137 197842 156203 197845
rect 149102 197840 156203 197842
rect 149102 197784 156142 197840
rect 156198 197784 156203 197840
rect 149102 197782 156203 197784
rect 135161 197706 135227 197709
rect 135294 197706 135300 197708
rect 135161 197704 135300 197706
rect 135161 197648 135166 197704
rect 135222 197648 135300 197704
rect 135161 197646 135300 197648
rect 135161 197643 135227 197646
rect 135294 197644 135300 197646
rect 135364 197644 135370 197708
rect 147254 197644 147260 197708
rect 147324 197706 147330 197708
rect 149102 197706 149162 197782
rect 156137 197779 156203 197782
rect 162393 197842 162459 197845
rect 162526 197842 162532 197844
rect 162393 197840 162532 197842
rect 162393 197784 162398 197840
rect 162454 197784 162532 197840
rect 162393 197782 162532 197784
rect 162393 197779 162459 197782
rect 162526 197780 162532 197782
rect 162596 197780 162602 197844
rect 164969 197842 165035 197845
rect 169293 197842 169359 197845
rect 164969 197840 169359 197842
rect 164969 197784 164974 197840
rect 165030 197784 169298 197840
rect 169354 197784 169359 197840
rect 164969 197782 169359 197784
rect 164969 197779 165035 197782
rect 169293 197779 169359 197782
rect 172421 197842 172487 197845
rect 172830 197842 172836 197844
rect 172421 197840 172836 197842
rect 172421 197784 172426 197840
rect 172482 197784 172836 197840
rect 172421 197782 172836 197784
rect 172421 197779 172487 197782
rect 172830 197780 172836 197782
rect 172900 197780 172906 197844
rect 173617 197842 173683 197845
rect 191966 197842 191972 197844
rect 173617 197840 191972 197842
rect 173617 197784 173622 197840
rect 173678 197784 191972 197840
rect 173617 197782 191972 197784
rect 173617 197779 173683 197782
rect 191966 197780 191972 197782
rect 192036 197780 192042 197844
rect 147324 197646 149162 197706
rect 147324 197644 147330 197646
rect 124765 197570 124831 197573
rect 135478 197570 135484 197572
rect 124765 197568 135484 197570
rect 124765 197512 124770 197568
rect 124826 197512 135484 197568
rect 124765 197510 135484 197512
rect 124765 197507 124831 197510
rect 135478 197508 135484 197510
rect 135548 197508 135554 197572
rect 140865 197570 140931 197573
rect 142102 197570 142108 197572
rect 140865 197568 142108 197570
rect 140865 197512 140870 197568
rect 140926 197512 142108 197568
rect 140865 197510 142108 197512
rect 140865 197507 140931 197510
rect 142102 197508 142108 197510
rect 142172 197508 142178 197572
rect 147070 197508 147076 197572
rect 147140 197570 147146 197572
rect 149513 197570 149579 197573
rect 147140 197568 149579 197570
rect 147140 197512 149518 197568
rect 149574 197512 149579 197568
rect 147140 197510 149579 197512
rect 147140 197508 147146 197510
rect 149513 197507 149579 197510
rect 134006 197372 134012 197436
rect 134076 197434 134082 197436
rect 134425 197434 134491 197437
rect 134076 197432 134491 197434
rect 134076 197376 134430 197432
rect 134486 197376 134491 197432
rect 134076 197374 134491 197376
rect 134076 197372 134082 197374
rect 134425 197371 134491 197374
rect 143942 197372 143948 197436
rect 144012 197434 144018 197436
rect 144637 197434 144703 197437
rect 144012 197432 144703 197434
rect 144012 197376 144642 197432
rect 144698 197376 144703 197432
rect 144012 197374 144703 197376
rect 144012 197372 144018 197374
rect 144637 197371 144703 197374
rect 166993 197434 167059 197437
rect 172513 197434 172579 197437
rect 166993 197432 172579 197434
rect 166993 197376 166998 197432
rect 167054 197376 172518 197432
rect 172574 197376 172579 197432
rect 166993 197374 172579 197376
rect 166993 197371 167059 197374
rect 172513 197371 172579 197374
rect 124949 197298 125015 197301
rect 150157 197298 150223 197301
rect 124949 197296 150223 197298
rect 124949 197240 124954 197296
rect 125010 197240 150162 197296
rect 150218 197240 150223 197296
rect 124949 197238 150223 197240
rect 124949 197235 125015 197238
rect 150157 197235 150223 197238
rect 165245 197298 165311 197301
rect 198774 197298 198780 197300
rect 165245 197296 198780 197298
rect 165245 197240 165250 197296
rect 165306 197240 198780 197296
rect 165245 197238 198780 197240
rect 165245 197235 165311 197238
rect 198774 197236 198780 197238
rect 198844 197236 198850 197300
rect 118509 197162 118575 197165
rect 147438 197162 147444 197164
rect 118509 197160 147444 197162
rect 118509 197104 118514 197160
rect 118570 197104 147444 197160
rect 118509 197102 147444 197104
rect 118509 197099 118575 197102
rect 147438 197100 147444 197102
rect 147508 197100 147514 197164
rect 164182 197100 164188 197164
rect 164252 197162 164258 197164
rect 197353 197162 197419 197165
rect 164252 197160 197419 197162
rect 164252 197104 197358 197160
rect 197414 197104 197419 197160
rect 164252 197102 197419 197104
rect 164252 197100 164258 197102
rect 197353 197099 197419 197102
rect 105537 197026 105603 197029
rect 136541 197026 136607 197029
rect 105537 197024 136607 197026
rect 105537 196968 105542 197024
rect 105598 196968 136546 197024
rect 136602 196968 136607 197024
rect 105537 196966 136607 196968
rect 105537 196963 105603 196966
rect 136541 196963 136607 196966
rect 147438 196964 147444 197028
rect 147508 197026 147514 197028
rect 148869 197026 148935 197029
rect 147508 197024 148935 197026
rect 147508 196968 148874 197024
rect 148930 196968 148935 197024
rect 147508 196966 148935 196968
rect 147508 196964 147514 196966
rect 148869 196963 148935 196966
rect 162209 197026 162275 197029
rect 196065 197026 196131 197029
rect 162209 197024 196131 197026
rect 162209 196968 162214 197024
rect 162270 196968 196070 197024
rect 196126 196968 196131 197024
rect 162209 196966 196131 196968
rect 162209 196963 162275 196966
rect 196065 196963 196131 196966
rect 108246 196828 108252 196892
rect 108316 196890 108322 196892
rect 138473 196890 138539 196893
rect 162209 196892 162275 196893
rect 108316 196888 138539 196890
rect 108316 196832 138478 196888
rect 138534 196832 138539 196888
rect 108316 196830 138539 196832
rect 108316 196828 108322 196830
rect 138473 196827 138539 196830
rect 162158 196828 162164 196892
rect 162228 196890 162275 196892
rect 162485 196890 162551 196893
rect 195973 196890 196039 196893
rect 162228 196888 162320 196890
rect 162270 196832 162320 196888
rect 162228 196830 162320 196832
rect 162485 196888 196039 196890
rect 162485 196832 162490 196888
rect 162546 196832 195978 196888
rect 196034 196832 196039 196888
rect 162485 196830 196039 196832
rect 162228 196828 162275 196830
rect 162209 196827 162275 196828
rect 162485 196827 162551 196830
rect 195973 196827 196039 196830
rect 101857 196754 101923 196757
rect 134057 196754 134123 196757
rect 101857 196752 134123 196754
rect 101857 196696 101862 196752
rect 101918 196696 134062 196752
rect 134118 196696 134123 196752
rect 101857 196694 134123 196696
rect 101857 196691 101923 196694
rect 134057 196691 134123 196694
rect 136582 196692 136588 196756
rect 136652 196754 136658 196756
rect 137277 196754 137343 196757
rect 136652 196752 137343 196754
rect 136652 196696 137282 196752
rect 137338 196696 137343 196752
rect 136652 196694 137343 196696
rect 136652 196692 136658 196694
rect 137277 196691 137343 196694
rect 139342 196692 139348 196756
rect 139412 196754 139418 196756
rect 139853 196754 139919 196757
rect 139412 196752 139919 196754
rect 139412 196696 139858 196752
rect 139914 196696 139919 196752
rect 139412 196694 139919 196696
rect 139412 196692 139418 196694
rect 139853 196691 139919 196694
rect 141509 196754 141575 196757
rect 143758 196754 143764 196756
rect 141509 196752 143764 196754
rect 141509 196696 141514 196752
rect 141570 196696 143764 196752
rect 141509 196694 143764 196696
rect 141509 196691 141575 196694
rect 143758 196692 143764 196694
rect 143828 196692 143834 196756
rect 166625 196754 166691 196757
rect 200205 196754 200271 196757
rect 166625 196752 200271 196754
rect 166625 196696 166630 196752
rect 166686 196696 200210 196752
rect 200266 196696 200271 196752
rect 166625 196694 200271 196696
rect 166625 196691 166691 196694
rect 200205 196691 200271 196694
rect 104341 196618 104407 196621
rect 137870 196618 137876 196620
rect 104341 196616 137876 196618
rect 104341 196560 104346 196616
rect 104402 196560 137876 196616
rect 104341 196558 137876 196560
rect 104341 196555 104407 196558
rect 137870 196556 137876 196558
rect 137940 196556 137946 196620
rect 164233 196618 164299 196621
rect 197537 196618 197603 196621
rect 164233 196616 197603 196618
rect 164233 196560 164238 196616
rect 164294 196560 197542 196616
rect 197598 196560 197603 196616
rect 164233 196558 197603 196560
rect 164233 196555 164299 196558
rect 197537 196555 197603 196558
rect 169661 196484 169727 196485
rect 169661 196482 169708 196484
rect 169616 196480 169708 196482
rect 169616 196424 169666 196480
rect 169616 196422 169708 196424
rect 169661 196420 169708 196422
rect 169772 196420 169778 196484
rect 170581 196482 170647 196485
rect 170806 196482 170812 196484
rect 170581 196480 170812 196482
rect 170581 196424 170586 196480
rect 170642 196424 170812 196480
rect 170581 196422 170812 196424
rect 169661 196419 169727 196420
rect 170581 196419 170647 196422
rect 170806 196420 170812 196422
rect 170876 196420 170882 196484
rect 172278 196420 172284 196484
rect 172348 196482 172354 196484
rect 173750 196482 173756 196484
rect 172348 196422 173756 196482
rect 172348 196420 172354 196422
rect 173750 196420 173756 196422
rect 173820 196420 173826 196484
rect 169385 196346 169451 196349
rect 169518 196346 169524 196348
rect 169385 196344 169524 196346
rect 169385 196288 169390 196344
rect 169446 196288 169524 196344
rect 169385 196286 169524 196288
rect 169385 196283 169451 196286
rect 169518 196284 169524 196286
rect 169588 196284 169594 196348
rect 134333 195938 134399 195941
rect 134742 195938 134748 195940
rect 134333 195936 134748 195938
rect 134333 195880 134338 195936
rect 134394 195880 134748 195936
rect 134333 195878 134748 195880
rect 134333 195875 134399 195878
rect 134742 195876 134748 195878
rect 134812 195876 134818 195940
rect 168741 195938 168807 195941
rect 169334 195938 169340 195940
rect 168741 195936 169340 195938
rect 168741 195880 168746 195936
rect 168802 195880 169340 195936
rect 168741 195878 169340 195880
rect 168741 195875 168807 195878
rect 169334 195876 169340 195878
rect 169404 195876 169410 195940
rect 176561 195938 176627 195941
rect 193806 195938 193812 195940
rect 176561 195936 193812 195938
rect 176561 195880 176566 195936
rect 176622 195880 193812 195936
rect 176561 195878 193812 195880
rect 176561 195875 176627 195878
rect 193806 195876 193812 195878
rect 193876 195876 193882 195940
rect 104525 195802 104591 195805
rect 138013 195802 138079 195805
rect 104525 195800 138079 195802
rect 104525 195744 104530 195800
rect 104586 195744 138018 195800
rect 138074 195744 138079 195800
rect 104525 195742 138079 195744
rect 104525 195739 104591 195742
rect 138013 195739 138079 195742
rect 157190 195740 157196 195804
rect 157260 195802 157266 195804
rect 180241 195802 180307 195805
rect 157260 195800 180307 195802
rect 157260 195744 180246 195800
rect 180302 195744 180307 195800
rect 157260 195742 180307 195744
rect 157260 195740 157266 195742
rect 180241 195739 180307 195742
rect 100334 195604 100340 195668
rect 100404 195666 100410 195668
rect 132677 195666 132743 195669
rect 100404 195664 132743 195666
rect 100404 195608 132682 195664
rect 132738 195608 132743 195664
rect 100404 195606 132743 195608
rect 100404 195604 100410 195606
rect 132677 195603 132743 195606
rect 150433 195666 150499 195669
rect 151169 195666 151235 195669
rect 150433 195664 151235 195666
rect 150433 195608 150438 195664
rect 150494 195608 151174 195664
rect 151230 195608 151235 195664
rect 150433 195606 151235 195608
rect 150433 195603 150499 195606
rect 151169 195603 151235 195606
rect 173382 195604 173388 195668
rect 173452 195666 173458 195668
rect 173801 195666 173867 195669
rect 173452 195664 173867 195666
rect 173452 195608 173806 195664
rect 173862 195608 173867 195664
rect 173452 195606 173867 195608
rect 173452 195604 173458 195606
rect 173801 195603 173867 195606
rect 175181 195666 175247 195669
rect 201718 195666 201724 195668
rect 175181 195664 201724 195666
rect 175181 195608 175186 195664
rect 175242 195608 201724 195664
rect 175181 195606 201724 195608
rect 175181 195603 175247 195606
rect 201718 195604 201724 195606
rect 201788 195604 201794 195668
rect 118366 195468 118372 195532
rect 118436 195530 118442 195532
rect 152917 195530 152983 195533
rect 118436 195528 152983 195530
rect 118436 195472 152922 195528
rect 152978 195472 152983 195528
rect 118436 195470 152983 195472
rect 118436 195468 118442 195470
rect 152917 195467 152983 195470
rect 156638 195468 156644 195532
rect 156708 195530 156714 195532
rect 190453 195530 190519 195533
rect 156708 195528 190519 195530
rect 156708 195472 190458 195528
rect 190514 195472 190519 195528
rect 156708 195470 190519 195472
rect 156708 195468 156714 195470
rect 190453 195467 190519 195470
rect 97717 195394 97783 195397
rect 150433 195394 150499 195397
rect 97717 195392 150499 195394
rect 97717 195336 97722 195392
rect 97778 195336 150438 195392
rect 150494 195336 150499 195392
rect 97717 195334 150499 195336
rect 97717 195331 97783 195334
rect 150433 195331 150499 195334
rect 161105 195394 161171 195397
rect 194777 195394 194843 195397
rect 161105 195392 194843 195394
rect 161105 195336 161110 195392
rect 161166 195336 194782 195392
rect 194838 195336 194843 195392
rect 161105 195334 194843 195336
rect 161105 195331 161171 195334
rect 194777 195331 194843 195334
rect 119838 195196 119844 195260
rect 119908 195258 119914 195260
rect 132033 195258 132099 195261
rect 119908 195256 132099 195258
rect 119908 195200 132038 195256
rect 132094 195200 132099 195256
rect 119908 195198 132099 195200
rect 119908 195196 119914 195198
rect 132033 195195 132099 195198
rect 133045 195258 133111 195261
rect 133822 195258 133828 195260
rect 133045 195256 133828 195258
rect 133045 195200 133050 195256
rect 133106 195200 133828 195256
rect 133045 195198 133828 195200
rect 133045 195195 133111 195198
rect 133822 195196 133828 195198
rect 133892 195196 133898 195260
rect 138105 195258 138171 195261
rect 138422 195258 138428 195260
rect 138105 195256 138428 195258
rect 138105 195200 138110 195256
rect 138166 195200 138428 195256
rect 138105 195198 138428 195200
rect 138105 195195 138171 195198
rect 138422 195196 138428 195198
rect 138492 195196 138498 195260
rect 158897 195258 158963 195261
rect 191782 195258 191788 195260
rect 158897 195256 191788 195258
rect 158897 195200 158902 195256
rect 158958 195200 191788 195256
rect 158897 195198 191788 195200
rect 158897 195195 158963 195198
rect 191782 195196 191788 195198
rect 191852 195196 191858 195260
rect 138054 195060 138060 195124
rect 138124 195122 138130 195124
rect 138841 195122 138907 195125
rect 138124 195120 138907 195122
rect 138124 195064 138846 195120
rect 138902 195064 138907 195120
rect 138124 195062 138907 195064
rect 138124 195060 138130 195062
rect 138841 195059 138907 195062
rect 177757 195122 177823 195125
rect 194542 195122 194548 195124
rect 177757 195120 194548 195122
rect 177757 195064 177762 195120
rect 177818 195064 194548 195120
rect 177757 195062 194548 195064
rect 177757 195059 177823 195062
rect 194542 195060 194548 195062
rect 194612 195060 194618 195124
rect 168833 194306 168899 194309
rect 203006 194306 203012 194308
rect 168833 194304 203012 194306
rect 168833 194248 168838 194304
rect 168894 194248 203012 194304
rect 168833 194246 203012 194248
rect 168833 194243 168899 194246
rect 203006 194244 203012 194246
rect 203076 194244 203082 194308
rect 173433 194170 173499 194173
rect 207013 194170 207079 194173
rect 173433 194168 207079 194170
rect 173433 194112 173438 194168
rect 173494 194112 207018 194168
rect 207074 194112 207079 194168
rect 173433 194110 207079 194112
rect 173433 194107 173499 194110
rect 207013 194107 207079 194110
rect 158897 194034 158963 194037
rect 159030 194034 159036 194036
rect 158897 194032 159036 194034
rect 158897 193976 158902 194032
rect 158958 193976 159036 194032
rect 158897 193974 159036 193976
rect 158897 193971 158963 193974
rect 159030 193972 159036 193974
rect 159100 193972 159106 194036
rect 176653 194034 176719 194037
rect 209814 194034 209820 194036
rect 176653 194032 209820 194034
rect 176653 193976 176658 194032
rect 176714 193976 209820 194032
rect 176653 193974 209820 193976
rect 176653 193971 176719 193974
rect 209814 193972 209820 193974
rect 209884 193972 209890 194036
rect 100518 193836 100524 193900
rect 100588 193898 100594 193900
rect 125133 193898 125199 193901
rect 100588 193896 125199 193898
rect 100588 193840 125138 193896
rect 125194 193840 125199 193896
rect 100588 193838 125199 193840
rect 100588 193836 100594 193838
rect 125133 193835 125199 193838
rect 151353 193898 151419 193901
rect 192661 193898 192727 193901
rect 151353 193896 192727 193898
rect 151353 193840 151358 193896
rect 151414 193840 192666 193896
rect 192722 193840 192727 193896
rect 151353 193838 192727 193840
rect 151353 193835 151419 193838
rect 192661 193835 192727 193838
rect 168097 193354 168163 193357
rect 168230 193354 168236 193356
rect 168097 193352 168236 193354
rect 168097 193296 168102 193352
rect 168158 193296 168236 193352
rect 168097 193294 168236 193296
rect 168097 193291 168163 193294
rect 168230 193292 168236 193294
rect 168300 193292 168306 193356
rect 170397 193218 170463 193221
rect 186998 193218 187004 193220
rect 170397 193216 187004 193218
rect 170397 193160 170402 193216
rect 170458 193160 187004 193216
rect 170397 193158 187004 193160
rect 170397 193155 170463 193158
rect 186998 193156 187004 193158
rect 187068 193156 187074 193220
rect 130469 193082 130535 193085
rect 147438 193082 147444 193084
rect 130469 193080 147444 193082
rect 130469 193024 130474 193080
rect 130530 193024 147444 193080
rect 130469 193022 147444 193024
rect 130469 193019 130535 193022
rect 147438 193020 147444 193022
rect 147508 193020 147514 193084
rect 172462 193020 172468 193084
rect 172532 193082 172538 193084
rect 205582 193082 205588 193084
rect 172532 193022 205588 193082
rect 172532 193020 172538 193022
rect 205582 193020 205588 193022
rect 205652 193020 205658 193084
rect 103278 192884 103284 192948
rect 103348 192946 103354 192948
rect 133597 192946 133663 192949
rect 103348 192944 133663 192946
rect 103348 192888 133602 192944
rect 133658 192888 133663 192944
rect 103348 192886 133663 192888
rect 103348 192884 103354 192886
rect 133597 192883 133663 192886
rect 133822 192884 133828 192948
rect 133892 192946 133898 192948
rect 134793 192946 134859 192949
rect 133892 192944 134859 192946
rect 133892 192888 134798 192944
rect 134854 192888 134859 192944
rect 133892 192886 134859 192888
rect 133892 192884 133898 192886
rect 134793 192883 134859 192886
rect 161054 192884 161060 192948
rect 161124 192946 161130 192948
rect 194685 192946 194751 192949
rect 161124 192944 194751 192946
rect 161124 192888 194690 192944
rect 194746 192888 194751 192944
rect 161124 192886 194751 192888
rect 161124 192884 161130 192886
rect 194685 192883 194751 192886
rect 104014 192748 104020 192812
rect 104084 192810 104090 192812
rect 125869 192810 125935 192813
rect 104084 192808 125935 192810
rect 104084 192752 125874 192808
rect 125930 192752 125935 192808
rect 104084 192750 125935 192752
rect 104084 192748 104090 192750
rect 125869 192747 125935 192750
rect 170438 192748 170444 192812
rect 170508 192810 170514 192812
rect 205173 192810 205239 192813
rect 170508 192808 205239 192810
rect 170508 192752 205178 192808
rect 205234 192752 205239 192808
rect 170508 192750 205239 192752
rect 170508 192748 170514 192750
rect 205173 192747 205239 192750
rect 113725 192674 113791 192677
rect 144310 192674 144316 192676
rect 113725 192672 144316 192674
rect 113725 192616 113730 192672
rect 113786 192616 144316 192672
rect 113725 192614 144316 192616
rect 113725 192611 113791 192614
rect 144310 192612 144316 192614
rect 144380 192612 144386 192676
rect 171777 192674 171843 192677
rect 205817 192674 205883 192677
rect 171777 192672 205883 192674
rect 171777 192616 171782 192672
rect 171838 192616 205822 192672
rect 205878 192616 205883 192672
rect 171777 192614 205883 192616
rect 171777 192611 171843 192614
rect 205817 192611 205883 192614
rect 124806 192476 124812 192540
rect 124876 192538 124882 192540
rect 156965 192538 157031 192541
rect 124876 192536 157031 192538
rect 124876 192480 156970 192536
rect 157026 192480 157031 192536
rect 124876 192478 157031 192480
rect 124876 192476 124882 192478
rect 156965 192475 157031 192478
rect 170990 192476 170996 192540
rect 171060 192538 171066 192540
rect 204805 192538 204871 192541
rect 171060 192536 204871 192538
rect 171060 192480 204810 192536
rect 204866 192480 204871 192536
rect 171060 192478 204871 192480
rect 171060 192476 171066 192478
rect 204805 192475 204871 192478
rect 580165 192538 580231 192541
rect 583520 192538 584960 192628
rect 580165 192536 584960 192538
rect 580165 192480 580170 192536
rect 580226 192480 584960 192536
rect 580165 192478 584960 192480
rect 580165 192475 580231 192478
rect 179413 192402 179479 192405
rect 187918 192402 187924 192404
rect 179413 192400 187924 192402
rect 179413 192344 179418 192400
rect 179474 192344 187924 192400
rect 179413 192342 187924 192344
rect 179413 192339 179479 192342
rect 187918 192340 187924 192342
rect 187988 192340 187994 192404
rect 583520 192388 584960 192478
rect 109534 191660 109540 191724
rect 109604 191722 109610 191724
rect 138790 191722 138796 191724
rect 109604 191662 138796 191722
rect 109604 191660 109610 191662
rect 138790 191660 138796 191662
rect 138860 191660 138866 191724
rect 100661 191586 100727 191589
rect 133822 191586 133828 191588
rect 100661 191584 133828 191586
rect 100661 191528 100666 191584
rect 100722 191528 133828 191584
rect 100661 191526 133828 191528
rect 100661 191523 100727 191526
rect 133822 191524 133828 191526
rect 133892 191524 133898 191588
rect 118550 191388 118556 191452
rect 118620 191450 118626 191452
rect 151813 191450 151879 191453
rect 118620 191448 151879 191450
rect 118620 191392 151818 191448
rect 151874 191392 151879 191448
rect 118620 191390 151879 191392
rect 118620 191388 118626 191390
rect 151813 191387 151879 191390
rect 102041 191314 102107 191317
rect 135478 191314 135484 191316
rect 102041 191312 135484 191314
rect 102041 191256 102046 191312
rect 102102 191256 135484 191312
rect 102041 191254 135484 191256
rect 102041 191251 102107 191254
rect 135478 191252 135484 191254
rect 135548 191252 135554 191316
rect 100569 191178 100635 191181
rect 134006 191178 134012 191180
rect 100569 191176 134012 191178
rect 100569 191120 100574 191176
rect 100630 191120 134012 191176
rect 100569 191118 134012 191120
rect 100569 191115 100635 191118
rect 134006 191116 134012 191118
rect 134076 191116 134082 191180
rect 101949 191042 102015 191045
rect 135294 191042 135300 191044
rect 101949 191040 135300 191042
rect 101949 190984 101954 191040
rect 102010 190984 135300 191040
rect 101949 190982 135300 190984
rect 101949 190979 102015 190982
rect 135294 190980 135300 190982
rect 135364 190980 135370 191044
rect 162301 191042 162367 191045
rect 186078 191042 186084 191044
rect 162301 191040 186084 191042
rect 162301 190984 162306 191040
rect 162362 190984 186084 191040
rect 162301 190982 186084 190984
rect 162301 190979 162367 190982
rect 186078 190980 186084 190982
rect 186148 190980 186154 191044
rect 106181 190226 106247 190229
rect 138422 190226 138428 190228
rect 106181 190224 138428 190226
rect 106181 190168 106186 190224
rect 106242 190168 138428 190224
rect 106181 190166 138428 190168
rect 106181 190163 106247 190166
rect 138422 190164 138428 190166
rect 138492 190164 138498 190228
rect 108481 190090 108547 190093
rect 142286 190090 142292 190092
rect 108481 190088 142292 190090
rect 108481 190032 108486 190088
rect 108542 190032 142292 190088
rect 108481 190030 142292 190032
rect 108481 190027 108547 190030
rect 142286 190028 142292 190030
rect 142356 190028 142362 190092
rect 160645 190090 160711 190093
rect 181294 190090 181300 190092
rect 160645 190088 181300 190090
rect 160645 190032 160650 190088
rect 160706 190032 181300 190088
rect 160645 190030 181300 190032
rect 160645 190027 160711 190030
rect 181294 190028 181300 190030
rect 181364 190028 181370 190092
rect 110045 189954 110111 189957
rect 143942 189954 143948 189956
rect 110045 189952 143948 189954
rect 110045 189896 110050 189952
rect 110106 189896 143948 189952
rect 110045 189894 143948 189896
rect 110045 189891 110111 189894
rect 143942 189892 143948 189894
rect 144012 189892 144018 189956
rect 176510 189892 176516 189956
rect 176580 189954 176586 189956
rect 209998 189954 210004 189956
rect 176580 189894 210004 189954
rect 176580 189892 176586 189894
rect 209998 189892 210004 189894
rect 210068 189892 210074 189956
rect 106825 189818 106891 189821
rect 142470 189818 142476 189820
rect 106825 189816 142476 189818
rect 106825 189760 106830 189816
rect 106886 189760 142476 189816
rect 106825 189758 142476 189760
rect 106825 189755 106891 189758
rect 142470 189756 142476 189758
rect 142540 189756 142546 189820
rect 174854 189756 174860 189820
rect 174924 189818 174930 189820
rect 208393 189818 208459 189821
rect 174924 189816 208459 189818
rect 174924 189760 208398 189816
rect 208454 189760 208459 189816
rect 174924 189758 208459 189760
rect 174924 189756 174930 189758
rect 208393 189755 208459 189758
rect 108205 189682 108271 189685
rect 143758 189682 143764 189684
rect 108205 189680 143764 189682
rect 108205 189624 108210 189680
rect 108266 189624 143764 189680
rect 108205 189622 143764 189624
rect 108205 189619 108271 189622
rect 143758 189620 143764 189622
rect 143828 189620 143834 189684
rect 154430 189620 154436 189684
rect 154500 189682 154506 189684
rect 218053 189682 218119 189685
rect 154500 189680 218119 189682
rect 154500 189624 218058 189680
rect 218114 189624 218119 189680
rect 154500 189622 218119 189624
rect 154500 189620 154506 189622
rect 218053 189619 218119 189622
rect -960 188866 480 188956
rect 3417 188866 3483 188869
rect -960 188864 3483 188866
rect -960 188808 3422 188864
rect 3478 188808 3483 188864
rect -960 188806 3483 188808
rect -960 188716 480 188806
rect 3417 188803 3483 188806
rect 115473 187642 115539 187645
rect 142102 187642 142108 187644
rect 115473 187640 142108 187642
rect 115473 187584 115478 187640
rect 115534 187584 142108 187640
rect 115473 187582 142108 187584
rect 115473 187579 115539 187582
rect 142102 187580 142108 187582
rect 142172 187580 142178 187644
rect 108430 187444 108436 187508
rect 108500 187506 108506 187508
rect 137277 187506 137343 187509
rect 108500 187504 137343 187506
rect 108500 187448 137282 187504
rect 137338 187448 137343 187504
rect 108500 187446 137343 187448
rect 108500 187444 108506 187446
rect 137277 187443 137343 187446
rect 107469 187370 107535 187373
rect 138238 187370 138244 187372
rect 107469 187368 138244 187370
rect 107469 187312 107474 187368
rect 107530 187312 138244 187368
rect 107469 187310 138244 187312
rect 107469 187307 107535 187310
rect 138238 187308 138244 187310
rect 138308 187308 138314 187372
rect 175038 187308 175044 187372
rect 175108 187370 175114 187372
rect 212625 187370 212691 187373
rect 175108 187368 212691 187370
rect 175108 187312 212630 187368
rect 212686 187312 212691 187368
rect 175108 187310 212691 187312
rect 175108 187308 175114 187310
rect 212625 187307 212691 187310
rect 106641 187234 106707 187237
rect 139526 187234 139532 187236
rect 106641 187232 139532 187234
rect 106641 187176 106646 187232
rect 106702 187176 139532 187232
rect 106641 187174 139532 187176
rect 106641 187171 106707 187174
rect 139526 187172 139532 187174
rect 139596 187172 139602 187236
rect 152958 187172 152964 187236
rect 153028 187234 153034 187236
rect 215293 187234 215359 187237
rect 153028 187232 215359 187234
rect 153028 187176 215298 187232
rect 215354 187176 215359 187232
rect 153028 187174 215359 187176
rect 153028 187172 153034 187174
rect 215293 187171 215359 187174
rect 104801 187098 104867 187101
rect 138054 187098 138060 187100
rect 104801 187096 138060 187098
rect 104801 187040 104806 187096
rect 104862 187040 138060 187096
rect 104801 187038 138060 187040
rect 104801 187035 104867 187038
rect 138054 187036 138060 187038
rect 138124 187036 138130 187100
rect 149830 187036 149836 187100
rect 149900 187098 149906 187100
rect 215753 187098 215819 187101
rect 149900 187096 215819 187098
rect 149900 187040 215758 187096
rect 215814 187040 215819 187096
rect 149900 187038 215819 187040
rect 149900 187036 149906 187038
rect 215753 187035 215819 187038
rect 99281 186962 99347 186965
rect 132534 186962 132540 186964
rect 99281 186960 132540 186962
rect 99281 186904 99286 186960
rect 99342 186904 132540 186960
rect 99281 186902 132540 186904
rect 99281 186899 99347 186902
rect 132534 186900 132540 186902
rect 132604 186900 132610 186964
rect 149646 186900 149652 186964
rect 149716 186962 149722 186964
rect 215569 186962 215635 186965
rect 149716 186960 215635 186962
rect 149716 186904 215574 186960
rect 215630 186904 215635 186960
rect 149716 186902 215635 186904
rect 149716 186900 149722 186902
rect 215569 186899 215635 186902
rect 580165 179210 580231 179213
rect 583520 179210 584960 179300
rect 580165 179208 584960 179210
rect 580165 179152 580170 179208
rect 580226 179152 584960 179208
rect 580165 179150 584960 179152
rect 580165 179147 580231 179150
rect 583520 179060 584960 179150
rect -960 175796 480 176036
rect 580165 165882 580231 165885
rect 583520 165882 584960 165972
rect 580165 165880 584960 165882
rect 580165 165824 580170 165880
rect 580226 165824 584960 165880
rect 580165 165822 584960 165824
rect 580165 165819 580231 165822
rect 583520 165732 584960 165822
rect -960 162890 480 162980
rect 3509 162890 3575 162893
rect -960 162888 3575 162890
rect -960 162832 3514 162888
rect 3570 162832 3575 162888
rect -960 162830 3575 162832
rect -960 162740 480 162830
rect 3509 162827 3575 162830
rect 148726 159292 148732 159356
rect 148796 159354 148802 159356
rect 210509 159354 210575 159357
rect 148796 159352 210575 159354
rect 148796 159296 210514 159352
rect 210570 159296 210575 159352
rect 148796 159294 210575 159296
rect 148796 159292 148802 159294
rect 210509 159291 210575 159294
rect 168230 156844 168236 156908
rect 168300 156906 168306 156908
rect 202413 156906 202479 156909
rect 168300 156904 202479 156906
rect 168300 156848 202418 156904
rect 202474 156848 202479 156904
rect 168300 156846 202479 156848
rect 168300 156844 168306 156846
rect 202413 156843 202479 156846
rect 169334 156708 169340 156772
rect 169404 156770 169410 156772
rect 203006 156770 203012 156772
rect 169404 156710 203012 156770
rect 169404 156708 169410 156710
rect 203006 156708 203012 156710
rect 203076 156708 203082 156772
rect 168741 156634 168807 156637
rect 203190 156634 203196 156636
rect 168741 156632 203196 156634
rect 168741 156576 168746 156632
rect 168802 156576 203196 156632
rect 168741 156574 203196 156576
rect 168741 156571 168807 156574
rect 203190 156572 203196 156574
rect 203260 156572 203266 156636
rect 177021 153914 177087 153917
rect 211286 153914 211292 153916
rect 177021 153912 211292 153914
rect 177021 153856 177026 153912
rect 177082 153856 211292 153912
rect 177021 153854 211292 153856
rect 177021 153851 177087 153854
rect 211286 153852 211292 153854
rect 211356 153852 211362 153916
rect 176837 153778 176903 153781
rect 211102 153778 211108 153780
rect 176837 153776 211108 153778
rect 176837 153720 176842 153776
rect 176898 153720 211108 153776
rect 176837 153718 211108 153720
rect 176837 153715 176903 153718
rect 211102 153716 211108 153718
rect 211172 153716 211178 153780
rect 579981 152690 580047 152693
rect 583520 152690 584960 152780
rect 579981 152688 584960 152690
rect 579981 152632 579986 152688
rect 580042 152632 584960 152688
rect 579981 152630 584960 152632
rect 579981 152627 580047 152630
rect 583520 152540 584960 152630
rect 177062 151404 177068 151468
rect 177132 151466 177138 151468
rect 207054 151466 207060 151468
rect 177132 151406 207060 151466
rect 177132 151404 177138 151406
rect 207054 151404 207060 151406
rect 207124 151404 207130 151468
rect 175457 151330 175523 151333
rect 205950 151330 205956 151332
rect 175457 151328 205956 151330
rect 175457 151272 175462 151328
rect 175518 151272 205956 151328
rect 175457 151270 205956 151272
rect 175457 151267 175523 151270
rect 205950 151268 205956 151270
rect 206020 151268 206026 151332
rect 122414 151132 122420 151196
rect 122484 151194 122490 151196
rect 139342 151194 139348 151196
rect 122484 151134 139348 151194
rect 122484 151132 122490 151134
rect 139342 151132 139348 151134
rect 139412 151132 139418 151196
rect 176653 151194 176719 151197
rect 207238 151194 207244 151196
rect 176653 151192 207244 151194
rect 176653 151136 176658 151192
rect 176714 151136 207244 151192
rect 176653 151134 207244 151136
rect 176653 151131 176719 151134
rect 207238 151132 207244 151134
rect 207308 151132 207314 151196
rect 122966 150996 122972 151060
rect 123036 151058 123042 151060
rect 139669 151058 139735 151061
rect 123036 151056 139735 151058
rect 123036 151000 139674 151056
rect 139730 151000 139735 151056
rect 123036 150998 139735 151000
rect 123036 150996 123042 150998
rect 139669 150995 139735 150998
rect 148910 150996 148916 151060
rect 148980 151058 148986 151060
rect 183645 151058 183711 151061
rect 148980 151056 183711 151058
rect 148980 151000 183650 151056
rect 183706 151000 183711 151056
rect 148980 150998 183711 151000
rect 148980 150996 148986 150998
rect 183645 150995 183711 150998
rect 122833 150514 122899 150517
rect 124070 150514 124076 150516
rect 122833 150512 124076 150514
rect 122833 150456 122838 150512
rect 122894 150456 124076 150512
rect 122833 150454 124076 150456
rect 122833 150451 122899 150454
rect 124070 150452 124076 150454
rect 124140 150514 124146 150516
rect 580257 150514 580323 150517
rect 124140 150512 580323 150514
rect 124140 150456 580262 150512
rect 580318 150456 580323 150512
rect 124140 150454 580323 150456
rect 124140 150452 124146 150454
rect 580257 150451 580323 150454
rect 168465 149970 168531 149973
rect 188286 149970 188292 149972
rect 168465 149968 188292 149970
rect -960 149834 480 149924
rect 168465 149912 168470 149968
rect 168526 149912 188292 149968
rect 168465 149910 188292 149912
rect 168465 149907 168531 149910
rect 188286 149908 188292 149910
rect 188356 149908 188362 149972
rect 3141 149834 3207 149837
rect -960 149832 3207 149834
rect -960 149776 3146 149832
rect 3202 149776 3207 149832
rect -960 149774 3207 149776
rect -960 149684 480 149774
rect 3141 149771 3207 149774
rect 167085 149834 167151 149837
rect 189390 149834 189396 149836
rect 167085 149832 189396 149834
rect 167085 149776 167090 149832
rect 167146 149776 189396 149832
rect 167085 149774 189396 149776
rect 167085 149771 167151 149774
rect 189390 149772 189396 149774
rect 189460 149772 189466 149836
rect 156822 149636 156828 149700
rect 156892 149698 156898 149700
rect 193765 149698 193831 149701
rect 156892 149696 193831 149698
rect 156892 149640 193770 149696
rect 193826 149640 193831 149696
rect 156892 149638 193831 149640
rect 156892 149636 156898 149638
rect 193765 149635 193831 149638
rect 197854 149092 197860 149156
rect 197924 149154 197930 149156
rect 198181 149154 198247 149157
rect 201033 149156 201099 149157
rect 200982 149154 200988 149156
rect 197924 149152 198247 149154
rect 197924 149096 198186 149152
rect 198242 149096 198247 149152
rect 197924 149094 198247 149096
rect 200942 149094 200988 149154
rect 201052 149152 201099 149156
rect 201094 149096 201099 149152
rect 197924 149092 197930 149094
rect 198181 149091 198247 149094
rect 200982 149092 200988 149094
rect 201052 149092 201099 149096
rect 201033 149091 201099 149092
rect 172513 149018 172579 149021
rect 197486 149018 197492 149020
rect 172513 149016 197492 149018
rect 172513 148960 172518 149016
rect 172574 148960 197492 149016
rect 172513 148958 197492 148960
rect 172513 148955 172579 148958
rect 197486 148956 197492 148958
rect 197556 148956 197562 149020
rect 175365 148882 175431 148885
rect 201902 148882 201908 148884
rect 175365 148880 201908 148882
rect 175365 148824 175370 148880
rect 175426 148824 201908 148880
rect 175365 148822 201908 148824
rect 175365 148819 175431 148822
rect 201902 148820 201908 148822
rect 201972 148820 201978 148884
rect 173750 148684 173756 148748
rect 173820 148746 173826 148748
rect 204897 148746 204963 148749
rect 173820 148744 204963 148746
rect 173820 148688 204902 148744
rect 204958 148688 204963 148744
rect 173820 148686 204963 148688
rect 173820 148684 173826 148686
rect 204897 148683 204963 148686
rect 103094 148548 103100 148612
rect 103164 148610 103170 148612
rect 135805 148610 135871 148613
rect 103164 148608 135871 148610
rect 103164 148552 135810 148608
rect 135866 148552 135871 148608
rect 103164 148550 135871 148552
rect 103164 148548 103170 148550
rect 135805 148547 135871 148550
rect 170622 148548 170628 148612
rect 170692 148610 170698 148612
rect 203374 148610 203380 148612
rect 170692 148550 203380 148610
rect 170692 148548 170698 148550
rect 203374 148548 203380 148550
rect 203444 148548 203450 148612
rect 104198 148412 104204 148476
rect 104268 148474 104274 148476
rect 136766 148474 136772 148476
rect 104268 148414 136772 148474
rect 104268 148412 104274 148414
rect 136766 148412 136772 148414
rect 136836 148412 136842 148476
rect 172697 148474 172763 148477
rect 205766 148474 205772 148476
rect 172697 148472 205772 148474
rect 172697 148416 172702 148472
rect 172758 148416 205772 148472
rect 172697 148414 205772 148416
rect 172697 148411 172763 148414
rect 205766 148412 205772 148414
rect 205836 148412 205842 148476
rect 119654 148276 119660 148340
rect 119724 148338 119730 148340
rect 153469 148338 153535 148341
rect 119724 148336 153535 148338
rect 119724 148280 153474 148336
rect 153530 148280 153535 148336
rect 119724 148278 153535 148280
rect 119724 148276 119730 148278
rect 153469 148275 153535 148278
rect 158478 148276 158484 148340
rect 158548 148338 158554 148340
rect 203609 148338 203675 148341
rect 158548 148336 203675 148338
rect 158548 148280 203614 148336
rect 203670 148280 203675 148336
rect 158548 148278 203675 148280
rect 158548 148276 158554 148278
rect 203609 148275 203675 148278
rect 172881 148202 172947 148205
rect 194726 148202 194732 148204
rect 172881 148200 194732 148202
rect 172881 148144 172886 148200
rect 172942 148144 194732 148200
rect 172881 148142 194732 148144
rect 172881 148139 172947 148142
rect 194726 148140 194732 148142
rect 194796 148140 194802 148204
rect 181437 147658 181503 147661
rect 199653 147658 199719 147661
rect 181437 147656 199719 147658
rect 181437 147600 181442 147656
rect 181498 147600 199658 147656
rect 199714 147600 199719 147656
rect 181437 147598 199719 147600
rect 181437 147595 181503 147598
rect 199653 147595 199719 147598
rect 112478 147460 112484 147524
rect 112548 147522 112554 147524
rect 131614 147522 131620 147524
rect 112548 147462 131620 147522
rect 112548 147460 112554 147462
rect 131614 147460 131620 147462
rect 131684 147460 131690 147524
rect 169845 147522 169911 147525
rect 196566 147522 196572 147524
rect 169845 147520 196572 147522
rect 169845 147464 169850 147520
rect 169906 147464 196572 147520
rect 169845 147462 196572 147464
rect 169845 147459 169911 147462
rect 196566 147460 196572 147462
rect 196636 147460 196642 147524
rect 113582 147324 113588 147388
rect 113652 147386 113658 147388
rect 137001 147386 137067 147389
rect 113652 147384 137067 147386
rect 113652 147328 137006 147384
rect 137062 147328 137067 147384
rect 113652 147326 137067 147328
rect 113652 147324 113658 147326
rect 137001 147323 137067 147326
rect 170857 147386 170923 147389
rect 210049 147386 210115 147389
rect 170857 147384 210115 147386
rect 170857 147328 170862 147384
rect 170918 147328 210054 147384
rect 210110 147328 210115 147384
rect 170857 147326 210115 147328
rect 170857 147323 170923 147326
rect 210049 147323 210115 147326
rect 115054 147188 115060 147252
rect 115124 147250 115130 147252
rect 138289 147250 138355 147253
rect 115124 147248 138355 147250
rect 115124 147192 138294 147248
rect 138350 147192 138355 147248
rect 115124 147190 138355 147192
rect 115124 147188 115130 147190
rect 138289 147187 138355 147190
rect 150014 147188 150020 147252
rect 150084 147250 150090 147252
rect 192661 147250 192727 147253
rect 150084 147248 192727 147250
rect 150084 147192 192666 147248
rect 192722 147192 192727 147248
rect 150084 147190 192727 147192
rect 150084 147188 150090 147190
rect 192661 147187 192727 147190
rect 122046 147052 122052 147116
rect 122116 147114 122122 147116
rect 147254 147114 147260 147116
rect 122116 147054 147260 147114
rect 122116 147052 122122 147054
rect 147254 147052 147260 147054
rect 147324 147052 147330 147116
rect 164233 147114 164299 147117
rect 207841 147114 207907 147117
rect 164233 147112 207907 147114
rect 164233 147056 164238 147112
rect 164294 147056 207846 147112
rect 207902 147056 207907 147112
rect 164233 147054 207907 147056
rect 164233 147051 164299 147054
rect 207841 147051 207907 147054
rect 102685 146978 102751 146981
rect 136582 146978 136588 146980
rect 102685 146976 136588 146978
rect 102685 146920 102690 146976
rect 102746 146920 136588 146976
rect 102685 146918 136588 146920
rect 102685 146915 102751 146918
rect 136582 146916 136588 146918
rect 136652 146916 136658 146980
rect 165705 146978 165771 146981
rect 214373 146978 214439 146981
rect 165705 146976 214439 146978
rect 165705 146920 165710 146976
rect 165766 146920 214378 146976
rect 214434 146920 214439 146976
rect 165705 146918 214439 146920
rect 165705 146915 165771 146918
rect 214373 146915 214439 146918
rect 115565 146298 115631 146301
rect 115790 146298 115796 146300
rect 115565 146296 115796 146298
rect 115565 146240 115570 146296
rect 115626 146240 115796 146296
rect 115565 146238 115796 146240
rect 115565 146235 115631 146238
rect 115790 146236 115796 146238
rect 115860 146236 115866 146300
rect 119429 146162 119495 146165
rect 146937 146162 147003 146165
rect 119429 146160 147003 146162
rect 119429 146104 119434 146160
rect 119490 146104 146942 146160
rect 146998 146104 147003 146160
rect 119429 146102 147003 146104
rect 119429 146099 119495 146102
rect 146937 146099 147003 146102
rect 180333 146162 180399 146165
rect 189758 146162 189764 146164
rect 180333 146160 189764 146162
rect 180333 146104 180338 146160
rect 180394 146104 189764 146160
rect 180333 146102 189764 146104
rect 180333 146099 180399 146102
rect 189758 146100 189764 146102
rect 189828 146100 189834 146164
rect 120758 145964 120764 146028
rect 120828 146026 120834 146028
rect 153377 146026 153443 146029
rect 120828 146024 153443 146026
rect 120828 145968 153382 146024
rect 153438 145968 153443 146024
rect 120828 145966 153443 145968
rect 120828 145964 120834 145966
rect 153377 145963 153443 145966
rect 180517 146026 180583 146029
rect 191598 146026 191604 146028
rect 180517 146024 191604 146026
rect 180517 145968 180522 146024
rect 180578 145968 191604 146024
rect 180517 145966 191604 145968
rect 180517 145963 180583 145966
rect 191598 145964 191604 145966
rect 191668 145964 191674 146028
rect 111006 145828 111012 145892
rect 111076 145890 111082 145892
rect 111241 145890 111307 145893
rect 111076 145888 111307 145890
rect 111076 145832 111246 145888
rect 111302 145832 111307 145888
rect 111076 145830 111307 145832
rect 111076 145828 111082 145830
rect 111241 145827 111307 145830
rect 112846 145828 112852 145892
rect 112916 145890 112922 145892
rect 147765 145890 147831 145893
rect 112916 145888 147831 145890
rect 112916 145832 147770 145888
rect 147826 145832 147831 145888
rect 112916 145830 147831 145832
rect 112916 145828 112922 145830
rect 147765 145827 147831 145830
rect 175273 145890 175339 145893
rect 187366 145890 187372 145892
rect 175273 145888 187372 145890
rect 175273 145832 175278 145888
rect 175334 145832 187372 145888
rect 175273 145830 187372 145832
rect 175273 145827 175339 145830
rect 187366 145828 187372 145830
rect 187436 145828 187442 145892
rect 112110 145692 112116 145756
rect 112180 145754 112186 145756
rect 151997 145754 152063 145757
rect 112180 145752 152063 145754
rect 112180 145696 152002 145752
rect 152058 145696 152063 145752
rect 112180 145694 152063 145696
rect 112180 145692 112186 145694
rect 151997 145691 152063 145694
rect 164233 145754 164299 145757
rect 196382 145754 196388 145756
rect 164233 145752 196388 145754
rect 164233 145696 164238 145752
rect 164294 145696 196388 145752
rect 164233 145694 196388 145696
rect 164233 145691 164299 145694
rect 196382 145692 196388 145694
rect 196452 145692 196458 145756
rect 115790 145556 115796 145620
rect 115860 145618 115866 145620
rect 156873 145618 156939 145621
rect 115860 145616 156939 145618
rect 115860 145560 156878 145616
rect 156934 145560 156939 145616
rect 115860 145558 156939 145560
rect 115860 145556 115866 145558
rect 156873 145555 156939 145558
rect 157333 145618 157399 145621
rect 192334 145618 192340 145620
rect 157333 145616 192340 145618
rect 157333 145560 157338 145616
rect 157394 145560 192340 145616
rect 157333 145558 192340 145560
rect 157333 145555 157399 145558
rect 192334 145556 192340 145558
rect 192404 145556 192410 145620
rect 112897 144802 112963 144805
rect 113030 144802 113036 144804
rect 112897 144800 113036 144802
rect 112897 144744 112902 144800
rect 112958 144744 113036 144800
rect 112897 144742 113036 144744
rect 112897 144739 112963 144742
rect 113030 144740 113036 144742
rect 113100 144740 113106 144804
rect 115606 144740 115612 144804
rect 115676 144802 115682 144804
rect 115841 144802 115907 144805
rect 115676 144800 115907 144802
rect 115676 144744 115846 144800
rect 115902 144744 115907 144800
rect 115676 144742 115907 144744
rect 115676 144740 115682 144742
rect 115841 144739 115907 144742
rect 116526 144740 116532 144804
rect 116596 144802 116602 144804
rect 117221 144802 117287 144805
rect 116596 144800 117287 144802
rect 116596 144744 117226 144800
rect 117282 144744 117287 144800
rect 116596 144742 117287 144744
rect 116596 144740 116602 144742
rect 117221 144739 117287 144742
rect 124765 144802 124831 144805
rect 125041 144802 125107 144805
rect 124765 144800 125107 144802
rect 124765 144744 124770 144800
rect 124826 144744 125046 144800
rect 125102 144744 125107 144800
rect 124765 144742 125107 144744
rect 124765 144739 124831 144742
rect 125041 144739 125107 144742
rect 165521 144802 165587 144805
rect 193622 144802 193628 144804
rect 165521 144800 193628 144802
rect 165521 144744 165526 144800
rect 165582 144744 193628 144800
rect 165521 144742 193628 144744
rect 165521 144739 165587 144742
rect 193622 144740 193628 144742
rect 193692 144740 193698 144804
rect 111558 144604 111564 144668
rect 111628 144666 111634 144668
rect 135897 144666 135963 144669
rect 111628 144664 135963 144666
rect 111628 144608 135902 144664
rect 135958 144608 135963 144664
rect 111628 144606 135963 144608
rect 111628 144604 111634 144606
rect 135897 144603 135963 144606
rect 162342 144604 162348 144668
rect 162412 144666 162418 144668
rect 194317 144666 194383 144669
rect 162412 144664 194383 144666
rect 162412 144608 194322 144664
rect 194378 144608 194383 144664
rect 162412 144606 194383 144608
rect 162412 144604 162418 144606
rect 194317 144603 194383 144606
rect 114134 144468 114140 144532
rect 114204 144530 114210 144532
rect 138657 144530 138723 144533
rect 114204 144528 138723 144530
rect 114204 144472 138662 144528
rect 138718 144472 138723 144528
rect 114204 144470 138723 144472
rect 114204 144468 114210 144470
rect 138657 144467 138723 144470
rect 156413 144530 156479 144533
rect 190494 144530 190500 144532
rect 156413 144528 190500 144530
rect 156413 144472 156418 144528
rect 156474 144472 190500 144528
rect 156413 144470 190500 144472
rect 156413 144467 156479 144470
rect 190494 144468 190500 144470
rect 190564 144468 190570 144532
rect 112662 144332 112668 144396
rect 112732 144394 112738 144396
rect 137553 144394 137619 144397
rect 112732 144392 137619 144394
rect 112732 144336 137558 144392
rect 137614 144336 137619 144392
rect 112732 144334 137619 144336
rect 112732 144332 112738 144334
rect 137553 144331 137619 144334
rect 154481 144394 154547 144397
rect 187693 144394 187759 144397
rect 154481 144392 187759 144394
rect 154481 144336 154486 144392
rect 154542 144336 187698 144392
rect 187754 144336 187759 144392
rect 154481 144334 187759 144336
rect 154481 144331 154547 144334
rect 187693 144331 187759 144334
rect 117589 144258 117655 144261
rect 147070 144258 147076 144260
rect 117589 144256 147076 144258
rect 117589 144200 117594 144256
rect 117650 144200 147076 144256
rect 117589 144198 147076 144200
rect 117589 144195 117655 144198
rect 147070 144196 147076 144198
rect 147140 144196 147146 144260
rect 152549 144258 152615 144261
rect 187141 144258 187207 144261
rect 152549 144256 187207 144258
rect 152549 144200 152554 144256
rect 152610 144200 187146 144256
rect 187202 144200 187207 144256
rect 152549 144198 187207 144200
rect 152549 144195 152615 144198
rect 187141 144195 187207 144198
rect 110873 144122 110939 144125
rect 143574 144122 143580 144124
rect 110873 144120 143580 144122
rect 110873 144064 110878 144120
rect 110934 144064 143580 144120
rect 110873 144062 143580 144064
rect 110873 144059 110939 144062
rect 143574 144060 143580 144062
rect 143644 144060 143650 144124
rect 153101 144122 153167 144125
rect 187509 144122 187575 144125
rect 153101 144120 187575 144122
rect 153101 144064 153106 144120
rect 153162 144064 187514 144120
rect 187570 144064 187575 144120
rect 153101 144062 187575 144064
rect 153101 144059 153167 144062
rect 187509 144059 187575 144062
rect 118141 143988 118207 143989
rect 118141 143984 118188 143988
rect 118252 143986 118258 143988
rect 138105 143986 138171 143989
rect 118141 143928 118146 143984
rect 118141 143924 118188 143928
rect 118252 143926 118298 143986
rect 122790 143984 138171 143986
rect 122790 143928 138110 143984
rect 138166 143928 138171 143984
rect 122790 143926 138171 143928
rect 118252 143924 118258 143926
rect 118141 143923 118207 143924
rect 116894 143788 116900 143852
rect 116964 143850 116970 143852
rect 122790 143850 122850 143926
rect 138105 143923 138171 143926
rect 116964 143790 122850 143850
rect 116964 143788 116970 143790
rect 124765 143578 124831 143581
rect 580349 143578 580415 143581
rect 124765 143576 580415 143578
rect 124765 143520 124770 143576
rect 124826 143520 580354 143576
rect 580410 143520 580415 143576
rect 124765 143518 580415 143520
rect 124765 143515 124831 143518
rect 580349 143515 580415 143518
rect 116710 143380 116716 143444
rect 116780 143442 116786 143444
rect 117221 143442 117287 143445
rect 116780 143440 117287 143442
rect 116780 143384 117226 143440
rect 117282 143384 117287 143440
rect 116780 143382 117287 143384
rect 116780 143380 116786 143382
rect 117221 143379 117287 143382
rect 183093 143442 183159 143445
rect 192334 143442 192340 143444
rect 183093 143440 192340 143442
rect 183093 143384 183098 143440
rect 183154 143384 192340 143440
rect 183093 143382 192340 143384
rect 183093 143379 183159 143382
rect 192334 143380 192340 143382
rect 192404 143380 192410 143444
rect 113950 143244 113956 143308
rect 114020 143306 114026 143308
rect 125685 143306 125751 143309
rect 114020 143304 125751 143306
rect 114020 143248 125690 143304
rect 125746 143248 125751 143304
rect 114020 143246 125751 143248
rect 114020 143244 114026 143246
rect 125685 143243 125751 143246
rect 184289 143306 184355 143309
rect 199009 143306 199075 143309
rect 184289 143304 199075 143306
rect 184289 143248 184294 143304
rect 184350 143248 199014 143304
rect 199070 143248 199075 143304
rect 184289 143246 199075 143248
rect 184289 143243 184355 143246
rect 199009 143243 199075 143246
rect 111190 143108 111196 143172
rect 111260 143170 111266 143172
rect 128261 143170 128327 143173
rect 111260 143168 128327 143170
rect 111260 143112 128266 143168
rect 128322 143112 128327 143168
rect 111260 143110 128327 143112
rect 111260 143108 111266 143110
rect 128261 143107 128327 143110
rect 183737 143170 183803 143173
rect 206093 143170 206159 143173
rect 183737 143168 206159 143170
rect 183737 143112 183742 143168
rect 183798 143112 206098 143168
rect 206154 143112 206159 143168
rect 183737 143110 206159 143112
rect 183737 143107 183803 143110
rect 206093 143107 206159 143110
rect 121126 142972 121132 143036
rect 121196 143034 121202 143036
rect 145005 143034 145071 143037
rect 121196 143032 145071 143034
rect 121196 142976 145010 143032
rect 145066 142976 145071 143032
rect 121196 142974 145071 142976
rect 121196 142972 121202 142974
rect 145005 142971 145071 142974
rect 161749 143034 161815 143037
rect 188889 143034 188955 143037
rect 161749 143032 188955 143034
rect 161749 142976 161754 143032
rect 161810 142976 188894 143032
rect 188950 142976 188955 143032
rect 161749 142974 188955 142976
rect 161749 142971 161815 142974
rect 188889 142971 188955 142974
rect 121310 142836 121316 142900
rect 121380 142898 121386 142900
rect 148041 142898 148107 142901
rect 121380 142896 148107 142898
rect 121380 142840 148046 142896
rect 148102 142840 148107 142896
rect 121380 142838 148107 142840
rect 121380 142836 121386 142838
rect 148041 142835 148107 142838
rect 156965 142898 157031 142901
rect 187734 142898 187740 142900
rect 156965 142896 187740 142898
rect 156965 142840 156970 142896
rect 157026 142840 187740 142896
rect 156965 142838 187740 142840
rect 156965 142835 157031 142838
rect 187734 142836 187740 142838
rect 187804 142836 187810 142900
rect 119705 142762 119771 142765
rect 146385 142762 146451 142765
rect 119705 142760 146451 142762
rect 119705 142704 119710 142760
rect 119766 142704 146390 142760
rect 146446 142704 146451 142760
rect 119705 142702 146451 142704
rect 119705 142699 119771 142702
rect 146385 142699 146451 142702
rect 178953 142762 179019 142765
rect 214097 142762 214163 142765
rect 178953 142760 214163 142762
rect 178953 142704 178958 142760
rect 179014 142704 214102 142760
rect 214158 142704 214163 142760
rect 178953 142702 214163 142704
rect 178953 142699 179019 142702
rect 214097 142699 214163 142702
rect 116526 142292 116532 142356
rect 116596 142354 116602 142356
rect 183737 142354 183803 142357
rect 116596 142352 183803 142354
rect 116596 142296 183742 142352
rect 183798 142296 183803 142352
rect 116596 142294 183803 142296
rect 116596 142292 116602 142294
rect 183737 142291 183803 142294
rect 111006 142156 111012 142220
rect 111076 142218 111082 142220
rect 184289 142218 184355 142221
rect 111076 142216 184355 142218
rect 111076 142160 184294 142216
rect 184350 142160 184355 142216
rect 111076 142158 184355 142160
rect 111076 142156 111082 142158
rect 184289 142155 184355 142158
rect 111374 142020 111380 142084
rect 111444 142082 111450 142084
rect 126145 142082 126211 142085
rect 111444 142080 126211 142082
rect 111444 142024 126150 142080
rect 126206 142024 126211 142080
rect 111444 142022 126211 142024
rect 111444 142020 111450 142022
rect 126145 142019 126211 142022
rect 157425 142082 157491 142085
rect 189206 142082 189212 142084
rect 157425 142080 189212 142082
rect 157425 142024 157430 142080
rect 157486 142024 189212 142080
rect 157425 142022 189212 142024
rect 157425 142019 157491 142022
rect 189206 142020 189212 142022
rect 189276 142020 189282 142084
rect 114134 141884 114140 141948
rect 114204 141946 114210 141948
rect 130469 141946 130535 141949
rect 114204 141944 130535 141946
rect 114204 141888 130474 141944
rect 130530 141888 130535 141944
rect 114204 141886 130535 141888
rect 114204 141884 114210 141886
rect 130469 141883 130535 141886
rect 108798 141748 108804 141812
rect 108868 141810 108874 141812
rect 139393 141810 139459 141813
rect 108868 141808 139459 141810
rect 108868 141752 139398 141808
rect 139454 141752 139459 141808
rect 108868 141750 139459 141752
rect 108868 141748 108874 141750
rect 139393 141747 139459 141750
rect 167453 141810 167519 141813
rect 192150 141810 192156 141812
rect 167453 141808 192156 141810
rect 167453 141752 167458 141808
rect 167514 141752 192156 141808
rect 167453 141750 192156 141752
rect 167453 141747 167519 141750
rect 192150 141748 192156 141750
rect 192220 141748 192226 141812
rect 121126 141612 121132 141676
rect 121196 141674 121202 141676
rect 153009 141674 153075 141677
rect 121196 141672 153075 141674
rect 121196 141616 153014 141672
rect 153070 141616 153075 141672
rect 121196 141614 153075 141616
rect 121196 141612 121202 141614
rect 153009 141611 153075 141614
rect 157149 141674 157215 141677
rect 189022 141674 189028 141676
rect 157149 141672 189028 141674
rect 157149 141616 157154 141672
rect 157210 141616 189028 141672
rect 157149 141614 189028 141616
rect 157149 141611 157215 141614
rect 189022 141612 189028 141614
rect 189092 141612 189098 141676
rect 116710 141476 116716 141540
rect 116780 141538 116786 141540
rect 155585 141538 155651 141541
rect 116780 141536 155651 141538
rect 116780 141480 155590 141536
rect 155646 141480 155651 141536
rect 116780 141478 155651 141480
rect 116780 141476 116786 141478
rect 155585 141475 155651 141478
rect 165470 141476 165476 141540
rect 165540 141538 165546 141540
rect 206093 141538 206159 141541
rect 165540 141536 206159 141538
rect 165540 141480 206098 141536
rect 206154 141480 206159 141536
rect 165540 141478 206159 141480
rect 165540 141476 165546 141478
rect 206093 141475 206159 141478
rect 117814 141340 117820 141404
rect 117884 141402 117890 141404
rect 177849 141402 177915 141405
rect 117884 141400 177915 141402
rect 117884 141344 177854 141400
rect 177910 141344 177915 141400
rect 117884 141342 177915 141344
rect 117884 141340 117890 141342
rect 177849 141339 177915 141342
rect 181897 141402 181963 141405
rect 190494 141402 190500 141404
rect 181897 141400 190500 141402
rect 181897 141344 181902 141400
rect 181958 141344 190500 141400
rect 181897 141342 190500 141344
rect 181897 141339 181963 141342
rect 190494 141340 190500 141342
rect 190564 141340 190570 141404
rect 113766 141204 113772 141268
rect 113836 141266 113842 141268
rect 126789 141266 126855 141269
rect 113836 141264 126855 141266
rect 113836 141208 126794 141264
rect 126850 141208 126855 141264
rect 113836 141206 126855 141208
rect 113836 141204 113842 141206
rect 126789 141203 126855 141206
rect 126789 140994 126855 140997
rect 464337 140994 464403 140997
rect 126789 140992 464403 140994
rect 126789 140936 126794 140992
rect 126850 140936 464342 140992
rect 464398 140936 464403 140992
rect 126789 140934 464403 140936
rect 126789 140931 126855 140934
rect 464337 140931 464403 140934
rect 126145 140858 126211 140861
rect 580625 140858 580691 140861
rect 126145 140856 580691 140858
rect 126145 140800 126150 140856
rect 126206 140800 580630 140856
rect 580686 140800 580691 140856
rect 126145 140798 580691 140800
rect 126145 140795 126211 140798
rect 580625 140795 580691 140798
rect 183001 140722 183067 140725
rect 193489 140724 193555 140725
rect 191046 140722 191052 140724
rect 183001 140720 191052 140722
rect 183001 140664 183006 140720
rect 183062 140664 191052 140720
rect 183001 140662 191052 140664
rect 183001 140659 183067 140662
rect 191046 140660 191052 140662
rect 191116 140660 191122 140724
rect 193438 140660 193444 140724
rect 193508 140722 193555 140724
rect 193508 140720 193600 140722
rect 193550 140664 193600 140720
rect 193508 140662 193600 140664
rect 193508 140660 193555 140662
rect 193489 140659 193555 140660
rect 119470 140524 119476 140588
rect 119540 140586 119546 140588
rect 126329 140586 126395 140589
rect 119540 140584 126395 140586
rect 119540 140528 126334 140584
rect 126390 140528 126395 140584
rect 119540 140526 126395 140528
rect 119540 140524 119546 140526
rect 126329 140523 126395 140526
rect 171133 140586 171199 140589
rect 185577 140586 185643 140589
rect 171133 140584 185643 140586
rect 171133 140528 171138 140584
rect 171194 140528 185582 140584
rect 185638 140528 185643 140584
rect 171133 140526 185643 140528
rect 171133 140523 171199 140526
rect 185577 140523 185643 140526
rect 189073 140586 189139 140589
rect 189574 140586 189580 140588
rect 189073 140584 189580 140586
rect 189073 140528 189078 140584
rect 189134 140528 189580 140584
rect 189073 140526 189580 140528
rect 189073 140523 189139 140526
rect 189574 140524 189580 140526
rect 189644 140524 189650 140588
rect 120942 140388 120948 140452
rect 121012 140450 121018 140452
rect 128997 140450 129063 140453
rect 121012 140448 129063 140450
rect 121012 140392 129002 140448
rect 129058 140392 129063 140448
rect 121012 140390 129063 140392
rect 121012 140388 121018 140390
rect 128997 140387 129063 140390
rect 169937 140450 170003 140453
rect 193438 140450 193444 140452
rect 169937 140448 193444 140450
rect 169937 140392 169942 140448
rect 169998 140392 193444 140448
rect 169937 140390 193444 140392
rect 169937 140387 170003 140390
rect 193438 140388 193444 140390
rect 193508 140388 193514 140452
rect 115606 140252 115612 140316
rect 115676 140314 115682 140316
rect 129457 140314 129523 140317
rect 115676 140312 129523 140314
rect 115676 140256 129462 140312
rect 129518 140256 129523 140312
rect 115676 140254 129523 140256
rect 115676 140252 115682 140254
rect 129457 140251 129523 140254
rect 169753 140314 169819 140317
rect 193622 140314 193628 140316
rect 169753 140312 193628 140314
rect 169753 140256 169758 140312
rect 169814 140256 193628 140312
rect 169753 140254 193628 140256
rect 169753 140251 169819 140254
rect 193622 140252 193628 140254
rect 193692 140252 193698 140316
rect 112294 140116 112300 140180
rect 112364 140178 112370 140180
rect 139945 140178 140011 140181
rect 112364 140176 140011 140178
rect 112364 140120 139950 140176
rect 140006 140120 140011 140176
rect 112364 140118 140011 140120
rect 112364 140116 112370 140118
rect 139945 140115 140011 140118
rect 161197 140178 161263 140181
rect 183369 140178 183435 140181
rect 185393 140180 185459 140181
rect 161197 140176 183435 140178
rect 161197 140120 161202 140176
rect 161258 140120 183374 140176
rect 183430 140120 183435 140176
rect 161197 140118 183435 140120
rect 161197 140115 161263 140118
rect 183369 140115 183435 140118
rect 185342 140116 185348 140180
rect 185412 140178 185459 140180
rect 185577 140178 185643 140181
rect 192150 140178 192156 140180
rect 185412 140176 185504 140178
rect 185454 140120 185504 140176
rect 185412 140118 185504 140120
rect 185577 140176 192156 140178
rect 185577 140120 185582 140176
rect 185638 140120 192156 140176
rect 185577 140118 192156 140120
rect 185412 140116 185459 140118
rect 185393 140115 185459 140116
rect 185577 140115 185643 140118
rect 192150 140116 192156 140118
rect 192220 140116 192226 140180
rect 122598 139980 122604 140044
rect 122668 140042 122674 140044
rect 124949 140042 125015 140045
rect 128905 140044 128971 140045
rect 130377 140044 130443 140045
rect 128854 140042 128860 140044
rect 122668 140040 125015 140042
rect 122668 139984 124954 140040
rect 125010 139984 125015 140040
rect 122668 139982 125015 139984
rect 128814 139982 128860 140042
rect 128924 140040 128971 140044
rect 130326 140042 130332 140044
rect 128966 139984 128971 140040
rect 122668 139980 122674 139982
rect 124949 139979 125015 139982
rect 128854 139980 128860 139982
rect 128924 139980 128971 139984
rect 130286 139982 130332 140042
rect 130396 140040 130443 140044
rect 177941 140042 178007 140045
rect 130438 139984 130443 140040
rect 130326 139980 130332 139982
rect 130396 139980 130443 139984
rect 128905 139979 128971 139980
rect 130377 139979 130443 139980
rect 132450 140040 178007 140042
rect 132450 139984 177946 140040
rect 178002 139984 178007 140040
rect 132450 139982 178007 139984
rect 120574 139844 120580 139908
rect 120644 139906 120650 139908
rect 132450 139906 132510 139982
rect 177941 139979 178007 139982
rect 180149 140042 180215 140045
rect 190678 140042 190684 140044
rect 180149 140040 190684 140042
rect 180149 139984 180154 140040
rect 180210 139984 190684 140040
rect 180149 139982 190684 139984
rect 180149 139979 180215 139982
rect 190678 139980 190684 139982
rect 190748 139980 190754 140044
rect 120644 139846 132510 139906
rect 183369 139906 183435 139909
rect 187182 139906 187188 139908
rect 183369 139904 187188 139906
rect 183369 139848 183374 139904
rect 183430 139848 187188 139904
rect 183369 139846 187188 139848
rect 120644 139844 120650 139846
rect 183369 139843 183435 139846
rect 187182 139844 187188 139846
rect 187252 139844 187258 139908
rect 181805 139770 181871 139773
rect 188102 139770 188108 139772
rect 181805 139768 188108 139770
rect 181805 139712 181810 139768
rect 181866 139712 188108 139768
rect 181805 139710 188108 139712
rect 181805 139707 181871 139710
rect 188102 139708 188108 139710
rect 188172 139708 188178 139772
rect 185577 139634 185643 139637
rect 187693 139636 187759 139637
rect 187693 139634 187740 139636
rect 185577 139632 187434 139634
rect 185577 139576 185582 139632
rect 185638 139576 187434 139632
rect 185577 139574 187434 139576
rect 187648 139632 187740 139634
rect 187648 139576 187698 139632
rect 187648 139574 187740 139576
rect 185577 139571 185643 139574
rect 118734 139436 118740 139500
rect 118804 139498 118810 139500
rect 119521 139498 119587 139501
rect 184381 139498 184447 139501
rect 186221 139498 186287 139501
rect 187374 139498 187434 139574
rect 187693 139572 187740 139574
rect 187804 139572 187810 139636
rect 187693 139571 187759 139572
rect 118804 139496 119587 139498
rect 118804 139440 119526 139496
rect 119582 139440 119587 139496
rect 118804 139438 119587 139440
rect 118804 139436 118810 139438
rect 119521 139435 119587 139438
rect 124078 139438 125794 139498
rect 111558 139300 111564 139364
rect 111628 139362 111634 139364
rect 123017 139362 123083 139365
rect 111628 139360 123083 139362
rect 111628 139304 123022 139360
rect 123078 139304 123083 139360
rect 111628 139302 123083 139304
rect 111628 139300 111634 139302
rect 123017 139299 123083 139302
rect 123150 139300 123156 139364
rect 123220 139362 123226 139364
rect 123937 139362 124003 139365
rect 123220 139360 124003 139362
rect 123220 139304 123942 139360
rect 123998 139304 124003 139360
rect 123220 139302 124003 139304
rect 123220 139300 123226 139302
rect 123937 139299 124003 139302
rect 116761 139226 116827 139229
rect 124078 139226 124138 139438
rect 125501 139362 125567 139365
rect 116761 139224 124138 139226
rect 116761 139168 116766 139224
rect 116822 139168 124138 139224
rect 116761 139166 124138 139168
rect 124446 139360 125567 139362
rect 124446 139304 125506 139360
rect 125562 139304 125567 139360
rect 124446 139302 125567 139304
rect 125734 139362 125794 139438
rect 169342 139438 169770 139498
rect 130561 139362 130627 139365
rect 125734 139360 130627 139362
rect 125734 139304 130566 139360
rect 130622 139304 130627 139360
rect 125734 139302 130627 139304
rect 116761 139163 116827 139166
rect 111190 139028 111196 139092
rect 111260 139090 111266 139092
rect 124446 139090 124506 139302
rect 125501 139299 125567 139302
rect 130561 139299 130627 139302
rect 130837 139362 130903 139365
rect 162301 139362 162367 139365
rect 169342 139362 169402 139438
rect 130837 139360 130946 139362
rect 130837 139304 130842 139360
rect 130898 139304 130946 139360
rect 130837 139299 130946 139304
rect 162301 139360 169402 139362
rect 162301 139304 162306 139360
rect 162362 139304 169402 139360
rect 162301 139302 169402 139304
rect 169477 139362 169543 139365
rect 169710 139362 169770 139438
rect 184381 139496 186146 139498
rect 184381 139440 184386 139496
rect 184442 139440 186146 139496
rect 184381 139438 186146 139440
rect 184381 139435 184447 139438
rect 173617 139362 173683 139365
rect 185894 139362 185900 139364
rect 169477 139360 169586 139362
rect 169477 139304 169482 139360
rect 169538 139304 169586 139360
rect 162301 139299 162367 139302
rect 169477 139299 169586 139304
rect 169710 139302 171150 139362
rect 111260 139030 124506 139090
rect 111260 139028 111266 139030
rect 115381 138954 115447 138957
rect 130886 138954 130946 139299
rect 115381 138952 130946 138954
rect 115381 138896 115386 138952
rect 115442 138896 130946 138952
rect 115381 138894 130946 138896
rect 115381 138891 115447 138894
rect 112345 138818 112411 138821
rect 130326 138818 130332 138820
rect 112345 138816 130332 138818
rect 112345 138760 112350 138816
rect 112406 138760 130332 138816
rect 112345 138758 130332 138760
rect 112345 138755 112411 138758
rect 130326 138756 130332 138758
rect 130396 138756 130402 138820
rect 169526 138818 169586 139299
rect 171090 138954 171150 139302
rect 173617 139360 185900 139362
rect 173617 139304 173622 139360
rect 173678 139304 185900 139360
rect 173617 139302 185900 139304
rect 173617 139299 173683 139302
rect 185894 139300 185900 139302
rect 185964 139300 185970 139364
rect 186086 139226 186146 139438
rect 186221 139496 187250 139498
rect 186221 139440 186226 139496
rect 186282 139440 187250 139496
rect 186221 139438 187250 139440
rect 187374 139438 188722 139498
rect 186221 139435 186287 139438
rect 186221 139362 186287 139365
rect 187049 139362 187115 139365
rect 186221 139360 187115 139362
rect 186221 139304 186226 139360
rect 186282 139304 187054 139360
rect 187110 139304 187115 139360
rect 186221 139302 187115 139304
rect 187190 139362 187250 139438
rect 188662 139362 188722 139438
rect 202086 139436 202092 139500
rect 202156 139498 202162 139500
rect 202505 139498 202571 139501
rect 202156 139496 202571 139498
rect 202156 139440 202510 139496
rect 202566 139440 202571 139496
rect 202156 139438 202571 139440
rect 202156 139436 202162 139438
rect 202505 139435 202571 139438
rect 192569 139362 192635 139365
rect 583520 139362 584960 139452
rect 187190 139302 188538 139362
rect 188662 139360 192635 139362
rect 188662 139304 192574 139360
rect 192630 139304 192635 139360
rect 188662 139302 192635 139304
rect 186221 139299 186287 139302
rect 187049 139299 187115 139302
rect 188245 139226 188311 139229
rect 186086 139224 188311 139226
rect 186086 139168 188250 139224
rect 188306 139168 188311 139224
rect 186086 139166 188311 139168
rect 188478 139226 188538 139302
rect 192569 139299 192635 139302
rect 583342 139302 584960 139362
rect 583342 139226 583402 139302
rect 583520 139226 584960 139302
rect 188478 139166 190470 139226
rect 583342 139212 584960 139226
rect 583342 139166 583586 139212
rect 188245 139163 188311 139166
rect 185342 139028 185348 139092
rect 185412 139090 185418 139092
rect 190410 139090 190470 139166
rect 193949 139090 194015 139093
rect 185412 139030 186514 139090
rect 190410 139088 194015 139090
rect 190410 139032 193954 139088
rect 194010 139032 194015 139088
rect 190410 139030 194015 139032
rect 185412 139028 185418 139030
rect 186262 138954 186268 138956
rect 171090 138894 186268 138954
rect 186262 138892 186268 138894
rect 186332 138892 186338 138956
rect 186454 138954 186514 139030
rect 193949 139027 194015 139030
rect 196617 138954 196683 138957
rect 186454 138952 196683 138954
rect 186454 138896 196622 138952
rect 196678 138896 196683 138952
rect 186454 138894 196683 138896
rect 196617 138891 196683 138894
rect 199377 138818 199443 138821
rect 169526 138816 199443 138818
rect 169526 138760 199382 138816
rect 199438 138760 199443 138816
rect 169526 138758 199443 138760
rect 199377 138755 199443 138758
rect 120717 138682 120783 138685
rect 146886 138682 146892 138684
rect 120717 138680 146892 138682
rect 120717 138624 120722 138680
rect 120778 138624 146892 138680
rect 120717 138622 146892 138624
rect 120717 138619 120783 138622
rect 146886 138620 146892 138622
rect 146956 138620 146962 138684
rect 169702 138620 169708 138684
rect 169772 138682 169778 138684
rect 201166 138682 201172 138684
rect 169772 138622 201172 138682
rect 169772 138620 169778 138622
rect 201166 138620 201172 138622
rect 201236 138620 201242 138684
rect 122230 138484 122236 138548
rect 122300 138546 122306 138548
rect 128854 138546 128860 138548
rect 122300 138486 128860 138546
rect 122300 138484 122306 138486
rect 128854 138484 128860 138486
rect 128924 138484 128930 138548
rect 122414 138138 122420 138140
rect 122238 138078 122420 138138
rect 116894 137940 116900 138004
rect 116964 138002 116970 138004
rect 122238 138002 122298 138078
rect 122414 138076 122420 138078
rect 122484 138076 122490 138140
rect 186446 138076 186452 138140
rect 186516 138138 186522 138140
rect 187601 138138 187667 138141
rect 186516 138136 187667 138138
rect 186516 138080 187606 138136
rect 187662 138080 187667 138136
rect 186516 138078 187667 138080
rect 186516 138076 186522 138078
rect 187601 138075 187667 138078
rect 187734 138076 187740 138140
rect 187804 138138 187810 138140
rect 583526 138138 583586 139166
rect 187804 138078 583586 138138
rect 187804 138076 187810 138078
rect 116964 137942 122298 138002
rect 116964 137940 116970 137942
rect 122414 137940 122420 138004
rect 122484 138002 122490 138004
rect 124806 138002 124812 138004
rect 122484 137942 124812 138002
rect 122484 137940 122490 137942
rect 124806 137940 124812 137942
rect 124876 137940 124882 138004
rect 181294 137940 181300 138004
rect 181364 138002 181370 138004
rect 181364 137942 190470 138002
rect 181364 137940 181370 137942
rect 185894 137804 185900 137868
rect 185964 137866 185970 137868
rect 190410 137866 190470 137942
rect 195421 137866 195487 137869
rect 185964 137806 186146 137866
rect 190410 137864 195487 137866
rect 190410 137808 195426 137864
rect 195482 137808 195487 137864
rect 190410 137806 195487 137808
rect 185964 137804 185970 137806
rect 118182 137396 118188 137460
rect 118252 137458 118258 137460
rect 122046 137458 122052 137460
rect 118252 137398 122052 137458
rect 118252 137396 118258 137398
rect 122046 137396 122052 137398
rect 122116 137396 122122 137460
rect 112846 137260 112852 137324
rect 112916 137322 112922 137324
rect 122966 137322 122972 137324
rect 112916 137262 122972 137322
rect 112916 137260 112922 137262
rect 122966 137260 122972 137262
rect 123036 137260 123042 137324
rect -960 136778 480 136868
rect 3233 136778 3299 136781
rect -960 136776 3299 136778
rect -960 136720 3238 136776
rect 3294 136720 3299 136776
rect -960 136718 3299 136720
rect -960 136628 480 136718
rect 3233 136715 3299 136718
rect 186086 136642 186146 137806
rect 195421 137803 195487 137806
rect 191189 136642 191255 136645
rect 186086 136640 191255 136642
rect 186086 136584 191194 136640
rect 191250 136584 191255 136640
rect 186086 136582 191255 136584
rect 191189 136579 191255 136582
rect 186262 135900 186268 135964
rect 186332 135962 186338 135964
rect 194041 135962 194107 135965
rect 186332 135960 194107 135962
rect 186332 135904 194046 135960
rect 194102 135904 194107 135960
rect 186332 135902 194107 135904
rect 186332 135900 186338 135902
rect 194041 135899 194107 135902
rect 121821 133922 121887 133925
rect 122966 133922 122972 133924
rect 121821 133920 122972 133922
rect 121821 133864 121826 133920
rect 121882 133864 122972 133920
rect 121821 133862 122972 133864
rect 121821 133859 121887 133862
rect 122966 133860 122972 133862
rect 123036 133860 123042 133924
rect 186078 131684 186084 131748
rect 186148 131684 186154 131748
rect 186086 131474 186146 131684
rect 186262 131474 186268 131476
rect 186086 131414 186268 131474
rect 186262 131412 186268 131414
rect 186332 131412 186338 131476
rect 580901 126034 580967 126037
rect 583520 126034 584960 126124
rect 580901 126032 584960 126034
rect 580901 125976 580906 126032
rect 580962 125976 584960 126032
rect 580901 125974 584960 125976
rect 580901 125971 580967 125974
rect 583520 125884 584960 125974
rect -960 123572 480 123812
rect 186078 117948 186084 118012
rect 186148 118010 186154 118012
rect 188429 118010 188495 118013
rect 186148 118008 188495 118010
rect 186148 117952 188434 118008
rect 188490 117952 188495 118008
rect 186148 117950 188495 117952
rect 186148 117948 186154 117950
rect 188429 117947 188495 117950
rect 580809 112842 580875 112845
rect 583520 112842 584960 112932
rect 580809 112840 584960 112842
rect 580809 112784 580814 112840
rect 580870 112784 584960 112840
rect 580809 112782 584960 112784
rect 580809 112779 580875 112782
rect 583520 112692 584960 112782
rect -960 110666 480 110756
rect 3049 110666 3115 110669
rect -960 110664 3115 110666
rect -960 110608 3054 110664
rect 3110 110608 3115 110664
rect -960 110606 3115 110608
rect -960 110516 480 110606
rect 3049 110603 3115 110606
rect 186262 104892 186268 104956
rect 186332 104954 186338 104956
rect 186630 104954 186636 104956
rect 186332 104894 186636 104954
rect 186332 104892 186338 104894
rect 186630 104892 186636 104894
rect 186700 104892 186706 104956
rect 580717 99514 580783 99517
rect 583520 99514 584960 99604
rect 580717 99512 584960 99514
rect 580717 99456 580722 99512
rect 580778 99456 584960 99512
rect 580717 99454 584960 99456
rect 580717 99451 580783 99454
rect 583520 99364 584960 99454
rect -960 97610 480 97700
rect -960 97550 674 97610
rect -960 97474 480 97550
rect 614 97474 674 97550
rect -960 97460 674 97474
rect 246 97414 674 97460
rect 246 96930 306 97414
rect 246 96870 6930 96930
rect 6870 96658 6930 96870
rect 118734 96658 118740 96660
rect 6870 96598 118740 96658
rect 118734 96596 118740 96598
rect 118804 96596 118810 96660
rect 186630 90340 186636 90404
rect 186700 90402 186706 90404
rect 189022 90402 189028 90404
rect 186700 90342 189028 90402
rect 186700 90340 186706 90342
rect 189022 90340 189028 90342
rect 189092 90340 189098 90404
rect 186078 86260 186084 86324
rect 186148 86322 186154 86324
rect 186630 86322 186636 86324
rect 186148 86262 186636 86322
rect 186148 86260 186154 86262
rect 186630 86260 186636 86262
rect 186700 86260 186706 86324
rect 120809 86186 120875 86189
rect 122966 86186 122972 86188
rect 120809 86184 122972 86186
rect 120809 86128 120814 86184
rect 120870 86128 122972 86184
rect 120809 86126 122972 86128
rect 120809 86123 120875 86126
rect 122966 86124 122972 86126
rect 123036 86124 123042 86188
rect 579613 86186 579679 86189
rect 583520 86186 584960 86276
rect 579613 86184 584960 86186
rect 579613 86128 579618 86184
rect 579674 86128 584960 86184
rect 579613 86126 584960 86128
rect 579613 86123 579679 86126
rect 121729 86050 121795 86053
rect 122966 86050 122972 86052
rect 121729 86048 122972 86050
rect 121729 85992 121734 86048
rect 121790 85992 122972 86048
rect 121729 85990 122972 85992
rect 121729 85987 121795 85990
rect 122966 85988 122972 85990
rect 123036 85988 123042 86052
rect 583520 86036 584960 86126
rect -960 84690 480 84780
rect -960 84630 6930 84690
rect -960 84540 480 84630
rect 6870 84282 6930 84630
rect 117814 84282 117820 84284
rect 6870 84222 117820 84282
rect 117814 84220 117820 84222
rect 117884 84220 117890 84284
rect 186078 82180 186084 82244
rect 186148 82242 186154 82244
rect 195421 82242 195487 82245
rect 186148 82240 195487 82242
rect 186148 82184 195426 82240
rect 195482 82184 195487 82240
rect 186148 82182 195487 82184
rect 186148 82180 186154 82182
rect 195421 82179 195487 82182
rect 186262 82044 186268 82108
rect 186332 82106 186338 82108
rect 191281 82106 191347 82109
rect 186332 82104 191347 82106
rect 186332 82048 191286 82104
rect 191342 82048 191347 82104
rect 186332 82046 191347 82048
rect 186332 82044 186338 82046
rect 191281 82043 191347 82046
rect 120717 81970 120783 81973
rect 122373 81970 122439 81973
rect 189809 81970 189875 81973
rect 120717 81968 122439 81970
rect 120717 81912 120722 81968
rect 120778 81912 122378 81968
rect 122434 81912 122439 81968
rect 120717 81910 122439 81912
rect 120717 81907 120783 81910
rect 122373 81907 122439 81910
rect 186086 81968 189875 81970
rect 186086 81912 189814 81968
rect 189870 81912 189875 81968
rect 186086 81910 189875 81912
rect 112110 81772 112116 81836
rect 112180 81834 112186 81836
rect 124070 81834 124076 81836
rect 112180 81774 124076 81834
rect 112180 81772 112186 81774
rect 124070 81772 124076 81774
rect 124140 81772 124146 81836
rect 184054 81772 184060 81836
rect 184124 81834 184130 81836
rect 186086 81834 186146 81910
rect 189809 81907 189875 81910
rect 184124 81774 186146 81834
rect 189533 81834 189599 81837
rect 196709 81834 196775 81837
rect 189533 81832 196775 81834
rect 189533 81776 189538 81832
rect 189594 81776 196714 81832
rect 196770 81776 196775 81832
rect 189533 81774 196775 81776
rect 184124 81772 184130 81774
rect 189533 81771 189599 81774
rect 196709 81771 196775 81774
rect 185342 81636 185348 81700
rect 185412 81698 185418 81700
rect 186630 81698 186636 81700
rect 185412 81638 186636 81698
rect 185412 81636 185418 81638
rect 186630 81636 186636 81638
rect 186700 81636 186706 81700
rect 178902 81500 178908 81564
rect 178972 81562 178978 81564
rect 189073 81562 189139 81565
rect 189574 81562 189580 81564
rect 178972 81502 183570 81562
rect 178972 81500 178978 81502
rect 183510 81426 183570 81502
rect 189073 81560 189580 81562
rect 189073 81504 189078 81560
rect 189134 81504 189580 81560
rect 189073 81502 189580 81504
rect 189073 81499 189139 81502
rect 189574 81500 189580 81502
rect 189644 81500 189650 81564
rect 196566 81500 196572 81564
rect 196636 81562 196642 81564
rect 196893 81562 196959 81565
rect 196636 81560 196959 81562
rect 196636 81504 196898 81560
rect 196954 81504 196959 81560
rect 196636 81502 196959 81504
rect 196636 81500 196642 81502
rect 196893 81499 196959 81502
rect 188521 81426 188587 81429
rect 183510 81424 188587 81426
rect 183510 81368 188526 81424
rect 188582 81368 188587 81424
rect 183510 81366 188587 81368
rect 188521 81363 188587 81366
rect 112253 81290 112319 81293
rect 121453 81290 121519 81293
rect 112253 81288 121519 81290
rect 112253 81232 112258 81288
rect 112314 81232 121458 81288
rect 121514 81232 121519 81288
rect 112253 81230 121519 81232
rect 112253 81227 112319 81230
rect 121453 81227 121519 81230
rect 175038 81228 175044 81292
rect 175108 81290 175114 81292
rect 197486 81290 197492 81292
rect 175108 81230 197492 81290
rect 175108 81228 175114 81230
rect 197486 81228 197492 81230
rect 197556 81228 197562 81292
rect 122189 81154 122255 81157
rect 146334 81154 146340 81156
rect 122189 81152 146340 81154
rect 122189 81096 122194 81152
rect 122250 81096 146340 81152
rect 122189 81094 146340 81096
rect 122189 81091 122255 81094
rect 146334 81092 146340 81094
rect 146404 81092 146410 81156
rect 175590 81092 175596 81156
rect 175660 81154 175666 81156
rect 205950 81154 205956 81156
rect 175660 81094 205956 81154
rect 175660 81092 175666 81094
rect 205950 81092 205956 81094
rect 206020 81092 206026 81156
rect 122281 81018 122347 81021
rect 149278 81018 149284 81020
rect 122281 81016 149284 81018
rect 122281 80960 122286 81016
rect 122342 80960 149284 81016
rect 122281 80958 149284 80960
rect 122281 80955 122347 80958
rect 149278 80956 149284 80958
rect 149348 80956 149354 81020
rect 177246 80956 177252 81020
rect 177316 81018 177322 81020
rect 202229 81018 202295 81021
rect 177316 81016 202295 81018
rect 177316 80960 202234 81016
rect 202290 80960 202295 81016
rect 177316 80958 202295 80960
rect 177316 80956 177322 80958
rect 202229 80955 202295 80958
rect 120441 80882 120507 80885
rect 148726 80882 148732 80884
rect 120441 80880 148732 80882
rect 120441 80824 120446 80880
rect 120502 80824 148732 80880
rect 120441 80822 148732 80824
rect 120441 80819 120507 80822
rect 148726 80820 148732 80822
rect 148796 80820 148802 80884
rect 206461 80882 206527 80885
rect 180520 80880 206527 80882
rect 180520 80824 206466 80880
rect 206522 80824 206527 80880
rect 180520 80822 206527 80824
rect 102593 80746 102659 80749
rect 102593 80744 131130 80746
rect 102593 80688 102598 80744
rect 102654 80688 131130 80744
rect 102593 80686 131130 80688
rect 102593 80683 102659 80686
rect 120809 80610 120875 80613
rect 122741 80610 122807 80613
rect 120809 80608 122807 80610
rect 120809 80552 120814 80608
rect 120870 80552 122746 80608
rect 122802 80552 122807 80608
rect 120809 80550 122807 80552
rect 131070 80610 131130 80686
rect 180520 80613 180580 80822
rect 206461 80819 206527 80822
rect 197302 80746 197308 80748
rect 186270 80686 197308 80746
rect 131941 80610 132007 80613
rect 131070 80608 132007 80610
rect 131070 80552 131946 80608
rect 132002 80552 132007 80608
rect 131070 80550 132007 80552
rect 120809 80547 120875 80550
rect 122741 80547 122807 80550
rect 131941 80547 132007 80550
rect 180517 80608 180583 80613
rect 186270 80610 186330 80686
rect 197302 80684 197308 80686
rect 197372 80746 197378 80748
rect 505093 80746 505159 80749
rect 197372 80744 505159 80746
rect 197372 80688 505098 80744
rect 505154 80688 505159 80744
rect 197372 80686 505159 80688
rect 197372 80684 197378 80686
rect 505093 80683 505159 80686
rect 180517 80552 180522 80608
rect 180578 80552 180583 80608
rect 180517 80547 180583 80552
rect 181486 80550 186330 80610
rect 117865 80474 117931 80477
rect 123937 80474 124003 80477
rect 181486 80474 181546 80550
rect 117865 80472 124003 80474
rect 117865 80416 117870 80472
rect 117926 80416 123942 80472
rect 123998 80416 124003 80472
rect 117865 80414 124003 80416
rect 117865 80411 117931 80414
rect 123937 80411 124003 80414
rect 171688 80414 181546 80474
rect 185761 80474 185827 80477
rect 192334 80474 192340 80476
rect 185761 80472 192340 80474
rect 185761 80416 185766 80472
rect 185822 80416 192340 80472
rect 185761 80414 192340 80416
rect 118182 80140 118188 80204
rect 118252 80202 118258 80204
rect 121821 80202 121887 80205
rect 118252 80200 121887 80202
rect 118252 80144 121826 80200
rect 121882 80144 121887 80200
rect 118252 80142 121887 80144
rect 118252 80140 118258 80142
rect 121821 80139 121887 80142
rect 131665 80202 131731 80205
rect 131665 80200 142354 80202
rect 131665 80144 131670 80200
rect 131726 80144 142354 80200
rect 131665 80142 142354 80144
rect 131665 80139 131731 80142
rect 128629 80066 128695 80069
rect 128629 80064 132740 80066
rect 128629 80008 128634 80064
rect 128690 80008 132740 80064
rect 128629 80006 132740 80008
rect 128629 80003 128695 80006
rect 126053 79930 126119 79933
rect 132539 79930 132605 79933
rect 126053 79928 132605 79930
rect 126053 79872 126058 79928
rect 126114 79872 132544 79928
rect 132600 79872 132605 79928
rect 126053 79870 132605 79872
rect 132680 79930 132740 80006
rect 142294 79967 142354 80142
rect 146518 80140 146524 80204
rect 146588 80202 146594 80204
rect 155718 80202 155724 80204
rect 146588 80142 147322 80202
rect 146588 80140 146594 80142
rect 147262 79967 147322 80142
rect 155220 80142 155724 80202
rect 155220 79967 155280 80142
rect 155718 80140 155724 80142
rect 155788 80140 155794 80204
rect 170806 80202 170812 80204
rect 170032 80142 170812 80202
rect 159030 80004 159036 80068
rect 159100 80066 159106 80068
rect 169518 80066 169524 80068
rect 159100 80006 160064 80066
rect 159100 80004 159106 80006
rect 133459 79962 133525 79967
rect 133091 79930 133157 79933
rect 132680 79928 133157 79930
rect 132680 79872 133096 79928
rect 133152 79872 133157 79928
rect 133459 79906 133464 79962
rect 133520 79906 133525 79962
rect 134747 79962 134813 79967
rect 138703 79964 138769 79967
rect 133459 79901 133525 79906
rect 132680 79870 133157 79872
rect 126053 79867 126119 79870
rect 132539 79867 132605 79870
rect 133091 79867 133157 79870
rect 133462 79797 133522 79901
rect 134006 79868 134012 79932
rect 134076 79930 134082 79932
rect 134471 79930 134537 79933
rect 134076 79928 134537 79930
rect 134076 79872 134476 79928
rect 134532 79872 134537 79928
rect 134747 79906 134752 79962
rect 134808 79906 134813 79962
rect 138430 79962 138769 79964
rect 135115 79932 135181 79933
rect 135110 79930 135116 79932
rect 134747 79901 134813 79906
rect 134076 79870 134537 79872
rect 134076 79868 134082 79870
rect 134471 79867 134537 79870
rect 132723 79794 132789 79797
rect 133270 79794 133276 79796
rect 132723 79792 133276 79794
rect 132723 79736 132728 79792
rect 132784 79736 133276 79792
rect 132723 79734 133276 79736
rect 132723 79731 132789 79734
rect 133270 79732 133276 79734
rect 133340 79732 133346 79796
rect 133462 79792 133571 79797
rect 133462 79736 133510 79792
rect 133566 79736 133571 79792
rect 133462 79734 133571 79736
rect 133505 79731 133571 79734
rect 133822 79732 133828 79796
rect 133892 79794 133898 79796
rect 134750 79794 134810 79901
rect 135024 79870 135116 79930
rect 135110 79868 135116 79870
rect 135180 79868 135186 79932
rect 135299 79930 135365 79933
rect 135478 79930 135484 79932
rect 135299 79928 135484 79930
rect 135299 79872 135304 79928
rect 135360 79872 135484 79928
rect 135299 79870 135484 79872
rect 135115 79867 135181 79868
rect 135299 79867 135365 79870
rect 135478 79868 135484 79870
rect 135548 79868 135554 79932
rect 135759 79930 135825 79933
rect 136030 79930 136036 79932
rect 135759 79928 136036 79930
rect 135759 79872 135764 79928
rect 135820 79872 136036 79928
rect 135759 79870 136036 79872
rect 135759 79867 135825 79870
rect 136030 79868 136036 79870
rect 136100 79868 136106 79932
rect 136771 79930 136837 79933
rect 137691 79932 137757 79933
rect 138059 79932 138125 79933
rect 138430 79932 138708 79962
rect 137502 79930 137508 79932
rect 136771 79928 137508 79930
rect 136771 79872 136776 79928
rect 136832 79872 137508 79928
rect 136771 79870 137508 79872
rect 136771 79867 136837 79870
rect 137502 79868 137508 79870
rect 137572 79868 137578 79932
rect 137686 79868 137692 79932
rect 137756 79930 137762 79932
rect 138054 79930 138060 79932
rect 137756 79870 137848 79930
rect 137968 79870 138060 79930
rect 137756 79868 137762 79870
rect 138054 79868 138060 79870
rect 138124 79868 138130 79932
rect 138422 79868 138428 79932
rect 138492 79906 138708 79932
rect 138764 79906 138769 79962
rect 139715 79962 139781 79967
rect 138492 79904 138769 79906
rect 138492 79868 138498 79904
rect 138703 79901 138769 79904
rect 138887 79930 138953 79933
rect 139158 79930 139164 79932
rect 138887 79928 139164 79930
rect 138887 79872 138892 79928
rect 138948 79872 139164 79928
rect 138887 79870 139164 79872
rect 137691 79867 137757 79868
rect 138059 79867 138125 79868
rect 138887 79867 138953 79870
rect 139158 79868 139164 79870
rect 139228 79868 139234 79932
rect 139715 79906 139720 79962
rect 139776 79930 139781 79962
rect 141095 79962 141161 79967
rect 139894 79930 139900 79932
rect 139776 79906 139900 79930
rect 139715 79901 139900 79906
rect 139718 79870 139900 79901
rect 139894 79868 139900 79870
rect 139964 79868 139970 79932
rect 140083 79928 140149 79933
rect 141095 79930 141100 79962
rect 140083 79872 140088 79928
rect 140144 79872 140149 79928
rect 140083 79867 140149 79872
rect 140638 79906 141100 79930
rect 141156 79906 141161 79962
rect 142291 79962 142357 79967
rect 143303 79964 143369 79967
rect 141555 79932 141621 79933
rect 140638 79901 141161 79906
rect 140638 79870 141158 79901
rect 133892 79734 134810 79794
rect 133892 79732 133898 79734
rect 135662 79732 135668 79796
rect 135732 79794 135738 79796
rect 136219 79794 136285 79797
rect 137139 79794 137205 79797
rect 135732 79792 136285 79794
rect 135732 79736 136224 79792
rect 136280 79736 136285 79792
rect 135732 79734 136285 79736
rect 135732 79732 135738 79734
rect 136219 79731 136285 79734
rect 136406 79792 137205 79794
rect 136406 79736 137144 79792
rect 137200 79736 137205 79792
rect 136406 79734 137205 79736
rect 133689 79658 133755 79661
rect 136406 79658 136466 79734
rect 137139 79731 137205 79734
rect 138238 79732 138244 79796
rect 138308 79794 138314 79796
rect 138611 79794 138677 79797
rect 138308 79792 138677 79794
rect 138308 79736 138616 79792
rect 138672 79736 138677 79792
rect 138308 79734 138677 79736
rect 138308 79732 138314 79734
rect 138611 79731 138677 79734
rect 139531 79794 139597 79797
rect 139894 79794 139900 79796
rect 139531 79792 139900 79794
rect 139531 79736 139536 79792
rect 139592 79736 139900 79792
rect 139531 79734 139900 79736
rect 139531 79731 139597 79734
rect 139894 79732 139900 79734
rect 139964 79732 139970 79796
rect 133689 79656 136466 79658
rect 133689 79600 133694 79656
rect 133750 79600 136466 79656
rect 133689 79598 136466 79600
rect 133689 79595 133755 79598
rect 136582 79596 136588 79660
rect 136652 79658 136658 79660
rect 136725 79658 136791 79661
rect 136652 79656 136791 79658
rect 136652 79600 136730 79656
rect 136786 79600 136791 79656
rect 136652 79598 136791 79600
rect 136652 79596 136658 79598
rect 136725 79595 136791 79598
rect 137553 79658 137619 79661
rect 140086 79658 140146 79867
rect 140267 79796 140333 79797
rect 140262 79732 140268 79796
rect 140332 79794 140338 79796
rect 140332 79734 140424 79794
rect 140332 79732 140338 79734
rect 140267 79731 140333 79732
rect 137553 79656 140146 79658
rect 137553 79600 137558 79656
rect 137614 79600 140146 79656
rect 137553 79598 140146 79600
rect 140313 79658 140379 79661
rect 140638 79658 140698 79870
rect 141550 79868 141556 79932
rect 141620 79930 141626 79932
rect 142107 79930 142173 79933
rect 141620 79870 141712 79930
rect 141926 79928 142173 79930
rect 141926 79872 142112 79928
rect 142168 79872 142173 79928
rect 142291 79906 142296 79962
rect 142352 79906 142357 79962
rect 143260 79962 143369 79964
rect 142291 79901 142357 79906
rect 141926 79870 142173 79872
rect 141620 79868 141626 79870
rect 141555 79867 141621 79868
rect 140865 79796 140931 79797
rect 140814 79794 140820 79796
rect 140774 79734 140820 79794
rect 140884 79792 140931 79796
rect 140926 79736 140931 79792
rect 140814 79732 140820 79734
rect 140884 79732 140931 79736
rect 140865 79731 140931 79732
rect 141509 79794 141575 79797
rect 141926 79794 141986 79870
rect 142107 79867 142173 79870
rect 142654 79868 142660 79932
rect 142724 79930 142730 79932
rect 143119 79930 143185 79933
rect 142724 79928 143185 79930
rect 142724 79872 143124 79928
rect 143180 79872 143185 79928
rect 142724 79870 143185 79872
rect 142724 79868 142730 79870
rect 143119 79867 143185 79870
rect 143260 79906 143308 79962
rect 143364 79906 143369 79962
rect 145235 79962 145301 79967
rect 146707 79964 146773 79967
rect 143260 79901 143369 79906
rect 142383 79826 142449 79831
rect 141509 79792 141986 79794
rect 141509 79736 141514 79792
rect 141570 79736 141986 79792
rect 141509 79734 141986 79736
rect 141509 79731 141575 79734
rect 142102 79732 142108 79796
rect 142172 79794 142178 79796
rect 142383 79794 142388 79826
rect 142172 79770 142388 79794
rect 142444 79770 142449 79826
rect 142172 79765 142449 79770
rect 142172 79734 142446 79765
rect 142172 79732 142178 79734
rect 143260 79661 143320 79901
rect 144126 79868 144132 79932
rect 144196 79930 144202 79932
rect 144591 79930 144657 79933
rect 145051 79930 145117 79933
rect 144196 79928 144657 79930
rect 144196 79872 144596 79928
rect 144652 79872 144657 79928
rect 144196 79870 144657 79872
rect 144196 79868 144202 79870
rect 144591 79867 144657 79870
rect 144870 79928 145117 79930
rect 144870 79872 145056 79928
rect 145112 79872 145117 79928
rect 145235 79906 145240 79962
rect 145296 79906 145301 79962
rect 146526 79962 146773 79964
rect 145235 79901 145301 79906
rect 145419 79928 145485 79933
rect 144870 79870 145117 79872
rect 143579 79796 143645 79797
rect 143574 79794 143580 79796
rect 143488 79734 143580 79794
rect 143574 79732 143580 79734
rect 143644 79732 143650 79796
rect 144545 79794 144611 79797
rect 144870 79794 144930 79870
rect 145051 79867 145117 79870
rect 144545 79792 144930 79794
rect 144545 79736 144550 79792
rect 144606 79736 144930 79792
rect 144545 79734 144930 79736
rect 143579 79731 143645 79732
rect 144545 79731 144611 79734
rect 140313 79656 140698 79658
rect 140313 79600 140318 79656
rect 140374 79600 140698 79656
rect 140313 79598 140698 79600
rect 140865 79658 140931 79661
rect 140998 79658 141004 79660
rect 140865 79656 141004 79658
rect 140865 79600 140870 79656
rect 140926 79600 141004 79656
rect 140865 79598 141004 79600
rect 137553 79595 137619 79598
rect 140313 79595 140379 79598
rect 140865 79595 140931 79598
rect 140998 79596 141004 79598
rect 141068 79596 141074 79660
rect 141877 79658 141943 79661
rect 142613 79658 142679 79661
rect 141877 79656 142679 79658
rect 141877 79600 141882 79656
rect 141938 79600 142618 79656
rect 142674 79600 142679 79656
rect 141877 79598 142679 79600
rect 141877 79595 141943 79598
rect 142613 79595 142679 79598
rect 143257 79656 143323 79661
rect 143257 79600 143262 79656
rect 143318 79600 143323 79656
rect 143257 79595 143323 79600
rect 135529 79522 135595 79525
rect 145238 79522 145298 79901
rect 145419 79872 145424 79928
rect 145480 79872 145485 79928
rect 145419 79867 145485 79872
rect 145598 79868 145604 79932
rect 145668 79930 145674 79932
rect 145879 79930 145945 79933
rect 145668 79928 145945 79930
rect 145668 79872 145884 79928
rect 145940 79872 145945 79928
rect 146526 79906 146712 79962
rect 146768 79906 146773 79962
rect 147259 79962 147325 79967
rect 146526 79904 146773 79906
rect 145668 79870 145945 79872
rect 145668 79868 145674 79870
rect 145879 79867 145945 79870
rect 146339 79894 146405 79899
rect 145422 79797 145482 79867
rect 146339 79838 146344 79894
rect 146400 79838 146405 79894
rect 146339 79833 146405 79838
rect 145422 79792 145531 79797
rect 145422 79736 145470 79792
rect 145526 79736 145531 79792
rect 145422 79734 145531 79736
rect 145465 79731 145531 79734
rect 146155 79792 146221 79797
rect 146155 79736 146160 79792
rect 146216 79736 146221 79792
rect 146155 79731 146221 79736
rect 145925 79658 145991 79661
rect 146158 79658 146218 79731
rect 146342 79661 146402 79833
rect 146526 79794 146586 79904
rect 146707 79901 146773 79904
rect 146886 79868 146892 79932
rect 146956 79930 146962 79932
rect 147075 79930 147141 79933
rect 146956 79928 147141 79930
rect 146956 79872 147080 79928
rect 147136 79872 147141 79928
rect 147259 79906 147264 79962
rect 147320 79906 147325 79962
rect 147259 79901 147325 79906
rect 147443 79962 147509 79967
rect 147443 79906 147448 79962
rect 147504 79906 147509 79962
rect 148547 79962 148613 79967
rect 149375 79964 149441 79967
rect 147627 79932 147693 79933
rect 147443 79901 147509 79906
rect 146956 79870 147141 79872
rect 146956 79868 146962 79870
rect 147075 79867 147141 79870
rect 146661 79794 146727 79797
rect 146526 79792 146727 79794
rect 146526 79736 146666 79792
rect 146722 79736 146727 79792
rect 146526 79734 146727 79736
rect 146661 79731 146727 79734
rect 147070 79732 147076 79796
rect 147140 79794 147146 79796
rect 147446 79794 147506 79901
rect 147622 79868 147628 79932
rect 147692 79930 147698 79932
rect 147692 79870 147784 79930
rect 148547 79906 148552 79962
rect 148608 79930 148613 79962
rect 149332 79962 149441 79964
rect 149332 79932 149380 79962
rect 148726 79930 148732 79932
rect 148608 79906 148732 79930
rect 148547 79901 148732 79906
rect 148550 79870 148732 79901
rect 147692 79868 147698 79870
rect 148726 79868 148732 79870
rect 148796 79868 148802 79932
rect 149278 79868 149284 79932
rect 149348 79906 149380 79932
rect 149436 79906 149441 79962
rect 150295 79964 150361 79967
rect 153607 79964 153673 79967
rect 150295 79962 150404 79964
rect 149348 79901 149441 79906
rect 149559 79930 149625 79933
rect 149830 79930 149836 79932
rect 149559 79928 149836 79930
rect 149348 79870 149392 79901
rect 149559 79872 149564 79928
rect 149620 79872 149836 79928
rect 149559 79870 149836 79872
rect 149348 79868 149354 79870
rect 147627 79867 147693 79868
rect 149559 79867 149625 79870
rect 149830 79868 149836 79870
rect 149900 79868 149906 79932
rect 150295 79906 150300 79962
rect 150356 79906 150404 79962
rect 153334 79962 153673 79964
rect 151215 79930 151281 79933
rect 151675 79932 151741 79933
rect 150295 79901 150404 79906
rect 147140 79734 147506 79794
rect 147140 79732 147146 79734
rect 147990 79732 147996 79796
rect 148060 79794 148066 79796
rect 148639 79794 148705 79797
rect 148060 79792 148705 79794
rect 148060 79736 148644 79792
rect 148700 79736 148705 79792
rect 148060 79734 148705 79736
rect 148060 79732 148066 79734
rect 148639 79731 148705 79734
rect 145925 79656 146218 79658
rect 145925 79600 145930 79656
rect 145986 79600 146218 79656
rect 145925 79598 146218 79600
rect 146293 79656 146402 79661
rect 146293 79600 146298 79656
rect 146354 79600 146402 79656
rect 146293 79598 146402 79600
rect 145925 79595 145991 79598
rect 146293 79595 146359 79598
rect 149646 79596 149652 79660
rect 149716 79658 149722 79660
rect 150344 79658 150404 79901
rect 150988 79928 151281 79930
rect 150988 79872 151220 79928
rect 151276 79872 151281 79928
rect 150988 79870 151281 79872
rect 150988 79661 151048 79870
rect 151215 79867 151281 79870
rect 151670 79868 151676 79932
rect 151740 79930 151746 79932
rect 152779 79930 152845 79933
rect 153142 79930 153148 79932
rect 151740 79870 151832 79930
rect 152779 79928 153148 79930
rect 152043 79894 152109 79899
rect 151740 79868 151746 79870
rect 151675 79867 151741 79868
rect 152043 79838 152048 79894
rect 152104 79838 152109 79894
rect 152779 79872 152784 79928
rect 152840 79872 153148 79928
rect 152779 79870 153148 79872
rect 152779 79867 152845 79870
rect 153142 79868 153148 79870
rect 153212 79868 153218 79932
rect 153334 79906 153612 79962
rect 153668 79906 153673 79962
rect 153334 79904 153673 79906
rect 152043 79833 152109 79838
rect 149716 79598 150404 79658
rect 150985 79656 151051 79661
rect 150985 79600 150990 79656
rect 151046 79600 151051 79656
rect 149716 79596 149722 79598
rect 150985 79595 151051 79600
rect 135529 79520 145298 79522
rect 135529 79464 135534 79520
rect 135590 79464 145298 79520
rect 135529 79462 145298 79464
rect 135529 79459 135595 79462
rect 146334 79460 146340 79524
rect 146404 79522 146410 79524
rect 146845 79522 146911 79525
rect 146404 79520 146911 79522
rect 146404 79464 146850 79520
rect 146906 79464 146911 79520
rect 146404 79462 146911 79464
rect 152046 79522 152106 79833
rect 153334 79794 153394 79904
rect 153607 79901 153673 79904
rect 153791 79962 153857 79967
rect 153975 79964 154041 79967
rect 153791 79906 153796 79962
rect 153852 79906 153857 79962
rect 153791 79901 153857 79906
rect 153932 79962 154041 79964
rect 153932 79906 153980 79962
rect 154036 79906 154041 79962
rect 154895 79964 154961 79967
rect 154895 79962 155004 79964
rect 153932 79901 154041 79906
rect 154159 79930 154225 79933
rect 154430 79930 154436 79932
rect 154159 79928 154436 79930
rect 153150 79734 153394 79794
rect 152590 79596 152596 79660
rect 152660 79658 152666 79660
rect 152733 79658 152799 79661
rect 152660 79656 152799 79658
rect 152660 79600 152738 79656
rect 152794 79600 152799 79656
rect 152660 79598 152799 79600
rect 152660 79596 152666 79598
rect 152733 79595 152799 79598
rect 152733 79522 152799 79525
rect 152046 79520 152799 79522
rect 152046 79464 152738 79520
rect 152794 79464 152799 79520
rect 152046 79462 152799 79464
rect 153150 79522 153210 79734
rect 153285 79658 153351 79661
rect 153794 79658 153854 79901
rect 153932 79797 153992 79901
rect 154159 79872 154164 79928
rect 154220 79872 154436 79928
rect 154159 79870 154436 79872
rect 154159 79867 154225 79870
rect 154430 79868 154436 79870
rect 154500 79868 154506 79932
rect 154895 79906 154900 79962
rect 154956 79932 155004 79962
rect 155220 79962 155329 79967
rect 154956 79906 154988 79932
rect 154895 79901 154988 79906
rect 154944 79870 154988 79901
rect 154982 79868 154988 79870
rect 155052 79868 155058 79932
rect 155220 79906 155268 79962
rect 155324 79906 155329 79962
rect 156459 79962 156525 79967
rect 155220 79904 155329 79906
rect 155263 79901 155329 79904
rect 155631 79930 155697 79933
rect 155902 79930 155908 79932
rect 155631 79928 155908 79930
rect 155631 79872 155636 79928
rect 155692 79872 155908 79928
rect 155631 79870 155908 79872
rect 155631 79867 155697 79870
rect 155902 79868 155908 79870
rect 155972 79868 155978 79932
rect 156459 79906 156464 79962
rect 156520 79906 156525 79962
rect 157563 79962 157629 79967
rect 156459 79901 156525 79906
rect 156091 79894 156157 79899
rect 156091 79838 156096 79894
rect 156152 79838 156157 79894
rect 156091 79833 156157 79838
rect 153929 79792 153995 79797
rect 153929 79736 153934 79792
rect 153990 79736 153995 79792
rect 153929 79731 153995 79736
rect 154205 79794 154271 79797
rect 154205 79792 154314 79794
rect 154205 79736 154210 79792
rect 154266 79736 154314 79792
rect 154205 79731 154314 79736
rect 153285 79656 153854 79658
rect 153285 79600 153290 79656
rect 153346 79600 153854 79656
rect 153285 79598 153854 79600
rect 153285 79595 153351 79598
rect 153561 79522 153627 79525
rect 153150 79520 153627 79522
rect 153150 79464 153566 79520
rect 153622 79464 153627 79520
rect 153150 79462 153627 79464
rect 146404 79460 146410 79462
rect 146845 79459 146911 79462
rect 152733 79459 152799 79462
rect 153561 79459 153627 79462
rect 153878 79460 153884 79524
rect 153948 79522 153954 79524
rect 154254 79522 154314 79731
rect 156094 79661 156154 79833
rect 156462 79794 156522 79901
rect 156638 79868 156644 79932
rect 156708 79930 156714 79932
rect 157287 79930 157353 79933
rect 156708 79928 157353 79930
rect 156708 79872 157292 79928
rect 157348 79872 157353 79928
rect 157563 79906 157568 79962
rect 157624 79906 157629 79962
rect 157563 79901 157629 79906
rect 158023 79964 158089 79967
rect 158023 79962 158132 79964
rect 158023 79906 158028 79962
rect 158084 79932 158132 79962
rect 158299 79962 158365 79967
rect 158575 79964 158641 79967
rect 158084 79906 158116 79932
rect 158023 79901 158116 79906
rect 156708 79870 157353 79872
rect 156708 79868 156714 79870
rect 157287 79867 157353 79870
rect 156822 79794 156828 79796
rect 156462 79734 156828 79794
rect 156822 79732 156828 79734
rect 156892 79732 156898 79796
rect 156045 79656 156154 79661
rect 156045 79600 156050 79656
rect 156106 79600 156154 79656
rect 156045 79598 156154 79600
rect 156597 79658 156663 79661
rect 157190 79658 157196 79660
rect 156597 79656 157196 79658
rect 156597 79600 156602 79656
rect 156658 79600 157196 79656
rect 156597 79598 157196 79600
rect 156045 79595 156111 79598
rect 156597 79595 156663 79598
rect 157190 79596 157196 79598
rect 157260 79596 157266 79660
rect 157566 79658 157626 79901
rect 158072 79870 158116 79901
rect 158110 79868 158116 79870
rect 158180 79868 158186 79932
rect 158299 79906 158304 79962
rect 158360 79906 158365 79962
rect 158532 79962 158641 79964
rect 158532 79932 158580 79962
rect 158299 79901 158365 79906
rect 158302 79794 158362 79901
rect 158478 79868 158484 79932
rect 158548 79906 158580 79932
rect 158636 79906 158641 79962
rect 158548 79901 158641 79906
rect 159127 79930 159193 79933
rect 159398 79930 159404 79932
rect 159127 79928 159404 79930
rect 158548 79870 158592 79901
rect 159127 79872 159132 79928
rect 159188 79872 159404 79928
rect 159127 79870 159404 79872
rect 158548 79868 158554 79870
rect 159127 79867 159193 79870
rect 159398 79868 159404 79870
rect 159468 79868 159474 79932
rect 160004 79831 160064 80006
rect 169204 80006 169524 80066
rect 162347 79962 162413 79967
rect 162623 79964 162689 79967
rect 160875 79930 160941 79933
rect 161054 79930 161060 79932
rect 160875 79928 161060 79930
rect 160875 79872 160880 79928
rect 160936 79872 161060 79928
rect 160875 79870 161060 79872
rect 160875 79867 160941 79870
rect 161054 79868 161060 79870
rect 161124 79868 161130 79932
rect 161427 79930 161493 79933
rect 161979 79932 162045 79933
rect 162347 79932 162352 79962
rect 162408 79932 162413 79962
rect 162580 79962 162689 79964
rect 161974 79930 161980 79932
rect 161384 79928 161493 79930
rect 161384 79872 161432 79928
rect 161488 79872 161493 79928
rect 161384 79867 161493 79872
rect 161888 79870 161980 79930
rect 161974 79868 161980 79870
rect 162044 79868 162050 79932
rect 162342 79868 162348 79932
rect 162412 79930 162418 79932
rect 162412 79870 162470 79930
rect 162580 79906 162628 79962
rect 162684 79930 162689 79962
rect 163451 79962 163517 79967
rect 162894 79930 162900 79932
rect 162684 79906 162900 79930
rect 162580 79870 162900 79906
rect 162412 79868 162418 79870
rect 162894 79868 162900 79870
rect 162964 79868 162970 79932
rect 163267 79928 163333 79933
rect 163267 79872 163272 79928
rect 163328 79872 163333 79928
rect 163451 79906 163456 79962
rect 163512 79930 163517 79962
rect 166395 79962 166461 79967
rect 167223 79964 167289 79967
rect 163512 79906 164388 79930
rect 163451 79901 164388 79906
rect 161979 79867 162045 79868
rect 163267 79867 163333 79872
rect 163454 79870 164388 79901
rect 160004 79826 160113 79831
rect 158662 79794 158668 79796
rect 158302 79734 158668 79794
rect 158662 79732 158668 79734
rect 158732 79732 158738 79796
rect 159403 79792 159469 79797
rect 159403 79736 159408 79792
rect 159464 79736 159469 79792
rect 160004 79770 160052 79826
rect 160108 79770 160113 79826
rect 160004 79768 160113 79770
rect 160047 79765 160113 79768
rect 159403 79731 159469 79736
rect 161238 79732 161244 79796
rect 161308 79794 161314 79796
rect 161384 79794 161444 79867
rect 161308 79734 161444 79794
rect 162531 79794 162597 79797
rect 162710 79794 162716 79796
rect 162531 79792 162716 79794
rect 162531 79736 162536 79792
rect 162592 79736 162716 79792
rect 162531 79734 162716 79736
rect 161308 79732 161314 79734
rect 162531 79731 162597 79734
rect 162710 79732 162716 79734
rect 162780 79732 162786 79796
rect 163078 79732 163084 79796
rect 163148 79794 163154 79796
rect 163270 79794 163330 79867
rect 163148 79734 163330 79794
rect 163405 79796 163471 79797
rect 163405 79792 163452 79796
rect 163516 79794 163522 79796
rect 163405 79736 163410 79792
rect 163148 79732 163154 79734
rect 163405 79732 163452 79736
rect 163516 79734 163562 79794
rect 163635 79792 163701 79797
rect 163635 79736 163640 79792
rect 163696 79736 163701 79792
rect 163516 79732 163522 79734
rect 163405 79731 163471 79732
rect 163635 79731 163701 79736
rect 158621 79658 158687 79661
rect 157566 79656 158687 79658
rect 157566 79600 158626 79656
rect 158682 79600 158687 79656
rect 157566 79598 158687 79600
rect 159406 79658 159466 79731
rect 162158 79658 162164 79660
rect 159406 79598 162164 79658
rect 158621 79595 158687 79598
rect 162158 79596 162164 79598
rect 162228 79596 162234 79660
rect 163262 79596 163268 79660
rect 163332 79658 163338 79660
rect 163638 79658 163698 79731
rect 164328 79661 164388 79870
rect 164555 79928 164621 79933
rect 164555 79872 164560 79928
rect 164616 79872 164621 79928
rect 164555 79867 164621 79872
rect 165015 79930 165081 79933
rect 165843 79930 165909 79933
rect 166206 79930 166212 79932
rect 165015 79928 165124 79930
rect 165015 79872 165020 79928
rect 165076 79872 165124 79928
rect 165015 79867 165124 79872
rect 165843 79928 166212 79930
rect 165843 79872 165848 79928
rect 165904 79872 166212 79928
rect 165843 79870 166212 79872
rect 165843 79867 165909 79870
rect 166206 79868 166212 79870
rect 166276 79868 166282 79932
rect 166395 79906 166400 79962
rect 166456 79930 166461 79962
rect 167180 79962 167289 79964
rect 166574 79930 166580 79932
rect 166456 79906 166580 79930
rect 166395 79901 166580 79906
rect 166398 79870 166580 79901
rect 166574 79868 166580 79870
rect 166644 79868 166650 79932
rect 167180 79906 167228 79962
rect 167284 79906 167289 79962
rect 167180 79901 167289 79906
rect 168051 79962 168117 79967
rect 168051 79906 168056 79962
rect 168112 79906 168117 79962
rect 168603 79962 168669 79967
rect 168051 79901 168117 79906
rect 168235 79928 168301 79933
rect 168603 79930 168608 79962
rect 167039 79896 167105 79899
rect 166904 79894 167105 79896
rect 163332 79598 163698 79658
rect 164325 79656 164391 79661
rect 164325 79600 164330 79656
rect 164386 79600 164391 79656
rect 163332 79596 163338 79598
rect 164325 79595 164391 79600
rect 164558 79658 164618 79867
rect 164785 79658 164851 79661
rect 164558 79656 164851 79658
rect 164558 79600 164790 79656
rect 164846 79600 164851 79656
rect 164558 79598 164851 79600
rect 165064 79660 165124 79867
rect 166904 79838 167044 79894
rect 167100 79838 167105 79894
rect 166904 79836 167105 79838
rect 165291 79796 165357 79797
rect 165475 79796 165541 79797
rect 165286 79794 165292 79796
rect 165200 79734 165292 79794
rect 165286 79732 165292 79734
rect 165356 79732 165362 79796
rect 165470 79732 165476 79796
rect 165540 79794 165546 79796
rect 166671 79794 166737 79797
rect 165540 79734 165632 79794
rect 166671 79792 166780 79794
rect 166671 79736 166676 79792
rect 166732 79736 166780 79792
rect 165540 79732 165546 79734
rect 165291 79731 165357 79732
rect 165475 79731 165541 79732
rect 166671 79731 166780 79736
rect 165064 79598 165108 79660
rect 164785 79595 164851 79598
rect 165102 79596 165108 79598
rect 165172 79596 165178 79660
rect 166073 79658 166139 79661
rect 166720 79660 166780 79731
rect 166904 79760 166964 79836
rect 167039 79833 167105 79836
rect 167180 79794 167240 79901
rect 167310 79794 167316 79796
rect 166904 79700 167010 79760
rect 167180 79734 167316 79794
rect 167310 79732 167316 79734
rect 167380 79732 167386 79796
rect 167499 79794 167565 79797
rect 167862 79794 167868 79796
rect 167499 79792 167868 79794
rect 167499 79736 167504 79792
rect 167560 79736 167868 79792
rect 167499 79734 167868 79736
rect 167499 79731 167565 79734
rect 167862 79732 167868 79734
rect 167932 79732 167938 79796
rect 166950 79661 167010 79700
rect 168054 79661 168114 79901
rect 168235 79872 168240 79928
rect 168296 79872 168301 79928
rect 168235 79867 168301 79872
rect 168422 79906 168608 79930
rect 168664 79906 168669 79962
rect 168422 79901 168669 79906
rect 168879 79964 168945 79967
rect 168879 79962 168988 79964
rect 168879 79906 168884 79962
rect 168940 79930 168988 79962
rect 169204 79930 169264 80006
rect 169518 80004 169524 80006
rect 169588 80004 169594 80068
rect 170032 79967 170092 80142
rect 170806 80140 170812 80142
rect 170876 80140 170882 80204
rect 171688 79967 171748 80414
rect 185761 80411 185827 80414
rect 192334 80412 192340 80414
rect 192404 80412 192410 80476
rect 177246 80338 177252 80340
rect 172286 80278 177252 80338
rect 172286 79967 172346 80278
rect 177246 80276 177252 80278
rect 177316 80276 177322 80340
rect 184238 80276 184244 80340
rect 184308 80338 184314 80340
rect 189717 80338 189783 80341
rect 184308 80336 189783 80338
rect 184308 80280 189722 80336
rect 189778 80280 189783 80336
rect 184308 80278 189783 80280
rect 184308 80276 184314 80278
rect 189717 80275 189783 80278
rect 184197 80202 184263 80205
rect 186446 80202 186452 80204
rect 176104 80200 186452 80202
rect 176104 80144 184202 80200
rect 184258 80144 186452 80200
rect 176104 80142 186452 80144
rect 173566 80004 173572 80068
rect 173636 80066 173642 80068
rect 173636 80004 173680 80066
rect 169983 79962 170092 79967
rect 169339 79932 169405 79933
rect 168940 79906 169264 79930
rect 168879 79901 169264 79906
rect 168422 79870 168666 79901
rect 168928 79870 169264 79901
rect 168238 79797 168298 79867
rect 168238 79792 168347 79797
rect 168238 79736 168286 79792
rect 168342 79736 168347 79792
rect 168238 79734 168347 79736
rect 168281 79731 168347 79734
rect 168422 79661 168482 79870
rect 169334 79868 169340 79932
rect 169404 79930 169410 79932
rect 169404 79870 169496 79930
rect 169983 79906 169988 79962
rect 170044 79906 170092 79962
rect 170535 79964 170601 79967
rect 170535 79962 170644 79964
rect 169983 79904 170092 79906
rect 170259 79928 170325 79933
rect 169983 79901 170049 79904
rect 170259 79872 170264 79928
rect 170320 79872 170325 79928
rect 170535 79906 170540 79962
rect 170596 79932 170644 79962
rect 170811 79962 170877 79967
rect 170596 79906 170628 79932
rect 170535 79901 170628 79906
rect 169404 79868 169410 79870
rect 169339 79867 169405 79868
rect 170259 79867 170325 79872
rect 170584 79870 170628 79901
rect 170622 79868 170628 79870
rect 170692 79868 170698 79932
rect 170811 79906 170816 79962
rect 170872 79906 170877 79962
rect 170811 79901 170877 79906
rect 171639 79962 171748 79967
rect 171639 79906 171644 79962
rect 171700 79906 171748 79962
rect 171639 79904 171748 79906
rect 171915 79962 171981 79967
rect 171915 79906 171920 79962
rect 171976 79906 171981 79962
rect 172283 79962 172349 79967
rect 171639 79901 171705 79904
rect 171915 79901 171981 79906
rect 170029 79792 170095 79797
rect 170029 79736 170034 79792
rect 170090 79736 170095 79792
rect 170029 79731 170095 79736
rect 170032 79661 170092 79731
rect 170262 79661 170322 79867
rect 170622 79732 170628 79796
rect 170692 79794 170698 79796
rect 170814 79794 170874 79901
rect 170692 79734 170874 79794
rect 171918 79794 171978 79901
rect 172094 79868 172100 79932
rect 172164 79930 172170 79932
rect 172283 79930 172288 79962
rect 172164 79906 172288 79930
rect 172344 79906 172349 79962
rect 172164 79901 172349 79906
rect 172743 79964 172809 79967
rect 172743 79962 172852 79964
rect 172743 79906 172748 79962
rect 172804 79906 172852 79962
rect 173203 79932 173269 79933
rect 173198 79930 173204 79932
rect 172743 79901 172852 79906
rect 172164 79870 172346 79901
rect 172164 79868 172170 79870
rect 172792 79797 172852 79901
rect 173112 79870 173204 79930
rect 173198 79868 173204 79870
rect 173268 79868 173274 79932
rect 173479 79930 173545 79933
rect 173620 79930 173680 80004
rect 176104 79967 176164 80142
rect 184197 80139 184263 80142
rect 186446 80140 186452 80142
rect 186516 80140 186522 80204
rect 185526 80004 185532 80068
rect 185596 80066 185602 80068
rect 186262 80066 186268 80068
rect 185596 80006 186268 80066
rect 185596 80004 185602 80006
rect 186262 80004 186268 80006
rect 186332 80004 186338 80068
rect 200798 80004 200804 80068
rect 200868 80066 200874 80068
rect 201033 80066 201099 80069
rect 200868 80064 201099 80066
rect 200868 80008 201038 80064
rect 201094 80008 201099 80064
rect 200868 80006 201099 80008
rect 200868 80004 200874 80006
rect 201033 80003 201099 80006
rect 173479 79928 173680 79930
rect 173479 79872 173484 79928
rect 173540 79872 173680 79928
rect 173755 79962 173821 79967
rect 173755 79906 173760 79962
rect 173816 79930 173821 79962
rect 174675 79962 174741 79967
rect 173934 79930 173940 79932
rect 173816 79906 173940 79930
rect 173755 79901 173940 79906
rect 173479 79870 173680 79872
rect 173758 79870 173940 79901
rect 173203 79867 173269 79868
rect 173479 79867 173545 79870
rect 173934 79868 173940 79870
rect 174004 79868 174010 79932
rect 174491 79930 174557 79933
rect 174126 79928 174557 79930
rect 174126 79872 174496 79928
rect 174552 79872 174557 79928
rect 174675 79906 174680 79962
rect 174736 79906 174741 79962
rect 174675 79901 174741 79906
rect 174951 79964 175017 79967
rect 174951 79962 175060 79964
rect 174951 79906 174956 79962
rect 175012 79906 175060 79962
rect 175779 79962 175845 79967
rect 174951 79901 175060 79906
rect 174126 79870 174557 79872
rect 172278 79794 172284 79796
rect 171918 79734 172284 79794
rect 170692 79732 170698 79734
rect 172278 79732 172284 79734
rect 172348 79732 172354 79796
rect 172651 79792 172717 79797
rect 172651 79736 172656 79792
rect 172712 79736 172717 79792
rect 172651 79731 172717 79736
rect 172789 79792 172855 79797
rect 172789 79736 172794 79792
rect 172850 79736 172855 79792
rect 172789 79731 172855 79736
rect 173019 79792 173085 79797
rect 173019 79736 173024 79792
rect 173080 79736 173085 79792
rect 173019 79731 173085 79736
rect 173249 79794 173315 79797
rect 173750 79794 173756 79796
rect 173249 79792 173756 79794
rect 173249 79736 173254 79792
rect 173310 79736 173756 79792
rect 173249 79734 173756 79736
rect 173249 79731 173315 79734
rect 173750 79732 173756 79734
rect 173820 79732 173826 79796
rect 172654 79661 172714 79731
rect 173022 79661 173082 79731
rect 166390 79658 166396 79660
rect 166073 79656 166396 79658
rect 166073 79600 166078 79656
rect 166134 79600 166396 79656
rect 166073 79598 166396 79600
rect 166073 79595 166139 79598
rect 166390 79596 166396 79598
rect 166460 79596 166466 79660
rect 166720 79598 166764 79660
rect 166758 79596 166764 79598
rect 166828 79596 166834 79660
rect 166950 79656 167059 79661
rect 166950 79600 166998 79656
rect 167054 79600 167059 79656
rect 166950 79598 167059 79600
rect 166993 79595 167059 79598
rect 167678 79596 167684 79660
rect 167748 79658 167754 79660
rect 167913 79658 167979 79661
rect 167748 79656 167979 79658
rect 167748 79600 167918 79656
rect 167974 79600 167979 79656
rect 167748 79598 167979 79600
rect 168054 79656 168163 79661
rect 168054 79600 168102 79656
rect 168158 79600 168163 79656
rect 168054 79598 168163 79600
rect 167748 79596 167754 79598
rect 167913 79595 167979 79598
rect 168097 79595 168163 79598
rect 168373 79656 168482 79661
rect 168373 79600 168378 79656
rect 168434 79600 168482 79656
rect 168373 79598 168482 79600
rect 170029 79656 170095 79661
rect 170029 79600 170034 79656
rect 170090 79600 170095 79656
rect 168373 79595 168439 79598
rect 170029 79595 170095 79600
rect 170262 79656 170371 79661
rect 170262 79600 170310 79656
rect 170366 79600 170371 79656
rect 170262 79598 170371 79600
rect 170305 79595 170371 79598
rect 170949 79660 171015 79661
rect 170949 79656 170996 79660
rect 171060 79658 171066 79660
rect 170949 79600 170954 79656
rect 170949 79596 170996 79600
rect 171060 79598 171106 79658
rect 171060 79596 171066 79598
rect 172094 79596 172100 79660
rect 172164 79658 172170 79660
rect 172421 79658 172487 79661
rect 172164 79656 172487 79658
rect 172164 79600 172426 79656
rect 172482 79600 172487 79656
rect 172164 79598 172487 79600
rect 172654 79656 172763 79661
rect 172654 79600 172702 79656
rect 172758 79600 172763 79656
rect 172654 79598 172763 79600
rect 173022 79656 173131 79661
rect 173022 79600 173070 79656
rect 173126 79600 173131 79656
rect 173022 79598 173131 79600
rect 172164 79596 172170 79598
rect 170949 79595 171015 79596
rect 172421 79595 172487 79598
rect 172697 79595 172763 79598
rect 173065 79595 173131 79598
rect 173249 79658 173315 79661
rect 173525 79658 173591 79661
rect 173249 79656 173591 79658
rect 173249 79600 173254 79656
rect 173310 79600 173530 79656
rect 173586 79600 173591 79656
rect 173249 79598 173591 79600
rect 173249 79595 173315 79598
rect 173525 79595 173591 79598
rect 173985 79658 174051 79661
rect 174126 79658 174186 79870
rect 174491 79867 174557 79870
rect 174537 79796 174603 79797
rect 174486 79794 174492 79796
rect 174446 79734 174492 79794
rect 174556 79792 174603 79796
rect 174598 79736 174603 79792
rect 174486 79732 174492 79734
rect 174556 79732 174603 79736
rect 174537 79731 174603 79732
rect 174678 79661 174738 79901
rect 174854 79732 174860 79796
rect 174924 79794 174930 79796
rect 175000 79794 175060 79901
rect 175319 79930 175385 79933
rect 175779 79932 175784 79962
rect 175840 79932 175845 79962
rect 176055 79962 176164 79967
rect 175319 79928 175428 79930
rect 175319 79872 175324 79928
rect 175380 79872 175428 79928
rect 175319 79867 175428 79872
rect 175774 79868 175780 79932
rect 175844 79930 175850 79932
rect 175844 79870 175902 79930
rect 176055 79906 176060 79962
rect 176116 79906 176164 79962
rect 176055 79904 176164 79906
rect 176239 79962 176305 79967
rect 176239 79906 176244 79962
rect 176300 79930 176305 79962
rect 177527 79964 177593 79967
rect 177527 79962 177636 79964
rect 176510 79930 176516 79932
rect 176300 79906 176516 79930
rect 176055 79901 176121 79904
rect 176239 79901 176516 79906
rect 176242 79870 176516 79901
rect 175844 79868 175850 79870
rect 176510 79868 176516 79870
rect 176580 79868 176586 79932
rect 176975 79930 177041 79933
rect 176975 79928 177314 79930
rect 176975 79872 176980 79928
rect 177036 79872 177314 79928
rect 177527 79906 177532 79962
rect 177588 79930 177636 79962
rect 180517 79930 180583 79933
rect 177588 79928 180583 79930
rect 177588 79906 180522 79928
rect 177527 79901 180522 79906
rect 176975 79870 177314 79872
rect 177576 79872 180522 79901
rect 180578 79872 180583 79928
rect 177576 79870 180583 79872
rect 176975 79867 177041 79870
rect 174924 79734 175060 79794
rect 175368 79794 175428 79867
rect 177021 79794 177087 79797
rect 177254 79794 177314 79870
rect 180517 79867 180583 79870
rect 185342 79868 185348 79932
rect 185412 79930 185418 79932
rect 187325 79930 187391 79933
rect 185412 79928 187391 79930
rect 185412 79872 187330 79928
rect 187386 79872 187391 79928
rect 185412 79870 187391 79872
rect 185412 79868 185418 79870
rect 187325 79867 187391 79870
rect 175368 79734 175980 79794
rect 174924 79732 174930 79734
rect 173985 79656 174186 79658
rect 173985 79600 173990 79656
rect 174046 79600 174186 79656
rect 173985 79598 174186 79600
rect 174629 79656 174738 79661
rect 174629 79600 174634 79656
rect 174690 79600 174738 79656
rect 174629 79598 174738 79600
rect 173985 79595 174051 79598
rect 174629 79595 174695 79598
rect 174854 79596 174860 79660
rect 174924 79658 174930 79660
rect 175181 79658 175247 79661
rect 174924 79656 175247 79658
rect 174924 79600 175186 79656
rect 175242 79600 175247 79656
rect 174924 79598 175247 79600
rect 174924 79596 174930 79598
rect 175181 79595 175247 79598
rect 175590 79596 175596 79660
rect 175660 79658 175666 79660
rect 175733 79658 175799 79661
rect 175660 79656 175799 79658
rect 175660 79600 175738 79656
rect 175794 79600 175799 79656
rect 175660 79598 175799 79600
rect 175920 79660 175980 79734
rect 177021 79792 177314 79794
rect 177021 79736 177026 79792
rect 177082 79736 177314 79792
rect 177021 79734 177314 79736
rect 177021 79731 177087 79734
rect 175920 79598 175964 79660
rect 175660 79596 175666 79598
rect 175733 79595 175799 79598
rect 175958 79596 175964 79598
rect 176028 79658 176034 79660
rect 179505 79658 179571 79661
rect 176028 79656 179571 79658
rect 176028 79600 179510 79656
rect 179566 79600 179571 79656
rect 176028 79598 179571 79600
rect 176028 79596 176034 79598
rect 179505 79595 179571 79598
rect 185342 79596 185348 79660
rect 185412 79658 185418 79660
rect 189533 79658 189599 79661
rect 185412 79656 189599 79658
rect 185412 79600 189538 79656
rect 189594 79600 189599 79656
rect 185412 79598 189599 79600
rect 185412 79596 185418 79598
rect 189533 79595 189599 79598
rect 153948 79462 154314 79522
rect 154849 79522 154915 79525
rect 288433 79522 288499 79525
rect 154849 79520 288499 79522
rect 154849 79464 154854 79520
rect 154910 79464 288438 79520
rect 288494 79464 288499 79520
rect 154849 79462 288499 79464
rect 153948 79460 153954 79462
rect 154849 79459 154915 79462
rect 288433 79459 288499 79462
rect 126237 79386 126303 79389
rect 136173 79386 136239 79389
rect 126237 79384 136239 79386
rect 126237 79328 126242 79384
rect 126298 79328 136178 79384
rect 136234 79328 136239 79384
rect 126237 79326 136239 79328
rect 126237 79323 126303 79326
rect 136173 79323 136239 79326
rect 148726 79324 148732 79388
rect 148796 79386 148802 79388
rect 148869 79386 148935 79389
rect 148796 79384 148935 79386
rect 148796 79328 148874 79384
rect 148930 79328 148935 79384
rect 148796 79326 148935 79328
rect 148796 79324 148802 79326
rect 148869 79323 148935 79326
rect 149094 79324 149100 79388
rect 149164 79386 149170 79388
rect 149605 79386 149671 79389
rect 149164 79384 149671 79386
rect 149164 79328 149610 79384
rect 149666 79328 149671 79384
rect 149164 79326 149671 79328
rect 149164 79324 149170 79326
rect 149605 79323 149671 79326
rect 165705 79384 165771 79389
rect 165705 79328 165710 79384
rect 165766 79328 165771 79384
rect 165705 79323 165771 79328
rect 165981 79386 166047 79389
rect 167085 79386 167151 79389
rect 165981 79384 167151 79386
rect 165981 79328 165986 79384
rect 166042 79328 167090 79384
rect 167146 79328 167151 79384
rect 165981 79326 167151 79328
rect 165981 79323 166047 79326
rect 167085 79323 167151 79326
rect 167453 79386 167519 79389
rect 168649 79386 168715 79389
rect 167453 79384 168715 79386
rect 167453 79328 167458 79384
rect 167514 79328 168654 79384
rect 168710 79328 168715 79384
rect 167453 79326 168715 79328
rect 167453 79323 167519 79326
rect 168649 79323 168715 79326
rect 169753 79386 169819 79389
rect 170622 79386 170628 79388
rect 169753 79384 170628 79386
rect 169753 79328 169758 79384
rect 169814 79328 170628 79384
rect 169753 79326 170628 79328
rect 169753 79323 169819 79326
rect 170622 79324 170628 79326
rect 170692 79324 170698 79388
rect 171133 79386 171199 79389
rect 171910 79386 171916 79388
rect 171133 79384 171916 79386
rect 171133 79328 171138 79384
rect 171194 79328 171916 79384
rect 171133 79326 171916 79328
rect 171133 79323 171199 79326
rect 171910 79324 171916 79326
rect 171980 79324 171986 79388
rect 173341 79386 173407 79389
rect 175038 79386 175044 79388
rect 173341 79384 175044 79386
rect 173341 79328 173346 79384
rect 173402 79328 175044 79384
rect 173341 79326 175044 79328
rect 173341 79323 173407 79326
rect 175038 79324 175044 79326
rect 175108 79324 175114 79388
rect 176653 79386 176719 79389
rect 193806 79386 193812 79388
rect 176653 79384 193812 79386
rect 176653 79328 176658 79384
rect 176714 79328 193812 79384
rect 176653 79326 193812 79328
rect 176653 79323 176719 79326
rect 193806 79324 193812 79326
rect 193876 79324 193882 79388
rect 118969 79250 119035 79253
rect 150525 79250 150591 79253
rect 151077 79250 151143 79253
rect 118969 79248 151143 79250
rect 118969 79192 118974 79248
rect 119030 79192 150530 79248
rect 150586 79192 151082 79248
rect 151138 79192 151143 79248
rect 118969 79190 151143 79192
rect 118969 79187 119035 79190
rect 150525 79187 150591 79190
rect 151077 79187 151143 79190
rect 152549 79250 152615 79253
rect 152774 79250 152780 79252
rect 152549 79248 152780 79250
rect 152549 79192 152554 79248
rect 152610 79192 152780 79248
rect 152549 79190 152780 79192
rect 152549 79187 152615 79190
rect 152774 79188 152780 79190
rect 152844 79188 152850 79252
rect 119337 79114 119403 79117
rect 150893 79114 150959 79117
rect 119337 79112 150959 79114
rect 119337 79056 119342 79112
rect 119398 79056 150898 79112
rect 150954 79056 150959 79112
rect 119337 79054 150959 79056
rect 119337 79051 119403 79054
rect 150893 79051 150959 79054
rect 120942 78916 120948 78980
rect 121012 78978 121018 78980
rect 154849 78978 154915 78981
rect 121012 78976 154915 78978
rect 121012 78920 154854 78976
rect 154910 78920 154915 78976
rect 121012 78918 154915 78920
rect 121012 78916 121018 78918
rect 154849 78915 154915 78918
rect 158110 78916 158116 78980
rect 158180 78978 158186 78980
rect 158805 78978 158871 78981
rect 158180 78976 158871 78978
rect 158180 78920 158810 78976
rect 158866 78920 158871 78976
rect 158180 78918 158871 78920
rect 158180 78916 158186 78918
rect 158805 78915 158871 78918
rect 164325 78978 164391 78981
rect 165708 78978 165768 79323
rect 166901 79250 166967 79253
rect 186998 79250 187004 79252
rect 166901 79248 187004 79250
rect 166901 79192 166906 79248
rect 166962 79192 187004 79248
rect 166901 79190 187004 79192
rect 166901 79187 166967 79190
rect 186998 79188 187004 79190
rect 187068 79188 187074 79252
rect 169385 79114 169451 79117
rect 191046 79114 191052 79116
rect 169385 79112 191052 79114
rect 169385 79056 169390 79112
rect 169446 79056 191052 79112
rect 169385 79054 191052 79056
rect 169385 79051 169451 79054
rect 191046 79052 191052 79054
rect 191116 79052 191122 79116
rect 187918 78978 187924 78980
rect 164325 78976 187924 78978
rect 164325 78920 164330 78976
rect 164386 78920 187924 78976
rect 164325 78918 187924 78920
rect 164325 78915 164391 78918
rect 187918 78916 187924 78918
rect 187988 78916 187994 78980
rect 100293 78842 100359 78845
rect 134149 78842 134215 78845
rect 153653 78842 153719 78845
rect 274633 78842 274699 78845
rect 100293 78840 134215 78842
rect 100293 78784 100298 78840
rect 100354 78784 134154 78840
rect 134210 78784 134215 78840
rect 100293 78782 134215 78784
rect 100293 78779 100359 78782
rect 134149 78779 134215 78782
rect 140730 78840 274699 78842
rect 140730 78784 153658 78840
rect 153714 78784 274638 78840
rect 274694 78784 274699 78840
rect 140730 78782 274699 78784
rect 119470 78644 119476 78708
rect 119540 78706 119546 78708
rect 140730 78706 140790 78782
rect 153653 78779 153719 78782
rect 274633 78779 274699 78782
rect 142613 78708 142679 78709
rect 142613 78706 142660 78708
rect 119540 78646 140790 78706
rect 142568 78704 142660 78706
rect 142568 78648 142618 78704
rect 142568 78646 142660 78648
rect 119540 78644 119546 78646
rect 142613 78644 142660 78646
rect 142724 78644 142730 78708
rect 146886 78644 146892 78708
rect 146956 78706 146962 78708
rect 147029 78706 147095 78709
rect 146956 78704 147095 78706
rect 146956 78648 147034 78704
rect 147090 78648 147095 78704
rect 146956 78646 147095 78648
rect 146956 78644 146962 78646
rect 142613 78643 142679 78644
rect 147029 78643 147095 78646
rect 151721 78706 151787 78709
rect 152406 78706 152412 78708
rect 151721 78704 152412 78706
rect 151721 78648 151726 78704
rect 151782 78648 152412 78704
rect 151721 78646 152412 78648
rect 151721 78643 151787 78646
rect 152406 78644 152412 78646
rect 152476 78644 152482 78708
rect 159173 78706 159239 78709
rect 160645 78708 160711 78709
rect 160921 78708 160987 78709
rect 159398 78706 159404 78708
rect 159173 78704 159404 78706
rect 159173 78648 159178 78704
rect 159234 78648 159404 78704
rect 159173 78646 159404 78648
rect 159173 78643 159239 78646
rect 159398 78644 159404 78646
rect 159468 78644 159474 78708
rect 160645 78706 160692 78708
rect 160600 78704 160692 78706
rect 160600 78648 160650 78704
rect 160600 78646 160692 78648
rect 160645 78644 160692 78646
rect 160756 78644 160762 78708
rect 160870 78706 160876 78708
rect 160830 78646 160876 78706
rect 160940 78704 160987 78708
rect 160982 78648 160987 78704
rect 160870 78644 160876 78646
rect 160940 78644 160987 78648
rect 160645 78643 160711 78644
rect 160921 78643 160987 78644
rect 170489 78706 170555 78709
rect 171726 78706 171732 78708
rect 170489 78704 171732 78706
rect 170489 78648 170494 78704
rect 170550 78648 171732 78704
rect 170489 78646 171732 78648
rect 170489 78643 170555 78646
rect 171726 78644 171732 78646
rect 171796 78644 171802 78708
rect 171910 78644 171916 78708
rect 171980 78706 171986 78708
rect 172145 78706 172211 78709
rect 171980 78704 172211 78706
rect 171980 78648 172150 78704
rect 172206 78648 172211 78704
rect 171980 78646 172211 78648
rect 171980 78644 171986 78646
rect 172145 78643 172211 78646
rect 175917 78706 175983 78709
rect 187366 78706 187372 78708
rect 175917 78704 187372 78706
rect 175917 78648 175922 78704
rect 175978 78648 187372 78704
rect 175917 78646 187372 78648
rect 175917 78643 175983 78646
rect 187366 78644 187372 78646
rect 187436 78644 187442 78708
rect 119838 78508 119844 78572
rect 119908 78570 119914 78572
rect 132033 78570 132099 78573
rect 119908 78568 132099 78570
rect 119908 78512 132038 78568
rect 132094 78512 132099 78568
rect 119908 78510 132099 78512
rect 119908 78508 119914 78510
rect 132033 78507 132099 78510
rect 149278 78508 149284 78572
rect 149348 78570 149354 78572
rect 149513 78570 149579 78573
rect 149348 78568 149579 78570
rect 149348 78512 149518 78568
rect 149574 78512 149579 78568
rect 149348 78510 149579 78512
rect 149348 78508 149354 78510
rect 149513 78507 149579 78510
rect 156505 78570 156571 78573
rect 157006 78570 157012 78572
rect 156505 78568 157012 78570
rect 156505 78512 156510 78568
rect 156566 78512 157012 78568
rect 156505 78510 157012 78512
rect 156505 78507 156571 78510
rect 157006 78508 157012 78510
rect 157076 78508 157082 78572
rect 158846 78508 158852 78572
rect 158916 78570 158922 78572
rect 159541 78570 159607 78573
rect 158916 78568 159607 78570
rect 158916 78512 159546 78568
rect 159602 78512 159607 78568
rect 158916 78510 159607 78512
rect 158916 78508 158922 78510
rect 159541 78507 159607 78510
rect 170029 78570 170095 78573
rect 170622 78570 170628 78572
rect 170029 78568 170628 78570
rect 170029 78512 170034 78568
rect 170090 78512 170628 78568
rect 170029 78510 170628 78512
rect 170029 78507 170095 78510
rect 170622 78508 170628 78510
rect 170692 78508 170698 78572
rect 122649 78434 122715 78437
rect 128997 78434 129063 78437
rect 131665 78434 131731 78437
rect 122649 78432 131731 78434
rect 122649 78376 122654 78432
rect 122710 78376 129002 78432
rect 129058 78376 131670 78432
rect 131726 78376 131731 78432
rect 122649 78374 131731 78376
rect 122649 78371 122715 78374
rect 128997 78371 129063 78374
rect 131665 78371 131731 78374
rect 132309 78434 132375 78437
rect 141550 78434 141556 78436
rect 132309 78432 141556 78434
rect 132309 78376 132314 78432
rect 132370 78376 141556 78432
rect 132309 78374 141556 78376
rect 132309 78371 132375 78374
rect 141550 78372 141556 78374
rect 141620 78372 141626 78436
rect 175273 78434 175339 78437
rect 175590 78434 175596 78436
rect 175273 78432 175596 78434
rect 175273 78376 175278 78432
rect 175334 78376 175596 78432
rect 175273 78374 175596 78376
rect 175273 78371 175339 78374
rect 175590 78372 175596 78374
rect 175660 78372 175666 78436
rect 180517 78434 180583 78437
rect 211286 78434 211292 78436
rect 180517 78432 211292 78434
rect 180517 78376 180522 78432
rect 180578 78376 211292 78432
rect 180517 78374 211292 78376
rect 180517 78371 180583 78374
rect 211286 78372 211292 78374
rect 211356 78434 211362 78436
rect 211356 78374 213562 78434
rect 211356 78372 211362 78374
rect 105261 78298 105327 78301
rect 123477 78298 123543 78301
rect 103470 78296 123543 78298
rect 103470 78240 105266 78296
rect 105322 78240 123482 78296
rect 123538 78240 123543 78296
rect 103470 78238 123543 78240
rect 20713 78162 20779 78165
rect 102174 78162 102180 78164
rect 20713 78160 102180 78162
rect 20713 78104 20718 78160
rect 20774 78104 102180 78160
rect 20713 78102 102180 78104
rect 20713 78099 20779 78102
rect 102174 78100 102180 78102
rect 102244 78100 102250 78164
rect 6913 78026 6979 78029
rect 103470 78026 103530 78238
rect 105261 78235 105327 78238
rect 123477 78235 123543 78238
rect 161473 78298 161539 78301
rect 162342 78298 162348 78300
rect 161473 78296 162348 78298
rect 161473 78240 161478 78296
rect 161534 78240 162348 78296
rect 161473 78238 162348 78240
rect 161473 78235 161539 78238
rect 162342 78236 162348 78238
rect 162412 78236 162418 78300
rect 173709 78298 173775 78301
rect 175038 78298 175044 78300
rect 173709 78296 175044 78298
rect 173709 78240 173714 78296
rect 173770 78240 175044 78296
rect 173709 78238 175044 78240
rect 173709 78235 173775 78238
rect 175038 78236 175044 78238
rect 175108 78236 175114 78300
rect 176142 78236 176148 78300
rect 176212 78298 176218 78300
rect 176377 78298 176443 78301
rect 176212 78296 176443 78298
rect 176212 78240 176382 78296
rect 176438 78240 176443 78296
rect 176212 78238 176443 78240
rect 176212 78236 176218 78238
rect 176377 78235 176443 78238
rect 177481 78298 177547 78301
rect 177481 78296 186330 78298
rect 177481 78240 177486 78296
rect 177542 78240 186330 78296
rect 177481 78238 186330 78240
rect 177481 78235 177547 78238
rect 124857 78162 124923 78165
rect 142337 78162 142403 78165
rect 124857 78160 142403 78162
rect 124857 78104 124862 78160
rect 124918 78104 142342 78160
rect 142398 78104 142403 78160
rect 124857 78102 142403 78104
rect 124857 78099 124923 78102
rect 142337 78099 142403 78102
rect 154982 78100 154988 78164
rect 155052 78162 155058 78164
rect 158069 78162 158135 78165
rect 155052 78160 158135 78162
rect 155052 78104 158074 78160
rect 158130 78104 158135 78160
rect 155052 78102 158135 78104
rect 155052 78100 155058 78102
rect 158069 78099 158135 78102
rect 173198 78100 173204 78164
rect 173268 78162 173274 78164
rect 173709 78162 173775 78165
rect 173268 78160 173775 78162
rect 173268 78104 173714 78160
rect 173770 78104 173775 78160
rect 173268 78102 173775 78104
rect 186270 78162 186330 78238
rect 190678 78236 190684 78300
rect 190748 78298 190754 78300
rect 190821 78298 190887 78301
rect 190748 78296 190887 78298
rect 190748 78240 190826 78296
rect 190882 78240 190887 78296
rect 190748 78238 190887 78240
rect 190748 78236 190754 78238
rect 190821 78235 190887 78238
rect 211102 78162 211108 78164
rect 186270 78102 211108 78162
rect 173268 78100 173274 78102
rect 173709 78099 173775 78102
rect 211102 78100 211108 78102
rect 211172 78162 211178 78164
rect 211172 78102 213378 78162
rect 211172 78100 211178 78102
rect 6913 78024 103530 78026
rect 6913 77968 6918 78024
rect 6974 77968 103530 78024
rect 6913 77966 103530 77968
rect 6913 77963 6979 77966
rect 134374 77964 134380 78028
rect 134444 78026 134450 78028
rect 134517 78026 134583 78029
rect 134444 78024 134583 78026
rect 134444 77968 134522 78024
rect 134578 77968 134583 78024
rect 134444 77966 134583 77968
rect 134444 77964 134450 77966
rect 134517 77963 134583 77966
rect 163078 77964 163084 78028
rect 163148 78026 163154 78028
rect 163221 78026 163287 78029
rect 163148 78024 163287 78026
rect 163148 77968 163226 78024
rect 163282 77968 163287 78024
rect 163148 77966 163287 77968
rect 163148 77964 163154 77966
rect 163221 77963 163287 77966
rect 167310 77964 167316 78028
rect 167380 78026 167386 78028
rect 167862 78026 167868 78028
rect 167380 77966 167868 78026
rect 167380 77964 167386 77966
rect 167862 77964 167868 77966
rect 167932 77964 167938 78028
rect 171409 78026 171475 78029
rect 178769 78026 178835 78029
rect 178902 78026 178908 78028
rect 171409 78024 176578 78026
rect 171409 77968 171414 78024
rect 171470 77968 176578 78024
rect 171409 77966 176578 77968
rect 171409 77963 171475 77966
rect 2773 77890 2839 77893
rect 134517 77890 134583 77893
rect 142061 77890 142127 77893
rect 2773 77888 103530 77890
rect 2773 77832 2778 77888
rect 2834 77832 103530 77888
rect 2773 77830 103530 77832
rect 2773 77827 2839 77830
rect 103470 77482 103530 77830
rect 134517 77888 142127 77890
rect 134517 77832 134522 77888
rect 134578 77832 142066 77888
rect 142122 77832 142127 77888
rect 134517 77830 142127 77832
rect 134517 77827 134583 77830
rect 142061 77827 142127 77830
rect 143942 77828 143948 77892
rect 144012 77890 144018 77892
rect 144453 77890 144519 77893
rect 144012 77888 144519 77890
rect 144012 77832 144458 77888
rect 144514 77832 144519 77888
rect 144012 77830 144519 77832
rect 144012 77828 144018 77830
rect 144453 77827 144519 77830
rect 163313 77890 163379 77893
rect 163446 77890 163452 77892
rect 163313 77888 163452 77890
rect 163313 77832 163318 77888
rect 163374 77832 163452 77888
rect 163313 77830 163452 77832
rect 163313 77827 163379 77830
rect 163446 77828 163452 77830
rect 163516 77828 163522 77892
rect 163630 77828 163636 77892
rect 163700 77890 163706 77892
rect 164141 77890 164207 77893
rect 163700 77888 164207 77890
rect 163700 77832 164146 77888
rect 164202 77832 164207 77888
rect 163700 77830 164207 77832
rect 176518 77890 176578 77966
rect 178769 78024 178908 78026
rect 178769 77968 178774 78024
rect 178830 77968 178908 78024
rect 178769 77966 178908 77968
rect 178769 77963 178835 77966
rect 178902 77964 178908 77966
rect 178972 77964 178978 78028
rect 179505 78026 179571 78029
rect 206369 78026 206435 78029
rect 179505 78024 206435 78026
rect 179505 77968 179510 78024
rect 179566 77968 206374 78024
rect 206430 77968 206435 78024
rect 179505 77966 206435 77968
rect 179505 77963 179571 77966
rect 206369 77963 206435 77966
rect 181621 77890 181687 77893
rect 182081 77890 182147 77893
rect 210601 77890 210667 77893
rect 176518 77830 181546 77890
rect 163700 77828 163706 77830
rect 164141 77827 164207 77830
rect 143574 77692 143580 77756
rect 143644 77754 143650 77756
rect 144453 77754 144519 77757
rect 143644 77752 144519 77754
rect 143644 77696 144458 77752
rect 144514 77696 144519 77752
rect 143644 77694 144519 77696
rect 143644 77692 143650 77694
rect 144453 77691 144519 77694
rect 163446 77692 163452 77756
rect 163516 77754 163522 77756
rect 163865 77754 163931 77757
rect 163516 77752 163931 77754
rect 163516 77696 163870 77752
rect 163926 77696 163931 77752
rect 163516 77694 163931 77696
rect 181486 77754 181546 77830
rect 181621 77888 210667 77890
rect 181621 77832 181626 77888
rect 181682 77832 182086 77888
rect 182142 77832 210606 77888
rect 210662 77832 210667 77888
rect 181621 77830 210667 77832
rect 213318 77890 213378 78102
rect 213502 78026 213562 78374
rect 213821 78162 213887 78165
rect 500953 78162 501019 78165
rect 213821 78160 501019 78162
rect 213821 78104 213826 78160
rect 213882 78104 500958 78160
rect 501014 78104 501019 78160
rect 213821 78102 501019 78104
rect 213821 78099 213887 78102
rect 500953 78099 501019 78102
rect 581085 78026 581151 78029
rect 213502 78024 581151 78026
rect 213502 77968 581090 78024
rect 581146 77968 581151 78024
rect 213502 77966 581151 77968
rect 581085 77963 581151 77966
rect 580993 77890 581059 77893
rect 213318 77888 581059 77890
rect 213318 77832 580998 77888
rect 581054 77832 581059 77888
rect 213318 77830 581059 77832
rect 181621 77827 181687 77830
rect 182081 77827 182147 77830
rect 210601 77827 210667 77830
rect 580993 77827 581059 77830
rect 181486 77694 186330 77754
rect 163516 77692 163522 77694
rect 163865 77691 163931 77694
rect 121453 77618 121519 77621
rect 130837 77618 130903 77621
rect 144177 77618 144243 77621
rect 121453 77616 144243 77618
rect 121453 77560 121458 77616
rect 121514 77560 130842 77616
rect 130898 77560 144182 77616
rect 144238 77560 144243 77616
rect 121453 77558 144243 77560
rect 121453 77555 121519 77558
rect 130837 77555 130903 77558
rect 144177 77555 144243 77558
rect 175958 77556 175964 77620
rect 176028 77618 176034 77620
rect 176101 77618 176167 77621
rect 176028 77616 176167 77618
rect 176028 77560 176106 77616
rect 176162 77560 176167 77616
rect 176028 77558 176167 77560
rect 186270 77618 186330 77694
rect 212993 77618 213059 77621
rect 213821 77618 213887 77621
rect 186270 77616 213887 77618
rect 186270 77560 212998 77616
rect 213054 77560 213826 77616
rect 213882 77560 213887 77616
rect 186270 77558 213887 77560
rect 176028 77556 176034 77558
rect 176101 77555 176167 77558
rect 212993 77555 213059 77558
rect 213821 77555 213887 77558
rect 107326 77482 107332 77484
rect 103470 77422 107332 77482
rect 107326 77420 107332 77422
rect 107396 77482 107402 77484
rect 126053 77482 126119 77485
rect 107396 77480 126119 77482
rect 107396 77424 126058 77480
rect 126114 77424 126119 77480
rect 107396 77422 126119 77424
rect 107396 77420 107402 77422
rect 126053 77419 126119 77422
rect 141233 77482 141299 77485
rect 142102 77482 142108 77484
rect 141233 77480 142108 77482
rect 141233 77424 141238 77480
rect 141294 77424 142108 77480
rect 141233 77422 142108 77424
rect 141233 77419 141299 77422
rect 142102 77420 142108 77422
rect 142172 77420 142178 77484
rect 148409 77482 148475 77485
rect 148910 77482 148916 77484
rect 148409 77480 148916 77482
rect 148409 77424 148414 77480
rect 148470 77424 148916 77480
rect 148409 77422 148916 77424
rect 148409 77419 148475 77422
rect 148910 77420 148916 77422
rect 148980 77420 148986 77484
rect 153837 77482 153903 77485
rect 175733 77484 175799 77485
rect 154430 77482 154436 77484
rect 153837 77480 154436 77482
rect 153837 77424 153842 77480
rect 153898 77424 154436 77480
rect 153837 77422 154436 77424
rect 153837 77419 153903 77422
rect 154430 77420 154436 77422
rect 154500 77420 154506 77484
rect 175733 77482 175780 77484
rect 175688 77480 175780 77482
rect 175688 77424 175738 77480
rect 175688 77422 175780 77424
rect 175733 77420 175780 77422
rect 175844 77420 175850 77484
rect 176377 77482 176443 77485
rect 210141 77482 210207 77485
rect 176377 77480 210207 77482
rect 176377 77424 176382 77480
rect 176438 77424 210146 77480
rect 210202 77424 210207 77480
rect 176377 77422 210207 77424
rect 175733 77419 175799 77420
rect 176377 77419 176443 77422
rect 210141 77419 210207 77422
rect 102174 77284 102180 77348
rect 102244 77346 102250 77348
rect 103278 77346 103284 77348
rect 102244 77286 103284 77346
rect 102244 77284 102250 77286
rect 103278 77284 103284 77286
rect 103348 77346 103354 77348
rect 133873 77346 133939 77349
rect 103348 77344 133939 77346
rect 103348 77288 133878 77344
rect 133934 77288 133939 77344
rect 103348 77286 133939 77288
rect 103348 77284 103354 77286
rect 133873 77283 133939 77286
rect 147806 77284 147812 77348
rect 147876 77346 147882 77348
rect 148593 77346 148659 77349
rect 147876 77344 148659 77346
rect 147876 77288 148598 77344
rect 148654 77288 148659 77344
rect 147876 77286 148659 77288
rect 147876 77284 147882 77286
rect 148593 77283 148659 77286
rect 150014 77284 150020 77348
rect 150084 77346 150090 77348
rect 150249 77346 150315 77349
rect 150084 77344 150315 77346
rect 150084 77288 150254 77344
rect 150310 77288 150315 77344
rect 150084 77286 150315 77288
rect 150084 77284 150090 77286
rect 150249 77283 150315 77286
rect 150801 77346 150867 77349
rect 151118 77346 151124 77348
rect 150801 77344 151124 77346
rect 150801 77288 150806 77344
rect 150862 77288 151124 77344
rect 150801 77286 151124 77288
rect 150801 77283 150867 77286
rect 151118 77284 151124 77286
rect 151188 77284 151194 77348
rect 152590 77284 152596 77348
rect 152660 77346 152666 77348
rect 152660 77286 153210 77346
rect 152660 77284 152666 77286
rect 99833 77210 99899 77213
rect 133505 77210 133571 77213
rect 99833 77208 133571 77210
rect 99833 77152 99838 77208
rect 99894 77152 133510 77208
rect 133566 77152 133571 77208
rect 99833 77150 133571 77152
rect 99833 77147 99899 77150
rect 133505 77147 133571 77150
rect 148358 77148 148364 77212
rect 148428 77210 148434 77212
rect 148961 77210 149027 77213
rect 148428 77208 149027 77210
rect 148428 77152 148966 77208
rect 149022 77152 149027 77208
rect 148428 77150 149027 77152
rect 153150 77210 153210 77286
rect 154062 77284 154068 77348
rect 154132 77346 154138 77348
rect 154481 77346 154547 77349
rect 154132 77344 154547 77346
rect 154132 77288 154486 77344
rect 154542 77288 154547 77344
rect 154132 77286 154547 77288
rect 154132 77284 154138 77286
rect 154481 77283 154547 77286
rect 155534 77284 155540 77348
rect 155604 77346 155610 77348
rect 155861 77346 155927 77349
rect 162485 77348 162551 77349
rect 155604 77344 155927 77346
rect 155604 77288 155866 77344
rect 155922 77288 155927 77344
rect 155604 77286 155927 77288
rect 155604 77284 155610 77286
rect 155861 77283 155927 77286
rect 161974 77284 161980 77348
rect 162044 77346 162050 77348
rect 162342 77346 162348 77348
rect 162044 77286 162348 77346
rect 162044 77284 162050 77286
rect 162342 77284 162348 77286
rect 162412 77284 162418 77348
rect 162485 77344 162532 77348
rect 162596 77346 162602 77348
rect 162485 77288 162490 77344
rect 162485 77284 162532 77288
rect 162596 77286 162642 77346
rect 162596 77284 162602 77286
rect 162894 77284 162900 77348
rect 162964 77346 162970 77348
rect 163497 77346 163563 77349
rect 162964 77344 163563 77346
rect 162964 77288 163502 77344
rect 163558 77288 163563 77344
rect 162964 77286 163563 77288
rect 162964 77284 162970 77286
rect 162485 77283 162551 77284
rect 163497 77283 163563 77286
rect 163681 77346 163747 77349
rect 164734 77346 164740 77348
rect 163681 77344 164740 77346
rect 163681 77288 163686 77344
rect 163742 77288 164740 77344
rect 163681 77286 164740 77288
rect 163681 77283 163747 77286
rect 164734 77284 164740 77286
rect 164804 77284 164810 77348
rect 167177 77346 167243 77349
rect 167494 77346 167500 77348
rect 167177 77344 167500 77346
rect 167177 77288 167182 77344
rect 167238 77288 167500 77344
rect 167177 77286 167500 77288
rect 167177 77283 167243 77286
rect 167494 77284 167500 77286
rect 167564 77284 167570 77348
rect 175641 77346 175707 77349
rect 175958 77346 175964 77348
rect 175641 77344 175964 77346
rect 175641 77288 175646 77344
rect 175702 77288 175964 77344
rect 175641 77286 175964 77288
rect 175641 77283 175707 77286
rect 175958 77284 175964 77286
rect 176028 77284 176034 77348
rect 214189 77210 214255 77213
rect 153150 77208 219450 77210
rect 153150 77152 214194 77208
rect 214250 77152 219450 77208
rect 153150 77150 219450 77152
rect 148428 77148 148434 77150
rect 148961 77147 149027 77150
rect 214189 77147 214255 77150
rect 101489 77074 101555 77077
rect 134977 77074 135043 77077
rect 84150 77072 135043 77074
rect 84150 77016 101494 77072
rect 101550 77016 134982 77072
rect 135038 77016 135043 77072
rect 84150 77014 135043 77016
rect 34513 76530 34579 76533
rect 84150 76530 84210 77014
rect 101489 77011 101555 77014
rect 134977 77011 135043 77014
rect 135294 77012 135300 77076
rect 135364 77074 135370 77076
rect 135897 77074 135963 77077
rect 135364 77072 135963 77074
rect 135364 77016 135902 77072
rect 135958 77016 135963 77072
rect 135364 77014 135963 77016
rect 135364 77012 135370 77014
rect 135897 77011 135963 77014
rect 138054 77012 138060 77076
rect 138124 77074 138130 77076
rect 138606 77074 138612 77076
rect 138124 77014 138612 77074
rect 138124 77012 138130 77014
rect 138606 77012 138612 77014
rect 138676 77012 138682 77076
rect 176469 77074 176535 77077
rect 210325 77074 210391 77077
rect 176469 77072 213194 77074
rect 176469 77016 176474 77072
rect 176530 77016 210330 77072
rect 210386 77016 213194 77072
rect 176469 77014 213194 77016
rect 176469 77011 176535 77014
rect 210325 77011 210391 77014
rect 118325 76938 118391 76941
rect 145833 76938 145899 76941
rect 118325 76936 145899 76938
rect 118325 76880 118330 76936
rect 118386 76880 145838 76936
rect 145894 76880 145899 76936
rect 118325 76878 145899 76880
rect 118325 76875 118391 76878
rect 145833 76875 145899 76878
rect 154665 76938 154731 76941
rect 155902 76938 155908 76940
rect 154665 76936 155908 76938
rect 154665 76880 154670 76936
rect 154726 76880 155908 76936
rect 154665 76878 155908 76880
rect 154665 76875 154731 76878
rect 155902 76876 155908 76878
rect 155972 76876 155978 76940
rect 173709 76938 173775 76941
rect 175917 76938 175983 76941
rect 173709 76936 175983 76938
rect 173709 76880 173714 76936
rect 173770 76880 175922 76936
rect 175978 76880 175983 76936
rect 173709 76878 175983 76880
rect 173709 76875 173775 76878
rect 175917 76875 175983 76878
rect 177849 76938 177915 76941
rect 210233 76938 210299 76941
rect 177849 76936 210299 76938
rect 177849 76880 177854 76936
rect 177910 76880 210238 76936
rect 210294 76880 210299 76936
rect 177849 76878 210299 76880
rect 177849 76875 177915 76878
rect 210233 76875 210299 76878
rect 99373 76802 99439 76805
rect 113766 76802 113772 76804
rect 99373 76800 113772 76802
rect 99373 76744 99378 76800
rect 99434 76744 113772 76800
rect 99373 76742 113772 76744
rect 99373 76739 99439 76742
rect 113766 76740 113772 76742
rect 113836 76802 113842 76804
rect 114001 76802 114067 76805
rect 113836 76800 114067 76802
rect 113836 76744 114006 76800
rect 114062 76744 114067 76800
rect 113836 76742 114067 76744
rect 113836 76740 113842 76742
rect 114001 76739 114067 76742
rect 116945 76802 117011 76805
rect 141693 76802 141759 76805
rect 116945 76800 141759 76802
rect 116945 76744 116950 76800
rect 117006 76744 141698 76800
rect 141754 76744 141759 76800
rect 116945 76742 141759 76744
rect 116945 76739 117011 76742
rect 141693 76739 141759 76742
rect 170673 76802 170739 76805
rect 193622 76802 193628 76804
rect 170673 76800 193628 76802
rect 170673 76744 170678 76800
rect 170734 76744 193628 76800
rect 170673 76742 193628 76744
rect 170673 76739 170739 76742
rect 193622 76740 193628 76742
rect 193692 76740 193698 76804
rect 99097 76666 99163 76669
rect 131573 76666 131639 76669
rect 99097 76664 131639 76666
rect 99097 76608 99102 76664
rect 99158 76608 131578 76664
rect 131634 76608 131639 76664
rect 99097 76606 131639 76608
rect 99097 76603 99163 76606
rect 131573 76603 131639 76606
rect 132585 76666 132651 76669
rect 133454 76666 133460 76668
rect 132585 76664 133460 76666
rect 132585 76608 132590 76664
rect 132646 76608 133460 76664
rect 132585 76606 133460 76608
rect 132585 76603 132651 76606
rect 133454 76604 133460 76606
rect 133524 76604 133530 76668
rect 134057 76666 134123 76669
rect 134190 76666 134196 76668
rect 134057 76664 134196 76666
rect 134057 76608 134062 76664
rect 134118 76608 134196 76664
rect 134057 76606 134196 76608
rect 134057 76603 134123 76606
rect 134190 76604 134196 76606
rect 134260 76604 134266 76668
rect 138054 76604 138060 76668
rect 138124 76666 138130 76668
rect 139158 76666 139164 76668
rect 138124 76606 139164 76666
rect 138124 76604 138130 76606
rect 139158 76604 139164 76606
rect 139228 76604 139234 76668
rect 139342 76604 139348 76668
rect 139412 76666 139418 76668
rect 139577 76666 139643 76669
rect 139412 76664 139643 76666
rect 139412 76608 139582 76664
rect 139638 76608 139643 76664
rect 139412 76606 139643 76608
rect 139412 76604 139418 76606
rect 139577 76603 139643 76606
rect 143574 76604 143580 76668
rect 143644 76666 143650 76668
rect 144821 76666 144887 76669
rect 143644 76664 144887 76666
rect 143644 76608 144826 76664
rect 144882 76608 144887 76664
rect 143644 76606 144887 76608
rect 143644 76604 143650 76606
rect 144821 76603 144887 76606
rect 145598 76604 145604 76668
rect 145668 76666 145674 76668
rect 145833 76666 145899 76669
rect 145668 76664 145899 76666
rect 145668 76608 145838 76664
rect 145894 76608 145899 76664
rect 145668 76606 145899 76608
rect 145668 76604 145674 76606
rect 145833 76603 145899 76606
rect 146702 76604 146708 76668
rect 146772 76666 146778 76668
rect 146937 76666 147003 76669
rect 146772 76664 147003 76666
rect 146772 76608 146942 76664
rect 146998 76608 147003 76664
rect 146772 76606 147003 76608
rect 146772 76604 146778 76606
rect 146937 76603 147003 76606
rect 173525 76666 173591 76669
rect 194726 76666 194732 76668
rect 173525 76664 194732 76666
rect 173525 76608 173530 76664
rect 173586 76608 194732 76664
rect 173525 76606 194732 76608
rect 173525 76603 173591 76606
rect 194726 76604 194732 76606
rect 194796 76604 194802 76668
rect 34513 76528 84210 76530
rect 34513 76472 34518 76528
rect 34574 76472 84210 76528
rect 34513 76470 84210 76472
rect 34513 76467 34579 76470
rect 139526 76468 139532 76532
rect 139596 76530 139602 76532
rect 140262 76530 140268 76532
rect 139596 76470 140268 76530
rect 139596 76468 139602 76470
rect 140262 76468 140268 76470
rect 140332 76468 140338 76532
rect 151629 76530 151695 76533
rect 193121 76530 193187 76533
rect 209221 76530 209287 76533
rect 151629 76528 209287 76530
rect 151629 76472 151634 76528
rect 151690 76472 193126 76528
rect 193182 76472 209226 76528
rect 209282 76472 209287 76528
rect 151629 76470 209287 76472
rect 213134 76530 213194 77014
rect 219390 76666 219450 77150
rect 260097 76666 260163 76669
rect 219390 76664 260163 76666
rect 219390 76608 260102 76664
rect 260158 76608 260163 76664
rect 219390 76606 260163 76608
rect 260097 76603 260163 76606
rect 566457 76530 566523 76533
rect 213134 76528 566523 76530
rect 213134 76472 566462 76528
rect 566518 76472 566523 76528
rect 213134 76470 566523 76472
rect 151629 76467 151695 76470
rect 193121 76467 193187 76470
rect 209221 76467 209287 76470
rect 566457 76467 566523 76470
rect 173617 76394 173683 76397
rect 173934 76394 173940 76396
rect 173617 76392 173940 76394
rect 173617 76336 173622 76392
rect 173678 76336 173940 76392
rect 173617 76334 173940 76336
rect 173617 76331 173683 76334
rect 173934 76332 173940 76334
rect 174004 76332 174010 76396
rect 170489 75986 170555 75989
rect 170673 75986 170739 75989
rect 170489 75984 170739 75986
rect 170489 75928 170494 75984
rect 170550 75928 170678 75984
rect 170734 75928 170739 75984
rect 170489 75926 170739 75928
rect 170489 75923 170555 75926
rect 170673 75923 170739 75926
rect 99465 75850 99531 75853
rect 99925 75850 99991 75853
rect 135110 75850 135116 75852
rect 99465 75848 135116 75850
rect 99465 75792 99470 75848
rect 99526 75792 99930 75848
rect 99986 75792 135116 75848
rect 99465 75790 135116 75792
rect 99465 75787 99531 75790
rect 99925 75787 99991 75790
rect 135110 75788 135116 75790
rect 135180 75788 135186 75852
rect 205582 75788 205588 75852
rect 205652 75850 205658 75852
rect 206369 75850 206435 75853
rect 205652 75848 206435 75850
rect 205652 75792 206374 75848
rect 206430 75792 206435 75848
rect 205652 75790 206435 75792
rect 205652 75788 205658 75790
rect 206369 75787 206435 75790
rect 103973 75714 104039 75717
rect 137686 75714 137692 75716
rect 84150 75712 137692 75714
rect 84150 75656 103978 75712
rect 104034 75656 137692 75712
rect 84150 75654 137692 75656
rect 71037 75442 71103 75445
rect 84150 75442 84210 75654
rect 103973 75651 104039 75654
rect 137686 75652 137692 75654
rect 137756 75652 137762 75716
rect 170990 75652 170996 75716
rect 171060 75714 171066 75716
rect 171060 75654 200130 75714
rect 171060 75652 171066 75654
rect 102777 75578 102843 75581
rect 133965 75578 134031 75581
rect 102777 75576 134031 75578
rect 102777 75520 102782 75576
rect 102838 75520 133970 75576
rect 134026 75520 134031 75576
rect 102777 75518 134031 75520
rect 102777 75515 102843 75518
rect 133965 75515 134031 75518
rect 167637 75578 167703 75581
rect 191598 75578 191604 75580
rect 167637 75576 191604 75578
rect 167637 75520 167642 75576
rect 167698 75520 191604 75576
rect 167637 75518 191604 75520
rect 167637 75515 167703 75518
rect 191598 75516 191604 75518
rect 191668 75516 191674 75580
rect 71037 75440 84210 75442
rect 71037 75384 71042 75440
rect 71098 75384 84210 75440
rect 71037 75382 84210 75384
rect 167545 75442 167611 75445
rect 189758 75442 189764 75444
rect 167545 75440 189764 75442
rect 167545 75384 167550 75440
rect 167606 75384 189764 75440
rect 167545 75382 189764 75384
rect 71037 75379 71103 75382
rect 167545 75379 167611 75382
rect 189758 75380 189764 75382
rect 189828 75380 189834 75444
rect 35893 75306 35959 75309
rect 99465 75306 99531 75309
rect 35893 75304 99531 75306
rect 35893 75248 35898 75304
rect 35954 75248 99470 75304
rect 99526 75248 99531 75304
rect 35893 75246 99531 75248
rect 35893 75243 35959 75246
rect 99465 75243 99531 75246
rect 113449 75306 113515 75309
rect 129733 75306 129799 75309
rect 135621 75306 135687 75309
rect 113449 75304 135687 75306
rect 113449 75248 113454 75304
rect 113510 75248 129738 75304
rect 129794 75248 135626 75304
rect 135682 75248 135687 75304
rect 113449 75246 135687 75248
rect 113449 75243 113515 75246
rect 129733 75243 129799 75246
rect 135621 75243 135687 75246
rect 169569 75306 169635 75309
rect 178953 75306 179019 75309
rect 188286 75306 188292 75308
rect 169569 75304 188292 75306
rect 169569 75248 169574 75304
rect 169630 75248 178958 75304
rect 179014 75248 188292 75304
rect 169569 75246 188292 75248
rect 169569 75243 169635 75246
rect 178953 75243 179019 75246
rect 188286 75244 188292 75246
rect 188356 75244 188362 75308
rect 200070 75306 200130 75654
rect 204805 75306 204871 75309
rect 454677 75306 454743 75309
rect 200070 75304 454743 75306
rect 200070 75248 204810 75304
rect 204866 75248 454682 75304
rect 454738 75248 454743 75304
rect 200070 75246 454743 75248
rect 204805 75243 204871 75246
rect 454677 75243 454743 75246
rect 7557 75170 7623 75173
rect 119838 75170 119844 75172
rect 7557 75168 119844 75170
rect 7557 75112 7562 75168
rect 7618 75112 119844 75168
rect 7557 75110 119844 75112
rect 7557 75107 7623 75110
rect 119838 75108 119844 75110
rect 119908 75108 119914 75172
rect 168281 75170 168347 75173
rect 179045 75170 179111 75173
rect 189390 75170 189396 75172
rect 168281 75168 189396 75170
rect 168281 75112 168286 75168
rect 168342 75112 179050 75168
rect 179106 75112 189396 75168
rect 168281 75110 189396 75112
rect 168281 75107 168347 75110
rect 179045 75107 179111 75110
rect 189390 75108 189396 75110
rect 189460 75108 189466 75172
rect 521653 75170 521719 75173
rect 209730 75168 521719 75170
rect 209730 75112 521658 75168
rect 521714 75112 521719 75168
rect 209730 75110 521719 75112
rect 177481 75034 177547 75037
rect 207933 75034 207999 75037
rect 209730 75034 209790 75110
rect 521653 75107 521719 75110
rect 177481 75032 209790 75034
rect 177481 74976 177486 75032
rect 177542 74976 207938 75032
rect 207994 74976 209790 75032
rect 177481 74974 209790 74976
rect 177481 74971 177547 74974
rect 207933 74971 207999 74974
rect 135253 74762 135319 74765
rect 136030 74762 136036 74764
rect 135253 74760 136036 74762
rect 135253 74704 135258 74760
rect 135314 74704 136036 74760
rect 135253 74702 136036 74704
rect 135253 74699 135319 74702
rect 136030 74700 136036 74702
rect 136100 74700 136106 74764
rect 143758 74700 143764 74764
rect 143828 74762 143834 74764
rect 144637 74762 144703 74765
rect 143828 74760 144703 74762
rect 143828 74704 144642 74760
rect 144698 74704 144703 74760
rect 143828 74702 144703 74704
rect 143828 74700 143834 74702
rect 144637 74699 144703 74702
rect 133086 74564 133092 74628
rect 133156 74626 133162 74628
rect 133321 74626 133387 74629
rect 133156 74624 133387 74626
rect 133156 74568 133326 74624
rect 133382 74568 133387 74624
rect 133156 74566 133387 74568
rect 133156 74564 133162 74566
rect 133321 74563 133387 74566
rect 118366 74428 118372 74492
rect 118436 74490 118442 74492
rect 151905 74490 151971 74493
rect 153009 74490 153075 74493
rect 118436 74488 153075 74490
rect 118436 74432 151910 74488
rect 151966 74432 153014 74488
rect 153070 74432 153075 74488
rect 118436 74430 153075 74432
rect 118436 74428 118442 74430
rect 151905 74427 151971 74430
rect 153009 74427 153075 74430
rect 170213 74490 170279 74493
rect 170581 74490 170647 74493
rect 170213 74488 170647 74490
rect 170213 74432 170218 74488
rect 170274 74432 170586 74488
rect 170642 74432 170647 74488
rect 170213 74430 170647 74432
rect 170213 74427 170279 74430
rect 170581 74427 170647 74430
rect 122230 74292 122236 74356
rect 122300 74354 122306 74356
rect 155493 74354 155559 74357
rect 122300 74352 155559 74354
rect 122300 74296 155498 74352
rect 155554 74296 155559 74352
rect 122300 74294 155559 74296
rect 122300 74292 122306 74294
rect 155493 74291 155559 74294
rect 218421 74354 218487 74357
rect 237373 74354 237439 74357
rect 218421 74352 237439 74354
rect 218421 74296 218426 74352
rect 218482 74296 237378 74352
rect 237434 74296 237439 74352
rect 218421 74294 237439 74296
rect 218421 74291 218487 74294
rect 237373 74291 237439 74294
rect 115289 74218 115355 74221
rect 147070 74218 147076 74220
rect 115289 74216 147076 74218
rect 115289 74160 115294 74216
rect 115350 74160 147076 74216
rect 115289 74158 147076 74160
rect 115289 74155 115355 74158
rect 147070 74156 147076 74158
rect 147140 74156 147146 74220
rect 149646 74156 149652 74220
rect 149716 74218 149722 74220
rect 215753 74218 215819 74221
rect 149716 74216 215819 74218
rect 149716 74160 215758 74216
rect 215814 74160 215819 74216
rect 149716 74158 215819 74160
rect 149716 74156 149722 74158
rect 215753 74155 215819 74158
rect 218237 74218 218303 74221
rect 248413 74218 248479 74221
rect 218237 74216 248479 74218
rect 218237 74160 218242 74216
rect 218298 74160 248418 74216
rect 248474 74160 248479 74216
rect 218237 74158 248479 74160
rect 218237 74155 218303 74158
rect 248413 74155 248479 74158
rect 106825 74084 106891 74085
rect 106774 74082 106780 74084
rect 106734 74022 106780 74082
rect 106844 74080 106891 74084
rect 106886 74024 106891 74080
rect 106774 74020 106780 74022
rect 106844 74020 106891 74024
rect 106825 74019 106891 74020
rect 122373 74082 122439 74085
rect 149605 74082 149671 74085
rect 150341 74082 150407 74085
rect 122373 74080 150407 74082
rect 122373 74024 122378 74080
rect 122434 74024 149610 74080
rect 149666 74024 150346 74080
rect 150402 74024 150407 74080
rect 122373 74022 150407 74024
rect 122373 74019 122439 74022
rect 149605 74019 149671 74022
rect 150341 74019 150407 74022
rect 153142 74020 153148 74084
rect 153212 74082 153218 74084
rect 218329 74082 218395 74085
rect 153212 74080 219450 74082
rect 153212 74024 218334 74080
rect 218390 74024 219450 74080
rect 153212 74022 219450 74024
rect 153212 74020 153218 74022
rect 218329 74019 218395 74022
rect 113582 73884 113588 73948
rect 113652 73946 113658 73948
rect 136725 73946 136791 73949
rect 113652 73944 136791 73946
rect 113652 73888 136730 73944
rect 136786 73888 136791 73944
rect 113652 73886 136791 73888
rect 113652 73884 113658 73886
rect 136725 73883 136791 73886
rect 149462 73884 149468 73948
rect 149532 73946 149538 73948
rect 211797 73946 211863 73949
rect 149532 73944 211863 73946
rect 149532 73888 211802 73944
rect 211858 73888 211863 73944
rect 149532 73886 211863 73888
rect 219390 73946 219450 74022
rect 261477 73946 261543 73949
rect 219390 73944 261543 73946
rect 219390 73888 261482 73944
rect 261538 73888 261543 73944
rect 219390 73886 261543 73888
rect 149532 73884 149538 73886
rect 211797 73883 211863 73886
rect 261477 73883 261543 73886
rect 54477 73810 54543 73813
rect 106825 73810 106891 73813
rect 54477 73808 106891 73810
rect 54477 73752 54482 73808
rect 54538 73752 106830 73808
rect 106886 73752 106891 73808
rect 54477 73750 106891 73752
rect 54477 73747 54543 73750
rect 106825 73747 106891 73750
rect 162158 73748 162164 73812
rect 162228 73810 162234 73812
rect 216857 73810 216923 73813
rect 347773 73810 347839 73813
rect 162228 73808 347839 73810
rect 162228 73752 216862 73808
rect 216918 73752 347778 73808
rect 347834 73752 347839 73808
rect 162228 73750 347839 73752
rect 162228 73748 162234 73750
rect 216857 73747 216923 73750
rect 347773 73747 347839 73750
rect 106273 73674 106339 73677
rect 111793 73674 111859 73677
rect 112294 73674 112300 73676
rect 106273 73672 112300 73674
rect 106273 73616 106278 73672
rect 106334 73616 111798 73672
rect 111854 73616 112300 73672
rect 106273 73614 112300 73616
rect 106273 73611 106339 73614
rect 111793 73611 111859 73614
rect 112294 73612 112300 73614
rect 112364 73612 112370 73676
rect 170581 73674 170647 73677
rect 193438 73674 193444 73676
rect 170581 73672 193444 73674
rect 170581 73616 170586 73672
rect 170642 73616 193444 73672
rect 170581 73614 193444 73616
rect 170581 73611 170647 73614
rect 193438 73612 193444 73614
rect 193508 73612 193514 73676
rect 215753 73674 215819 73677
rect 224217 73674 224283 73677
rect 215753 73672 224283 73674
rect 215753 73616 215758 73672
rect 215814 73616 224222 73672
rect 224278 73616 224283 73672
rect 215753 73614 224283 73616
rect 215753 73611 215819 73614
rect 224217 73611 224283 73614
rect 151118 73476 151124 73540
rect 151188 73538 151194 73540
rect 218421 73538 218487 73541
rect 151188 73536 218487 73538
rect 151188 73480 218426 73536
rect 218482 73480 218487 73536
rect 151188 73478 218487 73480
rect 151188 73476 151194 73478
rect 218421 73475 218487 73478
rect 151670 73340 151676 73404
rect 151740 73402 151746 73404
rect 218237 73402 218303 73405
rect 151740 73400 218303 73402
rect 151740 73344 218242 73400
rect 218298 73344 218303 73400
rect 151740 73342 218303 73344
rect 151740 73340 151746 73342
rect 218237 73339 218303 73342
rect 108297 73132 108363 73133
rect 108246 73130 108252 73132
rect 108206 73070 108252 73130
rect 108316 73128 108363 73132
rect 108358 73072 108363 73128
rect 108246 73068 108252 73070
rect 108316 73068 108363 73072
rect 117078 73068 117084 73132
rect 117148 73130 117154 73132
rect 150801 73130 150867 73133
rect 151537 73130 151603 73133
rect 117148 73128 151603 73130
rect 117148 73072 150806 73128
rect 150862 73072 151542 73128
rect 151598 73072 151603 73128
rect 117148 73070 151603 73072
rect 117148 73068 117154 73070
rect 108297 73067 108363 73068
rect 150801 73067 150867 73070
rect 151537 73067 151603 73070
rect 158662 73068 158668 73132
rect 158732 73130 158738 73132
rect 218145 73130 218211 73133
rect 158732 73128 218211 73130
rect 158732 73072 218150 73128
rect 218206 73072 218211 73128
rect 158732 73070 218211 73072
rect 158732 73068 158738 73070
rect 218145 73067 218211 73070
rect 111609 72994 111675 72997
rect 145414 72994 145420 72996
rect 111609 72992 145420 72994
rect 111609 72936 111614 72992
rect 111670 72936 145420 72992
rect 111609 72934 145420 72936
rect 111609 72931 111675 72934
rect 145414 72932 145420 72934
rect 145484 72932 145490 72996
rect 171593 72994 171659 72997
rect 172329 72994 172395 72997
rect 203517 72994 203583 72997
rect 171593 72992 203583 72994
rect 171593 72936 171598 72992
rect 171654 72936 172334 72992
rect 172390 72936 203522 72992
rect 203578 72936 203583 72992
rect 171593 72934 203583 72936
rect 171593 72931 171659 72934
rect 172329 72931 172395 72934
rect 203517 72931 203583 72934
rect 580165 72994 580231 72997
rect 583520 72994 584960 73084
rect 580165 72992 584960 72994
rect 580165 72936 580170 72992
rect 580226 72936 584960 72992
rect 580165 72934 584960 72936
rect 580165 72931 580231 72934
rect 115749 72858 115815 72861
rect 148358 72858 148364 72860
rect 115749 72856 148364 72858
rect 115749 72800 115754 72856
rect 115810 72800 148364 72856
rect 115749 72798 148364 72800
rect 115749 72795 115815 72798
rect 148358 72796 148364 72798
rect 148428 72796 148434 72860
rect 175825 72858 175891 72861
rect 176561 72858 176627 72861
rect 181621 72858 181687 72861
rect 205081 72858 205147 72861
rect 175825 72856 181687 72858
rect 175825 72800 175830 72856
rect 175886 72800 176566 72856
rect 176622 72800 181626 72856
rect 181682 72800 181687 72856
rect 175825 72798 181687 72800
rect 175825 72795 175891 72798
rect 176561 72795 176627 72798
rect 181621 72795 181687 72798
rect 186270 72856 205147 72858
rect 186270 72800 205086 72856
rect 205142 72800 205147 72856
rect 583520 72844 584960 72934
rect 186270 72798 205147 72800
rect 118509 72722 118575 72725
rect 147438 72722 147444 72724
rect 118509 72720 147444 72722
rect 118509 72664 118514 72720
rect 118570 72664 147444 72720
rect 118509 72662 147444 72664
rect 118509 72659 118575 72662
rect 147438 72660 147444 72662
rect 147508 72660 147514 72724
rect 176193 72722 176259 72725
rect 176561 72722 176627 72725
rect 186270 72722 186330 72798
rect 205081 72795 205147 72798
rect 201902 72722 201908 72724
rect 176193 72720 186330 72722
rect 176193 72664 176198 72720
rect 176254 72664 176566 72720
rect 176622 72664 186330 72720
rect 176193 72662 186330 72664
rect 190410 72662 201908 72722
rect 176193 72659 176259 72662
rect 176561 72659 176627 72662
rect 165153 72586 165219 72589
rect 181437 72586 181503 72589
rect 165153 72584 181503 72586
rect 165153 72528 165158 72584
rect 165214 72528 181442 72584
rect 181498 72528 181503 72584
rect 165153 72526 181503 72528
rect 165153 72523 165219 72526
rect 181437 72523 181503 72526
rect 181621 72586 181687 72589
rect 190410 72586 190470 72662
rect 201902 72660 201908 72662
rect 201972 72660 201978 72724
rect 181621 72584 190470 72586
rect 181621 72528 181626 72584
rect 181682 72528 190470 72584
rect 181621 72526 190470 72528
rect 181621 72523 181687 72526
rect 78673 72450 78739 72453
rect 108297 72450 108363 72453
rect 78673 72448 108363 72450
rect 78673 72392 78678 72448
rect 78734 72392 108302 72448
rect 108358 72392 108363 72448
rect 78673 72390 108363 72392
rect 78673 72387 78739 72390
rect 108297 72387 108363 72390
rect 172421 72450 172487 72453
rect 192150 72450 192156 72452
rect 172421 72448 192156 72450
rect 172421 72392 172426 72448
rect 172482 72392 192156 72448
rect 172421 72390 192156 72392
rect 172421 72387 172487 72390
rect 192150 72388 192156 72390
rect 192220 72388 192226 72452
rect 218145 72450 218211 72453
rect 332593 72450 332659 72453
rect 218145 72448 332659 72450
rect 218145 72392 218150 72448
rect 218206 72392 332598 72448
rect 332654 72392 332659 72448
rect 218145 72390 332659 72392
rect 218145 72387 218211 72390
rect 332593 72387 332659 72390
rect 181437 72314 181503 72317
rect 188102 72314 188108 72316
rect 181437 72312 188108 72314
rect 181437 72256 181442 72312
rect 181498 72256 188108 72312
rect 181437 72254 188108 72256
rect 181437 72251 181503 72254
rect 188102 72252 188108 72254
rect 188172 72252 188178 72316
rect 97809 71770 97875 71773
rect 144126 71770 144132 71772
rect 97809 71768 144132 71770
rect -960 71634 480 71724
rect 97809 71712 97814 71768
rect 97870 71712 144132 71768
rect 97809 71710 144132 71712
rect 97809 71707 97875 71710
rect 144126 71708 144132 71710
rect 144196 71708 144202 71772
rect 167913 71770 167979 71773
rect 168281 71770 168347 71773
rect 171225 71770 171291 71773
rect 209037 71770 209103 71773
rect 167913 71768 171058 71770
rect 167913 71712 167918 71768
rect 167974 71712 168286 71768
rect 168342 71712 171058 71768
rect 167913 71710 171058 71712
rect 167913 71707 167979 71710
rect 168281 71707 168347 71710
rect 3509 71634 3575 71637
rect 101213 71634 101279 71637
rect 135713 71634 135779 71637
rect -960 71632 3575 71634
rect -960 71576 3514 71632
rect 3570 71576 3575 71632
rect -960 71574 3575 71576
rect -960 71484 480 71574
rect 3509 71571 3575 71574
rect 84150 71632 135779 71634
rect 84150 71576 101218 71632
rect 101274 71576 135718 71632
rect 135774 71576 135779 71632
rect 84150 71574 135779 71576
rect 52453 71226 52519 71229
rect 84150 71226 84210 71574
rect 101213 71571 101279 71574
rect 135713 71571 135779 71574
rect 167729 71634 167795 71637
rect 168189 71634 168255 71637
rect 170998 71634 171058 71710
rect 171225 71768 209103 71770
rect 171225 71712 171230 71768
rect 171286 71712 209042 71768
rect 209098 71712 209103 71768
rect 171225 71710 209103 71712
rect 171225 71707 171291 71710
rect 209037 71707 209103 71710
rect 200849 71634 200915 71637
rect 167729 71632 170874 71634
rect 167729 71576 167734 71632
rect 167790 71576 168194 71632
rect 168250 71576 170874 71632
rect 167729 71574 170874 71576
rect 170998 71632 200915 71634
rect 170998 71576 200854 71632
rect 200910 71576 200915 71632
rect 170998 71574 200915 71576
rect 167729 71571 167795 71574
rect 168189 71571 168255 71574
rect 115606 71436 115612 71500
rect 115676 71498 115682 71500
rect 149881 71498 149947 71501
rect 115676 71496 149947 71498
rect 115676 71440 149886 71496
rect 149942 71440 149947 71496
rect 115676 71438 149947 71440
rect 170814 71498 170874 71574
rect 200849 71571 200915 71574
rect 171225 71498 171291 71501
rect 170814 71496 171291 71498
rect 170814 71440 171230 71496
rect 171286 71440 171291 71496
rect 170814 71438 171291 71440
rect 115676 71436 115682 71438
rect 149881 71435 149947 71438
rect 171225 71435 171291 71438
rect 173341 71498 173407 71501
rect 205766 71498 205772 71500
rect 173341 71496 205772 71498
rect 173341 71440 173346 71496
rect 173402 71440 205772 71496
rect 173341 71438 205772 71440
rect 173341 71435 173407 71438
rect 205766 71436 205772 71438
rect 205836 71436 205842 71500
rect 100017 71362 100083 71365
rect 134057 71362 134123 71365
rect 100017 71360 134123 71362
rect 100017 71304 100022 71360
rect 100078 71304 134062 71360
rect 134118 71304 134123 71360
rect 100017 71302 134123 71304
rect 100017 71299 100083 71302
rect 134057 71299 134123 71302
rect 170949 71362 171015 71365
rect 196198 71362 196204 71364
rect 170949 71360 196204 71362
rect 170949 71304 170954 71360
rect 171010 71304 196204 71360
rect 170949 71302 196204 71304
rect 170949 71299 171015 71302
rect 196198 71300 196204 71302
rect 196268 71362 196274 71364
rect 498193 71362 498259 71365
rect 196268 71360 498259 71362
rect 196268 71304 498198 71360
rect 498254 71304 498259 71360
rect 196268 71302 498259 71304
rect 196268 71300 196274 71302
rect 498193 71299 498259 71302
rect 107510 71226 107516 71228
rect 52453 71224 84210 71226
rect 52453 71168 52458 71224
rect 52514 71168 84210 71224
rect 52453 71166 84210 71168
rect 103470 71166 107516 71226
rect 52453 71163 52519 71166
rect 17217 71090 17283 71093
rect 103470 71090 103530 71166
rect 107510 71164 107516 71166
rect 107580 71226 107586 71228
rect 128169 71226 128235 71229
rect 107580 71224 128235 71226
rect 107580 71168 128174 71224
rect 128230 71168 128235 71224
rect 107580 71166 128235 71168
rect 107580 71164 107586 71166
rect 128169 71163 128235 71166
rect 175181 71226 175247 71229
rect 175181 71224 200130 71226
rect 175181 71168 175186 71224
rect 175242 71168 200130 71224
rect 175181 71166 200130 71168
rect 175181 71163 175247 71166
rect 17217 71088 103530 71090
rect 17217 71032 17222 71088
rect 17278 71032 103530 71088
rect 17217 71030 103530 71032
rect 169201 71090 169267 71093
rect 181805 71090 181871 71093
rect 169201 71088 181871 71090
rect 169201 71032 169206 71088
rect 169262 71032 181810 71088
rect 181866 71032 181871 71088
rect 169201 71030 181871 71032
rect 200070 71090 200130 71166
rect 205766 71164 205772 71228
rect 205836 71226 205842 71228
rect 531313 71226 531379 71229
rect 205836 71224 531379 71226
rect 205836 71168 531318 71224
rect 531374 71168 531379 71224
rect 205836 71166 531379 71168
rect 205836 71164 205842 71166
rect 531313 71163 531379 71166
rect 201718 71090 201724 71092
rect 200070 71030 201724 71090
rect 17217 71027 17283 71030
rect 169201 71027 169267 71030
rect 181805 71027 181871 71030
rect 201718 71028 201724 71030
rect 201788 71090 201794 71092
rect 549897 71090 549963 71093
rect 201788 71088 549963 71090
rect 201788 71032 549902 71088
rect 549958 71032 549963 71088
rect 201788 71030 549963 71032
rect 201788 71028 201794 71030
rect 549897 71027 549963 71030
rect 185393 70410 185459 70413
rect 185526 70410 185532 70412
rect 185393 70408 185532 70410
rect 185393 70352 185398 70408
rect 185454 70352 185532 70408
rect 185393 70350 185532 70352
rect 185393 70347 185459 70350
rect 185526 70348 185532 70350
rect 185596 70348 185602 70412
rect 112345 70274 112411 70277
rect 146518 70274 146524 70276
rect 112345 70272 146524 70274
rect 112345 70216 112350 70272
rect 112406 70216 146524 70272
rect 112345 70214 146524 70216
rect 112345 70211 112411 70214
rect 146518 70212 146524 70214
rect 146588 70212 146594 70276
rect 120022 70076 120028 70140
rect 120092 70138 120098 70140
rect 154113 70138 154179 70141
rect 120092 70136 154179 70138
rect 120092 70080 154118 70136
rect 154174 70080 154179 70136
rect 120092 70078 154179 70080
rect 120092 70076 120098 70078
rect 154113 70075 154179 70078
rect 166206 70076 166212 70140
rect 166276 70138 166282 70140
rect 166276 70078 200130 70138
rect 166276 70076 166282 70078
rect 120758 69940 120764 70004
rect 120828 70002 120834 70004
rect 154021 70002 154087 70005
rect 190494 70002 190500 70004
rect 120828 70000 154087 70002
rect 120828 69944 154026 70000
rect 154082 69944 154087 70000
rect 120828 69942 154087 69944
rect 120828 69940 120834 69942
rect 154021 69939 154087 69942
rect 171090 69942 190500 70002
rect 121126 69804 121132 69868
rect 121196 69866 121202 69868
rect 152089 69866 152155 69869
rect 121196 69864 152155 69866
rect 121196 69808 152094 69864
rect 152150 69808 152155 69864
rect 121196 69806 152155 69808
rect 121196 69804 121202 69806
rect 152089 69803 152155 69806
rect 163221 69866 163287 69869
rect 164141 69866 164207 69869
rect 171090 69866 171150 69942
rect 190494 69940 190500 69942
rect 190564 69940 190570 70004
rect 163221 69864 171150 69866
rect 163221 69808 163226 69864
rect 163282 69808 164146 69864
rect 164202 69808 171150 69864
rect 163221 69806 171150 69808
rect 175733 69866 175799 69869
rect 175733 69864 190470 69866
rect 175733 69808 175738 69864
rect 175794 69808 190470 69864
rect 175733 69806 190470 69808
rect 163221 69803 163287 69806
rect 164141 69803 164207 69806
rect 175733 69803 175799 69806
rect 122598 69668 122604 69732
rect 122668 69730 122674 69732
rect 153653 69730 153719 69733
rect 122668 69728 153719 69730
rect 122668 69672 153658 69728
rect 153714 69672 153719 69728
rect 122668 69670 153719 69672
rect 122668 69668 122674 69670
rect 153653 69667 153719 69670
rect 117037 69594 117103 69597
rect 146702 69594 146708 69596
rect 117037 69592 146708 69594
rect 117037 69536 117042 69592
rect 117098 69536 146708 69592
rect 117037 69534 146708 69536
rect 117037 69531 117103 69534
rect 146702 69532 146708 69534
rect 146772 69594 146778 69596
rect 147254 69594 147260 69596
rect 146772 69534 147260 69594
rect 146772 69532 146778 69534
rect 147254 69532 147260 69534
rect 147324 69532 147330 69596
rect 172973 69594 173039 69597
rect 173617 69594 173683 69597
rect 190410 69594 190470 69806
rect 200070 69730 200130 70078
rect 200481 69730 200547 69733
rect 430573 69730 430639 69733
rect 200070 69728 430639 69730
rect 200070 69672 200486 69728
rect 200542 69672 430578 69728
rect 430634 69672 430639 69728
rect 200070 69670 430639 69672
rect 200481 69667 200547 69670
rect 430573 69667 430639 69670
rect 200614 69594 200620 69596
rect 172973 69592 180810 69594
rect 172973 69536 172978 69592
rect 173034 69536 173622 69592
rect 173678 69536 180810 69592
rect 172973 69534 180810 69536
rect 190410 69534 200620 69594
rect 172973 69531 173039 69534
rect 173617 69531 173683 69534
rect 180750 69458 180810 69534
rect 200614 69532 200620 69534
rect 200684 69594 200690 69596
rect 557533 69594 557599 69597
rect 200684 69592 557599 69594
rect 200684 69536 557538 69592
rect 557594 69536 557599 69592
rect 200684 69534 557599 69536
rect 200684 69532 200690 69534
rect 557533 69531 557599 69534
rect 207197 69458 207263 69461
rect 180750 69456 207263 69458
rect 180750 69400 207202 69456
rect 207258 69400 207263 69456
rect 180750 69398 207263 69400
rect 207197 69395 207263 69398
rect 112437 68914 112503 68917
rect 115473 68914 115539 68917
rect 140998 68914 141004 68916
rect 112437 68912 141004 68914
rect 112437 68856 112442 68912
rect 112498 68856 115478 68912
rect 115534 68856 141004 68912
rect 112437 68854 141004 68856
rect 112437 68851 112503 68854
rect 115473 68851 115539 68854
rect 140998 68852 141004 68854
rect 141068 68852 141074 68916
rect 149830 68852 149836 68916
rect 149900 68914 149906 68916
rect 215569 68914 215635 68917
rect 220813 68914 220879 68917
rect 149900 68912 220879 68914
rect 149900 68856 215574 68912
rect 215630 68856 220818 68912
rect 220874 68856 220879 68912
rect 149900 68854 220879 68856
rect 149900 68852 149906 68854
rect 215569 68851 215635 68854
rect 220813 68851 220879 68854
rect 116710 68716 116716 68780
rect 116780 68778 116786 68780
rect 155217 68778 155283 68781
rect 116780 68776 155283 68778
rect 116780 68720 155222 68776
rect 155278 68720 155283 68776
rect 116780 68718 155283 68720
rect 116780 68716 116786 68718
rect 155217 68715 155283 68718
rect 161841 68778 161907 68781
rect 189022 68778 189028 68780
rect 161841 68776 189028 68778
rect 161841 68720 161846 68776
rect 161902 68720 189028 68776
rect 161841 68718 189028 68720
rect 161841 68715 161907 68718
rect 189022 68716 189028 68718
rect 189092 68716 189098 68780
rect 122414 68580 122420 68644
rect 122484 68642 122490 68644
rect 156873 68642 156939 68645
rect 122484 68640 156939 68642
rect 122484 68584 156878 68640
rect 156934 68584 156939 68640
rect 122484 68582 156939 68584
rect 122484 68580 122490 68582
rect 156873 68579 156939 68582
rect 161657 68642 161723 68645
rect 162761 68642 162827 68645
rect 185342 68642 185348 68644
rect 161657 68640 185348 68642
rect 161657 68584 161662 68640
rect 161718 68584 162766 68640
rect 162822 68584 185348 68640
rect 161657 68582 185348 68584
rect 161657 68579 161723 68582
rect 162761 68579 162827 68582
rect 185342 68580 185348 68582
rect 185412 68580 185418 68644
rect 111517 68506 111583 68509
rect 143942 68506 143948 68508
rect 111517 68504 143948 68506
rect 111517 68448 111522 68504
rect 111578 68448 143948 68504
rect 111517 68446 143948 68448
rect 111517 68443 111583 68446
rect 143942 68444 143948 68446
rect 144012 68506 144018 68508
rect 144494 68506 144500 68508
rect 144012 68446 144500 68506
rect 144012 68444 144018 68446
rect 144494 68444 144500 68446
rect 144564 68444 144570 68508
rect 177021 68506 177087 68509
rect 177021 68504 180810 68506
rect 177021 68448 177026 68504
rect 177082 68448 180810 68504
rect 177021 68446 180810 68448
rect 177021 68443 177087 68446
rect 111558 68308 111564 68372
rect 111628 68370 111634 68372
rect 138289 68370 138355 68373
rect 111628 68368 138355 68370
rect 111628 68312 138294 68368
rect 138350 68312 138355 68368
rect 111628 68310 138355 68312
rect 111628 68308 111634 68310
rect 138289 68307 138355 68310
rect 145598 68172 145604 68236
rect 145668 68234 145674 68236
rect 178033 68234 178099 68237
rect 145668 68232 178099 68234
rect 145668 68176 178038 68232
rect 178094 68176 178099 68232
rect 145668 68174 178099 68176
rect 180750 68234 180810 68446
rect 194542 68234 194548 68236
rect 180750 68174 194548 68234
rect 145668 68172 145674 68174
rect 178033 68171 178099 68174
rect 194542 68172 194548 68174
rect 194612 68234 194618 68236
rect 574737 68234 574803 68237
rect 194612 68232 574803 68234
rect 194612 68176 574742 68232
rect 574798 68176 574803 68232
rect 194612 68174 574803 68176
rect 194612 68172 194618 68174
rect 574737 68171 574803 68174
rect 110229 68098 110295 68101
rect 143758 68098 143764 68100
rect 110229 68096 143764 68098
rect 110229 68040 110234 68096
rect 110290 68040 143764 68096
rect 110229 68038 143764 68040
rect 110229 68035 110295 68038
rect 143758 68036 143764 68038
rect 143828 68098 143834 68100
rect 144310 68098 144316 68100
rect 143828 68038 144316 68098
rect 143828 68036 143834 68038
rect 144310 68036 144316 68038
rect 144380 68036 144386 68100
rect 156597 67690 156663 67693
rect 156873 67690 156939 67693
rect 156597 67688 156939 67690
rect 156597 67632 156602 67688
rect 156658 67632 156878 67688
rect 156934 67632 156939 67688
rect 156597 67630 156939 67632
rect 156597 67627 156663 67630
rect 156873 67627 156939 67630
rect 110045 67554 110111 67557
rect 143574 67554 143580 67556
rect 110045 67552 143580 67554
rect 110045 67496 110050 67552
rect 110106 67496 143580 67552
rect 110045 67494 143580 67496
rect 110045 67491 110111 67494
rect 143574 67492 143580 67494
rect 143644 67554 143650 67556
rect 144678 67554 144684 67556
rect 143644 67494 144684 67554
rect 143644 67492 143650 67494
rect 144678 67492 144684 67494
rect 144748 67492 144754 67556
rect 154941 67554 155007 67557
rect 155769 67554 155835 67557
rect 154941 67552 161490 67554
rect 154941 67496 154946 67552
rect 155002 67496 155774 67552
rect 155830 67496 161490 67552
rect 154941 67494 161490 67496
rect 154941 67491 155007 67494
rect 155769 67491 155835 67494
rect 114134 67356 114140 67420
rect 114204 67418 114210 67420
rect 147806 67418 147812 67420
rect 114204 67358 147812 67418
rect 114204 67356 114210 67358
rect 147806 67356 147812 67358
rect 147876 67418 147882 67420
rect 148174 67418 148180 67420
rect 147876 67358 148180 67418
rect 147876 67356 147882 67358
rect 148174 67356 148180 67358
rect 148244 67356 148250 67420
rect 161430 67418 161490 67494
rect 193254 67492 193260 67556
rect 193324 67554 193330 67556
rect 193397 67554 193463 67557
rect 193324 67552 193463 67554
rect 193324 67496 193402 67552
rect 193458 67496 193463 67552
rect 193324 67494 193463 67496
rect 193324 67492 193330 67494
rect 193397 67491 193463 67494
rect 201534 67492 201540 67556
rect 201604 67554 201610 67556
rect 201677 67554 201743 67557
rect 201604 67552 201743 67554
rect 201604 67496 201682 67552
rect 201738 67496 201743 67552
rect 201604 67494 201743 67496
rect 201604 67492 201610 67494
rect 201677 67491 201743 67494
rect 184238 67418 184244 67420
rect 161430 67358 184244 67418
rect 184238 67356 184244 67358
rect 184308 67356 184314 67420
rect 116761 67282 116827 67285
rect 147990 67282 147996 67284
rect 116761 67280 147996 67282
rect 116761 67224 116766 67280
rect 116822 67224 147996 67280
rect 116761 67222 147996 67224
rect 116761 67219 116827 67222
rect 147990 67220 147996 67222
rect 148060 67282 148066 67284
rect 148358 67282 148364 67284
rect 148060 67222 148364 67282
rect 148060 67220 148066 67222
rect 148358 67220 148364 67222
rect 148428 67220 148434 67284
rect 160369 67282 160435 67285
rect 161197 67282 161263 67285
rect 186078 67282 186084 67284
rect 160369 67280 186084 67282
rect 160369 67224 160374 67280
rect 160430 67224 161202 67280
rect 161258 67224 186084 67280
rect 160369 67222 186084 67224
rect 160369 67219 160435 67222
rect 161197 67219 161263 67222
rect 186078 67220 186084 67222
rect 186148 67220 186154 67284
rect 160553 67146 160619 67149
rect 161013 67146 161079 67149
rect 184054 67146 184060 67148
rect 160553 67144 184060 67146
rect 160553 67088 160558 67144
rect 160614 67088 161018 67144
rect 161074 67088 184060 67144
rect 160553 67086 184060 67088
rect 160553 67083 160619 67086
rect 161013 67083 161079 67086
rect 184054 67084 184060 67086
rect 184124 67084 184130 67148
rect 150014 66948 150020 67012
rect 150084 67010 150090 67012
rect 215477 67010 215543 67013
rect 227713 67010 227779 67013
rect 150084 67008 227779 67010
rect 150084 66952 215482 67008
rect 215538 66952 227718 67008
rect 227774 66952 227779 67008
rect 150084 66950 227779 66952
rect 150084 66948 150090 66950
rect 215477 66947 215543 66950
rect 227713 66947 227779 66950
rect 77293 66874 77359 66877
rect 109033 66874 109099 66877
rect 109534 66874 109540 66876
rect 77293 66872 109540 66874
rect 77293 66816 77298 66872
rect 77354 66816 109038 66872
rect 109094 66816 109540 66872
rect 77293 66814 109540 66816
rect 77293 66811 77359 66814
rect 109033 66811 109099 66814
rect 109534 66812 109540 66814
rect 109604 66812 109610 66876
rect 148910 66812 148916 66876
rect 148980 66874 148986 66876
rect 204161 66874 204227 66877
rect 148980 66872 204227 66874
rect 148980 66816 204166 66872
rect 204222 66816 204227 66872
rect 148980 66814 204227 66816
rect 148980 66812 148986 66814
rect 204161 66811 204227 66814
rect 199193 66468 199259 66469
rect 199142 66404 199148 66468
rect 199212 66466 199259 66468
rect 199212 66464 199304 66466
rect 199254 66408 199304 66464
rect 199212 66406 199304 66408
rect 199212 66404 199259 66406
rect 199193 66403 199259 66404
rect 115790 66132 115796 66196
rect 115860 66194 115866 66196
rect 156689 66194 156755 66197
rect 115860 66192 156755 66194
rect 115860 66136 156694 66192
rect 156750 66136 156755 66192
rect 115860 66134 156755 66136
rect 115860 66132 115866 66134
rect 156689 66131 156755 66134
rect 196014 66132 196020 66196
rect 196084 66194 196090 66196
rect 196157 66194 196223 66197
rect 196084 66192 196223 66194
rect 196084 66136 196162 66192
rect 196218 66136 196223 66192
rect 196084 66134 196223 66136
rect 196084 66132 196090 66134
rect 196157 66131 196223 66134
rect 118550 65996 118556 66060
rect 118620 66058 118626 66060
rect 152825 66058 152891 66061
rect 118620 66056 152891 66058
rect 118620 66000 152830 66056
rect 152886 66000 152891 66056
rect 118620 65998 152891 66000
rect 118620 65996 118626 65998
rect 152825 65995 152891 65998
rect 164734 65996 164740 66060
rect 164804 66058 164810 66060
rect 164804 65998 200130 66058
rect 164804 65996 164810 65998
rect 124070 65860 124076 65924
rect 124140 65922 124146 65924
rect 152641 65922 152707 65925
rect 124140 65920 152707 65922
rect 124140 65864 152646 65920
rect 152702 65864 152707 65920
rect 124140 65862 152707 65864
rect 124140 65860 124146 65862
rect 152641 65859 152707 65862
rect 93117 65650 93183 65653
rect 108297 65650 108363 65653
rect 108430 65650 108436 65652
rect 93117 65648 108436 65650
rect 93117 65592 93122 65648
rect 93178 65592 108302 65648
rect 108358 65592 108436 65648
rect 93117 65590 108436 65592
rect 93117 65587 93183 65590
rect 108297 65587 108363 65590
rect 108430 65588 108436 65590
rect 108500 65588 108506 65652
rect 8293 65514 8359 65517
rect 104014 65514 104020 65516
rect 8293 65512 104020 65514
rect 8293 65456 8298 65512
rect 8354 65456 104020 65512
rect 8293 65454 104020 65456
rect 8293 65451 8359 65454
rect 104014 65452 104020 65454
rect 104084 65514 104090 65516
rect 104617 65514 104683 65517
rect 104084 65512 104683 65514
rect 104084 65456 104622 65512
rect 104678 65456 104683 65512
rect 104084 65454 104683 65456
rect 200070 65514 200130 65998
rect 213085 65514 213151 65517
rect 402973 65514 403039 65517
rect 200070 65512 403039 65514
rect 200070 65456 213090 65512
rect 213146 65456 402978 65512
rect 403034 65456 403039 65512
rect 200070 65454 403039 65456
rect 104084 65452 104090 65454
rect 104617 65451 104683 65454
rect 213085 65451 213151 65454
rect 402973 65451 403039 65454
rect 198917 64836 198983 64837
rect 198917 64832 198964 64836
rect 199028 64834 199034 64836
rect 198917 64776 198922 64832
rect 198917 64772 198964 64776
rect 199028 64774 199074 64834
rect 199028 64772 199034 64774
rect 198917 64771 198983 64772
rect 171910 64636 171916 64700
rect 171980 64698 171986 64700
rect 212717 64698 212783 64701
rect 171980 64696 212783 64698
rect 171980 64640 212722 64696
rect 212778 64640 212783 64696
rect 171980 64638 212783 64640
rect 171980 64636 171986 64638
rect 212717 64635 212783 64638
rect 160686 64500 160692 64564
rect 160756 64562 160762 64564
rect 194869 64562 194935 64565
rect 160756 64560 194935 64562
rect 160756 64504 194874 64560
rect 194930 64504 194935 64560
rect 160756 64502 194935 64504
rect 160756 64500 160762 64502
rect 194869 64499 194935 64502
rect 152774 64364 152780 64428
rect 152844 64426 152850 64428
rect 215385 64426 215451 64429
rect 242157 64426 242223 64429
rect 152844 64424 242223 64426
rect 152844 64368 215390 64424
rect 215446 64368 242162 64424
rect 242218 64368 242223 64424
rect 152844 64366 242223 64368
rect 152844 64364 152850 64366
rect 215385 64363 215451 64366
rect 242157 64363 242223 64366
rect 194869 64290 194935 64293
rect 362953 64290 363019 64293
rect 194869 64288 363019 64290
rect 194869 64232 194874 64288
rect 194930 64232 362958 64288
rect 363014 64232 363019 64288
rect 194869 64230 363019 64232
rect 194869 64227 194935 64230
rect 362953 64227 363019 64230
rect 97993 64154 98059 64157
rect 111241 64156 111307 64157
rect 111190 64154 111196 64156
rect 97993 64152 111196 64154
rect 111260 64154 111307 64156
rect 111260 64152 111388 64154
rect 97993 64096 97998 64152
rect 98054 64096 111196 64152
rect 111302 64096 111388 64152
rect 97993 64094 111196 64096
rect 97993 64091 98059 64094
rect 111190 64092 111196 64094
rect 111260 64094 111388 64096
rect 111260 64092 111307 64094
rect 147438 64092 147444 64156
rect 147508 64154 147514 64156
rect 188337 64154 188403 64157
rect 147508 64152 188403 64154
rect 147508 64096 188342 64152
rect 188398 64096 188403 64152
rect 147508 64094 188403 64096
rect 147508 64092 147514 64094
rect 111241 64091 111307 64092
rect 188337 64091 188403 64094
rect 212717 64154 212783 64157
rect 511993 64154 512059 64157
rect 212717 64152 512059 64154
rect 212717 64096 212722 64152
rect 212778 64096 511998 64152
rect 512054 64096 512059 64152
rect 212717 64094 512059 64096
rect 212717 64091 212783 64094
rect 511993 64091 512059 64094
rect 187233 63476 187299 63477
rect 100334 63412 100340 63476
rect 100404 63474 100410 63476
rect 133454 63474 133460 63476
rect 100404 63414 133460 63474
rect 100404 63412 100410 63414
rect 133454 63412 133460 63414
rect 133524 63412 133530 63476
rect 187182 63474 187188 63476
rect 187142 63414 187188 63474
rect 187252 63472 187299 63476
rect 187294 63416 187299 63472
rect 187182 63412 187188 63414
rect 187252 63412 187299 63416
rect 187233 63411 187299 63412
rect 115105 63340 115171 63341
rect 115054 63338 115060 63340
rect 115014 63278 115060 63338
rect 115124 63336 115171 63340
rect 115166 63280 115171 63336
rect 115054 63276 115060 63278
rect 115124 63276 115171 63280
rect 167494 63276 167500 63340
rect 167564 63338 167570 63340
rect 201769 63338 201835 63341
rect 202781 63338 202847 63341
rect 167564 63336 202847 63338
rect 167564 63280 201774 63336
rect 201830 63280 202786 63336
rect 202842 63280 202847 63336
rect 167564 63278 202847 63280
rect 167564 63276 167570 63278
rect 115105 63275 115171 63276
rect 201769 63275 201835 63278
rect 202781 63275 202847 63278
rect 88333 62930 88399 62933
rect 115105 62930 115171 62933
rect 88333 62928 115171 62930
rect 88333 62872 88338 62928
rect 88394 62872 115110 62928
rect 115166 62872 115171 62928
rect 88333 62870 115171 62872
rect 88333 62867 88399 62870
rect 115105 62867 115171 62870
rect 148542 62868 148548 62932
rect 148612 62930 148618 62932
rect 213913 62930 213979 62933
rect 148612 62928 213979 62930
rect 148612 62872 213918 62928
rect 213974 62872 213979 62928
rect 148612 62870 213979 62872
rect 148612 62868 148618 62870
rect 213913 62867 213979 62870
rect 2865 62794 2931 62797
rect 100334 62794 100340 62796
rect 2865 62792 100340 62794
rect 2865 62736 2870 62792
rect 2926 62736 100340 62792
rect 2865 62734 100340 62736
rect 2865 62731 2931 62734
rect 100334 62732 100340 62734
rect 100404 62732 100410 62796
rect 202781 62794 202847 62797
rect 446397 62794 446463 62797
rect 202781 62792 446463 62794
rect 202781 62736 202786 62792
rect 202842 62736 446402 62792
rect 446458 62736 446463 62792
rect 202781 62734 446463 62736
rect 202781 62731 202847 62734
rect 446397 62731 446463 62734
rect 100109 62114 100175 62117
rect 202137 62116 202203 62117
rect 134374 62114 134380 62116
rect 100109 62112 134380 62114
rect 100109 62056 100114 62112
rect 100170 62056 134380 62112
rect 100109 62054 134380 62056
rect 100109 62051 100175 62054
rect 134374 62052 134380 62054
rect 134444 62052 134450 62116
rect 167678 62052 167684 62116
rect 167748 62114 167754 62116
rect 202086 62114 202092 62116
rect 167748 62054 200130 62114
rect 202046 62054 202092 62114
rect 202156 62112 202203 62116
rect 202198 62056 202203 62112
rect 167748 62052 167754 62054
rect 106181 61978 106247 61981
rect 138606 61978 138612 61980
rect 103470 61976 138612 61978
rect 103470 61920 106186 61976
rect 106242 61920 138612 61976
rect 103470 61918 138612 61920
rect 75177 61570 75243 61573
rect 103470 61570 103530 61918
rect 106181 61915 106247 61918
rect 138606 61916 138612 61918
rect 138676 61916 138682 61980
rect 176142 61916 176148 61980
rect 176212 61978 176218 61980
rect 176212 61918 180810 61978
rect 176212 61916 176218 61918
rect 75177 61568 103530 61570
rect 75177 61512 75182 61568
rect 75238 61512 103530 61568
rect 75177 61510 103530 61512
rect 75177 61507 75243 61510
rect 27613 61434 27679 61437
rect 100109 61434 100175 61437
rect 27613 61432 100175 61434
rect 27613 61376 27618 61432
rect 27674 61376 100114 61432
rect 100170 61376 100175 61432
rect 27613 61374 100175 61376
rect 180750 61434 180810 61918
rect 200070 61570 200130 62054
rect 202086 62052 202092 62054
rect 202156 62052 202203 62056
rect 202137 62051 202203 62052
rect 202413 61570 202479 61573
rect 459553 61570 459619 61573
rect 200070 61568 459619 61570
rect 200070 61512 202418 61568
rect 202474 61512 459558 61568
rect 459614 61512 459619 61568
rect 200070 61510 459619 61512
rect 202413 61507 202479 61510
rect 459553 61507 459619 61510
rect 200982 61434 200988 61436
rect 180750 61374 200988 61434
rect 27613 61371 27679 61374
rect 100109 61371 100175 61374
rect 200982 61372 200988 61374
rect 201052 61434 201058 61436
rect 563697 61434 563763 61437
rect 201052 61432 563763 61434
rect 201052 61376 563702 61432
rect 563758 61376 563763 61432
rect 201052 61374 563763 61376
rect 201052 61372 201058 61374
rect 563697 61371 563763 61374
rect 98821 60618 98887 60621
rect 99281 60618 99347 60621
rect 133270 60618 133276 60620
rect 98821 60616 133276 60618
rect 98821 60560 98826 60616
rect 98882 60560 99286 60616
rect 99342 60560 133276 60616
rect 98821 60558 133276 60560
rect 98821 60555 98887 60558
rect 99281 60555 99347 60558
rect 133270 60556 133276 60558
rect 133340 60556 133346 60620
rect 170622 60556 170628 60620
rect 170692 60618 170698 60620
rect 170692 60558 200130 60618
rect 170692 60556 170698 60558
rect 105353 60482 105419 60485
rect 138422 60482 138428 60484
rect 103470 60480 138428 60482
rect 103470 60424 105358 60480
rect 105414 60424 138428 60480
rect 103470 60422 138428 60424
rect 81433 60074 81499 60077
rect 103470 60074 103530 60422
rect 105353 60419 105419 60422
rect 138422 60420 138428 60422
rect 138492 60420 138498 60484
rect 81433 60072 103530 60074
rect 81433 60016 81438 60072
rect 81494 60016 103530 60072
rect 81433 60014 103530 60016
rect 81433 60011 81499 60014
rect 4153 59938 4219 59941
rect 98821 59938 98887 59941
rect 4153 59936 98887 59938
rect 4153 59880 4158 59936
rect 4214 59880 98826 59936
rect 98882 59880 98887 59936
rect 4153 59878 98887 59880
rect 200070 59938 200130 60558
rect 203374 59938 203380 59940
rect 200070 59878 203380 59938
rect 4153 59875 4219 59878
rect 98821 59875 98887 59878
rect 203374 59876 203380 59878
rect 203444 59938 203450 59940
rect 484393 59938 484459 59941
rect 203444 59936 484459 59938
rect 203444 59880 484398 59936
rect 484454 59880 484459 59936
rect 203444 59878 484459 59880
rect 203444 59876 203450 59878
rect 484393 59875 484459 59878
rect 580625 59666 580691 59669
rect 583520 59666 584960 59756
rect 580625 59664 584960 59666
rect 580625 59608 580630 59664
rect 580686 59608 584960 59664
rect 580625 59606 584960 59608
rect 580625 59603 580691 59606
rect 583520 59516 584960 59606
rect 111742 59196 111748 59260
rect 111812 59258 111818 59260
rect 112846 59258 112852 59260
rect 111812 59198 112852 59258
rect 111812 59196 111818 59198
rect 112846 59196 112852 59198
rect 112916 59258 112922 59260
rect 139894 59258 139900 59260
rect 112916 59198 139900 59258
rect 112916 59196 112922 59198
rect 139894 59196 139900 59198
rect 139964 59196 139970 59260
rect 153878 59196 153884 59260
rect 153948 59258 153954 59260
rect 153948 59198 209790 59258
rect 153948 59196 153954 59198
rect 139710 59122 139716 59124
rect 113130 59062 139716 59122
rect 93853 58850 93919 58853
rect 112478 58850 112484 58852
rect 93853 58848 112484 58850
rect 93853 58792 93858 58848
rect 93914 58792 112484 58848
rect 93853 58790 112484 58792
rect 93853 58787 93919 58790
rect 112478 58788 112484 58790
rect 112548 58850 112554 58852
rect 113130 58850 113190 59062
rect 139710 59060 139716 59062
rect 139780 59060 139786 59124
rect 162342 59060 162348 59124
rect 162412 59122 162418 59124
rect 196249 59122 196315 59125
rect 162412 59120 204914 59122
rect 162412 59064 196254 59120
rect 196310 59064 204914 59120
rect 162412 59062 204914 59064
rect 162412 59060 162418 59062
rect 196249 59059 196315 59062
rect 167862 58924 167868 58988
rect 167932 58986 167938 58988
rect 167932 58926 200130 58986
rect 167932 58924 167938 58926
rect 112548 58790 113190 58850
rect 112548 58788 112554 58790
rect 172094 58788 172100 58852
rect 172164 58850 172170 58852
rect 172164 58790 180810 58850
rect 172164 58788 172170 58790
rect 92473 58714 92539 58717
rect 111742 58714 111748 58716
rect 92473 58712 111748 58714
rect -960 58578 480 58668
rect 92473 58656 92478 58712
rect 92534 58656 111748 58712
rect 92473 58654 111748 58656
rect 92473 58651 92539 58654
rect 111742 58652 111748 58654
rect 111812 58652 111818 58716
rect 97533 58578 97599 58581
rect 110505 58578 110571 58581
rect 140814 58578 140820 58580
rect -960 58518 674 58578
rect -960 58442 480 58518
rect 614 58442 674 58518
rect 97533 58576 140820 58578
rect 97533 58520 97538 58576
rect 97594 58520 110510 58576
rect 110566 58520 140820 58576
rect 97533 58518 140820 58520
rect 97533 58515 97599 58518
rect 110505 58515 110571 58518
rect 140814 58516 140820 58518
rect 140884 58516 140890 58580
rect 180750 58578 180810 58790
rect 200070 58714 200130 58926
rect 204854 58850 204914 59062
rect 209730 58986 209790 59198
rect 214005 58986 214071 58989
rect 281533 58986 281599 58989
rect 209730 58984 281599 58986
rect 209730 58928 214010 58984
rect 214066 58928 281538 58984
rect 281594 58928 281599 58984
rect 209730 58926 281599 58928
rect 214005 58923 214071 58926
rect 281533 58923 281599 58926
rect 380893 58850 380959 58853
rect 204854 58848 380959 58850
rect 204854 58792 380898 58848
rect 380954 58792 380959 58848
rect 204854 58790 380959 58792
rect 380893 58787 380959 58790
rect 201861 58714 201927 58717
rect 448513 58714 448579 58717
rect 200070 58712 448579 58714
rect 200070 58656 201866 58712
rect 201922 58656 448518 58712
rect 448574 58656 448579 58712
rect 200070 58654 448579 58656
rect 201861 58651 201927 58654
rect 448513 58651 448579 58654
rect 191966 58578 191972 58580
rect 180750 58518 191972 58578
rect 191966 58516 191972 58518
rect 192036 58578 192042 58580
rect 514017 58578 514083 58581
rect 192036 58576 514083 58578
rect 192036 58520 514022 58576
rect 514078 58520 514083 58576
rect 192036 58518 514083 58520
rect 192036 58516 192042 58518
rect 514017 58515 514083 58518
rect -960 58428 674 58442
rect 246 58382 674 58428
rect 246 58034 306 58382
rect 111006 58034 111012 58036
rect 246 57974 111012 58034
rect 111006 57972 111012 57974
rect 111076 57972 111082 58036
rect 100753 57898 100819 57901
rect 101857 57898 101923 57901
rect 134190 57898 134196 57900
rect 100753 57896 134196 57898
rect 100753 57840 100758 57896
rect 100814 57840 101862 57896
rect 101918 57840 134196 57896
rect 100753 57838 134196 57840
rect 100753 57835 100819 57838
rect 101857 57835 101923 57838
rect 134190 57836 134196 57838
rect 134260 57836 134266 57900
rect 158846 57836 158852 57900
rect 158916 57898 158922 57900
rect 193213 57898 193279 57901
rect 158916 57896 209790 57898
rect 158916 57840 193218 57896
rect 193274 57840 209790 57896
rect 158916 57838 209790 57840
rect 158916 57836 158922 57838
rect 193213 57835 193279 57838
rect 107469 57762 107535 57765
rect 138238 57762 138244 57764
rect 103470 57760 138244 57762
rect 103470 57704 107474 57760
rect 107530 57704 138244 57760
rect 103470 57702 138244 57704
rect 80053 57354 80119 57357
rect 103470 57354 103530 57702
rect 107469 57699 107535 57702
rect 138238 57700 138244 57702
rect 138308 57700 138314 57764
rect 165102 57700 165108 57764
rect 165172 57762 165178 57764
rect 198825 57762 198891 57765
rect 203241 57764 203307 57765
rect 203190 57762 203196 57764
rect 165172 57760 200130 57762
rect 165172 57704 198830 57760
rect 198886 57704 200130 57760
rect 165172 57702 200130 57704
rect 203150 57702 203196 57762
rect 203260 57760 203307 57764
rect 203302 57704 203307 57760
rect 165172 57700 165178 57702
rect 198825 57699 198891 57702
rect 197854 57564 197860 57628
rect 197924 57626 197930 57628
rect 197997 57626 198063 57629
rect 197924 57624 198063 57626
rect 197924 57568 198002 57624
rect 198058 57568 198063 57624
rect 197924 57566 198063 57568
rect 197924 57564 197930 57566
rect 197997 57563 198063 57566
rect 80053 57352 103530 57354
rect 80053 57296 80058 57352
rect 80114 57296 103530 57352
rect 80053 57294 103530 57296
rect 80053 57291 80119 57294
rect 25497 57218 25563 57221
rect 100753 57218 100819 57221
rect 25497 57216 100819 57218
rect 25497 57160 25502 57216
rect 25558 57160 100758 57216
rect 100814 57160 100819 57216
rect 25497 57158 100819 57160
rect 25497 57155 25563 57158
rect 100753 57155 100819 57158
rect 147254 57156 147260 57220
rect 147324 57218 147330 57220
rect 187693 57218 187759 57221
rect 147324 57216 187759 57218
rect 147324 57160 187698 57216
rect 187754 57160 187759 57216
rect 147324 57158 187759 57160
rect 200070 57218 200130 57702
rect 203190 57700 203196 57702
rect 203260 57700 203307 57704
rect 203241 57699 203307 57700
rect 209730 57354 209790 57838
rect 349153 57354 349219 57357
rect 209730 57352 349219 57354
rect 209730 57296 349158 57352
rect 349214 57296 349219 57352
rect 209730 57294 349219 57296
rect 349153 57291 349219 57294
rect 418797 57218 418863 57221
rect 200070 57216 418863 57218
rect 200070 57160 418802 57216
rect 418858 57160 418863 57216
rect 200070 57158 418863 57160
rect 147324 57156 147330 57158
rect 187693 57155 187759 57158
rect 418797 57155 418863 57158
rect 99414 56476 99420 56540
rect 99484 56538 99490 56540
rect 100518 56538 100524 56540
rect 99484 56478 100524 56538
rect 99484 56476 99490 56478
rect 100518 56476 100524 56478
rect 100588 56538 100594 56540
rect 133086 56538 133092 56540
rect 100588 56478 133092 56538
rect 100588 56476 100594 56478
rect 133086 56476 133092 56478
rect 133156 56476 133162 56540
rect 170806 56476 170812 56540
rect 170876 56538 170882 56540
rect 208577 56538 208643 56541
rect 208945 56538 209011 56541
rect 170876 56536 209011 56538
rect 170876 56480 208582 56536
rect 208638 56480 208950 56536
rect 209006 56480 209011 56536
rect 170876 56478 209011 56480
rect 170876 56476 170882 56478
rect 208577 56475 208643 56478
rect 208945 56475 209011 56478
rect 162526 56340 162532 56404
rect 162596 56402 162602 56404
rect 196065 56402 196131 56405
rect 162596 56400 196131 56402
rect 162596 56344 196070 56400
rect 196126 56344 196131 56400
rect 162596 56342 196131 56344
rect 162596 56340 162602 56342
rect 196065 56339 196131 56342
rect 154062 56204 154068 56268
rect 154132 56266 154138 56268
rect 186589 56266 186655 56269
rect 284293 56266 284359 56269
rect 154132 56264 284359 56266
rect 154132 56208 186594 56264
rect 186650 56208 284298 56264
rect 284354 56208 284359 56264
rect 154132 56206 284359 56208
rect 154132 56204 154138 56206
rect 186589 56203 186655 56206
rect 284293 56203 284359 56206
rect 196065 56130 196131 56133
rect 382917 56130 382983 56133
rect 196065 56128 382983 56130
rect 196065 56072 196070 56128
rect 196126 56072 382922 56128
rect 382978 56072 382983 56128
rect 196065 56070 382983 56072
rect 196065 56067 196131 56070
rect 382917 56067 382983 56070
rect 60825 55994 60891 55997
rect 104198 55994 104204 55996
rect 60825 55992 104204 55994
rect 60825 55936 60830 55992
rect 60886 55936 104204 55992
rect 60825 55934 104204 55936
rect 60825 55931 60891 55934
rect 104198 55932 104204 55934
rect 104268 55994 104274 55996
rect 104433 55994 104499 55997
rect 104268 55992 104499 55994
rect 104268 55936 104438 55992
rect 104494 55936 104499 55992
rect 104268 55934 104499 55936
rect 104268 55932 104274 55934
rect 104433 55931 104499 55934
rect 168046 55932 168052 55996
rect 168116 55994 168122 55996
rect 201585 55994 201651 55997
rect 450537 55994 450603 55997
rect 168116 55992 450603 55994
rect 168116 55936 201590 55992
rect 201646 55936 450542 55992
rect 450598 55936 450603 55992
rect 168116 55934 450603 55936
rect 168116 55932 168122 55934
rect 201585 55931 201651 55934
rect 450537 55931 450603 55934
rect 12433 55858 12499 55861
rect 99414 55858 99420 55860
rect 12433 55856 99420 55858
rect 12433 55800 12438 55856
rect 12494 55800 99420 55856
rect 12433 55798 99420 55800
rect 12433 55795 12499 55798
rect 99414 55796 99420 55798
rect 99484 55796 99490 55860
rect 208945 55858 209011 55861
rect 482277 55858 482343 55861
rect 208945 55856 482343 55858
rect 208945 55800 208950 55856
rect 209006 55800 482282 55856
rect 482338 55800 482343 55856
rect 208945 55798 482343 55800
rect 208945 55795 209011 55798
rect 482277 55795 482343 55798
rect 84193 55178 84259 55181
rect 104801 55178 104867 55181
rect 138054 55178 138060 55180
rect 84193 55176 138060 55178
rect 84193 55120 84198 55176
rect 84254 55120 104806 55176
rect 104862 55120 138060 55176
rect 84193 55118 138060 55120
rect 84193 55115 84259 55118
rect 104801 55115 104867 55118
rect 138054 55116 138060 55118
rect 138124 55116 138130 55180
rect 172278 55116 172284 55180
rect 172348 55178 172354 55180
rect 211337 55178 211403 55181
rect 172348 55176 211403 55178
rect 172348 55120 211342 55176
rect 211398 55120 211403 55176
rect 172348 55118 211403 55120
rect 172348 55116 172354 55118
rect 211337 55115 211403 55118
rect 105445 55042 105511 55045
rect 137502 55042 137508 55044
rect 105445 55040 137508 55042
rect 105445 54984 105450 55040
rect 105506 54984 137508 55040
rect 105445 54982 137508 54984
rect 105445 54979 105511 54982
rect 137502 54980 137508 54982
rect 137572 54980 137578 55044
rect 166390 54980 166396 55044
rect 166460 55042 166466 55044
rect 200389 55042 200455 55045
rect 201401 55042 201467 55045
rect 166460 55040 201467 55042
rect 166460 54984 200394 55040
rect 200450 54984 201406 55040
rect 201462 54984 201467 55040
rect 166460 54982 201467 54984
rect 166460 54980 166466 54982
rect 200389 54979 200455 54982
rect 201401 54979 201467 54982
rect 160870 54844 160876 54908
rect 160940 54906 160946 54908
rect 194777 54906 194843 54909
rect 369853 54906 369919 54909
rect 160940 54904 369919 54906
rect 160940 54848 194782 54904
rect 194838 54848 369858 54904
rect 369914 54848 369919 54904
rect 160940 54846 369919 54848
rect 160940 54844 160946 54846
rect 194777 54843 194843 54846
rect 369853 54843 369919 54846
rect 201401 54770 201467 54773
rect 432597 54770 432663 54773
rect 201401 54768 432663 54770
rect 201401 54712 201406 54768
rect 201462 54712 432602 54768
rect 432658 54712 432663 54768
rect 201401 54710 432663 54712
rect 201401 54707 201467 54710
rect 432597 54707 432663 54710
rect 176326 54572 176332 54636
rect 176396 54634 176402 54636
rect 211337 54634 211403 54637
rect 507853 54634 507919 54637
rect 176396 54574 200130 54634
rect 176396 54572 176402 54574
rect 56593 54498 56659 54501
rect 105445 54498 105511 54501
rect 56593 54496 105511 54498
rect 56593 54440 56598 54496
rect 56654 54440 105450 54496
rect 105506 54440 105511 54496
rect 56593 54438 105511 54440
rect 200070 54498 200130 54574
rect 211337 54632 507919 54634
rect 211337 54576 211342 54632
rect 211398 54576 507858 54632
rect 507914 54576 507919 54632
rect 211337 54574 507919 54576
rect 211337 54571 211403 54574
rect 507853 54571 507919 54574
rect 209814 54498 209820 54500
rect 200070 54438 209820 54498
rect 56593 54435 56659 54438
rect 105445 54435 105511 54438
rect 209814 54436 209820 54438
rect 209884 54498 209890 54500
rect 560937 54498 561003 54501
rect 209884 54496 561003 54498
rect 209884 54440 560942 54496
rect 560998 54440 561003 54496
rect 209884 54438 561003 54440
rect 209884 54436 209890 54438
rect 560937 54435 561003 54438
rect 103094 53818 103100 53820
rect 84150 53758 103100 53818
rect 49693 53138 49759 53141
rect 84150 53138 84210 53758
rect 103094 53756 103100 53758
rect 103164 53818 103170 53820
rect 135662 53818 135668 53820
rect 103164 53758 135668 53818
rect 103164 53756 103170 53758
rect 135662 53756 135668 53758
rect 135732 53756 135738 53820
rect 166574 53756 166580 53820
rect 166644 53818 166650 53820
rect 200297 53818 200363 53821
rect 201401 53818 201467 53821
rect 166644 53816 201467 53818
rect 166644 53760 200302 53816
rect 200358 53760 201406 53816
rect 201462 53760 201467 53816
rect 166644 53758 201467 53760
rect 166644 53756 166650 53758
rect 200297 53755 200363 53758
rect 201401 53755 201467 53758
rect 106641 53682 106707 53685
rect 139526 53682 139532 53684
rect 106641 53680 139532 53682
rect 106641 53624 106646 53680
rect 106702 53624 139532 53680
rect 106641 53622 139532 53624
rect 106641 53619 106707 53622
rect 139526 53620 139532 53622
rect 139596 53620 139602 53684
rect 161054 53620 161060 53684
rect 161124 53682 161130 53684
rect 194593 53682 194659 53685
rect 161124 53680 209790 53682
rect 161124 53624 194598 53680
rect 194654 53624 209790 53680
rect 161124 53622 209790 53624
rect 161124 53620 161130 53622
rect 194593 53619 194659 53622
rect 169334 53484 169340 53548
rect 169404 53546 169410 53548
rect 169404 53486 200130 53546
rect 169404 53484 169410 53486
rect 102133 53274 102199 53277
rect 106641 53274 106707 53277
rect 102133 53272 106707 53274
rect 102133 53216 102138 53272
rect 102194 53216 106646 53272
rect 106702 53216 106707 53272
rect 102133 53214 106707 53216
rect 102133 53211 102199 53214
rect 106641 53211 106707 53214
rect 49693 53136 84210 53138
rect 49693 53080 49698 53136
rect 49754 53080 84210 53136
rect 49693 53078 84210 53080
rect 200070 53138 200130 53486
rect 209730 53410 209790 53622
rect 364977 53410 365043 53413
rect 209730 53408 365043 53410
rect 209730 53352 364982 53408
rect 365038 53352 365043 53408
rect 209730 53350 365043 53352
rect 364977 53347 365043 53350
rect 201401 53274 201467 53277
rect 437473 53274 437539 53277
rect 201401 53272 437539 53274
rect 201401 53216 201406 53272
rect 201462 53216 437478 53272
rect 437534 53216 437539 53272
rect 201401 53214 437539 53216
rect 201401 53211 201467 53214
rect 437473 53211 437539 53214
rect 201166 53138 201172 53140
rect 200070 53078 201172 53138
rect 49693 53075 49759 53078
rect 201166 53076 201172 53078
rect 201236 53138 201242 53140
rect 474733 53138 474799 53141
rect 201236 53136 474799 53138
rect 201236 53080 474738 53136
rect 474794 53080 474799 53136
rect 201236 53078 474799 53080
rect 201236 53076 201242 53078
rect 474733 53075 474799 53078
rect 163262 52396 163268 52460
rect 163332 52458 163338 52460
rect 197629 52458 197695 52461
rect 198273 52458 198339 52461
rect 163332 52456 198339 52458
rect 163332 52400 197634 52456
rect 197690 52400 198278 52456
rect 198334 52400 198339 52456
rect 163332 52398 198339 52400
rect 163332 52396 163338 52398
rect 197629 52395 197695 52398
rect 198273 52395 198339 52398
rect 159030 52260 159036 52324
rect 159100 52322 159106 52324
rect 193305 52322 193371 52325
rect 194501 52322 194567 52325
rect 159100 52320 194567 52322
rect 159100 52264 193310 52320
rect 193366 52264 194506 52320
rect 194562 52264 194567 52320
rect 159100 52262 194567 52264
rect 159100 52260 159106 52262
rect 193305 52259 193371 52262
rect 194501 52259 194567 52262
rect 156638 52124 156644 52188
rect 156708 52186 156714 52188
rect 190729 52186 190795 52189
rect 320173 52186 320239 52189
rect 156708 52184 320239 52186
rect 156708 52128 190734 52184
rect 190790 52128 320178 52184
rect 320234 52128 320239 52184
rect 156708 52126 320239 52128
rect 156708 52124 156714 52126
rect 190729 52123 190795 52126
rect 320173 52123 320239 52126
rect 194501 52050 194567 52053
rect 356053 52050 356119 52053
rect 194501 52048 356119 52050
rect 194501 51992 194506 52048
rect 194562 51992 356058 52048
rect 356114 51992 356119 52048
rect 194501 51990 356119 51992
rect 194501 51987 194567 51990
rect 356053 51987 356119 51990
rect 198273 51914 198339 51917
rect 400857 51914 400923 51917
rect 198273 51912 400923 51914
rect 198273 51856 198278 51912
rect 198334 51856 400862 51912
rect 400918 51856 400923 51912
rect 198273 51854 400923 51856
rect 198273 51851 198339 51854
rect 400857 51851 400923 51854
rect 144678 51716 144684 51780
rect 144748 51778 144754 51780
rect 160185 51778 160251 51781
rect 144748 51776 160251 51778
rect 144748 51720 160190 51776
rect 160246 51720 160251 51776
rect 144748 51718 160251 51720
rect 144748 51716 144754 51718
rect 160185 51715 160251 51718
rect 174486 51716 174492 51780
rect 174556 51778 174562 51780
rect 208485 51778 208551 51781
rect 542353 51778 542419 51781
rect 174556 51776 542419 51778
rect 174556 51720 208490 51776
rect 208546 51720 542358 51776
rect 542414 51720 542419 51776
rect 174556 51718 542419 51720
rect 174556 51716 174562 51718
rect 208485 51715 208551 51718
rect 542353 51715 542419 51718
rect 99465 50962 99531 50965
rect 100569 50962 100635 50965
rect 134006 50962 134012 50964
rect 99465 50960 134012 50962
rect 99465 50904 99470 50960
rect 99526 50904 100574 50960
rect 100630 50904 134012 50960
rect 99465 50902 134012 50904
rect 99465 50899 99531 50902
rect 100569 50899 100635 50902
rect 134006 50900 134012 50902
rect 134076 50900 134082 50964
rect 152406 50900 152412 50964
rect 152476 50962 152482 50964
rect 215293 50962 215359 50965
rect 152476 50960 219450 50962
rect 152476 50904 215298 50960
rect 215354 50904 219450 50960
rect 152476 50902 219450 50904
rect 152476 50900 152482 50902
rect 215293 50899 215359 50902
rect 116894 50826 116900 50828
rect 103470 50766 116900 50826
rect 95233 50418 95299 50421
rect 103470 50418 103530 50766
rect 116894 50764 116900 50766
rect 116964 50826 116970 50828
rect 139342 50826 139348 50828
rect 116964 50766 139348 50826
rect 116964 50764 116970 50766
rect 139342 50764 139348 50766
rect 139412 50764 139418 50828
rect 158110 50764 158116 50828
rect 158180 50826 158186 50828
rect 191782 50826 191788 50828
rect 158180 50766 191788 50826
rect 158180 50764 158186 50766
rect 191782 50764 191788 50766
rect 191852 50826 191858 50828
rect 193070 50826 193076 50828
rect 191852 50766 193076 50826
rect 191852 50764 191858 50766
rect 193070 50764 193076 50766
rect 193140 50764 193146 50828
rect 175958 50628 175964 50692
rect 176028 50690 176034 50692
rect 209998 50690 210004 50692
rect 176028 50630 210004 50690
rect 176028 50628 176034 50630
rect 209998 50628 210004 50630
rect 210068 50690 210074 50692
rect 211102 50690 211108 50692
rect 210068 50630 211108 50690
rect 210068 50628 210074 50630
rect 211102 50628 211108 50630
rect 211172 50628 211178 50692
rect 219390 50690 219450 50902
rect 256693 50690 256759 50693
rect 219390 50688 256759 50690
rect 219390 50632 256698 50688
rect 256754 50632 256759 50688
rect 219390 50630 256759 50632
rect 256693 50627 256759 50630
rect 193070 50492 193076 50556
rect 193140 50554 193146 50556
rect 338113 50554 338179 50557
rect 193140 50552 338179 50554
rect 193140 50496 338118 50552
rect 338174 50496 338179 50552
rect 193140 50494 338179 50496
rect 193140 50492 193146 50494
rect 338113 50491 338179 50494
rect 95233 50416 103530 50418
rect 95233 50360 95238 50416
rect 95294 50360 103530 50416
rect 95233 50358 103530 50360
rect 95233 50355 95299 50358
rect 161238 50356 161244 50420
rect 161308 50418 161314 50420
rect 194685 50418 194751 50421
rect 373993 50418 374059 50421
rect 161308 50416 374059 50418
rect 161308 50360 194690 50416
rect 194746 50360 373998 50416
rect 374054 50360 374059 50416
rect 161308 50358 374059 50360
rect 161308 50356 161314 50358
rect 194685 50355 194751 50358
rect 373993 50355 374059 50358
rect 27705 50282 27771 50285
rect 99465 50282 99531 50285
rect 27705 50280 99531 50282
rect 27705 50224 27710 50280
rect 27766 50224 99470 50280
rect 99526 50224 99531 50280
rect 27705 50222 99531 50224
rect 27705 50219 27771 50222
rect 99465 50219 99531 50222
rect 147070 50220 147076 50284
rect 147140 50282 147146 50284
rect 193305 50282 193371 50285
rect 147140 50280 193371 50282
rect 147140 50224 193310 50280
rect 193366 50224 193371 50280
rect 147140 50222 193371 50224
rect 147140 50220 147146 50222
rect 193305 50219 193371 50222
rect 211102 50220 211108 50284
rect 211172 50282 211178 50284
rect 556153 50282 556219 50285
rect 211172 50280 556219 50282
rect 211172 50224 556158 50280
rect 556214 50224 556219 50280
rect 211172 50222 556219 50224
rect 211172 50220 211178 50222
rect 556153 50219 556219 50222
rect 99465 49602 99531 49605
rect 100661 49602 100727 49605
rect 133822 49602 133828 49604
rect 99465 49600 133828 49602
rect 99465 49544 99470 49600
rect 99526 49544 100666 49600
rect 100722 49544 133828 49600
rect 99465 49542 133828 49544
rect 99465 49539 99531 49542
rect 100661 49539 100727 49542
rect 133822 49540 133828 49542
rect 133892 49540 133898 49604
rect 174670 49540 174676 49604
rect 174740 49602 174746 49604
rect 212625 49602 212691 49605
rect 213821 49602 213887 49605
rect 174740 49600 213887 49602
rect 174740 49544 212630 49600
rect 212686 49544 213826 49600
rect 213882 49544 213887 49600
rect 174740 49542 213887 49544
rect 174740 49540 174746 49542
rect 212625 49539 212691 49542
rect 213821 49539 213887 49542
rect 162710 49404 162716 49468
rect 162780 49466 162786 49468
rect 195973 49466 196039 49469
rect 196433 49466 196499 49469
rect 162780 49464 196499 49466
rect 162780 49408 195978 49464
rect 196034 49408 196438 49464
rect 196494 49408 196499 49464
rect 162780 49406 196499 49408
rect 162780 49404 162786 49406
rect 195973 49403 196039 49406
rect 196433 49403 196499 49406
rect 171726 49268 171732 49332
rect 171796 49330 171802 49332
rect 204989 49330 205055 49333
rect 171796 49328 205055 49330
rect 171796 49272 204994 49328
rect 205050 49272 205055 49328
rect 171796 49270 205055 49272
rect 171796 49268 171802 49270
rect 204989 49267 205055 49270
rect 196433 49194 196499 49197
rect 387793 49194 387859 49197
rect 196433 49192 387859 49194
rect 196433 49136 196438 49192
rect 196494 49136 387798 49192
rect 387854 49136 387859 49192
rect 196433 49134 387859 49136
rect 196433 49131 196499 49134
rect 387793 49131 387859 49134
rect 204989 49058 205055 49061
rect 489913 49058 489979 49061
rect 204989 49056 489979 49058
rect 204989 49000 204994 49056
rect 205050 49000 489918 49056
rect 489974 49000 489979 49056
rect 204989 48998 489979 49000
rect 204989 48995 205055 48998
rect 489913 48995 489979 48998
rect 30373 48922 30439 48925
rect 99465 48922 99531 48925
rect 30373 48920 99531 48922
rect 30373 48864 30378 48920
rect 30434 48864 99470 48920
rect 99526 48864 99531 48920
rect 30373 48862 99531 48864
rect 30373 48859 30439 48862
rect 99465 48859 99531 48862
rect 213821 48922 213887 48925
rect 547873 48922 547939 48925
rect 213821 48920 547939 48922
rect 213821 48864 213826 48920
rect 213882 48864 547878 48920
rect 547934 48864 547939 48920
rect 213821 48862 547939 48864
rect 213821 48859 213887 48862
rect 547873 48859 547939 48862
rect 100753 48242 100819 48245
rect 101949 48242 102015 48245
rect 203057 48244 203123 48245
rect 135478 48242 135484 48244
rect 100753 48240 135484 48242
rect 100753 48184 100758 48240
rect 100814 48184 101954 48240
rect 102010 48184 135484 48240
rect 100753 48182 135484 48184
rect 100753 48179 100819 48182
rect 101949 48179 102015 48182
rect 135478 48180 135484 48182
rect 135548 48180 135554 48244
rect 203006 48242 203012 48244
rect 202966 48182 203012 48242
rect 203076 48240 203123 48244
rect 203118 48184 203123 48240
rect 203006 48180 203012 48182
rect 203076 48180 203123 48184
rect 203057 48179 203123 48180
rect 163446 48044 163452 48108
rect 163516 48106 163522 48108
rect 197537 48106 197603 48109
rect 163516 48104 197603 48106
rect 163516 48048 197542 48104
rect 197598 48048 197603 48104
rect 163516 48046 197603 48048
rect 163516 48044 163522 48046
rect 197537 48043 197603 48046
rect 169518 47908 169524 47972
rect 169588 47970 169594 47972
rect 202822 47970 202828 47972
rect 169588 47910 202828 47970
rect 169588 47908 169594 47910
rect 202822 47908 202828 47910
rect 202892 47970 202898 47972
rect 204110 47970 204116 47972
rect 202892 47910 204116 47970
rect 202892 47908 202898 47910
rect 204110 47908 204116 47910
rect 204180 47908 204186 47972
rect 197537 47834 197603 47837
rect 405733 47834 405799 47837
rect 197537 47832 405799 47834
rect 197537 47776 197542 47832
rect 197598 47776 405738 47832
rect 405794 47776 405799 47832
rect 197537 47774 405799 47776
rect 197537 47771 197603 47774
rect 405733 47771 405799 47774
rect 204110 47636 204116 47700
rect 204180 47698 204186 47700
rect 468477 47698 468543 47701
rect 204180 47696 468543 47698
rect 204180 47640 468482 47696
rect 468538 47640 468543 47696
rect 204180 47638 468543 47640
rect 204180 47636 204186 47638
rect 468477 47635 468543 47638
rect 39297 47562 39363 47565
rect 100753 47562 100819 47565
rect 39297 47560 100819 47562
rect 39297 47504 39302 47560
rect 39358 47504 100758 47560
rect 100814 47504 100819 47560
rect 39297 47502 100819 47504
rect 39297 47499 39363 47502
rect 100753 47499 100819 47502
rect 170438 47500 170444 47564
rect 170508 47562 170514 47564
rect 209957 47562 210023 47565
rect 490005 47562 490071 47565
rect 170508 47560 490071 47562
rect 170508 47504 209962 47560
rect 210018 47504 490010 47560
rect 490066 47504 490071 47560
rect 170508 47502 490071 47504
rect 170508 47500 170514 47502
rect 209957 47499 210023 47502
rect 490005 47499 490071 47502
rect 100753 46882 100819 46885
rect 102041 46882 102107 46885
rect 135294 46882 135300 46884
rect 100753 46880 135300 46882
rect 100753 46824 100758 46880
rect 100814 46824 102046 46880
rect 102102 46824 135300 46880
rect 100753 46822 135300 46824
rect 100753 46819 100819 46822
rect 102041 46819 102107 46822
rect 135294 46820 135300 46822
rect 135364 46820 135370 46884
rect 165286 46820 165292 46884
rect 165356 46882 165362 46884
rect 198774 46882 198780 46884
rect 165356 46822 198780 46882
rect 165356 46820 165362 46822
rect 198774 46820 198780 46822
rect 198844 46882 198850 46884
rect 198844 46822 200130 46882
rect 198844 46820 198850 46822
rect 44173 46202 44239 46205
rect 100753 46202 100819 46205
rect 44173 46200 100819 46202
rect 44173 46144 44178 46200
rect 44234 46144 100758 46200
rect 100814 46144 100819 46200
rect 44173 46142 100819 46144
rect 44173 46139 44239 46142
rect 100753 46139 100819 46142
rect 146886 46140 146892 46204
rect 146956 46202 146962 46204
rect 191833 46202 191899 46205
rect 146956 46200 191899 46202
rect 146956 46144 191838 46200
rect 191894 46144 191899 46200
rect 146956 46142 191899 46144
rect 200070 46202 200130 46822
rect 207105 46610 207171 46613
rect 207238 46610 207244 46612
rect 207105 46608 207244 46610
rect 207105 46552 207110 46608
rect 207166 46552 207244 46608
rect 207105 46550 207244 46552
rect 207105 46547 207171 46550
rect 207238 46548 207244 46550
rect 207308 46610 207314 46612
rect 207841 46610 207907 46613
rect 207308 46608 207907 46610
rect 207308 46552 207846 46608
rect 207902 46552 207907 46608
rect 207308 46550 207907 46552
rect 207308 46548 207314 46550
rect 207841 46547 207907 46550
rect 580533 46338 580599 46341
rect 583520 46338 584960 46428
rect 580533 46336 584960 46338
rect 580533 46280 580538 46336
rect 580594 46280 584960 46336
rect 580533 46278 584960 46280
rect 580533 46275 580599 46278
rect 423765 46202 423831 46205
rect 200070 46200 423831 46202
rect 200070 46144 423770 46200
rect 423826 46144 423831 46200
rect 583520 46188 584960 46278
rect 200070 46142 423831 46144
rect 146956 46140 146962 46142
rect 191833 46139 191899 46142
rect 423765 46139 423831 46142
rect -960 45522 480 45612
rect -960 45462 674 45522
rect -960 45386 480 45462
rect 614 45386 674 45462
rect 154246 45460 154252 45524
rect 154316 45522 154322 45524
rect 218053 45522 218119 45525
rect 154316 45520 219450 45522
rect 154316 45464 218058 45520
rect 218114 45464 219450 45520
rect 154316 45462 219450 45464
rect 154316 45460 154322 45462
rect 218053 45459 218119 45462
rect -960 45372 674 45386
rect 246 45326 674 45372
rect 246 44842 306 45326
rect 166758 45324 166764 45388
rect 166828 45386 166834 45388
rect 200205 45386 200271 45389
rect 166828 45384 209790 45386
rect 166828 45328 200210 45384
rect 200266 45328 209790 45384
rect 166828 45326 209790 45328
rect 166828 45324 166834 45326
rect 200205 45323 200271 45326
rect 173566 45188 173572 45252
rect 173636 45250 173642 45252
rect 207013 45250 207079 45253
rect 173636 45248 207079 45250
rect 173636 45192 207018 45248
rect 207074 45192 207079 45248
rect 173636 45190 207079 45192
rect 173636 45188 173642 45190
rect 207013 45187 207079 45190
rect 209730 45114 209790 45326
rect 219390 45250 219450 45462
rect 279417 45250 279483 45253
rect 219390 45248 279483 45250
rect 219390 45192 279422 45248
rect 279478 45192 279483 45248
rect 219390 45190 279483 45192
rect 279417 45187 279483 45190
rect 440233 45114 440299 45117
rect 209730 45112 440299 45114
rect 209730 45056 440238 45112
rect 440294 45056 440299 45112
rect 209730 45054 440299 45056
rect 440233 45051 440299 45054
rect 173750 44916 173756 44980
rect 173820 44978 173826 44980
rect 204529 44978 204595 44981
rect 520917 44978 520983 44981
rect 173820 44976 520983 44978
rect 173820 44920 204534 44976
rect 204590 44920 520922 44976
rect 520978 44920 520983 44976
rect 173820 44918 520983 44920
rect 173820 44916 173826 44918
rect 204529 44915 204595 44918
rect 520917 44915 520983 44918
rect 207013 44842 207079 44845
rect 528553 44842 528619 44845
rect 246 44782 6930 44842
rect 6870 44298 6930 44782
rect 207013 44840 528619 44842
rect 207013 44784 207018 44840
rect 207074 44784 528558 44840
rect 528614 44784 528619 44840
rect 207013 44782 528619 44784
rect 207013 44779 207079 44782
rect 528553 44779 528619 44782
rect 116526 44298 116532 44300
rect 6870 44238 116532 44298
rect 116526 44236 116532 44238
rect 116596 44236 116602 44300
rect 102225 44162 102291 44165
rect 102685 44162 102751 44165
rect 136582 44162 136588 44164
rect 102225 44160 136588 44162
rect 102225 44104 102230 44160
rect 102286 44104 102690 44160
rect 102746 44104 136588 44160
rect 102225 44102 136588 44104
rect 102225 44099 102291 44102
rect 102685 44099 102751 44102
rect 136582 44100 136588 44102
rect 136652 44100 136658 44164
rect 163630 44100 163636 44164
rect 163700 44162 163706 44164
rect 197353 44162 197419 44165
rect 163700 44160 197419 44162
rect 163700 44104 197358 44160
rect 197414 44104 197419 44160
rect 163700 44102 197419 44104
rect 163700 44100 163706 44102
rect 197353 44099 197419 44102
rect 207013 44164 207079 44165
rect 207013 44160 207060 44164
rect 207124 44162 207130 44164
rect 207013 44104 207018 44160
rect 207013 44100 207060 44104
rect 207124 44102 207170 44162
rect 207124 44100 207130 44102
rect 207013 44099 207079 44100
rect 156822 43964 156828 44028
rect 156892 44026 156898 44028
rect 190453 44026 190519 44029
rect 191741 44026 191807 44029
rect 156892 44024 191807 44026
rect 156892 43968 190458 44024
rect 190514 43968 191746 44024
rect 191802 43968 191807 44024
rect 156892 43966 191807 43968
rect 156892 43964 156898 43966
rect 190453 43963 190519 43966
rect 191741 43963 191807 43966
rect 148358 43828 148364 43892
rect 148428 43890 148434 43892
rect 209865 43890 209931 43893
rect 148428 43888 209931 43890
rect 148428 43832 209870 43888
rect 209926 43832 209931 43888
rect 148428 43830 209931 43832
rect 148428 43828 148434 43830
rect 209865 43827 209931 43830
rect 191741 43754 191807 43757
rect 309133 43754 309199 43757
rect 191741 43752 309199 43754
rect 191741 43696 191746 43752
rect 191802 43696 309138 43752
rect 309194 43696 309199 43752
rect 191741 43694 309199 43696
rect 191741 43691 191807 43694
rect 309133 43691 309199 43694
rect 197353 43618 197419 43621
rect 408493 43618 408559 43621
rect 197353 43616 408559 43618
rect 197353 43560 197358 43616
rect 197414 43560 408498 43616
rect 408554 43560 408559 43616
rect 197353 43558 408559 43560
rect 197353 43555 197419 43558
rect 408493 43555 408559 43558
rect 63493 43482 63559 43485
rect 102225 43482 102291 43485
rect 63493 43480 102291 43482
rect 63493 43424 63498 43480
rect 63554 43424 102230 43480
rect 102286 43424 102291 43480
rect 63493 43422 102291 43424
rect 63493 43419 63559 43422
rect 102225 43419 102291 43422
rect 174854 43420 174860 43484
rect 174924 43482 174930 43484
rect 208393 43482 208459 43485
rect 534717 43482 534783 43485
rect 174924 43480 534783 43482
rect 174924 43424 208398 43480
rect 208454 43424 534722 43480
rect 534778 43424 534783 43480
rect 174924 43422 534783 43424
rect 174924 43420 174930 43422
rect 208393 43419 208459 43422
rect 534717 43419 534783 43422
rect 155534 42740 155540 42804
rect 155604 42802 155610 42804
rect 210693 42802 210759 42805
rect 211061 42802 211127 42805
rect 155604 42800 211127 42802
rect 155604 42744 210698 42800
rect 210754 42744 211066 42800
rect 211122 42744 211127 42800
rect 155604 42742 211127 42744
rect 155604 42740 155610 42742
rect 210693 42739 210759 42742
rect 211061 42739 211127 42742
rect 211061 42122 211127 42125
rect 300853 42122 300919 42125
rect 211061 42120 300919 42122
rect 211061 42064 211066 42120
rect 211122 42064 300858 42120
rect 300914 42064 300919 42120
rect 211061 42062 300919 42064
rect 211061 42059 211127 42062
rect 300853 42059 300919 42062
rect 154430 38524 154436 38588
rect 154500 38586 154506 38588
rect 187785 38586 187851 38589
rect 154500 38584 187851 38586
rect 154500 38528 187790 38584
rect 187846 38528 187851 38584
rect 154500 38526 187851 38528
rect 154500 38524 154506 38526
rect 187785 38523 187851 38526
rect 144494 37844 144500 37908
rect 144564 37906 144570 37908
rect 155953 37906 156019 37909
rect 144564 37904 156019 37906
rect 144564 37848 155958 37904
rect 156014 37848 156019 37904
rect 144564 37846 156019 37848
rect 144564 37844 144570 37846
rect 155953 37843 156019 37846
rect 187785 37906 187851 37909
rect 275277 37906 275343 37909
rect 187785 37904 275343 37906
rect 187785 37848 187790 37904
rect 187846 37848 275282 37904
rect 275338 37848 275343 37904
rect 187785 37846 275343 37848
rect 187785 37843 187851 37846
rect 275277 37843 275343 37846
rect 175038 37164 175044 37228
rect 175108 37226 175114 37228
rect 214097 37226 214163 37229
rect 214373 37226 214439 37229
rect 175108 37224 214439 37226
rect 175108 37168 214102 37224
rect 214158 37168 214378 37224
rect 214434 37168 214439 37224
rect 175108 37166 214439 37168
rect 175108 37164 175114 37166
rect 214097 37163 214163 37166
rect 214373 37163 214439 37166
rect 214373 36546 214439 36549
rect 534073 36546 534139 36549
rect 214373 36544 534139 36546
rect 214373 36488 214378 36544
rect 214434 36488 534078 36544
rect 534134 36488 534139 36544
rect 214373 36486 534139 36488
rect 214373 36483 214439 36486
rect 534073 36483 534139 36486
rect 165470 35804 165476 35868
rect 165540 35866 165546 35868
rect 206093 35866 206159 35869
rect 165540 35864 206159 35866
rect 165540 35808 206098 35864
rect 206154 35808 206159 35864
rect 165540 35806 206159 35808
rect 165540 35804 165546 35806
rect 206093 35803 206159 35806
rect 145414 35124 145420 35188
rect 145484 35186 145490 35188
rect 170397 35186 170463 35189
rect 145484 35184 170463 35186
rect 145484 35128 170402 35184
rect 170458 35128 170463 35184
rect 145484 35126 170463 35128
rect 145484 35124 145490 35126
rect 170397 35123 170463 35126
rect 206093 35186 206159 35189
rect 425053 35186 425119 35189
rect 206093 35184 425119 35186
rect 206093 35128 206098 35184
rect 206154 35128 425058 35184
rect 425114 35128 425119 35184
rect 206093 35126 425119 35128
rect 206093 35123 206159 35126
rect 425053 35123 425119 35126
rect 580441 33146 580507 33149
rect 583520 33146 584960 33236
rect 580441 33144 584960 33146
rect 580441 33088 580446 33144
rect 580502 33088 584960 33144
rect 580441 33086 584960 33088
rect 580441 33083 580507 33086
rect 583520 32996 584960 33086
rect -960 32466 480 32556
rect -960 32406 674 32466
rect -960 32330 480 32406
rect 614 32330 674 32406
rect -960 32316 674 32330
rect 246 32270 674 32316
rect 246 31786 306 32270
rect 120574 31786 120580 31788
rect 246 31726 120580 31786
rect 120574 31724 120580 31726
rect 120644 31724 120650 31788
rect 157006 28868 157012 28932
rect 157076 28930 157082 28932
rect 211245 28930 211311 28933
rect 212441 28930 212507 28933
rect 157076 28928 212507 28930
rect 157076 28872 211250 28928
rect 211306 28872 212446 28928
rect 212502 28872 212507 28928
rect 157076 28870 212507 28872
rect 157076 28868 157082 28870
rect 211245 28867 211311 28870
rect 212441 28867 212507 28870
rect 144310 28188 144316 28252
rect 144380 28250 144386 28252
rect 157977 28250 158043 28253
rect 144380 28248 158043 28250
rect 144380 28192 157982 28248
rect 158038 28192 158043 28248
rect 144380 28190 158043 28192
rect 144380 28188 144386 28190
rect 157977 28187 158043 28190
rect 212441 28250 212507 28253
rect 307017 28250 307083 28253
rect 212441 28248 307083 28250
rect 212441 28192 212446 28248
rect 212502 28192 307022 28248
rect 307078 28192 307083 28248
rect 212441 28190 307083 28192
rect 212441 28187 212507 28190
rect 307017 28187 307083 28190
rect 157190 24788 157196 24852
rect 157260 24850 157266 24852
rect 210049 24850 210115 24853
rect 211061 24850 211127 24853
rect 157260 24848 211127 24850
rect 157260 24792 210054 24848
rect 210110 24792 211066 24848
rect 211122 24792 211127 24848
rect 157260 24790 211127 24792
rect 157260 24788 157266 24790
rect 210049 24787 210115 24790
rect 211061 24787 211127 24790
rect 211061 24170 211127 24173
rect 310513 24170 310579 24173
rect 211061 24168 310579 24170
rect 211061 24112 211066 24168
rect 211122 24112 310518 24168
rect 310574 24112 310579 24168
rect 211061 24110 310579 24112
rect 211061 24107 211127 24110
rect 310513 24107 310579 24110
rect 158478 21932 158484 21996
rect 158548 21994 158554 21996
rect 212533 21994 212599 21997
rect 213821 21994 213887 21997
rect 158548 21992 213887 21994
rect 158548 21936 212538 21992
rect 212594 21936 213826 21992
rect 213882 21936 213887 21992
rect 158548 21934 213887 21936
rect 158548 21932 158554 21934
rect 212533 21931 212599 21934
rect 213821 21931 213887 21934
rect 158294 21796 158300 21860
rect 158364 21858 158370 21860
rect 158364 21798 200130 21858
rect 158364 21796 158370 21798
rect 200070 21450 200130 21798
rect 211153 21450 211219 21453
rect 329097 21450 329163 21453
rect 200070 21448 329163 21450
rect 200070 21392 211158 21448
rect 211214 21392 329102 21448
rect 329158 21392 329163 21448
rect 200070 21390 329163 21392
rect 211153 21387 211219 21390
rect 329097 21387 329163 21390
rect 213821 21314 213887 21317
rect 336733 21314 336799 21317
rect 213821 21312 336799 21314
rect 213821 21256 213826 21312
rect 213882 21256 336738 21312
rect 336794 21256 336799 21312
rect 213821 21254 336799 21256
rect 213821 21251 213887 21254
rect 336733 21251 336799 21254
rect 155718 20572 155724 20636
rect 155788 20634 155794 20636
rect 209773 20634 209839 20637
rect 211061 20634 211127 20637
rect 155788 20632 211127 20634
rect 155788 20576 209778 20632
rect 209834 20576 211066 20632
rect 211122 20576 211127 20632
rect 155788 20574 211127 20576
rect 155788 20572 155794 20574
rect 209773 20571 209839 20574
rect 211061 20571 211127 20574
rect 211061 19954 211127 19957
rect 293953 19954 294019 19957
rect 211061 19952 294019 19954
rect 211061 19896 211066 19952
rect 211122 19896 293958 19952
rect 294014 19896 294019 19952
rect 211061 19894 294019 19896
rect 211061 19891 211127 19894
rect 293953 19891 294019 19894
rect 580349 19818 580415 19821
rect 583520 19818 584960 19908
rect 580349 19816 584960 19818
rect 580349 19760 580354 19816
rect 580410 19760 584960 19816
rect 580349 19758 584960 19760
rect 580349 19755 580415 19758
rect 583520 19668 584960 19758
rect -960 19410 480 19500
rect 3417 19410 3483 19413
rect -960 19408 3483 19410
rect -960 19352 3422 19408
rect 3478 19352 3483 19408
rect -960 19350 3483 19352
rect -960 19260 480 19350
rect 3417 19347 3483 19350
rect 144126 10236 144132 10300
rect 144196 10298 144202 10300
rect 157793 10298 157859 10301
rect 144196 10296 157859 10298
rect 144196 10240 157798 10296
rect 157854 10240 157859 10296
rect 144196 10238 157859 10240
rect 144196 10236 144202 10238
rect 157793 10235 157859 10238
rect 148174 8876 148180 8940
rect 148244 8938 148250 8940
rect 213361 8938 213427 8941
rect 148244 8936 213427 8938
rect 148244 8880 213366 8936
rect 213422 8880 213427 8936
rect 148244 8878 213427 8880
rect 148244 8876 148250 8878
rect 213361 8875 213427 8878
rect 580257 6626 580323 6629
rect 583520 6626 584960 6716
rect 580257 6624 584960 6626
rect -960 6490 480 6580
rect 580257 6568 580262 6624
rect 580318 6568 584960 6624
rect 580257 6566 584960 6568
rect 580257 6563 580323 6566
rect 3417 6490 3483 6493
rect -960 6488 3483 6490
rect -960 6432 3422 6488
rect 3478 6432 3483 6488
rect 583520 6476 584960 6566
rect -960 6430 3483 6432
rect -960 6340 480 6430
rect 3417 6427 3483 6430
<< via3 >>
rect 187740 278020 187804 278084
rect 187740 277476 187804 277540
rect 111564 265100 111628 265164
rect 192156 265100 192220 265164
rect 108804 264964 108868 265028
rect 196388 264964 196452 265028
rect 116900 263740 116964 263804
rect 113036 263604 113100 263668
rect 111196 263060 111260 263124
rect 191788 263060 191852 263124
rect 111012 262924 111076 262988
rect 112852 262788 112916 262852
rect 115796 262652 115860 262716
rect 193628 262652 193692 262716
rect 114140 262516 114204 262580
rect 111380 262380 111444 262444
rect 190500 262380 190564 262444
rect 191788 262380 191852 262444
rect 192340 262244 192404 262308
rect 112668 261020 112732 261084
rect 193444 260884 193508 260948
rect 122788 260748 122852 260812
rect 116716 260476 116780 260540
rect 115612 260340 115676 260404
rect 121132 260204 121196 260268
rect 116532 260068 116596 260132
rect 121316 259932 121380 259996
rect 118188 259796 118252 259860
rect 189028 259796 189092 259860
rect 113956 259524 114020 259588
rect 189212 259660 189276 259724
rect 124076 259524 124140 259588
rect 122972 259388 123036 259452
rect 186084 259388 186148 259452
rect 186084 213828 186148 213892
rect 131620 201452 131684 201516
rect 139532 201452 139596 201516
rect 154620 200636 154684 200700
rect 173572 200636 173636 200700
rect 150940 200500 151004 200564
rect 163084 200500 163148 200564
rect 106780 200364 106844 200428
rect 122788 200092 122852 200156
rect 132724 199858 132728 199884
rect 132728 199858 132784 199884
rect 132784 199858 132788 199884
rect 132724 199820 132788 199858
rect 133828 199880 133892 199884
rect 133828 199824 133832 199880
rect 133832 199824 133888 199880
rect 133888 199824 133892 199880
rect 133828 199820 133892 199824
rect 134748 199820 134812 199884
rect 133644 199722 133648 199748
rect 133648 199722 133704 199748
rect 133704 199722 133708 199748
rect 133644 199684 133708 199722
rect 171180 200364 171244 200428
rect 135484 199880 135548 199884
rect 135484 199824 135488 199880
rect 135488 199824 135544 199880
rect 135544 199824 135548 199880
rect 135484 199820 135548 199824
rect 135852 199858 135856 199884
rect 135856 199858 135912 199884
rect 135912 199858 135916 199884
rect 135852 199820 135916 199858
rect 142292 200092 142356 200156
rect 150020 200092 150084 200156
rect 137140 199744 137204 199748
rect 137140 199688 137144 199744
rect 137144 199688 137200 199744
rect 137200 199688 137204 199744
rect 137140 199684 137204 199688
rect 138244 199820 138308 199884
rect 137876 199684 137940 199748
rect 139532 199684 139596 199748
rect 139532 199548 139596 199612
rect 141556 199858 141560 199884
rect 141560 199858 141616 199884
rect 141616 199858 141620 199884
rect 141556 199820 141620 199858
rect 142108 199858 142112 199884
rect 142112 199858 142168 199884
rect 142168 199858 142172 199884
rect 142108 199820 142172 199858
rect 141740 199684 141804 199748
rect 142660 199820 142724 199884
rect 143212 199820 143276 199884
rect 143396 199820 143460 199884
rect 142476 199548 142540 199612
rect 143028 199684 143092 199748
rect 146156 199820 146220 199884
rect 147444 199548 147508 199612
rect 151860 199858 151864 199884
rect 151864 199858 151920 199884
rect 151920 199858 151924 199884
rect 151860 199820 151924 199858
rect 150940 199548 151004 199612
rect 117084 199412 117148 199476
rect 154620 199820 154684 199884
rect 157380 199858 157384 199884
rect 157384 199858 157440 199884
rect 157440 199858 157444 199884
rect 157380 199820 157444 199858
rect 159036 199820 159100 199884
rect 135162 199004 135226 199068
rect 137140 199004 137204 199068
rect 141556 199200 141620 199204
rect 141556 199144 141570 199200
rect 141570 199144 141620 199200
rect 141556 199140 141620 199144
rect 141740 199200 141804 199204
rect 141740 199144 141754 199200
rect 141754 199144 141804 199200
rect 141740 199140 141804 199144
rect 142108 199200 142172 199204
rect 142108 199144 142158 199200
rect 142158 199144 142172 199200
rect 142108 199140 142172 199144
rect 143212 199140 143276 199204
rect 156828 199412 156892 199476
rect 161060 199820 161124 199884
rect 162164 199858 162168 199884
rect 162168 199858 162224 199884
rect 162224 199858 162228 199884
rect 162164 199820 162228 199858
rect 162532 199820 162596 199884
rect 163084 199744 163148 199748
rect 163084 199688 163134 199744
rect 163134 199688 163148 199744
rect 163084 199684 163148 199688
rect 164188 199880 164252 199884
rect 164188 199824 164192 199880
rect 164192 199824 164248 199880
rect 164248 199824 164252 199880
rect 164188 199820 164252 199824
rect 166764 199858 166768 199884
rect 166768 199858 166824 199884
rect 166824 199858 166828 199884
rect 166764 199820 166828 199858
rect 166212 199684 166276 199748
rect 169708 199684 169772 199748
rect 172284 200092 172348 200156
rect 172836 200092 172900 200156
rect 170444 199820 170508 199884
rect 170812 199820 170876 199884
rect 171180 199548 171244 199612
rect 172652 199684 172716 199748
rect 173572 199820 173636 199884
rect 173756 199880 173820 199884
rect 173756 199824 173760 199880
rect 173760 199824 173816 199880
rect 173816 199824 173820 199880
rect 173756 199820 173820 199824
rect 174124 199858 174128 199884
rect 174128 199858 174184 199884
rect 174184 199858 174188 199884
rect 174124 199820 174188 199858
rect 173388 199684 173452 199748
rect 175228 199820 175292 199884
rect 176700 199956 176764 200020
rect 176148 199820 176212 199884
rect 177436 199880 177500 199884
rect 177436 199824 177486 199880
rect 177486 199824 177500 199880
rect 177436 199820 177500 199824
rect 173572 199548 173636 199612
rect 175044 199684 175108 199748
rect 200804 199276 200868 199340
rect 198964 199140 199028 199204
rect 151860 199004 151924 199068
rect 173756 199004 173820 199068
rect 200620 199004 200684 199068
rect 176148 198868 176212 198932
rect 122972 198732 123036 198796
rect 143580 198596 143644 198660
rect 144316 198596 144380 198660
rect 148732 198596 148796 198660
rect 170996 198656 171060 198660
rect 174124 198732 174188 198796
rect 201540 198868 201604 198932
rect 177068 198732 177132 198796
rect 177436 198792 177500 198796
rect 177436 198736 177450 198792
rect 177450 198736 177500 198792
rect 177436 198732 177500 198736
rect 170996 198600 171010 198656
rect 171010 198600 171060 198656
rect 170996 198596 171060 198600
rect 196020 198596 196084 198660
rect 135116 198460 135180 198524
rect 142660 198460 142724 198524
rect 143028 198460 143092 198524
rect 143396 198520 143460 198524
rect 143396 198464 143410 198520
rect 143410 198464 143460 198520
rect 143396 198460 143460 198464
rect 146156 198460 146220 198524
rect 165476 198460 165540 198524
rect 193260 198460 193324 198524
rect 107516 198324 107580 198388
rect 148916 198324 148980 198388
rect 158484 198324 158548 198388
rect 173572 198324 173636 198388
rect 107332 198188 107396 198252
rect 146892 198188 146956 198252
rect 157380 198248 157444 198252
rect 157380 198192 157394 198248
rect 157394 198192 157444 198248
rect 157380 198188 157444 198192
rect 162348 198248 162412 198252
rect 162348 198192 162362 198248
rect 162362 198192 162412 198248
rect 162348 198188 162412 198192
rect 170444 198248 170508 198252
rect 170444 198192 170494 198248
rect 170494 198192 170508 198248
rect 170444 198188 170508 198192
rect 197308 198324 197372 198388
rect 136772 198052 136836 198116
rect 138796 198052 138860 198116
rect 149652 198112 149716 198116
rect 149652 198056 149666 198112
rect 149666 198056 149716 198112
rect 149652 198052 149716 198056
rect 149836 198052 149900 198116
rect 152964 198052 153028 198116
rect 154436 198052 154500 198116
rect 156644 198052 156708 198116
rect 157196 198112 157260 198116
rect 157196 198056 157246 198112
rect 157246 198056 157260 198112
rect 157196 198052 157260 198056
rect 166764 198112 166828 198116
rect 166764 198056 166778 198112
rect 166778 198056 166828 198112
rect 166764 198052 166828 198056
rect 199148 198188 199212 198252
rect 196204 198052 196268 198116
rect 133644 197916 133708 197980
rect 166212 197916 166276 197980
rect 135300 197644 135364 197708
rect 147260 197644 147324 197708
rect 162532 197780 162596 197844
rect 172836 197780 172900 197844
rect 191972 197780 192036 197844
rect 135484 197508 135548 197572
rect 142108 197508 142172 197572
rect 147076 197508 147140 197572
rect 134012 197372 134076 197436
rect 143948 197372 144012 197436
rect 198780 197236 198844 197300
rect 147444 197100 147508 197164
rect 164188 197100 164252 197164
rect 147444 196964 147508 197028
rect 108252 196828 108316 196892
rect 162164 196888 162228 196892
rect 162164 196832 162214 196888
rect 162214 196832 162228 196888
rect 162164 196828 162228 196832
rect 136588 196692 136652 196756
rect 139348 196692 139412 196756
rect 143764 196692 143828 196756
rect 137876 196556 137940 196620
rect 169708 196480 169772 196484
rect 169708 196424 169722 196480
rect 169722 196424 169772 196480
rect 169708 196420 169772 196424
rect 170812 196420 170876 196484
rect 172284 196420 172348 196484
rect 173756 196420 173820 196484
rect 169524 196284 169588 196348
rect 134748 195876 134812 195940
rect 169340 195876 169404 195940
rect 193812 195876 193876 195940
rect 157196 195740 157260 195804
rect 100340 195604 100404 195668
rect 173388 195604 173452 195668
rect 201724 195604 201788 195668
rect 118372 195468 118436 195532
rect 156644 195468 156708 195532
rect 119844 195196 119908 195260
rect 133828 195196 133892 195260
rect 138428 195196 138492 195260
rect 191788 195196 191852 195260
rect 138060 195060 138124 195124
rect 194548 195060 194612 195124
rect 203012 194244 203076 194308
rect 159036 193972 159100 194036
rect 209820 193972 209884 194036
rect 100524 193836 100588 193900
rect 168236 193292 168300 193356
rect 187004 193156 187068 193220
rect 147444 193020 147508 193084
rect 172468 193020 172532 193084
rect 205588 193020 205652 193084
rect 103284 192884 103348 192948
rect 133828 192884 133892 192948
rect 161060 192884 161124 192948
rect 104020 192748 104084 192812
rect 170444 192748 170508 192812
rect 144316 192612 144380 192676
rect 124812 192476 124876 192540
rect 170996 192476 171060 192540
rect 187924 192340 187988 192404
rect 109540 191660 109604 191724
rect 138796 191660 138860 191724
rect 133828 191524 133892 191588
rect 118556 191388 118620 191452
rect 135484 191252 135548 191316
rect 134012 191116 134076 191180
rect 135300 190980 135364 191044
rect 186084 190980 186148 191044
rect 138428 190164 138492 190228
rect 142292 190028 142356 190092
rect 181300 190028 181364 190092
rect 143948 189892 144012 189956
rect 176516 189892 176580 189956
rect 210004 189892 210068 189956
rect 142476 189756 142540 189820
rect 174860 189756 174924 189820
rect 143764 189620 143828 189684
rect 154436 189620 154500 189684
rect 142108 187580 142172 187644
rect 108436 187444 108500 187508
rect 138244 187308 138308 187372
rect 175044 187308 175108 187372
rect 139532 187172 139596 187236
rect 152964 187172 153028 187236
rect 138060 187036 138124 187100
rect 149836 187036 149900 187100
rect 132540 186900 132604 186964
rect 149652 186900 149716 186964
rect 148732 159292 148796 159356
rect 168236 156844 168300 156908
rect 169340 156708 169404 156772
rect 203012 156708 203076 156772
rect 203196 156572 203260 156636
rect 211292 153852 211356 153916
rect 211108 153716 211172 153780
rect 177068 151404 177132 151468
rect 207060 151404 207124 151468
rect 205956 151268 206020 151332
rect 122420 151132 122484 151196
rect 139348 151132 139412 151196
rect 207244 151132 207308 151196
rect 122972 150996 123036 151060
rect 148916 150996 148980 151060
rect 124076 150452 124140 150516
rect 188292 149908 188356 149972
rect 189396 149772 189460 149836
rect 156828 149636 156892 149700
rect 197860 149092 197924 149156
rect 200988 149152 201052 149156
rect 200988 149096 201038 149152
rect 201038 149096 201052 149152
rect 200988 149092 201052 149096
rect 197492 148956 197556 149020
rect 201908 148820 201972 148884
rect 173756 148684 173820 148748
rect 103100 148548 103164 148612
rect 170628 148548 170692 148612
rect 203380 148548 203444 148612
rect 104204 148412 104268 148476
rect 136772 148412 136836 148476
rect 205772 148412 205836 148476
rect 119660 148276 119724 148340
rect 158484 148276 158548 148340
rect 194732 148140 194796 148204
rect 112484 147460 112548 147524
rect 131620 147460 131684 147524
rect 196572 147460 196636 147524
rect 113588 147324 113652 147388
rect 115060 147188 115124 147252
rect 150020 147188 150084 147252
rect 122052 147052 122116 147116
rect 147260 147052 147324 147116
rect 136588 146916 136652 146980
rect 115796 146236 115860 146300
rect 189764 146100 189828 146164
rect 120764 145964 120828 146028
rect 191604 145964 191668 146028
rect 111012 145828 111076 145892
rect 112852 145828 112916 145892
rect 187372 145828 187436 145892
rect 112116 145692 112180 145756
rect 196388 145692 196452 145756
rect 115796 145556 115860 145620
rect 192340 145556 192404 145620
rect 113036 144740 113100 144804
rect 115612 144740 115676 144804
rect 116532 144740 116596 144804
rect 193628 144740 193692 144804
rect 111564 144604 111628 144668
rect 162348 144604 162412 144668
rect 114140 144468 114204 144532
rect 190500 144468 190564 144532
rect 112668 144332 112732 144396
rect 147076 144196 147140 144260
rect 143580 144060 143644 144124
rect 118188 143984 118252 143988
rect 118188 143928 118202 143984
rect 118202 143928 118252 143984
rect 118188 143924 118252 143928
rect 116900 143788 116964 143852
rect 116716 143380 116780 143444
rect 192340 143380 192404 143444
rect 113956 143244 114020 143308
rect 111196 143108 111260 143172
rect 121132 142972 121196 143036
rect 121316 142836 121380 142900
rect 187740 142836 187804 142900
rect 116532 142292 116596 142356
rect 111012 142156 111076 142220
rect 111380 142020 111444 142084
rect 189212 142020 189276 142084
rect 114140 141884 114204 141948
rect 108804 141748 108868 141812
rect 192156 141748 192220 141812
rect 121132 141612 121196 141676
rect 189028 141612 189092 141676
rect 116716 141476 116780 141540
rect 165476 141476 165540 141540
rect 117820 141340 117884 141404
rect 190500 141340 190564 141404
rect 113772 141204 113836 141268
rect 191052 140660 191116 140724
rect 193444 140720 193508 140724
rect 193444 140664 193494 140720
rect 193494 140664 193508 140720
rect 193444 140660 193508 140664
rect 119476 140524 119540 140588
rect 189580 140524 189644 140588
rect 120948 140388 121012 140452
rect 193444 140388 193508 140452
rect 115612 140252 115676 140316
rect 193628 140252 193692 140316
rect 112300 140116 112364 140180
rect 185348 140176 185412 140180
rect 185348 140120 185398 140176
rect 185398 140120 185412 140176
rect 185348 140116 185412 140120
rect 192156 140116 192220 140180
rect 122604 139980 122668 140044
rect 128860 140040 128924 140044
rect 128860 139984 128910 140040
rect 128910 139984 128924 140040
rect 128860 139980 128924 139984
rect 130332 140040 130396 140044
rect 130332 139984 130382 140040
rect 130382 139984 130396 140040
rect 130332 139980 130396 139984
rect 120580 139844 120644 139908
rect 190684 139980 190748 140044
rect 187188 139844 187252 139908
rect 188108 139708 188172 139772
rect 187740 139632 187804 139636
rect 187740 139576 187754 139632
rect 187754 139576 187804 139632
rect 118740 139436 118804 139500
rect 187740 139572 187804 139576
rect 111564 139300 111628 139364
rect 123156 139300 123220 139364
rect 111196 139028 111260 139092
rect 130332 138756 130396 138820
rect 185900 139300 185964 139364
rect 202092 139436 202156 139500
rect 185348 139028 185412 139092
rect 186268 138892 186332 138956
rect 146892 138620 146956 138684
rect 169708 138620 169772 138684
rect 201172 138620 201236 138684
rect 122236 138484 122300 138548
rect 128860 138484 128924 138548
rect 116900 137940 116964 138004
rect 122420 138076 122484 138140
rect 186452 138076 186516 138140
rect 187740 138076 187804 138140
rect 122420 137940 122484 138004
rect 124812 137940 124876 138004
rect 181300 137940 181364 138004
rect 185900 137804 185964 137868
rect 118188 137396 118252 137460
rect 122052 137396 122116 137460
rect 112852 137260 112916 137324
rect 122972 137260 123036 137324
rect 186268 135900 186332 135964
rect 122972 133860 123036 133924
rect 186084 131684 186148 131748
rect 186268 131412 186332 131476
rect 186084 117948 186148 118012
rect 186268 104892 186332 104956
rect 186636 104892 186700 104956
rect 118740 96596 118804 96660
rect 186636 90340 186700 90404
rect 189028 90340 189092 90404
rect 186084 86260 186148 86324
rect 186636 86260 186700 86324
rect 122972 86124 123036 86188
rect 122972 85988 123036 86052
rect 117820 84220 117884 84284
rect 186084 82180 186148 82244
rect 186268 82044 186332 82108
rect 112116 81772 112180 81836
rect 124076 81772 124140 81836
rect 184060 81772 184124 81836
rect 185348 81636 185412 81700
rect 186636 81636 186700 81700
rect 178908 81500 178972 81564
rect 189580 81500 189644 81564
rect 196572 81500 196636 81564
rect 175044 81228 175108 81292
rect 197492 81228 197556 81292
rect 146340 81092 146404 81156
rect 175596 81092 175660 81156
rect 205956 81092 206020 81156
rect 149284 80956 149348 81020
rect 177252 80956 177316 81020
rect 148732 80820 148796 80884
rect 197308 80684 197372 80748
rect 118188 80140 118252 80204
rect 146524 80140 146588 80204
rect 155724 80140 155788 80204
rect 159036 80004 159100 80068
rect 134012 79868 134076 79932
rect 133276 79732 133340 79796
rect 133828 79732 133892 79796
rect 135116 79928 135180 79932
rect 135116 79872 135120 79928
rect 135120 79872 135176 79928
rect 135176 79872 135180 79928
rect 135116 79868 135180 79872
rect 135484 79868 135548 79932
rect 136036 79868 136100 79932
rect 137508 79868 137572 79932
rect 137692 79928 137756 79932
rect 137692 79872 137696 79928
rect 137696 79872 137752 79928
rect 137752 79872 137756 79928
rect 137692 79868 137756 79872
rect 138060 79928 138124 79932
rect 138060 79872 138064 79928
rect 138064 79872 138120 79928
rect 138120 79872 138124 79928
rect 138060 79868 138124 79872
rect 138428 79868 138492 79932
rect 139164 79868 139228 79932
rect 139900 79868 139964 79932
rect 135668 79732 135732 79796
rect 138244 79732 138308 79796
rect 139900 79732 139964 79796
rect 136588 79596 136652 79660
rect 140268 79792 140332 79796
rect 140268 79736 140272 79792
rect 140272 79736 140328 79792
rect 140328 79736 140332 79792
rect 140268 79732 140332 79736
rect 141556 79928 141620 79932
rect 141556 79872 141560 79928
rect 141560 79872 141616 79928
rect 141616 79872 141620 79928
rect 141556 79868 141620 79872
rect 140820 79792 140884 79796
rect 140820 79736 140870 79792
rect 140870 79736 140884 79792
rect 140820 79732 140884 79736
rect 142660 79868 142724 79932
rect 142108 79732 142172 79796
rect 144132 79868 144196 79932
rect 143580 79792 143644 79796
rect 143580 79736 143584 79792
rect 143584 79736 143640 79792
rect 143640 79736 143644 79792
rect 143580 79732 143644 79736
rect 141004 79596 141068 79660
rect 145604 79868 145668 79932
rect 146892 79868 146956 79932
rect 147076 79732 147140 79796
rect 147628 79928 147692 79932
rect 147628 79872 147632 79928
rect 147632 79872 147688 79928
rect 147688 79872 147692 79928
rect 147628 79868 147692 79872
rect 148732 79868 148796 79932
rect 149284 79868 149348 79932
rect 149836 79868 149900 79932
rect 147996 79732 148060 79796
rect 149652 79596 149716 79660
rect 151676 79928 151740 79932
rect 151676 79872 151680 79928
rect 151680 79872 151736 79928
rect 151736 79872 151740 79928
rect 151676 79868 151740 79872
rect 153148 79868 153212 79932
rect 146340 79460 146404 79524
rect 152596 79596 152660 79660
rect 154436 79868 154500 79932
rect 154988 79868 155052 79932
rect 155908 79868 155972 79932
rect 153884 79460 153948 79524
rect 156644 79868 156708 79932
rect 156828 79732 156892 79796
rect 157196 79596 157260 79660
rect 158116 79868 158180 79932
rect 158484 79868 158548 79932
rect 159404 79868 159468 79932
rect 161060 79868 161124 79932
rect 161980 79928 162044 79932
rect 161980 79872 161984 79928
rect 161984 79872 162040 79928
rect 162040 79872 162044 79928
rect 161980 79868 162044 79872
rect 162348 79906 162352 79932
rect 162352 79906 162408 79932
rect 162408 79906 162412 79932
rect 162348 79868 162412 79906
rect 162900 79868 162964 79932
rect 158668 79732 158732 79796
rect 161244 79732 161308 79796
rect 162716 79732 162780 79796
rect 163084 79732 163148 79796
rect 163452 79792 163516 79796
rect 163452 79736 163466 79792
rect 163466 79736 163516 79792
rect 163452 79732 163516 79736
rect 162164 79596 162228 79660
rect 163268 79596 163332 79660
rect 166212 79868 166276 79932
rect 166580 79868 166644 79932
rect 165292 79792 165356 79796
rect 165292 79736 165296 79792
rect 165296 79736 165352 79792
rect 165352 79736 165356 79792
rect 165292 79732 165356 79736
rect 165476 79792 165540 79796
rect 165476 79736 165480 79792
rect 165480 79736 165536 79792
rect 165536 79736 165540 79792
rect 165476 79732 165540 79736
rect 165108 79596 165172 79660
rect 167316 79732 167380 79796
rect 167868 79732 167932 79796
rect 169524 80004 169588 80068
rect 170812 80140 170876 80204
rect 192340 80412 192404 80476
rect 177252 80276 177316 80340
rect 184244 80276 184308 80340
rect 173572 80004 173636 80068
rect 169340 79928 169404 79932
rect 169340 79872 169344 79928
rect 169344 79872 169400 79928
rect 169400 79872 169404 79928
rect 169340 79868 169404 79872
rect 170628 79868 170692 79932
rect 170628 79732 170692 79796
rect 172100 79868 172164 79932
rect 173204 79928 173268 79932
rect 173204 79872 173208 79928
rect 173208 79872 173264 79928
rect 173264 79872 173268 79928
rect 173204 79868 173268 79872
rect 186452 80140 186516 80204
rect 185532 80004 185596 80068
rect 186268 80004 186332 80068
rect 200804 80004 200868 80068
rect 173940 79868 174004 79932
rect 172284 79732 172348 79796
rect 173756 79732 173820 79796
rect 166396 79596 166460 79660
rect 166764 79596 166828 79660
rect 167684 79596 167748 79660
rect 170996 79656 171060 79660
rect 170996 79600 171010 79656
rect 171010 79600 171060 79656
rect 170996 79596 171060 79600
rect 172100 79596 172164 79660
rect 174492 79792 174556 79796
rect 174492 79736 174542 79792
rect 174542 79736 174556 79792
rect 174492 79732 174556 79736
rect 174860 79732 174924 79796
rect 175780 79906 175784 79932
rect 175784 79906 175840 79932
rect 175840 79906 175844 79932
rect 175780 79868 175844 79906
rect 176516 79868 176580 79932
rect 185348 79868 185412 79932
rect 174860 79596 174924 79660
rect 175596 79596 175660 79660
rect 175964 79596 176028 79660
rect 185348 79596 185412 79660
rect 148732 79324 148796 79388
rect 149100 79324 149164 79388
rect 170628 79324 170692 79388
rect 171916 79324 171980 79388
rect 175044 79324 175108 79388
rect 193812 79324 193876 79388
rect 152780 79188 152844 79252
rect 120948 78916 121012 78980
rect 158116 78916 158180 78980
rect 187004 79188 187068 79252
rect 191052 79052 191116 79116
rect 187924 78916 187988 78980
rect 119476 78644 119540 78708
rect 142660 78704 142724 78708
rect 142660 78648 142674 78704
rect 142674 78648 142724 78704
rect 142660 78644 142724 78648
rect 146892 78644 146956 78708
rect 152412 78644 152476 78708
rect 159404 78644 159468 78708
rect 160692 78704 160756 78708
rect 160692 78648 160706 78704
rect 160706 78648 160756 78704
rect 160692 78644 160756 78648
rect 160876 78704 160940 78708
rect 160876 78648 160926 78704
rect 160926 78648 160940 78704
rect 160876 78644 160940 78648
rect 171732 78644 171796 78708
rect 171916 78644 171980 78708
rect 187372 78644 187436 78708
rect 119844 78508 119908 78572
rect 149284 78508 149348 78572
rect 157012 78508 157076 78572
rect 158852 78508 158916 78572
rect 170628 78508 170692 78572
rect 141556 78372 141620 78436
rect 175596 78372 175660 78436
rect 211292 78372 211356 78436
rect 102180 78100 102244 78164
rect 162348 78236 162412 78300
rect 175044 78236 175108 78300
rect 176148 78236 176212 78300
rect 154988 78100 155052 78164
rect 173204 78100 173268 78164
rect 190684 78236 190748 78300
rect 211108 78100 211172 78164
rect 134380 77964 134444 78028
rect 163084 77964 163148 78028
rect 167316 77964 167380 78028
rect 167868 77964 167932 78028
rect 143948 77828 144012 77892
rect 163452 77828 163516 77892
rect 163636 77828 163700 77892
rect 178908 77964 178972 78028
rect 143580 77692 143644 77756
rect 163452 77692 163516 77756
rect 175964 77556 176028 77620
rect 107332 77420 107396 77484
rect 142108 77420 142172 77484
rect 148916 77420 148980 77484
rect 154436 77420 154500 77484
rect 175780 77480 175844 77484
rect 175780 77424 175794 77480
rect 175794 77424 175844 77480
rect 175780 77420 175844 77424
rect 102180 77284 102244 77348
rect 103284 77284 103348 77348
rect 147812 77284 147876 77348
rect 150020 77284 150084 77348
rect 151124 77284 151188 77348
rect 152596 77284 152660 77348
rect 148364 77148 148428 77212
rect 154068 77284 154132 77348
rect 155540 77284 155604 77348
rect 161980 77284 162044 77348
rect 162348 77284 162412 77348
rect 162532 77344 162596 77348
rect 162532 77288 162546 77344
rect 162546 77288 162596 77344
rect 162532 77284 162596 77288
rect 162900 77284 162964 77348
rect 164740 77284 164804 77348
rect 167500 77284 167564 77348
rect 175964 77284 176028 77348
rect 135300 77012 135364 77076
rect 138060 77012 138124 77076
rect 138612 77012 138676 77076
rect 155908 76876 155972 76940
rect 113772 76740 113836 76804
rect 193628 76740 193692 76804
rect 133460 76604 133524 76668
rect 134196 76604 134260 76668
rect 138060 76604 138124 76668
rect 139164 76604 139228 76668
rect 139348 76604 139412 76668
rect 143580 76604 143644 76668
rect 145604 76604 145668 76668
rect 146708 76604 146772 76668
rect 194732 76604 194796 76668
rect 139532 76468 139596 76532
rect 140268 76468 140332 76532
rect 173940 76332 174004 76396
rect 135116 75788 135180 75852
rect 205588 75788 205652 75852
rect 137692 75652 137756 75716
rect 170996 75652 171060 75716
rect 191604 75516 191668 75580
rect 189764 75380 189828 75444
rect 188292 75244 188356 75308
rect 119844 75108 119908 75172
rect 189396 75108 189460 75172
rect 136036 74700 136100 74764
rect 143764 74700 143828 74764
rect 133092 74564 133156 74628
rect 118372 74428 118436 74492
rect 122236 74292 122300 74356
rect 147076 74156 147140 74220
rect 149652 74156 149716 74220
rect 106780 74080 106844 74084
rect 106780 74024 106830 74080
rect 106830 74024 106844 74080
rect 106780 74020 106844 74024
rect 153148 74020 153212 74084
rect 113588 73884 113652 73948
rect 149468 73884 149532 73948
rect 162164 73748 162228 73812
rect 112300 73612 112364 73676
rect 193444 73612 193508 73676
rect 151124 73476 151188 73540
rect 151676 73340 151740 73404
rect 108252 73128 108316 73132
rect 108252 73072 108302 73128
rect 108302 73072 108316 73128
rect 108252 73068 108316 73072
rect 117084 73068 117148 73132
rect 158668 73068 158732 73132
rect 145420 72932 145484 72996
rect 148364 72796 148428 72860
rect 147444 72660 147508 72724
rect 201908 72660 201972 72724
rect 192156 72388 192220 72452
rect 188108 72252 188172 72316
rect 144132 71708 144196 71772
rect 115612 71436 115676 71500
rect 205772 71436 205836 71500
rect 196204 71300 196268 71364
rect 107516 71164 107580 71228
rect 205772 71164 205836 71228
rect 201724 71028 201788 71092
rect 185532 70348 185596 70412
rect 146524 70212 146588 70276
rect 120028 70076 120092 70140
rect 166212 70076 166276 70140
rect 120764 69940 120828 70004
rect 121132 69804 121196 69868
rect 190500 69940 190564 70004
rect 122604 69668 122668 69732
rect 146708 69532 146772 69596
rect 147260 69532 147324 69596
rect 200620 69532 200684 69596
rect 141004 68852 141068 68916
rect 149836 68852 149900 68916
rect 116716 68716 116780 68780
rect 189028 68716 189092 68780
rect 122420 68580 122484 68644
rect 185348 68580 185412 68644
rect 143948 68444 144012 68508
rect 144500 68444 144564 68508
rect 111564 68308 111628 68372
rect 145604 68172 145668 68236
rect 194548 68172 194612 68236
rect 143764 68036 143828 68100
rect 144316 68036 144380 68100
rect 143580 67492 143644 67556
rect 144684 67492 144748 67556
rect 114140 67356 114204 67420
rect 147812 67356 147876 67420
rect 148180 67356 148244 67420
rect 193260 67492 193324 67556
rect 201540 67492 201604 67556
rect 184244 67356 184308 67420
rect 147996 67220 148060 67284
rect 148364 67220 148428 67284
rect 186084 67220 186148 67284
rect 184060 67084 184124 67148
rect 150020 66948 150084 67012
rect 109540 66812 109604 66876
rect 148916 66812 148980 66876
rect 199148 66464 199212 66468
rect 199148 66408 199198 66464
rect 199198 66408 199212 66464
rect 199148 66404 199212 66408
rect 115796 66132 115860 66196
rect 196020 66132 196084 66196
rect 118556 65996 118620 66060
rect 164740 65996 164804 66060
rect 124076 65860 124140 65924
rect 108436 65588 108500 65652
rect 104020 65452 104084 65516
rect 198964 64832 199028 64836
rect 198964 64776 198978 64832
rect 198978 64776 199028 64832
rect 198964 64772 199028 64776
rect 171916 64636 171980 64700
rect 160692 64500 160756 64564
rect 152780 64364 152844 64428
rect 111196 64152 111260 64156
rect 111196 64096 111246 64152
rect 111246 64096 111260 64152
rect 111196 64092 111260 64096
rect 147444 64092 147508 64156
rect 100340 63412 100404 63476
rect 133460 63412 133524 63476
rect 187188 63472 187252 63476
rect 187188 63416 187238 63472
rect 187238 63416 187252 63472
rect 187188 63412 187252 63416
rect 115060 63336 115124 63340
rect 115060 63280 115110 63336
rect 115110 63280 115124 63336
rect 115060 63276 115124 63280
rect 167500 63276 167564 63340
rect 148548 62868 148612 62932
rect 100340 62732 100404 62796
rect 134380 62052 134444 62116
rect 167684 62052 167748 62116
rect 202092 62112 202156 62116
rect 202092 62056 202142 62112
rect 202142 62056 202156 62112
rect 138612 61916 138676 61980
rect 176148 61916 176212 61980
rect 202092 62052 202156 62056
rect 200988 61372 201052 61436
rect 133276 60556 133340 60620
rect 170628 60556 170692 60620
rect 138428 60420 138492 60484
rect 203380 59876 203444 59940
rect 111748 59196 111812 59260
rect 112852 59196 112916 59260
rect 139900 59196 139964 59260
rect 153884 59196 153948 59260
rect 112484 58788 112548 58852
rect 139716 59060 139780 59124
rect 162348 59060 162412 59124
rect 167868 58924 167932 58988
rect 172100 58788 172164 58852
rect 111748 58652 111812 58716
rect 140820 58516 140884 58580
rect 191972 58516 192036 58580
rect 111012 57972 111076 58036
rect 134196 57836 134260 57900
rect 158852 57836 158916 57900
rect 138244 57700 138308 57764
rect 165108 57700 165172 57764
rect 203196 57760 203260 57764
rect 203196 57704 203246 57760
rect 203246 57704 203260 57760
rect 197860 57564 197924 57628
rect 147260 57156 147324 57220
rect 203196 57700 203260 57704
rect 99420 56476 99484 56540
rect 100524 56476 100588 56540
rect 133092 56476 133156 56540
rect 170812 56476 170876 56540
rect 162532 56340 162596 56404
rect 154068 56204 154132 56268
rect 104204 55932 104268 55996
rect 168052 55932 168116 55996
rect 99420 55796 99484 55860
rect 138060 55116 138124 55180
rect 172284 55116 172348 55180
rect 137508 54980 137572 55044
rect 166396 54980 166460 55044
rect 160876 54844 160940 54908
rect 176332 54572 176396 54636
rect 209820 54436 209884 54500
rect 103100 53756 103164 53820
rect 135668 53756 135732 53820
rect 166580 53756 166644 53820
rect 139532 53620 139596 53684
rect 161060 53620 161124 53684
rect 169340 53484 169404 53548
rect 201172 53076 201236 53140
rect 163268 52396 163332 52460
rect 159036 52260 159100 52324
rect 156644 52124 156708 52188
rect 144684 51716 144748 51780
rect 174492 51716 174556 51780
rect 134012 50900 134076 50964
rect 152412 50900 152476 50964
rect 116900 50764 116964 50828
rect 139348 50764 139412 50828
rect 158116 50764 158180 50828
rect 191788 50764 191852 50828
rect 193076 50764 193140 50828
rect 175964 50628 176028 50692
rect 210004 50628 210068 50692
rect 211108 50628 211172 50692
rect 193076 50492 193140 50556
rect 161244 50356 161308 50420
rect 147076 50220 147140 50284
rect 211108 50220 211172 50284
rect 133828 49540 133892 49604
rect 174676 49540 174740 49604
rect 162716 49404 162780 49468
rect 171732 49268 171796 49332
rect 135484 48180 135548 48244
rect 203012 48240 203076 48244
rect 203012 48184 203062 48240
rect 203062 48184 203076 48240
rect 203012 48180 203076 48184
rect 163452 48044 163516 48108
rect 169524 47908 169588 47972
rect 202828 47908 202892 47972
rect 204116 47908 204180 47972
rect 204116 47636 204180 47700
rect 170444 47500 170508 47564
rect 135300 46820 135364 46884
rect 165292 46820 165356 46884
rect 198780 46820 198844 46884
rect 146892 46140 146956 46204
rect 207244 46548 207308 46612
rect 154252 45460 154316 45524
rect 166764 45324 166828 45388
rect 173572 45188 173636 45252
rect 173756 44916 173820 44980
rect 116532 44236 116596 44300
rect 136588 44100 136652 44164
rect 163636 44100 163700 44164
rect 207060 44160 207124 44164
rect 207060 44104 207074 44160
rect 207074 44104 207124 44160
rect 207060 44100 207124 44104
rect 156828 43964 156892 44028
rect 148364 43828 148428 43892
rect 174860 43420 174924 43484
rect 155540 42740 155604 42804
rect 154436 38524 154500 38588
rect 144500 37844 144564 37908
rect 175044 37164 175108 37228
rect 165476 35804 165540 35868
rect 145420 35124 145484 35188
rect 120580 31724 120644 31788
rect 157012 28868 157076 28932
rect 144316 28188 144380 28252
rect 157196 24788 157260 24852
rect 158484 21932 158548 21996
rect 158300 21796 158364 21860
rect 155724 20572 155788 20636
rect 144132 10236 144196 10300
rect 148180 8876 148244 8940
<< metal4 >>
rect -8726 711558 -8106 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 -8106 711558
rect -8726 711238 -8106 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 -8106 711238
rect -8726 682954 -8106 711002
rect -8726 682718 -8694 682954
rect -8458 682718 -8374 682954
rect -8138 682718 -8106 682954
rect -8726 682634 -8106 682718
rect -8726 682398 -8694 682634
rect -8458 682398 -8374 682634
rect -8138 682398 -8106 682634
rect -8726 646954 -8106 682398
rect -8726 646718 -8694 646954
rect -8458 646718 -8374 646954
rect -8138 646718 -8106 646954
rect -8726 646634 -8106 646718
rect -8726 646398 -8694 646634
rect -8458 646398 -8374 646634
rect -8138 646398 -8106 646634
rect -8726 610954 -8106 646398
rect -8726 610718 -8694 610954
rect -8458 610718 -8374 610954
rect -8138 610718 -8106 610954
rect -8726 610634 -8106 610718
rect -8726 610398 -8694 610634
rect -8458 610398 -8374 610634
rect -8138 610398 -8106 610634
rect -8726 574954 -8106 610398
rect -8726 574718 -8694 574954
rect -8458 574718 -8374 574954
rect -8138 574718 -8106 574954
rect -8726 574634 -8106 574718
rect -8726 574398 -8694 574634
rect -8458 574398 -8374 574634
rect -8138 574398 -8106 574634
rect -8726 538954 -8106 574398
rect -8726 538718 -8694 538954
rect -8458 538718 -8374 538954
rect -8138 538718 -8106 538954
rect -8726 538634 -8106 538718
rect -8726 538398 -8694 538634
rect -8458 538398 -8374 538634
rect -8138 538398 -8106 538634
rect -8726 502954 -8106 538398
rect -8726 502718 -8694 502954
rect -8458 502718 -8374 502954
rect -8138 502718 -8106 502954
rect -8726 502634 -8106 502718
rect -8726 502398 -8694 502634
rect -8458 502398 -8374 502634
rect -8138 502398 -8106 502634
rect -8726 466954 -8106 502398
rect -8726 466718 -8694 466954
rect -8458 466718 -8374 466954
rect -8138 466718 -8106 466954
rect -8726 466634 -8106 466718
rect -8726 466398 -8694 466634
rect -8458 466398 -8374 466634
rect -8138 466398 -8106 466634
rect -8726 430954 -8106 466398
rect -8726 430718 -8694 430954
rect -8458 430718 -8374 430954
rect -8138 430718 -8106 430954
rect -8726 430634 -8106 430718
rect -8726 430398 -8694 430634
rect -8458 430398 -8374 430634
rect -8138 430398 -8106 430634
rect -8726 394954 -8106 430398
rect -8726 394718 -8694 394954
rect -8458 394718 -8374 394954
rect -8138 394718 -8106 394954
rect -8726 394634 -8106 394718
rect -8726 394398 -8694 394634
rect -8458 394398 -8374 394634
rect -8138 394398 -8106 394634
rect -8726 358954 -8106 394398
rect -8726 358718 -8694 358954
rect -8458 358718 -8374 358954
rect -8138 358718 -8106 358954
rect -8726 358634 -8106 358718
rect -8726 358398 -8694 358634
rect -8458 358398 -8374 358634
rect -8138 358398 -8106 358634
rect -8726 322954 -8106 358398
rect -8726 322718 -8694 322954
rect -8458 322718 -8374 322954
rect -8138 322718 -8106 322954
rect -8726 322634 -8106 322718
rect -8726 322398 -8694 322634
rect -8458 322398 -8374 322634
rect -8138 322398 -8106 322634
rect -8726 286954 -8106 322398
rect -8726 286718 -8694 286954
rect -8458 286718 -8374 286954
rect -8138 286718 -8106 286954
rect -8726 286634 -8106 286718
rect -8726 286398 -8694 286634
rect -8458 286398 -8374 286634
rect -8138 286398 -8106 286634
rect -8726 250954 -8106 286398
rect -8726 250718 -8694 250954
rect -8458 250718 -8374 250954
rect -8138 250718 -8106 250954
rect -8726 250634 -8106 250718
rect -8726 250398 -8694 250634
rect -8458 250398 -8374 250634
rect -8138 250398 -8106 250634
rect -8726 214954 -8106 250398
rect -8726 214718 -8694 214954
rect -8458 214718 -8374 214954
rect -8138 214718 -8106 214954
rect -8726 214634 -8106 214718
rect -8726 214398 -8694 214634
rect -8458 214398 -8374 214634
rect -8138 214398 -8106 214634
rect -8726 178954 -8106 214398
rect -8726 178718 -8694 178954
rect -8458 178718 -8374 178954
rect -8138 178718 -8106 178954
rect -8726 178634 -8106 178718
rect -8726 178398 -8694 178634
rect -8458 178398 -8374 178634
rect -8138 178398 -8106 178634
rect -8726 142954 -8106 178398
rect -8726 142718 -8694 142954
rect -8458 142718 -8374 142954
rect -8138 142718 -8106 142954
rect -8726 142634 -8106 142718
rect -8726 142398 -8694 142634
rect -8458 142398 -8374 142634
rect -8138 142398 -8106 142634
rect -8726 106954 -8106 142398
rect -8726 106718 -8694 106954
rect -8458 106718 -8374 106954
rect -8138 106718 -8106 106954
rect -8726 106634 -8106 106718
rect -8726 106398 -8694 106634
rect -8458 106398 -8374 106634
rect -8138 106398 -8106 106634
rect -8726 70954 -8106 106398
rect -8726 70718 -8694 70954
rect -8458 70718 -8374 70954
rect -8138 70718 -8106 70954
rect -8726 70634 -8106 70718
rect -8726 70398 -8694 70634
rect -8458 70398 -8374 70634
rect -8138 70398 -8106 70634
rect -8726 34954 -8106 70398
rect -8726 34718 -8694 34954
rect -8458 34718 -8374 34954
rect -8138 34718 -8106 34954
rect -8726 34634 -8106 34718
rect -8726 34398 -8694 34634
rect -8458 34398 -8374 34634
rect -8138 34398 -8106 34634
rect -8726 -7066 -8106 34398
rect -7766 710598 -7146 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 -7146 710598
rect -7766 710278 -7146 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 -7146 710278
rect -7766 678454 -7146 710042
rect -7766 678218 -7734 678454
rect -7498 678218 -7414 678454
rect -7178 678218 -7146 678454
rect -7766 678134 -7146 678218
rect -7766 677898 -7734 678134
rect -7498 677898 -7414 678134
rect -7178 677898 -7146 678134
rect -7766 642454 -7146 677898
rect -7766 642218 -7734 642454
rect -7498 642218 -7414 642454
rect -7178 642218 -7146 642454
rect -7766 642134 -7146 642218
rect -7766 641898 -7734 642134
rect -7498 641898 -7414 642134
rect -7178 641898 -7146 642134
rect -7766 606454 -7146 641898
rect -7766 606218 -7734 606454
rect -7498 606218 -7414 606454
rect -7178 606218 -7146 606454
rect -7766 606134 -7146 606218
rect -7766 605898 -7734 606134
rect -7498 605898 -7414 606134
rect -7178 605898 -7146 606134
rect -7766 570454 -7146 605898
rect -7766 570218 -7734 570454
rect -7498 570218 -7414 570454
rect -7178 570218 -7146 570454
rect -7766 570134 -7146 570218
rect -7766 569898 -7734 570134
rect -7498 569898 -7414 570134
rect -7178 569898 -7146 570134
rect -7766 534454 -7146 569898
rect -7766 534218 -7734 534454
rect -7498 534218 -7414 534454
rect -7178 534218 -7146 534454
rect -7766 534134 -7146 534218
rect -7766 533898 -7734 534134
rect -7498 533898 -7414 534134
rect -7178 533898 -7146 534134
rect -7766 498454 -7146 533898
rect -7766 498218 -7734 498454
rect -7498 498218 -7414 498454
rect -7178 498218 -7146 498454
rect -7766 498134 -7146 498218
rect -7766 497898 -7734 498134
rect -7498 497898 -7414 498134
rect -7178 497898 -7146 498134
rect -7766 462454 -7146 497898
rect -7766 462218 -7734 462454
rect -7498 462218 -7414 462454
rect -7178 462218 -7146 462454
rect -7766 462134 -7146 462218
rect -7766 461898 -7734 462134
rect -7498 461898 -7414 462134
rect -7178 461898 -7146 462134
rect -7766 426454 -7146 461898
rect -7766 426218 -7734 426454
rect -7498 426218 -7414 426454
rect -7178 426218 -7146 426454
rect -7766 426134 -7146 426218
rect -7766 425898 -7734 426134
rect -7498 425898 -7414 426134
rect -7178 425898 -7146 426134
rect -7766 390454 -7146 425898
rect -7766 390218 -7734 390454
rect -7498 390218 -7414 390454
rect -7178 390218 -7146 390454
rect -7766 390134 -7146 390218
rect -7766 389898 -7734 390134
rect -7498 389898 -7414 390134
rect -7178 389898 -7146 390134
rect -7766 354454 -7146 389898
rect -7766 354218 -7734 354454
rect -7498 354218 -7414 354454
rect -7178 354218 -7146 354454
rect -7766 354134 -7146 354218
rect -7766 353898 -7734 354134
rect -7498 353898 -7414 354134
rect -7178 353898 -7146 354134
rect -7766 318454 -7146 353898
rect -7766 318218 -7734 318454
rect -7498 318218 -7414 318454
rect -7178 318218 -7146 318454
rect -7766 318134 -7146 318218
rect -7766 317898 -7734 318134
rect -7498 317898 -7414 318134
rect -7178 317898 -7146 318134
rect -7766 282454 -7146 317898
rect -7766 282218 -7734 282454
rect -7498 282218 -7414 282454
rect -7178 282218 -7146 282454
rect -7766 282134 -7146 282218
rect -7766 281898 -7734 282134
rect -7498 281898 -7414 282134
rect -7178 281898 -7146 282134
rect -7766 246454 -7146 281898
rect -7766 246218 -7734 246454
rect -7498 246218 -7414 246454
rect -7178 246218 -7146 246454
rect -7766 246134 -7146 246218
rect -7766 245898 -7734 246134
rect -7498 245898 -7414 246134
rect -7178 245898 -7146 246134
rect -7766 210454 -7146 245898
rect -7766 210218 -7734 210454
rect -7498 210218 -7414 210454
rect -7178 210218 -7146 210454
rect -7766 210134 -7146 210218
rect -7766 209898 -7734 210134
rect -7498 209898 -7414 210134
rect -7178 209898 -7146 210134
rect -7766 174454 -7146 209898
rect -7766 174218 -7734 174454
rect -7498 174218 -7414 174454
rect -7178 174218 -7146 174454
rect -7766 174134 -7146 174218
rect -7766 173898 -7734 174134
rect -7498 173898 -7414 174134
rect -7178 173898 -7146 174134
rect -7766 138454 -7146 173898
rect -7766 138218 -7734 138454
rect -7498 138218 -7414 138454
rect -7178 138218 -7146 138454
rect -7766 138134 -7146 138218
rect -7766 137898 -7734 138134
rect -7498 137898 -7414 138134
rect -7178 137898 -7146 138134
rect -7766 102454 -7146 137898
rect -7766 102218 -7734 102454
rect -7498 102218 -7414 102454
rect -7178 102218 -7146 102454
rect -7766 102134 -7146 102218
rect -7766 101898 -7734 102134
rect -7498 101898 -7414 102134
rect -7178 101898 -7146 102134
rect -7766 66454 -7146 101898
rect -7766 66218 -7734 66454
rect -7498 66218 -7414 66454
rect -7178 66218 -7146 66454
rect -7766 66134 -7146 66218
rect -7766 65898 -7734 66134
rect -7498 65898 -7414 66134
rect -7178 65898 -7146 66134
rect -7766 30454 -7146 65898
rect -7766 30218 -7734 30454
rect -7498 30218 -7414 30454
rect -7178 30218 -7146 30454
rect -7766 30134 -7146 30218
rect -7766 29898 -7734 30134
rect -7498 29898 -7414 30134
rect -7178 29898 -7146 30134
rect -7766 -6106 -7146 29898
rect -6806 709638 -6186 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 -6186 709638
rect -6806 709318 -6186 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 -6186 709318
rect -6806 673954 -6186 709082
rect -6806 673718 -6774 673954
rect -6538 673718 -6454 673954
rect -6218 673718 -6186 673954
rect -6806 673634 -6186 673718
rect -6806 673398 -6774 673634
rect -6538 673398 -6454 673634
rect -6218 673398 -6186 673634
rect -6806 637954 -6186 673398
rect -6806 637718 -6774 637954
rect -6538 637718 -6454 637954
rect -6218 637718 -6186 637954
rect -6806 637634 -6186 637718
rect -6806 637398 -6774 637634
rect -6538 637398 -6454 637634
rect -6218 637398 -6186 637634
rect -6806 601954 -6186 637398
rect -6806 601718 -6774 601954
rect -6538 601718 -6454 601954
rect -6218 601718 -6186 601954
rect -6806 601634 -6186 601718
rect -6806 601398 -6774 601634
rect -6538 601398 -6454 601634
rect -6218 601398 -6186 601634
rect -6806 565954 -6186 601398
rect -6806 565718 -6774 565954
rect -6538 565718 -6454 565954
rect -6218 565718 -6186 565954
rect -6806 565634 -6186 565718
rect -6806 565398 -6774 565634
rect -6538 565398 -6454 565634
rect -6218 565398 -6186 565634
rect -6806 529954 -6186 565398
rect -6806 529718 -6774 529954
rect -6538 529718 -6454 529954
rect -6218 529718 -6186 529954
rect -6806 529634 -6186 529718
rect -6806 529398 -6774 529634
rect -6538 529398 -6454 529634
rect -6218 529398 -6186 529634
rect -6806 493954 -6186 529398
rect -6806 493718 -6774 493954
rect -6538 493718 -6454 493954
rect -6218 493718 -6186 493954
rect -6806 493634 -6186 493718
rect -6806 493398 -6774 493634
rect -6538 493398 -6454 493634
rect -6218 493398 -6186 493634
rect -6806 457954 -6186 493398
rect -6806 457718 -6774 457954
rect -6538 457718 -6454 457954
rect -6218 457718 -6186 457954
rect -6806 457634 -6186 457718
rect -6806 457398 -6774 457634
rect -6538 457398 -6454 457634
rect -6218 457398 -6186 457634
rect -6806 421954 -6186 457398
rect -6806 421718 -6774 421954
rect -6538 421718 -6454 421954
rect -6218 421718 -6186 421954
rect -6806 421634 -6186 421718
rect -6806 421398 -6774 421634
rect -6538 421398 -6454 421634
rect -6218 421398 -6186 421634
rect -6806 385954 -6186 421398
rect -6806 385718 -6774 385954
rect -6538 385718 -6454 385954
rect -6218 385718 -6186 385954
rect -6806 385634 -6186 385718
rect -6806 385398 -6774 385634
rect -6538 385398 -6454 385634
rect -6218 385398 -6186 385634
rect -6806 349954 -6186 385398
rect -6806 349718 -6774 349954
rect -6538 349718 -6454 349954
rect -6218 349718 -6186 349954
rect -6806 349634 -6186 349718
rect -6806 349398 -6774 349634
rect -6538 349398 -6454 349634
rect -6218 349398 -6186 349634
rect -6806 313954 -6186 349398
rect -6806 313718 -6774 313954
rect -6538 313718 -6454 313954
rect -6218 313718 -6186 313954
rect -6806 313634 -6186 313718
rect -6806 313398 -6774 313634
rect -6538 313398 -6454 313634
rect -6218 313398 -6186 313634
rect -6806 277954 -6186 313398
rect -6806 277718 -6774 277954
rect -6538 277718 -6454 277954
rect -6218 277718 -6186 277954
rect -6806 277634 -6186 277718
rect -6806 277398 -6774 277634
rect -6538 277398 -6454 277634
rect -6218 277398 -6186 277634
rect -6806 241954 -6186 277398
rect -6806 241718 -6774 241954
rect -6538 241718 -6454 241954
rect -6218 241718 -6186 241954
rect -6806 241634 -6186 241718
rect -6806 241398 -6774 241634
rect -6538 241398 -6454 241634
rect -6218 241398 -6186 241634
rect -6806 205954 -6186 241398
rect -6806 205718 -6774 205954
rect -6538 205718 -6454 205954
rect -6218 205718 -6186 205954
rect -6806 205634 -6186 205718
rect -6806 205398 -6774 205634
rect -6538 205398 -6454 205634
rect -6218 205398 -6186 205634
rect -6806 169954 -6186 205398
rect -6806 169718 -6774 169954
rect -6538 169718 -6454 169954
rect -6218 169718 -6186 169954
rect -6806 169634 -6186 169718
rect -6806 169398 -6774 169634
rect -6538 169398 -6454 169634
rect -6218 169398 -6186 169634
rect -6806 133954 -6186 169398
rect -6806 133718 -6774 133954
rect -6538 133718 -6454 133954
rect -6218 133718 -6186 133954
rect -6806 133634 -6186 133718
rect -6806 133398 -6774 133634
rect -6538 133398 -6454 133634
rect -6218 133398 -6186 133634
rect -6806 97954 -6186 133398
rect -6806 97718 -6774 97954
rect -6538 97718 -6454 97954
rect -6218 97718 -6186 97954
rect -6806 97634 -6186 97718
rect -6806 97398 -6774 97634
rect -6538 97398 -6454 97634
rect -6218 97398 -6186 97634
rect -6806 61954 -6186 97398
rect -6806 61718 -6774 61954
rect -6538 61718 -6454 61954
rect -6218 61718 -6186 61954
rect -6806 61634 -6186 61718
rect -6806 61398 -6774 61634
rect -6538 61398 -6454 61634
rect -6218 61398 -6186 61634
rect -6806 25954 -6186 61398
rect -6806 25718 -6774 25954
rect -6538 25718 -6454 25954
rect -6218 25718 -6186 25954
rect -6806 25634 -6186 25718
rect -6806 25398 -6774 25634
rect -6538 25398 -6454 25634
rect -6218 25398 -6186 25634
rect -6806 -5146 -6186 25398
rect -5846 708678 -5226 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 -5226 708678
rect -5846 708358 -5226 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 -5226 708358
rect -5846 669454 -5226 708122
rect -5846 669218 -5814 669454
rect -5578 669218 -5494 669454
rect -5258 669218 -5226 669454
rect -5846 669134 -5226 669218
rect -5846 668898 -5814 669134
rect -5578 668898 -5494 669134
rect -5258 668898 -5226 669134
rect -5846 633454 -5226 668898
rect -5846 633218 -5814 633454
rect -5578 633218 -5494 633454
rect -5258 633218 -5226 633454
rect -5846 633134 -5226 633218
rect -5846 632898 -5814 633134
rect -5578 632898 -5494 633134
rect -5258 632898 -5226 633134
rect -5846 597454 -5226 632898
rect -5846 597218 -5814 597454
rect -5578 597218 -5494 597454
rect -5258 597218 -5226 597454
rect -5846 597134 -5226 597218
rect -5846 596898 -5814 597134
rect -5578 596898 -5494 597134
rect -5258 596898 -5226 597134
rect -5846 561454 -5226 596898
rect -5846 561218 -5814 561454
rect -5578 561218 -5494 561454
rect -5258 561218 -5226 561454
rect -5846 561134 -5226 561218
rect -5846 560898 -5814 561134
rect -5578 560898 -5494 561134
rect -5258 560898 -5226 561134
rect -5846 525454 -5226 560898
rect -5846 525218 -5814 525454
rect -5578 525218 -5494 525454
rect -5258 525218 -5226 525454
rect -5846 525134 -5226 525218
rect -5846 524898 -5814 525134
rect -5578 524898 -5494 525134
rect -5258 524898 -5226 525134
rect -5846 489454 -5226 524898
rect -5846 489218 -5814 489454
rect -5578 489218 -5494 489454
rect -5258 489218 -5226 489454
rect -5846 489134 -5226 489218
rect -5846 488898 -5814 489134
rect -5578 488898 -5494 489134
rect -5258 488898 -5226 489134
rect -5846 453454 -5226 488898
rect -5846 453218 -5814 453454
rect -5578 453218 -5494 453454
rect -5258 453218 -5226 453454
rect -5846 453134 -5226 453218
rect -5846 452898 -5814 453134
rect -5578 452898 -5494 453134
rect -5258 452898 -5226 453134
rect -5846 417454 -5226 452898
rect -5846 417218 -5814 417454
rect -5578 417218 -5494 417454
rect -5258 417218 -5226 417454
rect -5846 417134 -5226 417218
rect -5846 416898 -5814 417134
rect -5578 416898 -5494 417134
rect -5258 416898 -5226 417134
rect -5846 381454 -5226 416898
rect -5846 381218 -5814 381454
rect -5578 381218 -5494 381454
rect -5258 381218 -5226 381454
rect -5846 381134 -5226 381218
rect -5846 380898 -5814 381134
rect -5578 380898 -5494 381134
rect -5258 380898 -5226 381134
rect -5846 345454 -5226 380898
rect -5846 345218 -5814 345454
rect -5578 345218 -5494 345454
rect -5258 345218 -5226 345454
rect -5846 345134 -5226 345218
rect -5846 344898 -5814 345134
rect -5578 344898 -5494 345134
rect -5258 344898 -5226 345134
rect -5846 309454 -5226 344898
rect -5846 309218 -5814 309454
rect -5578 309218 -5494 309454
rect -5258 309218 -5226 309454
rect -5846 309134 -5226 309218
rect -5846 308898 -5814 309134
rect -5578 308898 -5494 309134
rect -5258 308898 -5226 309134
rect -5846 273454 -5226 308898
rect -5846 273218 -5814 273454
rect -5578 273218 -5494 273454
rect -5258 273218 -5226 273454
rect -5846 273134 -5226 273218
rect -5846 272898 -5814 273134
rect -5578 272898 -5494 273134
rect -5258 272898 -5226 273134
rect -5846 237454 -5226 272898
rect -5846 237218 -5814 237454
rect -5578 237218 -5494 237454
rect -5258 237218 -5226 237454
rect -5846 237134 -5226 237218
rect -5846 236898 -5814 237134
rect -5578 236898 -5494 237134
rect -5258 236898 -5226 237134
rect -5846 201454 -5226 236898
rect -5846 201218 -5814 201454
rect -5578 201218 -5494 201454
rect -5258 201218 -5226 201454
rect -5846 201134 -5226 201218
rect -5846 200898 -5814 201134
rect -5578 200898 -5494 201134
rect -5258 200898 -5226 201134
rect -5846 165454 -5226 200898
rect -5846 165218 -5814 165454
rect -5578 165218 -5494 165454
rect -5258 165218 -5226 165454
rect -5846 165134 -5226 165218
rect -5846 164898 -5814 165134
rect -5578 164898 -5494 165134
rect -5258 164898 -5226 165134
rect -5846 129454 -5226 164898
rect -5846 129218 -5814 129454
rect -5578 129218 -5494 129454
rect -5258 129218 -5226 129454
rect -5846 129134 -5226 129218
rect -5846 128898 -5814 129134
rect -5578 128898 -5494 129134
rect -5258 128898 -5226 129134
rect -5846 93454 -5226 128898
rect -5846 93218 -5814 93454
rect -5578 93218 -5494 93454
rect -5258 93218 -5226 93454
rect -5846 93134 -5226 93218
rect -5846 92898 -5814 93134
rect -5578 92898 -5494 93134
rect -5258 92898 -5226 93134
rect -5846 57454 -5226 92898
rect -5846 57218 -5814 57454
rect -5578 57218 -5494 57454
rect -5258 57218 -5226 57454
rect -5846 57134 -5226 57218
rect -5846 56898 -5814 57134
rect -5578 56898 -5494 57134
rect -5258 56898 -5226 57134
rect -5846 21454 -5226 56898
rect -5846 21218 -5814 21454
rect -5578 21218 -5494 21454
rect -5258 21218 -5226 21454
rect -5846 21134 -5226 21218
rect -5846 20898 -5814 21134
rect -5578 20898 -5494 21134
rect -5258 20898 -5226 21134
rect -5846 -4186 -5226 20898
rect -4886 707718 -4266 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 -4266 707718
rect -4886 707398 -4266 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 -4266 707398
rect -4886 700954 -4266 707162
rect -4886 700718 -4854 700954
rect -4618 700718 -4534 700954
rect -4298 700718 -4266 700954
rect -4886 700634 -4266 700718
rect -4886 700398 -4854 700634
rect -4618 700398 -4534 700634
rect -4298 700398 -4266 700634
rect -4886 664954 -4266 700398
rect -4886 664718 -4854 664954
rect -4618 664718 -4534 664954
rect -4298 664718 -4266 664954
rect -4886 664634 -4266 664718
rect -4886 664398 -4854 664634
rect -4618 664398 -4534 664634
rect -4298 664398 -4266 664634
rect -4886 628954 -4266 664398
rect -4886 628718 -4854 628954
rect -4618 628718 -4534 628954
rect -4298 628718 -4266 628954
rect -4886 628634 -4266 628718
rect -4886 628398 -4854 628634
rect -4618 628398 -4534 628634
rect -4298 628398 -4266 628634
rect -4886 592954 -4266 628398
rect -4886 592718 -4854 592954
rect -4618 592718 -4534 592954
rect -4298 592718 -4266 592954
rect -4886 592634 -4266 592718
rect -4886 592398 -4854 592634
rect -4618 592398 -4534 592634
rect -4298 592398 -4266 592634
rect -4886 556954 -4266 592398
rect -4886 556718 -4854 556954
rect -4618 556718 -4534 556954
rect -4298 556718 -4266 556954
rect -4886 556634 -4266 556718
rect -4886 556398 -4854 556634
rect -4618 556398 -4534 556634
rect -4298 556398 -4266 556634
rect -4886 520954 -4266 556398
rect -4886 520718 -4854 520954
rect -4618 520718 -4534 520954
rect -4298 520718 -4266 520954
rect -4886 520634 -4266 520718
rect -4886 520398 -4854 520634
rect -4618 520398 -4534 520634
rect -4298 520398 -4266 520634
rect -4886 484954 -4266 520398
rect -4886 484718 -4854 484954
rect -4618 484718 -4534 484954
rect -4298 484718 -4266 484954
rect -4886 484634 -4266 484718
rect -4886 484398 -4854 484634
rect -4618 484398 -4534 484634
rect -4298 484398 -4266 484634
rect -4886 448954 -4266 484398
rect -4886 448718 -4854 448954
rect -4618 448718 -4534 448954
rect -4298 448718 -4266 448954
rect -4886 448634 -4266 448718
rect -4886 448398 -4854 448634
rect -4618 448398 -4534 448634
rect -4298 448398 -4266 448634
rect -4886 412954 -4266 448398
rect -4886 412718 -4854 412954
rect -4618 412718 -4534 412954
rect -4298 412718 -4266 412954
rect -4886 412634 -4266 412718
rect -4886 412398 -4854 412634
rect -4618 412398 -4534 412634
rect -4298 412398 -4266 412634
rect -4886 376954 -4266 412398
rect -4886 376718 -4854 376954
rect -4618 376718 -4534 376954
rect -4298 376718 -4266 376954
rect -4886 376634 -4266 376718
rect -4886 376398 -4854 376634
rect -4618 376398 -4534 376634
rect -4298 376398 -4266 376634
rect -4886 340954 -4266 376398
rect -4886 340718 -4854 340954
rect -4618 340718 -4534 340954
rect -4298 340718 -4266 340954
rect -4886 340634 -4266 340718
rect -4886 340398 -4854 340634
rect -4618 340398 -4534 340634
rect -4298 340398 -4266 340634
rect -4886 304954 -4266 340398
rect -4886 304718 -4854 304954
rect -4618 304718 -4534 304954
rect -4298 304718 -4266 304954
rect -4886 304634 -4266 304718
rect -4886 304398 -4854 304634
rect -4618 304398 -4534 304634
rect -4298 304398 -4266 304634
rect -4886 268954 -4266 304398
rect -4886 268718 -4854 268954
rect -4618 268718 -4534 268954
rect -4298 268718 -4266 268954
rect -4886 268634 -4266 268718
rect -4886 268398 -4854 268634
rect -4618 268398 -4534 268634
rect -4298 268398 -4266 268634
rect -4886 232954 -4266 268398
rect -4886 232718 -4854 232954
rect -4618 232718 -4534 232954
rect -4298 232718 -4266 232954
rect -4886 232634 -4266 232718
rect -4886 232398 -4854 232634
rect -4618 232398 -4534 232634
rect -4298 232398 -4266 232634
rect -4886 196954 -4266 232398
rect -4886 196718 -4854 196954
rect -4618 196718 -4534 196954
rect -4298 196718 -4266 196954
rect -4886 196634 -4266 196718
rect -4886 196398 -4854 196634
rect -4618 196398 -4534 196634
rect -4298 196398 -4266 196634
rect -4886 160954 -4266 196398
rect -4886 160718 -4854 160954
rect -4618 160718 -4534 160954
rect -4298 160718 -4266 160954
rect -4886 160634 -4266 160718
rect -4886 160398 -4854 160634
rect -4618 160398 -4534 160634
rect -4298 160398 -4266 160634
rect -4886 124954 -4266 160398
rect -4886 124718 -4854 124954
rect -4618 124718 -4534 124954
rect -4298 124718 -4266 124954
rect -4886 124634 -4266 124718
rect -4886 124398 -4854 124634
rect -4618 124398 -4534 124634
rect -4298 124398 -4266 124634
rect -4886 88954 -4266 124398
rect -4886 88718 -4854 88954
rect -4618 88718 -4534 88954
rect -4298 88718 -4266 88954
rect -4886 88634 -4266 88718
rect -4886 88398 -4854 88634
rect -4618 88398 -4534 88634
rect -4298 88398 -4266 88634
rect -4886 52954 -4266 88398
rect -4886 52718 -4854 52954
rect -4618 52718 -4534 52954
rect -4298 52718 -4266 52954
rect -4886 52634 -4266 52718
rect -4886 52398 -4854 52634
rect -4618 52398 -4534 52634
rect -4298 52398 -4266 52634
rect -4886 16954 -4266 52398
rect -4886 16718 -4854 16954
rect -4618 16718 -4534 16954
rect -4298 16718 -4266 16954
rect -4886 16634 -4266 16718
rect -4886 16398 -4854 16634
rect -4618 16398 -4534 16634
rect -4298 16398 -4266 16634
rect -4886 -3226 -4266 16398
rect -3926 706758 -3306 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 -3306 706758
rect -3926 706438 -3306 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 -3306 706438
rect -3926 696454 -3306 706202
rect -3926 696218 -3894 696454
rect -3658 696218 -3574 696454
rect -3338 696218 -3306 696454
rect -3926 696134 -3306 696218
rect -3926 695898 -3894 696134
rect -3658 695898 -3574 696134
rect -3338 695898 -3306 696134
rect -3926 660454 -3306 695898
rect -3926 660218 -3894 660454
rect -3658 660218 -3574 660454
rect -3338 660218 -3306 660454
rect -3926 660134 -3306 660218
rect -3926 659898 -3894 660134
rect -3658 659898 -3574 660134
rect -3338 659898 -3306 660134
rect -3926 624454 -3306 659898
rect -3926 624218 -3894 624454
rect -3658 624218 -3574 624454
rect -3338 624218 -3306 624454
rect -3926 624134 -3306 624218
rect -3926 623898 -3894 624134
rect -3658 623898 -3574 624134
rect -3338 623898 -3306 624134
rect -3926 588454 -3306 623898
rect -3926 588218 -3894 588454
rect -3658 588218 -3574 588454
rect -3338 588218 -3306 588454
rect -3926 588134 -3306 588218
rect -3926 587898 -3894 588134
rect -3658 587898 -3574 588134
rect -3338 587898 -3306 588134
rect -3926 552454 -3306 587898
rect -3926 552218 -3894 552454
rect -3658 552218 -3574 552454
rect -3338 552218 -3306 552454
rect -3926 552134 -3306 552218
rect -3926 551898 -3894 552134
rect -3658 551898 -3574 552134
rect -3338 551898 -3306 552134
rect -3926 516454 -3306 551898
rect -3926 516218 -3894 516454
rect -3658 516218 -3574 516454
rect -3338 516218 -3306 516454
rect -3926 516134 -3306 516218
rect -3926 515898 -3894 516134
rect -3658 515898 -3574 516134
rect -3338 515898 -3306 516134
rect -3926 480454 -3306 515898
rect -3926 480218 -3894 480454
rect -3658 480218 -3574 480454
rect -3338 480218 -3306 480454
rect -3926 480134 -3306 480218
rect -3926 479898 -3894 480134
rect -3658 479898 -3574 480134
rect -3338 479898 -3306 480134
rect -3926 444454 -3306 479898
rect -3926 444218 -3894 444454
rect -3658 444218 -3574 444454
rect -3338 444218 -3306 444454
rect -3926 444134 -3306 444218
rect -3926 443898 -3894 444134
rect -3658 443898 -3574 444134
rect -3338 443898 -3306 444134
rect -3926 408454 -3306 443898
rect -3926 408218 -3894 408454
rect -3658 408218 -3574 408454
rect -3338 408218 -3306 408454
rect -3926 408134 -3306 408218
rect -3926 407898 -3894 408134
rect -3658 407898 -3574 408134
rect -3338 407898 -3306 408134
rect -3926 372454 -3306 407898
rect -3926 372218 -3894 372454
rect -3658 372218 -3574 372454
rect -3338 372218 -3306 372454
rect -3926 372134 -3306 372218
rect -3926 371898 -3894 372134
rect -3658 371898 -3574 372134
rect -3338 371898 -3306 372134
rect -3926 336454 -3306 371898
rect -3926 336218 -3894 336454
rect -3658 336218 -3574 336454
rect -3338 336218 -3306 336454
rect -3926 336134 -3306 336218
rect -3926 335898 -3894 336134
rect -3658 335898 -3574 336134
rect -3338 335898 -3306 336134
rect -3926 300454 -3306 335898
rect -3926 300218 -3894 300454
rect -3658 300218 -3574 300454
rect -3338 300218 -3306 300454
rect -3926 300134 -3306 300218
rect -3926 299898 -3894 300134
rect -3658 299898 -3574 300134
rect -3338 299898 -3306 300134
rect -3926 264454 -3306 299898
rect -3926 264218 -3894 264454
rect -3658 264218 -3574 264454
rect -3338 264218 -3306 264454
rect -3926 264134 -3306 264218
rect -3926 263898 -3894 264134
rect -3658 263898 -3574 264134
rect -3338 263898 -3306 264134
rect -3926 228454 -3306 263898
rect -3926 228218 -3894 228454
rect -3658 228218 -3574 228454
rect -3338 228218 -3306 228454
rect -3926 228134 -3306 228218
rect -3926 227898 -3894 228134
rect -3658 227898 -3574 228134
rect -3338 227898 -3306 228134
rect -3926 192454 -3306 227898
rect -3926 192218 -3894 192454
rect -3658 192218 -3574 192454
rect -3338 192218 -3306 192454
rect -3926 192134 -3306 192218
rect -3926 191898 -3894 192134
rect -3658 191898 -3574 192134
rect -3338 191898 -3306 192134
rect -3926 156454 -3306 191898
rect -3926 156218 -3894 156454
rect -3658 156218 -3574 156454
rect -3338 156218 -3306 156454
rect -3926 156134 -3306 156218
rect -3926 155898 -3894 156134
rect -3658 155898 -3574 156134
rect -3338 155898 -3306 156134
rect -3926 120454 -3306 155898
rect -3926 120218 -3894 120454
rect -3658 120218 -3574 120454
rect -3338 120218 -3306 120454
rect -3926 120134 -3306 120218
rect -3926 119898 -3894 120134
rect -3658 119898 -3574 120134
rect -3338 119898 -3306 120134
rect -3926 84454 -3306 119898
rect -3926 84218 -3894 84454
rect -3658 84218 -3574 84454
rect -3338 84218 -3306 84454
rect -3926 84134 -3306 84218
rect -3926 83898 -3894 84134
rect -3658 83898 -3574 84134
rect -3338 83898 -3306 84134
rect -3926 48454 -3306 83898
rect -3926 48218 -3894 48454
rect -3658 48218 -3574 48454
rect -3338 48218 -3306 48454
rect -3926 48134 -3306 48218
rect -3926 47898 -3894 48134
rect -3658 47898 -3574 48134
rect -3338 47898 -3306 48134
rect -3926 12454 -3306 47898
rect -3926 12218 -3894 12454
rect -3658 12218 -3574 12454
rect -3338 12218 -3306 12454
rect -3926 12134 -3306 12218
rect -3926 11898 -3894 12134
rect -3658 11898 -3574 12134
rect -3338 11898 -3306 12134
rect -3926 -2266 -3306 11898
rect -2966 705798 -2346 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 -2346 705798
rect -2966 705478 -2346 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 -2346 705478
rect -2966 691954 -2346 705242
rect -2966 691718 -2934 691954
rect -2698 691718 -2614 691954
rect -2378 691718 -2346 691954
rect -2966 691634 -2346 691718
rect -2966 691398 -2934 691634
rect -2698 691398 -2614 691634
rect -2378 691398 -2346 691634
rect -2966 655954 -2346 691398
rect -2966 655718 -2934 655954
rect -2698 655718 -2614 655954
rect -2378 655718 -2346 655954
rect -2966 655634 -2346 655718
rect -2966 655398 -2934 655634
rect -2698 655398 -2614 655634
rect -2378 655398 -2346 655634
rect -2966 619954 -2346 655398
rect -2966 619718 -2934 619954
rect -2698 619718 -2614 619954
rect -2378 619718 -2346 619954
rect -2966 619634 -2346 619718
rect -2966 619398 -2934 619634
rect -2698 619398 -2614 619634
rect -2378 619398 -2346 619634
rect -2966 583954 -2346 619398
rect -2966 583718 -2934 583954
rect -2698 583718 -2614 583954
rect -2378 583718 -2346 583954
rect -2966 583634 -2346 583718
rect -2966 583398 -2934 583634
rect -2698 583398 -2614 583634
rect -2378 583398 -2346 583634
rect -2966 547954 -2346 583398
rect -2966 547718 -2934 547954
rect -2698 547718 -2614 547954
rect -2378 547718 -2346 547954
rect -2966 547634 -2346 547718
rect -2966 547398 -2934 547634
rect -2698 547398 -2614 547634
rect -2378 547398 -2346 547634
rect -2966 511954 -2346 547398
rect -2966 511718 -2934 511954
rect -2698 511718 -2614 511954
rect -2378 511718 -2346 511954
rect -2966 511634 -2346 511718
rect -2966 511398 -2934 511634
rect -2698 511398 -2614 511634
rect -2378 511398 -2346 511634
rect -2966 475954 -2346 511398
rect -2966 475718 -2934 475954
rect -2698 475718 -2614 475954
rect -2378 475718 -2346 475954
rect -2966 475634 -2346 475718
rect -2966 475398 -2934 475634
rect -2698 475398 -2614 475634
rect -2378 475398 -2346 475634
rect -2966 439954 -2346 475398
rect -2966 439718 -2934 439954
rect -2698 439718 -2614 439954
rect -2378 439718 -2346 439954
rect -2966 439634 -2346 439718
rect -2966 439398 -2934 439634
rect -2698 439398 -2614 439634
rect -2378 439398 -2346 439634
rect -2966 403954 -2346 439398
rect -2966 403718 -2934 403954
rect -2698 403718 -2614 403954
rect -2378 403718 -2346 403954
rect -2966 403634 -2346 403718
rect -2966 403398 -2934 403634
rect -2698 403398 -2614 403634
rect -2378 403398 -2346 403634
rect -2966 367954 -2346 403398
rect -2966 367718 -2934 367954
rect -2698 367718 -2614 367954
rect -2378 367718 -2346 367954
rect -2966 367634 -2346 367718
rect -2966 367398 -2934 367634
rect -2698 367398 -2614 367634
rect -2378 367398 -2346 367634
rect -2966 331954 -2346 367398
rect -2966 331718 -2934 331954
rect -2698 331718 -2614 331954
rect -2378 331718 -2346 331954
rect -2966 331634 -2346 331718
rect -2966 331398 -2934 331634
rect -2698 331398 -2614 331634
rect -2378 331398 -2346 331634
rect -2966 295954 -2346 331398
rect -2966 295718 -2934 295954
rect -2698 295718 -2614 295954
rect -2378 295718 -2346 295954
rect -2966 295634 -2346 295718
rect -2966 295398 -2934 295634
rect -2698 295398 -2614 295634
rect -2378 295398 -2346 295634
rect -2966 259954 -2346 295398
rect -2966 259718 -2934 259954
rect -2698 259718 -2614 259954
rect -2378 259718 -2346 259954
rect -2966 259634 -2346 259718
rect -2966 259398 -2934 259634
rect -2698 259398 -2614 259634
rect -2378 259398 -2346 259634
rect -2966 223954 -2346 259398
rect -2966 223718 -2934 223954
rect -2698 223718 -2614 223954
rect -2378 223718 -2346 223954
rect -2966 223634 -2346 223718
rect -2966 223398 -2934 223634
rect -2698 223398 -2614 223634
rect -2378 223398 -2346 223634
rect -2966 187954 -2346 223398
rect -2966 187718 -2934 187954
rect -2698 187718 -2614 187954
rect -2378 187718 -2346 187954
rect -2966 187634 -2346 187718
rect -2966 187398 -2934 187634
rect -2698 187398 -2614 187634
rect -2378 187398 -2346 187634
rect -2966 151954 -2346 187398
rect -2966 151718 -2934 151954
rect -2698 151718 -2614 151954
rect -2378 151718 -2346 151954
rect -2966 151634 -2346 151718
rect -2966 151398 -2934 151634
rect -2698 151398 -2614 151634
rect -2378 151398 -2346 151634
rect -2966 115954 -2346 151398
rect -2966 115718 -2934 115954
rect -2698 115718 -2614 115954
rect -2378 115718 -2346 115954
rect -2966 115634 -2346 115718
rect -2966 115398 -2934 115634
rect -2698 115398 -2614 115634
rect -2378 115398 -2346 115634
rect -2966 79954 -2346 115398
rect -2966 79718 -2934 79954
rect -2698 79718 -2614 79954
rect -2378 79718 -2346 79954
rect -2966 79634 -2346 79718
rect -2966 79398 -2934 79634
rect -2698 79398 -2614 79634
rect -2378 79398 -2346 79634
rect -2966 43954 -2346 79398
rect -2966 43718 -2934 43954
rect -2698 43718 -2614 43954
rect -2378 43718 -2346 43954
rect -2966 43634 -2346 43718
rect -2966 43398 -2934 43634
rect -2698 43398 -2614 43634
rect -2378 43398 -2346 43634
rect -2966 7954 -2346 43398
rect -2966 7718 -2934 7954
rect -2698 7718 -2614 7954
rect -2378 7718 -2346 7954
rect -2966 7634 -2346 7718
rect -2966 7398 -2934 7634
rect -2698 7398 -2614 7634
rect -2378 7398 -2346 7634
rect -2966 -1306 -2346 7398
rect -2006 704838 -1386 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 -1386 704838
rect -2006 704518 -1386 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 -1386 704518
rect -2006 687454 -1386 704282
rect -2006 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 -1386 687454
rect -2006 687134 -1386 687218
rect -2006 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 -1386 687134
rect -2006 651454 -1386 686898
rect -2006 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 -1386 651454
rect -2006 651134 -1386 651218
rect -2006 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 -1386 651134
rect -2006 615454 -1386 650898
rect -2006 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 -1386 615454
rect -2006 615134 -1386 615218
rect -2006 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 -1386 615134
rect -2006 579454 -1386 614898
rect -2006 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 -1386 579454
rect -2006 579134 -1386 579218
rect -2006 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 -1386 579134
rect -2006 543454 -1386 578898
rect -2006 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 -1386 543454
rect -2006 543134 -1386 543218
rect -2006 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 -1386 543134
rect -2006 507454 -1386 542898
rect -2006 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 -1386 507454
rect -2006 507134 -1386 507218
rect -2006 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 -1386 507134
rect -2006 471454 -1386 506898
rect -2006 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 -1386 471454
rect -2006 471134 -1386 471218
rect -2006 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 -1386 471134
rect -2006 435454 -1386 470898
rect -2006 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 -1386 435454
rect -2006 435134 -1386 435218
rect -2006 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 -1386 435134
rect -2006 399454 -1386 434898
rect -2006 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 -1386 399454
rect -2006 399134 -1386 399218
rect -2006 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 -1386 399134
rect -2006 363454 -1386 398898
rect -2006 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 -1386 363454
rect -2006 363134 -1386 363218
rect -2006 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 -1386 363134
rect -2006 327454 -1386 362898
rect -2006 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 -1386 327454
rect -2006 327134 -1386 327218
rect -2006 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 -1386 327134
rect -2006 291454 -1386 326898
rect -2006 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 -1386 291454
rect -2006 291134 -1386 291218
rect -2006 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 -1386 291134
rect -2006 255454 -1386 290898
rect -2006 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 -1386 255454
rect -2006 255134 -1386 255218
rect -2006 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 -1386 255134
rect -2006 219454 -1386 254898
rect -2006 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 -1386 219454
rect -2006 219134 -1386 219218
rect -2006 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 -1386 219134
rect -2006 183454 -1386 218898
rect -2006 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 -1386 183454
rect -2006 183134 -1386 183218
rect -2006 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 -1386 183134
rect -2006 147454 -1386 182898
rect -2006 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 -1386 147454
rect -2006 147134 -1386 147218
rect -2006 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 -1386 147134
rect -2006 111454 -1386 146898
rect -2006 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 -1386 111454
rect -2006 111134 -1386 111218
rect -2006 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 -1386 111134
rect -2006 75454 -1386 110898
rect -2006 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 -1386 75454
rect -2006 75134 -1386 75218
rect -2006 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 -1386 75134
rect -2006 39454 -1386 74898
rect -2006 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 -1386 39454
rect -2006 39134 -1386 39218
rect -2006 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 -1386 39134
rect -2006 3454 -1386 38898
rect -2006 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 -1386 3454
rect -2006 3134 -1386 3218
rect -2006 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 -1386 3134
rect -2006 -346 -1386 2898
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 -1386 -346
rect -2006 -666 -1386 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 -1386 -666
rect -2006 -934 -1386 -902
rect 1794 704838 2414 711590
rect 1794 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 2414 704838
rect 1794 704518 2414 704602
rect 1794 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 2414 704518
rect 1794 687454 2414 704282
rect 1794 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 2414 687454
rect 1794 687134 2414 687218
rect 1794 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 2414 687134
rect 1794 651454 2414 686898
rect 1794 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 2414 651454
rect 1794 651134 2414 651218
rect 1794 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 2414 651134
rect 1794 615454 2414 650898
rect 1794 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 2414 615454
rect 1794 615134 2414 615218
rect 1794 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 2414 615134
rect 1794 579454 2414 614898
rect 1794 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 2414 579454
rect 1794 579134 2414 579218
rect 1794 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 2414 579134
rect 1794 543454 2414 578898
rect 1794 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 2414 543454
rect 1794 543134 2414 543218
rect 1794 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 2414 543134
rect 1794 507454 2414 542898
rect 1794 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 2414 507454
rect 1794 507134 2414 507218
rect 1794 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 2414 507134
rect 1794 471454 2414 506898
rect 1794 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 2414 471454
rect 1794 471134 2414 471218
rect 1794 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 2414 471134
rect 1794 435454 2414 470898
rect 1794 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 2414 435454
rect 1794 435134 2414 435218
rect 1794 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 2414 435134
rect 1794 399454 2414 434898
rect 1794 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 2414 399454
rect 1794 399134 2414 399218
rect 1794 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 2414 399134
rect 1794 363454 2414 398898
rect 1794 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 2414 363454
rect 1794 363134 2414 363218
rect 1794 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 2414 363134
rect 1794 327454 2414 362898
rect 1794 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 2414 327454
rect 1794 327134 2414 327218
rect 1794 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 2414 327134
rect 1794 291454 2414 326898
rect 1794 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 2414 291454
rect 1794 291134 2414 291218
rect 1794 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 2414 291134
rect 1794 255454 2414 290898
rect 1794 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 2414 255454
rect 1794 255134 2414 255218
rect 1794 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 2414 255134
rect 1794 219454 2414 254898
rect 1794 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 2414 219454
rect 1794 219134 2414 219218
rect 1794 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 2414 219134
rect 1794 183454 2414 218898
rect 1794 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 2414 183454
rect 1794 183134 2414 183218
rect 1794 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 2414 183134
rect 1794 147454 2414 182898
rect 1794 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 2414 147454
rect 1794 147134 2414 147218
rect 1794 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 2414 147134
rect 1794 111454 2414 146898
rect 1794 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 2414 111454
rect 1794 111134 2414 111218
rect 1794 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 2414 111134
rect 1794 75454 2414 110898
rect 1794 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 2414 75454
rect 1794 75134 2414 75218
rect 1794 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 2414 75134
rect 1794 39454 2414 74898
rect 1794 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 2414 39454
rect 1794 39134 2414 39218
rect 1794 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 2414 39134
rect 1794 3454 2414 38898
rect 1794 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 2414 3454
rect 1794 3134 2414 3218
rect 1794 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 2414 3134
rect 1794 -346 2414 2898
rect 1794 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 2414 -346
rect 1794 -666 2414 -582
rect 1794 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 2414 -666
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 -2346 -1306
rect -2966 -1626 -2346 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 -2346 -1626
rect -2966 -1894 -2346 -1862
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 -3306 -2266
rect -3926 -2586 -3306 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 -3306 -2586
rect -3926 -2854 -3306 -2822
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 -4266 -3226
rect -4886 -3546 -4266 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 -4266 -3546
rect -4886 -3814 -4266 -3782
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 -5226 -4186
rect -5846 -4506 -5226 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 -5226 -4506
rect -5846 -4774 -5226 -4742
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 -6186 -5146
rect -6806 -5466 -6186 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 -6186 -5466
rect -6806 -5734 -6186 -5702
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 -7146 -6106
rect -7766 -6426 -7146 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 -7146 -6426
rect -7766 -6694 -7146 -6662
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 -8106 -7066
rect -8726 -7386 -8106 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 -8106 -7386
rect -8726 -7654 -8106 -7622
rect 1794 -7654 2414 -902
rect 6294 705798 6914 711590
rect 6294 705562 6326 705798
rect 6562 705562 6646 705798
rect 6882 705562 6914 705798
rect 6294 705478 6914 705562
rect 6294 705242 6326 705478
rect 6562 705242 6646 705478
rect 6882 705242 6914 705478
rect 6294 691954 6914 705242
rect 6294 691718 6326 691954
rect 6562 691718 6646 691954
rect 6882 691718 6914 691954
rect 6294 691634 6914 691718
rect 6294 691398 6326 691634
rect 6562 691398 6646 691634
rect 6882 691398 6914 691634
rect 6294 655954 6914 691398
rect 6294 655718 6326 655954
rect 6562 655718 6646 655954
rect 6882 655718 6914 655954
rect 6294 655634 6914 655718
rect 6294 655398 6326 655634
rect 6562 655398 6646 655634
rect 6882 655398 6914 655634
rect 6294 619954 6914 655398
rect 6294 619718 6326 619954
rect 6562 619718 6646 619954
rect 6882 619718 6914 619954
rect 6294 619634 6914 619718
rect 6294 619398 6326 619634
rect 6562 619398 6646 619634
rect 6882 619398 6914 619634
rect 6294 583954 6914 619398
rect 6294 583718 6326 583954
rect 6562 583718 6646 583954
rect 6882 583718 6914 583954
rect 6294 583634 6914 583718
rect 6294 583398 6326 583634
rect 6562 583398 6646 583634
rect 6882 583398 6914 583634
rect 6294 547954 6914 583398
rect 6294 547718 6326 547954
rect 6562 547718 6646 547954
rect 6882 547718 6914 547954
rect 6294 547634 6914 547718
rect 6294 547398 6326 547634
rect 6562 547398 6646 547634
rect 6882 547398 6914 547634
rect 6294 511954 6914 547398
rect 6294 511718 6326 511954
rect 6562 511718 6646 511954
rect 6882 511718 6914 511954
rect 6294 511634 6914 511718
rect 6294 511398 6326 511634
rect 6562 511398 6646 511634
rect 6882 511398 6914 511634
rect 6294 475954 6914 511398
rect 6294 475718 6326 475954
rect 6562 475718 6646 475954
rect 6882 475718 6914 475954
rect 6294 475634 6914 475718
rect 6294 475398 6326 475634
rect 6562 475398 6646 475634
rect 6882 475398 6914 475634
rect 6294 439954 6914 475398
rect 6294 439718 6326 439954
rect 6562 439718 6646 439954
rect 6882 439718 6914 439954
rect 6294 439634 6914 439718
rect 6294 439398 6326 439634
rect 6562 439398 6646 439634
rect 6882 439398 6914 439634
rect 6294 403954 6914 439398
rect 6294 403718 6326 403954
rect 6562 403718 6646 403954
rect 6882 403718 6914 403954
rect 6294 403634 6914 403718
rect 6294 403398 6326 403634
rect 6562 403398 6646 403634
rect 6882 403398 6914 403634
rect 6294 367954 6914 403398
rect 6294 367718 6326 367954
rect 6562 367718 6646 367954
rect 6882 367718 6914 367954
rect 6294 367634 6914 367718
rect 6294 367398 6326 367634
rect 6562 367398 6646 367634
rect 6882 367398 6914 367634
rect 6294 331954 6914 367398
rect 6294 331718 6326 331954
rect 6562 331718 6646 331954
rect 6882 331718 6914 331954
rect 6294 331634 6914 331718
rect 6294 331398 6326 331634
rect 6562 331398 6646 331634
rect 6882 331398 6914 331634
rect 6294 295954 6914 331398
rect 6294 295718 6326 295954
rect 6562 295718 6646 295954
rect 6882 295718 6914 295954
rect 6294 295634 6914 295718
rect 6294 295398 6326 295634
rect 6562 295398 6646 295634
rect 6882 295398 6914 295634
rect 6294 259954 6914 295398
rect 6294 259718 6326 259954
rect 6562 259718 6646 259954
rect 6882 259718 6914 259954
rect 6294 259634 6914 259718
rect 6294 259398 6326 259634
rect 6562 259398 6646 259634
rect 6882 259398 6914 259634
rect 6294 223954 6914 259398
rect 6294 223718 6326 223954
rect 6562 223718 6646 223954
rect 6882 223718 6914 223954
rect 6294 223634 6914 223718
rect 6294 223398 6326 223634
rect 6562 223398 6646 223634
rect 6882 223398 6914 223634
rect 6294 187954 6914 223398
rect 6294 187718 6326 187954
rect 6562 187718 6646 187954
rect 6882 187718 6914 187954
rect 6294 187634 6914 187718
rect 6294 187398 6326 187634
rect 6562 187398 6646 187634
rect 6882 187398 6914 187634
rect 6294 151954 6914 187398
rect 6294 151718 6326 151954
rect 6562 151718 6646 151954
rect 6882 151718 6914 151954
rect 6294 151634 6914 151718
rect 6294 151398 6326 151634
rect 6562 151398 6646 151634
rect 6882 151398 6914 151634
rect 6294 115954 6914 151398
rect 6294 115718 6326 115954
rect 6562 115718 6646 115954
rect 6882 115718 6914 115954
rect 6294 115634 6914 115718
rect 6294 115398 6326 115634
rect 6562 115398 6646 115634
rect 6882 115398 6914 115634
rect 6294 79954 6914 115398
rect 6294 79718 6326 79954
rect 6562 79718 6646 79954
rect 6882 79718 6914 79954
rect 6294 79634 6914 79718
rect 6294 79398 6326 79634
rect 6562 79398 6646 79634
rect 6882 79398 6914 79634
rect 6294 43954 6914 79398
rect 6294 43718 6326 43954
rect 6562 43718 6646 43954
rect 6882 43718 6914 43954
rect 6294 43634 6914 43718
rect 6294 43398 6326 43634
rect 6562 43398 6646 43634
rect 6882 43398 6914 43634
rect 6294 7954 6914 43398
rect 6294 7718 6326 7954
rect 6562 7718 6646 7954
rect 6882 7718 6914 7954
rect 6294 7634 6914 7718
rect 6294 7398 6326 7634
rect 6562 7398 6646 7634
rect 6882 7398 6914 7634
rect 6294 -1306 6914 7398
rect 6294 -1542 6326 -1306
rect 6562 -1542 6646 -1306
rect 6882 -1542 6914 -1306
rect 6294 -1626 6914 -1542
rect 6294 -1862 6326 -1626
rect 6562 -1862 6646 -1626
rect 6882 -1862 6914 -1626
rect 6294 -7654 6914 -1862
rect 10794 706758 11414 711590
rect 10794 706522 10826 706758
rect 11062 706522 11146 706758
rect 11382 706522 11414 706758
rect 10794 706438 11414 706522
rect 10794 706202 10826 706438
rect 11062 706202 11146 706438
rect 11382 706202 11414 706438
rect 10794 696454 11414 706202
rect 10794 696218 10826 696454
rect 11062 696218 11146 696454
rect 11382 696218 11414 696454
rect 10794 696134 11414 696218
rect 10794 695898 10826 696134
rect 11062 695898 11146 696134
rect 11382 695898 11414 696134
rect 10794 660454 11414 695898
rect 10794 660218 10826 660454
rect 11062 660218 11146 660454
rect 11382 660218 11414 660454
rect 10794 660134 11414 660218
rect 10794 659898 10826 660134
rect 11062 659898 11146 660134
rect 11382 659898 11414 660134
rect 10794 624454 11414 659898
rect 10794 624218 10826 624454
rect 11062 624218 11146 624454
rect 11382 624218 11414 624454
rect 10794 624134 11414 624218
rect 10794 623898 10826 624134
rect 11062 623898 11146 624134
rect 11382 623898 11414 624134
rect 10794 588454 11414 623898
rect 10794 588218 10826 588454
rect 11062 588218 11146 588454
rect 11382 588218 11414 588454
rect 10794 588134 11414 588218
rect 10794 587898 10826 588134
rect 11062 587898 11146 588134
rect 11382 587898 11414 588134
rect 10794 552454 11414 587898
rect 10794 552218 10826 552454
rect 11062 552218 11146 552454
rect 11382 552218 11414 552454
rect 10794 552134 11414 552218
rect 10794 551898 10826 552134
rect 11062 551898 11146 552134
rect 11382 551898 11414 552134
rect 10794 516454 11414 551898
rect 10794 516218 10826 516454
rect 11062 516218 11146 516454
rect 11382 516218 11414 516454
rect 10794 516134 11414 516218
rect 10794 515898 10826 516134
rect 11062 515898 11146 516134
rect 11382 515898 11414 516134
rect 10794 480454 11414 515898
rect 10794 480218 10826 480454
rect 11062 480218 11146 480454
rect 11382 480218 11414 480454
rect 10794 480134 11414 480218
rect 10794 479898 10826 480134
rect 11062 479898 11146 480134
rect 11382 479898 11414 480134
rect 10794 444454 11414 479898
rect 10794 444218 10826 444454
rect 11062 444218 11146 444454
rect 11382 444218 11414 444454
rect 10794 444134 11414 444218
rect 10794 443898 10826 444134
rect 11062 443898 11146 444134
rect 11382 443898 11414 444134
rect 10794 408454 11414 443898
rect 10794 408218 10826 408454
rect 11062 408218 11146 408454
rect 11382 408218 11414 408454
rect 10794 408134 11414 408218
rect 10794 407898 10826 408134
rect 11062 407898 11146 408134
rect 11382 407898 11414 408134
rect 10794 372454 11414 407898
rect 10794 372218 10826 372454
rect 11062 372218 11146 372454
rect 11382 372218 11414 372454
rect 10794 372134 11414 372218
rect 10794 371898 10826 372134
rect 11062 371898 11146 372134
rect 11382 371898 11414 372134
rect 10794 336454 11414 371898
rect 10794 336218 10826 336454
rect 11062 336218 11146 336454
rect 11382 336218 11414 336454
rect 10794 336134 11414 336218
rect 10794 335898 10826 336134
rect 11062 335898 11146 336134
rect 11382 335898 11414 336134
rect 10794 300454 11414 335898
rect 10794 300218 10826 300454
rect 11062 300218 11146 300454
rect 11382 300218 11414 300454
rect 10794 300134 11414 300218
rect 10794 299898 10826 300134
rect 11062 299898 11146 300134
rect 11382 299898 11414 300134
rect 10794 264454 11414 299898
rect 10794 264218 10826 264454
rect 11062 264218 11146 264454
rect 11382 264218 11414 264454
rect 10794 264134 11414 264218
rect 10794 263898 10826 264134
rect 11062 263898 11146 264134
rect 11382 263898 11414 264134
rect 10794 228454 11414 263898
rect 10794 228218 10826 228454
rect 11062 228218 11146 228454
rect 11382 228218 11414 228454
rect 10794 228134 11414 228218
rect 10794 227898 10826 228134
rect 11062 227898 11146 228134
rect 11382 227898 11414 228134
rect 10794 192454 11414 227898
rect 10794 192218 10826 192454
rect 11062 192218 11146 192454
rect 11382 192218 11414 192454
rect 10794 192134 11414 192218
rect 10794 191898 10826 192134
rect 11062 191898 11146 192134
rect 11382 191898 11414 192134
rect 10794 156454 11414 191898
rect 10794 156218 10826 156454
rect 11062 156218 11146 156454
rect 11382 156218 11414 156454
rect 10794 156134 11414 156218
rect 10794 155898 10826 156134
rect 11062 155898 11146 156134
rect 11382 155898 11414 156134
rect 10794 120454 11414 155898
rect 10794 120218 10826 120454
rect 11062 120218 11146 120454
rect 11382 120218 11414 120454
rect 10794 120134 11414 120218
rect 10794 119898 10826 120134
rect 11062 119898 11146 120134
rect 11382 119898 11414 120134
rect 10794 84454 11414 119898
rect 10794 84218 10826 84454
rect 11062 84218 11146 84454
rect 11382 84218 11414 84454
rect 10794 84134 11414 84218
rect 10794 83898 10826 84134
rect 11062 83898 11146 84134
rect 11382 83898 11414 84134
rect 10794 48454 11414 83898
rect 10794 48218 10826 48454
rect 11062 48218 11146 48454
rect 11382 48218 11414 48454
rect 10794 48134 11414 48218
rect 10794 47898 10826 48134
rect 11062 47898 11146 48134
rect 11382 47898 11414 48134
rect 10794 12454 11414 47898
rect 10794 12218 10826 12454
rect 11062 12218 11146 12454
rect 11382 12218 11414 12454
rect 10794 12134 11414 12218
rect 10794 11898 10826 12134
rect 11062 11898 11146 12134
rect 11382 11898 11414 12134
rect 10794 -2266 11414 11898
rect 10794 -2502 10826 -2266
rect 11062 -2502 11146 -2266
rect 11382 -2502 11414 -2266
rect 10794 -2586 11414 -2502
rect 10794 -2822 10826 -2586
rect 11062 -2822 11146 -2586
rect 11382 -2822 11414 -2586
rect 10794 -7654 11414 -2822
rect 15294 707718 15914 711590
rect 15294 707482 15326 707718
rect 15562 707482 15646 707718
rect 15882 707482 15914 707718
rect 15294 707398 15914 707482
rect 15294 707162 15326 707398
rect 15562 707162 15646 707398
rect 15882 707162 15914 707398
rect 15294 700954 15914 707162
rect 15294 700718 15326 700954
rect 15562 700718 15646 700954
rect 15882 700718 15914 700954
rect 15294 700634 15914 700718
rect 15294 700398 15326 700634
rect 15562 700398 15646 700634
rect 15882 700398 15914 700634
rect 15294 664954 15914 700398
rect 15294 664718 15326 664954
rect 15562 664718 15646 664954
rect 15882 664718 15914 664954
rect 15294 664634 15914 664718
rect 15294 664398 15326 664634
rect 15562 664398 15646 664634
rect 15882 664398 15914 664634
rect 15294 628954 15914 664398
rect 15294 628718 15326 628954
rect 15562 628718 15646 628954
rect 15882 628718 15914 628954
rect 15294 628634 15914 628718
rect 15294 628398 15326 628634
rect 15562 628398 15646 628634
rect 15882 628398 15914 628634
rect 15294 592954 15914 628398
rect 15294 592718 15326 592954
rect 15562 592718 15646 592954
rect 15882 592718 15914 592954
rect 15294 592634 15914 592718
rect 15294 592398 15326 592634
rect 15562 592398 15646 592634
rect 15882 592398 15914 592634
rect 15294 556954 15914 592398
rect 15294 556718 15326 556954
rect 15562 556718 15646 556954
rect 15882 556718 15914 556954
rect 15294 556634 15914 556718
rect 15294 556398 15326 556634
rect 15562 556398 15646 556634
rect 15882 556398 15914 556634
rect 15294 520954 15914 556398
rect 15294 520718 15326 520954
rect 15562 520718 15646 520954
rect 15882 520718 15914 520954
rect 15294 520634 15914 520718
rect 15294 520398 15326 520634
rect 15562 520398 15646 520634
rect 15882 520398 15914 520634
rect 15294 484954 15914 520398
rect 15294 484718 15326 484954
rect 15562 484718 15646 484954
rect 15882 484718 15914 484954
rect 15294 484634 15914 484718
rect 15294 484398 15326 484634
rect 15562 484398 15646 484634
rect 15882 484398 15914 484634
rect 15294 448954 15914 484398
rect 15294 448718 15326 448954
rect 15562 448718 15646 448954
rect 15882 448718 15914 448954
rect 15294 448634 15914 448718
rect 15294 448398 15326 448634
rect 15562 448398 15646 448634
rect 15882 448398 15914 448634
rect 15294 412954 15914 448398
rect 15294 412718 15326 412954
rect 15562 412718 15646 412954
rect 15882 412718 15914 412954
rect 15294 412634 15914 412718
rect 15294 412398 15326 412634
rect 15562 412398 15646 412634
rect 15882 412398 15914 412634
rect 15294 376954 15914 412398
rect 15294 376718 15326 376954
rect 15562 376718 15646 376954
rect 15882 376718 15914 376954
rect 15294 376634 15914 376718
rect 15294 376398 15326 376634
rect 15562 376398 15646 376634
rect 15882 376398 15914 376634
rect 15294 340954 15914 376398
rect 15294 340718 15326 340954
rect 15562 340718 15646 340954
rect 15882 340718 15914 340954
rect 15294 340634 15914 340718
rect 15294 340398 15326 340634
rect 15562 340398 15646 340634
rect 15882 340398 15914 340634
rect 15294 304954 15914 340398
rect 15294 304718 15326 304954
rect 15562 304718 15646 304954
rect 15882 304718 15914 304954
rect 15294 304634 15914 304718
rect 15294 304398 15326 304634
rect 15562 304398 15646 304634
rect 15882 304398 15914 304634
rect 15294 268954 15914 304398
rect 15294 268718 15326 268954
rect 15562 268718 15646 268954
rect 15882 268718 15914 268954
rect 15294 268634 15914 268718
rect 15294 268398 15326 268634
rect 15562 268398 15646 268634
rect 15882 268398 15914 268634
rect 15294 232954 15914 268398
rect 15294 232718 15326 232954
rect 15562 232718 15646 232954
rect 15882 232718 15914 232954
rect 15294 232634 15914 232718
rect 15294 232398 15326 232634
rect 15562 232398 15646 232634
rect 15882 232398 15914 232634
rect 15294 196954 15914 232398
rect 15294 196718 15326 196954
rect 15562 196718 15646 196954
rect 15882 196718 15914 196954
rect 15294 196634 15914 196718
rect 15294 196398 15326 196634
rect 15562 196398 15646 196634
rect 15882 196398 15914 196634
rect 15294 160954 15914 196398
rect 15294 160718 15326 160954
rect 15562 160718 15646 160954
rect 15882 160718 15914 160954
rect 15294 160634 15914 160718
rect 15294 160398 15326 160634
rect 15562 160398 15646 160634
rect 15882 160398 15914 160634
rect 15294 124954 15914 160398
rect 15294 124718 15326 124954
rect 15562 124718 15646 124954
rect 15882 124718 15914 124954
rect 15294 124634 15914 124718
rect 15294 124398 15326 124634
rect 15562 124398 15646 124634
rect 15882 124398 15914 124634
rect 15294 88954 15914 124398
rect 15294 88718 15326 88954
rect 15562 88718 15646 88954
rect 15882 88718 15914 88954
rect 15294 88634 15914 88718
rect 15294 88398 15326 88634
rect 15562 88398 15646 88634
rect 15882 88398 15914 88634
rect 15294 52954 15914 88398
rect 15294 52718 15326 52954
rect 15562 52718 15646 52954
rect 15882 52718 15914 52954
rect 15294 52634 15914 52718
rect 15294 52398 15326 52634
rect 15562 52398 15646 52634
rect 15882 52398 15914 52634
rect 15294 16954 15914 52398
rect 15294 16718 15326 16954
rect 15562 16718 15646 16954
rect 15882 16718 15914 16954
rect 15294 16634 15914 16718
rect 15294 16398 15326 16634
rect 15562 16398 15646 16634
rect 15882 16398 15914 16634
rect 15294 -3226 15914 16398
rect 15294 -3462 15326 -3226
rect 15562 -3462 15646 -3226
rect 15882 -3462 15914 -3226
rect 15294 -3546 15914 -3462
rect 15294 -3782 15326 -3546
rect 15562 -3782 15646 -3546
rect 15882 -3782 15914 -3546
rect 15294 -7654 15914 -3782
rect 19794 708678 20414 711590
rect 19794 708442 19826 708678
rect 20062 708442 20146 708678
rect 20382 708442 20414 708678
rect 19794 708358 20414 708442
rect 19794 708122 19826 708358
rect 20062 708122 20146 708358
rect 20382 708122 20414 708358
rect 19794 669454 20414 708122
rect 19794 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 20414 669454
rect 19794 669134 20414 669218
rect 19794 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 20414 669134
rect 19794 633454 20414 668898
rect 19794 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 20414 633454
rect 19794 633134 20414 633218
rect 19794 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 20414 633134
rect 19794 597454 20414 632898
rect 19794 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 20414 597454
rect 19794 597134 20414 597218
rect 19794 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 20414 597134
rect 19794 561454 20414 596898
rect 19794 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 20414 561454
rect 19794 561134 20414 561218
rect 19794 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 20414 561134
rect 19794 525454 20414 560898
rect 19794 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 20414 525454
rect 19794 525134 20414 525218
rect 19794 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 20414 525134
rect 19794 489454 20414 524898
rect 19794 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 20414 489454
rect 19794 489134 20414 489218
rect 19794 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 20414 489134
rect 19794 453454 20414 488898
rect 19794 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 20414 453454
rect 19794 453134 20414 453218
rect 19794 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 20414 453134
rect 19794 417454 20414 452898
rect 19794 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 20414 417454
rect 19794 417134 20414 417218
rect 19794 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 20414 417134
rect 19794 381454 20414 416898
rect 19794 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 20414 381454
rect 19794 381134 20414 381218
rect 19794 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 20414 381134
rect 19794 345454 20414 380898
rect 19794 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 20414 345454
rect 19794 345134 20414 345218
rect 19794 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 20414 345134
rect 19794 309454 20414 344898
rect 19794 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 20414 309454
rect 19794 309134 20414 309218
rect 19794 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 20414 309134
rect 19794 273454 20414 308898
rect 19794 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 20414 273454
rect 19794 273134 20414 273218
rect 19794 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 20414 273134
rect 19794 237454 20414 272898
rect 19794 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 20414 237454
rect 19794 237134 20414 237218
rect 19794 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 20414 237134
rect 19794 201454 20414 236898
rect 19794 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 20414 201454
rect 19794 201134 20414 201218
rect 19794 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 20414 201134
rect 19794 165454 20414 200898
rect 19794 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 20414 165454
rect 19794 165134 20414 165218
rect 19794 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 20414 165134
rect 19794 129454 20414 164898
rect 19794 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 20414 129454
rect 19794 129134 20414 129218
rect 19794 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 20414 129134
rect 19794 93454 20414 128898
rect 19794 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 20414 93454
rect 19794 93134 20414 93218
rect 19794 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 20414 93134
rect 19794 57454 20414 92898
rect 19794 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 20414 57454
rect 19794 57134 20414 57218
rect 19794 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 20414 57134
rect 19794 21454 20414 56898
rect 19794 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 20414 21454
rect 19794 21134 20414 21218
rect 19794 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 20414 21134
rect 19794 -4186 20414 20898
rect 19794 -4422 19826 -4186
rect 20062 -4422 20146 -4186
rect 20382 -4422 20414 -4186
rect 19794 -4506 20414 -4422
rect 19794 -4742 19826 -4506
rect 20062 -4742 20146 -4506
rect 20382 -4742 20414 -4506
rect 19794 -7654 20414 -4742
rect 24294 709638 24914 711590
rect 24294 709402 24326 709638
rect 24562 709402 24646 709638
rect 24882 709402 24914 709638
rect 24294 709318 24914 709402
rect 24294 709082 24326 709318
rect 24562 709082 24646 709318
rect 24882 709082 24914 709318
rect 24294 673954 24914 709082
rect 24294 673718 24326 673954
rect 24562 673718 24646 673954
rect 24882 673718 24914 673954
rect 24294 673634 24914 673718
rect 24294 673398 24326 673634
rect 24562 673398 24646 673634
rect 24882 673398 24914 673634
rect 24294 637954 24914 673398
rect 24294 637718 24326 637954
rect 24562 637718 24646 637954
rect 24882 637718 24914 637954
rect 24294 637634 24914 637718
rect 24294 637398 24326 637634
rect 24562 637398 24646 637634
rect 24882 637398 24914 637634
rect 24294 601954 24914 637398
rect 24294 601718 24326 601954
rect 24562 601718 24646 601954
rect 24882 601718 24914 601954
rect 24294 601634 24914 601718
rect 24294 601398 24326 601634
rect 24562 601398 24646 601634
rect 24882 601398 24914 601634
rect 24294 565954 24914 601398
rect 24294 565718 24326 565954
rect 24562 565718 24646 565954
rect 24882 565718 24914 565954
rect 24294 565634 24914 565718
rect 24294 565398 24326 565634
rect 24562 565398 24646 565634
rect 24882 565398 24914 565634
rect 24294 529954 24914 565398
rect 24294 529718 24326 529954
rect 24562 529718 24646 529954
rect 24882 529718 24914 529954
rect 24294 529634 24914 529718
rect 24294 529398 24326 529634
rect 24562 529398 24646 529634
rect 24882 529398 24914 529634
rect 24294 493954 24914 529398
rect 24294 493718 24326 493954
rect 24562 493718 24646 493954
rect 24882 493718 24914 493954
rect 24294 493634 24914 493718
rect 24294 493398 24326 493634
rect 24562 493398 24646 493634
rect 24882 493398 24914 493634
rect 24294 457954 24914 493398
rect 24294 457718 24326 457954
rect 24562 457718 24646 457954
rect 24882 457718 24914 457954
rect 24294 457634 24914 457718
rect 24294 457398 24326 457634
rect 24562 457398 24646 457634
rect 24882 457398 24914 457634
rect 24294 421954 24914 457398
rect 24294 421718 24326 421954
rect 24562 421718 24646 421954
rect 24882 421718 24914 421954
rect 24294 421634 24914 421718
rect 24294 421398 24326 421634
rect 24562 421398 24646 421634
rect 24882 421398 24914 421634
rect 24294 385954 24914 421398
rect 24294 385718 24326 385954
rect 24562 385718 24646 385954
rect 24882 385718 24914 385954
rect 24294 385634 24914 385718
rect 24294 385398 24326 385634
rect 24562 385398 24646 385634
rect 24882 385398 24914 385634
rect 24294 349954 24914 385398
rect 24294 349718 24326 349954
rect 24562 349718 24646 349954
rect 24882 349718 24914 349954
rect 24294 349634 24914 349718
rect 24294 349398 24326 349634
rect 24562 349398 24646 349634
rect 24882 349398 24914 349634
rect 24294 313954 24914 349398
rect 24294 313718 24326 313954
rect 24562 313718 24646 313954
rect 24882 313718 24914 313954
rect 24294 313634 24914 313718
rect 24294 313398 24326 313634
rect 24562 313398 24646 313634
rect 24882 313398 24914 313634
rect 24294 277954 24914 313398
rect 24294 277718 24326 277954
rect 24562 277718 24646 277954
rect 24882 277718 24914 277954
rect 24294 277634 24914 277718
rect 24294 277398 24326 277634
rect 24562 277398 24646 277634
rect 24882 277398 24914 277634
rect 24294 241954 24914 277398
rect 24294 241718 24326 241954
rect 24562 241718 24646 241954
rect 24882 241718 24914 241954
rect 24294 241634 24914 241718
rect 24294 241398 24326 241634
rect 24562 241398 24646 241634
rect 24882 241398 24914 241634
rect 24294 205954 24914 241398
rect 24294 205718 24326 205954
rect 24562 205718 24646 205954
rect 24882 205718 24914 205954
rect 24294 205634 24914 205718
rect 24294 205398 24326 205634
rect 24562 205398 24646 205634
rect 24882 205398 24914 205634
rect 24294 169954 24914 205398
rect 24294 169718 24326 169954
rect 24562 169718 24646 169954
rect 24882 169718 24914 169954
rect 24294 169634 24914 169718
rect 24294 169398 24326 169634
rect 24562 169398 24646 169634
rect 24882 169398 24914 169634
rect 24294 133954 24914 169398
rect 24294 133718 24326 133954
rect 24562 133718 24646 133954
rect 24882 133718 24914 133954
rect 24294 133634 24914 133718
rect 24294 133398 24326 133634
rect 24562 133398 24646 133634
rect 24882 133398 24914 133634
rect 24294 97954 24914 133398
rect 24294 97718 24326 97954
rect 24562 97718 24646 97954
rect 24882 97718 24914 97954
rect 24294 97634 24914 97718
rect 24294 97398 24326 97634
rect 24562 97398 24646 97634
rect 24882 97398 24914 97634
rect 24294 61954 24914 97398
rect 24294 61718 24326 61954
rect 24562 61718 24646 61954
rect 24882 61718 24914 61954
rect 24294 61634 24914 61718
rect 24294 61398 24326 61634
rect 24562 61398 24646 61634
rect 24882 61398 24914 61634
rect 24294 25954 24914 61398
rect 24294 25718 24326 25954
rect 24562 25718 24646 25954
rect 24882 25718 24914 25954
rect 24294 25634 24914 25718
rect 24294 25398 24326 25634
rect 24562 25398 24646 25634
rect 24882 25398 24914 25634
rect 24294 -5146 24914 25398
rect 24294 -5382 24326 -5146
rect 24562 -5382 24646 -5146
rect 24882 -5382 24914 -5146
rect 24294 -5466 24914 -5382
rect 24294 -5702 24326 -5466
rect 24562 -5702 24646 -5466
rect 24882 -5702 24914 -5466
rect 24294 -7654 24914 -5702
rect 28794 710598 29414 711590
rect 28794 710362 28826 710598
rect 29062 710362 29146 710598
rect 29382 710362 29414 710598
rect 28794 710278 29414 710362
rect 28794 710042 28826 710278
rect 29062 710042 29146 710278
rect 29382 710042 29414 710278
rect 28794 678454 29414 710042
rect 28794 678218 28826 678454
rect 29062 678218 29146 678454
rect 29382 678218 29414 678454
rect 28794 678134 29414 678218
rect 28794 677898 28826 678134
rect 29062 677898 29146 678134
rect 29382 677898 29414 678134
rect 28794 642454 29414 677898
rect 28794 642218 28826 642454
rect 29062 642218 29146 642454
rect 29382 642218 29414 642454
rect 28794 642134 29414 642218
rect 28794 641898 28826 642134
rect 29062 641898 29146 642134
rect 29382 641898 29414 642134
rect 28794 606454 29414 641898
rect 28794 606218 28826 606454
rect 29062 606218 29146 606454
rect 29382 606218 29414 606454
rect 28794 606134 29414 606218
rect 28794 605898 28826 606134
rect 29062 605898 29146 606134
rect 29382 605898 29414 606134
rect 28794 570454 29414 605898
rect 28794 570218 28826 570454
rect 29062 570218 29146 570454
rect 29382 570218 29414 570454
rect 28794 570134 29414 570218
rect 28794 569898 28826 570134
rect 29062 569898 29146 570134
rect 29382 569898 29414 570134
rect 28794 534454 29414 569898
rect 28794 534218 28826 534454
rect 29062 534218 29146 534454
rect 29382 534218 29414 534454
rect 28794 534134 29414 534218
rect 28794 533898 28826 534134
rect 29062 533898 29146 534134
rect 29382 533898 29414 534134
rect 28794 498454 29414 533898
rect 28794 498218 28826 498454
rect 29062 498218 29146 498454
rect 29382 498218 29414 498454
rect 28794 498134 29414 498218
rect 28794 497898 28826 498134
rect 29062 497898 29146 498134
rect 29382 497898 29414 498134
rect 28794 462454 29414 497898
rect 28794 462218 28826 462454
rect 29062 462218 29146 462454
rect 29382 462218 29414 462454
rect 28794 462134 29414 462218
rect 28794 461898 28826 462134
rect 29062 461898 29146 462134
rect 29382 461898 29414 462134
rect 28794 426454 29414 461898
rect 28794 426218 28826 426454
rect 29062 426218 29146 426454
rect 29382 426218 29414 426454
rect 28794 426134 29414 426218
rect 28794 425898 28826 426134
rect 29062 425898 29146 426134
rect 29382 425898 29414 426134
rect 28794 390454 29414 425898
rect 28794 390218 28826 390454
rect 29062 390218 29146 390454
rect 29382 390218 29414 390454
rect 28794 390134 29414 390218
rect 28794 389898 28826 390134
rect 29062 389898 29146 390134
rect 29382 389898 29414 390134
rect 28794 354454 29414 389898
rect 28794 354218 28826 354454
rect 29062 354218 29146 354454
rect 29382 354218 29414 354454
rect 28794 354134 29414 354218
rect 28794 353898 28826 354134
rect 29062 353898 29146 354134
rect 29382 353898 29414 354134
rect 28794 318454 29414 353898
rect 28794 318218 28826 318454
rect 29062 318218 29146 318454
rect 29382 318218 29414 318454
rect 28794 318134 29414 318218
rect 28794 317898 28826 318134
rect 29062 317898 29146 318134
rect 29382 317898 29414 318134
rect 28794 282454 29414 317898
rect 28794 282218 28826 282454
rect 29062 282218 29146 282454
rect 29382 282218 29414 282454
rect 28794 282134 29414 282218
rect 28794 281898 28826 282134
rect 29062 281898 29146 282134
rect 29382 281898 29414 282134
rect 28794 246454 29414 281898
rect 28794 246218 28826 246454
rect 29062 246218 29146 246454
rect 29382 246218 29414 246454
rect 28794 246134 29414 246218
rect 28794 245898 28826 246134
rect 29062 245898 29146 246134
rect 29382 245898 29414 246134
rect 28794 210454 29414 245898
rect 28794 210218 28826 210454
rect 29062 210218 29146 210454
rect 29382 210218 29414 210454
rect 28794 210134 29414 210218
rect 28794 209898 28826 210134
rect 29062 209898 29146 210134
rect 29382 209898 29414 210134
rect 28794 174454 29414 209898
rect 28794 174218 28826 174454
rect 29062 174218 29146 174454
rect 29382 174218 29414 174454
rect 28794 174134 29414 174218
rect 28794 173898 28826 174134
rect 29062 173898 29146 174134
rect 29382 173898 29414 174134
rect 28794 138454 29414 173898
rect 28794 138218 28826 138454
rect 29062 138218 29146 138454
rect 29382 138218 29414 138454
rect 28794 138134 29414 138218
rect 28794 137898 28826 138134
rect 29062 137898 29146 138134
rect 29382 137898 29414 138134
rect 28794 102454 29414 137898
rect 28794 102218 28826 102454
rect 29062 102218 29146 102454
rect 29382 102218 29414 102454
rect 28794 102134 29414 102218
rect 28794 101898 28826 102134
rect 29062 101898 29146 102134
rect 29382 101898 29414 102134
rect 28794 66454 29414 101898
rect 28794 66218 28826 66454
rect 29062 66218 29146 66454
rect 29382 66218 29414 66454
rect 28794 66134 29414 66218
rect 28794 65898 28826 66134
rect 29062 65898 29146 66134
rect 29382 65898 29414 66134
rect 28794 30454 29414 65898
rect 28794 30218 28826 30454
rect 29062 30218 29146 30454
rect 29382 30218 29414 30454
rect 28794 30134 29414 30218
rect 28794 29898 28826 30134
rect 29062 29898 29146 30134
rect 29382 29898 29414 30134
rect 28794 -6106 29414 29898
rect 28794 -6342 28826 -6106
rect 29062 -6342 29146 -6106
rect 29382 -6342 29414 -6106
rect 28794 -6426 29414 -6342
rect 28794 -6662 28826 -6426
rect 29062 -6662 29146 -6426
rect 29382 -6662 29414 -6426
rect 28794 -7654 29414 -6662
rect 33294 711558 33914 711590
rect 33294 711322 33326 711558
rect 33562 711322 33646 711558
rect 33882 711322 33914 711558
rect 33294 711238 33914 711322
rect 33294 711002 33326 711238
rect 33562 711002 33646 711238
rect 33882 711002 33914 711238
rect 33294 682954 33914 711002
rect 33294 682718 33326 682954
rect 33562 682718 33646 682954
rect 33882 682718 33914 682954
rect 33294 682634 33914 682718
rect 33294 682398 33326 682634
rect 33562 682398 33646 682634
rect 33882 682398 33914 682634
rect 33294 646954 33914 682398
rect 33294 646718 33326 646954
rect 33562 646718 33646 646954
rect 33882 646718 33914 646954
rect 33294 646634 33914 646718
rect 33294 646398 33326 646634
rect 33562 646398 33646 646634
rect 33882 646398 33914 646634
rect 33294 610954 33914 646398
rect 33294 610718 33326 610954
rect 33562 610718 33646 610954
rect 33882 610718 33914 610954
rect 33294 610634 33914 610718
rect 33294 610398 33326 610634
rect 33562 610398 33646 610634
rect 33882 610398 33914 610634
rect 33294 574954 33914 610398
rect 33294 574718 33326 574954
rect 33562 574718 33646 574954
rect 33882 574718 33914 574954
rect 33294 574634 33914 574718
rect 33294 574398 33326 574634
rect 33562 574398 33646 574634
rect 33882 574398 33914 574634
rect 33294 538954 33914 574398
rect 33294 538718 33326 538954
rect 33562 538718 33646 538954
rect 33882 538718 33914 538954
rect 33294 538634 33914 538718
rect 33294 538398 33326 538634
rect 33562 538398 33646 538634
rect 33882 538398 33914 538634
rect 33294 502954 33914 538398
rect 33294 502718 33326 502954
rect 33562 502718 33646 502954
rect 33882 502718 33914 502954
rect 33294 502634 33914 502718
rect 33294 502398 33326 502634
rect 33562 502398 33646 502634
rect 33882 502398 33914 502634
rect 33294 466954 33914 502398
rect 33294 466718 33326 466954
rect 33562 466718 33646 466954
rect 33882 466718 33914 466954
rect 33294 466634 33914 466718
rect 33294 466398 33326 466634
rect 33562 466398 33646 466634
rect 33882 466398 33914 466634
rect 33294 430954 33914 466398
rect 33294 430718 33326 430954
rect 33562 430718 33646 430954
rect 33882 430718 33914 430954
rect 33294 430634 33914 430718
rect 33294 430398 33326 430634
rect 33562 430398 33646 430634
rect 33882 430398 33914 430634
rect 33294 394954 33914 430398
rect 33294 394718 33326 394954
rect 33562 394718 33646 394954
rect 33882 394718 33914 394954
rect 33294 394634 33914 394718
rect 33294 394398 33326 394634
rect 33562 394398 33646 394634
rect 33882 394398 33914 394634
rect 33294 358954 33914 394398
rect 33294 358718 33326 358954
rect 33562 358718 33646 358954
rect 33882 358718 33914 358954
rect 33294 358634 33914 358718
rect 33294 358398 33326 358634
rect 33562 358398 33646 358634
rect 33882 358398 33914 358634
rect 33294 322954 33914 358398
rect 33294 322718 33326 322954
rect 33562 322718 33646 322954
rect 33882 322718 33914 322954
rect 33294 322634 33914 322718
rect 33294 322398 33326 322634
rect 33562 322398 33646 322634
rect 33882 322398 33914 322634
rect 33294 286954 33914 322398
rect 33294 286718 33326 286954
rect 33562 286718 33646 286954
rect 33882 286718 33914 286954
rect 33294 286634 33914 286718
rect 33294 286398 33326 286634
rect 33562 286398 33646 286634
rect 33882 286398 33914 286634
rect 33294 250954 33914 286398
rect 33294 250718 33326 250954
rect 33562 250718 33646 250954
rect 33882 250718 33914 250954
rect 33294 250634 33914 250718
rect 33294 250398 33326 250634
rect 33562 250398 33646 250634
rect 33882 250398 33914 250634
rect 33294 214954 33914 250398
rect 33294 214718 33326 214954
rect 33562 214718 33646 214954
rect 33882 214718 33914 214954
rect 33294 214634 33914 214718
rect 33294 214398 33326 214634
rect 33562 214398 33646 214634
rect 33882 214398 33914 214634
rect 33294 178954 33914 214398
rect 33294 178718 33326 178954
rect 33562 178718 33646 178954
rect 33882 178718 33914 178954
rect 33294 178634 33914 178718
rect 33294 178398 33326 178634
rect 33562 178398 33646 178634
rect 33882 178398 33914 178634
rect 33294 142954 33914 178398
rect 33294 142718 33326 142954
rect 33562 142718 33646 142954
rect 33882 142718 33914 142954
rect 33294 142634 33914 142718
rect 33294 142398 33326 142634
rect 33562 142398 33646 142634
rect 33882 142398 33914 142634
rect 33294 106954 33914 142398
rect 33294 106718 33326 106954
rect 33562 106718 33646 106954
rect 33882 106718 33914 106954
rect 33294 106634 33914 106718
rect 33294 106398 33326 106634
rect 33562 106398 33646 106634
rect 33882 106398 33914 106634
rect 33294 70954 33914 106398
rect 33294 70718 33326 70954
rect 33562 70718 33646 70954
rect 33882 70718 33914 70954
rect 33294 70634 33914 70718
rect 33294 70398 33326 70634
rect 33562 70398 33646 70634
rect 33882 70398 33914 70634
rect 33294 34954 33914 70398
rect 33294 34718 33326 34954
rect 33562 34718 33646 34954
rect 33882 34718 33914 34954
rect 33294 34634 33914 34718
rect 33294 34398 33326 34634
rect 33562 34398 33646 34634
rect 33882 34398 33914 34634
rect 33294 -7066 33914 34398
rect 33294 -7302 33326 -7066
rect 33562 -7302 33646 -7066
rect 33882 -7302 33914 -7066
rect 33294 -7386 33914 -7302
rect 33294 -7622 33326 -7386
rect 33562 -7622 33646 -7386
rect 33882 -7622 33914 -7386
rect 33294 -7654 33914 -7622
rect 37794 704838 38414 711590
rect 37794 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 38414 704838
rect 37794 704518 38414 704602
rect 37794 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 38414 704518
rect 37794 687454 38414 704282
rect 37794 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 38414 687454
rect 37794 687134 38414 687218
rect 37794 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 38414 687134
rect 37794 651454 38414 686898
rect 37794 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 38414 651454
rect 37794 651134 38414 651218
rect 37794 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 38414 651134
rect 37794 615454 38414 650898
rect 37794 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 38414 615454
rect 37794 615134 38414 615218
rect 37794 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 38414 615134
rect 37794 579454 38414 614898
rect 37794 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 38414 579454
rect 37794 579134 38414 579218
rect 37794 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 38414 579134
rect 37794 543454 38414 578898
rect 37794 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 38414 543454
rect 37794 543134 38414 543218
rect 37794 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 38414 543134
rect 37794 507454 38414 542898
rect 37794 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 38414 507454
rect 37794 507134 38414 507218
rect 37794 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 38414 507134
rect 37794 471454 38414 506898
rect 37794 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 38414 471454
rect 37794 471134 38414 471218
rect 37794 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 38414 471134
rect 37794 435454 38414 470898
rect 37794 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 38414 435454
rect 37794 435134 38414 435218
rect 37794 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 38414 435134
rect 37794 399454 38414 434898
rect 37794 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 38414 399454
rect 37794 399134 38414 399218
rect 37794 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 38414 399134
rect 37794 363454 38414 398898
rect 37794 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 38414 363454
rect 37794 363134 38414 363218
rect 37794 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 38414 363134
rect 37794 327454 38414 362898
rect 37794 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 38414 327454
rect 37794 327134 38414 327218
rect 37794 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 38414 327134
rect 37794 291454 38414 326898
rect 37794 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 38414 291454
rect 37794 291134 38414 291218
rect 37794 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 38414 291134
rect 37794 255454 38414 290898
rect 37794 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 38414 255454
rect 37794 255134 38414 255218
rect 37794 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 38414 255134
rect 37794 219454 38414 254898
rect 37794 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 38414 219454
rect 37794 219134 38414 219218
rect 37794 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 38414 219134
rect 37794 183454 38414 218898
rect 37794 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 38414 183454
rect 37794 183134 38414 183218
rect 37794 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 38414 183134
rect 37794 147454 38414 182898
rect 37794 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 38414 147454
rect 37794 147134 38414 147218
rect 37794 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 38414 147134
rect 37794 111454 38414 146898
rect 37794 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 38414 111454
rect 37794 111134 38414 111218
rect 37794 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 38414 111134
rect 37794 75454 38414 110898
rect 37794 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 38414 75454
rect 37794 75134 38414 75218
rect 37794 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 38414 75134
rect 37794 39454 38414 74898
rect 37794 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 38414 39454
rect 37794 39134 38414 39218
rect 37794 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 38414 39134
rect 37794 3454 38414 38898
rect 37794 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 38414 3454
rect 37794 3134 38414 3218
rect 37794 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 38414 3134
rect 37794 -346 38414 2898
rect 37794 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 38414 -346
rect 37794 -666 38414 -582
rect 37794 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 38414 -666
rect 37794 -7654 38414 -902
rect 42294 705798 42914 711590
rect 42294 705562 42326 705798
rect 42562 705562 42646 705798
rect 42882 705562 42914 705798
rect 42294 705478 42914 705562
rect 42294 705242 42326 705478
rect 42562 705242 42646 705478
rect 42882 705242 42914 705478
rect 42294 691954 42914 705242
rect 42294 691718 42326 691954
rect 42562 691718 42646 691954
rect 42882 691718 42914 691954
rect 42294 691634 42914 691718
rect 42294 691398 42326 691634
rect 42562 691398 42646 691634
rect 42882 691398 42914 691634
rect 42294 655954 42914 691398
rect 42294 655718 42326 655954
rect 42562 655718 42646 655954
rect 42882 655718 42914 655954
rect 42294 655634 42914 655718
rect 42294 655398 42326 655634
rect 42562 655398 42646 655634
rect 42882 655398 42914 655634
rect 42294 619954 42914 655398
rect 42294 619718 42326 619954
rect 42562 619718 42646 619954
rect 42882 619718 42914 619954
rect 42294 619634 42914 619718
rect 42294 619398 42326 619634
rect 42562 619398 42646 619634
rect 42882 619398 42914 619634
rect 42294 583954 42914 619398
rect 42294 583718 42326 583954
rect 42562 583718 42646 583954
rect 42882 583718 42914 583954
rect 42294 583634 42914 583718
rect 42294 583398 42326 583634
rect 42562 583398 42646 583634
rect 42882 583398 42914 583634
rect 42294 547954 42914 583398
rect 42294 547718 42326 547954
rect 42562 547718 42646 547954
rect 42882 547718 42914 547954
rect 42294 547634 42914 547718
rect 42294 547398 42326 547634
rect 42562 547398 42646 547634
rect 42882 547398 42914 547634
rect 42294 511954 42914 547398
rect 42294 511718 42326 511954
rect 42562 511718 42646 511954
rect 42882 511718 42914 511954
rect 42294 511634 42914 511718
rect 42294 511398 42326 511634
rect 42562 511398 42646 511634
rect 42882 511398 42914 511634
rect 42294 475954 42914 511398
rect 42294 475718 42326 475954
rect 42562 475718 42646 475954
rect 42882 475718 42914 475954
rect 42294 475634 42914 475718
rect 42294 475398 42326 475634
rect 42562 475398 42646 475634
rect 42882 475398 42914 475634
rect 42294 439954 42914 475398
rect 42294 439718 42326 439954
rect 42562 439718 42646 439954
rect 42882 439718 42914 439954
rect 42294 439634 42914 439718
rect 42294 439398 42326 439634
rect 42562 439398 42646 439634
rect 42882 439398 42914 439634
rect 42294 403954 42914 439398
rect 42294 403718 42326 403954
rect 42562 403718 42646 403954
rect 42882 403718 42914 403954
rect 42294 403634 42914 403718
rect 42294 403398 42326 403634
rect 42562 403398 42646 403634
rect 42882 403398 42914 403634
rect 42294 367954 42914 403398
rect 42294 367718 42326 367954
rect 42562 367718 42646 367954
rect 42882 367718 42914 367954
rect 42294 367634 42914 367718
rect 42294 367398 42326 367634
rect 42562 367398 42646 367634
rect 42882 367398 42914 367634
rect 42294 331954 42914 367398
rect 42294 331718 42326 331954
rect 42562 331718 42646 331954
rect 42882 331718 42914 331954
rect 42294 331634 42914 331718
rect 42294 331398 42326 331634
rect 42562 331398 42646 331634
rect 42882 331398 42914 331634
rect 42294 295954 42914 331398
rect 42294 295718 42326 295954
rect 42562 295718 42646 295954
rect 42882 295718 42914 295954
rect 42294 295634 42914 295718
rect 42294 295398 42326 295634
rect 42562 295398 42646 295634
rect 42882 295398 42914 295634
rect 42294 259954 42914 295398
rect 42294 259718 42326 259954
rect 42562 259718 42646 259954
rect 42882 259718 42914 259954
rect 42294 259634 42914 259718
rect 42294 259398 42326 259634
rect 42562 259398 42646 259634
rect 42882 259398 42914 259634
rect 42294 223954 42914 259398
rect 42294 223718 42326 223954
rect 42562 223718 42646 223954
rect 42882 223718 42914 223954
rect 42294 223634 42914 223718
rect 42294 223398 42326 223634
rect 42562 223398 42646 223634
rect 42882 223398 42914 223634
rect 42294 187954 42914 223398
rect 42294 187718 42326 187954
rect 42562 187718 42646 187954
rect 42882 187718 42914 187954
rect 42294 187634 42914 187718
rect 42294 187398 42326 187634
rect 42562 187398 42646 187634
rect 42882 187398 42914 187634
rect 42294 151954 42914 187398
rect 42294 151718 42326 151954
rect 42562 151718 42646 151954
rect 42882 151718 42914 151954
rect 42294 151634 42914 151718
rect 42294 151398 42326 151634
rect 42562 151398 42646 151634
rect 42882 151398 42914 151634
rect 42294 115954 42914 151398
rect 42294 115718 42326 115954
rect 42562 115718 42646 115954
rect 42882 115718 42914 115954
rect 42294 115634 42914 115718
rect 42294 115398 42326 115634
rect 42562 115398 42646 115634
rect 42882 115398 42914 115634
rect 42294 79954 42914 115398
rect 42294 79718 42326 79954
rect 42562 79718 42646 79954
rect 42882 79718 42914 79954
rect 42294 79634 42914 79718
rect 42294 79398 42326 79634
rect 42562 79398 42646 79634
rect 42882 79398 42914 79634
rect 42294 43954 42914 79398
rect 42294 43718 42326 43954
rect 42562 43718 42646 43954
rect 42882 43718 42914 43954
rect 42294 43634 42914 43718
rect 42294 43398 42326 43634
rect 42562 43398 42646 43634
rect 42882 43398 42914 43634
rect 42294 7954 42914 43398
rect 42294 7718 42326 7954
rect 42562 7718 42646 7954
rect 42882 7718 42914 7954
rect 42294 7634 42914 7718
rect 42294 7398 42326 7634
rect 42562 7398 42646 7634
rect 42882 7398 42914 7634
rect 42294 -1306 42914 7398
rect 42294 -1542 42326 -1306
rect 42562 -1542 42646 -1306
rect 42882 -1542 42914 -1306
rect 42294 -1626 42914 -1542
rect 42294 -1862 42326 -1626
rect 42562 -1862 42646 -1626
rect 42882 -1862 42914 -1626
rect 42294 -7654 42914 -1862
rect 46794 706758 47414 711590
rect 46794 706522 46826 706758
rect 47062 706522 47146 706758
rect 47382 706522 47414 706758
rect 46794 706438 47414 706522
rect 46794 706202 46826 706438
rect 47062 706202 47146 706438
rect 47382 706202 47414 706438
rect 46794 696454 47414 706202
rect 46794 696218 46826 696454
rect 47062 696218 47146 696454
rect 47382 696218 47414 696454
rect 46794 696134 47414 696218
rect 46794 695898 46826 696134
rect 47062 695898 47146 696134
rect 47382 695898 47414 696134
rect 46794 660454 47414 695898
rect 46794 660218 46826 660454
rect 47062 660218 47146 660454
rect 47382 660218 47414 660454
rect 46794 660134 47414 660218
rect 46794 659898 46826 660134
rect 47062 659898 47146 660134
rect 47382 659898 47414 660134
rect 46794 624454 47414 659898
rect 46794 624218 46826 624454
rect 47062 624218 47146 624454
rect 47382 624218 47414 624454
rect 46794 624134 47414 624218
rect 46794 623898 46826 624134
rect 47062 623898 47146 624134
rect 47382 623898 47414 624134
rect 46794 588454 47414 623898
rect 46794 588218 46826 588454
rect 47062 588218 47146 588454
rect 47382 588218 47414 588454
rect 46794 588134 47414 588218
rect 46794 587898 46826 588134
rect 47062 587898 47146 588134
rect 47382 587898 47414 588134
rect 46794 552454 47414 587898
rect 46794 552218 46826 552454
rect 47062 552218 47146 552454
rect 47382 552218 47414 552454
rect 46794 552134 47414 552218
rect 46794 551898 46826 552134
rect 47062 551898 47146 552134
rect 47382 551898 47414 552134
rect 46794 516454 47414 551898
rect 46794 516218 46826 516454
rect 47062 516218 47146 516454
rect 47382 516218 47414 516454
rect 46794 516134 47414 516218
rect 46794 515898 46826 516134
rect 47062 515898 47146 516134
rect 47382 515898 47414 516134
rect 46794 480454 47414 515898
rect 46794 480218 46826 480454
rect 47062 480218 47146 480454
rect 47382 480218 47414 480454
rect 46794 480134 47414 480218
rect 46794 479898 46826 480134
rect 47062 479898 47146 480134
rect 47382 479898 47414 480134
rect 46794 444454 47414 479898
rect 46794 444218 46826 444454
rect 47062 444218 47146 444454
rect 47382 444218 47414 444454
rect 46794 444134 47414 444218
rect 46794 443898 46826 444134
rect 47062 443898 47146 444134
rect 47382 443898 47414 444134
rect 46794 408454 47414 443898
rect 46794 408218 46826 408454
rect 47062 408218 47146 408454
rect 47382 408218 47414 408454
rect 46794 408134 47414 408218
rect 46794 407898 46826 408134
rect 47062 407898 47146 408134
rect 47382 407898 47414 408134
rect 46794 372454 47414 407898
rect 46794 372218 46826 372454
rect 47062 372218 47146 372454
rect 47382 372218 47414 372454
rect 46794 372134 47414 372218
rect 46794 371898 46826 372134
rect 47062 371898 47146 372134
rect 47382 371898 47414 372134
rect 46794 336454 47414 371898
rect 46794 336218 46826 336454
rect 47062 336218 47146 336454
rect 47382 336218 47414 336454
rect 46794 336134 47414 336218
rect 46794 335898 46826 336134
rect 47062 335898 47146 336134
rect 47382 335898 47414 336134
rect 46794 300454 47414 335898
rect 46794 300218 46826 300454
rect 47062 300218 47146 300454
rect 47382 300218 47414 300454
rect 46794 300134 47414 300218
rect 46794 299898 46826 300134
rect 47062 299898 47146 300134
rect 47382 299898 47414 300134
rect 46794 264454 47414 299898
rect 46794 264218 46826 264454
rect 47062 264218 47146 264454
rect 47382 264218 47414 264454
rect 46794 264134 47414 264218
rect 46794 263898 46826 264134
rect 47062 263898 47146 264134
rect 47382 263898 47414 264134
rect 46794 228454 47414 263898
rect 46794 228218 46826 228454
rect 47062 228218 47146 228454
rect 47382 228218 47414 228454
rect 46794 228134 47414 228218
rect 46794 227898 46826 228134
rect 47062 227898 47146 228134
rect 47382 227898 47414 228134
rect 46794 192454 47414 227898
rect 46794 192218 46826 192454
rect 47062 192218 47146 192454
rect 47382 192218 47414 192454
rect 46794 192134 47414 192218
rect 46794 191898 46826 192134
rect 47062 191898 47146 192134
rect 47382 191898 47414 192134
rect 46794 156454 47414 191898
rect 46794 156218 46826 156454
rect 47062 156218 47146 156454
rect 47382 156218 47414 156454
rect 46794 156134 47414 156218
rect 46794 155898 46826 156134
rect 47062 155898 47146 156134
rect 47382 155898 47414 156134
rect 46794 120454 47414 155898
rect 46794 120218 46826 120454
rect 47062 120218 47146 120454
rect 47382 120218 47414 120454
rect 46794 120134 47414 120218
rect 46794 119898 46826 120134
rect 47062 119898 47146 120134
rect 47382 119898 47414 120134
rect 46794 84454 47414 119898
rect 46794 84218 46826 84454
rect 47062 84218 47146 84454
rect 47382 84218 47414 84454
rect 46794 84134 47414 84218
rect 46794 83898 46826 84134
rect 47062 83898 47146 84134
rect 47382 83898 47414 84134
rect 46794 48454 47414 83898
rect 46794 48218 46826 48454
rect 47062 48218 47146 48454
rect 47382 48218 47414 48454
rect 46794 48134 47414 48218
rect 46794 47898 46826 48134
rect 47062 47898 47146 48134
rect 47382 47898 47414 48134
rect 46794 12454 47414 47898
rect 46794 12218 46826 12454
rect 47062 12218 47146 12454
rect 47382 12218 47414 12454
rect 46794 12134 47414 12218
rect 46794 11898 46826 12134
rect 47062 11898 47146 12134
rect 47382 11898 47414 12134
rect 46794 -2266 47414 11898
rect 46794 -2502 46826 -2266
rect 47062 -2502 47146 -2266
rect 47382 -2502 47414 -2266
rect 46794 -2586 47414 -2502
rect 46794 -2822 46826 -2586
rect 47062 -2822 47146 -2586
rect 47382 -2822 47414 -2586
rect 46794 -7654 47414 -2822
rect 51294 707718 51914 711590
rect 51294 707482 51326 707718
rect 51562 707482 51646 707718
rect 51882 707482 51914 707718
rect 51294 707398 51914 707482
rect 51294 707162 51326 707398
rect 51562 707162 51646 707398
rect 51882 707162 51914 707398
rect 51294 700954 51914 707162
rect 51294 700718 51326 700954
rect 51562 700718 51646 700954
rect 51882 700718 51914 700954
rect 51294 700634 51914 700718
rect 51294 700398 51326 700634
rect 51562 700398 51646 700634
rect 51882 700398 51914 700634
rect 51294 664954 51914 700398
rect 51294 664718 51326 664954
rect 51562 664718 51646 664954
rect 51882 664718 51914 664954
rect 51294 664634 51914 664718
rect 51294 664398 51326 664634
rect 51562 664398 51646 664634
rect 51882 664398 51914 664634
rect 51294 628954 51914 664398
rect 51294 628718 51326 628954
rect 51562 628718 51646 628954
rect 51882 628718 51914 628954
rect 51294 628634 51914 628718
rect 51294 628398 51326 628634
rect 51562 628398 51646 628634
rect 51882 628398 51914 628634
rect 51294 592954 51914 628398
rect 51294 592718 51326 592954
rect 51562 592718 51646 592954
rect 51882 592718 51914 592954
rect 51294 592634 51914 592718
rect 51294 592398 51326 592634
rect 51562 592398 51646 592634
rect 51882 592398 51914 592634
rect 51294 556954 51914 592398
rect 51294 556718 51326 556954
rect 51562 556718 51646 556954
rect 51882 556718 51914 556954
rect 51294 556634 51914 556718
rect 51294 556398 51326 556634
rect 51562 556398 51646 556634
rect 51882 556398 51914 556634
rect 51294 520954 51914 556398
rect 51294 520718 51326 520954
rect 51562 520718 51646 520954
rect 51882 520718 51914 520954
rect 51294 520634 51914 520718
rect 51294 520398 51326 520634
rect 51562 520398 51646 520634
rect 51882 520398 51914 520634
rect 51294 484954 51914 520398
rect 51294 484718 51326 484954
rect 51562 484718 51646 484954
rect 51882 484718 51914 484954
rect 51294 484634 51914 484718
rect 51294 484398 51326 484634
rect 51562 484398 51646 484634
rect 51882 484398 51914 484634
rect 51294 448954 51914 484398
rect 51294 448718 51326 448954
rect 51562 448718 51646 448954
rect 51882 448718 51914 448954
rect 51294 448634 51914 448718
rect 51294 448398 51326 448634
rect 51562 448398 51646 448634
rect 51882 448398 51914 448634
rect 51294 412954 51914 448398
rect 51294 412718 51326 412954
rect 51562 412718 51646 412954
rect 51882 412718 51914 412954
rect 51294 412634 51914 412718
rect 51294 412398 51326 412634
rect 51562 412398 51646 412634
rect 51882 412398 51914 412634
rect 51294 376954 51914 412398
rect 51294 376718 51326 376954
rect 51562 376718 51646 376954
rect 51882 376718 51914 376954
rect 51294 376634 51914 376718
rect 51294 376398 51326 376634
rect 51562 376398 51646 376634
rect 51882 376398 51914 376634
rect 51294 340954 51914 376398
rect 51294 340718 51326 340954
rect 51562 340718 51646 340954
rect 51882 340718 51914 340954
rect 51294 340634 51914 340718
rect 51294 340398 51326 340634
rect 51562 340398 51646 340634
rect 51882 340398 51914 340634
rect 51294 304954 51914 340398
rect 51294 304718 51326 304954
rect 51562 304718 51646 304954
rect 51882 304718 51914 304954
rect 51294 304634 51914 304718
rect 51294 304398 51326 304634
rect 51562 304398 51646 304634
rect 51882 304398 51914 304634
rect 51294 268954 51914 304398
rect 51294 268718 51326 268954
rect 51562 268718 51646 268954
rect 51882 268718 51914 268954
rect 51294 268634 51914 268718
rect 51294 268398 51326 268634
rect 51562 268398 51646 268634
rect 51882 268398 51914 268634
rect 51294 232954 51914 268398
rect 51294 232718 51326 232954
rect 51562 232718 51646 232954
rect 51882 232718 51914 232954
rect 51294 232634 51914 232718
rect 51294 232398 51326 232634
rect 51562 232398 51646 232634
rect 51882 232398 51914 232634
rect 51294 196954 51914 232398
rect 51294 196718 51326 196954
rect 51562 196718 51646 196954
rect 51882 196718 51914 196954
rect 51294 196634 51914 196718
rect 51294 196398 51326 196634
rect 51562 196398 51646 196634
rect 51882 196398 51914 196634
rect 51294 160954 51914 196398
rect 51294 160718 51326 160954
rect 51562 160718 51646 160954
rect 51882 160718 51914 160954
rect 51294 160634 51914 160718
rect 51294 160398 51326 160634
rect 51562 160398 51646 160634
rect 51882 160398 51914 160634
rect 51294 124954 51914 160398
rect 51294 124718 51326 124954
rect 51562 124718 51646 124954
rect 51882 124718 51914 124954
rect 51294 124634 51914 124718
rect 51294 124398 51326 124634
rect 51562 124398 51646 124634
rect 51882 124398 51914 124634
rect 51294 88954 51914 124398
rect 51294 88718 51326 88954
rect 51562 88718 51646 88954
rect 51882 88718 51914 88954
rect 51294 88634 51914 88718
rect 51294 88398 51326 88634
rect 51562 88398 51646 88634
rect 51882 88398 51914 88634
rect 51294 52954 51914 88398
rect 51294 52718 51326 52954
rect 51562 52718 51646 52954
rect 51882 52718 51914 52954
rect 51294 52634 51914 52718
rect 51294 52398 51326 52634
rect 51562 52398 51646 52634
rect 51882 52398 51914 52634
rect 51294 16954 51914 52398
rect 51294 16718 51326 16954
rect 51562 16718 51646 16954
rect 51882 16718 51914 16954
rect 51294 16634 51914 16718
rect 51294 16398 51326 16634
rect 51562 16398 51646 16634
rect 51882 16398 51914 16634
rect 51294 -3226 51914 16398
rect 51294 -3462 51326 -3226
rect 51562 -3462 51646 -3226
rect 51882 -3462 51914 -3226
rect 51294 -3546 51914 -3462
rect 51294 -3782 51326 -3546
rect 51562 -3782 51646 -3546
rect 51882 -3782 51914 -3546
rect 51294 -7654 51914 -3782
rect 55794 708678 56414 711590
rect 55794 708442 55826 708678
rect 56062 708442 56146 708678
rect 56382 708442 56414 708678
rect 55794 708358 56414 708442
rect 55794 708122 55826 708358
rect 56062 708122 56146 708358
rect 56382 708122 56414 708358
rect 55794 669454 56414 708122
rect 55794 669218 55826 669454
rect 56062 669218 56146 669454
rect 56382 669218 56414 669454
rect 55794 669134 56414 669218
rect 55794 668898 55826 669134
rect 56062 668898 56146 669134
rect 56382 668898 56414 669134
rect 55794 633454 56414 668898
rect 55794 633218 55826 633454
rect 56062 633218 56146 633454
rect 56382 633218 56414 633454
rect 55794 633134 56414 633218
rect 55794 632898 55826 633134
rect 56062 632898 56146 633134
rect 56382 632898 56414 633134
rect 55794 597454 56414 632898
rect 55794 597218 55826 597454
rect 56062 597218 56146 597454
rect 56382 597218 56414 597454
rect 55794 597134 56414 597218
rect 55794 596898 55826 597134
rect 56062 596898 56146 597134
rect 56382 596898 56414 597134
rect 55794 561454 56414 596898
rect 55794 561218 55826 561454
rect 56062 561218 56146 561454
rect 56382 561218 56414 561454
rect 55794 561134 56414 561218
rect 55794 560898 55826 561134
rect 56062 560898 56146 561134
rect 56382 560898 56414 561134
rect 55794 525454 56414 560898
rect 55794 525218 55826 525454
rect 56062 525218 56146 525454
rect 56382 525218 56414 525454
rect 55794 525134 56414 525218
rect 55794 524898 55826 525134
rect 56062 524898 56146 525134
rect 56382 524898 56414 525134
rect 55794 489454 56414 524898
rect 55794 489218 55826 489454
rect 56062 489218 56146 489454
rect 56382 489218 56414 489454
rect 55794 489134 56414 489218
rect 55794 488898 55826 489134
rect 56062 488898 56146 489134
rect 56382 488898 56414 489134
rect 55794 453454 56414 488898
rect 55794 453218 55826 453454
rect 56062 453218 56146 453454
rect 56382 453218 56414 453454
rect 55794 453134 56414 453218
rect 55794 452898 55826 453134
rect 56062 452898 56146 453134
rect 56382 452898 56414 453134
rect 55794 417454 56414 452898
rect 55794 417218 55826 417454
rect 56062 417218 56146 417454
rect 56382 417218 56414 417454
rect 55794 417134 56414 417218
rect 55794 416898 55826 417134
rect 56062 416898 56146 417134
rect 56382 416898 56414 417134
rect 55794 381454 56414 416898
rect 55794 381218 55826 381454
rect 56062 381218 56146 381454
rect 56382 381218 56414 381454
rect 55794 381134 56414 381218
rect 55794 380898 55826 381134
rect 56062 380898 56146 381134
rect 56382 380898 56414 381134
rect 55794 345454 56414 380898
rect 55794 345218 55826 345454
rect 56062 345218 56146 345454
rect 56382 345218 56414 345454
rect 55794 345134 56414 345218
rect 55794 344898 55826 345134
rect 56062 344898 56146 345134
rect 56382 344898 56414 345134
rect 55794 309454 56414 344898
rect 55794 309218 55826 309454
rect 56062 309218 56146 309454
rect 56382 309218 56414 309454
rect 55794 309134 56414 309218
rect 55794 308898 55826 309134
rect 56062 308898 56146 309134
rect 56382 308898 56414 309134
rect 55794 273454 56414 308898
rect 55794 273218 55826 273454
rect 56062 273218 56146 273454
rect 56382 273218 56414 273454
rect 55794 273134 56414 273218
rect 55794 272898 55826 273134
rect 56062 272898 56146 273134
rect 56382 272898 56414 273134
rect 55794 237454 56414 272898
rect 55794 237218 55826 237454
rect 56062 237218 56146 237454
rect 56382 237218 56414 237454
rect 55794 237134 56414 237218
rect 55794 236898 55826 237134
rect 56062 236898 56146 237134
rect 56382 236898 56414 237134
rect 55794 201454 56414 236898
rect 55794 201218 55826 201454
rect 56062 201218 56146 201454
rect 56382 201218 56414 201454
rect 55794 201134 56414 201218
rect 55794 200898 55826 201134
rect 56062 200898 56146 201134
rect 56382 200898 56414 201134
rect 55794 165454 56414 200898
rect 55794 165218 55826 165454
rect 56062 165218 56146 165454
rect 56382 165218 56414 165454
rect 55794 165134 56414 165218
rect 55794 164898 55826 165134
rect 56062 164898 56146 165134
rect 56382 164898 56414 165134
rect 55794 129454 56414 164898
rect 55794 129218 55826 129454
rect 56062 129218 56146 129454
rect 56382 129218 56414 129454
rect 55794 129134 56414 129218
rect 55794 128898 55826 129134
rect 56062 128898 56146 129134
rect 56382 128898 56414 129134
rect 55794 93454 56414 128898
rect 55794 93218 55826 93454
rect 56062 93218 56146 93454
rect 56382 93218 56414 93454
rect 55794 93134 56414 93218
rect 55794 92898 55826 93134
rect 56062 92898 56146 93134
rect 56382 92898 56414 93134
rect 55794 57454 56414 92898
rect 55794 57218 55826 57454
rect 56062 57218 56146 57454
rect 56382 57218 56414 57454
rect 55794 57134 56414 57218
rect 55794 56898 55826 57134
rect 56062 56898 56146 57134
rect 56382 56898 56414 57134
rect 55794 21454 56414 56898
rect 55794 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 56414 21454
rect 55794 21134 56414 21218
rect 55794 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 56414 21134
rect 55794 -4186 56414 20898
rect 55794 -4422 55826 -4186
rect 56062 -4422 56146 -4186
rect 56382 -4422 56414 -4186
rect 55794 -4506 56414 -4422
rect 55794 -4742 55826 -4506
rect 56062 -4742 56146 -4506
rect 56382 -4742 56414 -4506
rect 55794 -7654 56414 -4742
rect 60294 709638 60914 711590
rect 60294 709402 60326 709638
rect 60562 709402 60646 709638
rect 60882 709402 60914 709638
rect 60294 709318 60914 709402
rect 60294 709082 60326 709318
rect 60562 709082 60646 709318
rect 60882 709082 60914 709318
rect 60294 673954 60914 709082
rect 60294 673718 60326 673954
rect 60562 673718 60646 673954
rect 60882 673718 60914 673954
rect 60294 673634 60914 673718
rect 60294 673398 60326 673634
rect 60562 673398 60646 673634
rect 60882 673398 60914 673634
rect 60294 637954 60914 673398
rect 60294 637718 60326 637954
rect 60562 637718 60646 637954
rect 60882 637718 60914 637954
rect 60294 637634 60914 637718
rect 60294 637398 60326 637634
rect 60562 637398 60646 637634
rect 60882 637398 60914 637634
rect 60294 601954 60914 637398
rect 60294 601718 60326 601954
rect 60562 601718 60646 601954
rect 60882 601718 60914 601954
rect 60294 601634 60914 601718
rect 60294 601398 60326 601634
rect 60562 601398 60646 601634
rect 60882 601398 60914 601634
rect 60294 565954 60914 601398
rect 60294 565718 60326 565954
rect 60562 565718 60646 565954
rect 60882 565718 60914 565954
rect 60294 565634 60914 565718
rect 60294 565398 60326 565634
rect 60562 565398 60646 565634
rect 60882 565398 60914 565634
rect 60294 529954 60914 565398
rect 60294 529718 60326 529954
rect 60562 529718 60646 529954
rect 60882 529718 60914 529954
rect 60294 529634 60914 529718
rect 60294 529398 60326 529634
rect 60562 529398 60646 529634
rect 60882 529398 60914 529634
rect 60294 493954 60914 529398
rect 60294 493718 60326 493954
rect 60562 493718 60646 493954
rect 60882 493718 60914 493954
rect 60294 493634 60914 493718
rect 60294 493398 60326 493634
rect 60562 493398 60646 493634
rect 60882 493398 60914 493634
rect 60294 457954 60914 493398
rect 60294 457718 60326 457954
rect 60562 457718 60646 457954
rect 60882 457718 60914 457954
rect 60294 457634 60914 457718
rect 60294 457398 60326 457634
rect 60562 457398 60646 457634
rect 60882 457398 60914 457634
rect 60294 421954 60914 457398
rect 60294 421718 60326 421954
rect 60562 421718 60646 421954
rect 60882 421718 60914 421954
rect 60294 421634 60914 421718
rect 60294 421398 60326 421634
rect 60562 421398 60646 421634
rect 60882 421398 60914 421634
rect 60294 385954 60914 421398
rect 60294 385718 60326 385954
rect 60562 385718 60646 385954
rect 60882 385718 60914 385954
rect 60294 385634 60914 385718
rect 60294 385398 60326 385634
rect 60562 385398 60646 385634
rect 60882 385398 60914 385634
rect 60294 349954 60914 385398
rect 60294 349718 60326 349954
rect 60562 349718 60646 349954
rect 60882 349718 60914 349954
rect 60294 349634 60914 349718
rect 60294 349398 60326 349634
rect 60562 349398 60646 349634
rect 60882 349398 60914 349634
rect 60294 313954 60914 349398
rect 60294 313718 60326 313954
rect 60562 313718 60646 313954
rect 60882 313718 60914 313954
rect 60294 313634 60914 313718
rect 60294 313398 60326 313634
rect 60562 313398 60646 313634
rect 60882 313398 60914 313634
rect 60294 277954 60914 313398
rect 60294 277718 60326 277954
rect 60562 277718 60646 277954
rect 60882 277718 60914 277954
rect 60294 277634 60914 277718
rect 60294 277398 60326 277634
rect 60562 277398 60646 277634
rect 60882 277398 60914 277634
rect 60294 241954 60914 277398
rect 60294 241718 60326 241954
rect 60562 241718 60646 241954
rect 60882 241718 60914 241954
rect 60294 241634 60914 241718
rect 60294 241398 60326 241634
rect 60562 241398 60646 241634
rect 60882 241398 60914 241634
rect 60294 205954 60914 241398
rect 60294 205718 60326 205954
rect 60562 205718 60646 205954
rect 60882 205718 60914 205954
rect 60294 205634 60914 205718
rect 60294 205398 60326 205634
rect 60562 205398 60646 205634
rect 60882 205398 60914 205634
rect 60294 169954 60914 205398
rect 60294 169718 60326 169954
rect 60562 169718 60646 169954
rect 60882 169718 60914 169954
rect 60294 169634 60914 169718
rect 60294 169398 60326 169634
rect 60562 169398 60646 169634
rect 60882 169398 60914 169634
rect 60294 133954 60914 169398
rect 60294 133718 60326 133954
rect 60562 133718 60646 133954
rect 60882 133718 60914 133954
rect 60294 133634 60914 133718
rect 60294 133398 60326 133634
rect 60562 133398 60646 133634
rect 60882 133398 60914 133634
rect 60294 97954 60914 133398
rect 60294 97718 60326 97954
rect 60562 97718 60646 97954
rect 60882 97718 60914 97954
rect 60294 97634 60914 97718
rect 60294 97398 60326 97634
rect 60562 97398 60646 97634
rect 60882 97398 60914 97634
rect 60294 61954 60914 97398
rect 60294 61718 60326 61954
rect 60562 61718 60646 61954
rect 60882 61718 60914 61954
rect 60294 61634 60914 61718
rect 60294 61398 60326 61634
rect 60562 61398 60646 61634
rect 60882 61398 60914 61634
rect 60294 25954 60914 61398
rect 60294 25718 60326 25954
rect 60562 25718 60646 25954
rect 60882 25718 60914 25954
rect 60294 25634 60914 25718
rect 60294 25398 60326 25634
rect 60562 25398 60646 25634
rect 60882 25398 60914 25634
rect 60294 -5146 60914 25398
rect 60294 -5382 60326 -5146
rect 60562 -5382 60646 -5146
rect 60882 -5382 60914 -5146
rect 60294 -5466 60914 -5382
rect 60294 -5702 60326 -5466
rect 60562 -5702 60646 -5466
rect 60882 -5702 60914 -5466
rect 60294 -7654 60914 -5702
rect 64794 710598 65414 711590
rect 64794 710362 64826 710598
rect 65062 710362 65146 710598
rect 65382 710362 65414 710598
rect 64794 710278 65414 710362
rect 64794 710042 64826 710278
rect 65062 710042 65146 710278
rect 65382 710042 65414 710278
rect 64794 678454 65414 710042
rect 64794 678218 64826 678454
rect 65062 678218 65146 678454
rect 65382 678218 65414 678454
rect 64794 678134 65414 678218
rect 64794 677898 64826 678134
rect 65062 677898 65146 678134
rect 65382 677898 65414 678134
rect 64794 642454 65414 677898
rect 64794 642218 64826 642454
rect 65062 642218 65146 642454
rect 65382 642218 65414 642454
rect 64794 642134 65414 642218
rect 64794 641898 64826 642134
rect 65062 641898 65146 642134
rect 65382 641898 65414 642134
rect 64794 606454 65414 641898
rect 64794 606218 64826 606454
rect 65062 606218 65146 606454
rect 65382 606218 65414 606454
rect 64794 606134 65414 606218
rect 64794 605898 64826 606134
rect 65062 605898 65146 606134
rect 65382 605898 65414 606134
rect 64794 570454 65414 605898
rect 64794 570218 64826 570454
rect 65062 570218 65146 570454
rect 65382 570218 65414 570454
rect 64794 570134 65414 570218
rect 64794 569898 64826 570134
rect 65062 569898 65146 570134
rect 65382 569898 65414 570134
rect 64794 534454 65414 569898
rect 64794 534218 64826 534454
rect 65062 534218 65146 534454
rect 65382 534218 65414 534454
rect 64794 534134 65414 534218
rect 64794 533898 64826 534134
rect 65062 533898 65146 534134
rect 65382 533898 65414 534134
rect 64794 498454 65414 533898
rect 64794 498218 64826 498454
rect 65062 498218 65146 498454
rect 65382 498218 65414 498454
rect 64794 498134 65414 498218
rect 64794 497898 64826 498134
rect 65062 497898 65146 498134
rect 65382 497898 65414 498134
rect 64794 462454 65414 497898
rect 64794 462218 64826 462454
rect 65062 462218 65146 462454
rect 65382 462218 65414 462454
rect 64794 462134 65414 462218
rect 64794 461898 64826 462134
rect 65062 461898 65146 462134
rect 65382 461898 65414 462134
rect 64794 426454 65414 461898
rect 64794 426218 64826 426454
rect 65062 426218 65146 426454
rect 65382 426218 65414 426454
rect 64794 426134 65414 426218
rect 64794 425898 64826 426134
rect 65062 425898 65146 426134
rect 65382 425898 65414 426134
rect 64794 390454 65414 425898
rect 64794 390218 64826 390454
rect 65062 390218 65146 390454
rect 65382 390218 65414 390454
rect 64794 390134 65414 390218
rect 64794 389898 64826 390134
rect 65062 389898 65146 390134
rect 65382 389898 65414 390134
rect 64794 354454 65414 389898
rect 64794 354218 64826 354454
rect 65062 354218 65146 354454
rect 65382 354218 65414 354454
rect 64794 354134 65414 354218
rect 64794 353898 64826 354134
rect 65062 353898 65146 354134
rect 65382 353898 65414 354134
rect 64794 318454 65414 353898
rect 64794 318218 64826 318454
rect 65062 318218 65146 318454
rect 65382 318218 65414 318454
rect 64794 318134 65414 318218
rect 64794 317898 64826 318134
rect 65062 317898 65146 318134
rect 65382 317898 65414 318134
rect 64794 282454 65414 317898
rect 64794 282218 64826 282454
rect 65062 282218 65146 282454
rect 65382 282218 65414 282454
rect 64794 282134 65414 282218
rect 64794 281898 64826 282134
rect 65062 281898 65146 282134
rect 65382 281898 65414 282134
rect 64794 246454 65414 281898
rect 64794 246218 64826 246454
rect 65062 246218 65146 246454
rect 65382 246218 65414 246454
rect 64794 246134 65414 246218
rect 64794 245898 64826 246134
rect 65062 245898 65146 246134
rect 65382 245898 65414 246134
rect 64794 210454 65414 245898
rect 64794 210218 64826 210454
rect 65062 210218 65146 210454
rect 65382 210218 65414 210454
rect 64794 210134 65414 210218
rect 64794 209898 64826 210134
rect 65062 209898 65146 210134
rect 65382 209898 65414 210134
rect 64794 174454 65414 209898
rect 64794 174218 64826 174454
rect 65062 174218 65146 174454
rect 65382 174218 65414 174454
rect 64794 174134 65414 174218
rect 64794 173898 64826 174134
rect 65062 173898 65146 174134
rect 65382 173898 65414 174134
rect 64794 138454 65414 173898
rect 64794 138218 64826 138454
rect 65062 138218 65146 138454
rect 65382 138218 65414 138454
rect 64794 138134 65414 138218
rect 64794 137898 64826 138134
rect 65062 137898 65146 138134
rect 65382 137898 65414 138134
rect 64794 102454 65414 137898
rect 64794 102218 64826 102454
rect 65062 102218 65146 102454
rect 65382 102218 65414 102454
rect 64794 102134 65414 102218
rect 64794 101898 64826 102134
rect 65062 101898 65146 102134
rect 65382 101898 65414 102134
rect 64794 66454 65414 101898
rect 64794 66218 64826 66454
rect 65062 66218 65146 66454
rect 65382 66218 65414 66454
rect 64794 66134 65414 66218
rect 64794 65898 64826 66134
rect 65062 65898 65146 66134
rect 65382 65898 65414 66134
rect 64794 30454 65414 65898
rect 64794 30218 64826 30454
rect 65062 30218 65146 30454
rect 65382 30218 65414 30454
rect 64794 30134 65414 30218
rect 64794 29898 64826 30134
rect 65062 29898 65146 30134
rect 65382 29898 65414 30134
rect 64794 -6106 65414 29898
rect 64794 -6342 64826 -6106
rect 65062 -6342 65146 -6106
rect 65382 -6342 65414 -6106
rect 64794 -6426 65414 -6342
rect 64794 -6662 64826 -6426
rect 65062 -6662 65146 -6426
rect 65382 -6662 65414 -6426
rect 64794 -7654 65414 -6662
rect 69294 711558 69914 711590
rect 69294 711322 69326 711558
rect 69562 711322 69646 711558
rect 69882 711322 69914 711558
rect 69294 711238 69914 711322
rect 69294 711002 69326 711238
rect 69562 711002 69646 711238
rect 69882 711002 69914 711238
rect 69294 682954 69914 711002
rect 69294 682718 69326 682954
rect 69562 682718 69646 682954
rect 69882 682718 69914 682954
rect 69294 682634 69914 682718
rect 69294 682398 69326 682634
rect 69562 682398 69646 682634
rect 69882 682398 69914 682634
rect 69294 646954 69914 682398
rect 69294 646718 69326 646954
rect 69562 646718 69646 646954
rect 69882 646718 69914 646954
rect 69294 646634 69914 646718
rect 69294 646398 69326 646634
rect 69562 646398 69646 646634
rect 69882 646398 69914 646634
rect 69294 610954 69914 646398
rect 69294 610718 69326 610954
rect 69562 610718 69646 610954
rect 69882 610718 69914 610954
rect 69294 610634 69914 610718
rect 69294 610398 69326 610634
rect 69562 610398 69646 610634
rect 69882 610398 69914 610634
rect 69294 574954 69914 610398
rect 69294 574718 69326 574954
rect 69562 574718 69646 574954
rect 69882 574718 69914 574954
rect 69294 574634 69914 574718
rect 69294 574398 69326 574634
rect 69562 574398 69646 574634
rect 69882 574398 69914 574634
rect 69294 538954 69914 574398
rect 69294 538718 69326 538954
rect 69562 538718 69646 538954
rect 69882 538718 69914 538954
rect 69294 538634 69914 538718
rect 69294 538398 69326 538634
rect 69562 538398 69646 538634
rect 69882 538398 69914 538634
rect 69294 502954 69914 538398
rect 69294 502718 69326 502954
rect 69562 502718 69646 502954
rect 69882 502718 69914 502954
rect 69294 502634 69914 502718
rect 69294 502398 69326 502634
rect 69562 502398 69646 502634
rect 69882 502398 69914 502634
rect 69294 466954 69914 502398
rect 69294 466718 69326 466954
rect 69562 466718 69646 466954
rect 69882 466718 69914 466954
rect 69294 466634 69914 466718
rect 69294 466398 69326 466634
rect 69562 466398 69646 466634
rect 69882 466398 69914 466634
rect 69294 430954 69914 466398
rect 69294 430718 69326 430954
rect 69562 430718 69646 430954
rect 69882 430718 69914 430954
rect 69294 430634 69914 430718
rect 69294 430398 69326 430634
rect 69562 430398 69646 430634
rect 69882 430398 69914 430634
rect 69294 394954 69914 430398
rect 69294 394718 69326 394954
rect 69562 394718 69646 394954
rect 69882 394718 69914 394954
rect 69294 394634 69914 394718
rect 69294 394398 69326 394634
rect 69562 394398 69646 394634
rect 69882 394398 69914 394634
rect 69294 358954 69914 394398
rect 69294 358718 69326 358954
rect 69562 358718 69646 358954
rect 69882 358718 69914 358954
rect 69294 358634 69914 358718
rect 69294 358398 69326 358634
rect 69562 358398 69646 358634
rect 69882 358398 69914 358634
rect 69294 322954 69914 358398
rect 69294 322718 69326 322954
rect 69562 322718 69646 322954
rect 69882 322718 69914 322954
rect 69294 322634 69914 322718
rect 69294 322398 69326 322634
rect 69562 322398 69646 322634
rect 69882 322398 69914 322634
rect 69294 286954 69914 322398
rect 69294 286718 69326 286954
rect 69562 286718 69646 286954
rect 69882 286718 69914 286954
rect 69294 286634 69914 286718
rect 69294 286398 69326 286634
rect 69562 286398 69646 286634
rect 69882 286398 69914 286634
rect 69294 250954 69914 286398
rect 69294 250718 69326 250954
rect 69562 250718 69646 250954
rect 69882 250718 69914 250954
rect 69294 250634 69914 250718
rect 69294 250398 69326 250634
rect 69562 250398 69646 250634
rect 69882 250398 69914 250634
rect 69294 214954 69914 250398
rect 69294 214718 69326 214954
rect 69562 214718 69646 214954
rect 69882 214718 69914 214954
rect 69294 214634 69914 214718
rect 69294 214398 69326 214634
rect 69562 214398 69646 214634
rect 69882 214398 69914 214634
rect 69294 178954 69914 214398
rect 69294 178718 69326 178954
rect 69562 178718 69646 178954
rect 69882 178718 69914 178954
rect 69294 178634 69914 178718
rect 69294 178398 69326 178634
rect 69562 178398 69646 178634
rect 69882 178398 69914 178634
rect 69294 142954 69914 178398
rect 69294 142718 69326 142954
rect 69562 142718 69646 142954
rect 69882 142718 69914 142954
rect 69294 142634 69914 142718
rect 69294 142398 69326 142634
rect 69562 142398 69646 142634
rect 69882 142398 69914 142634
rect 69294 106954 69914 142398
rect 69294 106718 69326 106954
rect 69562 106718 69646 106954
rect 69882 106718 69914 106954
rect 69294 106634 69914 106718
rect 69294 106398 69326 106634
rect 69562 106398 69646 106634
rect 69882 106398 69914 106634
rect 69294 70954 69914 106398
rect 69294 70718 69326 70954
rect 69562 70718 69646 70954
rect 69882 70718 69914 70954
rect 69294 70634 69914 70718
rect 69294 70398 69326 70634
rect 69562 70398 69646 70634
rect 69882 70398 69914 70634
rect 69294 34954 69914 70398
rect 69294 34718 69326 34954
rect 69562 34718 69646 34954
rect 69882 34718 69914 34954
rect 69294 34634 69914 34718
rect 69294 34398 69326 34634
rect 69562 34398 69646 34634
rect 69882 34398 69914 34634
rect 69294 -7066 69914 34398
rect 69294 -7302 69326 -7066
rect 69562 -7302 69646 -7066
rect 69882 -7302 69914 -7066
rect 69294 -7386 69914 -7302
rect 69294 -7622 69326 -7386
rect 69562 -7622 69646 -7386
rect 69882 -7622 69914 -7386
rect 69294 -7654 69914 -7622
rect 73794 704838 74414 711590
rect 73794 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 74414 704838
rect 73794 704518 74414 704602
rect 73794 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 74414 704518
rect 73794 687454 74414 704282
rect 73794 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 74414 687454
rect 73794 687134 74414 687218
rect 73794 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 74414 687134
rect 73794 651454 74414 686898
rect 73794 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 74414 651454
rect 73794 651134 74414 651218
rect 73794 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 74414 651134
rect 73794 615454 74414 650898
rect 73794 615218 73826 615454
rect 74062 615218 74146 615454
rect 74382 615218 74414 615454
rect 73794 615134 74414 615218
rect 73794 614898 73826 615134
rect 74062 614898 74146 615134
rect 74382 614898 74414 615134
rect 73794 579454 74414 614898
rect 73794 579218 73826 579454
rect 74062 579218 74146 579454
rect 74382 579218 74414 579454
rect 73794 579134 74414 579218
rect 73794 578898 73826 579134
rect 74062 578898 74146 579134
rect 74382 578898 74414 579134
rect 73794 543454 74414 578898
rect 73794 543218 73826 543454
rect 74062 543218 74146 543454
rect 74382 543218 74414 543454
rect 73794 543134 74414 543218
rect 73794 542898 73826 543134
rect 74062 542898 74146 543134
rect 74382 542898 74414 543134
rect 73794 507454 74414 542898
rect 73794 507218 73826 507454
rect 74062 507218 74146 507454
rect 74382 507218 74414 507454
rect 73794 507134 74414 507218
rect 73794 506898 73826 507134
rect 74062 506898 74146 507134
rect 74382 506898 74414 507134
rect 73794 471454 74414 506898
rect 73794 471218 73826 471454
rect 74062 471218 74146 471454
rect 74382 471218 74414 471454
rect 73794 471134 74414 471218
rect 73794 470898 73826 471134
rect 74062 470898 74146 471134
rect 74382 470898 74414 471134
rect 73794 435454 74414 470898
rect 73794 435218 73826 435454
rect 74062 435218 74146 435454
rect 74382 435218 74414 435454
rect 73794 435134 74414 435218
rect 73794 434898 73826 435134
rect 74062 434898 74146 435134
rect 74382 434898 74414 435134
rect 73794 399454 74414 434898
rect 73794 399218 73826 399454
rect 74062 399218 74146 399454
rect 74382 399218 74414 399454
rect 73794 399134 74414 399218
rect 73794 398898 73826 399134
rect 74062 398898 74146 399134
rect 74382 398898 74414 399134
rect 73794 363454 74414 398898
rect 73794 363218 73826 363454
rect 74062 363218 74146 363454
rect 74382 363218 74414 363454
rect 73794 363134 74414 363218
rect 73794 362898 73826 363134
rect 74062 362898 74146 363134
rect 74382 362898 74414 363134
rect 73794 327454 74414 362898
rect 73794 327218 73826 327454
rect 74062 327218 74146 327454
rect 74382 327218 74414 327454
rect 73794 327134 74414 327218
rect 73794 326898 73826 327134
rect 74062 326898 74146 327134
rect 74382 326898 74414 327134
rect 73794 291454 74414 326898
rect 73794 291218 73826 291454
rect 74062 291218 74146 291454
rect 74382 291218 74414 291454
rect 73794 291134 74414 291218
rect 73794 290898 73826 291134
rect 74062 290898 74146 291134
rect 74382 290898 74414 291134
rect 73794 255454 74414 290898
rect 73794 255218 73826 255454
rect 74062 255218 74146 255454
rect 74382 255218 74414 255454
rect 73794 255134 74414 255218
rect 73794 254898 73826 255134
rect 74062 254898 74146 255134
rect 74382 254898 74414 255134
rect 73794 219454 74414 254898
rect 73794 219218 73826 219454
rect 74062 219218 74146 219454
rect 74382 219218 74414 219454
rect 73794 219134 74414 219218
rect 73794 218898 73826 219134
rect 74062 218898 74146 219134
rect 74382 218898 74414 219134
rect 73794 183454 74414 218898
rect 73794 183218 73826 183454
rect 74062 183218 74146 183454
rect 74382 183218 74414 183454
rect 73794 183134 74414 183218
rect 73794 182898 73826 183134
rect 74062 182898 74146 183134
rect 74382 182898 74414 183134
rect 73794 147454 74414 182898
rect 73794 147218 73826 147454
rect 74062 147218 74146 147454
rect 74382 147218 74414 147454
rect 73794 147134 74414 147218
rect 73794 146898 73826 147134
rect 74062 146898 74146 147134
rect 74382 146898 74414 147134
rect 73794 111454 74414 146898
rect 73794 111218 73826 111454
rect 74062 111218 74146 111454
rect 74382 111218 74414 111454
rect 73794 111134 74414 111218
rect 73794 110898 73826 111134
rect 74062 110898 74146 111134
rect 74382 110898 74414 111134
rect 73794 75454 74414 110898
rect 73794 75218 73826 75454
rect 74062 75218 74146 75454
rect 74382 75218 74414 75454
rect 73794 75134 74414 75218
rect 73794 74898 73826 75134
rect 74062 74898 74146 75134
rect 74382 74898 74414 75134
rect 73794 39454 74414 74898
rect 73794 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 74414 39454
rect 73794 39134 74414 39218
rect 73794 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 74414 39134
rect 73794 3454 74414 38898
rect 73794 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 74414 3454
rect 73794 3134 74414 3218
rect 73794 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 74414 3134
rect 73794 -346 74414 2898
rect 73794 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 74414 -346
rect 73794 -666 74414 -582
rect 73794 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 74414 -666
rect 73794 -7654 74414 -902
rect 78294 705798 78914 711590
rect 78294 705562 78326 705798
rect 78562 705562 78646 705798
rect 78882 705562 78914 705798
rect 78294 705478 78914 705562
rect 78294 705242 78326 705478
rect 78562 705242 78646 705478
rect 78882 705242 78914 705478
rect 78294 691954 78914 705242
rect 78294 691718 78326 691954
rect 78562 691718 78646 691954
rect 78882 691718 78914 691954
rect 78294 691634 78914 691718
rect 78294 691398 78326 691634
rect 78562 691398 78646 691634
rect 78882 691398 78914 691634
rect 78294 655954 78914 691398
rect 78294 655718 78326 655954
rect 78562 655718 78646 655954
rect 78882 655718 78914 655954
rect 78294 655634 78914 655718
rect 78294 655398 78326 655634
rect 78562 655398 78646 655634
rect 78882 655398 78914 655634
rect 78294 619954 78914 655398
rect 78294 619718 78326 619954
rect 78562 619718 78646 619954
rect 78882 619718 78914 619954
rect 78294 619634 78914 619718
rect 78294 619398 78326 619634
rect 78562 619398 78646 619634
rect 78882 619398 78914 619634
rect 78294 583954 78914 619398
rect 78294 583718 78326 583954
rect 78562 583718 78646 583954
rect 78882 583718 78914 583954
rect 78294 583634 78914 583718
rect 78294 583398 78326 583634
rect 78562 583398 78646 583634
rect 78882 583398 78914 583634
rect 78294 547954 78914 583398
rect 78294 547718 78326 547954
rect 78562 547718 78646 547954
rect 78882 547718 78914 547954
rect 78294 547634 78914 547718
rect 78294 547398 78326 547634
rect 78562 547398 78646 547634
rect 78882 547398 78914 547634
rect 78294 511954 78914 547398
rect 78294 511718 78326 511954
rect 78562 511718 78646 511954
rect 78882 511718 78914 511954
rect 78294 511634 78914 511718
rect 78294 511398 78326 511634
rect 78562 511398 78646 511634
rect 78882 511398 78914 511634
rect 78294 475954 78914 511398
rect 78294 475718 78326 475954
rect 78562 475718 78646 475954
rect 78882 475718 78914 475954
rect 78294 475634 78914 475718
rect 78294 475398 78326 475634
rect 78562 475398 78646 475634
rect 78882 475398 78914 475634
rect 78294 439954 78914 475398
rect 78294 439718 78326 439954
rect 78562 439718 78646 439954
rect 78882 439718 78914 439954
rect 78294 439634 78914 439718
rect 78294 439398 78326 439634
rect 78562 439398 78646 439634
rect 78882 439398 78914 439634
rect 78294 403954 78914 439398
rect 78294 403718 78326 403954
rect 78562 403718 78646 403954
rect 78882 403718 78914 403954
rect 78294 403634 78914 403718
rect 78294 403398 78326 403634
rect 78562 403398 78646 403634
rect 78882 403398 78914 403634
rect 78294 367954 78914 403398
rect 78294 367718 78326 367954
rect 78562 367718 78646 367954
rect 78882 367718 78914 367954
rect 78294 367634 78914 367718
rect 78294 367398 78326 367634
rect 78562 367398 78646 367634
rect 78882 367398 78914 367634
rect 78294 331954 78914 367398
rect 78294 331718 78326 331954
rect 78562 331718 78646 331954
rect 78882 331718 78914 331954
rect 78294 331634 78914 331718
rect 78294 331398 78326 331634
rect 78562 331398 78646 331634
rect 78882 331398 78914 331634
rect 78294 295954 78914 331398
rect 78294 295718 78326 295954
rect 78562 295718 78646 295954
rect 78882 295718 78914 295954
rect 78294 295634 78914 295718
rect 78294 295398 78326 295634
rect 78562 295398 78646 295634
rect 78882 295398 78914 295634
rect 78294 259954 78914 295398
rect 78294 259718 78326 259954
rect 78562 259718 78646 259954
rect 78882 259718 78914 259954
rect 78294 259634 78914 259718
rect 78294 259398 78326 259634
rect 78562 259398 78646 259634
rect 78882 259398 78914 259634
rect 78294 223954 78914 259398
rect 78294 223718 78326 223954
rect 78562 223718 78646 223954
rect 78882 223718 78914 223954
rect 78294 223634 78914 223718
rect 78294 223398 78326 223634
rect 78562 223398 78646 223634
rect 78882 223398 78914 223634
rect 78294 187954 78914 223398
rect 78294 187718 78326 187954
rect 78562 187718 78646 187954
rect 78882 187718 78914 187954
rect 78294 187634 78914 187718
rect 78294 187398 78326 187634
rect 78562 187398 78646 187634
rect 78882 187398 78914 187634
rect 78294 151954 78914 187398
rect 78294 151718 78326 151954
rect 78562 151718 78646 151954
rect 78882 151718 78914 151954
rect 78294 151634 78914 151718
rect 78294 151398 78326 151634
rect 78562 151398 78646 151634
rect 78882 151398 78914 151634
rect 78294 115954 78914 151398
rect 78294 115718 78326 115954
rect 78562 115718 78646 115954
rect 78882 115718 78914 115954
rect 78294 115634 78914 115718
rect 78294 115398 78326 115634
rect 78562 115398 78646 115634
rect 78882 115398 78914 115634
rect 78294 79954 78914 115398
rect 78294 79718 78326 79954
rect 78562 79718 78646 79954
rect 78882 79718 78914 79954
rect 78294 79634 78914 79718
rect 78294 79398 78326 79634
rect 78562 79398 78646 79634
rect 78882 79398 78914 79634
rect 78294 43954 78914 79398
rect 78294 43718 78326 43954
rect 78562 43718 78646 43954
rect 78882 43718 78914 43954
rect 78294 43634 78914 43718
rect 78294 43398 78326 43634
rect 78562 43398 78646 43634
rect 78882 43398 78914 43634
rect 78294 7954 78914 43398
rect 78294 7718 78326 7954
rect 78562 7718 78646 7954
rect 78882 7718 78914 7954
rect 78294 7634 78914 7718
rect 78294 7398 78326 7634
rect 78562 7398 78646 7634
rect 78882 7398 78914 7634
rect 78294 -1306 78914 7398
rect 78294 -1542 78326 -1306
rect 78562 -1542 78646 -1306
rect 78882 -1542 78914 -1306
rect 78294 -1626 78914 -1542
rect 78294 -1862 78326 -1626
rect 78562 -1862 78646 -1626
rect 78882 -1862 78914 -1626
rect 78294 -7654 78914 -1862
rect 82794 706758 83414 711590
rect 82794 706522 82826 706758
rect 83062 706522 83146 706758
rect 83382 706522 83414 706758
rect 82794 706438 83414 706522
rect 82794 706202 82826 706438
rect 83062 706202 83146 706438
rect 83382 706202 83414 706438
rect 82794 696454 83414 706202
rect 82794 696218 82826 696454
rect 83062 696218 83146 696454
rect 83382 696218 83414 696454
rect 82794 696134 83414 696218
rect 82794 695898 82826 696134
rect 83062 695898 83146 696134
rect 83382 695898 83414 696134
rect 82794 660454 83414 695898
rect 82794 660218 82826 660454
rect 83062 660218 83146 660454
rect 83382 660218 83414 660454
rect 82794 660134 83414 660218
rect 82794 659898 82826 660134
rect 83062 659898 83146 660134
rect 83382 659898 83414 660134
rect 82794 624454 83414 659898
rect 82794 624218 82826 624454
rect 83062 624218 83146 624454
rect 83382 624218 83414 624454
rect 82794 624134 83414 624218
rect 82794 623898 82826 624134
rect 83062 623898 83146 624134
rect 83382 623898 83414 624134
rect 82794 588454 83414 623898
rect 82794 588218 82826 588454
rect 83062 588218 83146 588454
rect 83382 588218 83414 588454
rect 82794 588134 83414 588218
rect 82794 587898 82826 588134
rect 83062 587898 83146 588134
rect 83382 587898 83414 588134
rect 82794 552454 83414 587898
rect 82794 552218 82826 552454
rect 83062 552218 83146 552454
rect 83382 552218 83414 552454
rect 82794 552134 83414 552218
rect 82794 551898 82826 552134
rect 83062 551898 83146 552134
rect 83382 551898 83414 552134
rect 82794 516454 83414 551898
rect 82794 516218 82826 516454
rect 83062 516218 83146 516454
rect 83382 516218 83414 516454
rect 82794 516134 83414 516218
rect 82794 515898 82826 516134
rect 83062 515898 83146 516134
rect 83382 515898 83414 516134
rect 82794 480454 83414 515898
rect 82794 480218 82826 480454
rect 83062 480218 83146 480454
rect 83382 480218 83414 480454
rect 82794 480134 83414 480218
rect 82794 479898 82826 480134
rect 83062 479898 83146 480134
rect 83382 479898 83414 480134
rect 82794 444454 83414 479898
rect 82794 444218 82826 444454
rect 83062 444218 83146 444454
rect 83382 444218 83414 444454
rect 82794 444134 83414 444218
rect 82794 443898 82826 444134
rect 83062 443898 83146 444134
rect 83382 443898 83414 444134
rect 82794 408454 83414 443898
rect 82794 408218 82826 408454
rect 83062 408218 83146 408454
rect 83382 408218 83414 408454
rect 82794 408134 83414 408218
rect 82794 407898 82826 408134
rect 83062 407898 83146 408134
rect 83382 407898 83414 408134
rect 82794 372454 83414 407898
rect 82794 372218 82826 372454
rect 83062 372218 83146 372454
rect 83382 372218 83414 372454
rect 82794 372134 83414 372218
rect 82794 371898 82826 372134
rect 83062 371898 83146 372134
rect 83382 371898 83414 372134
rect 82794 336454 83414 371898
rect 82794 336218 82826 336454
rect 83062 336218 83146 336454
rect 83382 336218 83414 336454
rect 82794 336134 83414 336218
rect 82794 335898 82826 336134
rect 83062 335898 83146 336134
rect 83382 335898 83414 336134
rect 82794 300454 83414 335898
rect 82794 300218 82826 300454
rect 83062 300218 83146 300454
rect 83382 300218 83414 300454
rect 82794 300134 83414 300218
rect 82794 299898 82826 300134
rect 83062 299898 83146 300134
rect 83382 299898 83414 300134
rect 82794 264454 83414 299898
rect 82794 264218 82826 264454
rect 83062 264218 83146 264454
rect 83382 264218 83414 264454
rect 82794 264134 83414 264218
rect 82794 263898 82826 264134
rect 83062 263898 83146 264134
rect 83382 263898 83414 264134
rect 82794 228454 83414 263898
rect 82794 228218 82826 228454
rect 83062 228218 83146 228454
rect 83382 228218 83414 228454
rect 82794 228134 83414 228218
rect 82794 227898 82826 228134
rect 83062 227898 83146 228134
rect 83382 227898 83414 228134
rect 82794 192454 83414 227898
rect 82794 192218 82826 192454
rect 83062 192218 83146 192454
rect 83382 192218 83414 192454
rect 82794 192134 83414 192218
rect 82794 191898 82826 192134
rect 83062 191898 83146 192134
rect 83382 191898 83414 192134
rect 82794 156454 83414 191898
rect 82794 156218 82826 156454
rect 83062 156218 83146 156454
rect 83382 156218 83414 156454
rect 82794 156134 83414 156218
rect 82794 155898 82826 156134
rect 83062 155898 83146 156134
rect 83382 155898 83414 156134
rect 82794 120454 83414 155898
rect 82794 120218 82826 120454
rect 83062 120218 83146 120454
rect 83382 120218 83414 120454
rect 82794 120134 83414 120218
rect 82794 119898 82826 120134
rect 83062 119898 83146 120134
rect 83382 119898 83414 120134
rect 82794 84454 83414 119898
rect 82794 84218 82826 84454
rect 83062 84218 83146 84454
rect 83382 84218 83414 84454
rect 82794 84134 83414 84218
rect 82794 83898 82826 84134
rect 83062 83898 83146 84134
rect 83382 83898 83414 84134
rect 82794 48454 83414 83898
rect 82794 48218 82826 48454
rect 83062 48218 83146 48454
rect 83382 48218 83414 48454
rect 82794 48134 83414 48218
rect 82794 47898 82826 48134
rect 83062 47898 83146 48134
rect 83382 47898 83414 48134
rect 82794 12454 83414 47898
rect 82794 12218 82826 12454
rect 83062 12218 83146 12454
rect 83382 12218 83414 12454
rect 82794 12134 83414 12218
rect 82794 11898 82826 12134
rect 83062 11898 83146 12134
rect 83382 11898 83414 12134
rect 82794 -2266 83414 11898
rect 82794 -2502 82826 -2266
rect 83062 -2502 83146 -2266
rect 83382 -2502 83414 -2266
rect 82794 -2586 83414 -2502
rect 82794 -2822 82826 -2586
rect 83062 -2822 83146 -2586
rect 83382 -2822 83414 -2586
rect 82794 -7654 83414 -2822
rect 87294 707718 87914 711590
rect 87294 707482 87326 707718
rect 87562 707482 87646 707718
rect 87882 707482 87914 707718
rect 87294 707398 87914 707482
rect 87294 707162 87326 707398
rect 87562 707162 87646 707398
rect 87882 707162 87914 707398
rect 87294 700954 87914 707162
rect 87294 700718 87326 700954
rect 87562 700718 87646 700954
rect 87882 700718 87914 700954
rect 87294 700634 87914 700718
rect 87294 700398 87326 700634
rect 87562 700398 87646 700634
rect 87882 700398 87914 700634
rect 87294 664954 87914 700398
rect 87294 664718 87326 664954
rect 87562 664718 87646 664954
rect 87882 664718 87914 664954
rect 87294 664634 87914 664718
rect 87294 664398 87326 664634
rect 87562 664398 87646 664634
rect 87882 664398 87914 664634
rect 87294 628954 87914 664398
rect 87294 628718 87326 628954
rect 87562 628718 87646 628954
rect 87882 628718 87914 628954
rect 87294 628634 87914 628718
rect 87294 628398 87326 628634
rect 87562 628398 87646 628634
rect 87882 628398 87914 628634
rect 87294 592954 87914 628398
rect 87294 592718 87326 592954
rect 87562 592718 87646 592954
rect 87882 592718 87914 592954
rect 87294 592634 87914 592718
rect 87294 592398 87326 592634
rect 87562 592398 87646 592634
rect 87882 592398 87914 592634
rect 87294 556954 87914 592398
rect 87294 556718 87326 556954
rect 87562 556718 87646 556954
rect 87882 556718 87914 556954
rect 87294 556634 87914 556718
rect 87294 556398 87326 556634
rect 87562 556398 87646 556634
rect 87882 556398 87914 556634
rect 87294 520954 87914 556398
rect 87294 520718 87326 520954
rect 87562 520718 87646 520954
rect 87882 520718 87914 520954
rect 87294 520634 87914 520718
rect 87294 520398 87326 520634
rect 87562 520398 87646 520634
rect 87882 520398 87914 520634
rect 87294 484954 87914 520398
rect 87294 484718 87326 484954
rect 87562 484718 87646 484954
rect 87882 484718 87914 484954
rect 87294 484634 87914 484718
rect 87294 484398 87326 484634
rect 87562 484398 87646 484634
rect 87882 484398 87914 484634
rect 87294 448954 87914 484398
rect 87294 448718 87326 448954
rect 87562 448718 87646 448954
rect 87882 448718 87914 448954
rect 87294 448634 87914 448718
rect 87294 448398 87326 448634
rect 87562 448398 87646 448634
rect 87882 448398 87914 448634
rect 87294 412954 87914 448398
rect 87294 412718 87326 412954
rect 87562 412718 87646 412954
rect 87882 412718 87914 412954
rect 87294 412634 87914 412718
rect 87294 412398 87326 412634
rect 87562 412398 87646 412634
rect 87882 412398 87914 412634
rect 87294 376954 87914 412398
rect 87294 376718 87326 376954
rect 87562 376718 87646 376954
rect 87882 376718 87914 376954
rect 87294 376634 87914 376718
rect 87294 376398 87326 376634
rect 87562 376398 87646 376634
rect 87882 376398 87914 376634
rect 87294 340954 87914 376398
rect 87294 340718 87326 340954
rect 87562 340718 87646 340954
rect 87882 340718 87914 340954
rect 87294 340634 87914 340718
rect 87294 340398 87326 340634
rect 87562 340398 87646 340634
rect 87882 340398 87914 340634
rect 87294 304954 87914 340398
rect 87294 304718 87326 304954
rect 87562 304718 87646 304954
rect 87882 304718 87914 304954
rect 87294 304634 87914 304718
rect 87294 304398 87326 304634
rect 87562 304398 87646 304634
rect 87882 304398 87914 304634
rect 87294 268954 87914 304398
rect 87294 268718 87326 268954
rect 87562 268718 87646 268954
rect 87882 268718 87914 268954
rect 87294 268634 87914 268718
rect 87294 268398 87326 268634
rect 87562 268398 87646 268634
rect 87882 268398 87914 268634
rect 87294 232954 87914 268398
rect 87294 232718 87326 232954
rect 87562 232718 87646 232954
rect 87882 232718 87914 232954
rect 87294 232634 87914 232718
rect 87294 232398 87326 232634
rect 87562 232398 87646 232634
rect 87882 232398 87914 232634
rect 87294 196954 87914 232398
rect 87294 196718 87326 196954
rect 87562 196718 87646 196954
rect 87882 196718 87914 196954
rect 87294 196634 87914 196718
rect 87294 196398 87326 196634
rect 87562 196398 87646 196634
rect 87882 196398 87914 196634
rect 87294 160954 87914 196398
rect 87294 160718 87326 160954
rect 87562 160718 87646 160954
rect 87882 160718 87914 160954
rect 87294 160634 87914 160718
rect 87294 160398 87326 160634
rect 87562 160398 87646 160634
rect 87882 160398 87914 160634
rect 87294 124954 87914 160398
rect 87294 124718 87326 124954
rect 87562 124718 87646 124954
rect 87882 124718 87914 124954
rect 87294 124634 87914 124718
rect 87294 124398 87326 124634
rect 87562 124398 87646 124634
rect 87882 124398 87914 124634
rect 87294 88954 87914 124398
rect 87294 88718 87326 88954
rect 87562 88718 87646 88954
rect 87882 88718 87914 88954
rect 87294 88634 87914 88718
rect 87294 88398 87326 88634
rect 87562 88398 87646 88634
rect 87882 88398 87914 88634
rect 87294 52954 87914 88398
rect 87294 52718 87326 52954
rect 87562 52718 87646 52954
rect 87882 52718 87914 52954
rect 87294 52634 87914 52718
rect 87294 52398 87326 52634
rect 87562 52398 87646 52634
rect 87882 52398 87914 52634
rect 87294 16954 87914 52398
rect 87294 16718 87326 16954
rect 87562 16718 87646 16954
rect 87882 16718 87914 16954
rect 87294 16634 87914 16718
rect 87294 16398 87326 16634
rect 87562 16398 87646 16634
rect 87882 16398 87914 16634
rect 87294 -3226 87914 16398
rect 87294 -3462 87326 -3226
rect 87562 -3462 87646 -3226
rect 87882 -3462 87914 -3226
rect 87294 -3546 87914 -3462
rect 87294 -3782 87326 -3546
rect 87562 -3782 87646 -3546
rect 87882 -3782 87914 -3546
rect 87294 -7654 87914 -3782
rect 91794 708678 92414 711590
rect 91794 708442 91826 708678
rect 92062 708442 92146 708678
rect 92382 708442 92414 708678
rect 91794 708358 92414 708442
rect 91794 708122 91826 708358
rect 92062 708122 92146 708358
rect 92382 708122 92414 708358
rect 91794 669454 92414 708122
rect 91794 669218 91826 669454
rect 92062 669218 92146 669454
rect 92382 669218 92414 669454
rect 91794 669134 92414 669218
rect 91794 668898 91826 669134
rect 92062 668898 92146 669134
rect 92382 668898 92414 669134
rect 91794 633454 92414 668898
rect 91794 633218 91826 633454
rect 92062 633218 92146 633454
rect 92382 633218 92414 633454
rect 91794 633134 92414 633218
rect 91794 632898 91826 633134
rect 92062 632898 92146 633134
rect 92382 632898 92414 633134
rect 91794 597454 92414 632898
rect 91794 597218 91826 597454
rect 92062 597218 92146 597454
rect 92382 597218 92414 597454
rect 91794 597134 92414 597218
rect 91794 596898 91826 597134
rect 92062 596898 92146 597134
rect 92382 596898 92414 597134
rect 91794 561454 92414 596898
rect 91794 561218 91826 561454
rect 92062 561218 92146 561454
rect 92382 561218 92414 561454
rect 91794 561134 92414 561218
rect 91794 560898 91826 561134
rect 92062 560898 92146 561134
rect 92382 560898 92414 561134
rect 91794 525454 92414 560898
rect 91794 525218 91826 525454
rect 92062 525218 92146 525454
rect 92382 525218 92414 525454
rect 91794 525134 92414 525218
rect 91794 524898 91826 525134
rect 92062 524898 92146 525134
rect 92382 524898 92414 525134
rect 91794 489454 92414 524898
rect 91794 489218 91826 489454
rect 92062 489218 92146 489454
rect 92382 489218 92414 489454
rect 91794 489134 92414 489218
rect 91794 488898 91826 489134
rect 92062 488898 92146 489134
rect 92382 488898 92414 489134
rect 91794 453454 92414 488898
rect 91794 453218 91826 453454
rect 92062 453218 92146 453454
rect 92382 453218 92414 453454
rect 91794 453134 92414 453218
rect 91794 452898 91826 453134
rect 92062 452898 92146 453134
rect 92382 452898 92414 453134
rect 91794 417454 92414 452898
rect 91794 417218 91826 417454
rect 92062 417218 92146 417454
rect 92382 417218 92414 417454
rect 91794 417134 92414 417218
rect 91794 416898 91826 417134
rect 92062 416898 92146 417134
rect 92382 416898 92414 417134
rect 91794 381454 92414 416898
rect 91794 381218 91826 381454
rect 92062 381218 92146 381454
rect 92382 381218 92414 381454
rect 91794 381134 92414 381218
rect 91794 380898 91826 381134
rect 92062 380898 92146 381134
rect 92382 380898 92414 381134
rect 91794 345454 92414 380898
rect 91794 345218 91826 345454
rect 92062 345218 92146 345454
rect 92382 345218 92414 345454
rect 91794 345134 92414 345218
rect 91794 344898 91826 345134
rect 92062 344898 92146 345134
rect 92382 344898 92414 345134
rect 91794 309454 92414 344898
rect 91794 309218 91826 309454
rect 92062 309218 92146 309454
rect 92382 309218 92414 309454
rect 91794 309134 92414 309218
rect 91794 308898 91826 309134
rect 92062 308898 92146 309134
rect 92382 308898 92414 309134
rect 91794 273454 92414 308898
rect 91794 273218 91826 273454
rect 92062 273218 92146 273454
rect 92382 273218 92414 273454
rect 91794 273134 92414 273218
rect 91794 272898 91826 273134
rect 92062 272898 92146 273134
rect 92382 272898 92414 273134
rect 91794 237454 92414 272898
rect 91794 237218 91826 237454
rect 92062 237218 92146 237454
rect 92382 237218 92414 237454
rect 91794 237134 92414 237218
rect 91794 236898 91826 237134
rect 92062 236898 92146 237134
rect 92382 236898 92414 237134
rect 91794 201454 92414 236898
rect 91794 201218 91826 201454
rect 92062 201218 92146 201454
rect 92382 201218 92414 201454
rect 91794 201134 92414 201218
rect 91794 200898 91826 201134
rect 92062 200898 92146 201134
rect 92382 200898 92414 201134
rect 91794 165454 92414 200898
rect 91794 165218 91826 165454
rect 92062 165218 92146 165454
rect 92382 165218 92414 165454
rect 91794 165134 92414 165218
rect 91794 164898 91826 165134
rect 92062 164898 92146 165134
rect 92382 164898 92414 165134
rect 91794 129454 92414 164898
rect 91794 129218 91826 129454
rect 92062 129218 92146 129454
rect 92382 129218 92414 129454
rect 91794 129134 92414 129218
rect 91794 128898 91826 129134
rect 92062 128898 92146 129134
rect 92382 128898 92414 129134
rect 91794 93454 92414 128898
rect 91794 93218 91826 93454
rect 92062 93218 92146 93454
rect 92382 93218 92414 93454
rect 91794 93134 92414 93218
rect 91794 92898 91826 93134
rect 92062 92898 92146 93134
rect 92382 92898 92414 93134
rect 91794 57454 92414 92898
rect 91794 57218 91826 57454
rect 92062 57218 92146 57454
rect 92382 57218 92414 57454
rect 91794 57134 92414 57218
rect 91794 56898 91826 57134
rect 92062 56898 92146 57134
rect 92382 56898 92414 57134
rect 91794 21454 92414 56898
rect 91794 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 92414 21454
rect 91794 21134 92414 21218
rect 91794 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 92414 21134
rect 91794 -4186 92414 20898
rect 91794 -4422 91826 -4186
rect 92062 -4422 92146 -4186
rect 92382 -4422 92414 -4186
rect 91794 -4506 92414 -4422
rect 91794 -4742 91826 -4506
rect 92062 -4742 92146 -4506
rect 92382 -4742 92414 -4506
rect 91794 -7654 92414 -4742
rect 96294 709638 96914 711590
rect 96294 709402 96326 709638
rect 96562 709402 96646 709638
rect 96882 709402 96914 709638
rect 96294 709318 96914 709402
rect 96294 709082 96326 709318
rect 96562 709082 96646 709318
rect 96882 709082 96914 709318
rect 96294 673954 96914 709082
rect 96294 673718 96326 673954
rect 96562 673718 96646 673954
rect 96882 673718 96914 673954
rect 96294 673634 96914 673718
rect 96294 673398 96326 673634
rect 96562 673398 96646 673634
rect 96882 673398 96914 673634
rect 96294 637954 96914 673398
rect 96294 637718 96326 637954
rect 96562 637718 96646 637954
rect 96882 637718 96914 637954
rect 96294 637634 96914 637718
rect 96294 637398 96326 637634
rect 96562 637398 96646 637634
rect 96882 637398 96914 637634
rect 96294 601954 96914 637398
rect 96294 601718 96326 601954
rect 96562 601718 96646 601954
rect 96882 601718 96914 601954
rect 96294 601634 96914 601718
rect 96294 601398 96326 601634
rect 96562 601398 96646 601634
rect 96882 601398 96914 601634
rect 96294 565954 96914 601398
rect 96294 565718 96326 565954
rect 96562 565718 96646 565954
rect 96882 565718 96914 565954
rect 96294 565634 96914 565718
rect 96294 565398 96326 565634
rect 96562 565398 96646 565634
rect 96882 565398 96914 565634
rect 96294 529954 96914 565398
rect 96294 529718 96326 529954
rect 96562 529718 96646 529954
rect 96882 529718 96914 529954
rect 96294 529634 96914 529718
rect 96294 529398 96326 529634
rect 96562 529398 96646 529634
rect 96882 529398 96914 529634
rect 96294 493954 96914 529398
rect 96294 493718 96326 493954
rect 96562 493718 96646 493954
rect 96882 493718 96914 493954
rect 96294 493634 96914 493718
rect 96294 493398 96326 493634
rect 96562 493398 96646 493634
rect 96882 493398 96914 493634
rect 96294 457954 96914 493398
rect 96294 457718 96326 457954
rect 96562 457718 96646 457954
rect 96882 457718 96914 457954
rect 96294 457634 96914 457718
rect 96294 457398 96326 457634
rect 96562 457398 96646 457634
rect 96882 457398 96914 457634
rect 96294 421954 96914 457398
rect 96294 421718 96326 421954
rect 96562 421718 96646 421954
rect 96882 421718 96914 421954
rect 96294 421634 96914 421718
rect 96294 421398 96326 421634
rect 96562 421398 96646 421634
rect 96882 421398 96914 421634
rect 96294 385954 96914 421398
rect 96294 385718 96326 385954
rect 96562 385718 96646 385954
rect 96882 385718 96914 385954
rect 96294 385634 96914 385718
rect 96294 385398 96326 385634
rect 96562 385398 96646 385634
rect 96882 385398 96914 385634
rect 96294 349954 96914 385398
rect 96294 349718 96326 349954
rect 96562 349718 96646 349954
rect 96882 349718 96914 349954
rect 96294 349634 96914 349718
rect 96294 349398 96326 349634
rect 96562 349398 96646 349634
rect 96882 349398 96914 349634
rect 96294 313954 96914 349398
rect 96294 313718 96326 313954
rect 96562 313718 96646 313954
rect 96882 313718 96914 313954
rect 96294 313634 96914 313718
rect 96294 313398 96326 313634
rect 96562 313398 96646 313634
rect 96882 313398 96914 313634
rect 96294 277954 96914 313398
rect 96294 277718 96326 277954
rect 96562 277718 96646 277954
rect 96882 277718 96914 277954
rect 96294 277634 96914 277718
rect 96294 277398 96326 277634
rect 96562 277398 96646 277634
rect 96882 277398 96914 277634
rect 96294 241954 96914 277398
rect 96294 241718 96326 241954
rect 96562 241718 96646 241954
rect 96882 241718 96914 241954
rect 96294 241634 96914 241718
rect 96294 241398 96326 241634
rect 96562 241398 96646 241634
rect 96882 241398 96914 241634
rect 96294 205954 96914 241398
rect 96294 205718 96326 205954
rect 96562 205718 96646 205954
rect 96882 205718 96914 205954
rect 96294 205634 96914 205718
rect 96294 205398 96326 205634
rect 96562 205398 96646 205634
rect 96882 205398 96914 205634
rect 96294 169954 96914 205398
rect 100794 710598 101414 711590
rect 100794 710362 100826 710598
rect 101062 710362 101146 710598
rect 101382 710362 101414 710598
rect 100794 710278 101414 710362
rect 100794 710042 100826 710278
rect 101062 710042 101146 710278
rect 101382 710042 101414 710278
rect 100794 678454 101414 710042
rect 100794 678218 100826 678454
rect 101062 678218 101146 678454
rect 101382 678218 101414 678454
rect 100794 678134 101414 678218
rect 100794 677898 100826 678134
rect 101062 677898 101146 678134
rect 101382 677898 101414 678134
rect 100794 642454 101414 677898
rect 100794 642218 100826 642454
rect 101062 642218 101146 642454
rect 101382 642218 101414 642454
rect 100794 642134 101414 642218
rect 100794 641898 100826 642134
rect 101062 641898 101146 642134
rect 101382 641898 101414 642134
rect 100794 606454 101414 641898
rect 100794 606218 100826 606454
rect 101062 606218 101146 606454
rect 101382 606218 101414 606454
rect 100794 606134 101414 606218
rect 100794 605898 100826 606134
rect 101062 605898 101146 606134
rect 101382 605898 101414 606134
rect 100794 570454 101414 605898
rect 100794 570218 100826 570454
rect 101062 570218 101146 570454
rect 101382 570218 101414 570454
rect 100794 570134 101414 570218
rect 100794 569898 100826 570134
rect 101062 569898 101146 570134
rect 101382 569898 101414 570134
rect 100794 534454 101414 569898
rect 100794 534218 100826 534454
rect 101062 534218 101146 534454
rect 101382 534218 101414 534454
rect 100794 534134 101414 534218
rect 100794 533898 100826 534134
rect 101062 533898 101146 534134
rect 101382 533898 101414 534134
rect 100794 498454 101414 533898
rect 100794 498218 100826 498454
rect 101062 498218 101146 498454
rect 101382 498218 101414 498454
rect 100794 498134 101414 498218
rect 100794 497898 100826 498134
rect 101062 497898 101146 498134
rect 101382 497898 101414 498134
rect 100794 462454 101414 497898
rect 100794 462218 100826 462454
rect 101062 462218 101146 462454
rect 101382 462218 101414 462454
rect 100794 462134 101414 462218
rect 100794 461898 100826 462134
rect 101062 461898 101146 462134
rect 101382 461898 101414 462134
rect 100794 426454 101414 461898
rect 100794 426218 100826 426454
rect 101062 426218 101146 426454
rect 101382 426218 101414 426454
rect 100794 426134 101414 426218
rect 100794 425898 100826 426134
rect 101062 425898 101146 426134
rect 101382 425898 101414 426134
rect 100794 390454 101414 425898
rect 100794 390218 100826 390454
rect 101062 390218 101146 390454
rect 101382 390218 101414 390454
rect 100794 390134 101414 390218
rect 100794 389898 100826 390134
rect 101062 389898 101146 390134
rect 101382 389898 101414 390134
rect 100794 354454 101414 389898
rect 100794 354218 100826 354454
rect 101062 354218 101146 354454
rect 101382 354218 101414 354454
rect 100794 354134 101414 354218
rect 100794 353898 100826 354134
rect 101062 353898 101146 354134
rect 101382 353898 101414 354134
rect 100794 318454 101414 353898
rect 100794 318218 100826 318454
rect 101062 318218 101146 318454
rect 101382 318218 101414 318454
rect 100794 318134 101414 318218
rect 100794 317898 100826 318134
rect 101062 317898 101146 318134
rect 101382 317898 101414 318134
rect 100794 282454 101414 317898
rect 100794 282218 100826 282454
rect 101062 282218 101146 282454
rect 101382 282218 101414 282454
rect 100794 282134 101414 282218
rect 100794 281898 100826 282134
rect 101062 281898 101146 282134
rect 101382 281898 101414 282134
rect 100794 246454 101414 281898
rect 100794 246218 100826 246454
rect 101062 246218 101146 246454
rect 101382 246218 101414 246454
rect 100794 246134 101414 246218
rect 100794 245898 100826 246134
rect 101062 245898 101146 246134
rect 101382 245898 101414 246134
rect 100794 210454 101414 245898
rect 100794 210218 100826 210454
rect 101062 210218 101146 210454
rect 101382 210218 101414 210454
rect 100794 210134 101414 210218
rect 100794 209898 100826 210134
rect 101062 209898 101146 210134
rect 101382 209898 101414 210134
rect 100339 195668 100405 195669
rect 100339 195604 100340 195668
rect 100404 195604 100405 195668
rect 100339 195603 100405 195604
rect 96294 169718 96326 169954
rect 96562 169718 96646 169954
rect 96882 169718 96914 169954
rect 96294 169634 96914 169718
rect 96294 169398 96326 169634
rect 96562 169398 96646 169634
rect 96882 169398 96914 169634
rect 96294 133954 96914 169398
rect 96294 133718 96326 133954
rect 96562 133718 96646 133954
rect 96882 133718 96914 133954
rect 96294 133634 96914 133718
rect 96294 133398 96326 133634
rect 96562 133398 96646 133634
rect 96882 133398 96914 133634
rect 96294 97954 96914 133398
rect 96294 97718 96326 97954
rect 96562 97718 96646 97954
rect 96882 97718 96914 97954
rect 96294 97634 96914 97718
rect 96294 97398 96326 97634
rect 96562 97398 96646 97634
rect 96882 97398 96914 97634
rect 96294 61954 96914 97398
rect 100342 63477 100402 195603
rect 100523 193900 100589 193901
rect 100523 193836 100524 193900
rect 100588 193836 100589 193900
rect 100523 193835 100589 193836
rect 100339 63476 100405 63477
rect 100339 63412 100340 63476
rect 100404 63412 100405 63476
rect 100339 63411 100405 63412
rect 100342 62797 100402 63411
rect 100339 62796 100405 62797
rect 100339 62732 100340 62796
rect 100404 62732 100405 62796
rect 100339 62731 100405 62732
rect 96294 61718 96326 61954
rect 96562 61718 96646 61954
rect 96882 61718 96914 61954
rect 96294 61634 96914 61718
rect 96294 61398 96326 61634
rect 96562 61398 96646 61634
rect 96882 61398 96914 61634
rect 96294 25954 96914 61398
rect 100526 56541 100586 193835
rect 100794 174454 101414 209898
rect 105294 711558 105914 711590
rect 105294 711322 105326 711558
rect 105562 711322 105646 711558
rect 105882 711322 105914 711558
rect 105294 711238 105914 711322
rect 105294 711002 105326 711238
rect 105562 711002 105646 711238
rect 105882 711002 105914 711238
rect 105294 682954 105914 711002
rect 105294 682718 105326 682954
rect 105562 682718 105646 682954
rect 105882 682718 105914 682954
rect 105294 682634 105914 682718
rect 105294 682398 105326 682634
rect 105562 682398 105646 682634
rect 105882 682398 105914 682634
rect 105294 646954 105914 682398
rect 105294 646718 105326 646954
rect 105562 646718 105646 646954
rect 105882 646718 105914 646954
rect 105294 646634 105914 646718
rect 105294 646398 105326 646634
rect 105562 646398 105646 646634
rect 105882 646398 105914 646634
rect 105294 610954 105914 646398
rect 105294 610718 105326 610954
rect 105562 610718 105646 610954
rect 105882 610718 105914 610954
rect 105294 610634 105914 610718
rect 105294 610398 105326 610634
rect 105562 610398 105646 610634
rect 105882 610398 105914 610634
rect 105294 574954 105914 610398
rect 105294 574718 105326 574954
rect 105562 574718 105646 574954
rect 105882 574718 105914 574954
rect 105294 574634 105914 574718
rect 105294 574398 105326 574634
rect 105562 574398 105646 574634
rect 105882 574398 105914 574634
rect 105294 538954 105914 574398
rect 105294 538718 105326 538954
rect 105562 538718 105646 538954
rect 105882 538718 105914 538954
rect 105294 538634 105914 538718
rect 105294 538398 105326 538634
rect 105562 538398 105646 538634
rect 105882 538398 105914 538634
rect 105294 502954 105914 538398
rect 105294 502718 105326 502954
rect 105562 502718 105646 502954
rect 105882 502718 105914 502954
rect 105294 502634 105914 502718
rect 105294 502398 105326 502634
rect 105562 502398 105646 502634
rect 105882 502398 105914 502634
rect 105294 466954 105914 502398
rect 105294 466718 105326 466954
rect 105562 466718 105646 466954
rect 105882 466718 105914 466954
rect 105294 466634 105914 466718
rect 105294 466398 105326 466634
rect 105562 466398 105646 466634
rect 105882 466398 105914 466634
rect 105294 430954 105914 466398
rect 105294 430718 105326 430954
rect 105562 430718 105646 430954
rect 105882 430718 105914 430954
rect 105294 430634 105914 430718
rect 105294 430398 105326 430634
rect 105562 430398 105646 430634
rect 105882 430398 105914 430634
rect 105294 394954 105914 430398
rect 105294 394718 105326 394954
rect 105562 394718 105646 394954
rect 105882 394718 105914 394954
rect 105294 394634 105914 394718
rect 105294 394398 105326 394634
rect 105562 394398 105646 394634
rect 105882 394398 105914 394634
rect 105294 358954 105914 394398
rect 105294 358718 105326 358954
rect 105562 358718 105646 358954
rect 105882 358718 105914 358954
rect 105294 358634 105914 358718
rect 105294 358398 105326 358634
rect 105562 358398 105646 358634
rect 105882 358398 105914 358634
rect 105294 322954 105914 358398
rect 105294 322718 105326 322954
rect 105562 322718 105646 322954
rect 105882 322718 105914 322954
rect 105294 322634 105914 322718
rect 105294 322398 105326 322634
rect 105562 322398 105646 322634
rect 105882 322398 105914 322634
rect 105294 286954 105914 322398
rect 105294 286718 105326 286954
rect 105562 286718 105646 286954
rect 105882 286718 105914 286954
rect 105294 286634 105914 286718
rect 105294 286398 105326 286634
rect 105562 286398 105646 286634
rect 105882 286398 105914 286634
rect 105294 250954 105914 286398
rect 109794 704838 110414 711590
rect 109794 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 110414 704838
rect 109794 704518 110414 704602
rect 109794 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 110414 704518
rect 109794 687454 110414 704282
rect 109794 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 110414 687454
rect 109794 687134 110414 687218
rect 109794 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 110414 687134
rect 109794 651454 110414 686898
rect 109794 651218 109826 651454
rect 110062 651218 110146 651454
rect 110382 651218 110414 651454
rect 109794 651134 110414 651218
rect 109794 650898 109826 651134
rect 110062 650898 110146 651134
rect 110382 650898 110414 651134
rect 109794 615454 110414 650898
rect 109794 615218 109826 615454
rect 110062 615218 110146 615454
rect 110382 615218 110414 615454
rect 109794 615134 110414 615218
rect 109794 614898 109826 615134
rect 110062 614898 110146 615134
rect 110382 614898 110414 615134
rect 109794 579454 110414 614898
rect 109794 579218 109826 579454
rect 110062 579218 110146 579454
rect 110382 579218 110414 579454
rect 109794 579134 110414 579218
rect 109794 578898 109826 579134
rect 110062 578898 110146 579134
rect 110382 578898 110414 579134
rect 109794 543454 110414 578898
rect 109794 543218 109826 543454
rect 110062 543218 110146 543454
rect 110382 543218 110414 543454
rect 109794 543134 110414 543218
rect 109794 542898 109826 543134
rect 110062 542898 110146 543134
rect 110382 542898 110414 543134
rect 109794 507454 110414 542898
rect 109794 507218 109826 507454
rect 110062 507218 110146 507454
rect 110382 507218 110414 507454
rect 109794 507134 110414 507218
rect 109794 506898 109826 507134
rect 110062 506898 110146 507134
rect 110382 506898 110414 507134
rect 109794 471454 110414 506898
rect 109794 471218 109826 471454
rect 110062 471218 110146 471454
rect 110382 471218 110414 471454
rect 109794 471134 110414 471218
rect 109794 470898 109826 471134
rect 110062 470898 110146 471134
rect 110382 470898 110414 471134
rect 109794 435454 110414 470898
rect 109794 435218 109826 435454
rect 110062 435218 110146 435454
rect 110382 435218 110414 435454
rect 109794 435134 110414 435218
rect 109794 434898 109826 435134
rect 110062 434898 110146 435134
rect 110382 434898 110414 435134
rect 109794 399454 110414 434898
rect 109794 399218 109826 399454
rect 110062 399218 110146 399454
rect 110382 399218 110414 399454
rect 109794 399134 110414 399218
rect 109794 398898 109826 399134
rect 110062 398898 110146 399134
rect 110382 398898 110414 399134
rect 109794 363454 110414 398898
rect 109794 363218 109826 363454
rect 110062 363218 110146 363454
rect 110382 363218 110414 363454
rect 109794 363134 110414 363218
rect 109794 362898 109826 363134
rect 110062 362898 110146 363134
rect 110382 362898 110414 363134
rect 109794 327454 110414 362898
rect 109794 327218 109826 327454
rect 110062 327218 110146 327454
rect 110382 327218 110414 327454
rect 109794 327134 110414 327218
rect 109794 326898 109826 327134
rect 110062 326898 110146 327134
rect 110382 326898 110414 327134
rect 109794 291454 110414 326898
rect 109794 291218 109826 291454
rect 110062 291218 110146 291454
rect 110382 291218 110414 291454
rect 109794 291134 110414 291218
rect 109794 290898 109826 291134
rect 110062 290898 110146 291134
rect 110382 290898 110414 291134
rect 108803 265028 108869 265029
rect 108803 264964 108804 265028
rect 108868 264964 108869 265028
rect 108803 264963 108869 264964
rect 105294 250718 105326 250954
rect 105562 250718 105646 250954
rect 105882 250718 105914 250954
rect 105294 250634 105914 250718
rect 105294 250398 105326 250634
rect 105562 250398 105646 250634
rect 105882 250398 105914 250634
rect 105294 214954 105914 250398
rect 105294 214718 105326 214954
rect 105562 214718 105646 214954
rect 105882 214718 105914 214954
rect 105294 214634 105914 214718
rect 105294 214398 105326 214634
rect 105562 214398 105646 214634
rect 105882 214398 105914 214634
rect 103283 192948 103349 192949
rect 103283 192884 103284 192948
rect 103348 192884 103349 192948
rect 103283 192883 103349 192884
rect 100794 174218 100826 174454
rect 101062 174218 101146 174454
rect 101382 174218 101414 174454
rect 100794 174134 101414 174218
rect 100794 173898 100826 174134
rect 101062 173898 101146 174134
rect 101382 173898 101414 174134
rect 100794 138454 101414 173898
rect 103099 148612 103165 148613
rect 103099 148548 103100 148612
rect 103164 148548 103165 148612
rect 103099 148547 103165 148548
rect 100794 138218 100826 138454
rect 101062 138218 101146 138454
rect 101382 138218 101414 138454
rect 100794 138134 101414 138218
rect 100794 137898 100826 138134
rect 101062 137898 101146 138134
rect 101382 137898 101414 138134
rect 100794 102454 101414 137898
rect 100794 102218 100826 102454
rect 101062 102218 101146 102454
rect 101382 102218 101414 102454
rect 100794 102134 101414 102218
rect 100794 101898 100826 102134
rect 101062 101898 101146 102134
rect 101382 101898 101414 102134
rect 100794 66454 101414 101898
rect 102179 78164 102245 78165
rect 102179 78100 102180 78164
rect 102244 78100 102245 78164
rect 102179 78099 102245 78100
rect 102182 77349 102242 78099
rect 102179 77348 102245 77349
rect 102179 77284 102180 77348
rect 102244 77284 102245 77348
rect 102179 77283 102245 77284
rect 100794 66218 100826 66454
rect 101062 66218 101146 66454
rect 101382 66218 101414 66454
rect 100794 66134 101414 66218
rect 100794 65898 100826 66134
rect 101062 65898 101146 66134
rect 101382 65898 101414 66134
rect 99419 56540 99485 56541
rect 99419 56476 99420 56540
rect 99484 56476 99485 56540
rect 99419 56475 99485 56476
rect 100523 56540 100589 56541
rect 100523 56476 100524 56540
rect 100588 56476 100589 56540
rect 100523 56475 100589 56476
rect 99422 55861 99482 56475
rect 99419 55860 99485 55861
rect 99419 55796 99420 55860
rect 99484 55796 99485 55860
rect 99419 55795 99485 55796
rect 96294 25718 96326 25954
rect 96562 25718 96646 25954
rect 96882 25718 96914 25954
rect 96294 25634 96914 25718
rect 96294 25398 96326 25634
rect 96562 25398 96646 25634
rect 96882 25398 96914 25634
rect 96294 -5146 96914 25398
rect 96294 -5382 96326 -5146
rect 96562 -5382 96646 -5146
rect 96882 -5382 96914 -5146
rect 96294 -5466 96914 -5382
rect 96294 -5702 96326 -5466
rect 96562 -5702 96646 -5466
rect 96882 -5702 96914 -5466
rect 96294 -7654 96914 -5702
rect 100794 30454 101414 65898
rect 103102 53821 103162 148547
rect 103286 77349 103346 192883
rect 104019 192812 104085 192813
rect 104019 192748 104020 192812
rect 104084 192748 104085 192812
rect 104019 192747 104085 192748
rect 103283 77348 103349 77349
rect 103283 77284 103284 77348
rect 103348 77284 103349 77348
rect 103283 77283 103349 77284
rect 104022 65517 104082 192747
rect 105294 178954 105914 214398
rect 106779 200428 106845 200429
rect 106779 200364 106780 200428
rect 106844 200364 106845 200428
rect 106779 200363 106845 200364
rect 105294 178718 105326 178954
rect 105562 178718 105646 178954
rect 105882 178718 105914 178954
rect 105294 178634 105914 178718
rect 105294 178398 105326 178634
rect 105562 178398 105646 178634
rect 105882 178398 105914 178634
rect 104203 148476 104269 148477
rect 104203 148412 104204 148476
rect 104268 148412 104269 148476
rect 104203 148411 104269 148412
rect 104019 65516 104085 65517
rect 104019 65452 104020 65516
rect 104084 65452 104085 65516
rect 104019 65451 104085 65452
rect 104206 55997 104266 148411
rect 105294 142954 105914 178398
rect 105294 142718 105326 142954
rect 105562 142718 105646 142954
rect 105882 142718 105914 142954
rect 105294 142634 105914 142718
rect 105294 142398 105326 142634
rect 105562 142398 105646 142634
rect 105882 142398 105914 142634
rect 105294 106954 105914 142398
rect 105294 106718 105326 106954
rect 105562 106718 105646 106954
rect 105882 106718 105914 106954
rect 105294 106634 105914 106718
rect 105294 106398 105326 106634
rect 105562 106398 105646 106634
rect 105882 106398 105914 106634
rect 105294 70954 105914 106398
rect 106782 74085 106842 200363
rect 107515 198388 107581 198389
rect 107515 198324 107516 198388
rect 107580 198324 107581 198388
rect 107515 198323 107581 198324
rect 107331 198252 107397 198253
rect 107331 198188 107332 198252
rect 107396 198188 107397 198252
rect 107331 198187 107397 198188
rect 107334 77485 107394 198187
rect 107331 77484 107397 77485
rect 107331 77420 107332 77484
rect 107396 77420 107397 77484
rect 107331 77419 107397 77420
rect 106779 74084 106845 74085
rect 106779 74020 106780 74084
rect 106844 74020 106845 74084
rect 106779 74019 106845 74020
rect 107518 71229 107578 198323
rect 108251 196892 108317 196893
rect 108251 196828 108252 196892
rect 108316 196828 108317 196892
rect 108251 196827 108317 196828
rect 108254 73133 108314 196827
rect 108435 187508 108501 187509
rect 108435 187444 108436 187508
rect 108500 187444 108501 187508
rect 108435 187443 108501 187444
rect 108251 73132 108317 73133
rect 108251 73068 108252 73132
rect 108316 73068 108317 73132
rect 108251 73067 108317 73068
rect 107515 71228 107581 71229
rect 107515 71164 107516 71228
rect 107580 71164 107581 71228
rect 107515 71163 107581 71164
rect 105294 70718 105326 70954
rect 105562 70718 105646 70954
rect 105882 70718 105914 70954
rect 105294 70634 105914 70718
rect 105294 70398 105326 70634
rect 105562 70398 105646 70634
rect 105882 70398 105914 70634
rect 104203 55996 104269 55997
rect 104203 55932 104204 55996
rect 104268 55932 104269 55996
rect 104203 55931 104269 55932
rect 103099 53820 103165 53821
rect 103099 53756 103100 53820
rect 103164 53756 103165 53820
rect 103099 53755 103165 53756
rect 100794 30218 100826 30454
rect 101062 30218 101146 30454
rect 101382 30218 101414 30454
rect 100794 30134 101414 30218
rect 100794 29898 100826 30134
rect 101062 29898 101146 30134
rect 101382 29898 101414 30134
rect 100794 -6106 101414 29898
rect 100794 -6342 100826 -6106
rect 101062 -6342 101146 -6106
rect 101382 -6342 101414 -6106
rect 100794 -6426 101414 -6342
rect 100794 -6662 100826 -6426
rect 101062 -6662 101146 -6426
rect 101382 -6662 101414 -6426
rect 100794 -7654 101414 -6662
rect 105294 34954 105914 70398
rect 108438 65653 108498 187443
rect 108806 141813 108866 264963
rect 109794 255454 110414 290898
rect 114294 705798 114914 711590
rect 114294 705562 114326 705798
rect 114562 705562 114646 705798
rect 114882 705562 114914 705798
rect 114294 705478 114914 705562
rect 114294 705242 114326 705478
rect 114562 705242 114646 705478
rect 114882 705242 114914 705478
rect 114294 691954 114914 705242
rect 114294 691718 114326 691954
rect 114562 691718 114646 691954
rect 114882 691718 114914 691954
rect 114294 691634 114914 691718
rect 114294 691398 114326 691634
rect 114562 691398 114646 691634
rect 114882 691398 114914 691634
rect 114294 655954 114914 691398
rect 114294 655718 114326 655954
rect 114562 655718 114646 655954
rect 114882 655718 114914 655954
rect 114294 655634 114914 655718
rect 114294 655398 114326 655634
rect 114562 655398 114646 655634
rect 114882 655398 114914 655634
rect 114294 619954 114914 655398
rect 114294 619718 114326 619954
rect 114562 619718 114646 619954
rect 114882 619718 114914 619954
rect 114294 619634 114914 619718
rect 114294 619398 114326 619634
rect 114562 619398 114646 619634
rect 114882 619398 114914 619634
rect 114294 583954 114914 619398
rect 114294 583718 114326 583954
rect 114562 583718 114646 583954
rect 114882 583718 114914 583954
rect 114294 583634 114914 583718
rect 114294 583398 114326 583634
rect 114562 583398 114646 583634
rect 114882 583398 114914 583634
rect 114294 547954 114914 583398
rect 114294 547718 114326 547954
rect 114562 547718 114646 547954
rect 114882 547718 114914 547954
rect 114294 547634 114914 547718
rect 114294 547398 114326 547634
rect 114562 547398 114646 547634
rect 114882 547398 114914 547634
rect 114294 511954 114914 547398
rect 114294 511718 114326 511954
rect 114562 511718 114646 511954
rect 114882 511718 114914 511954
rect 114294 511634 114914 511718
rect 114294 511398 114326 511634
rect 114562 511398 114646 511634
rect 114882 511398 114914 511634
rect 114294 475954 114914 511398
rect 114294 475718 114326 475954
rect 114562 475718 114646 475954
rect 114882 475718 114914 475954
rect 114294 475634 114914 475718
rect 114294 475398 114326 475634
rect 114562 475398 114646 475634
rect 114882 475398 114914 475634
rect 114294 439954 114914 475398
rect 114294 439718 114326 439954
rect 114562 439718 114646 439954
rect 114882 439718 114914 439954
rect 114294 439634 114914 439718
rect 114294 439398 114326 439634
rect 114562 439398 114646 439634
rect 114882 439398 114914 439634
rect 114294 403954 114914 439398
rect 114294 403718 114326 403954
rect 114562 403718 114646 403954
rect 114882 403718 114914 403954
rect 114294 403634 114914 403718
rect 114294 403398 114326 403634
rect 114562 403398 114646 403634
rect 114882 403398 114914 403634
rect 114294 367954 114914 403398
rect 114294 367718 114326 367954
rect 114562 367718 114646 367954
rect 114882 367718 114914 367954
rect 114294 367634 114914 367718
rect 114294 367398 114326 367634
rect 114562 367398 114646 367634
rect 114882 367398 114914 367634
rect 114294 331954 114914 367398
rect 114294 331718 114326 331954
rect 114562 331718 114646 331954
rect 114882 331718 114914 331954
rect 114294 331634 114914 331718
rect 114294 331398 114326 331634
rect 114562 331398 114646 331634
rect 114882 331398 114914 331634
rect 114294 295954 114914 331398
rect 114294 295718 114326 295954
rect 114562 295718 114646 295954
rect 114882 295718 114914 295954
rect 114294 295634 114914 295718
rect 114294 295398 114326 295634
rect 114562 295398 114646 295634
rect 114882 295398 114914 295634
rect 111563 265164 111629 265165
rect 111563 265100 111564 265164
rect 111628 265100 111629 265164
rect 111563 265099 111629 265100
rect 111195 263124 111261 263125
rect 111195 263060 111196 263124
rect 111260 263060 111261 263124
rect 111195 263059 111261 263060
rect 111011 262988 111077 262989
rect 111011 262924 111012 262988
rect 111076 262924 111077 262988
rect 111011 262923 111077 262924
rect 109794 255218 109826 255454
rect 110062 255218 110146 255454
rect 110382 255218 110414 255454
rect 109794 255134 110414 255218
rect 109794 254898 109826 255134
rect 110062 254898 110146 255134
rect 110382 254898 110414 255134
rect 109794 219454 110414 254898
rect 109794 219218 109826 219454
rect 110062 219218 110146 219454
rect 110382 219218 110414 219454
rect 109794 219134 110414 219218
rect 109794 218898 109826 219134
rect 110062 218898 110146 219134
rect 110382 218898 110414 219134
rect 109539 191724 109605 191725
rect 109539 191660 109540 191724
rect 109604 191660 109605 191724
rect 109539 191659 109605 191660
rect 108803 141812 108869 141813
rect 108803 141748 108804 141812
rect 108868 141748 108869 141812
rect 108803 141747 108869 141748
rect 109542 66877 109602 191659
rect 109794 183454 110414 218898
rect 109794 183218 109826 183454
rect 110062 183218 110146 183454
rect 110382 183218 110414 183454
rect 109794 183134 110414 183218
rect 109794 182898 109826 183134
rect 110062 182898 110146 183134
rect 110382 182898 110414 183134
rect 109794 147454 110414 182898
rect 109794 147218 109826 147454
rect 110062 147218 110146 147454
rect 110382 147218 110414 147454
rect 109794 147134 110414 147218
rect 109794 146898 109826 147134
rect 110062 146898 110146 147134
rect 110382 146898 110414 147134
rect 109794 111454 110414 146898
rect 111014 145893 111074 262923
rect 111011 145892 111077 145893
rect 111011 145828 111012 145892
rect 111076 145828 111077 145892
rect 111011 145827 111077 145828
rect 111198 143173 111258 263059
rect 111379 262444 111445 262445
rect 111379 262380 111380 262444
rect 111444 262380 111445 262444
rect 111379 262379 111445 262380
rect 111195 143172 111261 143173
rect 111195 143108 111196 143172
rect 111260 143108 111261 143172
rect 111195 143107 111261 143108
rect 111011 142220 111077 142221
rect 111011 142156 111012 142220
rect 111076 142156 111077 142220
rect 111011 142155 111077 142156
rect 109794 111218 109826 111454
rect 110062 111218 110146 111454
rect 110382 111218 110414 111454
rect 109794 111134 110414 111218
rect 109794 110898 109826 111134
rect 110062 110898 110146 111134
rect 110382 110898 110414 111134
rect 109794 75454 110414 110898
rect 109794 75218 109826 75454
rect 110062 75218 110146 75454
rect 110382 75218 110414 75454
rect 109794 75134 110414 75218
rect 109794 74898 109826 75134
rect 110062 74898 110146 75134
rect 110382 74898 110414 75134
rect 109539 66876 109605 66877
rect 109539 66812 109540 66876
rect 109604 66812 109605 66876
rect 109539 66811 109605 66812
rect 108435 65652 108501 65653
rect 108435 65588 108436 65652
rect 108500 65588 108501 65652
rect 108435 65587 108501 65588
rect 105294 34718 105326 34954
rect 105562 34718 105646 34954
rect 105882 34718 105914 34954
rect 105294 34634 105914 34718
rect 105294 34398 105326 34634
rect 105562 34398 105646 34634
rect 105882 34398 105914 34634
rect 105294 -7066 105914 34398
rect 105294 -7302 105326 -7066
rect 105562 -7302 105646 -7066
rect 105882 -7302 105914 -7066
rect 105294 -7386 105914 -7302
rect 105294 -7622 105326 -7386
rect 105562 -7622 105646 -7386
rect 105882 -7622 105914 -7386
rect 105294 -7654 105914 -7622
rect 109794 39454 110414 74898
rect 111014 58037 111074 142155
rect 111382 142085 111442 262379
rect 111566 144669 111626 265099
rect 113035 263668 113101 263669
rect 113035 263604 113036 263668
rect 113100 263604 113101 263668
rect 113035 263603 113101 263604
rect 112851 262852 112917 262853
rect 112851 262788 112852 262852
rect 112916 262788 112917 262852
rect 112851 262787 112917 262788
rect 112667 261084 112733 261085
rect 112667 261020 112668 261084
rect 112732 261020 112733 261084
rect 112667 261019 112733 261020
rect 112483 147524 112549 147525
rect 112483 147460 112484 147524
rect 112548 147460 112549 147524
rect 112483 147459 112549 147460
rect 112115 145756 112181 145757
rect 112115 145692 112116 145756
rect 112180 145692 112181 145756
rect 112115 145691 112181 145692
rect 111563 144668 111629 144669
rect 111563 144604 111564 144668
rect 111628 144604 111629 144668
rect 111563 144603 111629 144604
rect 111379 142084 111445 142085
rect 111379 142020 111380 142084
rect 111444 142020 111445 142084
rect 111379 142019 111445 142020
rect 111563 139364 111629 139365
rect 111563 139300 111564 139364
rect 111628 139300 111629 139364
rect 111563 139299 111629 139300
rect 111195 139092 111261 139093
rect 111195 139028 111196 139092
rect 111260 139028 111261 139092
rect 111195 139027 111261 139028
rect 111198 64157 111258 139027
rect 111566 68373 111626 139299
rect 112118 81837 112178 145691
rect 112299 140180 112365 140181
rect 112299 140116 112300 140180
rect 112364 140116 112365 140180
rect 112299 140115 112365 140116
rect 112115 81836 112181 81837
rect 112115 81772 112116 81836
rect 112180 81772 112181 81836
rect 112115 81771 112181 81772
rect 112302 73677 112362 140115
rect 112299 73676 112365 73677
rect 112299 73612 112300 73676
rect 112364 73612 112365 73676
rect 112299 73611 112365 73612
rect 111563 68372 111629 68373
rect 111563 68308 111564 68372
rect 111628 68308 111629 68372
rect 111563 68307 111629 68308
rect 111195 64156 111261 64157
rect 111195 64092 111196 64156
rect 111260 64092 111261 64156
rect 111195 64091 111261 64092
rect 111747 59260 111813 59261
rect 111747 59196 111748 59260
rect 111812 59196 111813 59260
rect 111747 59195 111813 59196
rect 111750 58717 111810 59195
rect 112486 58853 112546 147459
rect 112670 144397 112730 261019
rect 112854 145893 112914 262787
rect 112851 145892 112917 145893
rect 112851 145828 112852 145892
rect 112916 145828 112917 145892
rect 112851 145827 112917 145828
rect 113038 144805 113098 263603
rect 114139 262580 114205 262581
rect 114139 262516 114140 262580
rect 114204 262516 114205 262580
rect 114139 262515 114205 262516
rect 113955 259588 114021 259589
rect 113955 259524 113956 259588
rect 114020 259524 114021 259588
rect 113955 259523 114021 259524
rect 113587 147388 113653 147389
rect 113587 147324 113588 147388
rect 113652 147324 113653 147388
rect 113587 147323 113653 147324
rect 113035 144804 113101 144805
rect 113035 144740 113036 144804
rect 113100 144740 113101 144804
rect 113035 144739 113101 144740
rect 112667 144396 112733 144397
rect 112667 144332 112668 144396
rect 112732 144332 112733 144396
rect 112667 144331 112733 144332
rect 112851 137324 112917 137325
rect 112851 137260 112852 137324
rect 112916 137260 112917 137324
rect 112851 137259 112917 137260
rect 112854 59261 112914 137259
rect 113590 73949 113650 147323
rect 113958 143309 114018 259523
rect 114142 144533 114202 262515
rect 114294 259954 114914 295398
rect 118794 706758 119414 711590
rect 118794 706522 118826 706758
rect 119062 706522 119146 706758
rect 119382 706522 119414 706758
rect 118794 706438 119414 706522
rect 118794 706202 118826 706438
rect 119062 706202 119146 706438
rect 119382 706202 119414 706438
rect 118794 696454 119414 706202
rect 118794 696218 118826 696454
rect 119062 696218 119146 696454
rect 119382 696218 119414 696454
rect 118794 696134 119414 696218
rect 118794 695898 118826 696134
rect 119062 695898 119146 696134
rect 119382 695898 119414 696134
rect 118794 660454 119414 695898
rect 118794 660218 118826 660454
rect 119062 660218 119146 660454
rect 119382 660218 119414 660454
rect 118794 660134 119414 660218
rect 118794 659898 118826 660134
rect 119062 659898 119146 660134
rect 119382 659898 119414 660134
rect 118794 624454 119414 659898
rect 118794 624218 118826 624454
rect 119062 624218 119146 624454
rect 119382 624218 119414 624454
rect 118794 624134 119414 624218
rect 118794 623898 118826 624134
rect 119062 623898 119146 624134
rect 119382 623898 119414 624134
rect 118794 588454 119414 623898
rect 118794 588218 118826 588454
rect 119062 588218 119146 588454
rect 119382 588218 119414 588454
rect 118794 588134 119414 588218
rect 118794 587898 118826 588134
rect 119062 587898 119146 588134
rect 119382 587898 119414 588134
rect 118794 552454 119414 587898
rect 118794 552218 118826 552454
rect 119062 552218 119146 552454
rect 119382 552218 119414 552454
rect 118794 552134 119414 552218
rect 118794 551898 118826 552134
rect 119062 551898 119146 552134
rect 119382 551898 119414 552134
rect 118794 516454 119414 551898
rect 118794 516218 118826 516454
rect 119062 516218 119146 516454
rect 119382 516218 119414 516454
rect 118794 516134 119414 516218
rect 118794 515898 118826 516134
rect 119062 515898 119146 516134
rect 119382 515898 119414 516134
rect 118794 480454 119414 515898
rect 118794 480218 118826 480454
rect 119062 480218 119146 480454
rect 119382 480218 119414 480454
rect 118794 480134 119414 480218
rect 118794 479898 118826 480134
rect 119062 479898 119146 480134
rect 119382 479898 119414 480134
rect 118794 444454 119414 479898
rect 118794 444218 118826 444454
rect 119062 444218 119146 444454
rect 119382 444218 119414 444454
rect 118794 444134 119414 444218
rect 118794 443898 118826 444134
rect 119062 443898 119146 444134
rect 119382 443898 119414 444134
rect 118794 408454 119414 443898
rect 118794 408218 118826 408454
rect 119062 408218 119146 408454
rect 119382 408218 119414 408454
rect 118794 408134 119414 408218
rect 118794 407898 118826 408134
rect 119062 407898 119146 408134
rect 119382 407898 119414 408134
rect 118794 372454 119414 407898
rect 118794 372218 118826 372454
rect 119062 372218 119146 372454
rect 119382 372218 119414 372454
rect 118794 372134 119414 372218
rect 118794 371898 118826 372134
rect 119062 371898 119146 372134
rect 119382 371898 119414 372134
rect 118794 336454 119414 371898
rect 118794 336218 118826 336454
rect 119062 336218 119146 336454
rect 119382 336218 119414 336454
rect 118794 336134 119414 336218
rect 118794 335898 118826 336134
rect 119062 335898 119146 336134
rect 119382 335898 119414 336134
rect 118794 300454 119414 335898
rect 118794 300218 118826 300454
rect 119062 300218 119146 300454
rect 119382 300218 119414 300454
rect 118794 300134 119414 300218
rect 118794 299898 118826 300134
rect 119062 299898 119146 300134
rect 119382 299898 119414 300134
rect 118794 264454 119414 299898
rect 118794 264218 118826 264454
rect 119062 264218 119146 264454
rect 119382 264218 119414 264454
rect 118794 264134 119414 264218
rect 118794 263898 118826 264134
rect 119062 263898 119146 264134
rect 119382 263898 119414 264134
rect 116899 263804 116965 263805
rect 116899 263740 116900 263804
rect 116964 263740 116965 263804
rect 116899 263739 116965 263740
rect 115795 262716 115861 262717
rect 115795 262652 115796 262716
rect 115860 262652 115861 262716
rect 115795 262651 115861 262652
rect 115611 260404 115677 260405
rect 115611 260340 115612 260404
rect 115676 260340 115677 260404
rect 115611 260339 115677 260340
rect 114294 259718 114326 259954
rect 114562 259718 114646 259954
rect 114882 259718 114914 259954
rect 114294 259634 114914 259718
rect 114294 259398 114326 259634
rect 114562 259398 114646 259634
rect 114882 259398 114914 259634
rect 114294 223954 114914 259398
rect 114294 223718 114326 223954
rect 114562 223718 114646 223954
rect 114882 223718 114914 223954
rect 114294 223634 114914 223718
rect 114294 223398 114326 223634
rect 114562 223398 114646 223634
rect 114882 223398 114914 223634
rect 114294 187954 114914 223398
rect 114294 187718 114326 187954
rect 114562 187718 114646 187954
rect 114882 187718 114914 187954
rect 114294 187634 114914 187718
rect 114294 187398 114326 187634
rect 114562 187398 114646 187634
rect 114882 187398 114914 187634
rect 114294 151954 114914 187398
rect 114294 151718 114326 151954
rect 114562 151718 114646 151954
rect 114882 151718 114914 151954
rect 114294 151634 114914 151718
rect 114294 151398 114326 151634
rect 114562 151398 114646 151634
rect 114882 151398 114914 151634
rect 114139 144532 114205 144533
rect 114139 144468 114140 144532
rect 114204 144468 114205 144532
rect 114139 144467 114205 144468
rect 113955 143308 114021 143309
rect 113955 143244 113956 143308
rect 114020 143244 114021 143308
rect 113955 143243 114021 143244
rect 114139 141948 114205 141949
rect 114139 141884 114140 141948
rect 114204 141884 114205 141948
rect 114139 141883 114205 141884
rect 113771 141268 113837 141269
rect 113771 141204 113772 141268
rect 113836 141204 113837 141268
rect 113771 141203 113837 141204
rect 113774 76805 113834 141203
rect 113771 76804 113837 76805
rect 113771 76740 113772 76804
rect 113836 76740 113837 76804
rect 113771 76739 113837 76740
rect 113587 73948 113653 73949
rect 113587 73884 113588 73948
rect 113652 73884 113653 73948
rect 113587 73883 113653 73884
rect 114142 67421 114202 141883
rect 114294 115954 114914 151398
rect 115059 147252 115125 147253
rect 115059 147188 115060 147252
rect 115124 147188 115125 147252
rect 115059 147187 115125 147188
rect 114294 115718 114326 115954
rect 114562 115718 114646 115954
rect 114882 115718 114914 115954
rect 114294 115634 114914 115718
rect 114294 115398 114326 115634
rect 114562 115398 114646 115634
rect 114882 115398 114914 115634
rect 114294 79954 114914 115398
rect 114294 79718 114326 79954
rect 114562 79718 114646 79954
rect 114882 79718 114914 79954
rect 114294 79634 114914 79718
rect 114294 79398 114326 79634
rect 114562 79398 114646 79634
rect 114882 79398 114914 79634
rect 114139 67420 114205 67421
rect 114139 67356 114140 67420
rect 114204 67356 114205 67420
rect 114139 67355 114205 67356
rect 112851 59260 112917 59261
rect 112851 59196 112852 59260
rect 112916 59196 112917 59260
rect 112851 59195 112917 59196
rect 112483 58852 112549 58853
rect 112483 58788 112484 58852
rect 112548 58788 112549 58852
rect 112483 58787 112549 58788
rect 111747 58716 111813 58717
rect 111747 58652 111748 58716
rect 111812 58652 111813 58716
rect 111747 58651 111813 58652
rect 111011 58036 111077 58037
rect 111011 57972 111012 58036
rect 111076 57972 111077 58036
rect 111011 57971 111077 57972
rect 109794 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 110414 39454
rect 109794 39134 110414 39218
rect 109794 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 110414 39134
rect 109794 3454 110414 38898
rect 109794 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 110414 3454
rect 109794 3134 110414 3218
rect 109794 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 110414 3134
rect 109794 -346 110414 2898
rect 109794 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 110414 -346
rect 109794 -666 110414 -582
rect 109794 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 110414 -666
rect 109794 -7654 110414 -902
rect 114294 43954 114914 79398
rect 115062 63341 115122 147187
rect 115614 144805 115674 260339
rect 115798 146301 115858 262651
rect 116715 260540 116781 260541
rect 116715 260476 116716 260540
rect 116780 260476 116781 260540
rect 116715 260475 116781 260476
rect 116531 260132 116597 260133
rect 116531 260068 116532 260132
rect 116596 260068 116597 260132
rect 116531 260067 116597 260068
rect 115795 146300 115861 146301
rect 115795 146236 115796 146300
rect 115860 146236 115861 146300
rect 115795 146235 115861 146236
rect 115795 145620 115861 145621
rect 115795 145556 115796 145620
rect 115860 145556 115861 145620
rect 115795 145555 115861 145556
rect 115611 144804 115677 144805
rect 115611 144740 115612 144804
rect 115676 144740 115677 144804
rect 115611 144739 115677 144740
rect 115611 140316 115677 140317
rect 115611 140252 115612 140316
rect 115676 140252 115677 140316
rect 115611 140251 115677 140252
rect 115614 71501 115674 140251
rect 115611 71500 115677 71501
rect 115611 71436 115612 71500
rect 115676 71436 115677 71500
rect 115611 71435 115677 71436
rect 115798 66197 115858 145555
rect 116534 144805 116594 260067
rect 116531 144804 116597 144805
rect 116531 144740 116532 144804
rect 116596 144740 116597 144804
rect 116531 144739 116597 144740
rect 116718 143445 116778 260475
rect 116902 143853 116962 263739
rect 118794 262000 119414 263898
rect 123294 707718 123914 711590
rect 123294 707482 123326 707718
rect 123562 707482 123646 707718
rect 123882 707482 123914 707718
rect 123294 707398 123914 707482
rect 123294 707162 123326 707398
rect 123562 707162 123646 707398
rect 123882 707162 123914 707398
rect 123294 700954 123914 707162
rect 123294 700718 123326 700954
rect 123562 700718 123646 700954
rect 123882 700718 123914 700954
rect 123294 700634 123914 700718
rect 123294 700398 123326 700634
rect 123562 700398 123646 700634
rect 123882 700398 123914 700634
rect 123294 664954 123914 700398
rect 123294 664718 123326 664954
rect 123562 664718 123646 664954
rect 123882 664718 123914 664954
rect 123294 664634 123914 664718
rect 123294 664398 123326 664634
rect 123562 664398 123646 664634
rect 123882 664398 123914 664634
rect 123294 628954 123914 664398
rect 123294 628718 123326 628954
rect 123562 628718 123646 628954
rect 123882 628718 123914 628954
rect 123294 628634 123914 628718
rect 123294 628398 123326 628634
rect 123562 628398 123646 628634
rect 123882 628398 123914 628634
rect 123294 592954 123914 628398
rect 123294 592718 123326 592954
rect 123562 592718 123646 592954
rect 123882 592718 123914 592954
rect 123294 592634 123914 592718
rect 123294 592398 123326 592634
rect 123562 592398 123646 592634
rect 123882 592398 123914 592634
rect 123294 556954 123914 592398
rect 123294 556718 123326 556954
rect 123562 556718 123646 556954
rect 123882 556718 123914 556954
rect 123294 556634 123914 556718
rect 123294 556398 123326 556634
rect 123562 556398 123646 556634
rect 123882 556398 123914 556634
rect 123294 520954 123914 556398
rect 123294 520718 123326 520954
rect 123562 520718 123646 520954
rect 123882 520718 123914 520954
rect 123294 520634 123914 520718
rect 123294 520398 123326 520634
rect 123562 520398 123646 520634
rect 123882 520398 123914 520634
rect 123294 484954 123914 520398
rect 123294 484718 123326 484954
rect 123562 484718 123646 484954
rect 123882 484718 123914 484954
rect 123294 484634 123914 484718
rect 123294 484398 123326 484634
rect 123562 484398 123646 484634
rect 123882 484398 123914 484634
rect 123294 448954 123914 484398
rect 123294 448718 123326 448954
rect 123562 448718 123646 448954
rect 123882 448718 123914 448954
rect 123294 448634 123914 448718
rect 123294 448398 123326 448634
rect 123562 448398 123646 448634
rect 123882 448398 123914 448634
rect 123294 412954 123914 448398
rect 123294 412718 123326 412954
rect 123562 412718 123646 412954
rect 123882 412718 123914 412954
rect 123294 412634 123914 412718
rect 123294 412398 123326 412634
rect 123562 412398 123646 412634
rect 123882 412398 123914 412634
rect 123294 376954 123914 412398
rect 123294 376718 123326 376954
rect 123562 376718 123646 376954
rect 123882 376718 123914 376954
rect 123294 376634 123914 376718
rect 123294 376398 123326 376634
rect 123562 376398 123646 376634
rect 123882 376398 123914 376634
rect 123294 340954 123914 376398
rect 123294 340718 123326 340954
rect 123562 340718 123646 340954
rect 123882 340718 123914 340954
rect 123294 340634 123914 340718
rect 123294 340398 123326 340634
rect 123562 340398 123646 340634
rect 123882 340398 123914 340634
rect 123294 304954 123914 340398
rect 123294 304718 123326 304954
rect 123562 304718 123646 304954
rect 123882 304718 123914 304954
rect 123294 304634 123914 304718
rect 123294 304398 123326 304634
rect 123562 304398 123646 304634
rect 123882 304398 123914 304634
rect 123294 268954 123914 304398
rect 123294 268718 123326 268954
rect 123562 268718 123646 268954
rect 123882 268718 123914 268954
rect 123294 268634 123914 268718
rect 123294 268398 123326 268634
rect 123562 268398 123646 268634
rect 123882 268398 123914 268634
rect 123294 262000 123914 268398
rect 127794 708678 128414 711590
rect 127794 708442 127826 708678
rect 128062 708442 128146 708678
rect 128382 708442 128414 708678
rect 127794 708358 128414 708442
rect 127794 708122 127826 708358
rect 128062 708122 128146 708358
rect 128382 708122 128414 708358
rect 127794 669454 128414 708122
rect 127794 669218 127826 669454
rect 128062 669218 128146 669454
rect 128382 669218 128414 669454
rect 127794 669134 128414 669218
rect 127794 668898 127826 669134
rect 128062 668898 128146 669134
rect 128382 668898 128414 669134
rect 127794 633454 128414 668898
rect 127794 633218 127826 633454
rect 128062 633218 128146 633454
rect 128382 633218 128414 633454
rect 127794 633134 128414 633218
rect 127794 632898 127826 633134
rect 128062 632898 128146 633134
rect 128382 632898 128414 633134
rect 127794 597454 128414 632898
rect 127794 597218 127826 597454
rect 128062 597218 128146 597454
rect 128382 597218 128414 597454
rect 127794 597134 128414 597218
rect 127794 596898 127826 597134
rect 128062 596898 128146 597134
rect 128382 596898 128414 597134
rect 127794 561454 128414 596898
rect 127794 561218 127826 561454
rect 128062 561218 128146 561454
rect 128382 561218 128414 561454
rect 127794 561134 128414 561218
rect 127794 560898 127826 561134
rect 128062 560898 128146 561134
rect 128382 560898 128414 561134
rect 127794 525454 128414 560898
rect 127794 525218 127826 525454
rect 128062 525218 128146 525454
rect 128382 525218 128414 525454
rect 127794 525134 128414 525218
rect 127794 524898 127826 525134
rect 128062 524898 128146 525134
rect 128382 524898 128414 525134
rect 127794 489454 128414 524898
rect 127794 489218 127826 489454
rect 128062 489218 128146 489454
rect 128382 489218 128414 489454
rect 127794 489134 128414 489218
rect 127794 488898 127826 489134
rect 128062 488898 128146 489134
rect 128382 488898 128414 489134
rect 127794 453454 128414 488898
rect 127794 453218 127826 453454
rect 128062 453218 128146 453454
rect 128382 453218 128414 453454
rect 127794 453134 128414 453218
rect 127794 452898 127826 453134
rect 128062 452898 128146 453134
rect 128382 452898 128414 453134
rect 127794 417454 128414 452898
rect 127794 417218 127826 417454
rect 128062 417218 128146 417454
rect 128382 417218 128414 417454
rect 127794 417134 128414 417218
rect 127794 416898 127826 417134
rect 128062 416898 128146 417134
rect 128382 416898 128414 417134
rect 127794 381454 128414 416898
rect 127794 381218 127826 381454
rect 128062 381218 128146 381454
rect 128382 381218 128414 381454
rect 127794 381134 128414 381218
rect 127794 380898 127826 381134
rect 128062 380898 128146 381134
rect 128382 380898 128414 381134
rect 127794 345454 128414 380898
rect 127794 345218 127826 345454
rect 128062 345218 128146 345454
rect 128382 345218 128414 345454
rect 127794 345134 128414 345218
rect 127794 344898 127826 345134
rect 128062 344898 128146 345134
rect 128382 344898 128414 345134
rect 127794 309454 128414 344898
rect 127794 309218 127826 309454
rect 128062 309218 128146 309454
rect 128382 309218 128414 309454
rect 127794 309134 128414 309218
rect 127794 308898 127826 309134
rect 128062 308898 128146 309134
rect 128382 308898 128414 309134
rect 127794 273454 128414 308898
rect 127794 273218 127826 273454
rect 128062 273218 128146 273454
rect 128382 273218 128414 273454
rect 127794 273134 128414 273218
rect 127794 272898 127826 273134
rect 128062 272898 128146 273134
rect 128382 272898 128414 273134
rect 127794 262000 128414 272898
rect 132294 709638 132914 711590
rect 132294 709402 132326 709638
rect 132562 709402 132646 709638
rect 132882 709402 132914 709638
rect 132294 709318 132914 709402
rect 132294 709082 132326 709318
rect 132562 709082 132646 709318
rect 132882 709082 132914 709318
rect 132294 673954 132914 709082
rect 132294 673718 132326 673954
rect 132562 673718 132646 673954
rect 132882 673718 132914 673954
rect 132294 673634 132914 673718
rect 132294 673398 132326 673634
rect 132562 673398 132646 673634
rect 132882 673398 132914 673634
rect 132294 637954 132914 673398
rect 132294 637718 132326 637954
rect 132562 637718 132646 637954
rect 132882 637718 132914 637954
rect 132294 637634 132914 637718
rect 132294 637398 132326 637634
rect 132562 637398 132646 637634
rect 132882 637398 132914 637634
rect 132294 601954 132914 637398
rect 132294 601718 132326 601954
rect 132562 601718 132646 601954
rect 132882 601718 132914 601954
rect 132294 601634 132914 601718
rect 132294 601398 132326 601634
rect 132562 601398 132646 601634
rect 132882 601398 132914 601634
rect 132294 565954 132914 601398
rect 132294 565718 132326 565954
rect 132562 565718 132646 565954
rect 132882 565718 132914 565954
rect 132294 565634 132914 565718
rect 132294 565398 132326 565634
rect 132562 565398 132646 565634
rect 132882 565398 132914 565634
rect 132294 529954 132914 565398
rect 132294 529718 132326 529954
rect 132562 529718 132646 529954
rect 132882 529718 132914 529954
rect 132294 529634 132914 529718
rect 132294 529398 132326 529634
rect 132562 529398 132646 529634
rect 132882 529398 132914 529634
rect 132294 493954 132914 529398
rect 132294 493718 132326 493954
rect 132562 493718 132646 493954
rect 132882 493718 132914 493954
rect 132294 493634 132914 493718
rect 132294 493398 132326 493634
rect 132562 493398 132646 493634
rect 132882 493398 132914 493634
rect 132294 457954 132914 493398
rect 132294 457718 132326 457954
rect 132562 457718 132646 457954
rect 132882 457718 132914 457954
rect 132294 457634 132914 457718
rect 132294 457398 132326 457634
rect 132562 457398 132646 457634
rect 132882 457398 132914 457634
rect 132294 421954 132914 457398
rect 132294 421718 132326 421954
rect 132562 421718 132646 421954
rect 132882 421718 132914 421954
rect 132294 421634 132914 421718
rect 132294 421398 132326 421634
rect 132562 421398 132646 421634
rect 132882 421398 132914 421634
rect 132294 385954 132914 421398
rect 132294 385718 132326 385954
rect 132562 385718 132646 385954
rect 132882 385718 132914 385954
rect 132294 385634 132914 385718
rect 132294 385398 132326 385634
rect 132562 385398 132646 385634
rect 132882 385398 132914 385634
rect 132294 349954 132914 385398
rect 132294 349718 132326 349954
rect 132562 349718 132646 349954
rect 132882 349718 132914 349954
rect 132294 349634 132914 349718
rect 132294 349398 132326 349634
rect 132562 349398 132646 349634
rect 132882 349398 132914 349634
rect 132294 313954 132914 349398
rect 132294 313718 132326 313954
rect 132562 313718 132646 313954
rect 132882 313718 132914 313954
rect 132294 313634 132914 313718
rect 132294 313398 132326 313634
rect 132562 313398 132646 313634
rect 132882 313398 132914 313634
rect 132294 277954 132914 313398
rect 132294 277718 132326 277954
rect 132562 277718 132646 277954
rect 132882 277718 132914 277954
rect 132294 277634 132914 277718
rect 132294 277398 132326 277634
rect 132562 277398 132646 277634
rect 132882 277398 132914 277634
rect 132294 262000 132914 277398
rect 136794 710598 137414 711590
rect 136794 710362 136826 710598
rect 137062 710362 137146 710598
rect 137382 710362 137414 710598
rect 136794 710278 137414 710362
rect 136794 710042 136826 710278
rect 137062 710042 137146 710278
rect 137382 710042 137414 710278
rect 136794 678454 137414 710042
rect 136794 678218 136826 678454
rect 137062 678218 137146 678454
rect 137382 678218 137414 678454
rect 136794 678134 137414 678218
rect 136794 677898 136826 678134
rect 137062 677898 137146 678134
rect 137382 677898 137414 678134
rect 136794 642454 137414 677898
rect 136794 642218 136826 642454
rect 137062 642218 137146 642454
rect 137382 642218 137414 642454
rect 136794 642134 137414 642218
rect 136794 641898 136826 642134
rect 137062 641898 137146 642134
rect 137382 641898 137414 642134
rect 136794 606454 137414 641898
rect 136794 606218 136826 606454
rect 137062 606218 137146 606454
rect 137382 606218 137414 606454
rect 136794 606134 137414 606218
rect 136794 605898 136826 606134
rect 137062 605898 137146 606134
rect 137382 605898 137414 606134
rect 136794 570454 137414 605898
rect 136794 570218 136826 570454
rect 137062 570218 137146 570454
rect 137382 570218 137414 570454
rect 136794 570134 137414 570218
rect 136794 569898 136826 570134
rect 137062 569898 137146 570134
rect 137382 569898 137414 570134
rect 136794 534454 137414 569898
rect 136794 534218 136826 534454
rect 137062 534218 137146 534454
rect 137382 534218 137414 534454
rect 136794 534134 137414 534218
rect 136794 533898 136826 534134
rect 137062 533898 137146 534134
rect 137382 533898 137414 534134
rect 136794 498454 137414 533898
rect 136794 498218 136826 498454
rect 137062 498218 137146 498454
rect 137382 498218 137414 498454
rect 136794 498134 137414 498218
rect 136794 497898 136826 498134
rect 137062 497898 137146 498134
rect 137382 497898 137414 498134
rect 136794 462454 137414 497898
rect 136794 462218 136826 462454
rect 137062 462218 137146 462454
rect 137382 462218 137414 462454
rect 136794 462134 137414 462218
rect 136794 461898 136826 462134
rect 137062 461898 137146 462134
rect 137382 461898 137414 462134
rect 136794 426454 137414 461898
rect 136794 426218 136826 426454
rect 137062 426218 137146 426454
rect 137382 426218 137414 426454
rect 136794 426134 137414 426218
rect 136794 425898 136826 426134
rect 137062 425898 137146 426134
rect 137382 425898 137414 426134
rect 136794 390454 137414 425898
rect 136794 390218 136826 390454
rect 137062 390218 137146 390454
rect 137382 390218 137414 390454
rect 136794 390134 137414 390218
rect 136794 389898 136826 390134
rect 137062 389898 137146 390134
rect 137382 389898 137414 390134
rect 136794 354454 137414 389898
rect 136794 354218 136826 354454
rect 137062 354218 137146 354454
rect 137382 354218 137414 354454
rect 136794 354134 137414 354218
rect 136794 353898 136826 354134
rect 137062 353898 137146 354134
rect 137382 353898 137414 354134
rect 136794 318454 137414 353898
rect 136794 318218 136826 318454
rect 137062 318218 137146 318454
rect 137382 318218 137414 318454
rect 136794 318134 137414 318218
rect 136794 317898 136826 318134
rect 137062 317898 137146 318134
rect 137382 317898 137414 318134
rect 136794 282454 137414 317898
rect 136794 282218 136826 282454
rect 137062 282218 137146 282454
rect 137382 282218 137414 282454
rect 136794 282134 137414 282218
rect 136794 281898 136826 282134
rect 137062 281898 137146 282134
rect 137382 281898 137414 282134
rect 136794 262000 137414 281898
rect 141294 711558 141914 711590
rect 141294 711322 141326 711558
rect 141562 711322 141646 711558
rect 141882 711322 141914 711558
rect 141294 711238 141914 711322
rect 141294 711002 141326 711238
rect 141562 711002 141646 711238
rect 141882 711002 141914 711238
rect 141294 682954 141914 711002
rect 141294 682718 141326 682954
rect 141562 682718 141646 682954
rect 141882 682718 141914 682954
rect 141294 682634 141914 682718
rect 141294 682398 141326 682634
rect 141562 682398 141646 682634
rect 141882 682398 141914 682634
rect 141294 646954 141914 682398
rect 141294 646718 141326 646954
rect 141562 646718 141646 646954
rect 141882 646718 141914 646954
rect 141294 646634 141914 646718
rect 141294 646398 141326 646634
rect 141562 646398 141646 646634
rect 141882 646398 141914 646634
rect 141294 610954 141914 646398
rect 141294 610718 141326 610954
rect 141562 610718 141646 610954
rect 141882 610718 141914 610954
rect 141294 610634 141914 610718
rect 141294 610398 141326 610634
rect 141562 610398 141646 610634
rect 141882 610398 141914 610634
rect 141294 574954 141914 610398
rect 141294 574718 141326 574954
rect 141562 574718 141646 574954
rect 141882 574718 141914 574954
rect 141294 574634 141914 574718
rect 141294 574398 141326 574634
rect 141562 574398 141646 574634
rect 141882 574398 141914 574634
rect 141294 538954 141914 574398
rect 141294 538718 141326 538954
rect 141562 538718 141646 538954
rect 141882 538718 141914 538954
rect 141294 538634 141914 538718
rect 141294 538398 141326 538634
rect 141562 538398 141646 538634
rect 141882 538398 141914 538634
rect 141294 502954 141914 538398
rect 141294 502718 141326 502954
rect 141562 502718 141646 502954
rect 141882 502718 141914 502954
rect 141294 502634 141914 502718
rect 141294 502398 141326 502634
rect 141562 502398 141646 502634
rect 141882 502398 141914 502634
rect 141294 466954 141914 502398
rect 141294 466718 141326 466954
rect 141562 466718 141646 466954
rect 141882 466718 141914 466954
rect 141294 466634 141914 466718
rect 141294 466398 141326 466634
rect 141562 466398 141646 466634
rect 141882 466398 141914 466634
rect 141294 430954 141914 466398
rect 141294 430718 141326 430954
rect 141562 430718 141646 430954
rect 141882 430718 141914 430954
rect 141294 430634 141914 430718
rect 141294 430398 141326 430634
rect 141562 430398 141646 430634
rect 141882 430398 141914 430634
rect 141294 394954 141914 430398
rect 141294 394718 141326 394954
rect 141562 394718 141646 394954
rect 141882 394718 141914 394954
rect 141294 394634 141914 394718
rect 141294 394398 141326 394634
rect 141562 394398 141646 394634
rect 141882 394398 141914 394634
rect 141294 358954 141914 394398
rect 141294 358718 141326 358954
rect 141562 358718 141646 358954
rect 141882 358718 141914 358954
rect 141294 358634 141914 358718
rect 141294 358398 141326 358634
rect 141562 358398 141646 358634
rect 141882 358398 141914 358634
rect 141294 322954 141914 358398
rect 141294 322718 141326 322954
rect 141562 322718 141646 322954
rect 141882 322718 141914 322954
rect 141294 322634 141914 322718
rect 141294 322398 141326 322634
rect 141562 322398 141646 322634
rect 141882 322398 141914 322634
rect 141294 286954 141914 322398
rect 141294 286718 141326 286954
rect 141562 286718 141646 286954
rect 141882 286718 141914 286954
rect 141294 286634 141914 286718
rect 141294 286398 141326 286634
rect 141562 286398 141646 286634
rect 141882 286398 141914 286634
rect 141294 262000 141914 286398
rect 145794 704838 146414 711590
rect 145794 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 146414 704838
rect 145794 704518 146414 704602
rect 145794 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 146414 704518
rect 145794 687454 146414 704282
rect 145794 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 146414 687454
rect 145794 687134 146414 687218
rect 145794 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 146414 687134
rect 145794 651454 146414 686898
rect 145794 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 146414 651454
rect 145794 651134 146414 651218
rect 145794 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 146414 651134
rect 145794 615454 146414 650898
rect 145794 615218 145826 615454
rect 146062 615218 146146 615454
rect 146382 615218 146414 615454
rect 145794 615134 146414 615218
rect 145794 614898 145826 615134
rect 146062 614898 146146 615134
rect 146382 614898 146414 615134
rect 145794 579454 146414 614898
rect 145794 579218 145826 579454
rect 146062 579218 146146 579454
rect 146382 579218 146414 579454
rect 145794 579134 146414 579218
rect 145794 578898 145826 579134
rect 146062 578898 146146 579134
rect 146382 578898 146414 579134
rect 145794 543454 146414 578898
rect 145794 543218 145826 543454
rect 146062 543218 146146 543454
rect 146382 543218 146414 543454
rect 145794 543134 146414 543218
rect 145794 542898 145826 543134
rect 146062 542898 146146 543134
rect 146382 542898 146414 543134
rect 145794 507454 146414 542898
rect 145794 507218 145826 507454
rect 146062 507218 146146 507454
rect 146382 507218 146414 507454
rect 145794 507134 146414 507218
rect 145794 506898 145826 507134
rect 146062 506898 146146 507134
rect 146382 506898 146414 507134
rect 145794 471454 146414 506898
rect 145794 471218 145826 471454
rect 146062 471218 146146 471454
rect 146382 471218 146414 471454
rect 145794 471134 146414 471218
rect 145794 470898 145826 471134
rect 146062 470898 146146 471134
rect 146382 470898 146414 471134
rect 145794 435454 146414 470898
rect 145794 435218 145826 435454
rect 146062 435218 146146 435454
rect 146382 435218 146414 435454
rect 145794 435134 146414 435218
rect 145794 434898 145826 435134
rect 146062 434898 146146 435134
rect 146382 434898 146414 435134
rect 145794 399454 146414 434898
rect 145794 399218 145826 399454
rect 146062 399218 146146 399454
rect 146382 399218 146414 399454
rect 145794 399134 146414 399218
rect 145794 398898 145826 399134
rect 146062 398898 146146 399134
rect 146382 398898 146414 399134
rect 145794 363454 146414 398898
rect 145794 363218 145826 363454
rect 146062 363218 146146 363454
rect 146382 363218 146414 363454
rect 145794 363134 146414 363218
rect 145794 362898 145826 363134
rect 146062 362898 146146 363134
rect 146382 362898 146414 363134
rect 145794 327454 146414 362898
rect 145794 327218 145826 327454
rect 146062 327218 146146 327454
rect 146382 327218 146414 327454
rect 145794 327134 146414 327218
rect 145794 326898 145826 327134
rect 146062 326898 146146 327134
rect 146382 326898 146414 327134
rect 145794 291454 146414 326898
rect 145794 291218 145826 291454
rect 146062 291218 146146 291454
rect 146382 291218 146414 291454
rect 145794 291134 146414 291218
rect 145794 290898 145826 291134
rect 146062 290898 146146 291134
rect 146382 290898 146414 291134
rect 145794 262000 146414 290898
rect 150294 705798 150914 711590
rect 150294 705562 150326 705798
rect 150562 705562 150646 705798
rect 150882 705562 150914 705798
rect 150294 705478 150914 705562
rect 150294 705242 150326 705478
rect 150562 705242 150646 705478
rect 150882 705242 150914 705478
rect 150294 691954 150914 705242
rect 150294 691718 150326 691954
rect 150562 691718 150646 691954
rect 150882 691718 150914 691954
rect 150294 691634 150914 691718
rect 150294 691398 150326 691634
rect 150562 691398 150646 691634
rect 150882 691398 150914 691634
rect 150294 655954 150914 691398
rect 150294 655718 150326 655954
rect 150562 655718 150646 655954
rect 150882 655718 150914 655954
rect 150294 655634 150914 655718
rect 150294 655398 150326 655634
rect 150562 655398 150646 655634
rect 150882 655398 150914 655634
rect 150294 619954 150914 655398
rect 150294 619718 150326 619954
rect 150562 619718 150646 619954
rect 150882 619718 150914 619954
rect 150294 619634 150914 619718
rect 150294 619398 150326 619634
rect 150562 619398 150646 619634
rect 150882 619398 150914 619634
rect 150294 583954 150914 619398
rect 150294 583718 150326 583954
rect 150562 583718 150646 583954
rect 150882 583718 150914 583954
rect 150294 583634 150914 583718
rect 150294 583398 150326 583634
rect 150562 583398 150646 583634
rect 150882 583398 150914 583634
rect 150294 547954 150914 583398
rect 150294 547718 150326 547954
rect 150562 547718 150646 547954
rect 150882 547718 150914 547954
rect 150294 547634 150914 547718
rect 150294 547398 150326 547634
rect 150562 547398 150646 547634
rect 150882 547398 150914 547634
rect 150294 511954 150914 547398
rect 150294 511718 150326 511954
rect 150562 511718 150646 511954
rect 150882 511718 150914 511954
rect 150294 511634 150914 511718
rect 150294 511398 150326 511634
rect 150562 511398 150646 511634
rect 150882 511398 150914 511634
rect 150294 475954 150914 511398
rect 150294 475718 150326 475954
rect 150562 475718 150646 475954
rect 150882 475718 150914 475954
rect 150294 475634 150914 475718
rect 150294 475398 150326 475634
rect 150562 475398 150646 475634
rect 150882 475398 150914 475634
rect 150294 439954 150914 475398
rect 150294 439718 150326 439954
rect 150562 439718 150646 439954
rect 150882 439718 150914 439954
rect 150294 439634 150914 439718
rect 150294 439398 150326 439634
rect 150562 439398 150646 439634
rect 150882 439398 150914 439634
rect 150294 403954 150914 439398
rect 150294 403718 150326 403954
rect 150562 403718 150646 403954
rect 150882 403718 150914 403954
rect 150294 403634 150914 403718
rect 150294 403398 150326 403634
rect 150562 403398 150646 403634
rect 150882 403398 150914 403634
rect 150294 367954 150914 403398
rect 150294 367718 150326 367954
rect 150562 367718 150646 367954
rect 150882 367718 150914 367954
rect 150294 367634 150914 367718
rect 150294 367398 150326 367634
rect 150562 367398 150646 367634
rect 150882 367398 150914 367634
rect 150294 331954 150914 367398
rect 150294 331718 150326 331954
rect 150562 331718 150646 331954
rect 150882 331718 150914 331954
rect 150294 331634 150914 331718
rect 150294 331398 150326 331634
rect 150562 331398 150646 331634
rect 150882 331398 150914 331634
rect 150294 295954 150914 331398
rect 150294 295718 150326 295954
rect 150562 295718 150646 295954
rect 150882 295718 150914 295954
rect 150294 295634 150914 295718
rect 150294 295398 150326 295634
rect 150562 295398 150646 295634
rect 150882 295398 150914 295634
rect 150294 262000 150914 295398
rect 154794 706758 155414 711590
rect 154794 706522 154826 706758
rect 155062 706522 155146 706758
rect 155382 706522 155414 706758
rect 154794 706438 155414 706522
rect 154794 706202 154826 706438
rect 155062 706202 155146 706438
rect 155382 706202 155414 706438
rect 154794 696454 155414 706202
rect 154794 696218 154826 696454
rect 155062 696218 155146 696454
rect 155382 696218 155414 696454
rect 154794 696134 155414 696218
rect 154794 695898 154826 696134
rect 155062 695898 155146 696134
rect 155382 695898 155414 696134
rect 154794 660454 155414 695898
rect 154794 660218 154826 660454
rect 155062 660218 155146 660454
rect 155382 660218 155414 660454
rect 154794 660134 155414 660218
rect 154794 659898 154826 660134
rect 155062 659898 155146 660134
rect 155382 659898 155414 660134
rect 154794 624454 155414 659898
rect 154794 624218 154826 624454
rect 155062 624218 155146 624454
rect 155382 624218 155414 624454
rect 154794 624134 155414 624218
rect 154794 623898 154826 624134
rect 155062 623898 155146 624134
rect 155382 623898 155414 624134
rect 154794 588454 155414 623898
rect 154794 588218 154826 588454
rect 155062 588218 155146 588454
rect 155382 588218 155414 588454
rect 154794 588134 155414 588218
rect 154794 587898 154826 588134
rect 155062 587898 155146 588134
rect 155382 587898 155414 588134
rect 154794 552454 155414 587898
rect 154794 552218 154826 552454
rect 155062 552218 155146 552454
rect 155382 552218 155414 552454
rect 154794 552134 155414 552218
rect 154794 551898 154826 552134
rect 155062 551898 155146 552134
rect 155382 551898 155414 552134
rect 154794 516454 155414 551898
rect 154794 516218 154826 516454
rect 155062 516218 155146 516454
rect 155382 516218 155414 516454
rect 154794 516134 155414 516218
rect 154794 515898 154826 516134
rect 155062 515898 155146 516134
rect 155382 515898 155414 516134
rect 154794 480454 155414 515898
rect 154794 480218 154826 480454
rect 155062 480218 155146 480454
rect 155382 480218 155414 480454
rect 154794 480134 155414 480218
rect 154794 479898 154826 480134
rect 155062 479898 155146 480134
rect 155382 479898 155414 480134
rect 154794 444454 155414 479898
rect 154794 444218 154826 444454
rect 155062 444218 155146 444454
rect 155382 444218 155414 444454
rect 154794 444134 155414 444218
rect 154794 443898 154826 444134
rect 155062 443898 155146 444134
rect 155382 443898 155414 444134
rect 154794 408454 155414 443898
rect 154794 408218 154826 408454
rect 155062 408218 155146 408454
rect 155382 408218 155414 408454
rect 154794 408134 155414 408218
rect 154794 407898 154826 408134
rect 155062 407898 155146 408134
rect 155382 407898 155414 408134
rect 154794 372454 155414 407898
rect 154794 372218 154826 372454
rect 155062 372218 155146 372454
rect 155382 372218 155414 372454
rect 154794 372134 155414 372218
rect 154794 371898 154826 372134
rect 155062 371898 155146 372134
rect 155382 371898 155414 372134
rect 154794 336454 155414 371898
rect 154794 336218 154826 336454
rect 155062 336218 155146 336454
rect 155382 336218 155414 336454
rect 154794 336134 155414 336218
rect 154794 335898 154826 336134
rect 155062 335898 155146 336134
rect 155382 335898 155414 336134
rect 154794 300454 155414 335898
rect 154794 300218 154826 300454
rect 155062 300218 155146 300454
rect 155382 300218 155414 300454
rect 154794 300134 155414 300218
rect 154794 299898 154826 300134
rect 155062 299898 155146 300134
rect 155382 299898 155414 300134
rect 154794 264454 155414 299898
rect 154794 264218 154826 264454
rect 155062 264218 155146 264454
rect 155382 264218 155414 264454
rect 154794 264134 155414 264218
rect 154794 263898 154826 264134
rect 155062 263898 155146 264134
rect 155382 263898 155414 264134
rect 154794 262000 155414 263898
rect 159294 707718 159914 711590
rect 159294 707482 159326 707718
rect 159562 707482 159646 707718
rect 159882 707482 159914 707718
rect 159294 707398 159914 707482
rect 159294 707162 159326 707398
rect 159562 707162 159646 707398
rect 159882 707162 159914 707398
rect 159294 700954 159914 707162
rect 159294 700718 159326 700954
rect 159562 700718 159646 700954
rect 159882 700718 159914 700954
rect 159294 700634 159914 700718
rect 159294 700398 159326 700634
rect 159562 700398 159646 700634
rect 159882 700398 159914 700634
rect 159294 664954 159914 700398
rect 159294 664718 159326 664954
rect 159562 664718 159646 664954
rect 159882 664718 159914 664954
rect 159294 664634 159914 664718
rect 159294 664398 159326 664634
rect 159562 664398 159646 664634
rect 159882 664398 159914 664634
rect 159294 628954 159914 664398
rect 159294 628718 159326 628954
rect 159562 628718 159646 628954
rect 159882 628718 159914 628954
rect 159294 628634 159914 628718
rect 159294 628398 159326 628634
rect 159562 628398 159646 628634
rect 159882 628398 159914 628634
rect 159294 592954 159914 628398
rect 159294 592718 159326 592954
rect 159562 592718 159646 592954
rect 159882 592718 159914 592954
rect 159294 592634 159914 592718
rect 159294 592398 159326 592634
rect 159562 592398 159646 592634
rect 159882 592398 159914 592634
rect 159294 556954 159914 592398
rect 159294 556718 159326 556954
rect 159562 556718 159646 556954
rect 159882 556718 159914 556954
rect 159294 556634 159914 556718
rect 159294 556398 159326 556634
rect 159562 556398 159646 556634
rect 159882 556398 159914 556634
rect 159294 520954 159914 556398
rect 159294 520718 159326 520954
rect 159562 520718 159646 520954
rect 159882 520718 159914 520954
rect 159294 520634 159914 520718
rect 159294 520398 159326 520634
rect 159562 520398 159646 520634
rect 159882 520398 159914 520634
rect 159294 484954 159914 520398
rect 159294 484718 159326 484954
rect 159562 484718 159646 484954
rect 159882 484718 159914 484954
rect 159294 484634 159914 484718
rect 159294 484398 159326 484634
rect 159562 484398 159646 484634
rect 159882 484398 159914 484634
rect 159294 448954 159914 484398
rect 159294 448718 159326 448954
rect 159562 448718 159646 448954
rect 159882 448718 159914 448954
rect 159294 448634 159914 448718
rect 159294 448398 159326 448634
rect 159562 448398 159646 448634
rect 159882 448398 159914 448634
rect 159294 412954 159914 448398
rect 159294 412718 159326 412954
rect 159562 412718 159646 412954
rect 159882 412718 159914 412954
rect 159294 412634 159914 412718
rect 159294 412398 159326 412634
rect 159562 412398 159646 412634
rect 159882 412398 159914 412634
rect 159294 376954 159914 412398
rect 159294 376718 159326 376954
rect 159562 376718 159646 376954
rect 159882 376718 159914 376954
rect 159294 376634 159914 376718
rect 159294 376398 159326 376634
rect 159562 376398 159646 376634
rect 159882 376398 159914 376634
rect 159294 340954 159914 376398
rect 159294 340718 159326 340954
rect 159562 340718 159646 340954
rect 159882 340718 159914 340954
rect 159294 340634 159914 340718
rect 159294 340398 159326 340634
rect 159562 340398 159646 340634
rect 159882 340398 159914 340634
rect 159294 304954 159914 340398
rect 159294 304718 159326 304954
rect 159562 304718 159646 304954
rect 159882 304718 159914 304954
rect 159294 304634 159914 304718
rect 159294 304398 159326 304634
rect 159562 304398 159646 304634
rect 159882 304398 159914 304634
rect 159294 268954 159914 304398
rect 159294 268718 159326 268954
rect 159562 268718 159646 268954
rect 159882 268718 159914 268954
rect 159294 268634 159914 268718
rect 159294 268398 159326 268634
rect 159562 268398 159646 268634
rect 159882 268398 159914 268634
rect 159294 262000 159914 268398
rect 163794 708678 164414 711590
rect 163794 708442 163826 708678
rect 164062 708442 164146 708678
rect 164382 708442 164414 708678
rect 163794 708358 164414 708442
rect 163794 708122 163826 708358
rect 164062 708122 164146 708358
rect 164382 708122 164414 708358
rect 163794 669454 164414 708122
rect 163794 669218 163826 669454
rect 164062 669218 164146 669454
rect 164382 669218 164414 669454
rect 163794 669134 164414 669218
rect 163794 668898 163826 669134
rect 164062 668898 164146 669134
rect 164382 668898 164414 669134
rect 163794 633454 164414 668898
rect 163794 633218 163826 633454
rect 164062 633218 164146 633454
rect 164382 633218 164414 633454
rect 163794 633134 164414 633218
rect 163794 632898 163826 633134
rect 164062 632898 164146 633134
rect 164382 632898 164414 633134
rect 163794 597454 164414 632898
rect 163794 597218 163826 597454
rect 164062 597218 164146 597454
rect 164382 597218 164414 597454
rect 163794 597134 164414 597218
rect 163794 596898 163826 597134
rect 164062 596898 164146 597134
rect 164382 596898 164414 597134
rect 163794 561454 164414 596898
rect 163794 561218 163826 561454
rect 164062 561218 164146 561454
rect 164382 561218 164414 561454
rect 163794 561134 164414 561218
rect 163794 560898 163826 561134
rect 164062 560898 164146 561134
rect 164382 560898 164414 561134
rect 163794 525454 164414 560898
rect 163794 525218 163826 525454
rect 164062 525218 164146 525454
rect 164382 525218 164414 525454
rect 163794 525134 164414 525218
rect 163794 524898 163826 525134
rect 164062 524898 164146 525134
rect 164382 524898 164414 525134
rect 163794 489454 164414 524898
rect 163794 489218 163826 489454
rect 164062 489218 164146 489454
rect 164382 489218 164414 489454
rect 163794 489134 164414 489218
rect 163794 488898 163826 489134
rect 164062 488898 164146 489134
rect 164382 488898 164414 489134
rect 163794 453454 164414 488898
rect 163794 453218 163826 453454
rect 164062 453218 164146 453454
rect 164382 453218 164414 453454
rect 163794 453134 164414 453218
rect 163794 452898 163826 453134
rect 164062 452898 164146 453134
rect 164382 452898 164414 453134
rect 163794 417454 164414 452898
rect 163794 417218 163826 417454
rect 164062 417218 164146 417454
rect 164382 417218 164414 417454
rect 163794 417134 164414 417218
rect 163794 416898 163826 417134
rect 164062 416898 164146 417134
rect 164382 416898 164414 417134
rect 163794 381454 164414 416898
rect 163794 381218 163826 381454
rect 164062 381218 164146 381454
rect 164382 381218 164414 381454
rect 163794 381134 164414 381218
rect 163794 380898 163826 381134
rect 164062 380898 164146 381134
rect 164382 380898 164414 381134
rect 163794 345454 164414 380898
rect 163794 345218 163826 345454
rect 164062 345218 164146 345454
rect 164382 345218 164414 345454
rect 163794 345134 164414 345218
rect 163794 344898 163826 345134
rect 164062 344898 164146 345134
rect 164382 344898 164414 345134
rect 163794 309454 164414 344898
rect 163794 309218 163826 309454
rect 164062 309218 164146 309454
rect 164382 309218 164414 309454
rect 163794 309134 164414 309218
rect 163794 308898 163826 309134
rect 164062 308898 164146 309134
rect 164382 308898 164414 309134
rect 163794 273454 164414 308898
rect 163794 273218 163826 273454
rect 164062 273218 164146 273454
rect 164382 273218 164414 273454
rect 163794 273134 164414 273218
rect 163794 272898 163826 273134
rect 164062 272898 164146 273134
rect 164382 272898 164414 273134
rect 163794 262000 164414 272898
rect 168294 709638 168914 711590
rect 168294 709402 168326 709638
rect 168562 709402 168646 709638
rect 168882 709402 168914 709638
rect 168294 709318 168914 709402
rect 168294 709082 168326 709318
rect 168562 709082 168646 709318
rect 168882 709082 168914 709318
rect 168294 673954 168914 709082
rect 168294 673718 168326 673954
rect 168562 673718 168646 673954
rect 168882 673718 168914 673954
rect 168294 673634 168914 673718
rect 168294 673398 168326 673634
rect 168562 673398 168646 673634
rect 168882 673398 168914 673634
rect 168294 637954 168914 673398
rect 168294 637718 168326 637954
rect 168562 637718 168646 637954
rect 168882 637718 168914 637954
rect 168294 637634 168914 637718
rect 168294 637398 168326 637634
rect 168562 637398 168646 637634
rect 168882 637398 168914 637634
rect 168294 601954 168914 637398
rect 168294 601718 168326 601954
rect 168562 601718 168646 601954
rect 168882 601718 168914 601954
rect 168294 601634 168914 601718
rect 168294 601398 168326 601634
rect 168562 601398 168646 601634
rect 168882 601398 168914 601634
rect 168294 565954 168914 601398
rect 168294 565718 168326 565954
rect 168562 565718 168646 565954
rect 168882 565718 168914 565954
rect 168294 565634 168914 565718
rect 168294 565398 168326 565634
rect 168562 565398 168646 565634
rect 168882 565398 168914 565634
rect 168294 529954 168914 565398
rect 168294 529718 168326 529954
rect 168562 529718 168646 529954
rect 168882 529718 168914 529954
rect 168294 529634 168914 529718
rect 168294 529398 168326 529634
rect 168562 529398 168646 529634
rect 168882 529398 168914 529634
rect 168294 493954 168914 529398
rect 168294 493718 168326 493954
rect 168562 493718 168646 493954
rect 168882 493718 168914 493954
rect 168294 493634 168914 493718
rect 168294 493398 168326 493634
rect 168562 493398 168646 493634
rect 168882 493398 168914 493634
rect 168294 457954 168914 493398
rect 168294 457718 168326 457954
rect 168562 457718 168646 457954
rect 168882 457718 168914 457954
rect 168294 457634 168914 457718
rect 168294 457398 168326 457634
rect 168562 457398 168646 457634
rect 168882 457398 168914 457634
rect 168294 421954 168914 457398
rect 168294 421718 168326 421954
rect 168562 421718 168646 421954
rect 168882 421718 168914 421954
rect 168294 421634 168914 421718
rect 168294 421398 168326 421634
rect 168562 421398 168646 421634
rect 168882 421398 168914 421634
rect 168294 385954 168914 421398
rect 168294 385718 168326 385954
rect 168562 385718 168646 385954
rect 168882 385718 168914 385954
rect 168294 385634 168914 385718
rect 168294 385398 168326 385634
rect 168562 385398 168646 385634
rect 168882 385398 168914 385634
rect 168294 349954 168914 385398
rect 168294 349718 168326 349954
rect 168562 349718 168646 349954
rect 168882 349718 168914 349954
rect 168294 349634 168914 349718
rect 168294 349398 168326 349634
rect 168562 349398 168646 349634
rect 168882 349398 168914 349634
rect 168294 313954 168914 349398
rect 168294 313718 168326 313954
rect 168562 313718 168646 313954
rect 168882 313718 168914 313954
rect 168294 313634 168914 313718
rect 168294 313398 168326 313634
rect 168562 313398 168646 313634
rect 168882 313398 168914 313634
rect 168294 277954 168914 313398
rect 168294 277718 168326 277954
rect 168562 277718 168646 277954
rect 168882 277718 168914 277954
rect 168294 277634 168914 277718
rect 168294 277398 168326 277634
rect 168562 277398 168646 277634
rect 168882 277398 168914 277634
rect 168294 262000 168914 277398
rect 172794 710598 173414 711590
rect 172794 710362 172826 710598
rect 173062 710362 173146 710598
rect 173382 710362 173414 710598
rect 172794 710278 173414 710362
rect 172794 710042 172826 710278
rect 173062 710042 173146 710278
rect 173382 710042 173414 710278
rect 172794 678454 173414 710042
rect 172794 678218 172826 678454
rect 173062 678218 173146 678454
rect 173382 678218 173414 678454
rect 172794 678134 173414 678218
rect 172794 677898 172826 678134
rect 173062 677898 173146 678134
rect 173382 677898 173414 678134
rect 172794 642454 173414 677898
rect 172794 642218 172826 642454
rect 173062 642218 173146 642454
rect 173382 642218 173414 642454
rect 172794 642134 173414 642218
rect 172794 641898 172826 642134
rect 173062 641898 173146 642134
rect 173382 641898 173414 642134
rect 172794 606454 173414 641898
rect 172794 606218 172826 606454
rect 173062 606218 173146 606454
rect 173382 606218 173414 606454
rect 172794 606134 173414 606218
rect 172794 605898 172826 606134
rect 173062 605898 173146 606134
rect 173382 605898 173414 606134
rect 172794 570454 173414 605898
rect 172794 570218 172826 570454
rect 173062 570218 173146 570454
rect 173382 570218 173414 570454
rect 172794 570134 173414 570218
rect 172794 569898 172826 570134
rect 173062 569898 173146 570134
rect 173382 569898 173414 570134
rect 172794 534454 173414 569898
rect 172794 534218 172826 534454
rect 173062 534218 173146 534454
rect 173382 534218 173414 534454
rect 172794 534134 173414 534218
rect 172794 533898 172826 534134
rect 173062 533898 173146 534134
rect 173382 533898 173414 534134
rect 172794 498454 173414 533898
rect 172794 498218 172826 498454
rect 173062 498218 173146 498454
rect 173382 498218 173414 498454
rect 172794 498134 173414 498218
rect 172794 497898 172826 498134
rect 173062 497898 173146 498134
rect 173382 497898 173414 498134
rect 172794 462454 173414 497898
rect 172794 462218 172826 462454
rect 173062 462218 173146 462454
rect 173382 462218 173414 462454
rect 172794 462134 173414 462218
rect 172794 461898 172826 462134
rect 173062 461898 173146 462134
rect 173382 461898 173414 462134
rect 172794 426454 173414 461898
rect 172794 426218 172826 426454
rect 173062 426218 173146 426454
rect 173382 426218 173414 426454
rect 172794 426134 173414 426218
rect 172794 425898 172826 426134
rect 173062 425898 173146 426134
rect 173382 425898 173414 426134
rect 172794 390454 173414 425898
rect 172794 390218 172826 390454
rect 173062 390218 173146 390454
rect 173382 390218 173414 390454
rect 172794 390134 173414 390218
rect 172794 389898 172826 390134
rect 173062 389898 173146 390134
rect 173382 389898 173414 390134
rect 172794 354454 173414 389898
rect 172794 354218 172826 354454
rect 173062 354218 173146 354454
rect 173382 354218 173414 354454
rect 172794 354134 173414 354218
rect 172794 353898 172826 354134
rect 173062 353898 173146 354134
rect 173382 353898 173414 354134
rect 172794 318454 173414 353898
rect 172794 318218 172826 318454
rect 173062 318218 173146 318454
rect 173382 318218 173414 318454
rect 172794 318134 173414 318218
rect 172794 317898 172826 318134
rect 173062 317898 173146 318134
rect 173382 317898 173414 318134
rect 172794 282454 173414 317898
rect 172794 282218 172826 282454
rect 173062 282218 173146 282454
rect 173382 282218 173414 282454
rect 172794 282134 173414 282218
rect 172794 281898 172826 282134
rect 173062 281898 173146 282134
rect 173382 281898 173414 282134
rect 172794 262000 173414 281898
rect 177294 711558 177914 711590
rect 177294 711322 177326 711558
rect 177562 711322 177646 711558
rect 177882 711322 177914 711558
rect 177294 711238 177914 711322
rect 177294 711002 177326 711238
rect 177562 711002 177646 711238
rect 177882 711002 177914 711238
rect 177294 682954 177914 711002
rect 177294 682718 177326 682954
rect 177562 682718 177646 682954
rect 177882 682718 177914 682954
rect 177294 682634 177914 682718
rect 177294 682398 177326 682634
rect 177562 682398 177646 682634
rect 177882 682398 177914 682634
rect 177294 646954 177914 682398
rect 177294 646718 177326 646954
rect 177562 646718 177646 646954
rect 177882 646718 177914 646954
rect 177294 646634 177914 646718
rect 177294 646398 177326 646634
rect 177562 646398 177646 646634
rect 177882 646398 177914 646634
rect 177294 610954 177914 646398
rect 177294 610718 177326 610954
rect 177562 610718 177646 610954
rect 177882 610718 177914 610954
rect 177294 610634 177914 610718
rect 177294 610398 177326 610634
rect 177562 610398 177646 610634
rect 177882 610398 177914 610634
rect 177294 574954 177914 610398
rect 177294 574718 177326 574954
rect 177562 574718 177646 574954
rect 177882 574718 177914 574954
rect 177294 574634 177914 574718
rect 177294 574398 177326 574634
rect 177562 574398 177646 574634
rect 177882 574398 177914 574634
rect 177294 538954 177914 574398
rect 177294 538718 177326 538954
rect 177562 538718 177646 538954
rect 177882 538718 177914 538954
rect 177294 538634 177914 538718
rect 177294 538398 177326 538634
rect 177562 538398 177646 538634
rect 177882 538398 177914 538634
rect 177294 502954 177914 538398
rect 177294 502718 177326 502954
rect 177562 502718 177646 502954
rect 177882 502718 177914 502954
rect 177294 502634 177914 502718
rect 177294 502398 177326 502634
rect 177562 502398 177646 502634
rect 177882 502398 177914 502634
rect 177294 466954 177914 502398
rect 177294 466718 177326 466954
rect 177562 466718 177646 466954
rect 177882 466718 177914 466954
rect 177294 466634 177914 466718
rect 177294 466398 177326 466634
rect 177562 466398 177646 466634
rect 177882 466398 177914 466634
rect 177294 430954 177914 466398
rect 177294 430718 177326 430954
rect 177562 430718 177646 430954
rect 177882 430718 177914 430954
rect 177294 430634 177914 430718
rect 177294 430398 177326 430634
rect 177562 430398 177646 430634
rect 177882 430398 177914 430634
rect 177294 394954 177914 430398
rect 177294 394718 177326 394954
rect 177562 394718 177646 394954
rect 177882 394718 177914 394954
rect 177294 394634 177914 394718
rect 177294 394398 177326 394634
rect 177562 394398 177646 394634
rect 177882 394398 177914 394634
rect 177294 358954 177914 394398
rect 177294 358718 177326 358954
rect 177562 358718 177646 358954
rect 177882 358718 177914 358954
rect 177294 358634 177914 358718
rect 177294 358398 177326 358634
rect 177562 358398 177646 358634
rect 177882 358398 177914 358634
rect 177294 322954 177914 358398
rect 177294 322718 177326 322954
rect 177562 322718 177646 322954
rect 177882 322718 177914 322954
rect 177294 322634 177914 322718
rect 177294 322398 177326 322634
rect 177562 322398 177646 322634
rect 177882 322398 177914 322634
rect 177294 286954 177914 322398
rect 177294 286718 177326 286954
rect 177562 286718 177646 286954
rect 177882 286718 177914 286954
rect 177294 286634 177914 286718
rect 177294 286398 177326 286634
rect 177562 286398 177646 286634
rect 177882 286398 177914 286634
rect 177294 262000 177914 286398
rect 181794 704838 182414 711590
rect 181794 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 182414 704838
rect 181794 704518 182414 704602
rect 181794 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 182414 704518
rect 181794 687454 182414 704282
rect 181794 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 182414 687454
rect 181794 687134 182414 687218
rect 181794 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 182414 687134
rect 181794 651454 182414 686898
rect 181794 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 182414 651454
rect 181794 651134 182414 651218
rect 181794 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 182414 651134
rect 181794 615454 182414 650898
rect 181794 615218 181826 615454
rect 182062 615218 182146 615454
rect 182382 615218 182414 615454
rect 181794 615134 182414 615218
rect 181794 614898 181826 615134
rect 182062 614898 182146 615134
rect 182382 614898 182414 615134
rect 181794 579454 182414 614898
rect 181794 579218 181826 579454
rect 182062 579218 182146 579454
rect 182382 579218 182414 579454
rect 181794 579134 182414 579218
rect 181794 578898 181826 579134
rect 182062 578898 182146 579134
rect 182382 578898 182414 579134
rect 181794 543454 182414 578898
rect 181794 543218 181826 543454
rect 182062 543218 182146 543454
rect 182382 543218 182414 543454
rect 181794 543134 182414 543218
rect 181794 542898 181826 543134
rect 182062 542898 182146 543134
rect 182382 542898 182414 543134
rect 181794 507454 182414 542898
rect 181794 507218 181826 507454
rect 182062 507218 182146 507454
rect 182382 507218 182414 507454
rect 181794 507134 182414 507218
rect 181794 506898 181826 507134
rect 182062 506898 182146 507134
rect 182382 506898 182414 507134
rect 181794 471454 182414 506898
rect 181794 471218 181826 471454
rect 182062 471218 182146 471454
rect 182382 471218 182414 471454
rect 181794 471134 182414 471218
rect 181794 470898 181826 471134
rect 182062 470898 182146 471134
rect 182382 470898 182414 471134
rect 181794 435454 182414 470898
rect 181794 435218 181826 435454
rect 182062 435218 182146 435454
rect 182382 435218 182414 435454
rect 181794 435134 182414 435218
rect 181794 434898 181826 435134
rect 182062 434898 182146 435134
rect 182382 434898 182414 435134
rect 181794 399454 182414 434898
rect 181794 399218 181826 399454
rect 182062 399218 182146 399454
rect 182382 399218 182414 399454
rect 181794 399134 182414 399218
rect 181794 398898 181826 399134
rect 182062 398898 182146 399134
rect 182382 398898 182414 399134
rect 181794 363454 182414 398898
rect 181794 363218 181826 363454
rect 182062 363218 182146 363454
rect 182382 363218 182414 363454
rect 181794 363134 182414 363218
rect 181794 362898 181826 363134
rect 182062 362898 182146 363134
rect 182382 362898 182414 363134
rect 181794 327454 182414 362898
rect 181794 327218 181826 327454
rect 182062 327218 182146 327454
rect 182382 327218 182414 327454
rect 181794 327134 182414 327218
rect 181794 326898 181826 327134
rect 182062 326898 182146 327134
rect 182382 326898 182414 327134
rect 181794 291454 182414 326898
rect 181794 291218 181826 291454
rect 182062 291218 182146 291454
rect 182382 291218 182414 291454
rect 181794 291134 182414 291218
rect 181794 290898 181826 291134
rect 182062 290898 182146 291134
rect 182382 290898 182414 291134
rect 181794 262000 182414 290898
rect 186294 705798 186914 711590
rect 186294 705562 186326 705798
rect 186562 705562 186646 705798
rect 186882 705562 186914 705798
rect 186294 705478 186914 705562
rect 186294 705242 186326 705478
rect 186562 705242 186646 705478
rect 186882 705242 186914 705478
rect 186294 691954 186914 705242
rect 186294 691718 186326 691954
rect 186562 691718 186646 691954
rect 186882 691718 186914 691954
rect 186294 691634 186914 691718
rect 186294 691398 186326 691634
rect 186562 691398 186646 691634
rect 186882 691398 186914 691634
rect 186294 655954 186914 691398
rect 186294 655718 186326 655954
rect 186562 655718 186646 655954
rect 186882 655718 186914 655954
rect 186294 655634 186914 655718
rect 186294 655398 186326 655634
rect 186562 655398 186646 655634
rect 186882 655398 186914 655634
rect 186294 619954 186914 655398
rect 186294 619718 186326 619954
rect 186562 619718 186646 619954
rect 186882 619718 186914 619954
rect 186294 619634 186914 619718
rect 186294 619398 186326 619634
rect 186562 619398 186646 619634
rect 186882 619398 186914 619634
rect 186294 583954 186914 619398
rect 186294 583718 186326 583954
rect 186562 583718 186646 583954
rect 186882 583718 186914 583954
rect 186294 583634 186914 583718
rect 186294 583398 186326 583634
rect 186562 583398 186646 583634
rect 186882 583398 186914 583634
rect 186294 547954 186914 583398
rect 186294 547718 186326 547954
rect 186562 547718 186646 547954
rect 186882 547718 186914 547954
rect 186294 547634 186914 547718
rect 186294 547398 186326 547634
rect 186562 547398 186646 547634
rect 186882 547398 186914 547634
rect 186294 511954 186914 547398
rect 186294 511718 186326 511954
rect 186562 511718 186646 511954
rect 186882 511718 186914 511954
rect 186294 511634 186914 511718
rect 186294 511398 186326 511634
rect 186562 511398 186646 511634
rect 186882 511398 186914 511634
rect 186294 475954 186914 511398
rect 186294 475718 186326 475954
rect 186562 475718 186646 475954
rect 186882 475718 186914 475954
rect 186294 475634 186914 475718
rect 186294 475398 186326 475634
rect 186562 475398 186646 475634
rect 186882 475398 186914 475634
rect 186294 439954 186914 475398
rect 186294 439718 186326 439954
rect 186562 439718 186646 439954
rect 186882 439718 186914 439954
rect 186294 439634 186914 439718
rect 186294 439398 186326 439634
rect 186562 439398 186646 439634
rect 186882 439398 186914 439634
rect 186294 403954 186914 439398
rect 186294 403718 186326 403954
rect 186562 403718 186646 403954
rect 186882 403718 186914 403954
rect 186294 403634 186914 403718
rect 186294 403398 186326 403634
rect 186562 403398 186646 403634
rect 186882 403398 186914 403634
rect 186294 367954 186914 403398
rect 186294 367718 186326 367954
rect 186562 367718 186646 367954
rect 186882 367718 186914 367954
rect 186294 367634 186914 367718
rect 186294 367398 186326 367634
rect 186562 367398 186646 367634
rect 186882 367398 186914 367634
rect 186294 331954 186914 367398
rect 186294 331718 186326 331954
rect 186562 331718 186646 331954
rect 186882 331718 186914 331954
rect 186294 331634 186914 331718
rect 186294 331398 186326 331634
rect 186562 331398 186646 331634
rect 186882 331398 186914 331634
rect 186294 295954 186914 331398
rect 186294 295718 186326 295954
rect 186562 295718 186646 295954
rect 186882 295718 186914 295954
rect 186294 295634 186914 295718
rect 186294 295398 186326 295634
rect 186562 295398 186646 295634
rect 186882 295398 186914 295634
rect 186294 262000 186914 295398
rect 190794 706758 191414 711590
rect 190794 706522 190826 706758
rect 191062 706522 191146 706758
rect 191382 706522 191414 706758
rect 190794 706438 191414 706522
rect 190794 706202 190826 706438
rect 191062 706202 191146 706438
rect 191382 706202 191414 706438
rect 190794 696454 191414 706202
rect 190794 696218 190826 696454
rect 191062 696218 191146 696454
rect 191382 696218 191414 696454
rect 190794 696134 191414 696218
rect 190794 695898 190826 696134
rect 191062 695898 191146 696134
rect 191382 695898 191414 696134
rect 190794 660454 191414 695898
rect 190794 660218 190826 660454
rect 191062 660218 191146 660454
rect 191382 660218 191414 660454
rect 190794 660134 191414 660218
rect 190794 659898 190826 660134
rect 191062 659898 191146 660134
rect 191382 659898 191414 660134
rect 190794 624454 191414 659898
rect 190794 624218 190826 624454
rect 191062 624218 191146 624454
rect 191382 624218 191414 624454
rect 190794 624134 191414 624218
rect 190794 623898 190826 624134
rect 191062 623898 191146 624134
rect 191382 623898 191414 624134
rect 190794 588454 191414 623898
rect 190794 588218 190826 588454
rect 191062 588218 191146 588454
rect 191382 588218 191414 588454
rect 190794 588134 191414 588218
rect 190794 587898 190826 588134
rect 191062 587898 191146 588134
rect 191382 587898 191414 588134
rect 190794 552454 191414 587898
rect 190794 552218 190826 552454
rect 191062 552218 191146 552454
rect 191382 552218 191414 552454
rect 190794 552134 191414 552218
rect 190794 551898 190826 552134
rect 191062 551898 191146 552134
rect 191382 551898 191414 552134
rect 190794 516454 191414 551898
rect 190794 516218 190826 516454
rect 191062 516218 191146 516454
rect 191382 516218 191414 516454
rect 190794 516134 191414 516218
rect 190794 515898 190826 516134
rect 191062 515898 191146 516134
rect 191382 515898 191414 516134
rect 190794 480454 191414 515898
rect 190794 480218 190826 480454
rect 191062 480218 191146 480454
rect 191382 480218 191414 480454
rect 190794 480134 191414 480218
rect 190794 479898 190826 480134
rect 191062 479898 191146 480134
rect 191382 479898 191414 480134
rect 190794 444454 191414 479898
rect 190794 444218 190826 444454
rect 191062 444218 191146 444454
rect 191382 444218 191414 444454
rect 190794 444134 191414 444218
rect 190794 443898 190826 444134
rect 191062 443898 191146 444134
rect 191382 443898 191414 444134
rect 190794 408454 191414 443898
rect 190794 408218 190826 408454
rect 191062 408218 191146 408454
rect 191382 408218 191414 408454
rect 190794 408134 191414 408218
rect 190794 407898 190826 408134
rect 191062 407898 191146 408134
rect 191382 407898 191414 408134
rect 190794 372454 191414 407898
rect 190794 372218 190826 372454
rect 191062 372218 191146 372454
rect 191382 372218 191414 372454
rect 190794 372134 191414 372218
rect 190794 371898 190826 372134
rect 191062 371898 191146 372134
rect 191382 371898 191414 372134
rect 190794 336454 191414 371898
rect 190794 336218 190826 336454
rect 191062 336218 191146 336454
rect 191382 336218 191414 336454
rect 190794 336134 191414 336218
rect 190794 335898 190826 336134
rect 191062 335898 191146 336134
rect 191382 335898 191414 336134
rect 190794 300454 191414 335898
rect 190794 300218 190826 300454
rect 191062 300218 191146 300454
rect 191382 300218 191414 300454
rect 190794 300134 191414 300218
rect 190794 299898 190826 300134
rect 191062 299898 191146 300134
rect 191382 299898 191414 300134
rect 187739 278084 187805 278085
rect 187739 278020 187740 278084
rect 187804 278020 187805 278084
rect 187739 278019 187805 278020
rect 187742 277541 187802 278019
rect 187739 277540 187805 277541
rect 187739 277476 187740 277540
rect 187804 277476 187805 277540
rect 187739 277475 187805 277476
rect 122787 260812 122853 260813
rect 122787 260810 122788 260812
rect 122606 260750 122788 260810
rect 121131 260268 121197 260269
rect 121131 260204 121132 260268
rect 121196 260204 121197 260268
rect 121131 260203 121197 260204
rect 118187 259860 118253 259861
rect 118187 259796 118188 259860
rect 118252 259796 118253 259860
rect 118187 259795 118253 259796
rect 117083 199476 117149 199477
rect 117083 199412 117084 199476
rect 117148 199412 117149 199476
rect 117083 199411 117149 199412
rect 116899 143852 116965 143853
rect 116899 143788 116900 143852
rect 116964 143788 116965 143852
rect 116899 143787 116965 143788
rect 116715 143444 116781 143445
rect 116715 143380 116716 143444
rect 116780 143380 116781 143444
rect 116715 143379 116781 143380
rect 116531 142356 116597 142357
rect 116531 142292 116532 142356
rect 116596 142292 116597 142356
rect 116531 142291 116597 142292
rect 115795 66196 115861 66197
rect 115795 66132 115796 66196
rect 115860 66132 115861 66196
rect 115795 66131 115861 66132
rect 115059 63340 115125 63341
rect 115059 63276 115060 63340
rect 115124 63276 115125 63340
rect 115059 63275 115125 63276
rect 116534 44301 116594 142291
rect 116715 141540 116781 141541
rect 116715 141476 116716 141540
rect 116780 141476 116781 141540
rect 116715 141475 116781 141476
rect 116718 68781 116778 141475
rect 116899 138004 116965 138005
rect 116899 137940 116900 138004
rect 116964 137940 116965 138004
rect 116899 137939 116965 137940
rect 116715 68780 116781 68781
rect 116715 68716 116716 68780
rect 116780 68716 116781 68780
rect 116715 68715 116781 68716
rect 116902 50829 116962 137939
rect 117086 73133 117146 199411
rect 118190 143989 118250 259795
rect 118371 195532 118437 195533
rect 118371 195468 118372 195532
rect 118436 195468 118437 195532
rect 118371 195467 118437 195468
rect 118187 143988 118253 143989
rect 118187 143924 118188 143988
rect 118252 143924 118253 143988
rect 118187 143923 118253 143924
rect 117819 141404 117885 141405
rect 117819 141340 117820 141404
rect 117884 141340 117885 141404
rect 117819 141339 117885 141340
rect 117822 84285 117882 141339
rect 118187 137460 118253 137461
rect 118187 137396 118188 137460
rect 118252 137396 118253 137460
rect 118187 137395 118253 137396
rect 117819 84284 117885 84285
rect 117819 84220 117820 84284
rect 117884 84220 117885 84284
rect 117819 84219 117885 84220
rect 118190 80205 118250 137395
rect 118187 80204 118253 80205
rect 118187 80140 118188 80204
rect 118252 80140 118253 80204
rect 118187 80139 118253 80140
rect 118374 74493 118434 195467
rect 118794 192454 119414 198000
rect 119843 195260 119909 195261
rect 119843 195196 119844 195260
rect 119908 195196 119909 195260
rect 119843 195195 119909 195196
rect 118794 192218 118826 192454
rect 119062 192218 119146 192454
rect 119382 192218 119414 192454
rect 118794 192134 119414 192218
rect 118794 191898 118826 192134
rect 119062 191898 119146 192134
rect 119382 191898 119414 192134
rect 118555 191452 118621 191453
rect 118555 191388 118556 191452
rect 118620 191388 118621 191452
rect 118555 191387 118621 191388
rect 118371 74492 118437 74493
rect 118371 74428 118372 74492
rect 118436 74428 118437 74492
rect 118371 74427 118437 74428
rect 117083 73132 117149 73133
rect 117083 73068 117084 73132
rect 117148 73068 117149 73132
rect 117083 73067 117149 73068
rect 118558 66061 118618 191387
rect 118794 156454 119414 191898
rect 118794 156218 118826 156454
rect 119062 156218 119146 156454
rect 119382 156218 119414 156454
rect 118794 156134 119414 156218
rect 118794 155898 118826 156134
rect 119062 155898 119146 156134
rect 119382 155898 119414 156134
rect 118794 142000 119414 155898
rect 119659 148340 119725 148341
rect 119659 148276 119660 148340
rect 119724 148276 119725 148340
rect 119659 148275 119725 148276
rect 119475 140588 119541 140589
rect 119475 140524 119476 140588
rect 119540 140524 119541 140588
rect 119475 140523 119541 140524
rect 118739 139500 118805 139501
rect 118739 139436 118740 139500
rect 118804 139436 118805 139500
rect 118739 139435 118805 139436
rect 118742 96661 118802 139435
rect 118739 96660 118805 96661
rect 118739 96596 118740 96660
rect 118804 96596 118805 96660
rect 118739 96595 118805 96596
rect 119478 78709 119538 140523
rect 119475 78708 119541 78709
rect 119475 78644 119476 78708
rect 119540 78644 119541 78708
rect 119475 78643 119541 78644
rect 118555 66060 118621 66061
rect 118555 65996 118556 66060
rect 118620 65996 118621 66060
rect 118555 65995 118621 65996
rect 116899 50828 116965 50829
rect 116899 50764 116900 50828
rect 116964 50764 116965 50828
rect 116899 50763 116965 50764
rect 118794 48454 119414 78000
rect 119662 70410 119722 148275
rect 119846 78573 119906 195195
rect 120763 146028 120829 146029
rect 120763 145964 120764 146028
rect 120828 145964 120829 146028
rect 120763 145963 120829 145964
rect 120579 139908 120645 139909
rect 120579 139844 120580 139908
rect 120644 139844 120645 139908
rect 120579 139843 120645 139844
rect 119843 78572 119909 78573
rect 119843 78508 119844 78572
rect 119908 78508 119909 78572
rect 119843 78507 119909 78508
rect 119846 75173 119906 78507
rect 119843 75172 119909 75173
rect 119843 75108 119844 75172
rect 119908 75108 119909 75172
rect 119843 75107 119909 75108
rect 119662 70350 120090 70410
rect 120030 70141 120090 70350
rect 120027 70140 120093 70141
rect 120027 70076 120028 70140
rect 120092 70076 120093 70140
rect 120027 70075 120093 70076
rect 118794 48218 118826 48454
rect 119062 48218 119146 48454
rect 119382 48218 119414 48454
rect 118794 48134 119414 48218
rect 118794 47898 118826 48134
rect 119062 47898 119146 48134
rect 119382 47898 119414 48134
rect 116531 44300 116597 44301
rect 116531 44236 116532 44300
rect 116596 44236 116597 44300
rect 116531 44235 116597 44236
rect 114294 43718 114326 43954
rect 114562 43718 114646 43954
rect 114882 43718 114914 43954
rect 114294 43634 114914 43718
rect 114294 43398 114326 43634
rect 114562 43398 114646 43634
rect 114882 43398 114914 43634
rect 114294 7954 114914 43398
rect 114294 7718 114326 7954
rect 114562 7718 114646 7954
rect 114882 7718 114914 7954
rect 114294 7634 114914 7718
rect 114294 7398 114326 7634
rect 114562 7398 114646 7634
rect 114882 7398 114914 7634
rect 114294 -1306 114914 7398
rect 114294 -1542 114326 -1306
rect 114562 -1542 114646 -1306
rect 114882 -1542 114914 -1306
rect 114294 -1626 114914 -1542
rect 114294 -1862 114326 -1626
rect 114562 -1862 114646 -1626
rect 114882 -1862 114914 -1626
rect 114294 -7654 114914 -1862
rect 118794 12454 119414 47898
rect 120582 31789 120642 139843
rect 120766 70005 120826 145963
rect 121134 143037 121194 260203
rect 121315 259996 121381 259997
rect 121315 259932 121316 259996
rect 121380 259932 121381 259996
rect 121315 259931 121381 259932
rect 121131 143036 121197 143037
rect 121131 142972 121132 143036
rect 121196 142972 121197 143036
rect 121131 142971 121197 142972
rect 121318 142901 121378 259931
rect 122606 200130 122666 260750
rect 122787 260748 122788 260750
rect 122852 260748 122853 260812
rect 122787 260747 122853 260748
rect 124075 259588 124141 259589
rect 124075 259524 124076 259588
rect 124140 259524 124141 259588
rect 124075 259523 124141 259524
rect 122971 259452 123037 259453
rect 122971 259388 122972 259452
rect 123036 259388 123037 259452
rect 122971 259387 123037 259388
rect 122787 200156 122853 200157
rect 122787 200130 122788 200156
rect 122606 200092 122788 200130
rect 122852 200092 122853 200156
rect 122606 200091 122853 200092
rect 122606 200070 122850 200091
rect 122974 198797 123034 259387
rect 122971 198796 123037 198797
rect 122971 198732 122972 198796
rect 123036 198732 123037 198796
rect 122971 198731 123037 198732
rect 123294 196954 123914 198000
rect 123294 196718 123326 196954
rect 123562 196718 123646 196954
rect 123882 196718 123914 196954
rect 123294 196634 123914 196718
rect 123294 196398 123326 196634
rect 123562 196398 123646 196634
rect 123882 196398 123914 196634
rect 123294 160954 123914 196398
rect 123294 160718 123326 160954
rect 123562 160718 123646 160954
rect 123882 160718 123914 160954
rect 123294 160634 123914 160718
rect 123294 160398 123326 160634
rect 123562 160398 123646 160634
rect 123882 160398 123914 160634
rect 122419 151196 122485 151197
rect 122419 151132 122420 151196
rect 122484 151132 122485 151196
rect 122419 151131 122485 151132
rect 122051 147116 122117 147117
rect 122051 147052 122052 147116
rect 122116 147052 122117 147116
rect 122051 147051 122117 147052
rect 121315 142900 121381 142901
rect 121315 142836 121316 142900
rect 121380 142836 121381 142900
rect 121315 142835 121381 142836
rect 121131 141676 121197 141677
rect 121131 141612 121132 141676
rect 121196 141612 121197 141676
rect 121131 141611 121197 141612
rect 120947 140452 121013 140453
rect 120947 140388 120948 140452
rect 121012 140388 121013 140452
rect 120947 140387 121013 140388
rect 120950 78981 121010 140387
rect 120947 78980 121013 78981
rect 120947 78916 120948 78980
rect 121012 78916 121013 78980
rect 120947 78915 121013 78916
rect 120763 70004 120829 70005
rect 120763 69940 120764 70004
rect 120828 69940 120829 70004
rect 120763 69939 120829 69940
rect 121134 69869 121194 141611
rect 122054 137461 122114 147051
rect 122235 138548 122301 138549
rect 122235 138484 122236 138548
rect 122300 138484 122301 138548
rect 122235 138483 122301 138484
rect 122051 137460 122117 137461
rect 122051 137396 122052 137460
rect 122116 137396 122117 137460
rect 122051 137395 122117 137396
rect 122238 74357 122298 138483
rect 122422 138141 122482 151131
rect 122971 151060 123037 151061
rect 122971 150996 122972 151060
rect 123036 150996 123037 151060
rect 122971 150995 123037 150996
rect 122603 140044 122669 140045
rect 122603 139980 122604 140044
rect 122668 139980 122669 140044
rect 122603 139979 122669 139980
rect 122419 138140 122485 138141
rect 122419 138076 122420 138140
rect 122484 138076 122485 138140
rect 122419 138075 122485 138076
rect 122419 138004 122485 138005
rect 122419 137940 122420 138004
rect 122484 137940 122485 138004
rect 122419 137939 122485 137940
rect 122235 74356 122301 74357
rect 122235 74292 122236 74356
rect 122300 74292 122301 74356
rect 122235 74291 122301 74292
rect 121131 69868 121197 69869
rect 121131 69804 121132 69868
rect 121196 69804 121197 69868
rect 121131 69803 121197 69804
rect 122422 68645 122482 137939
rect 122606 69733 122666 139979
rect 122974 137325 123034 150995
rect 123294 142000 123914 160398
rect 124078 150517 124138 259523
rect 186083 259452 186149 259453
rect 186083 259388 186084 259452
rect 186148 259388 186149 259452
rect 186083 259387 186149 259388
rect 124208 255454 124528 255486
rect 124208 255218 124250 255454
rect 124486 255218 124528 255454
rect 124208 255134 124528 255218
rect 124208 254898 124250 255134
rect 124486 254898 124528 255134
rect 124208 254866 124528 254898
rect 154928 255454 155248 255486
rect 154928 255218 154970 255454
rect 155206 255218 155248 255454
rect 154928 255134 155248 255218
rect 154928 254898 154970 255134
rect 155206 254898 155248 255134
rect 154928 254866 155248 254898
rect 185648 255454 185968 255486
rect 185648 255218 185690 255454
rect 185926 255218 185968 255454
rect 185648 255134 185968 255218
rect 185648 254898 185690 255134
rect 185926 254898 185968 255134
rect 185648 254866 185968 254898
rect 139568 223954 139888 223986
rect 139568 223718 139610 223954
rect 139846 223718 139888 223954
rect 139568 223634 139888 223718
rect 139568 223398 139610 223634
rect 139846 223398 139888 223634
rect 139568 223366 139888 223398
rect 170288 223954 170608 223986
rect 170288 223718 170330 223954
rect 170566 223718 170608 223954
rect 170288 223634 170608 223718
rect 170288 223398 170330 223634
rect 170566 223398 170608 223634
rect 170288 223366 170608 223398
rect 124208 219454 124528 219486
rect 124208 219218 124250 219454
rect 124486 219218 124528 219454
rect 124208 219134 124528 219218
rect 124208 218898 124250 219134
rect 124486 218898 124528 219134
rect 124208 218866 124528 218898
rect 154928 219454 155248 219486
rect 154928 219218 154970 219454
rect 155206 219218 155248 219454
rect 154928 219134 155248 219218
rect 154928 218898 154970 219134
rect 155206 218898 155248 219134
rect 154928 218866 155248 218898
rect 185648 219454 185968 219486
rect 185648 219218 185690 219454
rect 185926 219218 185968 219454
rect 185648 219134 185968 219218
rect 185648 218898 185690 219134
rect 185926 218898 185968 219134
rect 185648 218866 185968 218898
rect 186086 213893 186146 259387
rect 186083 213892 186149 213893
rect 186083 213828 186084 213892
rect 186148 213828 186149 213892
rect 186083 213827 186149 213828
rect 131619 201516 131685 201517
rect 131619 201452 131620 201516
rect 131684 201452 131685 201516
rect 131619 201451 131685 201452
rect 139531 201516 139597 201517
rect 139531 201452 139532 201516
rect 139596 201452 139597 201516
rect 139531 201451 139597 201452
rect 124811 192540 124877 192541
rect 124811 192476 124812 192540
rect 124876 192476 124877 192540
rect 124811 192475 124877 192476
rect 124075 150516 124141 150517
rect 124075 150452 124076 150516
rect 124140 150452 124141 150516
rect 124075 150451 124141 150452
rect 123155 139364 123221 139365
rect 123155 139300 123156 139364
rect 123220 139300 123221 139364
rect 123155 139299 123221 139300
rect 122971 137324 123037 137325
rect 122971 137260 122972 137324
rect 123036 137260 123037 137324
rect 122971 137259 123037 137260
rect 122971 133924 123037 133925
rect 122971 133860 122972 133924
rect 123036 133860 123037 133924
rect 122971 133859 123037 133860
rect 122974 86189 123034 133859
rect 122971 86188 123037 86189
rect 122971 86124 122972 86188
rect 123036 86124 123037 86188
rect 122971 86123 123037 86124
rect 122971 86052 123037 86053
rect 122971 85988 122972 86052
rect 123036 86050 123037 86052
rect 123158 86050 123218 139299
rect 124814 138005 124874 192475
rect 131622 147525 131682 201451
rect 132723 199884 132789 199885
rect 132723 199820 132724 199884
rect 132788 199820 132789 199884
rect 132723 199819 132789 199820
rect 133827 199884 133893 199885
rect 133827 199820 133828 199884
rect 133892 199820 133893 199884
rect 133827 199819 133893 199820
rect 134747 199884 134813 199885
rect 134747 199820 134748 199884
rect 134812 199820 134813 199884
rect 134747 199819 134813 199820
rect 135483 199884 135549 199885
rect 135483 199820 135484 199884
rect 135548 199820 135549 199884
rect 135483 199819 135549 199820
rect 135851 199884 135917 199885
rect 135851 199820 135852 199884
rect 135916 199820 135917 199884
rect 135851 199819 135917 199820
rect 138243 199884 138309 199885
rect 138243 199820 138244 199884
rect 138308 199820 138309 199884
rect 138243 199819 138309 199820
rect 132726 197370 132786 199819
rect 133643 199748 133709 199749
rect 133643 199684 133644 199748
rect 133708 199684 133709 199748
rect 133643 199683 133709 199684
rect 133646 197981 133706 199683
rect 133643 197980 133709 197981
rect 133643 197916 133644 197980
rect 133708 197916 133709 197980
rect 133643 197915 133709 197916
rect 132542 197310 132786 197370
rect 132542 186965 132602 197310
rect 133830 195261 133890 199819
rect 134011 197436 134077 197437
rect 134011 197372 134012 197436
rect 134076 197372 134077 197436
rect 134011 197371 134077 197372
rect 133827 195260 133893 195261
rect 133827 195196 133828 195260
rect 133892 195196 133893 195260
rect 133827 195195 133893 195196
rect 133827 192948 133893 192949
rect 133827 192884 133828 192948
rect 133892 192884 133893 192948
rect 133827 192883 133893 192884
rect 133830 191589 133890 192883
rect 133827 191588 133893 191589
rect 133827 191524 133828 191588
rect 133892 191524 133893 191588
rect 133827 191523 133893 191524
rect 134014 191181 134074 197371
rect 134750 195941 134810 199819
rect 135161 199068 135227 199069
rect 135161 199066 135162 199068
rect 135118 199004 135162 199066
rect 135226 199004 135227 199068
rect 135118 199003 135227 199004
rect 135118 198525 135178 199003
rect 135115 198524 135181 198525
rect 135115 198460 135116 198524
rect 135180 198460 135181 198524
rect 135115 198459 135181 198460
rect 135299 197708 135365 197709
rect 135299 197644 135300 197708
rect 135364 197644 135365 197708
rect 135299 197643 135365 197644
rect 134747 195940 134813 195941
rect 134747 195876 134748 195940
rect 134812 195876 134813 195940
rect 134747 195875 134813 195876
rect 134011 191180 134077 191181
rect 134011 191116 134012 191180
rect 134076 191116 134077 191180
rect 134011 191115 134077 191116
rect 135302 191045 135362 197643
rect 135486 197573 135546 199819
rect 135483 197572 135549 197573
rect 135483 197508 135484 197572
rect 135548 197508 135549 197572
rect 135483 197507 135549 197508
rect 135854 193230 135914 199819
rect 137139 199748 137205 199749
rect 137139 199684 137140 199748
rect 137204 199684 137205 199748
rect 137139 199683 137205 199684
rect 137875 199748 137941 199749
rect 137875 199684 137876 199748
rect 137940 199684 137941 199748
rect 137875 199683 137941 199684
rect 137142 199069 137202 199683
rect 137139 199068 137205 199069
rect 137139 199004 137140 199068
rect 137204 199004 137205 199068
rect 137139 199003 137205 199004
rect 136771 198116 136837 198117
rect 136771 198052 136772 198116
rect 136836 198052 136837 198116
rect 136771 198051 136837 198052
rect 136587 196756 136653 196757
rect 136587 196692 136588 196756
rect 136652 196692 136653 196756
rect 136587 196691 136653 196692
rect 135486 193170 135914 193230
rect 135486 191317 135546 193170
rect 135483 191316 135549 191317
rect 135483 191252 135484 191316
rect 135548 191252 135549 191316
rect 135483 191251 135549 191252
rect 135299 191044 135365 191045
rect 135299 190980 135300 191044
rect 135364 190980 135365 191044
rect 135299 190979 135365 190980
rect 132539 186964 132605 186965
rect 132539 186900 132540 186964
rect 132604 186900 132605 186964
rect 132539 186899 132605 186900
rect 131619 147524 131685 147525
rect 131619 147460 131620 147524
rect 131684 147460 131685 147524
rect 131619 147459 131685 147460
rect 136590 146981 136650 196691
rect 136774 148477 136834 198051
rect 137878 196621 137938 199683
rect 137875 196620 137941 196621
rect 137875 196556 137876 196620
rect 137940 196556 137941 196620
rect 137875 196555 137941 196556
rect 138059 195124 138125 195125
rect 138059 195060 138060 195124
rect 138124 195060 138125 195124
rect 138059 195059 138125 195060
rect 138062 187101 138122 195059
rect 138246 187373 138306 199819
rect 139534 199749 139594 201451
rect 154619 200700 154685 200701
rect 154619 200636 154620 200700
rect 154684 200636 154685 200700
rect 154619 200635 154685 200636
rect 173571 200700 173637 200701
rect 173571 200636 173572 200700
rect 173636 200636 173637 200700
rect 173571 200635 173637 200636
rect 150939 200564 151005 200565
rect 150939 200500 150940 200564
rect 151004 200500 151005 200564
rect 150939 200499 151005 200500
rect 142291 200156 142357 200157
rect 142291 200092 142292 200156
rect 142356 200092 142357 200156
rect 142291 200091 142357 200092
rect 150019 200156 150085 200157
rect 150019 200092 150020 200156
rect 150084 200092 150085 200156
rect 150019 200091 150085 200092
rect 141555 199884 141621 199885
rect 141555 199820 141556 199884
rect 141620 199820 141621 199884
rect 141555 199819 141621 199820
rect 142107 199884 142173 199885
rect 142107 199820 142108 199884
rect 142172 199820 142173 199884
rect 142107 199819 142173 199820
rect 139531 199748 139597 199749
rect 139531 199684 139532 199748
rect 139596 199684 139597 199748
rect 139531 199683 139597 199684
rect 139531 199612 139597 199613
rect 139531 199548 139532 199612
rect 139596 199548 139597 199612
rect 139531 199547 139597 199548
rect 138795 198116 138861 198117
rect 138795 198052 138796 198116
rect 138860 198052 138861 198116
rect 138795 198051 138861 198052
rect 138427 195260 138493 195261
rect 138427 195196 138428 195260
rect 138492 195196 138493 195260
rect 138427 195195 138493 195196
rect 138430 190229 138490 195195
rect 138798 191725 138858 198051
rect 139347 196756 139413 196757
rect 139347 196692 139348 196756
rect 139412 196692 139413 196756
rect 139347 196691 139413 196692
rect 138795 191724 138861 191725
rect 138795 191660 138796 191724
rect 138860 191660 138861 191724
rect 138795 191659 138861 191660
rect 138427 190228 138493 190229
rect 138427 190164 138428 190228
rect 138492 190164 138493 190228
rect 138427 190163 138493 190164
rect 138243 187372 138309 187373
rect 138243 187308 138244 187372
rect 138308 187308 138309 187372
rect 138243 187307 138309 187308
rect 138059 187100 138125 187101
rect 138059 187036 138060 187100
rect 138124 187036 138125 187100
rect 138059 187035 138125 187036
rect 139350 151197 139410 196691
rect 139534 187237 139594 199547
rect 141558 199205 141618 199819
rect 141739 199748 141805 199749
rect 141739 199684 141740 199748
rect 141804 199684 141805 199748
rect 141739 199683 141805 199684
rect 141742 199205 141802 199683
rect 142110 199205 142170 199819
rect 141555 199204 141621 199205
rect 141555 199140 141556 199204
rect 141620 199140 141621 199204
rect 141555 199139 141621 199140
rect 141739 199204 141805 199205
rect 141739 199140 141740 199204
rect 141804 199140 141805 199204
rect 141739 199139 141805 199140
rect 142107 199204 142173 199205
rect 142107 199140 142108 199204
rect 142172 199140 142173 199204
rect 142107 199139 142173 199140
rect 139531 187236 139597 187237
rect 139531 187172 139532 187236
rect 139596 187172 139597 187236
rect 139531 187171 139597 187172
rect 141294 178954 141914 198000
rect 142107 197572 142173 197573
rect 142107 197508 142108 197572
rect 142172 197508 142173 197572
rect 142107 197507 142173 197508
rect 142110 187645 142170 197507
rect 142294 190093 142354 200091
rect 142659 199884 142725 199885
rect 142659 199820 142660 199884
rect 142724 199820 142725 199884
rect 142659 199819 142725 199820
rect 143211 199884 143277 199885
rect 143211 199820 143212 199884
rect 143276 199820 143277 199884
rect 143211 199819 143277 199820
rect 143395 199884 143461 199885
rect 143395 199820 143396 199884
rect 143460 199820 143461 199884
rect 143395 199819 143461 199820
rect 146155 199884 146221 199885
rect 146155 199820 146156 199884
rect 146220 199820 146221 199884
rect 146155 199819 146221 199820
rect 142475 199612 142541 199613
rect 142475 199548 142476 199612
rect 142540 199548 142541 199612
rect 142475 199547 142541 199548
rect 142291 190092 142357 190093
rect 142291 190028 142292 190092
rect 142356 190028 142357 190092
rect 142291 190027 142357 190028
rect 142478 189821 142538 199547
rect 142662 198525 142722 199819
rect 143027 199748 143093 199749
rect 143027 199684 143028 199748
rect 143092 199684 143093 199748
rect 143027 199683 143093 199684
rect 143030 198525 143090 199683
rect 143214 199205 143274 199819
rect 143211 199204 143277 199205
rect 143211 199140 143212 199204
rect 143276 199140 143277 199204
rect 143211 199139 143277 199140
rect 143398 198525 143458 199819
rect 143579 198660 143645 198661
rect 143579 198596 143580 198660
rect 143644 198596 143645 198660
rect 143579 198595 143645 198596
rect 144315 198660 144381 198661
rect 144315 198596 144316 198660
rect 144380 198596 144381 198660
rect 144315 198595 144381 198596
rect 142659 198524 142725 198525
rect 142659 198460 142660 198524
rect 142724 198460 142725 198524
rect 142659 198459 142725 198460
rect 143027 198524 143093 198525
rect 143027 198460 143028 198524
rect 143092 198460 143093 198524
rect 143027 198459 143093 198460
rect 143395 198524 143461 198525
rect 143395 198460 143396 198524
rect 143460 198460 143461 198524
rect 143395 198459 143461 198460
rect 142475 189820 142541 189821
rect 142475 189756 142476 189820
rect 142540 189756 142541 189820
rect 142475 189755 142541 189756
rect 142107 187644 142173 187645
rect 142107 187580 142108 187644
rect 142172 187580 142173 187644
rect 142107 187579 142173 187580
rect 141294 178718 141326 178954
rect 141562 178718 141646 178954
rect 141882 178718 141914 178954
rect 141294 178634 141914 178718
rect 141294 178398 141326 178634
rect 141562 178398 141646 178634
rect 141882 178398 141914 178634
rect 139347 151196 139413 151197
rect 139347 151132 139348 151196
rect 139412 151132 139413 151196
rect 139347 151131 139413 151132
rect 136771 148476 136837 148477
rect 136771 148412 136772 148476
rect 136836 148412 136837 148476
rect 136771 148411 136837 148412
rect 136587 146980 136653 146981
rect 136587 146916 136588 146980
rect 136652 146916 136653 146980
rect 136587 146915 136653 146916
rect 141294 142954 141914 178398
rect 143582 144125 143642 198595
rect 143947 197436 144013 197437
rect 143947 197372 143948 197436
rect 144012 197372 144013 197436
rect 143947 197371 144013 197372
rect 143763 196756 143829 196757
rect 143763 196692 143764 196756
rect 143828 196692 143829 196756
rect 143763 196691 143829 196692
rect 143766 189685 143826 196691
rect 143950 189957 144010 197371
rect 144318 192677 144378 198595
rect 146158 198525 146218 199819
rect 147443 199612 147509 199613
rect 147443 199548 147444 199612
rect 147508 199548 147509 199612
rect 147443 199547 147509 199548
rect 146155 198524 146221 198525
rect 146155 198460 146156 198524
rect 146220 198460 146221 198524
rect 146155 198459 146221 198460
rect 146891 198252 146957 198253
rect 146891 198188 146892 198252
rect 146956 198188 146957 198252
rect 146891 198187 146957 198188
rect 144315 192676 144381 192677
rect 144315 192612 144316 192676
rect 144380 192612 144381 192676
rect 144315 192611 144381 192612
rect 143947 189956 144013 189957
rect 143947 189892 143948 189956
rect 144012 189892 144013 189956
rect 143947 189891 144013 189892
rect 143763 189684 143829 189685
rect 143763 189620 143764 189684
rect 143828 189620 143829 189684
rect 143763 189619 143829 189620
rect 145794 183454 146414 198000
rect 145794 183218 145826 183454
rect 146062 183218 146146 183454
rect 146382 183218 146414 183454
rect 145794 183134 146414 183218
rect 145794 182898 145826 183134
rect 146062 182898 146146 183134
rect 146382 182898 146414 183134
rect 145794 147454 146414 182898
rect 145794 147218 145826 147454
rect 146062 147218 146146 147454
rect 146382 147218 146414 147454
rect 145794 147134 146414 147218
rect 145794 146898 145826 147134
rect 146062 146898 146146 147134
rect 146382 146898 146414 147134
rect 143579 144124 143645 144125
rect 143579 144060 143580 144124
rect 143644 144060 143645 144124
rect 143579 144059 143645 144060
rect 141294 142718 141326 142954
rect 141562 142718 141646 142954
rect 141882 142718 141914 142954
rect 141294 142634 141914 142718
rect 141294 142398 141326 142634
rect 141562 142398 141646 142634
rect 141882 142398 141914 142634
rect 141294 142000 141914 142398
rect 145794 142000 146414 146898
rect 128859 140044 128925 140045
rect 128859 139980 128860 140044
rect 128924 139980 128925 140044
rect 128859 139979 128925 139980
rect 130331 140044 130397 140045
rect 130331 139980 130332 140044
rect 130396 139980 130397 140044
rect 130331 139979 130397 139980
rect 128862 138549 128922 139979
rect 130334 138821 130394 139979
rect 130331 138820 130397 138821
rect 130331 138756 130332 138820
rect 130396 138756 130397 138820
rect 130331 138755 130397 138756
rect 146894 138685 146954 198187
rect 147259 197708 147325 197709
rect 147259 197644 147260 197708
rect 147324 197644 147325 197708
rect 147259 197643 147325 197644
rect 147075 197572 147141 197573
rect 147075 197508 147076 197572
rect 147140 197508 147141 197572
rect 147075 197507 147141 197508
rect 147078 144261 147138 197507
rect 147262 147117 147322 197643
rect 147446 197165 147506 199547
rect 148731 198660 148797 198661
rect 148731 198596 148732 198660
rect 148796 198596 148797 198660
rect 148731 198595 148797 198596
rect 147443 197164 147509 197165
rect 147443 197100 147444 197164
rect 147508 197100 147509 197164
rect 147443 197099 147509 197100
rect 147443 197028 147509 197029
rect 147443 196964 147444 197028
rect 147508 196964 147509 197028
rect 147443 196963 147509 196964
rect 147446 193085 147506 196963
rect 147443 193084 147509 193085
rect 147443 193020 147444 193084
rect 147508 193020 147509 193084
rect 147443 193019 147509 193020
rect 148734 159357 148794 198595
rect 148915 198388 148981 198389
rect 148915 198324 148916 198388
rect 148980 198324 148981 198388
rect 148915 198323 148981 198324
rect 148731 159356 148797 159357
rect 148731 159292 148732 159356
rect 148796 159292 148797 159356
rect 148731 159291 148797 159292
rect 148918 151061 148978 198323
rect 149651 198116 149717 198117
rect 149651 198052 149652 198116
rect 149716 198052 149717 198116
rect 149651 198051 149717 198052
rect 149835 198116 149901 198117
rect 149835 198052 149836 198116
rect 149900 198052 149901 198116
rect 149835 198051 149901 198052
rect 149654 186965 149714 198051
rect 149838 187101 149898 198051
rect 149835 187100 149901 187101
rect 149835 187036 149836 187100
rect 149900 187036 149901 187100
rect 149835 187035 149901 187036
rect 149651 186964 149717 186965
rect 149651 186900 149652 186964
rect 149716 186900 149717 186964
rect 149651 186899 149717 186900
rect 148915 151060 148981 151061
rect 148915 150996 148916 151060
rect 148980 150996 148981 151060
rect 148915 150995 148981 150996
rect 150022 147253 150082 200091
rect 150942 199613 151002 200499
rect 154622 199885 154682 200635
rect 163083 200564 163149 200565
rect 163083 200500 163084 200564
rect 163148 200500 163149 200564
rect 163083 200499 163149 200500
rect 151859 199884 151925 199885
rect 151859 199820 151860 199884
rect 151924 199820 151925 199884
rect 151859 199819 151925 199820
rect 154619 199884 154685 199885
rect 154619 199820 154620 199884
rect 154684 199820 154685 199884
rect 154619 199819 154685 199820
rect 157379 199884 157445 199885
rect 157379 199820 157380 199884
rect 157444 199820 157445 199884
rect 157379 199819 157445 199820
rect 159035 199884 159101 199885
rect 159035 199820 159036 199884
rect 159100 199820 159101 199884
rect 159035 199819 159101 199820
rect 161059 199884 161125 199885
rect 161059 199820 161060 199884
rect 161124 199820 161125 199884
rect 161059 199819 161125 199820
rect 162163 199884 162229 199885
rect 162163 199820 162164 199884
rect 162228 199820 162229 199884
rect 162163 199819 162229 199820
rect 162531 199884 162597 199885
rect 162531 199820 162532 199884
rect 162596 199820 162597 199884
rect 162531 199819 162597 199820
rect 150939 199612 151005 199613
rect 150939 199548 150940 199612
rect 151004 199548 151005 199612
rect 150939 199547 151005 199548
rect 151862 199069 151922 199819
rect 156827 199476 156893 199477
rect 156827 199412 156828 199476
rect 156892 199412 156893 199476
rect 156827 199411 156893 199412
rect 151859 199068 151925 199069
rect 151859 199004 151860 199068
rect 151924 199004 151925 199068
rect 151859 199003 151925 199004
rect 152963 198116 153029 198117
rect 152963 198052 152964 198116
rect 153028 198052 153029 198116
rect 152963 198051 153029 198052
rect 154435 198116 154501 198117
rect 154435 198052 154436 198116
rect 154500 198052 154501 198116
rect 154435 198051 154501 198052
rect 156643 198116 156709 198117
rect 156643 198052 156644 198116
rect 156708 198052 156709 198116
rect 156643 198051 156709 198052
rect 150294 187954 150914 198000
rect 150294 187718 150326 187954
rect 150562 187718 150646 187954
rect 150882 187718 150914 187954
rect 150294 187634 150914 187718
rect 150294 187398 150326 187634
rect 150562 187398 150646 187634
rect 150882 187398 150914 187634
rect 150294 151954 150914 187398
rect 152966 187237 153026 198051
rect 154438 189685 154498 198051
rect 154794 192454 155414 198000
rect 156646 195533 156706 198051
rect 156643 195532 156709 195533
rect 156643 195468 156644 195532
rect 156708 195468 156709 195532
rect 156643 195467 156709 195468
rect 154794 192218 154826 192454
rect 155062 192218 155146 192454
rect 155382 192218 155414 192454
rect 154794 192134 155414 192218
rect 154794 191898 154826 192134
rect 155062 191898 155146 192134
rect 155382 191898 155414 192134
rect 154435 189684 154501 189685
rect 154435 189620 154436 189684
rect 154500 189620 154501 189684
rect 154435 189619 154501 189620
rect 152963 187236 153029 187237
rect 152963 187172 152964 187236
rect 153028 187172 153029 187236
rect 152963 187171 153029 187172
rect 150294 151718 150326 151954
rect 150562 151718 150646 151954
rect 150882 151718 150914 151954
rect 150294 151634 150914 151718
rect 150294 151398 150326 151634
rect 150562 151398 150646 151634
rect 150882 151398 150914 151634
rect 150019 147252 150085 147253
rect 150019 147188 150020 147252
rect 150084 147188 150085 147252
rect 150019 147187 150085 147188
rect 147259 147116 147325 147117
rect 147259 147052 147260 147116
rect 147324 147052 147325 147116
rect 147259 147051 147325 147052
rect 147075 144260 147141 144261
rect 147075 144196 147076 144260
rect 147140 144196 147141 144260
rect 147075 144195 147141 144196
rect 150294 142000 150914 151398
rect 154794 156454 155414 191898
rect 154794 156218 154826 156454
rect 155062 156218 155146 156454
rect 155382 156218 155414 156454
rect 154794 156134 155414 156218
rect 154794 155898 154826 156134
rect 155062 155898 155146 156134
rect 155382 155898 155414 156134
rect 154794 142000 155414 155898
rect 156830 149701 156890 199411
rect 157382 198253 157442 199819
rect 158483 198388 158549 198389
rect 158483 198324 158484 198388
rect 158548 198324 158549 198388
rect 158483 198323 158549 198324
rect 157379 198252 157445 198253
rect 157379 198188 157380 198252
rect 157444 198188 157445 198252
rect 157379 198187 157445 198188
rect 157195 198116 157261 198117
rect 157195 198052 157196 198116
rect 157260 198052 157261 198116
rect 157195 198051 157261 198052
rect 157198 195805 157258 198051
rect 157195 195804 157261 195805
rect 157195 195740 157196 195804
rect 157260 195740 157261 195804
rect 157195 195739 157261 195740
rect 156827 149700 156893 149701
rect 156827 149636 156828 149700
rect 156892 149636 156893 149700
rect 156827 149635 156893 149636
rect 158486 148341 158546 198323
rect 159038 194037 159098 199819
rect 159294 196954 159914 198000
rect 159294 196718 159326 196954
rect 159562 196718 159646 196954
rect 159882 196718 159914 196954
rect 159294 196634 159914 196718
rect 159294 196398 159326 196634
rect 159562 196398 159646 196634
rect 159882 196398 159914 196634
rect 159035 194036 159101 194037
rect 159035 193972 159036 194036
rect 159100 193972 159101 194036
rect 159035 193971 159101 193972
rect 159294 160954 159914 196398
rect 161062 192949 161122 199819
rect 162166 196893 162226 199819
rect 162347 198252 162413 198253
rect 162347 198188 162348 198252
rect 162412 198188 162413 198252
rect 162347 198187 162413 198188
rect 162163 196892 162229 196893
rect 162163 196828 162164 196892
rect 162228 196828 162229 196892
rect 162163 196827 162229 196828
rect 161059 192948 161125 192949
rect 161059 192884 161060 192948
rect 161124 192884 161125 192948
rect 161059 192883 161125 192884
rect 159294 160718 159326 160954
rect 159562 160718 159646 160954
rect 159882 160718 159914 160954
rect 159294 160634 159914 160718
rect 159294 160398 159326 160634
rect 159562 160398 159646 160634
rect 159882 160398 159914 160634
rect 158483 148340 158549 148341
rect 158483 148276 158484 148340
rect 158548 148276 158549 148340
rect 158483 148275 158549 148276
rect 159294 142000 159914 160398
rect 162350 144669 162410 198187
rect 162534 197845 162594 199819
rect 163086 199749 163146 200499
rect 171179 200428 171245 200429
rect 171179 200364 171180 200428
rect 171244 200364 171245 200428
rect 171179 200363 171245 200364
rect 164187 199884 164253 199885
rect 164187 199820 164188 199884
rect 164252 199820 164253 199884
rect 164187 199819 164253 199820
rect 166763 199884 166829 199885
rect 166763 199820 166764 199884
rect 166828 199820 166829 199884
rect 166763 199819 166829 199820
rect 170443 199884 170509 199885
rect 170443 199820 170444 199884
rect 170508 199882 170509 199884
rect 170811 199884 170877 199885
rect 170508 199822 170690 199882
rect 170508 199820 170509 199822
rect 170443 199819 170509 199820
rect 163083 199748 163149 199749
rect 163083 199684 163084 199748
rect 163148 199684 163149 199748
rect 163083 199683 163149 199684
rect 162531 197844 162597 197845
rect 162531 197780 162532 197844
rect 162596 197780 162597 197844
rect 162531 197779 162597 197780
rect 164190 197165 164250 199819
rect 166211 199748 166277 199749
rect 166211 199684 166212 199748
rect 166276 199684 166277 199748
rect 166211 199683 166277 199684
rect 165475 198524 165541 198525
rect 165475 198460 165476 198524
rect 165540 198460 165541 198524
rect 165475 198459 165541 198460
rect 164187 197164 164253 197165
rect 164187 197100 164188 197164
rect 164252 197100 164253 197164
rect 164187 197099 164253 197100
rect 162347 144668 162413 144669
rect 162347 144604 162348 144668
rect 162412 144604 162413 144668
rect 162347 144603 162413 144604
rect 165478 141541 165538 198459
rect 166214 197981 166274 199683
rect 166766 198117 166826 199819
rect 169707 199748 169773 199749
rect 169707 199684 169708 199748
rect 169772 199684 169773 199748
rect 169707 199683 169773 199684
rect 166763 198116 166829 198117
rect 166763 198052 166764 198116
rect 166828 198052 166829 198116
rect 166763 198051 166829 198052
rect 166211 197980 166277 197981
rect 166211 197916 166212 197980
rect 166276 197916 166277 197980
rect 166211 197915 166277 197916
rect 169710 196485 169770 199683
rect 170443 198252 170509 198253
rect 170443 198188 170444 198252
rect 170508 198188 170509 198252
rect 170443 198187 170509 198188
rect 169707 196484 169773 196485
rect 169707 196420 169708 196484
rect 169772 196420 169773 196484
rect 169707 196419 169773 196420
rect 169523 196348 169589 196349
rect 169523 196284 169524 196348
rect 169588 196284 169589 196348
rect 169523 196283 169589 196284
rect 169339 195940 169405 195941
rect 169339 195876 169340 195940
rect 169404 195876 169405 195940
rect 169339 195875 169405 195876
rect 168235 193356 168301 193357
rect 168235 193292 168236 193356
rect 168300 193292 168301 193356
rect 168235 193291 168301 193292
rect 168238 156909 168298 193291
rect 168235 156908 168301 156909
rect 168235 156844 168236 156908
rect 168300 156844 168301 156908
rect 168235 156843 168301 156844
rect 169342 156773 169402 195875
rect 169339 156772 169405 156773
rect 169339 156708 169340 156772
rect 169404 156708 169405 156772
rect 169339 156707 169405 156708
rect 169526 151830 169586 196283
rect 170446 192813 170506 198187
rect 170443 192812 170509 192813
rect 170443 192748 170444 192812
rect 170508 192748 170509 192812
rect 170443 192747 170509 192748
rect 169526 151770 169770 151830
rect 165475 141540 165541 141541
rect 165475 141476 165476 141540
rect 165540 141476 165541 141540
rect 165475 141475 165541 141476
rect 169710 138685 169770 151770
rect 170630 148613 170690 199822
rect 170811 199820 170812 199884
rect 170876 199820 170877 199884
rect 170811 199819 170877 199820
rect 170814 196485 170874 199819
rect 171182 199613 171242 200363
rect 172283 200156 172349 200157
rect 172283 200092 172284 200156
rect 172348 200092 172349 200156
rect 172283 200091 172349 200092
rect 172835 200156 172901 200157
rect 172835 200092 172836 200156
rect 172900 200092 172901 200156
rect 172835 200091 172901 200092
rect 171179 199612 171245 199613
rect 171179 199548 171180 199612
rect 171244 199548 171245 199612
rect 171179 199547 171245 199548
rect 170995 198660 171061 198661
rect 170995 198596 170996 198660
rect 171060 198596 171061 198660
rect 170995 198595 171061 198596
rect 170811 196484 170877 196485
rect 170811 196420 170812 196484
rect 170876 196420 170877 196484
rect 170811 196419 170877 196420
rect 170998 192541 171058 198595
rect 172286 196485 172346 200091
rect 172651 199748 172717 199749
rect 172651 199684 172652 199748
rect 172716 199684 172717 199748
rect 172651 199683 172717 199684
rect 172283 196484 172349 196485
rect 172283 196420 172284 196484
rect 172348 196420 172349 196484
rect 172283 196419 172349 196420
rect 172654 193230 172714 199683
rect 172838 197845 172898 200091
rect 173574 199885 173634 200635
rect 176699 200020 176765 200021
rect 176699 199956 176700 200020
rect 176764 199956 176765 200020
rect 176699 199955 176765 199956
rect 173571 199884 173637 199885
rect 173571 199820 173572 199884
rect 173636 199820 173637 199884
rect 173571 199819 173637 199820
rect 173755 199884 173821 199885
rect 173755 199820 173756 199884
rect 173820 199820 173821 199884
rect 173755 199819 173821 199820
rect 174123 199884 174189 199885
rect 174123 199820 174124 199884
rect 174188 199820 174189 199884
rect 175227 199884 175293 199885
rect 175227 199882 175228 199884
rect 174123 199819 174189 199820
rect 174862 199822 175228 199882
rect 173387 199748 173453 199749
rect 173387 199684 173388 199748
rect 173452 199684 173453 199748
rect 173387 199683 173453 199684
rect 172835 197844 172901 197845
rect 172835 197780 172836 197844
rect 172900 197780 172901 197844
rect 172835 197779 172901 197780
rect 173390 195669 173450 199683
rect 173571 199612 173637 199613
rect 173571 199548 173572 199612
rect 173636 199548 173637 199612
rect 173571 199547 173637 199548
rect 173574 198389 173634 199547
rect 173758 199069 173818 199819
rect 173755 199068 173821 199069
rect 173755 199004 173756 199068
rect 173820 199004 173821 199068
rect 173755 199003 173821 199004
rect 174126 198797 174186 199819
rect 174123 198796 174189 198797
rect 174123 198732 174124 198796
rect 174188 198732 174189 198796
rect 174123 198731 174189 198732
rect 173571 198388 173637 198389
rect 173571 198324 173572 198388
rect 173636 198324 173637 198388
rect 173571 198323 173637 198324
rect 173755 196484 173821 196485
rect 173755 196420 173756 196484
rect 173820 196420 173821 196484
rect 173755 196419 173821 196420
rect 173387 195668 173453 195669
rect 173387 195604 173388 195668
rect 173452 195604 173453 195668
rect 173387 195603 173453 195604
rect 172470 193170 172714 193230
rect 172470 193085 172530 193170
rect 172467 193084 172533 193085
rect 172467 193020 172468 193084
rect 172532 193020 172533 193084
rect 172467 193019 172533 193020
rect 170995 192540 171061 192541
rect 170995 192476 170996 192540
rect 171060 192476 171061 192540
rect 170995 192475 171061 192476
rect 173758 148749 173818 196419
rect 174862 189821 174922 199822
rect 175227 199820 175228 199822
rect 175292 199820 175293 199884
rect 175227 199819 175293 199820
rect 176147 199884 176213 199885
rect 176147 199820 176148 199884
rect 176212 199820 176213 199884
rect 176147 199819 176213 199820
rect 175043 199748 175109 199749
rect 175043 199684 175044 199748
rect 175108 199684 175109 199748
rect 175043 199683 175109 199684
rect 174859 189820 174925 189821
rect 174859 189756 174860 189820
rect 174924 189756 174925 189820
rect 174859 189755 174925 189756
rect 175046 187373 175106 199683
rect 176150 198933 176210 199819
rect 176147 198932 176213 198933
rect 176147 198868 176148 198932
rect 176212 198868 176213 198932
rect 176147 198867 176213 198868
rect 176702 194610 176762 199955
rect 177435 199884 177501 199885
rect 177435 199820 177436 199884
rect 177500 199820 177501 199884
rect 177435 199819 177501 199820
rect 177438 198797 177498 199819
rect 177067 198796 177133 198797
rect 177067 198732 177068 198796
rect 177132 198732 177133 198796
rect 177067 198731 177133 198732
rect 177435 198796 177501 198797
rect 177435 198732 177436 198796
rect 177500 198732 177501 198796
rect 177435 198731 177501 198732
rect 176518 194550 176762 194610
rect 176518 189957 176578 194550
rect 176515 189956 176581 189957
rect 176515 189892 176516 189956
rect 176580 189892 176581 189956
rect 176515 189891 176581 189892
rect 175043 187372 175109 187373
rect 175043 187308 175044 187372
rect 175108 187308 175109 187372
rect 175043 187307 175109 187308
rect 177070 151469 177130 198731
rect 177294 178954 177914 198000
rect 181299 190092 181365 190093
rect 181299 190028 181300 190092
rect 181364 190028 181365 190092
rect 181299 190027 181365 190028
rect 177294 178718 177326 178954
rect 177562 178718 177646 178954
rect 177882 178718 177914 178954
rect 177294 178634 177914 178718
rect 177294 178398 177326 178634
rect 177562 178398 177646 178634
rect 177882 178398 177914 178634
rect 177067 151468 177133 151469
rect 177067 151404 177068 151468
rect 177132 151404 177133 151468
rect 177067 151403 177133 151404
rect 173755 148748 173821 148749
rect 173755 148684 173756 148748
rect 173820 148684 173821 148748
rect 173755 148683 173821 148684
rect 170627 148612 170693 148613
rect 170627 148548 170628 148612
rect 170692 148548 170693 148612
rect 170627 148547 170693 148548
rect 177294 142954 177914 178398
rect 177294 142718 177326 142954
rect 177562 142718 177646 142954
rect 177882 142718 177914 142954
rect 177294 142634 177914 142718
rect 177294 142398 177326 142634
rect 177562 142398 177646 142634
rect 177882 142398 177914 142634
rect 177294 142000 177914 142398
rect 146891 138684 146957 138685
rect 146891 138620 146892 138684
rect 146956 138620 146957 138684
rect 146891 138619 146957 138620
rect 169707 138684 169773 138685
rect 169707 138620 169708 138684
rect 169772 138620 169773 138684
rect 169707 138619 169773 138620
rect 128859 138548 128925 138549
rect 128859 138484 128860 138548
rect 128924 138484 128925 138548
rect 128859 138483 128925 138484
rect 181302 138005 181362 190027
rect 181794 183454 182414 198000
rect 186083 191044 186149 191045
rect 186083 190980 186084 191044
rect 186148 190980 186149 191044
rect 186083 190979 186149 190980
rect 181794 183218 181826 183454
rect 182062 183218 182146 183454
rect 182382 183218 182414 183454
rect 181794 183134 182414 183218
rect 181794 182898 181826 183134
rect 182062 182898 182146 183134
rect 182382 182898 182414 183134
rect 181794 147454 182414 182898
rect 181794 147218 181826 147454
rect 182062 147218 182146 147454
rect 182382 147218 182414 147454
rect 181794 147134 182414 147218
rect 181794 146898 181826 147134
rect 182062 146898 182146 147134
rect 182382 146898 182414 147134
rect 181794 142000 182414 146898
rect 185347 140180 185413 140181
rect 185347 140116 185348 140180
rect 185412 140116 185413 140180
rect 185347 140115 185413 140116
rect 185350 139093 185410 140115
rect 185899 139364 185965 139365
rect 185899 139300 185900 139364
rect 185964 139300 185965 139364
rect 185899 139299 185965 139300
rect 185347 139092 185413 139093
rect 185347 139028 185348 139092
rect 185412 139028 185413 139092
rect 185347 139027 185413 139028
rect 124811 138004 124877 138005
rect 124811 137940 124812 138004
rect 124876 137940 124877 138004
rect 124811 137939 124877 137940
rect 181299 138004 181365 138005
rect 181299 137940 181300 138004
rect 181364 137940 181365 138004
rect 181299 137939 181365 137940
rect 185902 137869 185962 139299
rect 185899 137868 185965 137869
rect 185899 137804 185900 137868
rect 185964 137804 185965 137868
rect 185899 137803 185965 137804
rect 186086 131749 186146 190979
rect 186294 187954 186914 198000
rect 187003 193220 187069 193221
rect 187003 193156 187004 193220
rect 187068 193156 187069 193220
rect 187003 193155 187069 193156
rect 186294 187718 186326 187954
rect 186562 187718 186646 187954
rect 186882 187718 186914 187954
rect 186294 187634 186914 187718
rect 186294 187398 186326 187634
rect 186562 187398 186646 187634
rect 186882 187398 186914 187634
rect 186294 151954 186914 187398
rect 186294 151718 186326 151954
rect 186562 151718 186646 151954
rect 186882 151718 186914 151954
rect 186294 151634 186914 151718
rect 186294 151398 186326 151634
rect 186562 151398 186646 151634
rect 186882 151398 186914 151634
rect 186294 142000 186914 151398
rect 186267 138956 186333 138957
rect 186267 138892 186268 138956
rect 186332 138892 186333 138956
rect 186267 138891 186333 138892
rect 186270 135965 186330 138891
rect 186451 138140 186517 138141
rect 186451 138076 186452 138140
rect 186516 138076 186517 138140
rect 186451 138075 186517 138076
rect 186267 135964 186333 135965
rect 186267 135900 186268 135964
rect 186332 135900 186333 135964
rect 186267 135899 186333 135900
rect 186083 131748 186149 131749
rect 186083 131684 186084 131748
rect 186148 131684 186149 131748
rect 186083 131683 186149 131684
rect 186267 131476 186333 131477
rect 186267 131412 186268 131476
rect 186332 131412 186333 131476
rect 186267 131411 186333 131412
rect 186270 128370 186330 131411
rect 186086 128310 186330 128370
rect 186086 122850 186146 128310
rect 186086 122790 186330 122850
rect 186083 118012 186149 118013
rect 186083 117948 186084 118012
rect 186148 117948 186149 118012
rect 186083 117947 186149 117948
rect 139568 115954 139888 115986
rect 139568 115718 139610 115954
rect 139846 115718 139888 115954
rect 139568 115634 139888 115718
rect 139568 115398 139610 115634
rect 139846 115398 139888 115634
rect 139568 115366 139888 115398
rect 170288 115954 170608 115986
rect 170288 115718 170330 115954
rect 170566 115718 170608 115954
rect 170288 115634 170608 115718
rect 170288 115398 170330 115634
rect 170566 115398 170608 115634
rect 170288 115366 170608 115398
rect 124208 111454 124528 111486
rect 124208 111218 124250 111454
rect 124486 111218 124528 111454
rect 124208 111134 124528 111218
rect 124208 110898 124250 111134
rect 124486 110898 124528 111134
rect 124208 110866 124528 110898
rect 154928 111454 155248 111486
rect 154928 111218 154970 111454
rect 155206 111218 155248 111454
rect 154928 111134 155248 111218
rect 154928 110898 154970 111134
rect 155206 110898 155248 111134
rect 154928 110866 155248 110898
rect 185648 111454 185968 111486
rect 185648 111218 185690 111454
rect 185926 111218 185968 111454
rect 185648 111134 185968 111218
rect 185648 110898 185690 111134
rect 185926 110898 185968 111134
rect 185648 110866 185968 110898
rect 186086 86325 186146 117947
rect 186270 104957 186330 122790
rect 186267 104956 186333 104957
rect 186267 104892 186268 104956
rect 186332 104892 186333 104956
rect 186267 104891 186333 104892
rect 186083 86324 186149 86325
rect 186083 86260 186084 86324
rect 186148 86260 186149 86324
rect 186083 86259 186149 86260
rect 123036 85990 123218 86050
rect 123036 85988 123037 85990
rect 122971 85987 123037 85988
rect 186083 82244 186149 82245
rect 186083 82180 186084 82244
rect 186148 82180 186149 82244
rect 186083 82179 186149 82180
rect 186086 81970 186146 82179
rect 186267 82108 186333 82109
rect 186267 82044 186268 82108
rect 186332 82044 186333 82108
rect 186267 82043 186333 82044
rect 185902 81910 186146 81970
rect 124075 81836 124141 81837
rect 124075 81772 124076 81836
rect 124140 81772 124141 81836
rect 124075 81771 124141 81772
rect 184059 81836 184125 81837
rect 184059 81772 184060 81836
rect 184124 81772 184125 81836
rect 184059 81771 184125 81772
rect 122603 69732 122669 69733
rect 122603 69668 122604 69732
rect 122668 69668 122669 69732
rect 122603 69667 122669 69668
rect 122419 68644 122485 68645
rect 122419 68580 122420 68644
rect 122484 68580 122485 68644
rect 122419 68579 122485 68580
rect 123294 52954 123914 78000
rect 124078 65925 124138 81771
rect 178907 81564 178973 81565
rect 178907 81500 178908 81564
rect 178972 81500 178973 81564
rect 178907 81499 178973 81500
rect 175043 81292 175109 81293
rect 175043 81228 175044 81292
rect 175108 81228 175109 81292
rect 175043 81227 175109 81228
rect 146339 81156 146405 81157
rect 146339 81092 146340 81156
rect 146404 81092 146405 81156
rect 146339 81091 146405 81092
rect 134011 79932 134077 79933
rect 134011 79868 134012 79932
rect 134076 79868 134077 79932
rect 134011 79867 134077 79868
rect 135115 79932 135181 79933
rect 135115 79868 135116 79932
rect 135180 79868 135181 79932
rect 135115 79867 135181 79868
rect 135483 79932 135549 79933
rect 135483 79868 135484 79932
rect 135548 79868 135549 79932
rect 135483 79867 135549 79868
rect 136035 79932 136101 79933
rect 136035 79868 136036 79932
rect 136100 79868 136101 79932
rect 136035 79867 136101 79868
rect 137507 79932 137573 79933
rect 137507 79868 137508 79932
rect 137572 79868 137573 79932
rect 137507 79867 137573 79868
rect 137691 79932 137757 79933
rect 137691 79868 137692 79932
rect 137756 79868 137757 79932
rect 137691 79867 137757 79868
rect 138059 79932 138125 79933
rect 138059 79868 138060 79932
rect 138124 79868 138125 79932
rect 138059 79867 138125 79868
rect 138427 79932 138493 79933
rect 138427 79868 138428 79932
rect 138492 79868 138493 79932
rect 138427 79867 138493 79868
rect 139163 79932 139229 79933
rect 139163 79868 139164 79932
rect 139228 79868 139229 79932
rect 139899 79932 139965 79933
rect 139899 79930 139900 79932
rect 139163 79867 139229 79868
rect 139718 79870 139900 79930
rect 133275 79796 133341 79797
rect 133275 79732 133276 79796
rect 133340 79732 133341 79796
rect 133275 79731 133341 79732
rect 133827 79796 133893 79797
rect 133827 79732 133828 79796
rect 133892 79732 133893 79796
rect 133827 79731 133893 79732
rect 124075 65924 124141 65925
rect 124075 65860 124076 65924
rect 124140 65860 124141 65924
rect 124075 65859 124141 65860
rect 123294 52718 123326 52954
rect 123562 52718 123646 52954
rect 123882 52718 123914 52954
rect 123294 52634 123914 52718
rect 123294 52398 123326 52634
rect 123562 52398 123646 52634
rect 123882 52398 123914 52634
rect 120579 31788 120645 31789
rect 120579 31724 120580 31788
rect 120644 31724 120645 31788
rect 120579 31723 120645 31724
rect 118794 12218 118826 12454
rect 119062 12218 119146 12454
rect 119382 12218 119414 12454
rect 118794 12134 119414 12218
rect 118794 11898 118826 12134
rect 119062 11898 119146 12134
rect 119382 11898 119414 12134
rect 118794 -2266 119414 11898
rect 118794 -2502 118826 -2266
rect 119062 -2502 119146 -2266
rect 119382 -2502 119414 -2266
rect 118794 -2586 119414 -2502
rect 118794 -2822 118826 -2586
rect 119062 -2822 119146 -2586
rect 119382 -2822 119414 -2586
rect 118794 -7654 119414 -2822
rect 123294 16954 123914 52398
rect 123294 16718 123326 16954
rect 123562 16718 123646 16954
rect 123882 16718 123914 16954
rect 123294 16634 123914 16718
rect 123294 16398 123326 16634
rect 123562 16398 123646 16634
rect 123882 16398 123914 16634
rect 123294 -3226 123914 16398
rect 123294 -3462 123326 -3226
rect 123562 -3462 123646 -3226
rect 123882 -3462 123914 -3226
rect 123294 -3546 123914 -3462
rect 123294 -3782 123326 -3546
rect 123562 -3782 123646 -3546
rect 123882 -3782 123914 -3546
rect 123294 -7654 123914 -3782
rect 127794 57454 128414 78000
rect 127794 57218 127826 57454
rect 128062 57218 128146 57454
rect 128382 57218 128414 57454
rect 127794 57134 128414 57218
rect 127794 56898 127826 57134
rect 128062 56898 128146 57134
rect 128382 56898 128414 57134
rect 127794 21454 128414 56898
rect 127794 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 128414 21454
rect 127794 21134 128414 21218
rect 127794 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 128414 21134
rect 127794 -4186 128414 20898
rect 127794 -4422 127826 -4186
rect 128062 -4422 128146 -4186
rect 128382 -4422 128414 -4186
rect 127794 -4506 128414 -4422
rect 127794 -4742 127826 -4506
rect 128062 -4742 128146 -4506
rect 128382 -4742 128414 -4506
rect 127794 -7654 128414 -4742
rect 132294 61954 132914 78000
rect 133091 74628 133157 74629
rect 133091 74564 133092 74628
rect 133156 74564 133157 74628
rect 133091 74563 133157 74564
rect 132294 61718 132326 61954
rect 132562 61718 132646 61954
rect 132882 61718 132914 61954
rect 132294 61634 132914 61718
rect 132294 61398 132326 61634
rect 132562 61398 132646 61634
rect 132882 61398 132914 61634
rect 132294 25954 132914 61398
rect 133094 56541 133154 74563
rect 133278 60621 133338 79731
rect 133459 76668 133525 76669
rect 133459 76604 133460 76668
rect 133524 76604 133525 76668
rect 133459 76603 133525 76604
rect 133462 63477 133522 76603
rect 133459 63476 133525 63477
rect 133459 63412 133460 63476
rect 133524 63412 133525 63476
rect 133459 63411 133525 63412
rect 133275 60620 133341 60621
rect 133275 60556 133276 60620
rect 133340 60556 133341 60620
rect 133275 60555 133341 60556
rect 133091 56540 133157 56541
rect 133091 56476 133092 56540
rect 133156 56476 133157 56540
rect 133091 56475 133157 56476
rect 133830 49605 133890 79731
rect 134014 50965 134074 79867
rect 134379 78028 134445 78029
rect 134379 77964 134380 78028
rect 134444 77964 134445 78028
rect 134379 77963 134445 77964
rect 134195 76668 134261 76669
rect 134195 76604 134196 76668
rect 134260 76604 134261 76668
rect 134195 76603 134261 76604
rect 134198 57901 134258 76603
rect 134382 62117 134442 77963
rect 135118 75853 135178 79867
rect 135299 77076 135365 77077
rect 135299 77012 135300 77076
rect 135364 77012 135365 77076
rect 135299 77011 135365 77012
rect 135115 75852 135181 75853
rect 135115 75788 135116 75852
rect 135180 75788 135181 75852
rect 135115 75787 135181 75788
rect 134379 62116 134445 62117
rect 134379 62052 134380 62116
rect 134444 62052 134445 62116
rect 134379 62051 134445 62052
rect 134195 57900 134261 57901
rect 134195 57836 134196 57900
rect 134260 57836 134261 57900
rect 134195 57835 134261 57836
rect 134011 50964 134077 50965
rect 134011 50900 134012 50964
rect 134076 50900 134077 50964
rect 134011 50899 134077 50900
rect 133827 49604 133893 49605
rect 133827 49540 133828 49604
rect 133892 49540 133893 49604
rect 133827 49539 133893 49540
rect 135302 46885 135362 77011
rect 135486 48245 135546 79867
rect 135667 79796 135733 79797
rect 135667 79732 135668 79796
rect 135732 79732 135733 79796
rect 135667 79731 135733 79732
rect 135670 53821 135730 79731
rect 136038 74765 136098 79867
rect 136587 79660 136653 79661
rect 136587 79596 136588 79660
rect 136652 79596 136653 79660
rect 136587 79595 136653 79596
rect 136035 74764 136101 74765
rect 136035 74700 136036 74764
rect 136100 74700 136101 74764
rect 136035 74699 136101 74700
rect 135667 53820 135733 53821
rect 135667 53756 135668 53820
rect 135732 53756 135733 53820
rect 135667 53755 135733 53756
rect 135483 48244 135549 48245
rect 135483 48180 135484 48244
rect 135548 48180 135549 48244
rect 135483 48179 135549 48180
rect 135299 46884 135365 46885
rect 135299 46820 135300 46884
rect 135364 46820 135365 46884
rect 135299 46819 135365 46820
rect 136590 44165 136650 79595
rect 136794 66454 137414 78000
rect 136794 66218 136826 66454
rect 137062 66218 137146 66454
rect 137382 66218 137414 66454
rect 136794 66134 137414 66218
rect 136794 65898 136826 66134
rect 137062 65898 137146 66134
rect 137382 65898 137414 66134
rect 136587 44164 136653 44165
rect 136587 44100 136588 44164
rect 136652 44100 136653 44164
rect 136587 44099 136653 44100
rect 132294 25718 132326 25954
rect 132562 25718 132646 25954
rect 132882 25718 132914 25954
rect 132294 25634 132914 25718
rect 132294 25398 132326 25634
rect 132562 25398 132646 25634
rect 132882 25398 132914 25634
rect 132294 -5146 132914 25398
rect 132294 -5382 132326 -5146
rect 132562 -5382 132646 -5146
rect 132882 -5382 132914 -5146
rect 132294 -5466 132914 -5382
rect 132294 -5702 132326 -5466
rect 132562 -5702 132646 -5466
rect 132882 -5702 132914 -5466
rect 132294 -7654 132914 -5702
rect 136794 30454 137414 65898
rect 137510 55045 137570 79867
rect 137694 75717 137754 79867
rect 138062 77077 138122 79867
rect 138243 79796 138309 79797
rect 138243 79732 138244 79796
rect 138308 79732 138309 79796
rect 138243 79731 138309 79732
rect 138059 77076 138125 77077
rect 138059 77012 138060 77076
rect 138124 77012 138125 77076
rect 138059 77011 138125 77012
rect 138059 76668 138125 76669
rect 138059 76604 138060 76668
rect 138124 76604 138125 76668
rect 138059 76603 138125 76604
rect 137691 75716 137757 75717
rect 137691 75652 137692 75716
rect 137756 75652 137757 75716
rect 137691 75651 137757 75652
rect 138062 55181 138122 76603
rect 138246 57765 138306 79731
rect 138430 60485 138490 79867
rect 138611 77076 138677 77077
rect 138611 77012 138612 77076
rect 138676 77012 138677 77076
rect 138611 77011 138677 77012
rect 138614 61981 138674 77011
rect 139166 76669 139226 79867
rect 139163 76668 139229 76669
rect 139163 76604 139164 76668
rect 139228 76604 139229 76668
rect 139163 76603 139229 76604
rect 139347 76668 139413 76669
rect 139347 76604 139348 76668
rect 139412 76604 139413 76668
rect 139347 76603 139413 76604
rect 138611 61980 138677 61981
rect 138611 61916 138612 61980
rect 138676 61916 138677 61980
rect 138611 61915 138677 61916
rect 138427 60484 138493 60485
rect 138427 60420 138428 60484
rect 138492 60420 138493 60484
rect 138427 60419 138493 60420
rect 138243 57764 138309 57765
rect 138243 57700 138244 57764
rect 138308 57700 138309 57764
rect 138243 57699 138309 57700
rect 138059 55180 138125 55181
rect 138059 55116 138060 55180
rect 138124 55116 138125 55180
rect 138059 55115 138125 55116
rect 137507 55044 137573 55045
rect 137507 54980 137508 55044
rect 137572 54980 137573 55044
rect 137507 54979 137573 54980
rect 139350 50829 139410 76603
rect 139531 76532 139597 76533
rect 139531 76468 139532 76532
rect 139596 76468 139597 76532
rect 139531 76467 139597 76468
rect 139534 53685 139594 76467
rect 139718 59125 139778 79870
rect 139899 79868 139900 79870
rect 139964 79868 139965 79932
rect 139899 79867 139965 79868
rect 141555 79932 141621 79933
rect 141555 79868 141556 79932
rect 141620 79868 141621 79932
rect 141555 79867 141621 79868
rect 142659 79932 142725 79933
rect 142659 79868 142660 79932
rect 142724 79868 142725 79932
rect 142659 79867 142725 79868
rect 144131 79932 144197 79933
rect 144131 79868 144132 79932
rect 144196 79868 144197 79932
rect 145603 79932 145669 79933
rect 145603 79930 145604 79932
rect 144131 79867 144197 79868
rect 145422 79870 145604 79930
rect 139899 79796 139965 79797
rect 139899 79732 139900 79796
rect 139964 79732 139965 79796
rect 139899 79731 139965 79732
rect 140267 79796 140333 79797
rect 140267 79732 140268 79796
rect 140332 79732 140333 79796
rect 140267 79731 140333 79732
rect 140819 79796 140885 79797
rect 140819 79732 140820 79796
rect 140884 79732 140885 79796
rect 140819 79731 140885 79732
rect 139902 59261 139962 79731
rect 140270 76533 140330 79731
rect 140267 76532 140333 76533
rect 140267 76468 140268 76532
rect 140332 76468 140333 76532
rect 140267 76467 140333 76468
rect 139899 59260 139965 59261
rect 139899 59196 139900 59260
rect 139964 59196 139965 59260
rect 139899 59195 139965 59196
rect 139715 59124 139781 59125
rect 139715 59060 139716 59124
rect 139780 59060 139781 59124
rect 139715 59059 139781 59060
rect 140822 58581 140882 79731
rect 141003 79660 141069 79661
rect 141003 79596 141004 79660
rect 141068 79596 141069 79660
rect 141003 79595 141069 79596
rect 141006 68917 141066 79595
rect 141558 78437 141618 79867
rect 142107 79796 142173 79797
rect 142107 79732 142108 79796
rect 142172 79732 142173 79796
rect 142107 79731 142173 79732
rect 141555 78436 141621 78437
rect 141555 78372 141556 78436
rect 141620 78372 141621 78436
rect 141555 78371 141621 78372
rect 141294 70954 141914 78000
rect 142110 77485 142170 79731
rect 142662 78709 142722 79867
rect 143579 79796 143645 79797
rect 143579 79732 143580 79796
rect 143644 79732 143645 79796
rect 143579 79731 143645 79732
rect 142659 78708 142725 78709
rect 142659 78644 142660 78708
rect 142724 78644 142725 78708
rect 142659 78643 142725 78644
rect 143582 77757 143642 79731
rect 143947 77892 144013 77893
rect 143947 77828 143948 77892
rect 144012 77828 144013 77892
rect 143947 77827 144013 77828
rect 143579 77756 143645 77757
rect 143579 77692 143580 77756
rect 143644 77692 143645 77756
rect 143579 77691 143645 77692
rect 142107 77484 142173 77485
rect 142107 77420 142108 77484
rect 142172 77420 142173 77484
rect 142107 77419 142173 77420
rect 143579 76668 143645 76669
rect 143579 76604 143580 76668
rect 143644 76604 143645 76668
rect 143579 76603 143645 76604
rect 141294 70718 141326 70954
rect 141562 70718 141646 70954
rect 141882 70718 141914 70954
rect 141294 70634 141914 70718
rect 141294 70398 141326 70634
rect 141562 70398 141646 70634
rect 141882 70398 141914 70634
rect 141003 68916 141069 68917
rect 141003 68852 141004 68916
rect 141068 68852 141069 68916
rect 141003 68851 141069 68852
rect 140819 58580 140885 58581
rect 140819 58516 140820 58580
rect 140884 58516 140885 58580
rect 140819 58515 140885 58516
rect 139531 53684 139597 53685
rect 139531 53620 139532 53684
rect 139596 53620 139597 53684
rect 139531 53619 139597 53620
rect 139347 50828 139413 50829
rect 139347 50764 139348 50828
rect 139412 50764 139413 50828
rect 139347 50763 139413 50764
rect 136794 30218 136826 30454
rect 137062 30218 137146 30454
rect 137382 30218 137414 30454
rect 136794 30134 137414 30218
rect 136794 29898 136826 30134
rect 137062 29898 137146 30134
rect 137382 29898 137414 30134
rect 136794 -6106 137414 29898
rect 136794 -6342 136826 -6106
rect 137062 -6342 137146 -6106
rect 137382 -6342 137414 -6106
rect 136794 -6426 137414 -6342
rect 136794 -6662 136826 -6426
rect 137062 -6662 137146 -6426
rect 137382 -6662 137414 -6426
rect 136794 -7654 137414 -6662
rect 141294 34954 141914 70398
rect 143582 67557 143642 76603
rect 143763 74764 143829 74765
rect 143763 74700 143764 74764
rect 143828 74700 143829 74764
rect 143763 74699 143829 74700
rect 143766 68101 143826 74699
rect 143950 68509 144010 77827
rect 144134 71773 144194 79867
rect 145422 72997 145482 79870
rect 145603 79868 145604 79870
rect 145668 79868 145669 79932
rect 145603 79867 145669 79868
rect 146342 79525 146402 81091
rect 149283 81020 149349 81021
rect 149283 80956 149284 81020
rect 149348 80956 149349 81020
rect 149283 80955 149349 80956
rect 148731 80884 148797 80885
rect 148731 80820 148732 80884
rect 148796 80820 148797 80884
rect 148731 80819 148797 80820
rect 146523 80204 146589 80205
rect 146523 80140 146524 80204
rect 146588 80140 146589 80204
rect 146523 80139 146589 80140
rect 146339 79524 146405 79525
rect 146339 79460 146340 79524
rect 146404 79460 146405 79524
rect 146339 79459 146405 79460
rect 145603 76668 145669 76669
rect 145603 76604 145604 76668
rect 145668 76604 145669 76668
rect 145603 76603 145669 76604
rect 145419 72996 145485 72997
rect 145419 72932 145420 72996
rect 145484 72932 145485 72996
rect 145419 72931 145485 72932
rect 144131 71772 144197 71773
rect 144131 71708 144132 71772
rect 144196 71708 144197 71772
rect 144131 71707 144197 71708
rect 143947 68508 144013 68509
rect 143947 68444 143948 68508
rect 144012 68444 144013 68508
rect 143947 68443 144013 68444
rect 143763 68100 143829 68101
rect 143763 68036 143764 68100
rect 143828 68036 143829 68100
rect 143763 68035 143829 68036
rect 143579 67556 143645 67557
rect 143579 67492 143580 67556
rect 143644 67492 143645 67556
rect 143579 67491 143645 67492
rect 141294 34718 141326 34954
rect 141562 34718 141646 34954
rect 141882 34718 141914 34954
rect 141294 34634 141914 34718
rect 141294 34398 141326 34634
rect 141562 34398 141646 34634
rect 141882 34398 141914 34634
rect 141294 -7066 141914 34398
rect 144134 10301 144194 71707
rect 144499 68508 144565 68509
rect 144499 68444 144500 68508
rect 144564 68444 144565 68508
rect 144499 68443 144565 68444
rect 144315 68100 144381 68101
rect 144315 68036 144316 68100
rect 144380 68036 144381 68100
rect 144315 68035 144381 68036
rect 144318 28253 144378 68035
rect 144502 37909 144562 68443
rect 144683 67556 144749 67557
rect 144683 67492 144684 67556
rect 144748 67492 144749 67556
rect 144683 67491 144749 67492
rect 144686 51781 144746 67491
rect 144683 51780 144749 51781
rect 144683 51716 144684 51780
rect 144748 51716 144749 51780
rect 144683 51715 144749 51716
rect 144499 37908 144565 37909
rect 144499 37844 144500 37908
rect 144564 37844 144565 37908
rect 144499 37843 144565 37844
rect 145422 35189 145482 72931
rect 145606 68237 145666 76603
rect 145794 75454 146414 78000
rect 145794 75218 145826 75454
rect 146062 75218 146146 75454
rect 146382 75218 146414 75454
rect 145794 75134 146414 75218
rect 145794 74898 145826 75134
rect 146062 74898 146146 75134
rect 146382 74898 146414 75134
rect 145603 68236 145669 68237
rect 145603 68172 145604 68236
rect 145668 68172 145669 68236
rect 145603 68171 145669 68172
rect 145794 39454 146414 74898
rect 146526 70277 146586 80139
rect 148734 79933 148794 80819
rect 149286 79933 149346 80955
rect 155723 80204 155789 80205
rect 155723 80140 155724 80204
rect 155788 80140 155789 80204
rect 155723 80139 155789 80140
rect 170811 80204 170877 80205
rect 170811 80140 170812 80204
rect 170876 80140 170877 80204
rect 170811 80139 170877 80140
rect 146891 79932 146957 79933
rect 146891 79868 146892 79932
rect 146956 79868 146957 79932
rect 146891 79867 146957 79868
rect 147627 79932 147693 79933
rect 147627 79868 147628 79932
rect 147692 79868 147693 79932
rect 147627 79867 147693 79868
rect 148731 79932 148797 79933
rect 148731 79868 148732 79932
rect 148796 79868 148797 79932
rect 148731 79867 148797 79868
rect 149283 79932 149349 79933
rect 149283 79868 149284 79932
rect 149348 79868 149349 79932
rect 149283 79867 149349 79868
rect 149835 79932 149901 79933
rect 149835 79868 149836 79932
rect 149900 79868 149901 79932
rect 149835 79867 149901 79868
rect 151675 79932 151741 79933
rect 151675 79868 151676 79932
rect 151740 79868 151741 79932
rect 151675 79867 151741 79868
rect 153147 79932 153213 79933
rect 153147 79868 153148 79932
rect 153212 79868 153213 79932
rect 154435 79932 154501 79933
rect 154435 79930 154436 79932
rect 153147 79867 153213 79868
rect 154254 79870 154436 79930
rect 146894 78709 146954 79867
rect 147075 79796 147141 79797
rect 147075 79732 147076 79796
rect 147140 79732 147141 79796
rect 147075 79731 147141 79732
rect 146891 78708 146957 78709
rect 146891 78644 146892 78708
rect 146956 78644 146957 78708
rect 146891 78643 146957 78644
rect 146707 76668 146773 76669
rect 146707 76604 146708 76668
rect 146772 76604 146773 76668
rect 146707 76603 146773 76604
rect 146523 70276 146589 70277
rect 146523 70212 146524 70276
rect 146588 70212 146589 70276
rect 146523 70211 146589 70212
rect 146526 64890 146586 70211
rect 146710 69597 146770 76603
rect 147078 74221 147138 79731
rect 147630 77310 147690 79867
rect 147995 79796 148061 79797
rect 147995 79732 147996 79796
rect 148060 79732 148061 79796
rect 147995 79731 148061 79732
rect 147446 77250 147690 77310
rect 147811 77348 147877 77349
rect 147811 77284 147812 77348
rect 147876 77284 147877 77348
rect 147811 77283 147877 77284
rect 147075 74220 147141 74221
rect 147075 74156 147076 74220
rect 147140 74156 147141 74220
rect 147075 74155 147141 74156
rect 146707 69596 146773 69597
rect 146707 69532 146708 69596
rect 146772 69532 146773 69596
rect 146707 69531 146773 69532
rect 146526 64830 146954 64890
rect 146894 46205 146954 64830
rect 147078 50285 147138 74155
rect 147446 72725 147506 77250
rect 147443 72724 147509 72725
rect 147443 72660 147444 72724
rect 147508 72660 147509 72724
rect 147443 72659 147509 72660
rect 147259 69596 147325 69597
rect 147259 69532 147260 69596
rect 147324 69532 147325 69596
rect 147259 69531 147325 69532
rect 147262 57221 147322 69531
rect 147446 64157 147506 72659
rect 147814 67421 147874 77283
rect 147811 67420 147877 67421
rect 147811 67356 147812 67420
rect 147876 67356 147877 67420
rect 147811 67355 147877 67356
rect 147998 67285 148058 79731
rect 148734 79389 148794 79867
rect 148731 79388 148797 79389
rect 148731 79324 148732 79388
rect 148796 79324 148797 79388
rect 148731 79323 148797 79324
rect 149099 79388 149165 79389
rect 149099 79324 149100 79388
rect 149164 79324 149165 79388
rect 149099 79323 149165 79324
rect 148915 77484 148981 77485
rect 148915 77420 148916 77484
rect 148980 77420 148981 77484
rect 148915 77419 148981 77420
rect 148363 77212 148429 77213
rect 148363 77148 148364 77212
rect 148428 77148 148429 77212
rect 148363 77147 148429 77148
rect 148366 72861 148426 77147
rect 148363 72860 148429 72861
rect 148363 72796 148364 72860
rect 148428 72796 148429 72860
rect 148363 72795 148429 72796
rect 148366 70410 148426 72795
rect 148366 70350 148610 70410
rect 148179 67420 148245 67421
rect 148179 67356 148180 67420
rect 148244 67356 148245 67420
rect 148179 67355 148245 67356
rect 147995 67284 148061 67285
rect 147995 67220 147996 67284
rect 148060 67220 148061 67284
rect 147995 67219 148061 67220
rect 147443 64156 147509 64157
rect 147443 64092 147444 64156
rect 147508 64092 147509 64156
rect 147443 64091 147509 64092
rect 147259 57220 147325 57221
rect 147259 57156 147260 57220
rect 147324 57156 147325 57220
rect 147259 57155 147325 57156
rect 147075 50284 147141 50285
rect 147075 50220 147076 50284
rect 147140 50220 147141 50284
rect 147075 50219 147141 50220
rect 146891 46204 146957 46205
rect 146891 46140 146892 46204
rect 146956 46140 146957 46204
rect 146891 46139 146957 46140
rect 145794 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 146414 39454
rect 145794 39134 146414 39218
rect 145794 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 146414 39134
rect 145419 35188 145485 35189
rect 145419 35124 145420 35188
rect 145484 35124 145485 35188
rect 145419 35123 145485 35124
rect 144315 28252 144381 28253
rect 144315 28188 144316 28252
rect 144380 28188 144381 28252
rect 144315 28187 144381 28188
rect 144131 10300 144197 10301
rect 144131 10236 144132 10300
rect 144196 10236 144197 10300
rect 144131 10235 144197 10236
rect 141294 -7302 141326 -7066
rect 141562 -7302 141646 -7066
rect 141882 -7302 141914 -7066
rect 141294 -7386 141914 -7302
rect 141294 -7622 141326 -7386
rect 141562 -7622 141646 -7386
rect 141882 -7622 141914 -7386
rect 141294 -7654 141914 -7622
rect 145794 3454 146414 38898
rect 148182 8941 148242 67355
rect 148363 67284 148429 67285
rect 148363 67220 148364 67284
rect 148428 67220 148429 67284
rect 148363 67219 148429 67220
rect 148366 43893 148426 67219
rect 148550 62933 148610 70350
rect 148918 66877 148978 77419
rect 149102 74550 149162 79323
rect 149286 78573 149346 79867
rect 149651 79660 149717 79661
rect 149651 79596 149652 79660
rect 149716 79596 149717 79660
rect 149651 79595 149717 79596
rect 149283 78572 149349 78573
rect 149283 78508 149284 78572
rect 149348 78508 149349 78572
rect 149283 78507 149349 78508
rect 149102 74490 149530 74550
rect 149470 73949 149530 74490
rect 149654 74221 149714 79595
rect 149651 74220 149717 74221
rect 149651 74156 149652 74220
rect 149716 74156 149717 74220
rect 149651 74155 149717 74156
rect 149467 73948 149533 73949
rect 149467 73884 149468 73948
rect 149532 73884 149533 73948
rect 149467 73883 149533 73884
rect 149838 68917 149898 79867
rect 150019 77348 150085 77349
rect 150019 77284 150020 77348
rect 150084 77284 150085 77348
rect 150019 77283 150085 77284
rect 149835 68916 149901 68917
rect 149835 68852 149836 68916
rect 149900 68852 149901 68916
rect 149835 68851 149901 68852
rect 150022 67013 150082 77283
rect 150019 67012 150085 67013
rect 150019 66948 150020 67012
rect 150084 66948 150085 67012
rect 150019 66947 150085 66948
rect 148915 66876 148981 66877
rect 148915 66812 148916 66876
rect 148980 66812 148981 66876
rect 148915 66811 148981 66812
rect 148547 62932 148613 62933
rect 148547 62868 148548 62932
rect 148612 62868 148613 62932
rect 148547 62867 148613 62868
rect 150294 43954 150914 78000
rect 151123 77348 151189 77349
rect 151123 77284 151124 77348
rect 151188 77284 151189 77348
rect 151123 77283 151189 77284
rect 151126 73541 151186 77283
rect 151123 73540 151189 73541
rect 151123 73476 151124 73540
rect 151188 73476 151189 73540
rect 151123 73475 151189 73476
rect 151678 73405 151738 79867
rect 152595 79660 152661 79661
rect 152595 79596 152596 79660
rect 152660 79596 152661 79660
rect 152595 79595 152661 79596
rect 152411 78708 152477 78709
rect 152411 78644 152412 78708
rect 152476 78644 152477 78708
rect 152411 78643 152477 78644
rect 151675 73404 151741 73405
rect 151675 73340 151676 73404
rect 151740 73340 151741 73404
rect 151675 73339 151741 73340
rect 152414 50965 152474 78643
rect 152598 77349 152658 79595
rect 152779 79252 152845 79253
rect 152779 79188 152780 79252
rect 152844 79188 152845 79252
rect 152779 79187 152845 79188
rect 152595 77348 152661 77349
rect 152595 77284 152596 77348
rect 152660 77284 152661 77348
rect 152595 77283 152661 77284
rect 152782 64429 152842 79187
rect 153150 74085 153210 79867
rect 153883 79524 153949 79525
rect 153883 79460 153884 79524
rect 153948 79460 153949 79524
rect 153883 79459 153949 79460
rect 153147 74084 153213 74085
rect 153147 74020 153148 74084
rect 153212 74020 153213 74084
rect 153147 74019 153213 74020
rect 152779 64428 152845 64429
rect 152779 64364 152780 64428
rect 152844 64364 152845 64428
rect 152779 64363 152845 64364
rect 153886 59261 153946 79459
rect 154067 77348 154133 77349
rect 154067 77284 154068 77348
rect 154132 77284 154133 77348
rect 154067 77283 154133 77284
rect 153883 59260 153949 59261
rect 153883 59196 153884 59260
rect 153948 59196 153949 59260
rect 153883 59195 153949 59196
rect 154070 56269 154130 77283
rect 154067 56268 154133 56269
rect 154067 56204 154068 56268
rect 154132 56204 154133 56268
rect 154067 56203 154133 56204
rect 152411 50964 152477 50965
rect 152411 50900 152412 50964
rect 152476 50900 152477 50964
rect 152411 50899 152477 50900
rect 154254 45525 154314 79870
rect 154435 79868 154436 79870
rect 154500 79868 154501 79932
rect 154435 79867 154501 79868
rect 154987 79932 155053 79933
rect 154987 79868 154988 79932
rect 155052 79868 155053 79932
rect 154987 79867 155053 79868
rect 154990 78165 155050 79867
rect 154987 78164 155053 78165
rect 154987 78100 154988 78164
rect 155052 78100 155053 78164
rect 154987 78099 155053 78100
rect 154435 77484 154501 77485
rect 154435 77420 154436 77484
rect 154500 77420 154501 77484
rect 154435 77419 154501 77420
rect 154251 45524 154317 45525
rect 154251 45460 154252 45524
rect 154316 45460 154317 45524
rect 154251 45459 154317 45460
rect 148363 43892 148429 43893
rect 148363 43828 148364 43892
rect 148428 43828 148429 43892
rect 148363 43827 148429 43828
rect 150294 43718 150326 43954
rect 150562 43718 150646 43954
rect 150882 43718 150914 43954
rect 150294 43634 150914 43718
rect 150294 43398 150326 43634
rect 150562 43398 150646 43634
rect 150882 43398 150914 43634
rect 148179 8940 148245 8941
rect 148179 8876 148180 8940
rect 148244 8876 148245 8940
rect 148179 8875 148245 8876
rect 145794 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 146414 3454
rect 145794 3134 146414 3218
rect 145794 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 146414 3134
rect 145794 -346 146414 2898
rect 145794 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 146414 -346
rect 145794 -666 146414 -582
rect 145794 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 146414 -666
rect 145794 -7654 146414 -902
rect 150294 7954 150914 43398
rect 154438 38589 154498 77419
rect 154794 48454 155414 78000
rect 155539 77348 155605 77349
rect 155539 77284 155540 77348
rect 155604 77284 155605 77348
rect 155539 77283 155605 77284
rect 154794 48218 154826 48454
rect 155062 48218 155146 48454
rect 155382 48218 155414 48454
rect 154794 48134 155414 48218
rect 154794 47898 154826 48134
rect 155062 47898 155146 48134
rect 155382 47898 155414 48134
rect 154435 38588 154501 38589
rect 154435 38524 154436 38588
rect 154500 38524 154501 38588
rect 154435 38523 154501 38524
rect 150294 7718 150326 7954
rect 150562 7718 150646 7954
rect 150882 7718 150914 7954
rect 150294 7634 150914 7718
rect 150294 7398 150326 7634
rect 150562 7398 150646 7634
rect 150882 7398 150914 7634
rect 150294 -1306 150914 7398
rect 150294 -1542 150326 -1306
rect 150562 -1542 150646 -1306
rect 150882 -1542 150914 -1306
rect 150294 -1626 150914 -1542
rect 150294 -1862 150326 -1626
rect 150562 -1862 150646 -1626
rect 150882 -1862 150914 -1626
rect 150294 -7654 150914 -1862
rect 154794 12454 155414 47898
rect 155542 42805 155602 77283
rect 155539 42804 155605 42805
rect 155539 42740 155540 42804
rect 155604 42740 155605 42804
rect 155539 42739 155605 42740
rect 155726 20637 155786 80139
rect 159035 80068 159101 80069
rect 159035 80004 159036 80068
rect 159100 80004 159101 80068
rect 159035 80003 159101 80004
rect 169523 80068 169589 80069
rect 169523 80004 169524 80068
rect 169588 80004 169589 80068
rect 169523 80003 169589 80004
rect 155907 79932 155973 79933
rect 155907 79868 155908 79932
rect 155972 79868 155973 79932
rect 155907 79867 155973 79868
rect 156643 79932 156709 79933
rect 156643 79868 156644 79932
rect 156708 79868 156709 79932
rect 156643 79867 156709 79868
rect 158115 79932 158181 79933
rect 158115 79868 158116 79932
rect 158180 79930 158181 79932
rect 158483 79932 158549 79933
rect 158180 79870 158362 79930
rect 158180 79868 158181 79870
rect 158115 79867 158181 79868
rect 155910 76941 155970 79867
rect 155907 76940 155973 76941
rect 155907 76876 155908 76940
rect 155972 76876 155973 76940
rect 155907 76875 155973 76876
rect 156646 52189 156706 79867
rect 156827 79796 156893 79797
rect 156827 79732 156828 79796
rect 156892 79732 156893 79796
rect 156827 79731 156893 79732
rect 156643 52188 156709 52189
rect 156643 52124 156644 52188
rect 156708 52124 156709 52188
rect 156643 52123 156709 52124
rect 156830 44029 156890 79731
rect 157195 79660 157261 79661
rect 157195 79596 157196 79660
rect 157260 79596 157261 79660
rect 157195 79595 157261 79596
rect 157011 78572 157077 78573
rect 157011 78508 157012 78572
rect 157076 78508 157077 78572
rect 157011 78507 157077 78508
rect 156827 44028 156893 44029
rect 156827 43964 156828 44028
rect 156892 43964 156893 44028
rect 156827 43963 156893 43964
rect 157014 28933 157074 78507
rect 157011 28932 157077 28933
rect 157011 28868 157012 28932
rect 157076 28868 157077 28932
rect 157011 28867 157077 28868
rect 157198 24853 157258 79595
rect 158115 78980 158181 78981
rect 158115 78916 158116 78980
rect 158180 78916 158181 78980
rect 158115 78915 158181 78916
rect 158118 50829 158178 78915
rect 158115 50828 158181 50829
rect 158115 50764 158116 50828
rect 158180 50764 158181 50828
rect 158115 50763 158181 50764
rect 157195 24852 157261 24853
rect 157195 24788 157196 24852
rect 157260 24788 157261 24852
rect 157195 24787 157261 24788
rect 158302 21861 158362 79870
rect 158483 79868 158484 79932
rect 158548 79868 158549 79932
rect 158483 79867 158549 79868
rect 158486 21997 158546 79867
rect 158667 79796 158733 79797
rect 158667 79732 158668 79796
rect 158732 79732 158733 79796
rect 158667 79731 158733 79732
rect 158670 73133 158730 79731
rect 158851 78572 158917 78573
rect 158851 78508 158852 78572
rect 158916 78508 158917 78572
rect 158851 78507 158917 78508
rect 158667 73132 158733 73133
rect 158667 73068 158668 73132
rect 158732 73068 158733 73132
rect 158667 73067 158733 73068
rect 158854 57901 158914 78507
rect 158851 57900 158917 57901
rect 158851 57836 158852 57900
rect 158916 57836 158917 57900
rect 158851 57835 158917 57836
rect 159038 52325 159098 80003
rect 159403 79932 159469 79933
rect 159403 79868 159404 79932
rect 159468 79868 159469 79932
rect 159403 79867 159469 79868
rect 161059 79932 161125 79933
rect 161059 79868 161060 79932
rect 161124 79868 161125 79932
rect 161059 79867 161125 79868
rect 161979 79932 162045 79933
rect 161979 79868 161980 79932
rect 162044 79868 162045 79932
rect 161979 79867 162045 79868
rect 162347 79932 162413 79933
rect 162347 79868 162348 79932
rect 162412 79868 162413 79932
rect 162347 79867 162413 79868
rect 162899 79932 162965 79933
rect 162899 79868 162900 79932
rect 162964 79868 162965 79932
rect 162899 79867 162965 79868
rect 166211 79932 166277 79933
rect 166211 79868 166212 79932
rect 166276 79868 166277 79932
rect 166211 79867 166277 79868
rect 166579 79932 166645 79933
rect 166579 79868 166580 79932
rect 166644 79868 166645 79932
rect 166579 79867 166645 79868
rect 169339 79932 169405 79933
rect 169339 79868 169340 79932
rect 169404 79868 169405 79932
rect 169339 79867 169405 79868
rect 159406 78709 159466 79867
rect 159403 78708 159469 78709
rect 159403 78644 159404 78708
rect 159468 78644 159469 78708
rect 159403 78643 159469 78644
rect 160691 78708 160757 78709
rect 160691 78644 160692 78708
rect 160756 78644 160757 78708
rect 160691 78643 160757 78644
rect 160875 78708 160941 78709
rect 160875 78644 160876 78708
rect 160940 78644 160941 78708
rect 160875 78643 160941 78644
rect 159294 52954 159914 78000
rect 160694 64565 160754 78643
rect 160691 64564 160757 64565
rect 160691 64500 160692 64564
rect 160756 64500 160757 64564
rect 160691 64499 160757 64500
rect 160878 54909 160938 78643
rect 160875 54908 160941 54909
rect 160875 54844 160876 54908
rect 160940 54844 160941 54908
rect 160875 54843 160941 54844
rect 161062 53685 161122 79867
rect 161243 79796 161309 79797
rect 161243 79732 161244 79796
rect 161308 79732 161309 79796
rect 161243 79731 161309 79732
rect 161059 53684 161125 53685
rect 161059 53620 161060 53684
rect 161124 53620 161125 53684
rect 161059 53619 161125 53620
rect 159294 52718 159326 52954
rect 159562 52718 159646 52954
rect 159882 52718 159914 52954
rect 159294 52634 159914 52718
rect 159294 52398 159326 52634
rect 159562 52398 159646 52634
rect 159882 52398 159914 52634
rect 159035 52324 159101 52325
rect 159035 52260 159036 52324
rect 159100 52260 159101 52324
rect 159035 52259 159101 52260
rect 158483 21996 158549 21997
rect 158483 21932 158484 21996
rect 158548 21932 158549 21996
rect 158483 21931 158549 21932
rect 158299 21860 158365 21861
rect 158299 21796 158300 21860
rect 158364 21796 158365 21860
rect 158299 21795 158365 21796
rect 155723 20636 155789 20637
rect 155723 20572 155724 20636
rect 155788 20572 155789 20636
rect 155723 20571 155789 20572
rect 154794 12218 154826 12454
rect 155062 12218 155146 12454
rect 155382 12218 155414 12454
rect 154794 12134 155414 12218
rect 154794 11898 154826 12134
rect 155062 11898 155146 12134
rect 155382 11898 155414 12134
rect 154794 -2266 155414 11898
rect 154794 -2502 154826 -2266
rect 155062 -2502 155146 -2266
rect 155382 -2502 155414 -2266
rect 154794 -2586 155414 -2502
rect 154794 -2822 154826 -2586
rect 155062 -2822 155146 -2586
rect 155382 -2822 155414 -2586
rect 154794 -7654 155414 -2822
rect 159294 16954 159914 52398
rect 161246 50421 161306 79731
rect 161982 77349 162042 79867
rect 162163 79660 162229 79661
rect 162163 79596 162164 79660
rect 162228 79596 162229 79660
rect 162163 79595 162229 79596
rect 161979 77348 162045 77349
rect 161979 77284 161980 77348
rect 162044 77284 162045 77348
rect 161979 77283 162045 77284
rect 162166 73813 162226 79595
rect 162350 78301 162410 79867
rect 162715 79796 162781 79797
rect 162715 79732 162716 79796
rect 162780 79732 162781 79796
rect 162715 79731 162781 79732
rect 162347 78300 162413 78301
rect 162347 78236 162348 78300
rect 162412 78236 162413 78300
rect 162347 78235 162413 78236
rect 162347 77348 162413 77349
rect 162347 77284 162348 77348
rect 162412 77284 162413 77348
rect 162347 77283 162413 77284
rect 162531 77348 162597 77349
rect 162531 77284 162532 77348
rect 162596 77284 162597 77348
rect 162531 77283 162597 77284
rect 162163 73812 162229 73813
rect 162163 73748 162164 73812
rect 162228 73748 162229 73812
rect 162163 73747 162229 73748
rect 162350 59125 162410 77283
rect 162347 59124 162413 59125
rect 162347 59060 162348 59124
rect 162412 59060 162413 59124
rect 162347 59059 162413 59060
rect 162534 56405 162594 77283
rect 162531 56404 162597 56405
rect 162531 56340 162532 56404
rect 162596 56340 162597 56404
rect 162531 56339 162597 56340
rect 161243 50420 161309 50421
rect 161243 50356 161244 50420
rect 161308 50356 161309 50420
rect 161243 50355 161309 50356
rect 162718 49469 162778 79731
rect 162902 77349 162962 79867
rect 163083 79796 163149 79797
rect 163083 79732 163084 79796
rect 163148 79732 163149 79796
rect 163083 79731 163149 79732
rect 163451 79796 163517 79797
rect 163451 79732 163452 79796
rect 163516 79732 163517 79796
rect 163451 79731 163517 79732
rect 165291 79796 165357 79797
rect 165291 79732 165292 79796
rect 165356 79732 165357 79796
rect 165291 79731 165357 79732
rect 165475 79796 165541 79797
rect 165475 79732 165476 79796
rect 165540 79732 165541 79796
rect 165475 79731 165541 79732
rect 163086 78029 163146 79731
rect 163267 79660 163333 79661
rect 163267 79596 163268 79660
rect 163332 79596 163333 79660
rect 163267 79595 163333 79596
rect 163083 78028 163149 78029
rect 163083 77964 163084 78028
rect 163148 77964 163149 78028
rect 163083 77963 163149 77964
rect 162899 77348 162965 77349
rect 162899 77284 162900 77348
rect 162964 77284 162965 77348
rect 162899 77283 162965 77284
rect 163270 52461 163330 79595
rect 163454 77893 163514 79731
rect 165107 79660 165173 79661
rect 165107 79596 165108 79660
rect 165172 79596 165173 79660
rect 165107 79595 165173 79596
rect 163451 77892 163517 77893
rect 163451 77828 163452 77892
rect 163516 77828 163517 77892
rect 163451 77827 163517 77828
rect 163635 77892 163701 77893
rect 163635 77828 163636 77892
rect 163700 77828 163701 77892
rect 163635 77827 163701 77828
rect 163451 77756 163517 77757
rect 163451 77692 163452 77756
rect 163516 77692 163517 77756
rect 163451 77691 163517 77692
rect 163267 52460 163333 52461
rect 163267 52396 163268 52460
rect 163332 52396 163333 52460
rect 163267 52395 163333 52396
rect 162715 49468 162781 49469
rect 162715 49404 162716 49468
rect 162780 49404 162781 49468
rect 162715 49403 162781 49404
rect 163454 48109 163514 77691
rect 163451 48108 163517 48109
rect 163451 48044 163452 48108
rect 163516 48044 163517 48108
rect 163451 48043 163517 48044
rect 163638 44165 163698 77827
rect 163794 57454 164414 78000
rect 164739 77348 164805 77349
rect 164739 77284 164740 77348
rect 164804 77284 164805 77348
rect 164739 77283 164805 77284
rect 164742 66061 164802 77283
rect 164739 66060 164805 66061
rect 164739 65996 164740 66060
rect 164804 65996 164805 66060
rect 164739 65995 164805 65996
rect 165110 57765 165170 79595
rect 165107 57764 165173 57765
rect 165107 57700 165108 57764
rect 165172 57700 165173 57764
rect 165107 57699 165173 57700
rect 163794 57218 163826 57454
rect 164062 57218 164146 57454
rect 164382 57218 164414 57454
rect 163794 57134 164414 57218
rect 163794 56898 163826 57134
rect 164062 56898 164146 57134
rect 164382 56898 164414 57134
rect 163635 44164 163701 44165
rect 163635 44100 163636 44164
rect 163700 44100 163701 44164
rect 163635 44099 163701 44100
rect 159294 16718 159326 16954
rect 159562 16718 159646 16954
rect 159882 16718 159914 16954
rect 159294 16634 159914 16718
rect 159294 16398 159326 16634
rect 159562 16398 159646 16634
rect 159882 16398 159914 16634
rect 159294 -3226 159914 16398
rect 159294 -3462 159326 -3226
rect 159562 -3462 159646 -3226
rect 159882 -3462 159914 -3226
rect 159294 -3546 159914 -3462
rect 159294 -3782 159326 -3546
rect 159562 -3782 159646 -3546
rect 159882 -3782 159914 -3546
rect 159294 -7654 159914 -3782
rect 163794 21454 164414 56898
rect 165294 46885 165354 79731
rect 165291 46884 165357 46885
rect 165291 46820 165292 46884
rect 165356 46820 165357 46884
rect 165291 46819 165357 46820
rect 165478 35869 165538 79731
rect 166214 70141 166274 79867
rect 166395 79660 166461 79661
rect 166395 79596 166396 79660
rect 166460 79596 166461 79660
rect 166395 79595 166461 79596
rect 166211 70140 166277 70141
rect 166211 70076 166212 70140
rect 166276 70076 166277 70140
rect 166211 70075 166277 70076
rect 166398 55045 166458 79595
rect 166395 55044 166461 55045
rect 166395 54980 166396 55044
rect 166460 54980 166461 55044
rect 166395 54979 166461 54980
rect 166582 53821 166642 79867
rect 167315 79796 167381 79797
rect 167315 79732 167316 79796
rect 167380 79732 167381 79796
rect 167315 79731 167381 79732
rect 167867 79796 167933 79797
rect 167867 79732 167868 79796
rect 167932 79794 167933 79796
rect 167932 79734 168114 79794
rect 167932 79732 167933 79734
rect 167867 79731 167933 79732
rect 166763 79660 166829 79661
rect 166763 79596 166764 79660
rect 166828 79596 166829 79660
rect 166763 79595 166829 79596
rect 166579 53820 166645 53821
rect 166579 53756 166580 53820
rect 166644 53756 166645 53820
rect 166579 53755 166645 53756
rect 166766 45389 166826 79595
rect 167318 78029 167378 79731
rect 167683 79660 167749 79661
rect 167683 79596 167684 79660
rect 167748 79596 167749 79660
rect 167683 79595 167749 79596
rect 167315 78028 167381 78029
rect 167315 77964 167316 78028
rect 167380 77964 167381 78028
rect 167315 77963 167381 77964
rect 167499 77348 167565 77349
rect 167499 77284 167500 77348
rect 167564 77284 167565 77348
rect 167499 77283 167565 77284
rect 167502 63341 167562 77283
rect 167499 63340 167565 63341
rect 167499 63276 167500 63340
rect 167564 63276 167565 63340
rect 167499 63275 167565 63276
rect 167686 62117 167746 79595
rect 167867 78028 167933 78029
rect 167867 77964 167868 78028
rect 167932 77964 167933 78028
rect 167867 77963 167933 77964
rect 167683 62116 167749 62117
rect 167683 62052 167684 62116
rect 167748 62052 167749 62116
rect 167683 62051 167749 62052
rect 167870 58989 167930 77963
rect 167867 58988 167933 58989
rect 167867 58924 167868 58988
rect 167932 58924 167933 58988
rect 167867 58923 167933 58924
rect 168054 55997 168114 79734
rect 168294 61954 168914 78000
rect 168294 61718 168326 61954
rect 168562 61718 168646 61954
rect 168882 61718 168914 61954
rect 168294 61634 168914 61718
rect 168294 61398 168326 61634
rect 168562 61398 168646 61634
rect 168882 61398 168914 61634
rect 168051 55996 168117 55997
rect 168051 55932 168052 55996
rect 168116 55932 168117 55996
rect 168051 55931 168117 55932
rect 166763 45388 166829 45389
rect 166763 45324 166764 45388
rect 166828 45324 166829 45388
rect 166763 45323 166829 45324
rect 165475 35868 165541 35869
rect 165475 35804 165476 35868
rect 165540 35804 165541 35868
rect 165475 35803 165541 35804
rect 163794 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 164414 21454
rect 163794 21134 164414 21218
rect 163794 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 164414 21134
rect 163794 -4186 164414 20898
rect 163794 -4422 163826 -4186
rect 164062 -4422 164146 -4186
rect 164382 -4422 164414 -4186
rect 163794 -4506 164414 -4422
rect 163794 -4742 163826 -4506
rect 164062 -4742 164146 -4506
rect 164382 -4742 164414 -4506
rect 163794 -7654 164414 -4742
rect 168294 25954 168914 61398
rect 169342 53549 169402 79867
rect 169339 53548 169405 53549
rect 169339 53484 169340 53548
rect 169404 53484 169405 53548
rect 169339 53483 169405 53484
rect 169526 47973 169586 80003
rect 170627 79932 170693 79933
rect 170627 79930 170628 79932
rect 170446 79870 170628 79930
rect 169523 47972 169589 47973
rect 169523 47908 169524 47972
rect 169588 47908 169589 47972
rect 169523 47907 169589 47908
rect 170446 47565 170506 79870
rect 170627 79868 170628 79870
rect 170692 79868 170693 79932
rect 170627 79867 170693 79868
rect 170627 79796 170693 79797
rect 170627 79732 170628 79796
rect 170692 79732 170693 79796
rect 170627 79731 170693 79732
rect 170630 79389 170690 79731
rect 170627 79388 170693 79389
rect 170627 79324 170628 79388
rect 170692 79324 170693 79388
rect 170627 79323 170693 79324
rect 170627 78572 170693 78573
rect 170627 78508 170628 78572
rect 170692 78508 170693 78572
rect 170627 78507 170693 78508
rect 170630 60621 170690 78507
rect 170627 60620 170693 60621
rect 170627 60556 170628 60620
rect 170692 60556 170693 60620
rect 170627 60555 170693 60556
rect 170814 56541 170874 80139
rect 173571 80068 173637 80069
rect 173571 80004 173572 80068
rect 173636 80004 173637 80068
rect 173571 80003 173637 80004
rect 172099 79932 172165 79933
rect 172099 79930 172100 79932
rect 171918 79870 172100 79930
rect 170995 79660 171061 79661
rect 170995 79596 170996 79660
rect 171060 79596 171061 79660
rect 170995 79595 171061 79596
rect 170998 75717 171058 79595
rect 171918 79389 171978 79870
rect 172099 79868 172100 79870
rect 172164 79868 172165 79932
rect 172099 79867 172165 79868
rect 173203 79932 173269 79933
rect 173203 79868 173204 79932
rect 173268 79868 173269 79932
rect 173203 79867 173269 79868
rect 172283 79796 172349 79797
rect 172283 79732 172284 79796
rect 172348 79732 172349 79796
rect 172283 79731 172349 79732
rect 172099 79660 172165 79661
rect 172099 79596 172100 79660
rect 172164 79596 172165 79660
rect 172099 79595 172165 79596
rect 171915 79388 171981 79389
rect 171915 79324 171916 79388
rect 171980 79324 171981 79388
rect 171915 79323 171981 79324
rect 171731 78708 171797 78709
rect 171731 78644 171732 78708
rect 171796 78644 171797 78708
rect 171731 78643 171797 78644
rect 171915 78708 171981 78709
rect 171915 78644 171916 78708
rect 171980 78644 171981 78708
rect 171915 78643 171981 78644
rect 170995 75716 171061 75717
rect 170995 75652 170996 75716
rect 171060 75652 171061 75716
rect 170995 75651 171061 75652
rect 170811 56540 170877 56541
rect 170811 56476 170812 56540
rect 170876 56476 170877 56540
rect 170811 56475 170877 56476
rect 171734 49333 171794 78643
rect 171918 64701 171978 78643
rect 171915 64700 171981 64701
rect 171915 64636 171916 64700
rect 171980 64636 171981 64700
rect 171915 64635 171981 64636
rect 172102 58853 172162 79595
rect 172099 58852 172165 58853
rect 172099 58788 172100 58852
rect 172164 58788 172165 58852
rect 172099 58787 172165 58788
rect 172286 55181 172346 79731
rect 173206 78165 173266 79867
rect 173203 78164 173269 78165
rect 173203 78100 173204 78164
rect 173268 78100 173269 78164
rect 173203 78099 173269 78100
rect 172794 66454 173414 78000
rect 172794 66218 172826 66454
rect 173062 66218 173146 66454
rect 173382 66218 173414 66454
rect 172794 66134 173414 66218
rect 172794 65898 172826 66134
rect 173062 65898 173146 66134
rect 173382 65898 173414 66134
rect 172283 55180 172349 55181
rect 172283 55116 172284 55180
rect 172348 55116 172349 55180
rect 172283 55115 172349 55116
rect 171731 49332 171797 49333
rect 171731 49268 171732 49332
rect 171796 49268 171797 49332
rect 171731 49267 171797 49268
rect 170443 47564 170509 47565
rect 170443 47500 170444 47564
rect 170508 47500 170509 47564
rect 170443 47499 170509 47500
rect 168294 25718 168326 25954
rect 168562 25718 168646 25954
rect 168882 25718 168914 25954
rect 168294 25634 168914 25718
rect 168294 25398 168326 25634
rect 168562 25398 168646 25634
rect 168882 25398 168914 25634
rect 168294 -5146 168914 25398
rect 168294 -5382 168326 -5146
rect 168562 -5382 168646 -5146
rect 168882 -5382 168914 -5146
rect 168294 -5466 168914 -5382
rect 168294 -5702 168326 -5466
rect 168562 -5702 168646 -5466
rect 168882 -5702 168914 -5466
rect 168294 -7654 168914 -5702
rect 172794 30454 173414 65898
rect 173574 45253 173634 80003
rect 173939 79932 174005 79933
rect 173939 79868 173940 79932
rect 174004 79868 174005 79932
rect 173939 79867 174005 79868
rect 173755 79796 173821 79797
rect 173755 79732 173756 79796
rect 173820 79732 173821 79796
rect 173755 79731 173821 79732
rect 173571 45252 173637 45253
rect 173571 45188 173572 45252
rect 173636 45188 173637 45252
rect 173571 45187 173637 45188
rect 173758 44981 173818 79731
rect 173942 76397 174002 79867
rect 174491 79796 174557 79797
rect 174491 79732 174492 79796
rect 174556 79732 174557 79796
rect 174859 79796 174925 79797
rect 174859 79794 174860 79796
rect 174491 79731 174557 79732
rect 174678 79734 174860 79794
rect 173939 76396 174005 76397
rect 173939 76332 173940 76396
rect 174004 76332 174005 76396
rect 173939 76331 174005 76332
rect 174494 51781 174554 79731
rect 174491 51780 174557 51781
rect 174491 51716 174492 51780
rect 174556 51716 174557 51780
rect 174491 51715 174557 51716
rect 174678 49605 174738 79734
rect 174859 79732 174860 79734
rect 174924 79732 174925 79796
rect 174859 79731 174925 79732
rect 174859 79660 174925 79661
rect 174859 79596 174860 79660
rect 174924 79596 174925 79660
rect 174859 79595 174925 79596
rect 174675 49604 174741 49605
rect 174675 49540 174676 49604
rect 174740 49540 174741 49604
rect 174675 49539 174741 49540
rect 173755 44980 173821 44981
rect 173755 44916 173756 44980
rect 173820 44916 173821 44980
rect 173755 44915 173821 44916
rect 174862 43485 174922 79595
rect 175046 79389 175106 81227
rect 175595 81156 175661 81157
rect 175595 81092 175596 81156
rect 175660 81092 175661 81156
rect 175595 81091 175661 81092
rect 175598 79661 175658 81091
rect 177251 81020 177317 81021
rect 177251 80956 177252 81020
rect 177316 80956 177317 81020
rect 177251 80955 177317 80956
rect 177254 80341 177314 80955
rect 177251 80340 177317 80341
rect 177251 80276 177252 80340
rect 177316 80276 177317 80340
rect 177251 80275 177317 80276
rect 175779 79932 175845 79933
rect 175779 79868 175780 79932
rect 175844 79868 175845 79932
rect 175779 79867 175845 79868
rect 176515 79932 176581 79933
rect 176515 79868 176516 79932
rect 176580 79868 176581 79932
rect 176515 79867 176581 79868
rect 175595 79660 175661 79661
rect 175595 79596 175596 79660
rect 175660 79596 175661 79660
rect 175595 79595 175661 79596
rect 175043 79388 175109 79389
rect 175043 79324 175044 79388
rect 175108 79324 175109 79388
rect 175043 79323 175109 79324
rect 175598 78437 175658 79595
rect 175595 78436 175661 78437
rect 175595 78372 175596 78436
rect 175660 78372 175661 78436
rect 175595 78371 175661 78372
rect 175043 78300 175109 78301
rect 175043 78236 175044 78300
rect 175108 78236 175109 78300
rect 175043 78235 175109 78236
rect 174859 43484 174925 43485
rect 174859 43420 174860 43484
rect 174924 43420 174925 43484
rect 174859 43419 174925 43420
rect 175046 37229 175106 78235
rect 175782 77485 175842 79867
rect 175963 79660 176029 79661
rect 175963 79596 175964 79660
rect 176028 79596 176029 79660
rect 175963 79595 176029 79596
rect 175966 77621 176026 79595
rect 176147 78300 176213 78301
rect 176147 78236 176148 78300
rect 176212 78236 176213 78300
rect 176147 78235 176213 78236
rect 175963 77620 176029 77621
rect 175963 77556 175964 77620
rect 176028 77556 176029 77620
rect 175963 77555 176029 77556
rect 175779 77484 175845 77485
rect 175779 77420 175780 77484
rect 175844 77420 175845 77484
rect 175779 77419 175845 77420
rect 175963 77348 176029 77349
rect 175963 77284 175964 77348
rect 176028 77284 176029 77348
rect 175963 77283 176029 77284
rect 175966 50693 176026 77283
rect 176150 61981 176210 78235
rect 176518 74550 176578 79867
rect 178910 78029 178970 81499
rect 178907 78028 178973 78029
rect 176334 74490 176578 74550
rect 176147 61980 176213 61981
rect 176147 61916 176148 61980
rect 176212 61916 176213 61980
rect 176147 61915 176213 61916
rect 176334 54637 176394 74490
rect 177294 70954 177914 78000
rect 178907 77964 178908 78028
rect 178972 77964 178973 78028
rect 178907 77963 178973 77964
rect 177294 70718 177326 70954
rect 177562 70718 177646 70954
rect 177882 70718 177914 70954
rect 177294 70634 177914 70718
rect 177294 70398 177326 70634
rect 177562 70398 177646 70634
rect 177882 70398 177914 70634
rect 176331 54636 176397 54637
rect 176331 54572 176332 54636
rect 176396 54572 176397 54636
rect 176331 54571 176397 54572
rect 175963 50692 176029 50693
rect 175963 50628 175964 50692
rect 176028 50628 176029 50692
rect 175963 50627 176029 50628
rect 175043 37228 175109 37229
rect 175043 37164 175044 37228
rect 175108 37164 175109 37228
rect 175043 37163 175109 37164
rect 172794 30218 172826 30454
rect 173062 30218 173146 30454
rect 173382 30218 173414 30454
rect 172794 30134 173414 30218
rect 172794 29898 172826 30134
rect 173062 29898 173146 30134
rect 173382 29898 173414 30134
rect 172794 -6106 173414 29898
rect 172794 -6342 172826 -6106
rect 173062 -6342 173146 -6106
rect 173382 -6342 173414 -6106
rect 172794 -6426 173414 -6342
rect 172794 -6662 172826 -6426
rect 173062 -6662 173146 -6426
rect 173382 -6662 173414 -6426
rect 172794 -7654 173414 -6662
rect 177294 34954 177914 70398
rect 177294 34718 177326 34954
rect 177562 34718 177646 34954
rect 177882 34718 177914 34954
rect 177294 34634 177914 34718
rect 177294 34398 177326 34634
rect 177562 34398 177646 34634
rect 177882 34398 177914 34634
rect 177294 -7066 177914 34398
rect 177294 -7302 177326 -7066
rect 177562 -7302 177646 -7066
rect 177882 -7302 177914 -7066
rect 177294 -7386 177914 -7302
rect 177294 -7622 177326 -7386
rect 177562 -7622 177646 -7386
rect 177882 -7622 177914 -7386
rect 177294 -7654 177914 -7622
rect 181794 75454 182414 78000
rect 181794 75218 181826 75454
rect 182062 75218 182146 75454
rect 182382 75218 182414 75454
rect 181794 75134 182414 75218
rect 181794 74898 181826 75134
rect 182062 74898 182146 75134
rect 182382 74898 182414 75134
rect 181794 39454 182414 74898
rect 184062 67149 184122 81771
rect 185347 81700 185413 81701
rect 185347 81636 185348 81700
rect 185412 81636 185413 81700
rect 185347 81635 185413 81636
rect 184243 80340 184309 80341
rect 184243 80276 184244 80340
rect 184308 80276 184309 80340
rect 184243 80275 184309 80276
rect 184246 67421 184306 80275
rect 185350 79933 185410 81635
rect 185902 80070 185962 81910
rect 186270 81290 186330 82043
rect 186086 81230 186330 81290
rect 186086 80202 186146 81230
rect 186454 80205 186514 138075
rect 186635 104956 186701 104957
rect 186635 104892 186636 104956
rect 186700 104892 186701 104956
rect 186635 104891 186701 104892
rect 186638 90405 186698 104891
rect 186635 90404 186701 90405
rect 186635 90340 186636 90404
rect 186700 90340 186701 90404
rect 186635 90339 186701 90340
rect 186635 86324 186701 86325
rect 186635 86260 186636 86324
rect 186700 86260 186701 86324
rect 186635 86259 186701 86260
rect 186638 81701 186698 86259
rect 186635 81700 186701 81701
rect 186635 81636 186636 81700
rect 186700 81636 186701 81700
rect 186635 81635 186701 81636
rect 186451 80204 186517 80205
rect 186086 80142 186330 80202
rect 185531 80068 185597 80069
rect 185531 80004 185532 80068
rect 185596 80004 185597 80068
rect 185902 80010 186146 80070
rect 186270 80069 186330 80142
rect 186451 80140 186452 80204
rect 186516 80140 186517 80204
rect 186451 80139 186517 80140
rect 185531 80003 185597 80004
rect 185347 79932 185413 79933
rect 185347 79868 185348 79932
rect 185412 79868 185413 79932
rect 185347 79867 185413 79868
rect 185347 79660 185413 79661
rect 185347 79596 185348 79660
rect 185412 79596 185413 79660
rect 185347 79595 185413 79596
rect 185350 68645 185410 79595
rect 185534 70413 185594 80003
rect 185531 70412 185597 70413
rect 185531 70348 185532 70412
rect 185596 70348 185597 70412
rect 185531 70347 185597 70348
rect 185347 68644 185413 68645
rect 185347 68580 185348 68644
rect 185412 68580 185413 68644
rect 185347 68579 185413 68580
rect 184243 67420 184309 67421
rect 184243 67356 184244 67420
rect 184308 67356 184309 67420
rect 184243 67355 184309 67356
rect 186086 67285 186146 80010
rect 186267 80068 186333 80069
rect 186267 80004 186268 80068
rect 186332 80004 186333 80068
rect 186267 80003 186333 80004
rect 187006 79253 187066 193155
rect 187371 145892 187437 145893
rect 187371 145828 187372 145892
rect 187436 145828 187437 145892
rect 187371 145827 187437 145828
rect 187187 139908 187253 139909
rect 187187 139844 187188 139908
rect 187252 139844 187253 139908
rect 187187 139843 187253 139844
rect 187003 79252 187069 79253
rect 187003 79188 187004 79252
rect 187068 79188 187069 79252
rect 187003 79187 187069 79188
rect 186083 67284 186149 67285
rect 186083 67220 186084 67284
rect 186148 67220 186149 67284
rect 186083 67219 186149 67220
rect 184059 67148 184125 67149
rect 184059 67084 184060 67148
rect 184124 67084 184125 67148
rect 184059 67083 184125 67084
rect 181794 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 182414 39454
rect 181794 39134 182414 39218
rect 181794 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 182414 39134
rect 181794 3454 182414 38898
rect 181794 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 182414 3454
rect 181794 3134 182414 3218
rect 181794 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 182414 3134
rect 181794 -346 182414 2898
rect 181794 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 182414 -346
rect 181794 -666 182414 -582
rect 181794 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 182414 -666
rect 181794 -7654 182414 -902
rect 186294 43954 186914 78000
rect 187190 63477 187250 139843
rect 187374 78709 187434 145827
rect 187742 142901 187802 277475
rect 190794 264454 191414 299898
rect 195294 707718 195914 711590
rect 195294 707482 195326 707718
rect 195562 707482 195646 707718
rect 195882 707482 195914 707718
rect 195294 707398 195914 707482
rect 195294 707162 195326 707398
rect 195562 707162 195646 707398
rect 195882 707162 195914 707398
rect 195294 700954 195914 707162
rect 195294 700718 195326 700954
rect 195562 700718 195646 700954
rect 195882 700718 195914 700954
rect 195294 700634 195914 700718
rect 195294 700398 195326 700634
rect 195562 700398 195646 700634
rect 195882 700398 195914 700634
rect 195294 664954 195914 700398
rect 195294 664718 195326 664954
rect 195562 664718 195646 664954
rect 195882 664718 195914 664954
rect 195294 664634 195914 664718
rect 195294 664398 195326 664634
rect 195562 664398 195646 664634
rect 195882 664398 195914 664634
rect 195294 628954 195914 664398
rect 195294 628718 195326 628954
rect 195562 628718 195646 628954
rect 195882 628718 195914 628954
rect 195294 628634 195914 628718
rect 195294 628398 195326 628634
rect 195562 628398 195646 628634
rect 195882 628398 195914 628634
rect 195294 592954 195914 628398
rect 195294 592718 195326 592954
rect 195562 592718 195646 592954
rect 195882 592718 195914 592954
rect 195294 592634 195914 592718
rect 195294 592398 195326 592634
rect 195562 592398 195646 592634
rect 195882 592398 195914 592634
rect 195294 556954 195914 592398
rect 195294 556718 195326 556954
rect 195562 556718 195646 556954
rect 195882 556718 195914 556954
rect 195294 556634 195914 556718
rect 195294 556398 195326 556634
rect 195562 556398 195646 556634
rect 195882 556398 195914 556634
rect 195294 520954 195914 556398
rect 195294 520718 195326 520954
rect 195562 520718 195646 520954
rect 195882 520718 195914 520954
rect 195294 520634 195914 520718
rect 195294 520398 195326 520634
rect 195562 520398 195646 520634
rect 195882 520398 195914 520634
rect 195294 484954 195914 520398
rect 195294 484718 195326 484954
rect 195562 484718 195646 484954
rect 195882 484718 195914 484954
rect 195294 484634 195914 484718
rect 195294 484398 195326 484634
rect 195562 484398 195646 484634
rect 195882 484398 195914 484634
rect 195294 448954 195914 484398
rect 195294 448718 195326 448954
rect 195562 448718 195646 448954
rect 195882 448718 195914 448954
rect 195294 448634 195914 448718
rect 195294 448398 195326 448634
rect 195562 448398 195646 448634
rect 195882 448398 195914 448634
rect 195294 412954 195914 448398
rect 195294 412718 195326 412954
rect 195562 412718 195646 412954
rect 195882 412718 195914 412954
rect 195294 412634 195914 412718
rect 195294 412398 195326 412634
rect 195562 412398 195646 412634
rect 195882 412398 195914 412634
rect 195294 376954 195914 412398
rect 195294 376718 195326 376954
rect 195562 376718 195646 376954
rect 195882 376718 195914 376954
rect 195294 376634 195914 376718
rect 195294 376398 195326 376634
rect 195562 376398 195646 376634
rect 195882 376398 195914 376634
rect 195294 340954 195914 376398
rect 195294 340718 195326 340954
rect 195562 340718 195646 340954
rect 195882 340718 195914 340954
rect 195294 340634 195914 340718
rect 195294 340398 195326 340634
rect 195562 340398 195646 340634
rect 195882 340398 195914 340634
rect 195294 304954 195914 340398
rect 195294 304718 195326 304954
rect 195562 304718 195646 304954
rect 195882 304718 195914 304954
rect 195294 304634 195914 304718
rect 195294 304398 195326 304634
rect 195562 304398 195646 304634
rect 195882 304398 195914 304634
rect 195294 268954 195914 304398
rect 195294 268718 195326 268954
rect 195562 268718 195646 268954
rect 195882 268718 195914 268954
rect 195294 268634 195914 268718
rect 195294 268398 195326 268634
rect 195562 268398 195646 268634
rect 195882 268398 195914 268634
rect 192155 265164 192221 265165
rect 192155 265100 192156 265164
rect 192220 265100 192221 265164
rect 192155 265099 192221 265100
rect 190794 264218 190826 264454
rect 191062 264218 191146 264454
rect 191382 264218 191414 264454
rect 190794 264134 191414 264218
rect 190794 263898 190826 264134
rect 191062 263898 191146 264134
rect 191382 263898 191414 264134
rect 190499 262444 190565 262445
rect 190499 262380 190500 262444
rect 190564 262380 190565 262444
rect 190499 262379 190565 262380
rect 189027 259860 189093 259861
rect 189027 259796 189028 259860
rect 189092 259796 189093 259860
rect 189027 259795 189093 259796
rect 187923 192404 187989 192405
rect 187923 192340 187924 192404
rect 187988 192340 187989 192404
rect 187923 192339 187989 192340
rect 187739 142900 187805 142901
rect 187739 142836 187740 142900
rect 187804 142836 187805 142900
rect 187739 142835 187805 142836
rect 187739 139636 187805 139637
rect 187739 139572 187740 139636
rect 187804 139572 187805 139636
rect 187739 139571 187805 139572
rect 187742 138141 187802 139571
rect 187739 138140 187805 138141
rect 187739 138076 187740 138140
rect 187804 138076 187805 138140
rect 187739 138075 187805 138076
rect 187926 78981 187986 192339
rect 188291 149972 188357 149973
rect 188291 149908 188292 149972
rect 188356 149908 188357 149972
rect 188291 149907 188357 149908
rect 188107 139772 188173 139773
rect 188107 139708 188108 139772
rect 188172 139708 188173 139772
rect 188107 139707 188173 139708
rect 187923 78980 187989 78981
rect 187923 78916 187924 78980
rect 187988 78916 187989 78980
rect 187923 78915 187989 78916
rect 187371 78708 187437 78709
rect 187371 78644 187372 78708
rect 187436 78644 187437 78708
rect 187371 78643 187437 78644
rect 188110 72317 188170 139707
rect 188294 75309 188354 149907
rect 189030 141677 189090 259795
rect 189211 259724 189277 259725
rect 189211 259660 189212 259724
rect 189276 259660 189277 259724
rect 189211 259659 189277 259660
rect 189214 142085 189274 259659
rect 189395 149836 189461 149837
rect 189395 149772 189396 149836
rect 189460 149772 189461 149836
rect 189395 149771 189461 149772
rect 189211 142084 189277 142085
rect 189211 142020 189212 142084
rect 189276 142020 189277 142084
rect 189211 142019 189277 142020
rect 189027 141676 189093 141677
rect 189027 141612 189028 141676
rect 189092 141612 189093 141676
rect 189027 141611 189093 141612
rect 189027 90404 189093 90405
rect 189027 90340 189028 90404
rect 189092 90340 189093 90404
rect 189027 90339 189093 90340
rect 188291 75308 188357 75309
rect 188291 75244 188292 75308
rect 188356 75244 188357 75308
rect 188291 75243 188357 75244
rect 188107 72316 188173 72317
rect 188107 72252 188108 72316
rect 188172 72252 188173 72316
rect 188107 72251 188173 72252
rect 189030 68781 189090 90339
rect 189398 75173 189458 149771
rect 189763 146164 189829 146165
rect 189763 146100 189764 146164
rect 189828 146100 189829 146164
rect 189763 146099 189829 146100
rect 189579 140588 189645 140589
rect 189579 140524 189580 140588
rect 189644 140524 189645 140588
rect 189579 140523 189645 140524
rect 189582 81565 189642 140523
rect 189579 81564 189645 81565
rect 189579 81500 189580 81564
rect 189644 81500 189645 81564
rect 189579 81499 189645 81500
rect 189766 75445 189826 146099
rect 190502 144533 190562 262379
rect 190794 262000 191414 263898
rect 191787 263124 191853 263125
rect 191787 263060 191788 263124
rect 191852 263060 191853 263124
rect 191787 263059 191853 263060
rect 191790 262445 191850 263059
rect 191787 262444 191853 262445
rect 191787 262380 191788 262444
rect 191852 262380 191853 262444
rect 191787 262379 191853 262380
rect 190794 192454 191414 198000
rect 191971 197844 192037 197845
rect 191971 197780 191972 197844
rect 192036 197780 192037 197844
rect 191971 197779 192037 197780
rect 191787 195260 191853 195261
rect 191787 195196 191788 195260
rect 191852 195196 191853 195260
rect 191787 195195 191853 195196
rect 190794 192218 190826 192454
rect 191062 192218 191146 192454
rect 191382 192218 191414 192454
rect 190794 192134 191414 192218
rect 190794 191898 190826 192134
rect 191062 191898 191146 192134
rect 191382 191898 191414 192134
rect 190794 156454 191414 191898
rect 190794 156218 190826 156454
rect 191062 156218 191146 156454
rect 191382 156218 191414 156454
rect 190794 156134 191414 156218
rect 190794 155898 190826 156134
rect 191062 155898 191146 156134
rect 191382 155898 191414 156134
rect 190499 144532 190565 144533
rect 190499 144468 190500 144532
rect 190564 144468 190565 144532
rect 190499 144467 190565 144468
rect 190794 142000 191414 155898
rect 191603 146028 191669 146029
rect 191603 145964 191604 146028
rect 191668 145964 191669 146028
rect 191603 145963 191669 145964
rect 190499 141404 190565 141405
rect 190499 141340 190500 141404
rect 190564 141340 190565 141404
rect 190499 141339 190565 141340
rect 189763 75444 189829 75445
rect 189763 75380 189764 75444
rect 189828 75380 189829 75444
rect 189763 75379 189829 75380
rect 189395 75172 189461 75173
rect 189395 75108 189396 75172
rect 189460 75108 189461 75172
rect 189395 75107 189461 75108
rect 190502 70005 190562 141339
rect 191051 140724 191117 140725
rect 191051 140660 191052 140724
rect 191116 140660 191117 140724
rect 191051 140659 191117 140660
rect 190683 140044 190749 140045
rect 190683 139980 190684 140044
rect 190748 139980 190749 140044
rect 190683 139979 190749 139980
rect 190686 78301 190746 139979
rect 191054 79117 191114 140659
rect 191051 79116 191117 79117
rect 191051 79052 191052 79116
rect 191116 79052 191117 79116
rect 191051 79051 191117 79052
rect 190683 78300 190749 78301
rect 190683 78236 190684 78300
rect 190748 78236 190749 78300
rect 190683 78235 190749 78236
rect 190499 70004 190565 70005
rect 190499 69940 190500 70004
rect 190564 69940 190565 70004
rect 190499 69939 190565 69940
rect 189027 68780 189093 68781
rect 189027 68716 189028 68780
rect 189092 68716 189093 68780
rect 189027 68715 189093 68716
rect 187187 63476 187253 63477
rect 187187 63412 187188 63476
rect 187252 63412 187253 63476
rect 187187 63411 187253 63412
rect 186294 43718 186326 43954
rect 186562 43718 186646 43954
rect 186882 43718 186914 43954
rect 186294 43634 186914 43718
rect 186294 43398 186326 43634
rect 186562 43398 186646 43634
rect 186882 43398 186914 43634
rect 186294 7954 186914 43398
rect 186294 7718 186326 7954
rect 186562 7718 186646 7954
rect 186882 7718 186914 7954
rect 186294 7634 186914 7718
rect 186294 7398 186326 7634
rect 186562 7398 186646 7634
rect 186882 7398 186914 7634
rect 186294 -1306 186914 7398
rect 186294 -1542 186326 -1306
rect 186562 -1542 186646 -1306
rect 186882 -1542 186914 -1306
rect 186294 -1626 186914 -1542
rect 186294 -1862 186326 -1626
rect 186562 -1862 186646 -1626
rect 186882 -1862 186914 -1626
rect 186294 -7654 186914 -1862
rect 190794 48454 191414 78000
rect 191606 75581 191666 145963
rect 191603 75580 191669 75581
rect 191603 75516 191604 75580
rect 191668 75516 191669 75580
rect 191603 75515 191669 75516
rect 191790 50829 191850 195195
rect 191974 58581 192034 197779
rect 192158 141813 192218 265099
rect 193627 262716 193693 262717
rect 193627 262652 193628 262716
rect 193692 262652 193693 262716
rect 193627 262651 193693 262652
rect 192339 262308 192405 262309
rect 192339 262244 192340 262308
rect 192404 262244 192405 262308
rect 192339 262243 192405 262244
rect 192342 145621 192402 262243
rect 193443 260948 193509 260949
rect 193443 260884 193444 260948
rect 193508 260884 193509 260948
rect 193443 260883 193509 260884
rect 193259 198524 193325 198525
rect 193259 198460 193260 198524
rect 193324 198460 193325 198524
rect 193259 198459 193325 198460
rect 192339 145620 192405 145621
rect 192339 145556 192340 145620
rect 192404 145556 192405 145620
rect 192339 145555 192405 145556
rect 192339 143444 192405 143445
rect 192339 143380 192340 143444
rect 192404 143380 192405 143444
rect 192339 143379 192405 143380
rect 192155 141812 192221 141813
rect 192155 141748 192156 141812
rect 192220 141748 192221 141812
rect 192155 141747 192221 141748
rect 192155 140180 192221 140181
rect 192155 140116 192156 140180
rect 192220 140116 192221 140180
rect 192155 140115 192221 140116
rect 192158 72453 192218 140115
rect 192342 80477 192402 143379
rect 192339 80476 192405 80477
rect 192339 80412 192340 80476
rect 192404 80412 192405 80476
rect 192339 80411 192405 80412
rect 192155 72452 192221 72453
rect 192155 72388 192156 72452
rect 192220 72388 192221 72452
rect 192155 72387 192221 72388
rect 193262 67557 193322 198459
rect 193446 140725 193506 260883
rect 193630 144805 193690 262651
rect 195294 232954 195914 268398
rect 199794 708678 200414 711590
rect 199794 708442 199826 708678
rect 200062 708442 200146 708678
rect 200382 708442 200414 708678
rect 199794 708358 200414 708442
rect 199794 708122 199826 708358
rect 200062 708122 200146 708358
rect 200382 708122 200414 708358
rect 199794 669454 200414 708122
rect 199794 669218 199826 669454
rect 200062 669218 200146 669454
rect 200382 669218 200414 669454
rect 199794 669134 200414 669218
rect 199794 668898 199826 669134
rect 200062 668898 200146 669134
rect 200382 668898 200414 669134
rect 199794 633454 200414 668898
rect 199794 633218 199826 633454
rect 200062 633218 200146 633454
rect 200382 633218 200414 633454
rect 199794 633134 200414 633218
rect 199794 632898 199826 633134
rect 200062 632898 200146 633134
rect 200382 632898 200414 633134
rect 199794 597454 200414 632898
rect 199794 597218 199826 597454
rect 200062 597218 200146 597454
rect 200382 597218 200414 597454
rect 199794 597134 200414 597218
rect 199794 596898 199826 597134
rect 200062 596898 200146 597134
rect 200382 596898 200414 597134
rect 199794 561454 200414 596898
rect 199794 561218 199826 561454
rect 200062 561218 200146 561454
rect 200382 561218 200414 561454
rect 199794 561134 200414 561218
rect 199794 560898 199826 561134
rect 200062 560898 200146 561134
rect 200382 560898 200414 561134
rect 199794 525454 200414 560898
rect 199794 525218 199826 525454
rect 200062 525218 200146 525454
rect 200382 525218 200414 525454
rect 199794 525134 200414 525218
rect 199794 524898 199826 525134
rect 200062 524898 200146 525134
rect 200382 524898 200414 525134
rect 199794 489454 200414 524898
rect 199794 489218 199826 489454
rect 200062 489218 200146 489454
rect 200382 489218 200414 489454
rect 199794 489134 200414 489218
rect 199794 488898 199826 489134
rect 200062 488898 200146 489134
rect 200382 488898 200414 489134
rect 199794 453454 200414 488898
rect 199794 453218 199826 453454
rect 200062 453218 200146 453454
rect 200382 453218 200414 453454
rect 199794 453134 200414 453218
rect 199794 452898 199826 453134
rect 200062 452898 200146 453134
rect 200382 452898 200414 453134
rect 199794 417454 200414 452898
rect 199794 417218 199826 417454
rect 200062 417218 200146 417454
rect 200382 417218 200414 417454
rect 199794 417134 200414 417218
rect 199794 416898 199826 417134
rect 200062 416898 200146 417134
rect 200382 416898 200414 417134
rect 199794 381454 200414 416898
rect 199794 381218 199826 381454
rect 200062 381218 200146 381454
rect 200382 381218 200414 381454
rect 199794 381134 200414 381218
rect 199794 380898 199826 381134
rect 200062 380898 200146 381134
rect 200382 380898 200414 381134
rect 199794 345454 200414 380898
rect 199794 345218 199826 345454
rect 200062 345218 200146 345454
rect 200382 345218 200414 345454
rect 199794 345134 200414 345218
rect 199794 344898 199826 345134
rect 200062 344898 200146 345134
rect 200382 344898 200414 345134
rect 199794 309454 200414 344898
rect 199794 309218 199826 309454
rect 200062 309218 200146 309454
rect 200382 309218 200414 309454
rect 199794 309134 200414 309218
rect 199794 308898 199826 309134
rect 200062 308898 200146 309134
rect 200382 308898 200414 309134
rect 199794 273454 200414 308898
rect 199794 273218 199826 273454
rect 200062 273218 200146 273454
rect 200382 273218 200414 273454
rect 199794 273134 200414 273218
rect 199794 272898 199826 273134
rect 200062 272898 200146 273134
rect 200382 272898 200414 273134
rect 196387 265028 196453 265029
rect 196387 264964 196388 265028
rect 196452 264964 196453 265028
rect 196387 264963 196453 264964
rect 195294 232718 195326 232954
rect 195562 232718 195646 232954
rect 195882 232718 195914 232954
rect 195294 232634 195914 232718
rect 195294 232398 195326 232634
rect 195562 232398 195646 232634
rect 195882 232398 195914 232634
rect 195294 196954 195914 232398
rect 196019 198660 196085 198661
rect 196019 198596 196020 198660
rect 196084 198596 196085 198660
rect 196019 198595 196085 198596
rect 195294 196718 195326 196954
rect 195562 196718 195646 196954
rect 195882 196718 195914 196954
rect 195294 196634 195914 196718
rect 195294 196398 195326 196634
rect 195562 196398 195646 196634
rect 195882 196398 195914 196634
rect 193811 195940 193877 195941
rect 193811 195876 193812 195940
rect 193876 195876 193877 195940
rect 193811 195875 193877 195876
rect 193627 144804 193693 144805
rect 193627 144740 193628 144804
rect 193692 144740 193693 144804
rect 193627 144739 193693 144740
rect 193443 140724 193509 140725
rect 193443 140660 193444 140724
rect 193508 140660 193509 140724
rect 193443 140659 193509 140660
rect 193443 140452 193509 140453
rect 193443 140388 193444 140452
rect 193508 140388 193509 140452
rect 193443 140387 193509 140388
rect 193446 73677 193506 140387
rect 193627 140316 193693 140317
rect 193627 140252 193628 140316
rect 193692 140252 193693 140316
rect 193627 140251 193693 140252
rect 193630 76805 193690 140251
rect 193814 79389 193874 195875
rect 194547 195124 194613 195125
rect 194547 195060 194548 195124
rect 194612 195060 194613 195124
rect 194547 195059 194613 195060
rect 193811 79388 193877 79389
rect 193811 79324 193812 79388
rect 193876 79324 193877 79388
rect 193811 79323 193877 79324
rect 193627 76804 193693 76805
rect 193627 76740 193628 76804
rect 193692 76740 193693 76804
rect 193627 76739 193693 76740
rect 193443 73676 193509 73677
rect 193443 73612 193444 73676
rect 193508 73612 193509 73676
rect 193443 73611 193509 73612
rect 194550 68237 194610 195059
rect 195294 160954 195914 196398
rect 195294 160718 195326 160954
rect 195562 160718 195646 160954
rect 195882 160718 195914 160954
rect 195294 160634 195914 160718
rect 195294 160398 195326 160634
rect 195562 160398 195646 160634
rect 195882 160398 195914 160634
rect 194731 148204 194797 148205
rect 194731 148140 194732 148204
rect 194796 148140 194797 148204
rect 194731 148139 194797 148140
rect 194734 76669 194794 148139
rect 195294 124954 195914 160398
rect 195294 124718 195326 124954
rect 195562 124718 195646 124954
rect 195882 124718 195914 124954
rect 195294 124634 195914 124718
rect 195294 124398 195326 124634
rect 195562 124398 195646 124634
rect 195882 124398 195914 124634
rect 195294 88954 195914 124398
rect 195294 88718 195326 88954
rect 195562 88718 195646 88954
rect 195882 88718 195914 88954
rect 195294 88634 195914 88718
rect 195294 88398 195326 88634
rect 195562 88398 195646 88634
rect 195882 88398 195914 88634
rect 194731 76668 194797 76669
rect 194731 76604 194732 76668
rect 194796 76604 194797 76668
rect 194731 76603 194797 76604
rect 194547 68236 194613 68237
rect 194547 68172 194548 68236
rect 194612 68172 194613 68236
rect 194547 68171 194613 68172
rect 193259 67556 193325 67557
rect 193259 67492 193260 67556
rect 193324 67492 193325 67556
rect 193259 67491 193325 67492
rect 191971 58580 192037 58581
rect 191971 58516 191972 58580
rect 192036 58516 192037 58580
rect 191971 58515 192037 58516
rect 195294 52954 195914 88398
rect 196022 66197 196082 198595
rect 196203 198116 196269 198117
rect 196203 198052 196204 198116
rect 196268 198052 196269 198116
rect 196203 198051 196269 198052
rect 196206 71365 196266 198051
rect 196390 145757 196450 264963
rect 199794 237454 200414 272898
rect 199794 237218 199826 237454
rect 200062 237218 200146 237454
rect 200382 237218 200414 237454
rect 199794 237134 200414 237218
rect 199794 236898 199826 237134
rect 200062 236898 200146 237134
rect 200382 236898 200414 237134
rect 199794 201454 200414 236898
rect 199794 201218 199826 201454
rect 200062 201218 200146 201454
rect 200382 201218 200414 201454
rect 199794 201134 200414 201218
rect 199794 200898 199826 201134
rect 200062 200898 200146 201134
rect 200382 200898 200414 201134
rect 198963 199204 199029 199205
rect 198963 199140 198964 199204
rect 199028 199140 199029 199204
rect 198963 199139 199029 199140
rect 197307 198388 197373 198389
rect 197307 198324 197308 198388
rect 197372 198324 197373 198388
rect 197307 198323 197373 198324
rect 196571 147524 196637 147525
rect 196571 147460 196572 147524
rect 196636 147460 196637 147524
rect 196571 147459 196637 147460
rect 196387 145756 196453 145757
rect 196387 145692 196388 145756
rect 196452 145692 196453 145756
rect 196387 145691 196453 145692
rect 196574 81565 196634 147459
rect 196571 81564 196637 81565
rect 196571 81500 196572 81564
rect 196636 81500 196637 81564
rect 196571 81499 196637 81500
rect 197310 80749 197370 198323
rect 198779 197300 198845 197301
rect 198779 197236 198780 197300
rect 198844 197236 198845 197300
rect 198779 197235 198845 197236
rect 197859 149156 197925 149157
rect 197859 149092 197860 149156
rect 197924 149092 197925 149156
rect 197859 149091 197925 149092
rect 197491 149020 197557 149021
rect 197491 148956 197492 149020
rect 197556 148956 197557 149020
rect 197491 148955 197557 148956
rect 197494 81293 197554 148955
rect 197491 81292 197557 81293
rect 197491 81228 197492 81292
rect 197556 81228 197557 81292
rect 197491 81227 197557 81228
rect 197307 80748 197373 80749
rect 197307 80684 197308 80748
rect 197372 80684 197373 80748
rect 197307 80683 197373 80684
rect 196203 71364 196269 71365
rect 196203 71300 196204 71364
rect 196268 71300 196269 71364
rect 196203 71299 196269 71300
rect 196019 66196 196085 66197
rect 196019 66132 196020 66196
rect 196084 66132 196085 66196
rect 196019 66131 196085 66132
rect 197862 57629 197922 149091
rect 197859 57628 197925 57629
rect 197859 57564 197860 57628
rect 197924 57564 197925 57628
rect 197859 57563 197925 57564
rect 195294 52718 195326 52954
rect 195562 52718 195646 52954
rect 195882 52718 195914 52954
rect 195294 52634 195914 52718
rect 195294 52398 195326 52634
rect 195562 52398 195646 52634
rect 195882 52398 195914 52634
rect 191787 50828 191853 50829
rect 191787 50764 191788 50828
rect 191852 50764 191853 50828
rect 191787 50763 191853 50764
rect 193075 50828 193141 50829
rect 193075 50764 193076 50828
rect 193140 50764 193141 50828
rect 193075 50763 193141 50764
rect 193078 50557 193138 50763
rect 193075 50556 193141 50557
rect 193075 50492 193076 50556
rect 193140 50492 193141 50556
rect 193075 50491 193141 50492
rect 190794 48218 190826 48454
rect 191062 48218 191146 48454
rect 191382 48218 191414 48454
rect 190794 48134 191414 48218
rect 190794 47898 190826 48134
rect 191062 47898 191146 48134
rect 191382 47898 191414 48134
rect 190794 12454 191414 47898
rect 190794 12218 190826 12454
rect 191062 12218 191146 12454
rect 191382 12218 191414 12454
rect 190794 12134 191414 12218
rect 190794 11898 190826 12134
rect 191062 11898 191146 12134
rect 191382 11898 191414 12134
rect 190794 -2266 191414 11898
rect 190794 -2502 190826 -2266
rect 191062 -2502 191146 -2266
rect 191382 -2502 191414 -2266
rect 190794 -2586 191414 -2502
rect 190794 -2822 190826 -2586
rect 191062 -2822 191146 -2586
rect 191382 -2822 191414 -2586
rect 190794 -7654 191414 -2822
rect 195294 16954 195914 52398
rect 198782 46885 198842 197235
rect 198966 64837 199026 199139
rect 199147 198252 199213 198253
rect 199147 198188 199148 198252
rect 199212 198188 199213 198252
rect 199147 198187 199213 198188
rect 199150 66469 199210 198187
rect 199794 165454 200414 200898
rect 204294 709638 204914 711590
rect 204294 709402 204326 709638
rect 204562 709402 204646 709638
rect 204882 709402 204914 709638
rect 204294 709318 204914 709402
rect 204294 709082 204326 709318
rect 204562 709082 204646 709318
rect 204882 709082 204914 709318
rect 204294 673954 204914 709082
rect 204294 673718 204326 673954
rect 204562 673718 204646 673954
rect 204882 673718 204914 673954
rect 204294 673634 204914 673718
rect 204294 673398 204326 673634
rect 204562 673398 204646 673634
rect 204882 673398 204914 673634
rect 204294 637954 204914 673398
rect 204294 637718 204326 637954
rect 204562 637718 204646 637954
rect 204882 637718 204914 637954
rect 204294 637634 204914 637718
rect 204294 637398 204326 637634
rect 204562 637398 204646 637634
rect 204882 637398 204914 637634
rect 204294 601954 204914 637398
rect 204294 601718 204326 601954
rect 204562 601718 204646 601954
rect 204882 601718 204914 601954
rect 204294 601634 204914 601718
rect 204294 601398 204326 601634
rect 204562 601398 204646 601634
rect 204882 601398 204914 601634
rect 204294 565954 204914 601398
rect 204294 565718 204326 565954
rect 204562 565718 204646 565954
rect 204882 565718 204914 565954
rect 204294 565634 204914 565718
rect 204294 565398 204326 565634
rect 204562 565398 204646 565634
rect 204882 565398 204914 565634
rect 204294 529954 204914 565398
rect 204294 529718 204326 529954
rect 204562 529718 204646 529954
rect 204882 529718 204914 529954
rect 204294 529634 204914 529718
rect 204294 529398 204326 529634
rect 204562 529398 204646 529634
rect 204882 529398 204914 529634
rect 204294 493954 204914 529398
rect 204294 493718 204326 493954
rect 204562 493718 204646 493954
rect 204882 493718 204914 493954
rect 204294 493634 204914 493718
rect 204294 493398 204326 493634
rect 204562 493398 204646 493634
rect 204882 493398 204914 493634
rect 204294 457954 204914 493398
rect 204294 457718 204326 457954
rect 204562 457718 204646 457954
rect 204882 457718 204914 457954
rect 204294 457634 204914 457718
rect 204294 457398 204326 457634
rect 204562 457398 204646 457634
rect 204882 457398 204914 457634
rect 204294 421954 204914 457398
rect 204294 421718 204326 421954
rect 204562 421718 204646 421954
rect 204882 421718 204914 421954
rect 204294 421634 204914 421718
rect 204294 421398 204326 421634
rect 204562 421398 204646 421634
rect 204882 421398 204914 421634
rect 204294 385954 204914 421398
rect 204294 385718 204326 385954
rect 204562 385718 204646 385954
rect 204882 385718 204914 385954
rect 204294 385634 204914 385718
rect 204294 385398 204326 385634
rect 204562 385398 204646 385634
rect 204882 385398 204914 385634
rect 204294 349954 204914 385398
rect 204294 349718 204326 349954
rect 204562 349718 204646 349954
rect 204882 349718 204914 349954
rect 204294 349634 204914 349718
rect 204294 349398 204326 349634
rect 204562 349398 204646 349634
rect 204882 349398 204914 349634
rect 204294 313954 204914 349398
rect 204294 313718 204326 313954
rect 204562 313718 204646 313954
rect 204882 313718 204914 313954
rect 204294 313634 204914 313718
rect 204294 313398 204326 313634
rect 204562 313398 204646 313634
rect 204882 313398 204914 313634
rect 204294 277954 204914 313398
rect 204294 277718 204326 277954
rect 204562 277718 204646 277954
rect 204882 277718 204914 277954
rect 204294 277634 204914 277718
rect 204294 277398 204326 277634
rect 204562 277398 204646 277634
rect 204882 277398 204914 277634
rect 204294 241954 204914 277398
rect 204294 241718 204326 241954
rect 204562 241718 204646 241954
rect 204882 241718 204914 241954
rect 204294 241634 204914 241718
rect 204294 241398 204326 241634
rect 204562 241398 204646 241634
rect 204882 241398 204914 241634
rect 204294 205954 204914 241398
rect 204294 205718 204326 205954
rect 204562 205718 204646 205954
rect 204882 205718 204914 205954
rect 204294 205634 204914 205718
rect 204294 205398 204326 205634
rect 204562 205398 204646 205634
rect 204882 205398 204914 205634
rect 200803 199340 200869 199341
rect 200803 199276 200804 199340
rect 200868 199276 200869 199340
rect 200803 199275 200869 199276
rect 200619 199068 200685 199069
rect 200619 199004 200620 199068
rect 200684 199004 200685 199068
rect 200619 199003 200685 199004
rect 199794 165218 199826 165454
rect 200062 165218 200146 165454
rect 200382 165218 200414 165454
rect 199794 165134 200414 165218
rect 199794 164898 199826 165134
rect 200062 164898 200146 165134
rect 200382 164898 200414 165134
rect 199794 129454 200414 164898
rect 199794 129218 199826 129454
rect 200062 129218 200146 129454
rect 200382 129218 200414 129454
rect 199794 129134 200414 129218
rect 199794 128898 199826 129134
rect 200062 128898 200146 129134
rect 200382 128898 200414 129134
rect 199794 93454 200414 128898
rect 199794 93218 199826 93454
rect 200062 93218 200146 93454
rect 200382 93218 200414 93454
rect 199794 93134 200414 93218
rect 199794 92898 199826 93134
rect 200062 92898 200146 93134
rect 200382 92898 200414 93134
rect 199147 66468 199213 66469
rect 199147 66404 199148 66468
rect 199212 66404 199213 66468
rect 199147 66403 199213 66404
rect 198963 64836 199029 64837
rect 198963 64772 198964 64836
rect 199028 64772 199029 64836
rect 198963 64771 199029 64772
rect 199794 57454 200414 92898
rect 200622 69597 200682 199003
rect 200806 80069 200866 199275
rect 201539 198932 201605 198933
rect 201539 198868 201540 198932
rect 201604 198868 201605 198932
rect 201539 198867 201605 198868
rect 200987 149156 201053 149157
rect 200987 149092 200988 149156
rect 201052 149092 201053 149156
rect 200987 149091 201053 149092
rect 200803 80068 200869 80069
rect 200803 80004 200804 80068
rect 200868 80004 200869 80068
rect 200803 80003 200869 80004
rect 200619 69596 200685 69597
rect 200619 69532 200620 69596
rect 200684 69532 200685 69596
rect 200619 69531 200685 69532
rect 200990 61437 201050 149091
rect 201171 138684 201237 138685
rect 201171 138620 201172 138684
rect 201236 138620 201237 138684
rect 201171 138619 201237 138620
rect 200987 61436 201053 61437
rect 200987 61372 200988 61436
rect 201052 61372 201053 61436
rect 200987 61371 201053 61372
rect 199794 57218 199826 57454
rect 200062 57218 200146 57454
rect 200382 57218 200414 57454
rect 199794 57134 200414 57218
rect 199794 56898 199826 57134
rect 200062 56898 200146 57134
rect 200382 56898 200414 57134
rect 198779 46884 198845 46885
rect 198779 46820 198780 46884
rect 198844 46820 198845 46884
rect 198779 46819 198845 46820
rect 195294 16718 195326 16954
rect 195562 16718 195646 16954
rect 195882 16718 195914 16954
rect 195294 16634 195914 16718
rect 195294 16398 195326 16634
rect 195562 16398 195646 16634
rect 195882 16398 195914 16634
rect 195294 -3226 195914 16398
rect 195294 -3462 195326 -3226
rect 195562 -3462 195646 -3226
rect 195882 -3462 195914 -3226
rect 195294 -3546 195914 -3462
rect 195294 -3782 195326 -3546
rect 195562 -3782 195646 -3546
rect 195882 -3782 195914 -3546
rect 195294 -7654 195914 -3782
rect 199794 21454 200414 56898
rect 201174 53141 201234 138619
rect 201542 67557 201602 198867
rect 201723 195668 201789 195669
rect 201723 195604 201724 195668
rect 201788 195604 201789 195668
rect 201723 195603 201789 195604
rect 201726 71093 201786 195603
rect 203011 194308 203077 194309
rect 203011 194244 203012 194308
rect 203076 194244 203077 194308
rect 203011 194243 203077 194244
rect 203014 161490 203074 194243
rect 202830 161430 203074 161490
rect 204294 169954 204914 205398
rect 208794 710598 209414 711590
rect 208794 710362 208826 710598
rect 209062 710362 209146 710598
rect 209382 710362 209414 710598
rect 208794 710278 209414 710362
rect 208794 710042 208826 710278
rect 209062 710042 209146 710278
rect 209382 710042 209414 710278
rect 208794 678454 209414 710042
rect 208794 678218 208826 678454
rect 209062 678218 209146 678454
rect 209382 678218 209414 678454
rect 208794 678134 209414 678218
rect 208794 677898 208826 678134
rect 209062 677898 209146 678134
rect 209382 677898 209414 678134
rect 208794 642454 209414 677898
rect 208794 642218 208826 642454
rect 209062 642218 209146 642454
rect 209382 642218 209414 642454
rect 208794 642134 209414 642218
rect 208794 641898 208826 642134
rect 209062 641898 209146 642134
rect 209382 641898 209414 642134
rect 208794 606454 209414 641898
rect 208794 606218 208826 606454
rect 209062 606218 209146 606454
rect 209382 606218 209414 606454
rect 208794 606134 209414 606218
rect 208794 605898 208826 606134
rect 209062 605898 209146 606134
rect 209382 605898 209414 606134
rect 208794 570454 209414 605898
rect 208794 570218 208826 570454
rect 209062 570218 209146 570454
rect 209382 570218 209414 570454
rect 208794 570134 209414 570218
rect 208794 569898 208826 570134
rect 209062 569898 209146 570134
rect 209382 569898 209414 570134
rect 208794 534454 209414 569898
rect 208794 534218 208826 534454
rect 209062 534218 209146 534454
rect 209382 534218 209414 534454
rect 208794 534134 209414 534218
rect 208794 533898 208826 534134
rect 209062 533898 209146 534134
rect 209382 533898 209414 534134
rect 208794 498454 209414 533898
rect 208794 498218 208826 498454
rect 209062 498218 209146 498454
rect 209382 498218 209414 498454
rect 208794 498134 209414 498218
rect 208794 497898 208826 498134
rect 209062 497898 209146 498134
rect 209382 497898 209414 498134
rect 208794 462454 209414 497898
rect 208794 462218 208826 462454
rect 209062 462218 209146 462454
rect 209382 462218 209414 462454
rect 208794 462134 209414 462218
rect 208794 461898 208826 462134
rect 209062 461898 209146 462134
rect 209382 461898 209414 462134
rect 208794 426454 209414 461898
rect 208794 426218 208826 426454
rect 209062 426218 209146 426454
rect 209382 426218 209414 426454
rect 208794 426134 209414 426218
rect 208794 425898 208826 426134
rect 209062 425898 209146 426134
rect 209382 425898 209414 426134
rect 208794 390454 209414 425898
rect 208794 390218 208826 390454
rect 209062 390218 209146 390454
rect 209382 390218 209414 390454
rect 208794 390134 209414 390218
rect 208794 389898 208826 390134
rect 209062 389898 209146 390134
rect 209382 389898 209414 390134
rect 208794 354454 209414 389898
rect 208794 354218 208826 354454
rect 209062 354218 209146 354454
rect 209382 354218 209414 354454
rect 208794 354134 209414 354218
rect 208794 353898 208826 354134
rect 209062 353898 209146 354134
rect 209382 353898 209414 354134
rect 208794 318454 209414 353898
rect 208794 318218 208826 318454
rect 209062 318218 209146 318454
rect 209382 318218 209414 318454
rect 208794 318134 209414 318218
rect 208794 317898 208826 318134
rect 209062 317898 209146 318134
rect 209382 317898 209414 318134
rect 208794 282454 209414 317898
rect 208794 282218 208826 282454
rect 209062 282218 209146 282454
rect 209382 282218 209414 282454
rect 208794 282134 209414 282218
rect 208794 281898 208826 282134
rect 209062 281898 209146 282134
rect 209382 281898 209414 282134
rect 208794 246454 209414 281898
rect 208794 246218 208826 246454
rect 209062 246218 209146 246454
rect 209382 246218 209414 246454
rect 208794 246134 209414 246218
rect 208794 245898 208826 246134
rect 209062 245898 209146 246134
rect 209382 245898 209414 246134
rect 208794 210454 209414 245898
rect 208794 210218 208826 210454
rect 209062 210218 209146 210454
rect 209382 210218 209414 210454
rect 208794 210134 209414 210218
rect 208794 209898 208826 210134
rect 209062 209898 209146 210134
rect 209382 209898 209414 210134
rect 205587 193084 205653 193085
rect 205587 193020 205588 193084
rect 205652 193020 205653 193084
rect 205587 193019 205653 193020
rect 204294 169718 204326 169954
rect 204562 169718 204646 169954
rect 204882 169718 204914 169954
rect 204294 169634 204914 169718
rect 204294 169398 204326 169634
rect 204562 169398 204646 169634
rect 204882 169398 204914 169634
rect 201907 148884 201973 148885
rect 201907 148820 201908 148884
rect 201972 148820 201973 148884
rect 201907 148819 201973 148820
rect 201910 72725 201970 148819
rect 202091 139500 202157 139501
rect 202091 139436 202092 139500
rect 202156 139436 202157 139500
rect 202091 139435 202157 139436
rect 201907 72724 201973 72725
rect 201907 72660 201908 72724
rect 201972 72660 201973 72724
rect 201907 72659 201973 72660
rect 201723 71092 201789 71093
rect 201723 71028 201724 71092
rect 201788 71028 201789 71092
rect 201723 71027 201789 71028
rect 201539 67556 201605 67557
rect 201539 67492 201540 67556
rect 201604 67492 201605 67556
rect 201539 67491 201605 67492
rect 202094 62117 202154 139435
rect 202091 62116 202157 62117
rect 202091 62052 202092 62116
rect 202156 62052 202157 62116
rect 202091 62051 202157 62052
rect 201171 53140 201237 53141
rect 201171 53076 201172 53140
rect 201236 53076 201237 53140
rect 201171 53075 201237 53076
rect 202830 47973 202890 161430
rect 203011 156772 203077 156773
rect 203011 156708 203012 156772
rect 203076 156708 203077 156772
rect 203011 156707 203077 156708
rect 203014 48245 203074 156707
rect 203195 156636 203261 156637
rect 203195 156572 203196 156636
rect 203260 156572 203261 156636
rect 203195 156571 203261 156572
rect 203198 57765 203258 156571
rect 203379 148612 203445 148613
rect 203379 148548 203380 148612
rect 203444 148548 203445 148612
rect 203379 148547 203445 148548
rect 203382 59941 203442 148547
rect 204294 133954 204914 169398
rect 204294 133718 204326 133954
rect 204562 133718 204646 133954
rect 204882 133718 204914 133954
rect 204294 133634 204914 133718
rect 204294 133398 204326 133634
rect 204562 133398 204646 133634
rect 204882 133398 204914 133634
rect 204294 97954 204914 133398
rect 204294 97718 204326 97954
rect 204562 97718 204646 97954
rect 204882 97718 204914 97954
rect 204294 97634 204914 97718
rect 204294 97398 204326 97634
rect 204562 97398 204646 97634
rect 204882 97398 204914 97634
rect 204294 61954 204914 97398
rect 205590 75853 205650 193019
rect 208794 174454 209414 209898
rect 213294 711558 213914 711590
rect 213294 711322 213326 711558
rect 213562 711322 213646 711558
rect 213882 711322 213914 711558
rect 213294 711238 213914 711322
rect 213294 711002 213326 711238
rect 213562 711002 213646 711238
rect 213882 711002 213914 711238
rect 213294 682954 213914 711002
rect 213294 682718 213326 682954
rect 213562 682718 213646 682954
rect 213882 682718 213914 682954
rect 213294 682634 213914 682718
rect 213294 682398 213326 682634
rect 213562 682398 213646 682634
rect 213882 682398 213914 682634
rect 213294 646954 213914 682398
rect 213294 646718 213326 646954
rect 213562 646718 213646 646954
rect 213882 646718 213914 646954
rect 213294 646634 213914 646718
rect 213294 646398 213326 646634
rect 213562 646398 213646 646634
rect 213882 646398 213914 646634
rect 213294 610954 213914 646398
rect 213294 610718 213326 610954
rect 213562 610718 213646 610954
rect 213882 610718 213914 610954
rect 213294 610634 213914 610718
rect 213294 610398 213326 610634
rect 213562 610398 213646 610634
rect 213882 610398 213914 610634
rect 213294 574954 213914 610398
rect 213294 574718 213326 574954
rect 213562 574718 213646 574954
rect 213882 574718 213914 574954
rect 213294 574634 213914 574718
rect 213294 574398 213326 574634
rect 213562 574398 213646 574634
rect 213882 574398 213914 574634
rect 213294 538954 213914 574398
rect 213294 538718 213326 538954
rect 213562 538718 213646 538954
rect 213882 538718 213914 538954
rect 213294 538634 213914 538718
rect 213294 538398 213326 538634
rect 213562 538398 213646 538634
rect 213882 538398 213914 538634
rect 213294 502954 213914 538398
rect 213294 502718 213326 502954
rect 213562 502718 213646 502954
rect 213882 502718 213914 502954
rect 213294 502634 213914 502718
rect 213294 502398 213326 502634
rect 213562 502398 213646 502634
rect 213882 502398 213914 502634
rect 213294 466954 213914 502398
rect 213294 466718 213326 466954
rect 213562 466718 213646 466954
rect 213882 466718 213914 466954
rect 213294 466634 213914 466718
rect 213294 466398 213326 466634
rect 213562 466398 213646 466634
rect 213882 466398 213914 466634
rect 213294 430954 213914 466398
rect 213294 430718 213326 430954
rect 213562 430718 213646 430954
rect 213882 430718 213914 430954
rect 213294 430634 213914 430718
rect 213294 430398 213326 430634
rect 213562 430398 213646 430634
rect 213882 430398 213914 430634
rect 213294 394954 213914 430398
rect 213294 394718 213326 394954
rect 213562 394718 213646 394954
rect 213882 394718 213914 394954
rect 213294 394634 213914 394718
rect 213294 394398 213326 394634
rect 213562 394398 213646 394634
rect 213882 394398 213914 394634
rect 213294 358954 213914 394398
rect 213294 358718 213326 358954
rect 213562 358718 213646 358954
rect 213882 358718 213914 358954
rect 213294 358634 213914 358718
rect 213294 358398 213326 358634
rect 213562 358398 213646 358634
rect 213882 358398 213914 358634
rect 213294 322954 213914 358398
rect 213294 322718 213326 322954
rect 213562 322718 213646 322954
rect 213882 322718 213914 322954
rect 213294 322634 213914 322718
rect 213294 322398 213326 322634
rect 213562 322398 213646 322634
rect 213882 322398 213914 322634
rect 213294 286954 213914 322398
rect 213294 286718 213326 286954
rect 213562 286718 213646 286954
rect 213882 286718 213914 286954
rect 213294 286634 213914 286718
rect 213294 286398 213326 286634
rect 213562 286398 213646 286634
rect 213882 286398 213914 286634
rect 213294 250954 213914 286398
rect 213294 250718 213326 250954
rect 213562 250718 213646 250954
rect 213882 250718 213914 250954
rect 213294 250634 213914 250718
rect 213294 250398 213326 250634
rect 213562 250398 213646 250634
rect 213882 250398 213914 250634
rect 213294 214954 213914 250398
rect 213294 214718 213326 214954
rect 213562 214718 213646 214954
rect 213882 214718 213914 214954
rect 213294 214634 213914 214718
rect 213294 214398 213326 214634
rect 213562 214398 213646 214634
rect 213882 214398 213914 214634
rect 209819 194036 209885 194037
rect 209819 193972 209820 194036
rect 209884 193972 209885 194036
rect 209819 193971 209885 193972
rect 208794 174218 208826 174454
rect 209062 174218 209146 174454
rect 209382 174218 209414 174454
rect 208794 174134 209414 174218
rect 208794 173898 208826 174134
rect 209062 173898 209146 174134
rect 209382 173898 209414 174134
rect 207059 151468 207125 151469
rect 207059 151404 207060 151468
rect 207124 151404 207125 151468
rect 207059 151403 207125 151404
rect 205955 151332 206021 151333
rect 205955 151268 205956 151332
rect 206020 151268 206021 151332
rect 205955 151267 206021 151268
rect 205771 148476 205837 148477
rect 205771 148412 205772 148476
rect 205836 148412 205837 148476
rect 205771 148411 205837 148412
rect 205587 75852 205653 75853
rect 205587 75788 205588 75852
rect 205652 75788 205653 75852
rect 205587 75787 205653 75788
rect 205774 71501 205834 148411
rect 205958 81157 206018 151267
rect 205955 81156 206021 81157
rect 205955 81092 205956 81156
rect 206020 81092 206021 81156
rect 205955 81091 206021 81092
rect 205771 71500 205837 71501
rect 205771 71436 205772 71500
rect 205836 71436 205837 71500
rect 205771 71435 205837 71436
rect 205774 71229 205834 71435
rect 205771 71228 205837 71229
rect 205771 71164 205772 71228
rect 205836 71164 205837 71228
rect 205771 71163 205837 71164
rect 204294 61718 204326 61954
rect 204562 61718 204646 61954
rect 204882 61718 204914 61954
rect 204294 61634 204914 61718
rect 204294 61398 204326 61634
rect 204562 61398 204646 61634
rect 204882 61398 204914 61634
rect 203379 59940 203445 59941
rect 203379 59876 203380 59940
rect 203444 59876 203445 59940
rect 203379 59875 203445 59876
rect 203195 57764 203261 57765
rect 203195 57700 203196 57764
rect 203260 57700 203261 57764
rect 203195 57699 203261 57700
rect 203011 48244 203077 48245
rect 203011 48180 203012 48244
rect 203076 48180 203077 48244
rect 203011 48179 203077 48180
rect 202827 47972 202893 47973
rect 202827 47908 202828 47972
rect 202892 47908 202893 47972
rect 202827 47907 202893 47908
rect 204115 47972 204181 47973
rect 204115 47908 204116 47972
rect 204180 47908 204181 47972
rect 204115 47907 204181 47908
rect 204118 47701 204178 47907
rect 204115 47700 204181 47701
rect 204115 47636 204116 47700
rect 204180 47636 204181 47700
rect 204115 47635 204181 47636
rect 199794 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 200414 21454
rect 199794 21134 200414 21218
rect 199794 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 200414 21134
rect 199794 -4186 200414 20898
rect 199794 -4422 199826 -4186
rect 200062 -4422 200146 -4186
rect 200382 -4422 200414 -4186
rect 199794 -4506 200414 -4422
rect 199794 -4742 199826 -4506
rect 200062 -4742 200146 -4506
rect 200382 -4742 200414 -4506
rect 199794 -7654 200414 -4742
rect 204294 25954 204914 61398
rect 207062 44165 207122 151403
rect 207243 151196 207309 151197
rect 207243 151132 207244 151196
rect 207308 151132 207309 151196
rect 207243 151131 207309 151132
rect 207246 46613 207306 151131
rect 208794 138454 209414 173898
rect 208794 138218 208826 138454
rect 209062 138218 209146 138454
rect 209382 138218 209414 138454
rect 208794 138134 209414 138218
rect 208794 137898 208826 138134
rect 209062 137898 209146 138134
rect 209382 137898 209414 138134
rect 208794 102454 209414 137898
rect 208794 102218 208826 102454
rect 209062 102218 209146 102454
rect 209382 102218 209414 102454
rect 208794 102134 209414 102218
rect 208794 101898 208826 102134
rect 209062 101898 209146 102134
rect 209382 101898 209414 102134
rect 208794 66454 209414 101898
rect 208794 66218 208826 66454
rect 209062 66218 209146 66454
rect 209382 66218 209414 66454
rect 208794 66134 209414 66218
rect 208794 65898 208826 66134
rect 209062 65898 209146 66134
rect 209382 65898 209414 66134
rect 207243 46612 207309 46613
rect 207243 46548 207244 46612
rect 207308 46548 207309 46612
rect 207243 46547 207309 46548
rect 207059 44164 207125 44165
rect 207059 44100 207060 44164
rect 207124 44100 207125 44164
rect 207059 44099 207125 44100
rect 204294 25718 204326 25954
rect 204562 25718 204646 25954
rect 204882 25718 204914 25954
rect 204294 25634 204914 25718
rect 204294 25398 204326 25634
rect 204562 25398 204646 25634
rect 204882 25398 204914 25634
rect 204294 -5146 204914 25398
rect 204294 -5382 204326 -5146
rect 204562 -5382 204646 -5146
rect 204882 -5382 204914 -5146
rect 204294 -5466 204914 -5382
rect 204294 -5702 204326 -5466
rect 204562 -5702 204646 -5466
rect 204882 -5702 204914 -5466
rect 204294 -7654 204914 -5702
rect 208794 30454 209414 65898
rect 209822 54501 209882 193971
rect 210003 189956 210069 189957
rect 210003 189892 210004 189956
rect 210068 189892 210069 189956
rect 210003 189891 210069 189892
rect 209819 54500 209885 54501
rect 209819 54436 209820 54500
rect 209884 54436 209885 54500
rect 209819 54435 209885 54436
rect 210006 50693 210066 189891
rect 213294 178954 213914 214398
rect 213294 178718 213326 178954
rect 213562 178718 213646 178954
rect 213882 178718 213914 178954
rect 213294 178634 213914 178718
rect 213294 178398 213326 178634
rect 213562 178398 213646 178634
rect 213882 178398 213914 178634
rect 211291 153916 211357 153917
rect 211291 153852 211292 153916
rect 211356 153852 211357 153916
rect 211291 153851 211357 153852
rect 211107 153780 211173 153781
rect 211107 153716 211108 153780
rect 211172 153716 211173 153780
rect 211107 153715 211173 153716
rect 211110 78165 211170 153715
rect 211294 78437 211354 153851
rect 213294 142954 213914 178398
rect 213294 142718 213326 142954
rect 213562 142718 213646 142954
rect 213882 142718 213914 142954
rect 213294 142634 213914 142718
rect 213294 142398 213326 142634
rect 213562 142398 213646 142634
rect 213882 142398 213914 142634
rect 213294 106954 213914 142398
rect 213294 106718 213326 106954
rect 213562 106718 213646 106954
rect 213882 106718 213914 106954
rect 213294 106634 213914 106718
rect 213294 106398 213326 106634
rect 213562 106398 213646 106634
rect 213882 106398 213914 106634
rect 211291 78436 211357 78437
rect 211291 78372 211292 78436
rect 211356 78372 211357 78436
rect 211291 78371 211357 78372
rect 211107 78164 211173 78165
rect 211107 78100 211108 78164
rect 211172 78100 211173 78164
rect 211107 78099 211173 78100
rect 213294 70954 213914 106398
rect 213294 70718 213326 70954
rect 213562 70718 213646 70954
rect 213882 70718 213914 70954
rect 213294 70634 213914 70718
rect 213294 70398 213326 70634
rect 213562 70398 213646 70634
rect 213882 70398 213914 70634
rect 210003 50692 210069 50693
rect 210003 50628 210004 50692
rect 210068 50628 210069 50692
rect 210003 50627 210069 50628
rect 211107 50692 211173 50693
rect 211107 50628 211108 50692
rect 211172 50628 211173 50692
rect 211107 50627 211173 50628
rect 211110 50285 211170 50627
rect 211107 50284 211173 50285
rect 211107 50220 211108 50284
rect 211172 50220 211173 50284
rect 211107 50219 211173 50220
rect 208794 30218 208826 30454
rect 209062 30218 209146 30454
rect 209382 30218 209414 30454
rect 208794 30134 209414 30218
rect 208794 29898 208826 30134
rect 209062 29898 209146 30134
rect 209382 29898 209414 30134
rect 208794 -6106 209414 29898
rect 208794 -6342 208826 -6106
rect 209062 -6342 209146 -6106
rect 209382 -6342 209414 -6106
rect 208794 -6426 209414 -6342
rect 208794 -6662 208826 -6426
rect 209062 -6662 209146 -6426
rect 209382 -6662 209414 -6426
rect 208794 -7654 209414 -6662
rect 213294 34954 213914 70398
rect 213294 34718 213326 34954
rect 213562 34718 213646 34954
rect 213882 34718 213914 34954
rect 213294 34634 213914 34718
rect 213294 34398 213326 34634
rect 213562 34398 213646 34634
rect 213882 34398 213914 34634
rect 213294 -7066 213914 34398
rect 213294 -7302 213326 -7066
rect 213562 -7302 213646 -7066
rect 213882 -7302 213914 -7066
rect 213294 -7386 213914 -7302
rect 213294 -7622 213326 -7386
rect 213562 -7622 213646 -7386
rect 213882 -7622 213914 -7386
rect 213294 -7654 213914 -7622
rect 217794 704838 218414 711590
rect 217794 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 218414 704838
rect 217794 704518 218414 704602
rect 217794 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 218414 704518
rect 217794 687454 218414 704282
rect 217794 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 218414 687454
rect 217794 687134 218414 687218
rect 217794 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 218414 687134
rect 217794 651454 218414 686898
rect 217794 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 218414 651454
rect 217794 651134 218414 651218
rect 217794 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 218414 651134
rect 217794 615454 218414 650898
rect 217794 615218 217826 615454
rect 218062 615218 218146 615454
rect 218382 615218 218414 615454
rect 217794 615134 218414 615218
rect 217794 614898 217826 615134
rect 218062 614898 218146 615134
rect 218382 614898 218414 615134
rect 217794 579454 218414 614898
rect 217794 579218 217826 579454
rect 218062 579218 218146 579454
rect 218382 579218 218414 579454
rect 217794 579134 218414 579218
rect 217794 578898 217826 579134
rect 218062 578898 218146 579134
rect 218382 578898 218414 579134
rect 217794 543454 218414 578898
rect 217794 543218 217826 543454
rect 218062 543218 218146 543454
rect 218382 543218 218414 543454
rect 217794 543134 218414 543218
rect 217794 542898 217826 543134
rect 218062 542898 218146 543134
rect 218382 542898 218414 543134
rect 217794 507454 218414 542898
rect 217794 507218 217826 507454
rect 218062 507218 218146 507454
rect 218382 507218 218414 507454
rect 217794 507134 218414 507218
rect 217794 506898 217826 507134
rect 218062 506898 218146 507134
rect 218382 506898 218414 507134
rect 217794 471454 218414 506898
rect 217794 471218 217826 471454
rect 218062 471218 218146 471454
rect 218382 471218 218414 471454
rect 217794 471134 218414 471218
rect 217794 470898 217826 471134
rect 218062 470898 218146 471134
rect 218382 470898 218414 471134
rect 217794 435454 218414 470898
rect 217794 435218 217826 435454
rect 218062 435218 218146 435454
rect 218382 435218 218414 435454
rect 217794 435134 218414 435218
rect 217794 434898 217826 435134
rect 218062 434898 218146 435134
rect 218382 434898 218414 435134
rect 217794 399454 218414 434898
rect 217794 399218 217826 399454
rect 218062 399218 218146 399454
rect 218382 399218 218414 399454
rect 217794 399134 218414 399218
rect 217794 398898 217826 399134
rect 218062 398898 218146 399134
rect 218382 398898 218414 399134
rect 217794 363454 218414 398898
rect 217794 363218 217826 363454
rect 218062 363218 218146 363454
rect 218382 363218 218414 363454
rect 217794 363134 218414 363218
rect 217794 362898 217826 363134
rect 218062 362898 218146 363134
rect 218382 362898 218414 363134
rect 217794 327454 218414 362898
rect 217794 327218 217826 327454
rect 218062 327218 218146 327454
rect 218382 327218 218414 327454
rect 217794 327134 218414 327218
rect 217794 326898 217826 327134
rect 218062 326898 218146 327134
rect 218382 326898 218414 327134
rect 217794 291454 218414 326898
rect 217794 291218 217826 291454
rect 218062 291218 218146 291454
rect 218382 291218 218414 291454
rect 217794 291134 218414 291218
rect 217794 290898 217826 291134
rect 218062 290898 218146 291134
rect 218382 290898 218414 291134
rect 217794 255454 218414 290898
rect 217794 255218 217826 255454
rect 218062 255218 218146 255454
rect 218382 255218 218414 255454
rect 217794 255134 218414 255218
rect 217794 254898 217826 255134
rect 218062 254898 218146 255134
rect 218382 254898 218414 255134
rect 217794 219454 218414 254898
rect 217794 219218 217826 219454
rect 218062 219218 218146 219454
rect 218382 219218 218414 219454
rect 217794 219134 218414 219218
rect 217794 218898 217826 219134
rect 218062 218898 218146 219134
rect 218382 218898 218414 219134
rect 217794 183454 218414 218898
rect 217794 183218 217826 183454
rect 218062 183218 218146 183454
rect 218382 183218 218414 183454
rect 217794 183134 218414 183218
rect 217794 182898 217826 183134
rect 218062 182898 218146 183134
rect 218382 182898 218414 183134
rect 217794 147454 218414 182898
rect 217794 147218 217826 147454
rect 218062 147218 218146 147454
rect 218382 147218 218414 147454
rect 217794 147134 218414 147218
rect 217794 146898 217826 147134
rect 218062 146898 218146 147134
rect 218382 146898 218414 147134
rect 217794 111454 218414 146898
rect 217794 111218 217826 111454
rect 218062 111218 218146 111454
rect 218382 111218 218414 111454
rect 217794 111134 218414 111218
rect 217794 110898 217826 111134
rect 218062 110898 218146 111134
rect 218382 110898 218414 111134
rect 217794 75454 218414 110898
rect 217794 75218 217826 75454
rect 218062 75218 218146 75454
rect 218382 75218 218414 75454
rect 217794 75134 218414 75218
rect 217794 74898 217826 75134
rect 218062 74898 218146 75134
rect 218382 74898 218414 75134
rect 217794 39454 218414 74898
rect 217794 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 218414 39454
rect 217794 39134 218414 39218
rect 217794 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 218414 39134
rect 217794 3454 218414 38898
rect 217794 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 218414 3454
rect 217794 3134 218414 3218
rect 217794 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 218414 3134
rect 217794 -346 218414 2898
rect 217794 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 218414 -346
rect 217794 -666 218414 -582
rect 217794 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 218414 -666
rect 217794 -7654 218414 -902
rect 222294 705798 222914 711590
rect 222294 705562 222326 705798
rect 222562 705562 222646 705798
rect 222882 705562 222914 705798
rect 222294 705478 222914 705562
rect 222294 705242 222326 705478
rect 222562 705242 222646 705478
rect 222882 705242 222914 705478
rect 222294 691954 222914 705242
rect 222294 691718 222326 691954
rect 222562 691718 222646 691954
rect 222882 691718 222914 691954
rect 222294 691634 222914 691718
rect 222294 691398 222326 691634
rect 222562 691398 222646 691634
rect 222882 691398 222914 691634
rect 222294 655954 222914 691398
rect 222294 655718 222326 655954
rect 222562 655718 222646 655954
rect 222882 655718 222914 655954
rect 222294 655634 222914 655718
rect 222294 655398 222326 655634
rect 222562 655398 222646 655634
rect 222882 655398 222914 655634
rect 222294 619954 222914 655398
rect 222294 619718 222326 619954
rect 222562 619718 222646 619954
rect 222882 619718 222914 619954
rect 222294 619634 222914 619718
rect 222294 619398 222326 619634
rect 222562 619398 222646 619634
rect 222882 619398 222914 619634
rect 222294 583954 222914 619398
rect 222294 583718 222326 583954
rect 222562 583718 222646 583954
rect 222882 583718 222914 583954
rect 222294 583634 222914 583718
rect 222294 583398 222326 583634
rect 222562 583398 222646 583634
rect 222882 583398 222914 583634
rect 222294 547954 222914 583398
rect 222294 547718 222326 547954
rect 222562 547718 222646 547954
rect 222882 547718 222914 547954
rect 222294 547634 222914 547718
rect 222294 547398 222326 547634
rect 222562 547398 222646 547634
rect 222882 547398 222914 547634
rect 222294 511954 222914 547398
rect 222294 511718 222326 511954
rect 222562 511718 222646 511954
rect 222882 511718 222914 511954
rect 222294 511634 222914 511718
rect 222294 511398 222326 511634
rect 222562 511398 222646 511634
rect 222882 511398 222914 511634
rect 222294 475954 222914 511398
rect 222294 475718 222326 475954
rect 222562 475718 222646 475954
rect 222882 475718 222914 475954
rect 222294 475634 222914 475718
rect 222294 475398 222326 475634
rect 222562 475398 222646 475634
rect 222882 475398 222914 475634
rect 222294 439954 222914 475398
rect 222294 439718 222326 439954
rect 222562 439718 222646 439954
rect 222882 439718 222914 439954
rect 222294 439634 222914 439718
rect 222294 439398 222326 439634
rect 222562 439398 222646 439634
rect 222882 439398 222914 439634
rect 222294 403954 222914 439398
rect 222294 403718 222326 403954
rect 222562 403718 222646 403954
rect 222882 403718 222914 403954
rect 222294 403634 222914 403718
rect 222294 403398 222326 403634
rect 222562 403398 222646 403634
rect 222882 403398 222914 403634
rect 222294 367954 222914 403398
rect 222294 367718 222326 367954
rect 222562 367718 222646 367954
rect 222882 367718 222914 367954
rect 222294 367634 222914 367718
rect 222294 367398 222326 367634
rect 222562 367398 222646 367634
rect 222882 367398 222914 367634
rect 222294 331954 222914 367398
rect 222294 331718 222326 331954
rect 222562 331718 222646 331954
rect 222882 331718 222914 331954
rect 222294 331634 222914 331718
rect 222294 331398 222326 331634
rect 222562 331398 222646 331634
rect 222882 331398 222914 331634
rect 222294 295954 222914 331398
rect 222294 295718 222326 295954
rect 222562 295718 222646 295954
rect 222882 295718 222914 295954
rect 222294 295634 222914 295718
rect 222294 295398 222326 295634
rect 222562 295398 222646 295634
rect 222882 295398 222914 295634
rect 222294 259954 222914 295398
rect 222294 259718 222326 259954
rect 222562 259718 222646 259954
rect 222882 259718 222914 259954
rect 222294 259634 222914 259718
rect 222294 259398 222326 259634
rect 222562 259398 222646 259634
rect 222882 259398 222914 259634
rect 222294 223954 222914 259398
rect 222294 223718 222326 223954
rect 222562 223718 222646 223954
rect 222882 223718 222914 223954
rect 222294 223634 222914 223718
rect 222294 223398 222326 223634
rect 222562 223398 222646 223634
rect 222882 223398 222914 223634
rect 222294 187954 222914 223398
rect 222294 187718 222326 187954
rect 222562 187718 222646 187954
rect 222882 187718 222914 187954
rect 222294 187634 222914 187718
rect 222294 187398 222326 187634
rect 222562 187398 222646 187634
rect 222882 187398 222914 187634
rect 222294 151954 222914 187398
rect 222294 151718 222326 151954
rect 222562 151718 222646 151954
rect 222882 151718 222914 151954
rect 222294 151634 222914 151718
rect 222294 151398 222326 151634
rect 222562 151398 222646 151634
rect 222882 151398 222914 151634
rect 222294 115954 222914 151398
rect 222294 115718 222326 115954
rect 222562 115718 222646 115954
rect 222882 115718 222914 115954
rect 222294 115634 222914 115718
rect 222294 115398 222326 115634
rect 222562 115398 222646 115634
rect 222882 115398 222914 115634
rect 222294 79954 222914 115398
rect 222294 79718 222326 79954
rect 222562 79718 222646 79954
rect 222882 79718 222914 79954
rect 222294 79634 222914 79718
rect 222294 79398 222326 79634
rect 222562 79398 222646 79634
rect 222882 79398 222914 79634
rect 222294 43954 222914 79398
rect 222294 43718 222326 43954
rect 222562 43718 222646 43954
rect 222882 43718 222914 43954
rect 222294 43634 222914 43718
rect 222294 43398 222326 43634
rect 222562 43398 222646 43634
rect 222882 43398 222914 43634
rect 222294 7954 222914 43398
rect 222294 7718 222326 7954
rect 222562 7718 222646 7954
rect 222882 7718 222914 7954
rect 222294 7634 222914 7718
rect 222294 7398 222326 7634
rect 222562 7398 222646 7634
rect 222882 7398 222914 7634
rect 222294 -1306 222914 7398
rect 222294 -1542 222326 -1306
rect 222562 -1542 222646 -1306
rect 222882 -1542 222914 -1306
rect 222294 -1626 222914 -1542
rect 222294 -1862 222326 -1626
rect 222562 -1862 222646 -1626
rect 222882 -1862 222914 -1626
rect 222294 -7654 222914 -1862
rect 226794 706758 227414 711590
rect 226794 706522 226826 706758
rect 227062 706522 227146 706758
rect 227382 706522 227414 706758
rect 226794 706438 227414 706522
rect 226794 706202 226826 706438
rect 227062 706202 227146 706438
rect 227382 706202 227414 706438
rect 226794 696454 227414 706202
rect 226794 696218 226826 696454
rect 227062 696218 227146 696454
rect 227382 696218 227414 696454
rect 226794 696134 227414 696218
rect 226794 695898 226826 696134
rect 227062 695898 227146 696134
rect 227382 695898 227414 696134
rect 226794 660454 227414 695898
rect 226794 660218 226826 660454
rect 227062 660218 227146 660454
rect 227382 660218 227414 660454
rect 226794 660134 227414 660218
rect 226794 659898 226826 660134
rect 227062 659898 227146 660134
rect 227382 659898 227414 660134
rect 226794 624454 227414 659898
rect 226794 624218 226826 624454
rect 227062 624218 227146 624454
rect 227382 624218 227414 624454
rect 226794 624134 227414 624218
rect 226794 623898 226826 624134
rect 227062 623898 227146 624134
rect 227382 623898 227414 624134
rect 226794 588454 227414 623898
rect 226794 588218 226826 588454
rect 227062 588218 227146 588454
rect 227382 588218 227414 588454
rect 226794 588134 227414 588218
rect 226794 587898 226826 588134
rect 227062 587898 227146 588134
rect 227382 587898 227414 588134
rect 226794 552454 227414 587898
rect 226794 552218 226826 552454
rect 227062 552218 227146 552454
rect 227382 552218 227414 552454
rect 226794 552134 227414 552218
rect 226794 551898 226826 552134
rect 227062 551898 227146 552134
rect 227382 551898 227414 552134
rect 226794 516454 227414 551898
rect 226794 516218 226826 516454
rect 227062 516218 227146 516454
rect 227382 516218 227414 516454
rect 226794 516134 227414 516218
rect 226794 515898 226826 516134
rect 227062 515898 227146 516134
rect 227382 515898 227414 516134
rect 226794 480454 227414 515898
rect 226794 480218 226826 480454
rect 227062 480218 227146 480454
rect 227382 480218 227414 480454
rect 226794 480134 227414 480218
rect 226794 479898 226826 480134
rect 227062 479898 227146 480134
rect 227382 479898 227414 480134
rect 226794 444454 227414 479898
rect 226794 444218 226826 444454
rect 227062 444218 227146 444454
rect 227382 444218 227414 444454
rect 226794 444134 227414 444218
rect 226794 443898 226826 444134
rect 227062 443898 227146 444134
rect 227382 443898 227414 444134
rect 226794 408454 227414 443898
rect 226794 408218 226826 408454
rect 227062 408218 227146 408454
rect 227382 408218 227414 408454
rect 226794 408134 227414 408218
rect 226794 407898 226826 408134
rect 227062 407898 227146 408134
rect 227382 407898 227414 408134
rect 226794 372454 227414 407898
rect 226794 372218 226826 372454
rect 227062 372218 227146 372454
rect 227382 372218 227414 372454
rect 226794 372134 227414 372218
rect 226794 371898 226826 372134
rect 227062 371898 227146 372134
rect 227382 371898 227414 372134
rect 226794 336454 227414 371898
rect 226794 336218 226826 336454
rect 227062 336218 227146 336454
rect 227382 336218 227414 336454
rect 226794 336134 227414 336218
rect 226794 335898 226826 336134
rect 227062 335898 227146 336134
rect 227382 335898 227414 336134
rect 226794 300454 227414 335898
rect 226794 300218 226826 300454
rect 227062 300218 227146 300454
rect 227382 300218 227414 300454
rect 226794 300134 227414 300218
rect 226794 299898 226826 300134
rect 227062 299898 227146 300134
rect 227382 299898 227414 300134
rect 226794 264454 227414 299898
rect 226794 264218 226826 264454
rect 227062 264218 227146 264454
rect 227382 264218 227414 264454
rect 226794 264134 227414 264218
rect 226794 263898 226826 264134
rect 227062 263898 227146 264134
rect 227382 263898 227414 264134
rect 226794 228454 227414 263898
rect 226794 228218 226826 228454
rect 227062 228218 227146 228454
rect 227382 228218 227414 228454
rect 226794 228134 227414 228218
rect 226794 227898 226826 228134
rect 227062 227898 227146 228134
rect 227382 227898 227414 228134
rect 226794 192454 227414 227898
rect 226794 192218 226826 192454
rect 227062 192218 227146 192454
rect 227382 192218 227414 192454
rect 226794 192134 227414 192218
rect 226794 191898 226826 192134
rect 227062 191898 227146 192134
rect 227382 191898 227414 192134
rect 226794 156454 227414 191898
rect 226794 156218 226826 156454
rect 227062 156218 227146 156454
rect 227382 156218 227414 156454
rect 226794 156134 227414 156218
rect 226794 155898 226826 156134
rect 227062 155898 227146 156134
rect 227382 155898 227414 156134
rect 226794 120454 227414 155898
rect 226794 120218 226826 120454
rect 227062 120218 227146 120454
rect 227382 120218 227414 120454
rect 226794 120134 227414 120218
rect 226794 119898 226826 120134
rect 227062 119898 227146 120134
rect 227382 119898 227414 120134
rect 226794 84454 227414 119898
rect 226794 84218 226826 84454
rect 227062 84218 227146 84454
rect 227382 84218 227414 84454
rect 226794 84134 227414 84218
rect 226794 83898 226826 84134
rect 227062 83898 227146 84134
rect 227382 83898 227414 84134
rect 226794 48454 227414 83898
rect 226794 48218 226826 48454
rect 227062 48218 227146 48454
rect 227382 48218 227414 48454
rect 226794 48134 227414 48218
rect 226794 47898 226826 48134
rect 227062 47898 227146 48134
rect 227382 47898 227414 48134
rect 226794 12454 227414 47898
rect 226794 12218 226826 12454
rect 227062 12218 227146 12454
rect 227382 12218 227414 12454
rect 226794 12134 227414 12218
rect 226794 11898 226826 12134
rect 227062 11898 227146 12134
rect 227382 11898 227414 12134
rect 226794 -2266 227414 11898
rect 226794 -2502 226826 -2266
rect 227062 -2502 227146 -2266
rect 227382 -2502 227414 -2266
rect 226794 -2586 227414 -2502
rect 226794 -2822 226826 -2586
rect 227062 -2822 227146 -2586
rect 227382 -2822 227414 -2586
rect 226794 -7654 227414 -2822
rect 231294 707718 231914 711590
rect 231294 707482 231326 707718
rect 231562 707482 231646 707718
rect 231882 707482 231914 707718
rect 231294 707398 231914 707482
rect 231294 707162 231326 707398
rect 231562 707162 231646 707398
rect 231882 707162 231914 707398
rect 231294 700954 231914 707162
rect 231294 700718 231326 700954
rect 231562 700718 231646 700954
rect 231882 700718 231914 700954
rect 231294 700634 231914 700718
rect 231294 700398 231326 700634
rect 231562 700398 231646 700634
rect 231882 700398 231914 700634
rect 231294 664954 231914 700398
rect 231294 664718 231326 664954
rect 231562 664718 231646 664954
rect 231882 664718 231914 664954
rect 231294 664634 231914 664718
rect 231294 664398 231326 664634
rect 231562 664398 231646 664634
rect 231882 664398 231914 664634
rect 231294 628954 231914 664398
rect 231294 628718 231326 628954
rect 231562 628718 231646 628954
rect 231882 628718 231914 628954
rect 231294 628634 231914 628718
rect 231294 628398 231326 628634
rect 231562 628398 231646 628634
rect 231882 628398 231914 628634
rect 231294 592954 231914 628398
rect 231294 592718 231326 592954
rect 231562 592718 231646 592954
rect 231882 592718 231914 592954
rect 231294 592634 231914 592718
rect 231294 592398 231326 592634
rect 231562 592398 231646 592634
rect 231882 592398 231914 592634
rect 231294 556954 231914 592398
rect 231294 556718 231326 556954
rect 231562 556718 231646 556954
rect 231882 556718 231914 556954
rect 231294 556634 231914 556718
rect 231294 556398 231326 556634
rect 231562 556398 231646 556634
rect 231882 556398 231914 556634
rect 231294 520954 231914 556398
rect 231294 520718 231326 520954
rect 231562 520718 231646 520954
rect 231882 520718 231914 520954
rect 231294 520634 231914 520718
rect 231294 520398 231326 520634
rect 231562 520398 231646 520634
rect 231882 520398 231914 520634
rect 231294 484954 231914 520398
rect 231294 484718 231326 484954
rect 231562 484718 231646 484954
rect 231882 484718 231914 484954
rect 231294 484634 231914 484718
rect 231294 484398 231326 484634
rect 231562 484398 231646 484634
rect 231882 484398 231914 484634
rect 231294 448954 231914 484398
rect 231294 448718 231326 448954
rect 231562 448718 231646 448954
rect 231882 448718 231914 448954
rect 231294 448634 231914 448718
rect 231294 448398 231326 448634
rect 231562 448398 231646 448634
rect 231882 448398 231914 448634
rect 231294 412954 231914 448398
rect 231294 412718 231326 412954
rect 231562 412718 231646 412954
rect 231882 412718 231914 412954
rect 231294 412634 231914 412718
rect 231294 412398 231326 412634
rect 231562 412398 231646 412634
rect 231882 412398 231914 412634
rect 231294 376954 231914 412398
rect 231294 376718 231326 376954
rect 231562 376718 231646 376954
rect 231882 376718 231914 376954
rect 231294 376634 231914 376718
rect 231294 376398 231326 376634
rect 231562 376398 231646 376634
rect 231882 376398 231914 376634
rect 231294 340954 231914 376398
rect 231294 340718 231326 340954
rect 231562 340718 231646 340954
rect 231882 340718 231914 340954
rect 231294 340634 231914 340718
rect 231294 340398 231326 340634
rect 231562 340398 231646 340634
rect 231882 340398 231914 340634
rect 231294 304954 231914 340398
rect 231294 304718 231326 304954
rect 231562 304718 231646 304954
rect 231882 304718 231914 304954
rect 231294 304634 231914 304718
rect 231294 304398 231326 304634
rect 231562 304398 231646 304634
rect 231882 304398 231914 304634
rect 231294 268954 231914 304398
rect 231294 268718 231326 268954
rect 231562 268718 231646 268954
rect 231882 268718 231914 268954
rect 231294 268634 231914 268718
rect 231294 268398 231326 268634
rect 231562 268398 231646 268634
rect 231882 268398 231914 268634
rect 231294 232954 231914 268398
rect 231294 232718 231326 232954
rect 231562 232718 231646 232954
rect 231882 232718 231914 232954
rect 231294 232634 231914 232718
rect 231294 232398 231326 232634
rect 231562 232398 231646 232634
rect 231882 232398 231914 232634
rect 231294 196954 231914 232398
rect 231294 196718 231326 196954
rect 231562 196718 231646 196954
rect 231882 196718 231914 196954
rect 231294 196634 231914 196718
rect 231294 196398 231326 196634
rect 231562 196398 231646 196634
rect 231882 196398 231914 196634
rect 231294 160954 231914 196398
rect 231294 160718 231326 160954
rect 231562 160718 231646 160954
rect 231882 160718 231914 160954
rect 231294 160634 231914 160718
rect 231294 160398 231326 160634
rect 231562 160398 231646 160634
rect 231882 160398 231914 160634
rect 231294 124954 231914 160398
rect 231294 124718 231326 124954
rect 231562 124718 231646 124954
rect 231882 124718 231914 124954
rect 231294 124634 231914 124718
rect 231294 124398 231326 124634
rect 231562 124398 231646 124634
rect 231882 124398 231914 124634
rect 231294 88954 231914 124398
rect 231294 88718 231326 88954
rect 231562 88718 231646 88954
rect 231882 88718 231914 88954
rect 231294 88634 231914 88718
rect 231294 88398 231326 88634
rect 231562 88398 231646 88634
rect 231882 88398 231914 88634
rect 231294 52954 231914 88398
rect 231294 52718 231326 52954
rect 231562 52718 231646 52954
rect 231882 52718 231914 52954
rect 231294 52634 231914 52718
rect 231294 52398 231326 52634
rect 231562 52398 231646 52634
rect 231882 52398 231914 52634
rect 231294 16954 231914 52398
rect 231294 16718 231326 16954
rect 231562 16718 231646 16954
rect 231882 16718 231914 16954
rect 231294 16634 231914 16718
rect 231294 16398 231326 16634
rect 231562 16398 231646 16634
rect 231882 16398 231914 16634
rect 231294 -3226 231914 16398
rect 231294 -3462 231326 -3226
rect 231562 -3462 231646 -3226
rect 231882 -3462 231914 -3226
rect 231294 -3546 231914 -3462
rect 231294 -3782 231326 -3546
rect 231562 -3782 231646 -3546
rect 231882 -3782 231914 -3546
rect 231294 -7654 231914 -3782
rect 235794 708678 236414 711590
rect 235794 708442 235826 708678
rect 236062 708442 236146 708678
rect 236382 708442 236414 708678
rect 235794 708358 236414 708442
rect 235794 708122 235826 708358
rect 236062 708122 236146 708358
rect 236382 708122 236414 708358
rect 235794 669454 236414 708122
rect 235794 669218 235826 669454
rect 236062 669218 236146 669454
rect 236382 669218 236414 669454
rect 235794 669134 236414 669218
rect 235794 668898 235826 669134
rect 236062 668898 236146 669134
rect 236382 668898 236414 669134
rect 235794 633454 236414 668898
rect 235794 633218 235826 633454
rect 236062 633218 236146 633454
rect 236382 633218 236414 633454
rect 235794 633134 236414 633218
rect 235794 632898 235826 633134
rect 236062 632898 236146 633134
rect 236382 632898 236414 633134
rect 235794 597454 236414 632898
rect 235794 597218 235826 597454
rect 236062 597218 236146 597454
rect 236382 597218 236414 597454
rect 235794 597134 236414 597218
rect 235794 596898 235826 597134
rect 236062 596898 236146 597134
rect 236382 596898 236414 597134
rect 235794 561454 236414 596898
rect 235794 561218 235826 561454
rect 236062 561218 236146 561454
rect 236382 561218 236414 561454
rect 235794 561134 236414 561218
rect 235794 560898 235826 561134
rect 236062 560898 236146 561134
rect 236382 560898 236414 561134
rect 235794 525454 236414 560898
rect 235794 525218 235826 525454
rect 236062 525218 236146 525454
rect 236382 525218 236414 525454
rect 235794 525134 236414 525218
rect 235794 524898 235826 525134
rect 236062 524898 236146 525134
rect 236382 524898 236414 525134
rect 235794 489454 236414 524898
rect 235794 489218 235826 489454
rect 236062 489218 236146 489454
rect 236382 489218 236414 489454
rect 235794 489134 236414 489218
rect 235794 488898 235826 489134
rect 236062 488898 236146 489134
rect 236382 488898 236414 489134
rect 235794 453454 236414 488898
rect 235794 453218 235826 453454
rect 236062 453218 236146 453454
rect 236382 453218 236414 453454
rect 235794 453134 236414 453218
rect 235794 452898 235826 453134
rect 236062 452898 236146 453134
rect 236382 452898 236414 453134
rect 235794 417454 236414 452898
rect 235794 417218 235826 417454
rect 236062 417218 236146 417454
rect 236382 417218 236414 417454
rect 235794 417134 236414 417218
rect 235794 416898 235826 417134
rect 236062 416898 236146 417134
rect 236382 416898 236414 417134
rect 235794 381454 236414 416898
rect 235794 381218 235826 381454
rect 236062 381218 236146 381454
rect 236382 381218 236414 381454
rect 235794 381134 236414 381218
rect 235794 380898 235826 381134
rect 236062 380898 236146 381134
rect 236382 380898 236414 381134
rect 235794 345454 236414 380898
rect 235794 345218 235826 345454
rect 236062 345218 236146 345454
rect 236382 345218 236414 345454
rect 235794 345134 236414 345218
rect 235794 344898 235826 345134
rect 236062 344898 236146 345134
rect 236382 344898 236414 345134
rect 235794 309454 236414 344898
rect 235794 309218 235826 309454
rect 236062 309218 236146 309454
rect 236382 309218 236414 309454
rect 235794 309134 236414 309218
rect 235794 308898 235826 309134
rect 236062 308898 236146 309134
rect 236382 308898 236414 309134
rect 235794 273454 236414 308898
rect 235794 273218 235826 273454
rect 236062 273218 236146 273454
rect 236382 273218 236414 273454
rect 235794 273134 236414 273218
rect 235794 272898 235826 273134
rect 236062 272898 236146 273134
rect 236382 272898 236414 273134
rect 235794 237454 236414 272898
rect 235794 237218 235826 237454
rect 236062 237218 236146 237454
rect 236382 237218 236414 237454
rect 235794 237134 236414 237218
rect 235794 236898 235826 237134
rect 236062 236898 236146 237134
rect 236382 236898 236414 237134
rect 235794 201454 236414 236898
rect 235794 201218 235826 201454
rect 236062 201218 236146 201454
rect 236382 201218 236414 201454
rect 235794 201134 236414 201218
rect 235794 200898 235826 201134
rect 236062 200898 236146 201134
rect 236382 200898 236414 201134
rect 235794 165454 236414 200898
rect 235794 165218 235826 165454
rect 236062 165218 236146 165454
rect 236382 165218 236414 165454
rect 235794 165134 236414 165218
rect 235794 164898 235826 165134
rect 236062 164898 236146 165134
rect 236382 164898 236414 165134
rect 235794 129454 236414 164898
rect 235794 129218 235826 129454
rect 236062 129218 236146 129454
rect 236382 129218 236414 129454
rect 235794 129134 236414 129218
rect 235794 128898 235826 129134
rect 236062 128898 236146 129134
rect 236382 128898 236414 129134
rect 235794 93454 236414 128898
rect 235794 93218 235826 93454
rect 236062 93218 236146 93454
rect 236382 93218 236414 93454
rect 235794 93134 236414 93218
rect 235794 92898 235826 93134
rect 236062 92898 236146 93134
rect 236382 92898 236414 93134
rect 235794 57454 236414 92898
rect 235794 57218 235826 57454
rect 236062 57218 236146 57454
rect 236382 57218 236414 57454
rect 235794 57134 236414 57218
rect 235794 56898 235826 57134
rect 236062 56898 236146 57134
rect 236382 56898 236414 57134
rect 235794 21454 236414 56898
rect 235794 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 236414 21454
rect 235794 21134 236414 21218
rect 235794 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 236414 21134
rect 235794 -4186 236414 20898
rect 235794 -4422 235826 -4186
rect 236062 -4422 236146 -4186
rect 236382 -4422 236414 -4186
rect 235794 -4506 236414 -4422
rect 235794 -4742 235826 -4506
rect 236062 -4742 236146 -4506
rect 236382 -4742 236414 -4506
rect 235794 -7654 236414 -4742
rect 240294 709638 240914 711590
rect 240294 709402 240326 709638
rect 240562 709402 240646 709638
rect 240882 709402 240914 709638
rect 240294 709318 240914 709402
rect 240294 709082 240326 709318
rect 240562 709082 240646 709318
rect 240882 709082 240914 709318
rect 240294 673954 240914 709082
rect 240294 673718 240326 673954
rect 240562 673718 240646 673954
rect 240882 673718 240914 673954
rect 240294 673634 240914 673718
rect 240294 673398 240326 673634
rect 240562 673398 240646 673634
rect 240882 673398 240914 673634
rect 240294 637954 240914 673398
rect 240294 637718 240326 637954
rect 240562 637718 240646 637954
rect 240882 637718 240914 637954
rect 240294 637634 240914 637718
rect 240294 637398 240326 637634
rect 240562 637398 240646 637634
rect 240882 637398 240914 637634
rect 240294 601954 240914 637398
rect 240294 601718 240326 601954
rect 240562 601718 240646 601954
rect 240882 601718 240914 601954
rect 240294 601634 240914 601718
rect 240294 601398 240326 601634
rect 240562 601398 240646 601634
rect 240882 601398 240914 601634
rect 240294 565954 240914 601398
rect 240294 565718 240326 565954
rect 240562 565718 240646 565954
rect 240882 565718 240914 565954
rect 240294 565634 240914 565718
rect 240294 565398 240326 565634
rect 240562 565398 240646 565634
rect 240882 565398 240914 565634
rect 240294 529954 240914 565398
rect 240294 529718 240326 529954
rect 240562 529718 240646 529954
rect 240882 529718 240914 529954
rect 240294 529634 240914 529718
rect 240294 529398 240326 529634
rect 240562 529398 240646 529634
rect 240882 529398 240914 529634
rect 240294 493954 240914 529398
rect 240294 493718 240326 493954
rect 240562 493718 240646 493954
rect 240882 493718 240914 493954
rect 240294 493634 240914 493718
rect 240294 493398 240326 493634
rect 240562 493398 240646 493634
rect 240882 493398 240914 493634
rect 240294 457954 240914 493398
rect 240294 457718 240326 457954
rect 240562 457718 240646 457954
rect 240882 457718 240914 457954
rect 240294 457634 240914 457718
rect 240294 457398 240326 457634
rect 240562 457398 240646 457634
rect 240882 457398 240914 457634
rect 240294 421954 240914 457398
rect 240294 421718 240326 421954
rect 240562 421718 240646 421954
rect 240882 421718 240914 421954
rect 240294 421634 240914 421718
rect 240294 421398 240326 421634
rect 240562 421398 240646 421634
rect 240882 421398 240914 421634
rect 240294 385954 240914 421398
rect 240294 385718 240326 385954
rect 240562 385718 240646 385954
rect 240882 385718 240914 385954
rect 240294 385634 240914 385718
rect 240294 385398 240326 385634
rect 240562 385398 240646 385634
rect 240882 385398 240914 385634
rect 240294 349954 240914 385398
rect 240294 349718 240326 349954
rect 240562 349718 240646 349954
rect 240882 349718 240914 349954
rect 240294 349634 240914 349718
rect 240294 349398 240326 349634
rect 240562 349398 240646 349634
rect 240882 349398 240914 349634
rect 240294 313954 240914 349398
rect 240294 313718 240326 313954
rect 240562 313718 240646 313954
rect 240882 313718 240914 313954
rect 240294 313634 240914 313718
rect 240294 313398 240326 313634
rect 240562 313398 240646 313634
rect 240882 313398 240914 313634
rect 240294 277954 240914 313398
rect 240294 277718 240326 277954
rect 240562 277718 240646 277954
rect 240882 277718 240914 277954
rect 240294 277634 240914 277718
rect 240294 277398 240326 277634
rect 240562 277398 240646 277634
rect 240882 277398 240914 277634
rect 240294 241954 240914 277398
rect 240294 241718 240326 241954
rect 240562 241718 240646 241954
rect 240882 241718 240914 241954
rect 240294 241634 240914 241718
rect 240294 241398 240326 241634
rect 240562 241398 240646 241634
rect 240882 241398 240914 241634
rect 240294 205954 240914 241398
rect 240294 205718 240326 205954
rect 240562 205718 240646 205954
rect 240882 205718 240914 205954
rect 240294 205634 240914 205718
rect 240294 205398 240326 205634
rect 240562 205398 240646 205634
rect 240882 205398 240914 205634
rect 240294 169954 240914 205398
rect 240294 169718 240326 169954
rect 240562 169718 240646 169954
rect 240882 169718 240914 169954
rect 240294 169634 240914 169718
rect 240294 169398 240326 169634
rect 240562 169398 240646 169634
rect 240882 169398 240914 169634
rect 240294 133954 240914 169398
rect 240294 133718 240326 133954
rect 240562 133718 240646 133954
rect 240882 133718 240914 133954
rect 240294 133634 240914 133718
rect 240294 133398 240326 133634
rect 240562 133398 240646 133634
rect 240882 133398 240914 133634
rect 240294 97954 240914 133398
rect 240294 97718 240326 97954
rect 240562 97718 240646 97954
rect 240882 97718 240914 97954
rect 240294 97634 240914 97718
rect 240294 97398 240326 97634
rect 240562 97398 240646 97634
rect 240882 97398 240914 97634
rect 240294 61954 240914 97398
rect 240294 61718 240326 61954
rect 240562 61718 240646 61954
rect 240882 61718 240914 61954
rect 240294 61634 240914 61718
rect 240294 61398 240326 61634
rect 240562 61398 240646 61634
rect 240882 61398 240914 61634
rect 240294 25954 240914 61398
rect 240294 25718 240326 25954
rect 240562 25718 240646 25954
rect 240882 25718 240914 25954
rect 240294 25634 240914 25718
rect 240294 25398 240326 25634
rect 240562 25398 240646 25634
rect 240882 25398 240914 25634
rect 240294 -5146 240914 25398
rect 240294 -5382 240326 -5146
rect 240562 -5382 240646 -5146
rect 240882 -5382 240914 -5146
rect 240294 -5466 240914 -5382
rect 240294 -5702 240326 -5466
rect 240562 -5702 240646 -5466
rect 240882 -5702 240914 -5466
rect 240294 -7654 240914 -5702
rect 244794 710598 245414 711590
rect 244794 710362 244826 710598
rect 245062 710362 245146 710598
rect 245382 710362 245414 710598
rect 244794 710278 245414 710362
rect 244794 710042 244826 710278
rect 245062 710042 245146 710278
rect 245382 710042 245414 710278
rect 244794 678454 245414 710042
rect 244794 678218 244826 678454
rect 245062 678218 245146 678454
rect 245382 678218 245414 678454
rect 244794 678134 245414 678218
rect 244794 677898 244826 678134
rect 245062 677898 245146 678134
rect 245382 677898 245414 678134
rect 244794 642454 245414 677898
rect 244794 642218 244826 642454
rect 245062 642218 245146 642454
rect 245382 642218 245414 642454
rect 244794 642134 245414 642218
rect 244794 641898 244826 642134
rect 245062 641898 245146 642134
rect 245382 641898 245414 642134
rect 244794 606454 245414 641898
rect 244794 606218 244826 606454
rect 245062 606218 245146 606454
rect 245382 606218 245414 606454
rect 244794 606134 245414 606218
rect 244794 605898 244826 606134
rect 245062 605898 245146 606134
rect 245382 605898 245414 606134
rect 244794 570454 245414 605898
rect 244794 570218 244826 570454
rect 245062 570218 245146 570454
rect 245382 570218 245414 570454
rect 244794 570134 245414 570218
rect 244794 569898 244826 570134
rect 245062 569898 245146 570134
rect 245382 569898 245414 570134
rect 244794 534454 245414 569898
rect 244794 534218 244826 534454
rect 245062 534218 245146 534454
rect 245382 534218 245414 534454
rect 244794 534134 245414 534218
rect 244794 533898 244826 534134
rect 245062 533898 245146 534134
rect 245382 533898 245414 534134
rect 244794 498454 245414 533898
rect 244794 498218 244826 498454
rect 245062 498218 245146 498454
rect 245382 498218 245414 498454
rect 244794 498134 245414 498218
rect 244794 497898 244826 498134
rect 245062 497898 245146 498134
rect 245382 497898 245414 498134
rect 244794 462454 245414 497898
rect 244794 462218 244826 462454
rect 245062 462218 245146 462454
rect 245382 462218 245414 462454
rect 244794 462134 245414 462218
rect 244794 461898 244826 462134
rect 245062 461898 245146 462134
rect 245382 461898 245414 462134
rect 244794 426454 245414 461898
rect 244794 426218 244826 426454
rect 245062 426218 245146 426454
rect 245382 426218 245414 426454
rect 244794 426134 245414 426218
rect 244794 425898 244826 426134
rect 245062 425898 245146 426134
rect 245382 425898 245414 426134
rect 244794 390454 245414 425898
rect 244794 390218 244826 390454
rect 245062 390218 245146 390454
rect 245382 390218 245414 390454
rect 244794 390134 245414 390218
rect 244794 389898 244826 390134
rect 245062 389898 245146 390134
rect 245382 389898 245414 390134
rect 244794 354454 245414 389898
rect 244794 354218 244826 354454
rect 245062 354218 245146 354454
rect 245382 354218 245414 354454
rect 244794 354134 245414 354218
rect 244794 353898 244826 354134
rect 245062 353898 245146 354134
rect 245382 353898 245414 354134
rect 244794 318454 245414 353898
rect 244794 318218 244826 318454
rect 245062 318218 245146 318454
rect 245382 318218 245414 318454
rect 244794 318134 245414 318218
rect 244794 317898 244826 318134
rect 245062 317898 245146 318134
rect 245382 317898 245414 318134
rect 244794 282454 245414 317898
rect 244794 282218 244826 282454
rect 245062 282218 245146 282454
rect 245382 282218 245414 282454
rect 244794 282134 245414 282218
rect 244794 281898 244826 282134
rect 245062 281898 245146 282134
rect 245382 281898 245414 282134
rect 244794 246454 245414 281898
rect 244794 246218 244826 246454
rect 245062 246218 245146 246454
rect 245382 246218 245414 246454
rect 244794 246134 245414 246218
rect 244794 245898 244826 246134
rect 245062 245898 245146 246134
rect 245382 245898 245414 246134
rect 244794 210454 245414 245898
rect 244794 210218 244826 210454
rect 245062 210218 245146 210454
rect 245382 210218 245414 210454
rect 244794 210134 245414 210218
rect 244794 209898 244826 210134
rect 245062 209898 245146 210134
rect 245382 209898 245414 210134
rect 244794 174454 245414 209898
rect 244794 174218 244826 174454
rect 245062 174218 245146 174454
rect 245382 174218 245414 174454
rect 244794 174134 245414 174218
rect 244794 173898 244826 174134
rect 245062 173898 245146 174134
rect 245382 173898 245414 174134
rect 244794 138454 245414 173898
rect 244794 138218 244826 138454
rect 245062 138218 245146 138454
rect 245382 138218 245414 138454
rect 244794 138134 245414 138218
rect 244794 137898 244826 138134
rect 245062 137898 245146 138134
rect 245382 137898 245414 138134
rect 244794 102454 245414 137898
rect 244794 102218 244826 102454
rect 245062 102218 245146 102454
rect 245382 102218 245414 102454
rect 244794 102134 245414 102218
rect 244794 101898 244826 102134
rect 245062 101898 245146 102134
rect 245382 101898 245414 102134
rect 244794 66454 245414 101898
rect 244794 66218 244826 66454
rect 245062 66218 245146 66454
rect 245382 66218 245414 66454
rect 244794 66134 245414 66218
rect 244794 65898 244826 66134
rect 245062 65898 245146 66134
rect 245382 65898 245414 66134
rect 244794 30454 245414 65898
rect 244794 30218 244826 30454
rect 245062 30218 245146 30454
rect 245382 30218 245414 30454
rect 244794 30134 245414 30218
rect 244794 29898 244826 30134
rect 245062 29898 245146 30134
rect 245382 29898 245414 30134
rect 244794 -6106 245414 29898
rect 244794 -6342 244826 -6106
rect 245062 -6342 245146 -6106
rect 245382 -6342 245414 -6106
rect 244794 -6426 245414 -6342
rect 244794 -6662 244826 -6426
rect 245062 -6662 245146 -6426
rect 245382 -6662 245414 -6426
rect 244794 -7654 245414 -6662
rect 249294 711558 249914 711590
rect 249294 711322 249326 711558
rect 249562 711322 249646 711558
rect 249882 711322 249914 711558
rect 249294 711238 249914 711322
rect 249294 711002 249326 711238
rect 249562 711002 249646 711238
rect 249882 711002 249914 711238
rect 249294 682954 249914 711002
rect 249294 682718 249326 682954
rect 249562 682718 249646 682954
rect 249882 682718 249914 682954
rect 249294 682634 249914 682718
rect 249294 682398 249326 682634
rect 249562 682398 249646 682634
rect 249882 682398 249914 682634
rect 249294 646954 249914 682398
rect 249294 646718 249326 646954
rect 249562 646718 249646 646954
rect 249882 646718 249914 646954
rect 249294 646634 249914 646718
rect 249294 646398 249326 646634
rect 249562 646398 249646 646634
rect 249882 646398 249914 646634
rect 249294 610954 249914 646398
rect 249294 610718 249326 610954
rect 249562 610718 249646 610954
rect 249882 610718 249914 610954
rect 249294 610634 249914 610718
rect 249294 610398 249326 610634
rect 249562 610398 249646 610634
rect 249882 610398 249914 610634
rect 249294 574954 249914 610398
rect 249294 574718 249326 574954
rect 249562 574718 249646 574954
rect 249882 574718 249914 574954
rect 249294 574634 249914 574718
rect 249294 574398 249326 574634
rect 249562 574398 249646 574634
rect 249882 574398 249914 574634
rect 249294 538954 249914 574398
rect 249294 538718 249326 538954
rect 249562 538718 249646 538954
rect 249882 538718 249914 538954
rect 249294 538634 249914 538718
rect 249294 538398 249326 538634
rect 249562 538398 249646 538634
rect 249882 538398 249914 538634
rect 249294 502954 249914 538398
rect 249294 502718 249326 502954
rect 249562 502718 249646 502954
rect 249882 502718 249914 502954
rect 249294 502634 249914 502718
rect 249294 502398 249326 502634
rect 249562 502398 249646 502634
rect 249882 502398 249914 502634
rect 249294 466954 249914 502398
rect 249294 466718 249326 466954
rect 249562 466718 249646 466954
rect 249882 466718 249914 466954
rect 249294 466634 249914 466718
rect 249294 466398 249326 466634
rect 249562 466398 249646 466634
rect 249882 466398 249914 466634
rect 249294 430954 249914 466398
rect 249294 430718 249326 430954
rect 249562 430718 249646 430954
rect 249882 430718 249914 430954
rect 249294 430634 249914 430718
rect 249294 430398 249326 430634
rect 249562 430398 249646 430634
rect 249882 430398 249914 430634
rect 249294 394954 249914 430398
rect 249294 394718 249326 394954
rect 249562 394718 249646 394954
rect 249882 394718 249914 394954
rect 249294 394634 249914 394718
rect 249294 394398 249326 394634
rect 249562 394398 249646 394634
rect 249882 394398 249914 394634
rect 249294 358954 249914 394398
rect 249294 358718 249326 358954
rect 249562 358718 249646 358954
rect 249882 358718 249914 358954
rect 249294 358634 249914 358718
rect 249294 358398 249326 358634
rect 249562 358398 249646 358634
rect 249882 358398 249914 358634
rect 249294 322954 249914 358398
rect 249294 322718 249326 322954
rect 249562 322718 249646 322954
rect 249882 322718 249914 322954
rect 249294 322634 249914 322718
rect 249294 322398 249326 322634
rect 249562 322398 249646 322634
rect 249882 322398 249914 322634
rect 249294 286954 249914 322398
rect 249294 286718 249326 286954
rect 249562 286718 249646 286954
rect 249882 286718 249914 286954
rect 249294 286634 249914 286718
rect 249294 286398 249326 286634
rect 249562 286398 249646 286634
rect 249882 286398 249914 286634
rect 249294 250954 249914 286398
rect 249294 250718 249326 250954
rect 249562 250718 249646 250954
rect 249882 250718 249914 250954
rect 249294 250634 249914 250718
rect 249294 250398 249326 250634
rect 249562 250398 249646 250634
rect 249882 250398 249914 250634
rect 249294 214954 249914 250398
rect 249294 214718 249326 214954
rect 249562 214718 249646 214954
rect 249882 214718 249914 214954
rect 249294 214634 249914 214718
rect 249294 214398 249326 214634
rect 249562 214398 249646 214634
rect 249882 214398 249914 214634
rect 249294 178954 249914 214398
rect 249294 178718 249326 178954
rect 249562 178718 249646 178954
rect 249882 178718 249914 178954
rect 249294 178634 249914 178718
rect 249294 178398 249326 178634
rect 249562 178398 249646 178634
rect 249882 178398 249914 178634
rect 249294 142954 249914 178398
rect 249294 142718 249326 142954
rect 249562 142718 249646 142954
rect 249882 142718 249914 142954
rect 249294 142634 249914 142718
rect 249294 142398 249326 142634
rect 249562 142398 249646 142634
rect 249882 142398 249914 142634
rect 249294 106954 249914 142398
rect 249294 106718 249326 106954
rect 249562 106718 249646 106954
rect 249882 106718 249914 106954
rect 249294 106634 249914 106718
rect 249294 106398 249326 106634
rect 249562 106398 249646 106634
rect 249882 106398 249914 106634
rect 249294 70954 249914 106398
rect 249294 70718 249326 70954
rect 249562 70718 249646 70954
rect 249882 70718 249914 70954
rect 249294 70634 249914 70718
rect 249294 70398 249326 70634
rect 249562 70398 249646 70634
rect 249882 70398 249914 70634
rect 249294 34954 249914 70398
rect 249294 34718 249326 34954
rect 249562 34718 249646 34954
rect 249882 34718 249914 34954
rect 249294 34634 249914 34718
rect 249294 34398 249326 34634
rect 249562 34398 249646 34634
rect 249882 34398 249914 34634
rect 249294 -7066 249914 34398
rect 249294 -7302 249326 -7066
rect 249562 -7302 249646 -7066
rect 249882 -7302 249914 -7066
rect 249294 -7386 249914 -7302
rect 249294 -7622 249326 -7386
rect 249562 -7622 249646 -7386
rect 249882 -7622 249914 -7386
rect 249294 -7654 249914 -7622
rect 253794 704838 254414 711590
rect 253794 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 254414 704838
rect 253794 704518 254414 704602
rect 253794 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 254414 704518
rect 253794 687454 254414 704282
rect 253794 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 254414 687454
rect 253794 687134 254414 687218
rect 253794 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 254414 687134
rect 253794 651454 254414 686898
rect 253794 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 254414 651454
rect 253794 651134 254414 651218
rect 253794 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 254414 651134
rect 253794 615454 254414 650898
rect 253794 615218 253826 615454
rect 254062 615218 254146 615454
rect 254382 615218 254414 615454
rect 253794 615134 254414 615218
rect 253794 614898 253826 615134
rect 254062 614898 254146 615134
rect 254382 614898 254414 615134
rect 253794 579454 254414 614898
rect 253794 579218 253826 579454
rect 254062 579218 254146 579454
rect 254382 579218 254414 579454
rect 253794 579134 254414 579218
rect 253794 578898 253826 579134
rect 254062 578898 254146 579134
rect 254382 578898 254414 579134
rect 253794 543454 254414 578898
rect 253794 543218 253826 543454
rect 254062 543218 254146 543454
rect 254382 543218 254414 543454
rect 253794 543134 254414 543218
rect 253794 542898 253826 543134
rect 254062 542898 254146 543134
rect 254382 542898 254414 543134
rect 253794 507454 254414 542898
rect 253794 507218 253826 507454
rect 254062 507218 254146 507454
rect 254382 507218 254414 507454
rect 253794 507134 254414 507218
rect 253794 506898 253826 507134
rect 254062 506898 254146 507134
rect 254382 506898 254414 507134
rect 253794 471454 254414 506898
rect 253794 471218 253826 471454
rect 254062 471218 254146 471454
rect 254382 471218 254414 471454
rect 253794 471134 254414 471218
rect 253794 470898 253826 471134
rect 254062 470898 254146 471134
rect 254382 470898 254414 471134
rect 253794 435454 254414 470898
rect 253794 435218 253826 435454
rect 254062 435218 254146 435454
rect 254382 435218 254414 435454
rect 253794 435134 254414 435218
rect 253794 434898 253826 435134
rect 254062 434898 254146 435134
rect 254382 434898 254414 435134
rect 253794 399454 254414 434898
rect 253794 399218 253826 399454
rect 254062 399218 254146 399454
rect 254382 399218 254414 399454
rect 253794 399134 254414 399218
rect 253794 398898 253826 399134
rect 254062 398898 254146 399134
rect 254382 398898 254414 399134
rect 253794 363454 254414 398898
rect 253794 363218 253826 363454
rect 254062 363218 254146 363454
rect 254382 363218 254414 363454
rect 253794 363134 254414 363218
rect 253794 362898 253826 363134
rect 254062 362898 254146 363134
rect 254382 362898 254414 363134
rect 253794 327454 254414 362898
rect 253794 327218 253826 327454
rect 254062 327218 254146 327454
rect 254382 327218 254414 327454
rect 253794 327134 254414 327218
rect 253794 326898 253826 327134
rect 254062 326898 254146 327134
rect 254382 326898 254414 327134
rect 253794 291454 254414 326898
rect 253794 291218 253826 291454
rect 254062 291218 254146 291454
rect 254382 291218 254414 291454
rect 253794 291134 254414 291218
rect 253794 290898 253826 291134
rect 254062 290898 254146 291134
rect 254382 290898 254414 291134
rect 253794 255454 254414 290898
rect 253794 255218 253826 255454
rect 254062 255218 254146 255454
rect 254382 255218 254414 255454
rect 253794 255134 254414 255218
rect 253794 254898 253826 255134
rect 254062 254898 254146 255134
rect 254382 254898 254414 255134
rect 253794 219454 254414 254898
rect 253794 219218 253826 219454
rect 254062 219218 254146 219454
rect 254382 219218 254414 219454
rect 253794 219134 254414 219218
rect 253794 218898 253826 219134
rect 254062 218898 254146 219134
rect 254382 218898 254414 219134
rect 253794 183454 254414 218898
rect 253794 183218 253826 183454
rect 254062 183218 254146 183454
rect 254382 183218 254414 183454
rect 253794 183134 254414 183218
rect 253794 182898 253826 183134
rect 254062 182898 254146 183134
rect 254382 182898 254414 183134
rect 253794 147454 254414 182898
rect 253794 147218 253826 147454
rect 254062 147218 254146 147454
rect 254382 147218 254414 147454
rect 253794 147134 254414 147218
rect 253794 146898 253826 147134
rect 254062 146898 254146 147134
rect 254382 146898 254414 147134
rect 253794 111454 254414 146898
rect 253794 111218 253826 111454
rect 254062 111218 254146 111454
rect 254382 111218 254414 111454
rect 253794 111134 254414 111218
rect 253794 110898 253826 111134
rect 254062 110898 254146 111134
rect 254382 110898 254414 111134
rect 253794 75454 254414 110898
rect 253794 75218 253826 75454
rect 254062 75218 254146 75454
rect 254382 75218 254414 75454
rect 253794 75134 254414 75218
rect 253794 74898 253826 75134
rect 254062 74898 254146 75134
rect 254382 74898 254414 75134
rect 253794 39454 254414 74898
rect 253794 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 254414 39454
rect 253794 39134 254414 39218
rect 253794 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 254414 39134
rect 253794 3454 254414 38898
rect 253794 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 254414 3454
rect 253794 3134 254414 3218
rect 253794 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 254414 3134
rect 253794 -346 254414 2898
rect 253794 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 254414 -346
rect 253794 -666 254414 -582
rect 253794 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 254414 -666
rect 253794 -7654 254414 -902
rect 258294 705798 258914 711590
rect 258294 705562 258326 705798
rect 258562 705562 258646 705798
rect 258882 705562 258914 705798
rect 258294 705478 258914 705562
rect 258294 705242 258326 705478
rect 258562 705242 258646 705478
rect 258882 705242 258914 705478
rect 258294 691954 258914 705242
rect 258294 691718 258326 691954
rect 258562 691718 258646 691954
rect 258882 691718 258914 691954
rect 258294 691634 258914 691718
rect 258294 691398 258326 691634
rect 258562 691398 258646 691634
rect 258882 691398 258914 691634
rect 258294 655954 258914 691398
rect 258294 655718 258326 655954
rect 258562 655718 258646 655954
rect 258882 655718 258914 655954
rect 258294 655634 258914 655718
rect 258294 655398 258326 655634
rect 258562 655398 258646 655634
rect 258882 655398 258914 655634
rect 258294 619954 258914 655398
rect 258294 619718 258326 619954
rect 258562 619718 258646 619954
rect 258882 619718 258914 619954
rect 258294 619634 258914 619718
rect 258294 619398 258326 619634
rect 258562 619398 258646 619634
rect 258882 619398 258914 619634
rect 258294 583954 258914 619398
rect 258294 583718 258326 583954
rect 258562 583718 258646 583954
rect 258882 583718 258914 583954
rect 258294 583634 258914 583718
rect 258294 583398 258326 583634
rect 258562 583398 258646 583634
rect 258882 583398 258914 583634
rect 258294 547954 258914 583398
rect 258294 547718 258326 547954
rect 258562 547718 258646 547954
rect 258882 547718 258914 547954
rect 258294 547634 258914 547718
rect 258294 547398 258326 547634
rect 258562 547398 258646 547634
rect 258882 547398 258914 547634
rect 258294 511954 258914 547398
rect 258294 511718 258326 511954
rect 258562 511718 258646 511954
rect 258882 511718 258914 511954
rect 258294 511634 258914 511718
rect 258294 511398 258326 511634
rect 258562 511398 258646 511634
rect 258882 511398 258914 511634
rect 258294 475954 258914 511398
rect 258294 475718 258326 475954
rect 258562 475718 258646 475954
rect 258882 475718 258914 475954
rect 258294 475634 258914 475718
rect 258294 475398 258326 475634
rect 258562 475398 258646 475634
rect 258882 475398 258914 475634
rect 258294 439954 258914 475398
rect 258294 439718 258326 439954
rect 258562 439718 258646 439954
rect 258882 439718 258914 439954
rect 258294 439634 258914 439718
rect 258294 439398 258326 439634
rect 258562 439398 258646 439634
rect 258882 439398 258914 439634
rect 258294 403954 258914 439398
rect 258294 403718 258326 403954
rect 258562 403718 258646 403954
rect 258882 403718 258914 403954
rect 258294 403634 258914 403718
rect 258294 403398 258326 403634
rect 258562 403398 258646 403634
rect 258882 403398 258914 403634
rect 258294 367954 258914 403398
rect 258294 367718 258326 367954
rect 258562 367718 258646 367954
rect 258882 367718 258914 367954
rect 258294 367634 258914 367718
rect 258294 367398 258326 367634
rect 258562 367398 258646 367634
rect 258882 367398 258914 367634
rect 258294 331954 258914 367398
rect 258294 331718 258326 331954
rect 258562 331718 258646 331954
rect 258882 331718 258914 331954
rect 258294 331634 258914 331718
rect 258294 331398 258326 331634
rect 258562 331398 258646 331634
rect 258882 331398 258914 331634
rect 258294 295954 258914 331398
rect 258294 295718 258326 295954
rect 258562 295718 258646 295954
rect 258882 295718 258914 295954
rect 258294 295634 258914 295718
rect 258294 295398 258326 295634
rect 258562 295398 258646 295634
rect 258882 295398 258914 295634
rect 258294 259954 258914 295398
rect 258294 259718 258326 259954
rect 258562 259718 258646 259954
rect 258882 259718 258914 259954
rect 258294 259634 258914 259718
rect 258294 259398 258326 259634
rect 258562 259398 258646 259634
rect 258882 259398 258914 259634
rect 258294 223954 258914 259398
rect 258294 223718 258326 223954
rect 258562 223718 258646 223954
rect 258882 223718 258914 223954
rect 258294 223634 258914 223718
rect 258294 223398 258326 223634
rect 258562 223398 258646 223634
rect 258882 223398 258914 223634
rect 258294 187954 258914 223398
rect 258294 187718 258326 187954
rect 258562 187718 258646 187954
rect 258882 187718 258914 187954
rect 258294 187634 258914 187718
rect 258294 187398 258326 187634
rect 258562 187398 258646 187634
rect 258882 187398 258914 187634
rect 258294 151954 258914 187398
rect 258294 151718 258326 151954
rect 258562 151718 258646 151954
rect 258882 151718 258914 151954
rect 258294 151634 258914 151718
rect 258294 151398 258326 151634
rect 258562 151398 258646 151634
rect 258882 151398 258914 151634
rect 258294 115954 258914 151398
rect 258294 115718 258326 115954
rect 258562 115718 258646 115954
rect 258882 115718 258914 115954
rect 258294 115634 258914 115718
rect 258294 115398 258326 115634
rect 258562 115398 258646 115634
rect 258882 115398 258914 115634
rect 258294 79954 258914 115398
rect 258294 79718 258326 79954
rect 258562 79718 258646 79954
rect 258882 79718 258914 79954
rect 258294 79634 258914 79718
rect 258294 79398 258326 79634
rect 258562 79398 258646 79634
rect 258882 79398 258914 79634
rect 258294 43954 258914 79398
rect 258294 43718 258326 43954
rect 258562 43718 258646 43954
rect 258882 43718 258914 43954
rect 258294 43634 258914 43718
rect 258294 43398 258326 43634
rect 258562 43398 258646 43634
rect 258882 43398 258914 43634
rect 258294 7954 258914 43398
rect 258294 7718 258326 7954
rect 258562 7718 258646 7954
rect 258882 7718 258914 7954
rect 258294 7634 258914 7718
rect 258294 7398 258326 7634
rect 258562 7398 258646 7634
rect 258882 7398 258914 7634
rect 258294 -1306 258914 7398
rect 258294 -1542 258326 -1306
rect 258562 -1542 258646 -1306
rect 258882 -1542 258914 -1306
rect 258294 -1626 258914 -1542
rect 258294 -1862 258326 -1626
rect 258562 -1862 258646 -1626
rect 258882 -1862 258914 -1626
rect 258294 -7654 258914 -1862
rect 262794 706758 263414 711590
rect 262794 706522 262826 706758
rect 263062 706522 263146 706758
rect 263382 706522 263414 706758
rect 262794 706438 263414 706522
rect 262794 706202 262826 706438
rect 263062 706202 263146 706438
rect 263382 706202 263414 706438
rect 262794 696454 263414 706202
rect 262794 696218 262826 696454
rect 263062 696218 263146 696454
rect 263382 696218 263414 696454
rect 262794 696134 263414 696218
rect 262794 695898 262826 696134
rect 263062 695898 263146 696134
rect 263382 695898 263414 696134
rect 262794 660454 263414 695898
rect 262794 660218 262826 660454
rect 263062 660218 263146 660454
rect 263382 660218 263414 660454
rect 262794 660134 263414 660218
rect 262794 659898 262826 660134
rect 263062 659898 263146 660134
rect 263382 659898 263414 660134
rect 262794 624454 263414 659898
rect 262794 624218 262826 624454
rect 263062 624218 263146 624454
rect 263382 624218 263414 624454
rect 262794 624134 263414 624218
rect 262794 623898 262826 624134
rect 263062 623898 263146 624134
rect 263382 623898 263414 624134
rect 262794 588454 263414 623898
rect 262794 588218 262826 588454
rect 263062 588218 263146 588454
rect 263382 588218 263414 588454
rect 262794 588134 263414 588218
rect 262794 587898 262826 588134
rect 263062 587898 263146 588134
rect 263382 587898 263414 588134
rect 262794 552454 263414 587898
rect 262794 552218 262826 552454
rect 263062 552218 263146 552454
rect 263382 552218 263414 552454
rect 262794 552134 263414 552218
rect 262794 551898 262826 552134
rect 263062 551898 263146 552134
rect 263382 551898 263414 552134
rect 262794 516454 263414 551898
rect 262794 516218 262826 516454
rect 263062 516218 263146 516454
rect 263382 516218 263414 516454
rect 262794 516134 263414 516218
rect 262794 515898 262826 516134
rect 263062 515898 263146 516134
rect 263382 515898 263414 516134
rect 262794 480454 263414 515898
rect 262794 480218 262826 480454
rect 263062 480218 263146 480454
rect 263382 480218 263414 480454
rect 262794 480134 263414 480218
rect 262794 479898 262826 480134
rect 263062 479898 263146 480134
rect 263382 479898 263414 480134
rect 262794 444454 263414 479898
rect 262794 444218 262826 444454
rect 263062 444218 263146 444454
rect 263382 444218 263414 444454
rect 262794 444134 263414 444218
rect 262794 443898 262826 444134
rect 263062 443898 263146 444134
rect 263382 443898 263414 444134
rect 262794 408454 263414 443898
rect 262794 408218 262826 408454
rect 263062 408218 263146 408454
rect 263382 408218 263414 408454
rect 262794 408134 263414 408218
rect 262794 407898 262826 408134
rect 263062 407898 263146 408134
rect 263382 407898 263414 408134
rect 262794 372454 263414 407898
rect 262794 372218 262826 372454
rect 263062 372218 263146 372454
rect 263382 372218 263414 372454
rect 262794 372134 263414 372218
rect 262794 371898 262826 372134
rect 263062 371898 263146 372134
rect 263382 371898 263414 372134
rect 262794 336454 263414 371898
rect 262794 336218 262826 336454
rect 263062 336218 263146 336454
rect 263382 336218 263414 336454
rect 262794 336134 263414 336218
rect 262794 335898 262826 336134
rect 263062 335898 263146 336134
rect 263382 335898 263414 336134
rect 262794 300454 263414 335898
rect 262794 300218 262826 300454
rect 263062 300218 263146 300454
rect 263382 300218 263414 300454
rect 262794 300134 263414 300218
rect 262794 299898 262826 300134
rect 263062 299898 263146 300134
rect 263382 299898 263414 300134
rect 262794 264454 263414 299898
rect 262794 264218 262826 264454
rect 263062 264218 263146 264454
rect 263382 264218 263414 264454
rect 262794 264134 263414 264218
rect 262794 263898 262826 264134
rect 263062 263898 263146 264134
rect 263382 263898 263414 264134
rect 262794 228454 263414 263898
rect 262794 228218 262826 228454
rect 263062 228218 263146 228454
rect 263382 228218 263414 228454
rect 262794 228134 263414 228218
rect 262794 227898 262826 228134
rect 263062 227898 263146 228134
rect 263382 227898 263414 228134
rect 262794 192454 263414 227898
rect 262794 192218 262826 192454
rect 263062 192218 263146 192454
rect 263382 192218 263414 192454
rect 262794 192134 263414 192218
rect 262794 191898 262826 192134
rect 263062 191898 263146 192134
rect 263382 191898 263414 192134
rect 262794 156454 263414 191898
rect 262794 156218 262826 156454
rect 263062 156218 263146 156454
rect 263382 156218 263414 156454
rect 262794 156134 263414 156218
rect 262794 155898 262826 156134
rect 263062 155898 263146 156134
rect 263382 155898 263414 156134
rect 262794 120454 263414 155898
rect 262794 120218 262826 120454
rect 263062 120218 263146 120454
rect 263382 120218 263414 120454
rect 262794 120134 263414 120218
rect 262794 119898 262826 120134
rect 263062 119898 263146 120134
rect 263382 119898 263414 120134
rect 262794 84454 263414 119898
rect 262794 84218 262826 84454
rect 263062 84218 263146 84454
rect 263382 84218 263414 84454
rect 262794 84134 263414 84218
rect 262794 83898 262826 84134
rect 263062 83898 263146 84134
rect 263382 83898 263414 84134
rect 262794 48454 263414 83898
rect 262794 48218 262826 48454
rect 263062 48218 263146 48454
rect 263382 48218 263414 48454
rect 262794 48134 263414 48218
rect 262794 47898 262826 48134
rect 263062 47898 263146 48134
rect 263382 47898 263414 48134
rect 262794 12454 263414 47898
rect 262794 12218 262826 12454
rect 263062 12218 263146 12454
rect 263382 12218 263414 12454
rect 262794 12134 263414 12218
rect 262794 11898 262826 12134
rect 263062 11898 263146 12134
rect 263382 11898 263414 12134
rect 262794 -2266 263414 11898
rect 262794 -2502 262826 -2266
rect 263062 -2502 263146 -2266
rect 263382 -2502 263414 -2266
rect 262794 -2586 263414 -2502
rect 262794 -2822 262826 -2586
rect 263062 -2822 263146 -2586
rect 263382 -2822 263414 -2586
rect 262794 -7654 263414 -2822
rect 267294 707718 267914 711590
rect 267294 707482 267326 707718
rect 267562 707482 267646 707718
rect 267882 707482 267914 707718
rect 267294 707398 267914 707482
rect 267294 707162 267326 707398
rect 267562 707162 267646 707398
rect 267882 707162 267914 707398
rect 267294 700954 267914 707162
rect 267294 700718 267326 700954
rect 267562 700718 267646 700954
rect 267882 700718 267914 700954
rect 267294 700634 267914 700718
rect 267294 700398 267326 700634
rect 267562 700398 267646 700634
rect 267882 700398 267914 700634
rect 267294 664954 267914 700398
rect 267294 664718 267326 664954
rect 267562 664718 267646 664954
rect 267882 664718 267914 664954
rect 267294 664634 267914 664718
rect 267294 664398 267326 664634
rect 267562 664398 267646 664634
rect 267882 664398 267914 664634
rect 267294 628954 267914 664398
rect 267294 628718 267326 628954
rect 267562 628718 267646 628954
rect 267882 628718 267914 628954
rect 267294 628634 267914 628718
rect 267294 628398 267326 628634
rect 267562 628398 267646 628634
rect 267882 628398 267914 628634
rect 267294 592954 267914 628398
rect 267294 592718 267326 592954
rect 267562 592718 267646 592954
rect 267882 592718 267914 592954
rect 267294 592634 267914 592718
rect 267294 592398 267326 592634
rect 267562 592398 267646 592634
rect 267882 592398 267914 592634
rect 267294 556954 267914 592398
rect 267294 556718 267326 556954
rect 267562 556718 267646 556954
rect 267882 556718 267914 556954
rect 267294 556634 267914 556718
rect 267294 556398 267326 556634
rect 267562 556398 267646 556634
rect 267882 556398 267914 556634
rect 267294 520954 267914 556398
rect 267294 520718 267326 520954
rect 267562 520718 267646 520954
rect 267882 520718 267914 520954
rect 267294 520634 267914 520718
rect 267294 520398 267326 520634
rect 267562 520398 267646 520634
rect 267882 520398 267914 520634
rect 267294 484954 267914 520398
rect 267294 484718 267326 484954
rect 267562 484718 267646 484954
rect 267882 484718 267914 484954
rect 267294 484634 267914 484718
rect 267294 484398 267326 484634
rect 267562 484398 267646 484634
rect 267882 484398 267914 484634
rect 267294 448954 267914 484398
rect 267294 448718 267326 448954
rect 267562 448718 267646 448954
rect 267882 448718 267914 448954
rect 267294 448634 267914 448718
rect 267294 448398 267326 448634
rect 267562 448398 267646 448634
rect 267882 448398 267914 448634
rect 267294 412954 267914 448398
rect 267294 412718 267326 412954
rect 267562 412718 267646 412954
rect 267882 412718 267914 412954
rect 267294 412634 267914 412718
rect 267294 412398 267326 412634
rect 267562 412398 267646 412634
rect 267882 412398 267914 412634
rect 267294 376954 267914 412398
rect 267294 376718 267326 376954
rect 267562 376718 267646 376954
rect 267882 376718 267914 376954
rect 267294 376634 267914 376718
rect 267294 376398 267326 376634
rect 267562 376398 267646 376634
rect 267882 376398 267914 376634
rect 267294 340954 267914 376398
rect 267294 340718 267326 340954
rect 267562 340718 267646 340954
rect 267882 340718 267914 340954
rect 267294 340634 267914 340718
rect 267294 340398 267326 340634
rect 267562 340398 267646 340634
rect 267882 340398 267914 340634
rect 267294 304954 267914 340398
rect 267294 304718 267326 304954
rect 267562 304718 267646 304954
rect 267882 304718 267914 304954
rect 267294 304634 267914 304718
rect 267294 304398 267326 304634
rect 267562 304398 267646 304634
rect 267882 304398 267914 304634
rect 267294 268954 267914 304398
rect 267294 268718 267326 268954
rect 267562 268718 267646 268954
rect 267882 268718 267914 268954
rect 267294 268634 267914 268718
rect 267294 268398 267326 268634
rect 267562 268398 267646 268634
rect 267882 268398 267914 268634
rect 267294 232954 267914 268398
rect 267294 232718 267326 232954
rect 267562 232718 267646 232954
rect 267882 232718 267914 232954
rect 267294 232634 267914 232718
rect 267294 232398 267326 232634
rect 267562 232398 267646 232634
rect 267882 232398 267914 232634
rect 267294 196954 267914 232398
rect 267294 196718 267326 196954
rect 267562 196718 267646 196954
rect 267882 196718 267914 196954
rect 267294 196634 267914 196718
rect 267294 196398 267326 196634
rect 267562 196398 267646 196634
rect 267882 196398 267914 196634
rect 267294 160954 267914 196398
rect 267294 160718 267326 160954
rect 267562 160718 267646 160954
rect 267882 160718 267914 160954
rect 267294 160634 267914 160718
rect 267294 160398 267326 160634
rect 267562 160398 267646 160634
rect 267882 160398 267914 160634
rect 267294 124954 267914 160398
rect 267294 124718 267326 124954
rect 267562 124718 267646 124954
rect 267882 124718 267914 124954
rect 267294 124634 267914 124718
rect 267294 124398 267326 124634
rect 267562 124398 267646 124634
rect 267882 124398 267914 124634
rect 267294 88954 267914 124398
rect 267294 88718 267326 88954
rect 267562 88718 267646 88954
rect 267882 88718 267914 88954
rect 267294 88634 267914 88718
rect 267294 88398 267326 88634
rect 267562 88398 267646 88634
rect 267882 88398 267914 88634
rect 267294 52954 267914 88398
rect 267294 52718 267326 52954
rect 267562 52718 267646 52954
rect 267882 52718 267914 52954
rect 267294 52634 267914 52718
rect 267294 52398 267326 52634
rect 267562 52398 267646 52634
rect 267882 52398 267914 52634
rect 267294 16954 267914 52398
rect 267294 16718 267326 16954
rect 267562 16718 267646 16954
rect 267882 16718 267914 16954
rect 267294 16634 267914 16718
rect 267294 16398 267326 16634
rect 267562 16398 267646 16634
rect 267882 16398 267914 16634
rect 267294 -3226 267914 16398
rect 267294 -3462 267326 -3226
rect 267562 -3462 267646 -3226
rect 267882 -3462 267914 -3226
rect 267294 -3546 267914 -3462
rect 267294 -3782 267326 -3546
rect 267562 -3782 267646 -3546
rect 267882 -3782 267914 -3546
rect 267294 -7654 267914 -3782
rect 271794 708678 272414 711590
rect 271794 708442 271826 708678
rect 272062 708442 272146 708678
rect 272382 708442 272414 708678
rect 271794 708358 272414 708442
rect 271794 708122 271826 708358
rect 272062 708122 272146 708358
rect 272382 708122 272414 708358
rect 271794 669454 272414 708122
rect 271794 669218 271826 669454
rect 272062 669218 272146 669454
rect 272382 669218 272414 669454
rect 271794 669134 272414 669218
rect 271794 668898 271826 669134
rect 272062 668898 272146 669134
rect 272382 668898 272414 669134
rect 271794 633454 272414 668898
rect 271794 633218 271826 633454
rect 272062 633218 272146 633454
rect 272382 633218 272414 633454
rect 271794 633134 272414 633218
rect 271794 632898 271826 633134
rect 272062 632898 272146 633134
rect 272382 632898 272414 633134
rect 271794 597454 272414 632898
rect 271794 597218 271826 597454
rect 272062 597218 272146 597454
rect 272382 597218 272414 597454
rect 271794 597134 272414 597218
rect 271794 596898 271826 597134
rect 272062 596898 272146 597134
rect 272382 596898 272414 597134
rect 271794 561454 272414 596898
rect 271794 561218 271826 561454
rect 272062 561218 272146 561454
rect 272382 561218 272414 561454
rect 271794 561134 272414 561218
rect 271794 560898 271826 561134
rect 272062 560898 272146 561134
rect 272382 560898 272414 561134
rect 271794 525454 272414 560898
rect 271794 525218 271826 525454
rect 272062 525218 272146 525454
rect 272382 525218 272414 525454
rect 271794 525134 272414 525218
rect 271794 524898 271826 525134
rect 272062 524898 272146 525134
rect 272382 524898 272414 525134
rect 271794 489454 272414 524898
rect 271794 489218 271826 489454
rect 272062 489218 272146 489454
rect 272382 489218 272414 489454
rect 271794 489134 272414 489218
rect 271794 488898 271826 489134
rect 272062 488898 272146 489134
rect 272382 488898 272414 489134
rect 271794 453454 272414 488898
rect 271794 453218 271826 453454
rect 272062 453218 272146 453454
rect 272382 453218 272414 453454
rect 271794 453134 272414 453218
rect 271794 452898 271826 453134
rect 272062 452898 272146 453134
rect 272382 452898 272414 453134
rect 271794 417454 272414 452898
rect 271794 417218 271826 417454
rect 272062 417218 272146 417454
rect 272382 417218 272414 417454
rect 271794 417134 272414 417218
rect 271794 416898 271826 417134
rect 272062 416898 272146 417134
rect 272382 416898 272414 417134
rect 271794 381454 272414 416898
rect 271794 381218 271826 381454
rect 272062 381218 272146 381454
rect 272382 381218 272414 381454
rect 271794 381134 272414 381218
rect 271794 380898 271826 381134
rect 272062 380898 272146 381134
rect 272382 380898 272414 381134
rect 271794 345454 272414 380898
rect 271794 345218 271826 345454
rect 272062 345218 272146 345454
rect 272382 345218 272414 345454
rect 271794 345134 272414 345218
rect 271794 344898 271826 345134
rect 272062 344898 272146 345134
rect 272382 344898 272414 345134
rect 271794 309454 272414 344898
rect 271794 309218 271826 309454
rect 272062 309218 272146 309454
rect 272382 309218 272414 309454
rect 271794 309134 272414 309218
rect 271794 308898 271826 309134
rect 272062 308898 272146 309134
rect 272382 308898 272414 309134
rect 271794 273454 272414 308898
rect 271794 273218 271826 273454
rect 272062 273218 272146 273454
rect 272382 273218 272414 273454
rect 271794 273134 272414 273218
rect 271794 272898 271826 273134
rect 272062 272898 272146 273134
rect 272382 272898 272414 273134
rect 271794 237454 272414 272898
rect 271794 237218 271826 237454
rect 272062 237218 272146 237454
rect 272382 237218 272414 237454
rect 271794 237134 272414 237218
rect 271794 236898 271826 237134
rect 272062 236898 272146 237134
rect 272382 236898 272414 237134
rect 271794 201454 272414 236898
rect 271794 201218 271826 201454
rect 272062 201218 272146 201454
rect 272382 201218 272414 201454
rect 271794 201134 272414 201218
rect 271794 200898 271826 201134
rect 272062 200898 272146 201134
rect 272382 200898 272414 201134
rect 271794 165454 272414 200898
rect 271794 165218 271826 165454
rect 272062 165218 272146 165454
rect 272382 165218 272414 165454
rect 271794 165134 272414 165218
rect 271794 164898 271826 165134
rect 272062 164898 272146 165134
rect 272382 164898 272414 165134
rect 271794 129454 272414 164898
rect 271794 129218 271826 129454
rect 272062 129218 272146 129454
rect 272382 129218 272414 129454
rect 271794 129134 272414 129218
rect 271794 128898 271826 129134
rect 272062 128898 272146 129134
rect 272382 128898 272414 129134
rect 271794 93454 272414 128898
rect 271794 93218 271826 93454
rect 272062 93218 272146 93454
rect 272382 93218 272414 93454
rect 271794 93134 272414 93218
rect 271794 92898 271826 93134
rect 272062 92898 272146 93134
rect 272382 92898 272414 93134
rect 271794 57454 272414 92898
rect 271794 57218 271826 57454
rect 272062 57218 272146 57454
rect 272382 57218 272414 57454
rect 271794 57134 272414 57218
rect 271794 56898 271826 57134
rect 272062 56898 272146 57134
rect 272382 56898 272414 57134
rect 271794 21454 272414 56898
rect 271794 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 272414 21454
rect 271794 21134 272414 21218
rect 271794 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 272414 21134
rect 271794 -4186 272414 20898
rect 271794 -4422 271826 -4186
rect 272062 -4422 272146 -4186
rect 272382 -4422 272414 -4186
rect 271794 -4506 272414 -4422
rect 271794 -4742 271826 -4506
rect 272062 -4742 272146 -4506
rect 272382 -4742 272414 -4506
rect 271794 -7654 272414 -4742
rect 276294 709638 276914 711590
rect 276294 709402 276326 709638
rect 276562 709402 276646 709638
rect 276882 709402 276914 709638
rect 276294 709318 276914 709402
rect 276294 709082 276326 709318
rect 276562 709082 276646 709318
rect 276882 709082 276914 709318
rect 276294 673954 276914 709082
rect 276294 673718 276326 673954
rect 276562 673718 276646 673954
rect 276882 673718 276914 673954
rect 276294 673634 276914 673718
rect 276294 673398 276326 673634
rect 276562 673398 276646 673634
rect 276882 673398 276914 673634
rect 276294 637954 276914 673398
rect 276294 637718 276326 637954
rect 276562 637718 276646 637954
rect 276882 637718 276914 637954
rect 276294 637634 276914 637718
rect 276294 637398 276326 637634
rect 276562 637398 276646 637634
rect 276882 637398 276914 637634
rect 276294 601954 276914 637398
rect 276294 601718 276326 601954
rect 276562 601718 276646 601954
rect 276882 601718 276914 601954
rect 276294 601634 276914 601718
rect 276294 601398 276326 601634
rect 276562 601398 276646 601634
rect 276882 601398 276914 601634
rect 276294 565954 276914 601398
rect 276294 565718 276326 565954
rect 276562 565718 276646 565954
rect 276882 565718 276914 565954
rect 276294 565634 276914 565718
rect 276294 565398 276326 565634
rect 276562 565398 276646 565634
rect 276882 565398 276914 565634
rect 276294 529954 276914 565398
rect 276294 529718 276326 529954
rect 276562 529718 276646 529954
rect 276882 529718 276914 529954
rect 276294 529634 276914 529718
rect 276294 529398 276326 529634
rect 276562 529398 276646 529634
rect 276882 529398 276914 529634
rect 276294 493954 276914 529398
rect 276294 493718 276326 493954
rect 276562 493718 276646 493954
rect 276882 493718 276914 493954
rect 276294 493634 276914 493718
rect 276294 493398 276326 493634
rect 276562 493398 276646 493634
rect 276882 493398 276914 493634
rect 276294 457954 276914 493398
rect 276294 457718 276326 457954
rect 276562 457718 276646 457954
rect 276882 457718 276914 457954
rect 276294 457634 276914 457718
rect 276294 457398 276326 457634
rect 276562 457398 276646 457634
rect 276882 457398 276914 457634
rect 276294 421954 276914 457398
rect 276294 421718 276326 421954
rect 276562 421718 276646 421954
rect 276882 421718 276914 421954
rect 276294 421634 276914 421718
rect 276294 421398 276326 421634
rect 276562 421398 276646 421634
rect 276882 421398 276914 421634
rect 276294 385954 276914 421398
rect 276294 385718 276326 385954
rect 276562 385718 276646 385954
rect 276882 385718 276914 385954
rect 276294 385634 276914 385718
rect 276294 385398 276326 385634
rect 276562 385398 276646 385634
rect 276882 385398 276914 385634
rect 276294 349954 276914 385398
rect 276294 349718 276326 349954
rect 276562 349718 276646 349954
rect 276882 349718 276914 349954
rect 276294 349634 276914 349718
rect 276294 349398 276326 349634
rect 276562 349398 276646 349634
rect 276882 349398 276914 349634
rect 276294 313954 276914 349398
rect 276294 313718 276326 313954
rect 276562 313718 276646 313954
rect 276882 313718 276914 313954
rect 276294 313634 276914 313718
rect 276294 313398 276326 313634
rect 276562 313398 276646 313634
rect 276882 313398 276914 313634
rect 276294 277954 276914 313398
rect 276294 277718 276326 277954
rect 276562 277718 276646 277954
rect 276882 277718 276914 277954
rect 276294 277634 276914 277718
rect 276294 277398 276326 277634
rect 276562 277398 276646 277634
rect 276882 277398 276914 277634
rect 276294 241954 276914 277398
rect 276294 241718 276326 241954
rect 276562 241718 276646 241954
rect 276882 241718 276914 241954
rect 276294 241634 276914 241718
rect 276294 241398 276326 241634
rect 276562 241398 276646 241634
rect 276882 241398 276914 241634
rect 276294 205954 276914 241398
rect 276294 205718 276326 205954
rect 276562 205718 276646 205954
rect 276882 205718 276914 205954
rect 276294 205634 276914 205718
rect 276294 205398 276326 205634
rect 276562 205398 276646 205634
rect 276882 205398 276914 205634
rect 276294 169954 276914 205398
rect 276294 169718 276326 169954
rect 276562 169718 276646 169954
rect 276882 169718 276914 169954
rect 276294 169634 276914 169718
rect 276294 169398 276326 169634
rect 276562 169398 276646 169634
rect 276882 169398 276914 169634
rect 276294 133954 276914 169398
rect 276294 133718 276326 133954
rect 276562 133718 276646 133954
rect 276882 133718 276914 133954
rect 276294 133634 276914 133718
rect 276294 133398 276326 133634
rect 276562 133398 276646 133634
rect 276882 133398 276914 133634
rect 276294 97954 276914 133398
rect 276294 97718 276326 97954
rect 276562 97718 276646 97954
rect 276882 97718 276914 97954
rect 276294 97634 276914 97718
rect 276294 97398 276326 97634
rect 276562 97398 276646 97634
rect 276882 97398 276914 97634
rect 276294 61954 276914 97398
rect 276294 61718 276326 61954
rect 276562 61718 276646 61954
rect 276882 61718 276914 61954
rect 276294 61634 276914 61718
rect 276294 61398 276326 61634
rect 276562 61398 276646 61634
rect 276882 61398 276914 61634
rect 276294 25954 276914 61398
rect 276294 25718 276326 25954
rect 276562 25718 276646 25954
rect 276882 25718 276914 25954
rect 276294 25634 276914 25718
rect 276294 25398 276326 25634
rect 276562 25398 276646 25634
rect 276882 25398 276914 25634
rect 276294 -5146 276914 25398
rect 276294 -5382 276326 -5146
rect 276562 -5382 276646 -5146
rect 276882 -5382 276914 -5146
rect 276294 -5466 276914 -5382
rect 276294 -5702 276326 -5466
rect 276562 -5702 276646 -5466
rect 276882 -5702 276914 -5466
rect 276294 -7654 276914 -5702
rect 280794 710598 281414 711590
rect 280794 710362 280826 710598
rect 281062 710362 281146 710598
rect 281382 710362 281414 710598
rect 280794 710278 281414 710362
rect 280794 710042 280826 710278
rect 281062 710042 281146 710278
rect 281382 710042 281414 710278
rect 280794 678454 281414 710042
rect 280794 678218 280826 678454
rect 281062 678218 281146 678454
rect 281382 678218 281414 678454
rect 280794 678134 281414 678218
rect 280794 677898 280826 678134
rect 281062 677898 281146 678134
rect 281382 677898 281414 678134
rect 280794 642454 281414 677898
rect 280794 642218 280826 642454
rect 281062 642218 281146 642454
rect 281382 642218 281414 642454
rect 280794 642134 281414 642218
rect 280794 641898 280826 642134
rect 281062 641898 281146 642134
rect 281382 641898 281414 642134
rect 280794 606454 281414 641898
rect 280794 606218 280826 606454
rect 281062 606218 281146 606454
rect 281382 606218 281414 606454
rect 280794 606134 281414 606218
rect 280794 605898 280826 606134
rect 281062 605898 281146 606134
rect 281382 605898 281414 606134
rect 280794 570454 281414 605898
rect 280794 570218 280826 570454
rect 281062 570218 281146 570454
rect 281382 570218 281414 570454
rect 280794 570134 281414 570218
rect 280794 569898 280826 570134
rect 281062 569898 281146 570134
rect 281382 569898 281414 570134
rect 280794 534454 281414 569898
rect 280794 534218 280826 534454
rect 281062 534218 281146 534454
rect 281382 534218 281414 534454
rect 280794 534134 281414 534218
rect 280794 533898 280826 534134
rect 281062 533898 281146 534134
rect 281382 533898 281414 534134
rect 280794 498454 281414 533898
rect 280794 498218 280826 498454
rect 281062 498218 281146 498454
rect 281382 498218 281414 498454
rect 280794 498134 281414 498218
rect 280794 497898 280826 498134
rect 281062 497898 281146 498134
rect 281382 497898 281414 498134
rect 280794 462454 281414 497898
rect 280794 462218 280826 462454
rect 281062 462218 281146 462454
rect 281382 462218 281414 462454
rect 280794 462134 281414 462218
rect 280794 461898 280826 462134
rect 281062 461898 281146 462134
rect 281382 461898 281414 462134
rect 280794 426454 281414 461898
rect 280794 426218 280826 426454
rect 281062 426218 281146 426454
rect 281382 426218 281414 426454
rect 280794 426134 281414 426218
rect 280794 425898 280826 426134
rect 281062 425898 281146 426134
rect 281382 425898 281414 426134
rect 280794 390454 281414 425898
rect 280794 390218 280826 390454
rect 281062 390218 281146 390454
rect 281382 390218 281414 390454
rect 280794 390134 281414 390218
rect 280794 389898 280826 390134
rect 281062 389898 281146 390134
rect 281382 389898 281414 390134
rect 280794 354454 281414 389898
rect 280794 354218 280826 354454
rect 281062 354218 281146 354454
rect 281382 354218 281414 354454
rect 280794 354134 281414 354218
rect 280794 353898 280826 354134
rect 281062 353898 281146 354134
rect 281382 353898 281414 354134
rect 280794 318454 281414 353898
rect 280794 318218 280826 318454
rect 281062 318218 281146 318454
rect 281382 318218 281414 318454
rect 280794 318134 281414 318218
rect 280794 317898 280826 318134
rect 281062 317898 281146 318134
rect 281382 317898 281414 318134
rect 280794 282454 281414 317898
rect 280794 282218 280826 282454
rect 281062 282218 281146 282454
rect 281382 282218 281414 282454
rect 280794 282134 281414 282218
rect 280794 281898 280826 282134
rect 281062 281898 281146 282134
rect 281382 281898 281414 282134
rect 280794 246454 281414 281898
rect 280794 246218 280826 246454
rect 281062 246218 281146 246454
rect 281382 246218 281414 246454
rect 280794 246134 281414 246218
rect 280794 245898 280826 246134
rect 281062 245898 281146 246134
rect 281382 245898 281414 246134
rect 280794 210454 281414 245898
rect 280794 210218 280826 210454
rect 281062 210218 281146 210454
rect 281382 210218 281414 210454
rect 280794 210134 281414 210218
rect 280794 209898 280826 210134
rect 281062 209898 281146 210134
rect 281382 209898 281414 210134
rect 280794 174454 281414 209898
rect 280794 174218 280826 174454
rect 281062 174218 281146 174454
rect 281382 174218 281414 174454
rect 280794 174134 281414 174218
rect 280794 173898 280826 174134
rect 281062 173898 281146 174134
rect 281382 173898 281414 174134
rect 280794 138454 281414 173898
rect 280794 138218 280826 138454
rect 281062 138218 281146 138454
rect 281382 138218 281414 138454
rect 280794 138134 281414 138218
rect 280794 137898 280826 138134
rect 281062 137898 281146 138134
rect 281382 137898 281414 138134
rect 280794 102454 281414 137898
rect 280794 102218 280826 102454
rect 281062 102218 281146 102454
rect 281382 102218 281414 102454
rect 280794 102134 281414 102218
rect 280794 101898 280826 102134
rect 281062 101898 281146 102134
rect 281382 101898 281414 102134
rect 280794 66454 281414 101898
rect 280794 66218 280826 66454
rect 281062 66218 281146 66454
rect 281382 66218 281414 66454
rect 280794 66134 281414 66218
rect 280794 65898 280826 66134
rect 281062 65898 281146 66134
rect 281382 65898 281414 66134
rect 280794 30454 281414 65898
rect 280794 30218 280826 30454
rect 281062 30218 281146 30454
rect 281382 30218 281414 30454
rect 280794 30134 281414 30218
rect 280794 29898 280826 30134
rect 281062 29898 281146 30134
rect 281382 29898 281414 30134
rect 280794 -6106 281414 29898
rect 280794 -6342 280826 -6106
rect 281062 -6342 281146 -6106
rect 281382 -6342 281414 -6106
rect 280794 -6426 281414 -6342
rect 280794 -6662 280826 -6426
rect 281062 -6662 281146 -6426
rect 281382 -6662 281414 -6426
rect 280794 -7654 281414 -6662
rect 285294 711558 285914 711590
rect 285294 711322 285326 711558
rect 285562 711322 285646 711558
rect 285882 711322 285914 711558
rect 285294 711238 285914 711322
rect 285294 711002 285326 711238
rect 285562 711002 285646 711238
rect 285882 711002 285914 711238
rect 285294 682954 285914 711002
rect 285294 682718 285326 682954
rect 285562 682718 285646 682954
rect 285882 682718 285914 682954
rect 285294 682634 285914 682718
rect 285294 682398 285326 682634
rect 285562 682398 285646 682634
rect 285882 682398 285914 682634
rect 285294 646954 285914 682398
rect 285294 646718 285326 646954
rect 285562 646718 285646 646954
rect 285882 646718 285914 646954
rect 285294 646634 285914 646718
rect 285294 646398 285326 646634
rect 285562 646398 285646 646634
rect 285882 646398 285914 646634
rect 285294 610954 285914 646398
rect 285294 610718 285326 610954
rect 285562 610718 285646 610954
rect 285882 610718 285914 610954
rect 285294 610634 285914 610718
rect 285294 610398 285326 610634
rect 285562 610398 285646 610634
rect 285882 610398 285914 610634
rect 285294 574954 285914 610398
rect 285294 574718 285326 574954
rect 285562 574718 285646 574954
rect 285882 574718 285914 574954
rect 285294 574634 285914 574718
rect 285294 574398 285326 574634
rect 285562 574398 285646 574634
rect 285882 574398 285914 574634
rect 285294 538954 285914 574398
rect 285294 538718 285326 538954
rect 285562 538718 285646 538954
rect 285882 538718 285914 538954
rect 285294 538634 285914 538718
rect 285294 538398 285326 538634
rect 285562 538398 285646 538634
rect 285882 538398 285914 538634
rect 285294 502954 285914 538398
rect 285294 502718 285326 502954
rect 285562 502718 285646 502954
rect 285882 502718 285914 502954
rect 285294 502634 285914 502718
rect 285294 502398 285326 502634
rect 285562 502398 285646 502634
rect 285882 502398 285914 502634
rect 285294 466954 285914 502398
rect 285294 466718 285326 466954
rect 285562 466718 285646 466954
rect 285882 466718 285914 466954
rect 285294 466634 285914 466718
rect 285294 466398 285326 466634
rect 285562 466398 285646 466634
rect 285882 466398 285914 466634
rect 285294 430954 285914 466398
rect 285294 430718 285326 430954
rect 285562 430718 285646 430954
rect 285882 430718 285914 430954
rect 285294 430634 285914 430718
rect 285294 430398 285326 430634
rect 285562 430398 285646 430634
rect 285882 430398 285914 430634
rect 285294 394954 285914 430398
rect 285294 394718 285326 394954
rect 285562 394718 285646 394954
rect 285882 394718 285914 394954
rect 285294 394634 285914 394718
rect 285294 394398 285326 394634
rect 285562 394398 285646 394634
rect 285882 394398 285914 394634
rect 285294 358954 285914 394398
rect 285294 358718 285326 358954
rect 285562 358718 285646 358954
rect 285882 358718 285914 358954
rect 285294 358634 285914 358718
rect 285294 358398 285326 358634
rect 285562 358398 285646 358634
rect 285882 358398 285914 358634
rect 285294 322954 285914 358398
rect 285294 322718 285326 322954
rect 285562 322718 285646 322954
rect 285882 322718 285914 322954
rect 285294 322634 285914 322718
rect 285294 322398 285326 322634
rect 285562 322398 285646 322634
rect 285882 322398 285914 322634
rect 285294 286954 285914 322398
rect 285294 286718 285326 286954
rect 285562 286718 285646 286954
rect 285882 286718 285914 286954
rect 285294 286634 285914 286718
rect 285294 286398 285326 286634
rect 285562 286398 285646 286634
rect 285882 286398 285914 286634
rect 285294 250954 285914 286398
rect 285294 250718 285326 250954
rect 285562 250718 285646 250954
rect 285882 250718 285914 250954
rect 285294 250634 285914 250718
rect 285294 250398 285326 250634
rect 285562 250398 285646 250634
rect 285882 250398 285914 250634
rect 285294 214954 285914 250398
rect 285294 214718 285326 214954
rect 285562 214718 285646 214954
rect 285882 214718 285914 214954
rect 285294 214634 285914 214718
rect 285294 214398 285326 214634
rect 285562 214398 285646 214634
rect 285882 214398 285914 214634
rect 285294 178954 285914 214398
rect 285294 178718 285326 178954
rect 285562 178718 285646 178954
rect 285882 178718 285914 178954
rect 285294 178634 285914 178718
rect 285294 178398 285326 178634
rect 285562 178398 285646 178634
rect 285882 178398 285914 178634
rect 285294 142954 285914 178398
rect 285294 142718 285326 142954
rect 285562 142718 285646 142954
rect 285882 142718 285914 142954
rect 285294 142634 285914 142718
rect 285294 142398 285326 142634
rect 285562 142398 285646 142634
rect 285882 142398 285914 142634
rect 285294 106954 285914 142398
rect 285294 106718 285326 106954
rect 285562 106718 285646 106954
rect 285882 106718 285914 106954
rect 285294 106634 285914 106718
rect 285294 106398 285326 106634
rect 285562 106398 285646 106634
rect 285882 106398 285914 106634
rect 285294 70954 285914 106398
rect 285294 70718 285326 70954
rect 285562 70718 285646 70954
rect 285882 70718 285914 70954
rect 285294 70634 285914 70718
rect 285294 70398 285326 70634
rect 285562 70398 285646 70634
rect 285882 70398 285914 70634
rect 285294 34954 285914 70398
rect 285294 34718 285326 34954
rect 285562 34718 285646 34954
rect 285882 34718 285914 34954
rect 285294 34634 285914 34718
rect 285294 34398 285326 34634
rect 285562 34398 285646 34634
rect 285882 34398 285914 34634
rect 285294 -7066 285914 34398
rect 285294 -7302 285326 -7066
rect 285562 -7302 285646 -7066
rect 285882 -7302 285914 -7066
rect 285294 -7386 285914 -7302
rect 285294 -7622 285326 -7386
rect 285562 -7622 285646 -7386
rect 285882 -7622 285914 -7386
rect 285294 -7654 285914 -7622
rect 289794 704838 290414 711590
rect 289794 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 290414 704838
rect 289794 704518 290414 704602
rect 289794 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 290414 704518
rect 289794 687454 290414 704282
rect 289794 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 290414 687454
rect 289794 687134 290414 687218
rect 289794 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 290414 687134
rect 289794 651454 290414 686898
rect 289794 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 290414 651454
rect 289794 651134 290414 651218
rect 289794 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 290414 651134
rect 289794 615454 290414 650898
rect 289794 615218 289826 615454
rect 290062 615218 290146 615454
rect 290382 615218 290414 615454
rect 289794 615134 290414 615218
rect 289794 614898 289826 615134
rect 290062 614898 290146 615134
rect 290382 614898 290414 615134
rect 289794 579454 290414 614898
rect 289794 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 290414 579454
rect 289794 579134 290414 579218
rect 289794 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 290414 579134
rect 289794 543454 290414 578898
rect 289794 543218 289826 543454
rect 290062 543218 290146 543454
rect 290382 543218 290414 543454
rect 289794 543134 290414 543218
rect 289794 542898 289826 543134
rect 290062 542898 290146 543134
rect 290382 542898 290414 543134
rect 289794 507454 290414 542898
rect 289794 507218 289826 507454
rect 290062 507218 290146 507454
rect 290382 507218 290414 507454
rect 289794 507134 290414 507218
rect 289794 506898 289826 507134
rect 290062 506898 290146 507134
rect 290382 506898 290414 507134
rect 289794 471454 290414 506898
rect 289794 471218 289826 471454
rect 290062 471218 290146 471454
rect 290382 471218 290414 471454
rect 289794 471134 290414 471218
rect 289794 470898 289826 471134
rect 290062 470898 290146 471134
rect 290382 470898 290414 471134
rect 289794 435454 290414 470898
rect 289794 435218 289826 435454
rect 290062 435218 290146 435454
rect 290382 435218 290414 435454
rect 289794 435134 290414 435218
rect 289794 434898 289826 435134
rect 290062 434898 290146 435134
rect 290382 434898 290414 435134
rect 289794 399454 290414 434898
rect 289794 399218 289826 399454
rect 290062 399218 290146 399454
rect 290382 399218 290414 399454
rect 289794 399134 290414 399218
rect 289794 398898 289826 399134
rect 290062 398898 290146 399134
rect 290382 398898 290414 399134
rect 289794 363454 290414 398898
rect 289794 363218 289826 363454
rect 290062 363218 290146 363454
rect 290382 363218 290414 363454
rect 289794 363134 290414 363218
rect 289794 362898 289826 363134
rect 290062 362898 290146 363134
rect 290382 362898 290414 363134
rect 289794 327454 290414 362898
rect 289794 327218 289826 327454
rect 290062 327218 290146 327454
rect 290382 327218 290414 327454
rect 289794 327134 290414 327218
rect 289794 326898 289826 327134
rect 290062 326898 290146 327134
rect 290382 326898 290414 327134
rect 289794 291454 290414 326898
rect 289794 291218 289826 291454
rect 290062 291218 290146 291454
rect 290382 291218 290414 291454
rect 289794 291134 290414 291218
rect 289794 290898 289826 291134
rect 290062 290898 290146 291134
rect 290382 290898 290414 291134
rect 289794 255454 290414 290898
rect 289794 255218 289826 255454
rect 290062 255218 290146 255454
rect 290382 255218 290414 255454
rect 289794 255134 290414 255218
rect 289794 254898 289826 255134
rect 290062 254898 290146 255134
rect 290382 254898 290414 255134
rect 289794 219454 290414 254898
rect 289794 219218 289826 219454
rect 290062 219218 290146 219454
rect 290382 219218 290414 219454
rect 289794 219134 290414 219218
rect 289794 218898 289826 219134
rect 290062 218898 290146 219134
rect 290382 218898 290414 219134
rect 289794 183454 290414 218898
rect 289794 183218 289826 183454
rect 290062 183218 290146 183454
rect 290382 183218 290414 183454
rect 289794 183134 290414 183218
rect 289794 182898 289826 183134
rect 290062 182898 290146 183134
rect 290382 182898 290414 183134
rect 289794 147454 290414 182898
rect 289794 147218 289826 147454
rect 290062 147218 290146 147454
rect 290382 147218 290414 147454
rect 289794 147134 290414 147218
rect 289794 146898 289826 147134
rect 290062 146898 290146 147134
rect 290382 146898 290414 147134
rect 289794 111454 290414 146898
rect 289794 111218 289826 111454
rect 290062 111218 290146 111454
rect 290382 111218 290414 111454
rect 289794 111134 290414 111218
rect 289794 110898 289826 111134
rect 290062 110898 290146 111134
rect 290382 110898 290414 111134
rect 289794 75454 290414 110898
rect 289794 75218 289826 75454
rect 290062 75218 290146 75454
rect 290382 75218 290414 75454
rect 289794 75134 290414 75218
rect 289794 74898 289826 75134
rect 290062 74898 290146 75134
rect 290382 74898 290414 75134
rect 289794 39454 290414 74898
rect 289794 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 290414 39454
rect 289794 39134 290414 39218
rect 289794 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 290414 39134
rect 289794 3454 290414 38898
rect 289794 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 290414 3454
rect 289794 3134 290414 3218
rect 289794 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 290414 3134
rect 289794 -346 290414 2898
rect 289794 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 290414 -346
rect 289794 -666 290414 -582
rect 289794 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 290414 -666
rect 289794 -7654 290414 -902
rect 294294 705798 294914 711590
rect 294294 705562 294326 705798
rect 294562 705562 294646 705798
rect 294882 705562 294914 705798
rect 294294 705478 294914 705562
rect 294294 705242 294326 705478
rect 294562 705242 294646 705478
rect 294882 705242 294914 705478
rect 294294 691954 294914 705242
rect 294294 691718 294326 691954
rect 294562 691718 294646 691954
rect 294882 691718 294914 691954
rect 294294 691634 294914 691718
rect 294294 691398 294326 691634
rect 294562 691398 294646 691634
rect 294882 691398 294914 691634
rect 294294 655954 294914 691398
rect 294294 655718 294326 655954
rect 294562 655718 294646 655954
rect 294882 655718 294914 655954
rect 294294 655634 294914 655718
rect 294294 655398 294326 655634
rect 294562 655398 294646 655634
rect 294882 655398 294914 655634
rect 294294 619954 294914 655398
rect 294294 619718 294326 619954
rect 294562 619718 294646 619954
rect 294882 619718 294914 619954
rect 294294 619634 294914 619718
rect 294294 619398 294326 619634
rect 294562 619398 294646 619634
rect 294882 619398 294914 619634
rect 294294 583954 294914 619398
rect 294294 583718 294326 583954
rect 294562 583718 294646 583954
rect 294882 583718 294914 583954
rect 294294 583634 294914 583718
rect 294294 583398 294326 583634
rect 294562 583398 294646 583634
rect 294882 583398 294914 583634
rect 294294 547954 294914 583398
rect 294294 547718 294326 547954
rect 294562 547718 294646 547954
rect 294882 547718 294914 547954
rect 294294 547634 294914 547718
rect 294294 547398 294326 547634
rect 294562 547398 294646 547634
rect 294882 547398 294914 547634
rect 294294 511954 294914 547398
rect 294294 511718 294326 511954
rect 294562 511718 294646 511954
rect 294882 511718 294914 511954
rect 294294 511634 294914 511718
rect 294294 511398 294326 511634
rect 294562 511398 294646 511634
rect 294882 511398 294914 511634
rect 294294 475954 294914 511398
rect 294294 475718 294326 475954
rect 294562 475718 294646 475954
rect 294882 475718 294914 475954
rect 294294 475634 294914 475718
rect 294294 475398 294326 475634
rect 294562 475398 294646 475634
rect 294882 475398 294914 475634
rect 294294 439954 294914 475398
rect 294294 439718 294326 439954
rect 294562 439718 294646 439954
rect 294882 439718 294914 439954
rect 294294 439634 294914 439718
rect 294294 439398 294326 439634
rect 294562 439398 294646 439634
rect 294882 439398 294914 439634
rect 294294 403954 294914 439398
rect 294294 403718 294326 403954
rect 294562 403718 294646 403954
rect 294882 403718 294914 403954
rect 294294 403634 294914 403718
rect 294294 403398 294326 403634
rect 294562 403398 294646 403634
rect 294882 403398 294914 403634
rect 294294 367954 294914 403398
rect 294294 367718 294326 367954
rect 294562 367718 294646 367954
rect 294882 367718 294914 367954
rect 294294 367634 294914 367718
rect 294294 367398 294326 367634
rect 294562 367398 294646 367634
rect 294882 367398 294914 367634
rect 294294 331954 294914 367398
rect 294294 331718 294326 331954
rect 294562 331718 294646 331954
rect 294882 331718 294914 331954
rect 294294 331634 294914 331718
rect 294294 331398 294326 331634
rect 294562 331398 294646 331634
rect 294882 331398 294914 331634
rect 294294 295954 294914 331398
rect 294294 295718 294326 295954
rect 294562 295718 294646 295954
rect 294882 295718 294914 295954
rect 294294 295634 294914 295718
rect 294294 295398 294326 295634
rect 294562 295398 294646 295634
rect 294882 295398 294914 295634
rect 294294 259954 294914 295398
rect 294294 259718 294326 259954
rect 294562 259718 294646 259954
rect 294882 259718 294914 259954
rect 294294 259634 294914 259718
rect 294294 259398 294326 259634
rect 294562 259398 294646 259634
rect 294882 259398 294914 259634
rect 294294 223954 294914 259398
rect 294294 223718 294326 223954
rect 294562 223718 294646 223954
rect 294882 223718 294914 223954
rect 294294 223634 294914 223718
rect 294294 223398 294326 223634
rect 294562 223398 294646 223634
rect 294882 223398 294914 223634
rect 294294 187954 294914 223398
rect 294294 187718 294326 187954
rect 294562 187718 294646 187954
rect 294882 187718 294914 187954
rect 294294 187634 294914 187718
rect 294294 187398 294326 187634
rect 294562 187398 294646 187634
rect 294882 187398 294914 187634
rect 294294 151954 294914 187398
rect 294294 151718 294326 151954
rect 294562 151718 294646 151954
rect 294882 151718 294914 151954
rect 294294 151634 294914 151718
rect 294294 151398 294326 151634
rect 294562 151398 294646 151634
rect 294882 151398 294914 151634
rect 294294 115954 294914 151398
rect 294294 115718 294326 115954
rect 294562 115718 294646 115954
rect 294882 115718 294914 115954
rect 294294 115634 294914 115718
rect 294294 115398 294326 115634
rect 294562 115398 294646 115634
rect 294882 115398 294914 115634
rect 294294 79954 294914 115398
rect 294294 79718 294326 79954
rect 294562 79718 294646 79954
rect 294882 79718 294914 79954
rect 294294 79634 294914 79718
rect 294294 79398 294326 79634
rect 294562 79398 294646 79634
rect 294882 79398 294914 79634
rect 294294 43954 294914 79398
rect 294294 43718 294326 43954
rect 294562 43718 294646 43954
rect 294882 43718 294914 43954
rect 294294 43634 294914 43718
rect 294294 43398 294326 43634
rect 294562 43398 294646 43634
rect 294882 43398 294914 43634
rect 294294 7954 294914 43398
rect 294294 7718 294326 7954
rect 294562 7718 294646 7954
rect 294882 7718 294914 7954
rect 294294 7634 294914 7718
rect 294294 7398 294326 7634
rect 294562 7398 294646 7634
rect 294882 7398 294914 7634
rect 294294 -1306 294914 7398
rect 294294 -1542 294326 -1306
rect 294562 -1542 294646 -1306
rect 294882 -1542 294914 -1306
rect 294294 -1626 294914 -1542
rect 294294 -1862 294326 -1626
rect 294562 -1862 294646 -1626
rect 294882 -1862 294914 -1626
rect 294294 -7654 294914 -1862
rect 298794 706758 299414 711590
rect 298794 706522 298826 706758
rect 299062 706522 299146 706758
rect 299382 706522 299414 706758
rect 298794 706438 299414 706522
rect 298794 706202 298826 706438
rect 299062 706202 299146 706438
rect 299382 706202 299414 706438
rect 298794 696454 299414 706202
rect 298794 696218 298826 696454
rect 299062 696218 299146 696454
rect 299382 696218 299414 696454
rect 298794 696134 299414 696218
rect 298794 695898 298826 696134
rect 299062 695898 299146 696134
rect 299382 695898 299414 696134
rect 298794 660454 299414 695898
rect 298794 660218 298826 660454
rect 299062 660218 299146 660454
rect 299382 660218 299414 660454
rect 298794 660134 299414 660218
rect 298794 659898 298826 660134
rect 299062 659898 299146 660134
rect 299382 659898 299414 660134
rect 298794 624454 299414 659898
rect 298794 624218 298826 624454
rect 299062 624218 299146 624454
rect 299382 624218 299414 624454
rect 298794 624134 299414 624218
rect 298794 623898 298826 624134
rect 299062 623898 299146 624134
rect 299382 623898 299414 624134
rect 298794 588454 299414 623898
rect 298794 588218 298826 588454
rect 299062 588218 299146 588454
rect 299382 588218 299414 588454
rect 298794 588134 299414 588218
rect 298794 587898 298826 588134
rect 299062 587898 299146 588134
rect 299382 587898 299414 588134
rect 298794 552454 299414 587898
rect 298794 552218 298826 552454
rect 299062 552218 299146 552454
rect 299382 552218 299414 552454
rect 298794 552134 299414 552218
rect 298794 551898 298826 552134
rect 299062 551898 299146 552134
rect 299382 551898 299414 552134
rect 298794 516454 299414 551898
rect 298794 516218 298826 516454
rect 299062 516218 299146 516454
rect 299382 516218 299414 516454
rect 298794 516134 299414 516218
rect 298794 515898 298826 516134
rect 299062 515898 299146 516134
rect 299382 515898 299414 516134
rect 298794 480454 299414 515898
rect 298794 480218 298826 480454
rect 299062 480218 299146 480454
rect 299382 480218 299414 480454
rect 298794 480134 299414 480218
rect 298794 479898 298826 480134
rect 299062 479898 299146 480134
rect 299382 479898 299414 480134
rect 298794 444454 299414 479898
rect 298794 444218 298826 444454
rect 299062 444218 299146 444454
rect 299382 444218 299414 444454
rect 298794 444134 299414 444218
rect 298794 443898 298826 444134
rect 299062 443898 299146 444134
rect 299382 443898 299414 444134
rect 298794 408454 299414 443898
rect 298794 408218 298826 408454
rect 299062 408218 299146 408454
rect 299382 408218 299414 408454
rect 298794 408134 299414 408218
rect 298794 407898 298826 408134
rect 299062 407898 299146 408134
rect 299382 407898 299414 408134
rect 298794 372454 299414 407898
rect 298794 372218 298826 372454
rect 299062 372218 299146 372454
rect 299382 372218 299414 372454
rect 298794 372134 299414 372218
rect 298794 371898 298826 372134
rect 299062 371898 299146 372134
rect 299382 371898 299414 372134
rect 298794 336454 299414 371898
rect 298794 336218 298826 336454
rect 299062 336218 299146 336454
rect 299382 336218 299414 336454
rect 298794 336134 299414 336218
rect 298794 335898 298826 336134
rect 299062 335898 299146 336134
rect 299382 335898 299414 336134
rect 298794 300454 299414 335898
rect 298794 300218 298826 300454
rect 299062 300218 299146 300454
rect 299382 300218 299414 300454
rect 298794 300134 299414 300218
rect 298794 299898 298826 300134
rect 299062 299898 299146 300134
rect 299382 299898 299414 300134
rect 298794 264454 299414 299898
rect 298794 264218 298826 264454
rect 299062 264218 299146 264454
rect 299382 264218 299414 264454
rect 298794 264134 299414 264218
rect 298794 263898 298826 264134
rect 299062 263898 299146 264134
rect 299382 263898 299414 264134
rect 298794 228454 299414 263898
rect 298794 228218 298826 228454
rect 299062 228218 299146 228454
rect 299382 228218 299414 228454
rect 298794 228134 299414 228218
rect 298794 227898 298826 228134
rect 299062 227898 299146 228134
rect 299382 227898 299414 228134
rect 298794 192454 299414 227898
rect 298794 192218 298826 192454
rect 299062 192218 299146 192454
rect 299382 192218 299414 192454
rect 298794 192134 299414 192218
rect 298794 191898 298826 192134
rect 299062 191898 299146 192134
rect 299382 191898 299414 192134
rect 298794 156454 299414 191898
rect 298794 156218 298826 156454
rect 299062 156218 299146 156454
rect 299382 156218 299414 156454
rect 298794 156134 299414 156218
rect 298794 155898 298826 156134
rect 299062 155898 299146 156134
rect 299382 155898 299414 156134
rect 298794 120454 299414 155898
rect 298794 120218 298826 120454
rect 299062 120218 299146 120454
rect 299382 120218 299414 120454
rect 298794 120134 299414 120218
rect 298794 119898 298826 120134
rect 299062 119898 299146 120134
rect 299382 119898 299414 120134
rect 298794 84454 299414 119898
rect 298794 84218 298826 84454
rect 299062 84218 299146 84454
rect 299382 84218 299414 84454
rect 298794 84134 299414 84218
rect 298794 83898 298826 84134
rect 299062 83898 299146 84134
rect 299382 83898 299414 84134
rect 298794 48454 299414 83898
rect 298794 48218 298826 48454
rect 299062 48218 299146 48454
rect 299382 48218 299414 48454
rect 298794 48134 299414 48218
rect 298794 47898 298826 48134
rect 299062 47898 299146 48134
rect 299382 47898 299414 48134
rect 298794 12454 299414 47898
rect 298794 12218 298826 12454
rect 299062 12218 299146 12454
rect 299382 12218 299414 12454
rect 298794 12134 299414 12218
rect 298794 11898 298826 12134
rect 299062 11898 299146 12134
rect 299382 11898 299414 12134
rect 298794 -2266 299414 11898
rect 298794 -2502 298826 -2266
rect 299062 -2502 299146 -2266
rect 299382 -2502 299414 -2266
rect 298794 -2586 299414 -2502
rect 298794 -2822 298826 -2586
rect 299062 -2822 299146 -2586
rect 299382 -2822 299414 -2586
rect 298794 -7654 299414 -2822
rect 303294 707718 303914 711590
rect 303294 707482 303326 707718
rect 303562 707482 303646 707718
rect 303882 707482 303914 707718
rect 303294 707398 303914 707482
rect 303294 707162 303326 707398
rect 303562 707162 303646 707398
rect 303882 707162 303914 707398
rect 303294 700954 303914 707162
rect 303294 700718 303326 700954
rect 303562 700718 303646 700954
rect 303882 700718 303914 700954
rect 303294 700634 303914 700718
rect 303294 700398 303326 700634
rect 303562 700398 303646 700634
rect 303882 700398 303914 700634
rect 303294 664954 303914 700398
rect 303294 664718 303326 664954
rect 303562 664718 303646 664954
rect 303882 664718 303914 664954
rect 303294 664634 303914 664718
rect 303294 664398 303326 664634
rect 303562 664398 303646 664634
rect 303882 664398 303914 664634
rect 303294 628954 303914 664398
rect 303294 628718 303326 628954
rect 303562 628718 303646 628954
rect 303882 628718 303914 628954
rect 303294 628634 303914 628718
rect 303294 628398 303326 628634
rect 303562 628398 303646 628634
rect 303882 628398 303914 628634
rect 303294 592954 303914 628398
rect 303294 592718 303326 592954
rect 303562 592718 303646 592954
rect 303882 592718 303914 592954
rect 303294 592634 303914 592718
rect 303294 592398 303326 592634
rect 303562 592398 303646 592634
rect 303882 592398 303914 592634
rect 303294 556954 303914 592398
rect 303294 556718 303326 556954
rect 303562 556718 303646 556954
rect 303882 556718 303914 556954
rect 303294 556634 303914 556718
rect 303294 556398 303326 556634
rect 303562 556398 303646 556634
rect 303882 556398 303914 556634
rect 303294 520954 303914 556398
rect 303294 520718 303326 520954
rect 303562 520718 303646 520954
rect 303882 520718 303914 520954
rect 303294 520634 303914 520718
rect 303294 520398 303326 520634
rect 303562 520398 303646 520634
rect 303882 520398 303914 520634
rect 303294 484954 303914 520398
rect 303294 484718 303326 484954
rect 303562 484718 303646 484954
rect 303882 484718 303914 484954
rect 303294 484634 303914 484718
rect 303294 484398 303326 484634
rect 303562 484398 303646 484634
rect 303882 484398 303914 484634
rect 303294 448954 303914 484398
rect 303294 448718 303326 448954
rect 303562 448718 303646 448954
rect 303882 448718 303914 448954
rect 303294 448634 303914 448718
rect 303294 448398 303326 448634
rect 303562 448398 303646 448634
rect 303882 448398 303914 448634
rect 303294 412954 303914 448398
rect 303294 412718 303326 412954
rect 303562 412718 303646 412954
rect 303882 412718 303914 412954
rect 303294 412634 303914 412718
rect 303294 412398 303326 412634
rect 303562 412398 303646 412634
rect 303882 412398 303914 412634
rect 303294 376954 303914 412398
rect 303294 376718 303326 376954
rect 303562 376718 303646 376954
rect 303882 376718 303914 376954
rect 303294 376634 303914 376718
rect 303294 376398 303326 376634
rect 303562 376398 303646 376634
rect 303882 376398 303914 376634
rect 303294 340954 303914 376398
rect 303294 340718 303326 340954
rect 303562 340718 303646 340954
rect 303882 340718 303914 340954
rect 303294 340634 303914 340718
rect 303294 340398 303326 340634
rect 303562 340398 303646 340634
rect 303882 340398 303914 340634
rect 303294 304954 303914 340398
rect 303294 304718 303326 304954
rect 303562 304718 303646 304954
rect 303882 304718 303914 304954
rect 303294 304634 303914 304718
rect 303294 304398 303326 304634
rect 303562 304398 303646 304634
rect 303882 304398 303914 304634
rect 303294 268954 303914 304398
rect 303294 268718 303326 268954
rect 303562 268718 303646 268954
rect 303882 268718 303914 268954
rect 303294 268634 303914 268718
rect 303294 268398 303326 268634
rect 303562 268398 303646 268634
rect 303882 268398 303914 268634
rect 303294 232954 303914 268398
rect 303294 232718 303326 232954
rect 303562 232718 303646 232954
rect 303882 232718 303914 232954
rect 303294 232634 303914 232718
rect 303294 232398 303326 232634
rect 303562 232398 303646 232634
rect 303882 232398 303914 232634
rect 303294 196954 303914 232398
rect 303294 196718 303326 196954
rect 303562 196718 303646 196954
rect 303882 196718 303914 196954
rect 303294 196634 303914 196718
rect 303294 196398 303326 196634
rect 303562 196398 303646 196634
rect 303882 196398 303914 196634
rect 303294 160954 303914 196398
rect 303294 160718 303326 160954
rect 303562 160718 303646 160954
rect 303882 160718 303914 160954
rect 303294 160634 303914 160718
rect 303294 160398 303326 160634
rect 303562 160398 303646 160634
rect 303882 160398 303914 160634
rect 303294 124954 303914 160398
rect 303294 124718 303326 124954
rect 303562 124718 303646 124954
rect 303882 124718 303914 124954
rect 303294 124634 303914 124718
rect 303294 124398 303326 124634
rect 303562 124398 303646 124634
rect 303882 124398 303914 124634
rect 303294 88954 303914 124398
rect 303294 88718 303326 88954
rect 303562 88718 303646 88954
rect 303882 88718 303914 88954
rect 303294 88634 303914 88718
rect 303294 88398 303326 88634
rect 303562 88398 303646 88634
rect 303882 88398 303914 88634
rect 303294 52954 303914 88398
rect 303294 52718 303326 52954
rect 303562 52718 303646 52954
rect 303882 52718 303914 52954
rect 303294 52634 303914 52718
rect 303294 52398 303326 52634
rect 303562 52398 303646 52634
rect 303882 52398 303914 52634
rect 303294 16954 303914 52398
rect 303294 16718 303326 16954
rect 303562 16718 303646 16954
rect 303882 16718 303914 16954
rect 303294 16634 303914 16718
rect 303294 16398 303326 16634
rect 303562 16398 303646 16634
rect 303882 16398 303914 16634
rect 303294 -3226 303914 16398
rect 303294 -3462 303326 -3226
rect 303562 -3462 303646 -3226
rect 303882 -3462 303914 -3226
rect 303294 -3546 303914 -3462
rect 303294 -3782 303326 -3546
rect 303562 -3782 303646 -3546
rect 303882 -3782 303914 -3546
rect 303294 -7654 303914 -3782
rect 307794 708678 308414 711590
rect 307794 708442 307826 708678
rect 308062 708442 308146 708678
rect 308382 708442 308414 708678
rect 307794 708358 308414 708442
rect 307794 708122 307826 708358
rect 308062 708122 308146 708358
rect 308382 708122 308414 708358
rect 307794 669454 308414 708122
rect 307794 669218 307826 669454
rect 308062 669218 308146 669454
rect 308382 669218 308414 669454
rect 307794 669134 308414 669218
rect 307794 668898 307826 669134
rect 308062 668898 308146 669134
rect 308382 668898 308414 669134
rect 307794 633454 308414 668898
rect 307794 633218 307826 633454
rect 308062 633218 308146 633454
rect 308382 633218 308414 633454
rect 307794 633134 308414 633218
rect 307794 632898 307826 633134
rect 308062 632898 308146 633134
rect 308382 632898 308414 633134
rect 307794 597454 308414 632898
rect 307794 597218 307826 597454
rect 308062 597218 308146 597454
rect 308382 597218 308414 597454
rect 307794 597134 308414 597218
rect 307794 596898 307826 597134
rect 308062 596898 308146 597134
rect 308382 596898 308414 597134
rect 307794 561454 308414 596898
rect 307794 561218 307826 561454
rect 308062 561218 308146 561454
rect 308382 561218 308414 561454
rect 307794 561134 308414 561218
rect 307794 560898 307826 561134
rect 308062 560898 308146 561134
rect 308382 560898 308414 561134
rect 307794 525454 308414 560898
rect 307794 525218 307826 525454
rect 308062 525218 308146 525454
rect 308382 525218 308414 525454
rect 307794 525134 308414 525218
rect 307794 524898 307826 525134
rect 308062 524898 308146 525134
rect 308382 524898 308414 525134
rect 307794 489454 308414 524898
rect 307794 489218 307826 489454
rect 308062 489218 308146 489454
rect 308382 489218 308414 489454
rect 307794 489134 308414 489218
rect 307794 488898 307826 489134
rect 308062 488898 308146 489134
rect 308382 488898 308414 489134
rect 307794 453454 308414 488898
rect 307794 453218 307826 453454
rect 308062 453218 308146 453454
rect 308382 453218 308414 453454
rect 307794 453134 308414 453218
rect 307794 452898 307826 453134
rect 308062 452898 308146 453134
rect 308382 452898 308414 453134
rect 307794 417454 308414 452898
rect 307794 417218 307826 417454
rect 308062 417218 308146 417454
rect 308382 417218 308414 417454
rect 307794 417134 308414 417218
rect 307794 416898 307826 417134
rect 308062 416898 308146 417134
rect 308382 416898 308414 417134
rect 307794 381454 308414 416898
rect 307794 381218 307826 381454
rect 308062 381218 308146 381454
rect 308382 381218 308414 381454
rect 307794 381134 308414 381218
rect 307794 380898 307826 381134
rect 308062 380898 308146 381134
rect 308382 380898 308414 381134
rect 307794 345454 308414 380898
rect 307794 345218 307826 345454
rect 308062 345218 308146 345454
rect 308382 345218 308414 345454
rect 307794 345134 308414 345218
rect 307794 344898 307826 345134
rect 308062 344898 308146 345134
rect 308382 344898 308414 345134
rect 307794 309454 308414 344898
rect 307794 309218 307826 309454
rect 308062 309218 308146 309454
rect 308382 309218 308414 309454
rect 307794 309134 308414 309218
rect 307794 308898 307826 309134
rect 308062 308898 308146 309134
rect 308382 308898 308414 309134
rect 307794 273454 308414 308898
rect 307794 273218 307826 273454
rect 308062 273218 308146 273454
rect 308382 273218 308414 273454
rect 307794 273134 308414 273218
rect 307794 272898 307826 273134
rect 308062 272898 308146 273134
rect 308382 272898 308414 273134
rect 307794 237454 308414 272898
rect 307794 237218 307826 237454
rect 308062 237218 308146 237454
rect 308382 237218 308414 237454
rect 307794 237134 308414 237218
rect 307794 236898 307826 237134
rect 308062 236898 308146 237134
rect 308382 236898 308414 237134
rect 307794 201454 308414 236898
rect 307794 201218 307826 201454
rect 308062 201218 308146 201454
rect 308382 201218 308414 201454
rect 307794 201134 308414 201218
rect 307794 200898 307826 201134
rect 308062 200898 308146 201134
rect 308382 200898 308414 201134
rect 307794 165454 308414 200898
rect 307794 165218 307826 165454
rect 308062 165218 308146 165454
rect 308382 165218 308414 165454
rect 307794 165134 308414 165218
rect 307794 164898 307826 165134
rect 308062 164898 308146 165134
rect 308382 164898 308414 165134
rect 307794 129454 308414 164898
rect 307794 129218 307826 129454
rect 308062 129218 308146 129454
rect 308382 129218 308414 129454
rect 307794 129134 308414 129218
rect 307794 128898 307826 129134
rect 308062 128898 308146 129134
rect 308382 128898 308414 129134
rect 307794 93454 308414 128898
rect 307794 93218 307826 93454
rect 308062 93218 308146 93454
rect 308382 93218 308414 93454
rect 307794 93134 308414 93218
rect 307794 92898 307826 93134
rect 308062 92898 308146 93134
rect 308382 92898 308414 93134
rect 307794 57454 308414 92898
rect 307794 57218 307826 57454
rect 308062 57218 308146 57454
rect 308382 57218 308414 57454
rect 307794 57134 308414 57218
rect 307794 56898 307826 57134
rect 308062 56898 308146 57134
rect 308382 56898 308414 57134
rect 307794 21454 308414 56898
rect 307794 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 308414 21454
rect 307794 21134 308414 21218
rect 307794 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 308414 21134
rect 307794 -4186 308414 20898
rect 307794 -4422 307826 -4186
rect 308062 -4422 308146 -4186
rect 308382 -4422 308414 -4186
rect 307794 -4506 308414 -4422
rect 307794 -4742 307826 -4506
rect 308062 -4742 308146 -4506
rect 308382 -4742 308414 -4506
rect 307794 -7654 308414 -4742
rect 312294 709638 312914 711590
rect 312294 709402 312326 709638
rect 312562 709402 312646 709638
rect 312882 709402 312914 709638
rect 312294 709318 312914 709402
rect 312294 709082 312326 709318
rect 312562 709082 312646 709318
rect 312882 709082 312914 709318
rect 312294 673954 312914 709082
rect 312294 673718 312326 673954
rect 312562 673718 312646 673954
rect 312882 673718 312914 673954
rect 312294 673634 312914 673718
rect 312294 673398 312326 673634
rect 312562 673398 312646 673634
rect 312882 673398 312914 673634
rect 312294 637954 312914 673398
rect 312294 637718 312326 637954
rect 312562 637718 312646 637954
rect 312882 637718 312914 637954
rect 312294 637634 312914 637718
rect 312294 637398 312326 637634
rect 312562 637398 312646 637634
rect 312882 637398 312914 637634
rect 312294 601954 312914 637398
rect 312294 601718 312326 601954
rect 312562 601718 312646 601954
rect 312882 601718 312914 601954
rect 312294 601634 312914 601718
rect 312294 601398 312326 601634
rect 312562 601398 312646 601634
rect 312882 601398 312914 601634
rect 312294 565954 312914 601398
rect 312294 565718 312326 565954
rect 312562 565718 312646 565954
rect 312882 565718 312914 565954
rect 312294 565634 312914 565718
rect 312294 565398 312326 565634
rect 312562 565398 312646 565634
rect 312882 565398 312914 565634
rect 312294 529954 312914 565398
rect 312294 529718 312326 529954
rect 312562 529718 312646 529954
rect 312882 529718 312914 529954
rect 312294 529634 312914 529718
rect 312294 529398 312326 529634
rect 312562 529398 312646 529634
rect 312882 529398 312914 529634
rect 312294 493954 312914 529398
rect 312294 493718 312326 493954
rect 312562 493718 312646 493954
rect 312882 493718 312914 493954
rect 312294 493634 312914 493718
rect 312294 493398 312326 493634
rect 312562 493398 312646 493634
rect 312882 493398 312914 493634
rect 312294 457954 312914 493398
rect 312294 457718 312326 457954
rect 312562 457718 312646 457954
rect 312882 457718 312914 457954
rect 312294 457634 312914 457718
rect 312294 457398 312326 457634
rect 312562 457398 312646 457634
rect 312882 457398 312914 457634
rect 312294 421954 312914 457398
rect 312294 421718 312326 421954
rect 312562 421718 312646 421954
rect 312882 421718 312914 421954
rect 312294 421634 312914 421718
rect 312294 421398 312326 421634
rect 312562 421398 312646 421634
rect 312882 421398 312914 421634
rect 312294 385954 312914 421398
rect 312294 385718 312326 385954
rect 312562 385718 312646 385954
rect 312882 385718 312914 385954
rect 312294 385634 312914 385718
rect 312294 385398 312326 385634
rect 312562 385398 312646 385634
rect 312882 385398 312914 385634
rect 312294 349954 312914 385398
rect 312294 349718 312326 349954
rect 312562 349718 312646 349954
rect 312882 349718 312914 349954
rect 312294 349634 312914 349718
rect 312294 349398 312326 349634
rect 312562 349398 312646 349634
rect 312882 349398 312914 349634
rect 312294 313954 312914 349398
rect 312294 313718 312326 313954
rect 312562 313718 312646 313954
rect 312882 313718 312914 313954
rect 312294 313634 312914 313718
rect 312294 313398 312326 313634
rect 312562 313398 312646 313634
rect 312882 313398 312914 313634
rect 312294 277954 312914 313398
rect 312294 277718 312326 277954
rect 312562 277718 312646 277954
rect 312882 277718 312914 277954
rect 312294 277634 312914 277718
rect 312294 277398 312326 277634
rect 312562 277398 312646 277634
rect 312882 277398 312914 277634
rect 312294 241954 312914 277398
rect 312294 241718 312326 241954
rect 312562 241718 312646 241954
rect 312882 241718 312914 241954
rect 312294 241634 312914 241718
rect 312294 241398 312326 241634
rect 312562 241398 312646 241634
rect 312882 241398 312914 241634
rect 312294 205954 312914 241398
rect 312294 205718 312326 205954
rect 312562 205718 312646 205954
rect 312882 205718 312914 205954
rect 312294 205634 312914 205718
rect 312294 205398 312326 205634
rect 312562 205398 312646 205634
rect 312882 205398 312914 205634
rect 312294 169954 312914 205398
rect 312294 169718 312326 169954
rect 312562 169718 312646 169954
rect 312882 169718 312914 169954
rect 312294 169634 312914 169718
rect 312294 169398 312326 169634
rect 312562 169398 312646 169634
rect 312882 169398 312914 169634
rect 312294 133954 312914 169398
rect 312294 133718 312326 133954
rect 312562 133718 312646 133954
rect 312882 133718 312914 133954
rect 312294 133634 312914 133718
rect 312294 133398 312326 133634
rect 312562 133398 312646 133634
rect 312882 133398 312914 133634
rect 312294 97954 312914 133398
rect 312294 97718 312326 97954
rect 312562 97718 312646 97954
rect 312882 97718 312914 97954
rect 312294 97634 312914 97718
rect 312294 97398 312326 97634
rect 312562 97398 312646 97634
rect 312882 97398 312914 97634
rect 312294 61954 312914 97398
rect 312294 61718 312326 61954
rect 312562 61718 312646 61954
rect 312882 61718 312914 61954
rect 312294 61634 312914 61718
rect 312294 61398 312326 61634
rect 312562 61398 312646 61634
rect 312882 61398 312914 61634
rect 312294 25954 312914 61398
rect 312294 25718 312326 25954
rect 312562 25718 312646 25954
rect 312882 25718 312914 25954
rect 312294 25634 312914 25718
rect 312294 25398 312326 25634
rect 312562 25398 312646 25634
rect 312882 25398 312914 25634
rect 312294 -5146 312914 25398
rect 312294 -5382 312326 -5146
rect 312562 -5382 312646 -5146
rect 312882 -5382 312914 -5146
rect 312294 -5466 312914 -5382
rect 312294 -5702 312326 -5466
rect 312562 -5702 312646 -5466
rect 312882 -5702 312914 -5466
rect 312294 -7654 312914 -5702
rect 316794 710598 317414 711590
rect 316794 710362 316826 710598
rect 317062 710362 317146 710598
rect 317382 710362 317414 710598
rect 316794 710278 317414 710362
rect 316794 710042 316826 710278
rect 317062 710042 317146 710278
rect 317382 710042 317414 710278
rect 316794 678454 317414 710042
rect 316794 678218 316826 678454
rect 317062 678218 317146 678454
rect 317382 678218 317414 678454
rect 316794 678134 317414 678218
rect 316794 677898 316826 678134
rect 317062 677898 317146 678134
rect 317382 677898 317414 678134
rect 316794 642454 317414 677898
rect 316794 642218 316826 642454
rect 317062 642218 317146 642454
rect 317382 642218 317414 642454
rect 316794 642134 317414 642218
rect 316794 641898 316826 642134
rect 317062 641898 317146 642134
rect 317382 641898 317414 642134
rect 316794 606454 317414 641898
rect 316794 606218 316826 606454
rect 317062 606218 317146 606454
rect 317382 606218 317414 606454
rect 316794 606134 317414 606218
rect 316794 605898 316826 606134
rect 317062 605898 317146 606134
rect 317382 605898 317414 606134
rect 316794 570454 317414 605898
rect 316794 570218 316826 570454
rect 317062 570218 317146 570454
rect 317382 570218 317414 570454
rect 316794 570134 317414 570218
rect 316794 569898 316826 570134
rect 317062 569898 317146 570134
rect 317382 569898 317414 570134
rect 316794 534454 317414 569898
rect 316794 534218 316826 534454
rect 317062 534218 317146 534454
rect 317382 534218 317414 534454
rect 316794 534134 317414 534218
rect 316794 533898 316826 534134
rect 317062 533898 317146 534134
rect 317382 533898 317414 534134
rect 316794 498454 317414 533898
rect 316794 498218 316826 498454
rect 317062 498218 317146 498454
rect 317382 498218 317414 498454
rect 316794 498134 317414 498218
rect 316794 497898 316826 498134
rect 317062 497898 317146 498134
rect 317382 497898 317414 498134
rect 316794 462454 317414 497898
rect 316794 462218 316826 462454
rect 317062 462218 317146 462454
rect 317382 462218 317414 462454
rect 316794 462134 317414 462218
rect 316794 461898 316826 462134
rect 317062 461898 317146 462134
rect 317382 461898 317414 462134
rect 316794 426454 317414 461898
rect 316794 426218 316826 426454
rect 317062 426218 317146 426454
rect 317382 426218 317414 426454
rect 316794 426134 317414 426218
rect 316794 425898 316826 426134
rect 317062 425898 317146 426134
rect 317382 425898 317414 426134
rect 316794 390454 317414 425898
rect 316794 390218 316826 390454
rect 317062 390218 317146 390454
rect 317382 390218 317414 390454
rect 316794 390134 317414 390218
rect 316794 389898 316826 390134
rect 317062 389898 317146 390134
rect 317382 389898 317414 390134
rect 316794 354454 317414 389898
rect 316794 354218 316826 354454
rect 317062 354218 317146 354454
rect 317382 354218 317414 354454
rect 316794 354134 317414 354218
rect 316794 353898 316826 354134
rect 317062 353898 317146 354134
rect 317382 353898 317414 354134
rect 316794 318454 317414 353898
rect 316794 318218 316826 318454
rect 317062 318218 317146 318454
rect 317382 318218 317414 318454
rect 316794 318134 317414 318218
rect 316794 317898 316826 318134
rect 317062 317898 317146 318134
rect 317382 317898 317414 318134
rect 316794 282454 317414 317898
rect 316794 282218 316826 282454
rect 317062 282218 317146 282454
rect 317382 282218 317414 282454
rect 316794 282134 317414 282218
rect 316794 281898 316826 282134
rect 317062 281898 317146 282134
rect 317382 281898 317414 282134
rect 316794 246454 317414 281898
rect 316794 246218 316826 246454
rect 317062 246218 317146 246454
rect 317382 246218 317414 246454
rect 316794 246134 317414 246218
rect 316794 245898 316826 246134
rect 317062 245898 317146 246134
rect 317382 245898 317414 246134
rect 316794 210454 317414 245898
rect 316794 210218 316826 210454
rect 317062 210218 317146 210454
rect 317382 210218 317414 210454
rect 316794 210134 317414 210218
rect 316794 209898 316826 210134
rect 317062 209898 317146 210134
rect 317382 209898 317414 210134
rect 316794 174454 317414 209898
rect 316794 174218 316826 174454
rect 317062 174218 317146 174454
rect 317382 174218 317414 174454
rect 316794 174134 317414 174218
rect 316794 173898 316826 174134
rect 317062 173898 317146 174134
rect 317382 173898 317414 174134
rect 316794 138454 317414 173898
rect 316794 138218 316826 138454
rect 317062 138218 317146 138454
rect 317382 138218 317414 138454
rect 316794 138134 317414 138218
rect 316794 137898 316826 138134
rect 317062 137898 317146 138134
rect 317382 137898 317414 138134
rect 316794 102454 317414 137898
rect 316794 102218 316826 102454
rect 317062 102218 317146 102454
rect 317382 102218 317414 102454
rect 316794 102134 317414 102218
rect 316794 101898 316826 102134
rect 317062 101898 317146 102134
rect 317382 101898 317414 102134
rect 316794 66454 317414 101898
rect 316794 66218 316826 66454
rect 317062 66218 317146 66454
rect 317382 66218 317414 66454
rect 316794 66134 317414 66218
rect 316794 65898 316826 66134
rect 317062 65898 317146 66134
rect 317382 65898 317414 66134
rect 316794 30454 317414 65898
rect 316794 30218 316826 30454
rect 317062 30218 317146 30454
rect 317382 30218 317414 30454
rect 316794 30134 317414 30218
rect 316794 29898 316826 30134
rect 317062 29898 317146 30134
rect 317382 29898 317414 30134
rect 316794 -6106 317414 29898
rect 316794 -6342 316826 -6106
rect 317062 -6342 317146 -6106
rect 317382 -6342 317414 -6106
rect 316794 -6426 317414 -6342
rect 316794 -6662 316826 -6426
rect 317062 -6662 317146 -6426
rect 317382 -6662 317414 -6426
rect 316794 -7654 317414 -6662
rect 321294 711558 321914 711590
rect 321294 711322 321326 711558
rect 321562 711322 321646 711558
rect 321882 711322 321914 711558
rect 321294 711238 321914 711322
rect 321294 711002 321326 711238
rect 321562 711002 321646 711238
rect 321882 711002 321914 711238
rect 321294 682954 321914 711002
rect 321294 682718 321326 682954
rect 321562 682718 321646 682954
rect 321882 682718 321914 682954
rect 321294 682634 321914 682718
rect 321294 682398 321326 682634
rect 321562 682398 321646 682634
rect 321882 682398 321914 682634
rect 321294 646954 321914 682398
rect 321294 646718 321326 646954
rect 321562 646718 321646 646954
rect 321882 646718 321914 646954
rect 321294 646634 321914 646718
rect 321294 646398 321326 646634
rect 321562 646398 321646 646634
rect 321882 646398 321914 646634
rect 321294 610954 321914 646398
rect 321294 610718 321326 610954
rect 321562 610718 321646 610954
rect 321882 610718 321914 610954
rect 321294 610634 321914 610718
rect 321294 610398 321326 610634
rect 321562 610398 321646 610634
rect 321882 610398 321914 610634
rect 321294 574954 321914 610398
rect 321294 574718 321326 574954
rect 321562 574718 321646 574954
rect 321882 574718 321914 574954
rect 321294 574634 321914 574718
rect 321294 574398 321326 574634
rect 321562 574398 321646 574634
rect 321882 574398 321914 574634
rect 321294 538954 321914 574398
rect 321294 538718 321326 538954
rect 321562 538718 321646 538954
rect 321882 538718 321914 538954
rect 321294 538634 321914 538718
rect 321294 538398 321326 538634
rect 321562 538398 321646 538634
rect 321882 538398 321914 538634
rect 321294 502954 321914 538398
rect 321294 502718 321326 502954
rect 321562 502718 321646 502954
rect 321882 502718 321914 502954
rect 321294 502634 321914 502718
rect 321294 502398 321326 502634
rect 321562 502398 321646 502634
rect 321882 502398 321914 502634
rect 321294 466954 321914 502398
rect 321294 466718 321326 466954
rect 321562 466718 321646 466954
rect 321882 466718 321914 466954
rect 321294 466634 321914 466718
rect 321294 466398 321326 466634
rect 321562 466398 321646 466634
rect 321882 466398 321914 466634
rect 321294 430954 321914 466398
rect 321294 430718 321326 430954
rect 321562 430718 321646 430954
rect 321882 430718 321914 430954
rect 321294 430634 321914 430718
rect 321294 430398 321326 430634
rect 321562 430398 321646 430634
rect 321882 430398 321914 430634
rect 321294 394954 321914 430398
rect 321294 394718 321326 394954
rect 321562 394718 321646 394954
rect 321882 394718 321914 394954
rect 321294 394634 321914 394718
rect 321294 394398 321326 394634
rect 321562 394398 321646 394634
rect 321882 394398 321914 394634
rect 321294 358954 321914 394398
rect 321294 358718 321326 358954
rect 321562 358718 321646 358954
rect 321882 358718 321914 358954
rect 321294 358634 321914 358718
rect 321294 358398 321326 358634
rect 321562 358398 321646 358634
rect 321882 358398 321914 358634
rect 321294 322954 321914 358398
rect 321294 322718 321326 322954
rect 321562 322718 321646 322954
rect 321882 322718 321914 322954
rect 321294 322634 321914 322718
rect 321294 322398 321326 322634
rect 321562 322398 321646 322634
rect 321882 322398 321914 322634
rect 321294 286954 321914 322398
rect 321294 286718 321326 286954
rect 321562 286718 321646 286954
rect 321882 286718 321914 286954
rect 321294 286634 321914 286718
rect 321294 286398 321326 286634
rect 321562 286398 321646 286634
rect 321882 286398 321914 286634
rect 321294 250954 321914 286398
rect 321294 250718 321326 250954
rect 321562 250718 321646 250954
rect 321882 250718 321914 250954
rect 321294 250634 321914 250718
rect 321294 250398 321326 250634
rect 321562 250398 321646 250634
rect 321882 250398 321914 250634
rect 321294 214954 321914 250398
rect 321294 214718 321326 214954
rect 321562 214718 321646 214954
rect 321882 214718 321914 214954
rect 321294 214634 321914 214718
rect 321294 214398 321326 214634
rect 321562 214398 321646 214634
rect 321882 214398 321914 214634
rect 321294 178954 321914 214398
rect 321294 178718 321326 178954
rect 321562 178718 321646 178954
rect 321882 178718 321914 178954
rect 321294 178634 321914 178718
rect 321294 178398 321326 178634
rect 321562 178398 321646 178634
rect 321882 178398 321914 178634
rect 321294 142954 321914 178398
rect 321294 142718 321326 142954
rect 321562 142718 321646 142954
rect 321882 142718 321914 142954
rect 321294 142634 321914 142718
rect 321294 142398 321326 142634
rect 321562 142398 321646 142634
rect 321882 142398 321914 142634
rect 321294 106954 321914 142398
rect 321294 106718 321326 106954
rect 321562 106718 321646 106954
rect 321882 106718 321914 106954
rect 321294 106634 321914 106718
rect 321294 106398 321326 106634
rect 321562 106398 321646 106634
rect 321882 106398 321914 106634
rect 321294 70954 321914 106398
rect 321294 70718 321326 70954
rect 321562 70718 321646 70954
rect 321882 70718 321914 70954
rect 321294 70634 321914 70718
rect 321294 70398 321326 70634
rect 321562 70398 321646 70634
rect 321882 70398 321914 70634
rect 321294 34954 321914 70398
rect 321294 34718 321326 34954
rect 321562 34718 321646 34954
rect 321882 34718 321914 34954
rect 321294 34634 321914 34718
rect 321294 34398 321326 34634
rect 321562 34398 321646 34634
rect 321882 34398 321914 34634
rect 321294 -7066 321914 34398
rect 321294 -7302 321326 -7066
rect 321562 -7302 321646 -7066
rect 321882 -7302 321914 -7066
rect 321294 -7386 321914 -7302
rect 321294 -7622 321326 -7386
rect 321562 -7622 321646 -7386
rect 321882 -7622 321914 -7386
rect 321294 -7654 321914 -7622
rect 325794 704838 326414 711590
rect 325794 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 326414 704838
rect 325794 704518 326414 704602
rect 325794 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 326414 704518
rect 325794 687454 326414 704282
rect 325794 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 326414 687454
rect 325794 687134 326414 687218
rect 325794 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 326414 687134
rect 325794 651454 326414 686898
rect 325794 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 326414 651454
rect 325794 651134 326414 651218
rect 325794 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 326414 651134
rect 325794 615454 326414 650898
rect 325794 615218 325826 615454
rect 326062 615218 326146 615454
rect 326382 615218 326414 615454
rect 325794 615134 326414 615218
rect 325794 614898 325826 615134
rect 326062 614898 326146 615134
rect 326382 614898 326414 615134
rect 325794 579454 326414 614898
rect 325794 579218 325826 579454
rect 326062 579218 326146 579454
rect 326382 579218 326414 579454
rect 325794 579134 326414 579218
rect 325794 578898 325826 579134
rect 326062 578898 326146 579134
rect 326382 578898 326414 579134
rect 325794 543454 326414 578898
rect 325794 543218 325826 543454
rect 326062 543218 326146 543454
rect 326382 543218 326414 543454
rect 325794 543134 326414 543218
rect 325794 542898 325826 543134
rect 326062 542898 326146 543134
rect 326382 542898 326414 543134
rect 325794 507454 326414 542898
rect 325794 507218 325826 507454
rect 326062 507218 326146 507454
rect 326382 507218 326414 507454
rect 325794 507134 326414 507218
rect 325794 506898 325826 507134
rect 326062 506898 326146 507134
rect 326382 506898 326414 507134
rect 325794 471454 326414 506898
rect 325794 471218 325826 471454
rect 326062 471218 326146 471454
rect 326382 471218 326414 471454
rect 325794 471134 326414 471218
rect 325794 470898 325826 471134
rect 326062 470898 326146 471134
rect 326382 470898 326414 471134
rect 325794 435454 326414 470898
rect 325794 435218 325826 435454
rect 326062 435218 326146 435454
rect 326382 435218 326414 435454
rect 325794 435134 326414 435218
rect 325794 434898 325826 435134
rect 326062 434898 326146 435134
rect 326382 434898 326414 435134
rect 325794 399454 326414 434898
rect 325794 399218 325826 399454
rect 326062 399218 326146 399454
rect 326382 399218 326414 399454
rect 325794 399134 326414 399218
rect 325794 398898 325826 399134
rect 326062 398898 326146 399134
rect 326382 398898 326414 399134
rect 325794 363454 326414 398898
rect 325794 363218 325826 363454
rect 326062 363218 326146 363454
rect 326382 363218 326414 363454
rect 325794 363134 326414 363218
rect 325794 362898 325826 363134
rect 326062 362898 326146 363134
rect 326382 362898 326414 363134
rect 325794 327454 326414 362898
rect 325794 327218 325826 327454
rect 326062 327218 326146 327454
rect 326382 327218 326414 327454
rect 325794 327134 326414 327218
rect 325794 326898 325826 327134
rect 326062 326898 326146 327134
rect 326382 326898 326414 327134
rect 325794 291454 326414 326898
rect 325794 291218 325826 291454
rect 326062 291218 326146 291454
rect 326382 291218 326414 291454
rect 325794 291134 326414 291218
rect 325794 290898 325826 291134
rect 326062 290898 326146 291134
rect 326382 290898 326414 291134
rect 325794 255454 326414 290898
rect 325794 255218 325826 255454
rect 326062 255218 326146 255454
rect 326382 255218 326414 255454
rect 325794 255134 326414 255218
rect 325794 254898 325826 255134
rect 326062 254898 326146 255134
rect 326382 254898 326414 255134
rect 325794 219454 326414 254898
rect 325794 219218 325826 219454
rect 326062 219218 326146 219454
rect 326382 219218 326414 219454
rect 325794 219134 326414 219218
rect 325794 218898 325826 219134
rect 326062 218898 326146 219134
rect 326382 218898 326414 219134
rect 325794 183454 326414 218898
rect 325794 183218 325826 183454
rect 326062 183218 326146 183454
rect 326382 183218 326414 183454
rect 325794 183134 326414 183218
rect 325794 182898 325826 183134
rect 326062 182898 326146 183134
rect 326382 182898 326414 183134
rect 325794 147454 326414 182898
rect 325794 147218 325826 147454
rect 326062 147218 326146 147454
rect 326382 147218 326414 147454
rect 325794 147134 326414 147218
rect 325794 146898 325826 147134
rect 326062 146898 326146 147134
rect 326382 146898 326414 147134
rect 325794 111454 326414 146898
rect 325794 111218 325826 111454
rect 326062 111218 326146 111454
rect 326382 111218 326414 111454
rect 325794 111134 326414 111218
rect 325794 110898 325826 111134
rect 326062 110898 326146 111134
rect 326382 110898 326414 111134
rect 325794 75454 326414 110898
rect 325794 75218 325826 75454
rect 326062 75218 326146 75454
rect 326382 75218 326414 75454
rect 325794 75134 326414 75218
rect 325794 74898 325826 75134
rect 326062 74898 326146 75134
rect 326382 74898 326414 75134
rect 325794 39454 326414 74898
rect 325794 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 326414 39454
rect 325794 39134 326414 39218
rect 325794 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 326414 39134
rect 325794 3454 326414 38898
rect 325794 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 326414 3454
rect 325794 3134 326414 3218
rect 325794 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 326414 3134
rect 325794 -346 326414 2898
rect 325794 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 326414 -346
rect 325794 -666 326414 -582
rect 325794 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 326414 -666
rect 325794 -7654 326414 -902
rect 330294 705798 330914 711590
rect 330294 705562 330326 705798
rect 330562 705562 330646 705798
rect 330882 705562 330914 705798
rect 330294 705478 330914 705562
rect 330294 705242 330326 705478
rect 330562 705242 330646 705478
rect 330882 705242 330914 705478
rect 330294 691954 330914 705242
rect 330294 691718 330326 691954
rect 330562 691718 330646 691954
rect 330882 691718 330914 691954
rect 330294 691634 330914 691718
rect 330294 691398 330326 691634
rect 330562 691398 330646 691634
rect 330882 691398 330914 691634
rect 330294 655954 330914 691398
rect 330294 655718 330326 655954
rect 330562 655718 330646 655954
rect 330882 655718 330914 655954
rect 330294 655634 330914 655718
rect 330294 655398 330326 655634
rect 330562 655398 330646 655634
rect 330882 655398 330914 655634
rect 330294 619954 330914 655398
rect 330294 619718 330326 619954
rect 330562 619718 330646 619954
rect 330882 619718 330914 619954
rect 330294 619634 330914 619718
rect 330294 619398 330326 619634
rect 330562 619398 330646 619634
rect 330882 619398 330914 619634
rect 330294 583954 330914 619398
rect 330294 583718 330326 583954
rect 330562 583718 330646 583954
rect 330882 583718 330914 583954
rect 330294 583634 330914 583718
rect 330294 583398 330326 583634
rect 330562 583398 330646 583634
rect 330882 583398 330914 583634
rect 330294 547954 330914 583398
rect 330294 547718 330326 547954
rect 330562 547718 330646 547954
rect 330882 547718 330914 547954
rect 330294 547634 330914 547718
rect 330294 547398 330326 547634
rect 330562 547398 330646 547634
rect 330882 547398 330914 547634
rect 330294 511954 330914 547398
rect 330294 511718 330326 511954
rect 330562 511718 330646 511954
rect 330882 511718 330914 511954
rect 330294 511634 330914 511718
rect 330294 511398 330326 511634
rect 330562 511398 330646 511634
rect 330882 511398 330914 511634
rect 330294 475954 330914 511398
rect 330294 475718 330326 475954
rect 330562 475718 330646 475954
rect 330882 475718 330914 475954
rect 330294 475634 330914 475718
rect 330294 475398 330326 475634
rect 330562 475398 330646 475634
rect 330882 475398 330914 475634
rect 330294 439954 330914 475398
rect 330294 439718 330326 439954
rect 330562 439718 330646 439954
rect 330882 439718 330914 439954
rect 330294 439634 330914 439718
rect 330294 439398 330326 439634
rect 330562 439398 330646 439634
rect 330882 439398 330914 439634
rect 330294 403954 330914 439398
rect 330294 403718 330326 403954
rect 330562 403718 330646 403954
rect 330882 403718 330914 403954
rect 330294 403634 330914 403718
rect 330294 403398 330326 403634
rect 330562 403398 330646 403634
rect 330882 403398 330914 403634
rect 330294 367954 330914 403398
rect 330294 367718 330326 367954
rect 330562 367718 330646 367954
rect 330882 367718 330914 367954
rect 330294 367634 330914 367718
rect 330294 367398 330326 367634
rect 330562 367398 330646 367634
rect 330882 367398 330914 367634
rect 330294 331954 330914 367398
rect 330294 331718 330326 331954
rect 330562 331718 330646 331954
rect 330882 331718 330914 331954
rect 330294 331634 330914 331718
rect 330294 331398 330326 331634
rect 330562 331398 330646 331634
rect 330882 331398 330914 331634
rect 330294 295954 330914 331398
rect 330294 295718 330326 295954
rect 330562 295718 330646 295954
rect 330882 295718 330914 295954
rect 330294 295634 330914 295718
rect 330294 295398 330326 295634
rect 330562 295398 330646 295634
rect 330882 295398 330914 295634
rect 330294 259954 330914 295398
rect 330294 259718 330326 259954
rect 330562 259718 330646 259954
rect 330882 259718 330914 259954
rect 330294 259634 330914 259718
rect 330294 259398 330326 259634
rect 330562 259398 330646 259634
rect 330882 259398 330914 259634
rect 330294 223954 330914 259398
rect 330294 223718 330326 223954
rect 330562 223718 330646 223954
rect 330882 223718 330914 223954
rect 330294 223634 330914 223718
rect 330294 223398 330326 223634
rect 330562 223398 330646 223634
rect 330882 223398 330914 223634
rect 330294 187954 330914 223398
rect 330294 187718 330326 187954
rect 330562 187718 330646 187954
rect 330882 187718 330914 187954
rect 330294 187634 330914 187718
rect 330294 187398 330326 187634
rect 330562 187398 330646 187634
rect 330882 187398 330914 187634
rect 330294 151954 330914 187398
rect 330294 151718 330326 151954
rect 330562 151718 330646 151954
rect 330882 151718 330914 151954
rect 330294 151634 330914 151718
rect 330294 151398 330326 151634
rect 330562 151398 330646 151634
rect 330882 151398 330914 151634
rect 330294 115954 330914 151398
rect 330294 115718 330326 115954
rect 330562 115718 330646 115954
rect 330882 115718 330914 115954
rect 330294 115634 330914 115718
rect 330294 115398 330326 115634
rect 330562 115398 330646 115634
rect 330882 115398 330914 115634
rect 330294 79954 330914 115398
rect 330294 79718 330326 79954
rect 330562 79718 330646 79954
rect 330882 79718 330914 79954
rect 330294 79634 330914 79718
rect 330294 79398 330326 79634
rect 330562 79398 330646 79634
rect 330882 79398 330914 79634
rect 330294 43954 330914 79398
rect 330294 43718 330326 43954
rect 330562 43718 330646 43954
rect 330882 43718 330914 43954
rect 330294 43634 330914 43718
rect 330294 43398 330326 43634
rect 330562 43398 330646 43634
rect 330882 43398 330914 43634
rect 330294 7954 330914 43398
rect 330294 7718 330326 7954
rect 330562 7718 330646 7954
rect 330882 7718 330914 7954
rect 330294 7634 330914 7718
rect 330294 7398 330326 7634
rect 330562 7398 330646 7634
rect 330882 7398 330914 7634
rect 330294 -1306 330914 7398
rect 330294 -1542 330326 -1306
rect 330562 -1542 330646 -1306
rect 330882 -1542 330914 -1306
rect 330294 -1626 330914 -1542
rect 330294 -1862 330326 -1626
rect 330562 -1862 330646 -1626
rect 330882 -1862 330914 -1626
rect 330294 -7654 330914 -1862
rect 334794 706758 335414 711590
rect 334794 706522 334826 706758
rect 335062 706522 335146 706758
rect 335382 706522 335414 706758
rect 334794 706438 335414 706522
rect 334794 706202 334826 706438
rect 335062 706202 335146 706438
rect 335382 706202 335414 706438
rect 334794 696454 335414 706202
rect 334794 696218 334826 696454
rect 335062 696218 335146 696454
rect 335382 696218 335414 696454
rect 334794 696134 335414 696218
rect 334794 695898 334826 696134
rect 335062 695898 335146 696134
rect 335382 695898 335414 696134
rect 334794 660454 335414 695898
rect 334794 660218 334826 660454
rect 335062 660218 335146 660454
rect 335382 660218 335414 660454
rect 334794 660134 335414 660218
rect 334794 659898 334826 660134
rect 335062 659898 335146 660134
rect 335382 659898 335414 660134
rect 334794 624454 335414 659898
rect 334794 624218 334826 624454
rect 335062 624218 335146 624454
rect 335382 624218 335414 624454
rect 334794 624134 335414 624218
rect 334794 623898 334826 624134
rect 335062 623898 335146 624134
rect 335382 623898 335414 624134
rect 334794 588454 335414 623898
rect 334794 588218 334826 588454
rect 335062 588218 335146 588454
rect 335382 588218 335414 588454
rect 334794 588134 335414 588218
rect 334794 587898 334826 588134
rect 335062 587898 335146 588134
rect 335382 587898 335414 588134
rect 334794 552454 335414 587898
rect 334794 552218 334826 552454
rect 335062 552218 335146 552454
rect 335382 552218 335414 552454
rect 334794 552134 335414 552218
rect 334794 551898 334826 552134
rect 335062 551898 335146 552134
rect 335382 551898 335414 552134
rect 334794 516454 335414 551898
rect 334794 516218 334826 516454
rect 335062 516218 335146 516454
rect 335382 516218 335414 516454
rect 334794 516134 335414 516218
rect 334794 515898 334826 516134
rect 335062 515898 335146 516134
rect 335382 515898 335414 516134
rect 334794 480454 335414 515898
rect 334794 480218 334826 480454
rect 335062 480218 335146 480454
rect 335382 480218 335414 480454
rect 334794 480134 335414 480218
rect 334794 479898 334826 480134
rect 335062 479898 335146 480134
rect 335382 479898 335414 480134
rect 334794 444454 335414 479898
rect 334794 444218 334826 444454
rect 335062 444218 335146 444454
rect 335382 444218 335414 444454
rect 334794 444134 335414 444218
rect 334794 443898 334826 444134
rect 335062 443898 335146 444134
rect 335382 443898 335414 444134
rect 334794 408454 335414 443898
rect 334794 408218 334826 408454
rect 335062 408218 335146 408454
rect 335382 408218 335414 408454
rect 334794 408134 335414 408218
rect 334794 407898 334826 408134
rect 335062 407898 335146 408134
rect 335382 407898 335414 408134
rect 334794 372454 335414 407898
rect 334794 372218 334826 372454
rect 335062 372218 335146 372454
rect 335382 372218 335414 372454
rect 334794 372134 335414 372218
rect 334794 371898 334826 372134
rect 335062 371898 335146 372134
rect 335382 371898 335414 372134
rect 334794 336454 335414 371898
rect 334794 336218 334826 336454
rect 335062 336218 335146 336454
rect 335382 336218 335414 336454
rect 334794 336134 335414 336218
rect 334794 335898 334826 336134
rect 335062 335898 335146 336134
rect 335382 335898 335414 336134
rect 334794 300454 335414 335898
rect 334794 300218 334826 300454
rect 335062 300218 335146 300454
rect 335382 300218 335414 300454
rect 334794 300134 335414 300218
rect 334794 299898 334826 300134
rect 335062 299898 335146 300134
rect 335382 299898 335414 300134
rect 334794 264454 335414 299898
rect 334794 264218 334826 264454
rect 335062 264218 335146 264454
rect 335382 264218 335414 264454
rect 334794 264134 335414 264218
rect 334794 263898 334826 264134
rect 335062 263898 335146 264134
rect 335382 263898 335414 264134
rect 334794 228454 335414 263898
rect 334794 228218 334826 228454
rect 335062 228218 335146 228454
rect 335382 228218 335414 228454
rect 334794 228134 335414 228218
rect 334794 227898 334826 228134
rect 335062 227898 335146 228134
rect 335382 227898 335414 228134
rect 334794 192454 335414 227898
rect 334794 192218 334826 192454
rect 335062 192218 335146 192454
rect 335382 192218 335414 192454
rect 334794 192134 335414 192218
rect 334794 191898 334826 192134
rect 335062 191898 335146 192134
rect 335382 191898 335414 192134
rect 334794 156454 335414 191898
rect 334794 156218 334826 156454
rect 335062 156218 335146 156454
rect 335382 156218 335414 156454
rect 334794 156134 335414 156218
rect 334794 155898 334826 156134
rect 335062 155898 335146 156134
rect 335382 155898 335414 156134
rect 334794 120454 335414 155898
rect 334794 120218 334826 120454
rect 335062 120218 335146 120454
rect 335382 120218 335414 120454
rect 334794 120134 335414 120218
rect 334794 119898 334826 120134
rect 335062 119898 335146 120134
rect 335382 119898 335414 120134
rect 334794 84454 335414 119898
rect 334794 84218 334826 84454
rect 335062 84218 335146 84454
rect 335382 84218 335414 84454
rect 334794 84134 335414 84218
rect 334794 83898 334826 84134
rect 335062 83898 335146 84134
rect 335382 83898 335414 84134
rect 334794 48454 335414 83898
rect 334794 48218 334826 48454
rect 335062 48218 335146 48454
rect 335382 48218 335414 48454
rect 334794 48134 335414 48218
rect 334794 47898 334826 48134
rect 335062 47898 335146 48134
rect 335382 47898 335414 48134
rect 334794 12454 335414 47898
rect 334794 12218 334826 12454
rect 335062 12218 335146 12454
rect 335382 12218 335414 12454
rect 334794 12134 335414 12218
rect 334794 11898 334826 12134
rect 335062 11898 335146 12134
rect 335382 11898 335414 12134
rect 334794 -2266 335414 11898
rect 334794 -2502 334826 -2266
rect 335062 -2502 335146 -2266
rect 335382 -2502 335414 -2266
rect 334794 -2586 335414 -2502
rect 334794 -2822 334826 -2586
rect 335062 -2822 335146 -2586
rect 335382 -2822 335414 -2586
rect 334794 -7654 335414 -2822
rect 339294 707718 339914 711590
rect 339294 707482 339326 707718
rect 339562 707482 339646 707718
rect 339882 707482 339914 707718
rect 339294 707398 339914 707482
rect 339294 707162 339326 707398
rect 339562 707162 339646 707398
rect 339882 707162 339914 707398
rect 339294 700954 339914 707162
rect 339294 700718 339326 700954
rect 339562 700718 339646 700954
rect 339882 700718 339914 700954
rect 339294 700634 339914 700718
rect 339294 700398 339326 700634
rect 339562 700398 339646 700634
rect 339882 700398 339914 700634
rect 339294 664954 339914 700398
rect 339294 664718 339326 664954
rect 339562 664718 339646 664954
rect 339882 664718 339914 664954
rect 339294 664634 339914 664718
rect 339294 664398 339326 664634
rect 339562 664398 339646 664634
rect 339882 664398 339914 664634
rect 339294 628954 339914 664398
rect 339294 628718 339326 628954
rect 339562 628718 339646 628954
rect 339882 628718 339914 628954
rect 339294 628634 339914 628718
rect 339294 628398 339326 628634
rect 339562 628398 339646 628634
rect 339882 628398 339914 628634
rect 339294 592954 339914 628398
rect 339294 592718 339326 592954
rect 339562 592718 339646 592954
rect 339882 592718 339914 592954
rect 339294 592634 339914 592718
rect 339294 592398 339326 592634
rect 339562 592398 339646 592634
rect 339882 592398 339914 592634
rect 339294 556954 339914 592398
rect 339294 556718 339326 556954
rect 339562 556718 339646 556954
rect 339882 556718 339914 556954
rect 339294 556634 339914 556718
rect 339294 556398 339326 556634
rect 339562 556398 339646 556634
rect 339882 556398 339914 556634
rect 339294 520954 339914 556398
rect 339294 520718 339326 520954
rect 339562 520718 339646 520954
rect 339882 520718 339914 520954
rect 339294 520634 339914 520718
rect 339294 520398 339326 520634
rect 339562 520398 339646 520634
rect 339882 520398 339914 520634
rect 339294 484954 339914 520398
rect 339294 484718 339326 484954
rect 339562 484718 339646 484954
rect 339882 484718 339914 484954
rect 339294 484634 339914 484718
rect 339294 484398 339326 484634
rect 339562 484398 339646 484634
rect 339882 484398 339914 484634
rect 339294 448954 339914 484398
rect 339294 448718 339326 448954
rect 339562 448718 339646 448954
rect 339882 448718 339914 448954
rect 339294 448634 339914 448718
rect 339294 448398 339326 448634
rect 339562 448398 339646 448634
rect 339882 448398 339914 448634
rect 339294 412954 339914 448398
rect 339294 412718 339326 412954
rect 339562 412718 339646 412954
rect 339882 412718 339914 412954
rect 339294 412634 339914 412718
rect 339294 412398 339326 412634
rect 339562 412398 339646 412634
rect 339882 412398 339914 412634
rect 339294 376954 339914 412398
rect 339294 376718 339326 376954
rect 339562 376718 339646 376954
rect 339882 376718 339914 376954
rect 339294 376634 339914 376718
rect 339294 376398 339326 376634
rect 339562 376398 339646 376634
rect 339882 376398 339914 376634
rect 339294 340954 339914 376398
rect 339294 340718 339326 340954
rect 339562 340718 339646 340954
rect 339882 340718 339914 340954
rect 339294 340634 339914 340718
rect 339294 340398 339326 340634
rect 339562 340398 339646 340634
rect 339882 340398 339914 340634
rect 339294 304954 339914 340398
rect 339294 304718 339326 304954
rect 339562 304718 339646 304954
rect 339882 304718 339914 304954
rect 339294 304634 339914 304718
rect 339294 304398 339326 304634
rect 339562 304398 339646 304634
rect 339882 304398 339914 304634
rect 339294 268954 339914 304398
rect 339294 268718 339326 268954
rect 339562 268718 339646 268954
rect 339882 268718 339914 268954
rect 339294 268634 339914 268718
rect 339294 268398 339326 268634
rect 339562 268398 339646 268634
rect 339882 268398 339914 268634
rect 339294 232954 339914 268398
rect 339294 232718 339326 232954
rect 339562 232718 339646 232954
rect 339882 232718 339914 232954
rect 339294 232634 339914 232718
rect 339294 232398 339326 232634
rect 339562 232398 339646 232634
rect 339882 232398 339914 232634
rect 339294 196954 339914 232398
rect 339294 196718 339326 196954
rect 339562 196718 339646 196954
rect 339882 196718 339914 196954
rect 339294 196634 339914 196718
rect 339294 196398 339326 196634
rect 339562 196398 339646 196634
rect 339882 196398 339914 196634
rect 339294 160954 339914 196398
rect 339294 160718 339326 160954
rect 339562 160718 339646 160954
rect 339882 160718 339914 160954
rect 339294 160634 339914 160718
rect 339294 160398 339326 160634
rect 339562 160398 339646 160634
rect 339882 160398 339914 160634
rect 339294 124954 339914 160398
rect 339294 124718 339326 124954
rect 339562 124718 339646 124954
rect 339882 124718 339914 124954
rect 339294 124634 339914 124718
rect 339294 124398 339326 124634
rect 339562 124398 339646 124634
rect 339882 124398 339914 124634
rect 339294 88954 339914 124398
rect 339294 88718 339326 88954
rect 339562 88718 339646 88954
rect 339882 88718 339914 88954
rect 339294 88634 339914 88718
rect 339294 88398 339326 88634
rect 339562 88398 339646 88634
rect 339882 88398 339914 88634
rect 339294 52954 339914 88398
rect 339294 52718 339326 52954
rect 339562 52718 339646 52954
rect 339882 52718 339914 52954
rect 339294 52634 339914 52718
rect 339294 52398 339326 52634
rect 339562 52398 339646 52634
rect 339882 52398 339914 52634
rect 339294 16954 339914 52398
rect 339294 16718 339326 16954
rect 339562 16718 339646 16954
rect 339882 16718 339914 16954
rect 339294 16634 339914 16718
rect 339294 16398 339326 16634
rect 339562 16398 339646 16634
rect 339882 16398 339914 16634
rect 339294 -3226 339914 16398
rect 339294 -3462 339326 -3226
rect 339562 -3462 339646 -3226
rect 339882 -3462 339914 -3226
rect 339294 -3546 339914 -3462
rect 339294 -3782 339326 -3546
rect 339562 -3782 339646 -3546
rect 339882 -3782 339914 -3546
rect 339294 -7654 339914 -3782
rect 343794 708678 344414 711590
rect 343794 708442 343826 708678
rect 344062 708442 344146 708678
rect 344382 708442 344414 708678
rect 343794 708358 344414 708442
rect 343794 708122 343826 708358
rect 344062 708122 344146 708358
rect 344382 708122 344414 708358
rect 343794 669454 344414 708122
rect 343794 669218 343826 669454
rect 344062 669218 344146 669454
rect 344382 669218 344414 669454
rect 343794 669134 344414 669218
rect 343794 668898 343826 669134
rect 344062 668898 344146 669134
rect 344382 668898 344414 669134
rect 343794 633454 344414 668898
rect 343794 633218 343826 633454
rect 344062 633218 344146 633454
rect 344382 633218 344414 633454
rect 343794 633134 344414 633218
rect 343794 632898 343826 633134
rect 344062 632898 344146 633134
rect 344382 632898 344414 633134
rect 343794 597454 344414 632898
rect 343794 597218 343826 597454
rect 344062 597218 344146 597454
rect 344382 597218 344414 597454
rect 343794 597134 344414 597218
rect 343794 596898 343826 597134
rect 344062 596898 344146 597134
rect 344382 596898 344414 597134
rect 343794 561454 344414 596898
rect 343794 561218 343826 561454
rect 344062 561218 344146 561454
rect 344382 561218 344414 561454
rect 343794 561134 344414 561218
rect 343794 560898 343826 561134
rect 344062 560898 344146 561134
rect 344382 560898 344414 561134
rect 343794 525454 344414 560898
rect 343794 525218 343826 525454
rect 344062 525218 344146 525454
rect 344382 525218 344414 525454
rect 343794 525134 344414 525218
rect 343794 524898 343826 525134
rect 344062 524898 344146 525134
rect 344382 524898 344414 525134
rect 343794 489454 344414 524898
rect 343794 489218 343826 489454
rect 344062 489218 344146 489454
rect 344382 489218 344414 489454
rect 343794 489134 344414 489218
rect 343794 488898 343826 489134
rect 344062 488898 344146 489134
rect 344382 488898 344414 489134
rect 343794 453454 344414 488898
rect 343794 453218 343826 453454
rect 344062 453218 344146 453454
rect 344382 453218 344414 453454
rect 343794 453134 344414 453218
rect 343794 452898 343826 453134
rect 344062 452898 344146 453134
rect 344382 452898 344414 453134
rect 343794 417454 344414 452898
rect 343794 417218 343826 417454
rect 344062 417218 344146 417454
rect 344382 417218 344414 417454
rect 343794 417134 344414 417218
rect 343794 416898 343826 417134
rect 344062 416898 344146 417134
rect 344382 416898 344414 417134
rect 343794 381454 344414 416898
rect 343794 381218 343826 381454
rect 344062 381218 344146 381454
rect 344382 381218 344414 381454
rect 343794 381134 344414 381218
rect 343794 380898 343826 381134
rect 344062 380898 344146 381134
rect 344382 380898 344414 381134
rect 343794 345454 344414 380898
rect 343794 345218 343826 345454
rect 344062 345218 344146 345454
rect 344382 345218 344414 345454
rect 343794 345134 344414 345218
rect 343794 344898 343826 345134
rect 344062 344898 344146 345134
rect 344382 344898 344414 345134
rect 343794 309454 344414 344898
rect 343794 309218 343826 309454
rect 344062 309218 344146 309454
rect 344382 309218 344414 309454
rect 343794 309134 344414 309218
rect 343794 308898 343826 309134
rect 344062 308898 344146 309134
rect 344382 308898 344414 309134
rect 343794 273454 344414 308898
rect 343794 273218 343826 273454
rect 344062 273218 344146 273454
rect 344382 273218 344414 273454
rect 343794 273134 344414 273218
rect 343794 272898 343826 273134
rect 344062 272898 344146 273134
rect 344382 272898 344414 273134
rect 343794 237454 344414 272898
rect 343794 237218 343826 237454
rect 344062 237218 344146 237454
rect 344382 237218 344414 237454
rect 343794 237134 344414 237218
rect 343794 236898 343826 237134
rect 344062 236898 344146 237134
rect 344382 236898 344414 237134
rect 343794 201454 344414 236898
rect 343794 201218 343826 201454
rect 344062 201218 344146 201454
rect 344382 201218 344414 201454
rect 343794 201134 344414 201218
rect 343794 200898 343826 201134
rect 344062 200898 344146 201134
rect 344382 200898 344414 201134
rect 343794 165454 344414 200898
rect 343794 165218 343826 165454
rect 344062 165218 344146 165454
rect 344382 165218 344414 165454
rect 343794 165134 344414 165218
rect 343794 164898 343826 165134
rect 344062 164898 344146 165134
rect 344382 164898 344414 165134
rect 343794 129454 344414 164898
rect 343794 129218 343826 129454
rect 344062 129218 344146 129454
rect 344382 129218 344414 129454
rect 343794 129134 344414 129218
rect 343794 128898 343826 129134
rect 344062 128898 344146 129134
rect 344382 128898 344414 129134
rect 343794 93454 344414 128898
rect 343794 93218 343826 93454
rect 344062 93218 344146 93454
rect 344382 93218 344414 93454
rect 343794 93134 344414 93218
rect 343794 92898 343826 93134
rect 344062 92898 344146 93134
rect 344382 92898 344414 93134
rect 343794 57454 344414 92898
rect 343794 57218 343826 57454
rect 344062 57218 344146 57454
rect 344382 57218 344414 57454
rect 343794 57134 344414 57218
rect 343794 56898 343826 57134
rect 344062 56898 344146 57134
rect 344382 56898 344414 57134
rect 343794 21454 344414 56898
rect 343794 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 344414 21454
rect 343794 21134 344414 21218
rect 343794 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 344414 21134
rect 343794 -4186 344414 20898
rect 343794 -4422 343826 -4186
rect 344062 -4422 344146 -4186
rect 344382 -4422 344414 -4186
rect 343794 -4506 344414 -4422
rect 343794 -4742 343826 -4506
rect 344062 -4742 344146 -4506
rect 344382 -4742 344414 -4506
rect 343794 -7654 344414 -4742
rect 348294 709638 348914 711590
rect 348294 709402 348326 709638
rect 348562 709402 348646 709638
rect 348882 709402 348914 709638
rect 348294 709318 348914 709402
rect 348294 709082 348326 709318
rect 348562 709082 348646 709318
rect 348882 709082 348914 709318
rect 348294 673954 348914 709082
rect 348294 673718 348326 673954
rect 348562 673718 348646 673954
rect 348882 673718 348914 673954
rect 348294 673634 348914 673718
rect 348294 673398 348326 673634
rect 348562 673398 348646 673634
rect 348882 673398 348914 673634
rect 348294 637954 348914 673398
rect 348294 637718 348326 637954
rect 348562 637718 348646 637954
rect 348882 637718 348914 637954
rect 348294 637634 348914 637718
rect 348294 637398 348326 637634
rect 348562 637398 348646 637634
rect 348882 637398 348914 637634
rect 348294 601954 348914 637398
rect 348294 601718 348326 601954
rect 348562 601718 348646 601954
rect 348882 601718 348914 601954
rect 348294 601634 348914 601718
rect 348294 601398 348326 601634
rect 348562 601398 348646 601634
rect 348882 601398 348914 601634
rect 348294 565954 348914 601398
rect 348294 565718 348326 565954
rect 348562 565718 348646 565954
rect 348882 565718 348914 565954
rect 348294 565634 348914 565718
rect 348294 565398 348326 565634
rect 348562 565398 348646 565634
rect 348882 565398 348914 565634
rect 348294 529954 348914 565398
rect 348294 529718 348326 529954
rect 348562 529718 348646 529954
rect 348882 529718 348914 529954
rect 348294 529634 348914 529718
rect 348294 529398 348326 529634
rect 348562 529398 348646 529634
rect 348882 529398 348914 529634
rect 348294 493954 348914 529398
rect 348294 493718 348326 493954
rect 348562 493718 348646 493954
rect 348882 493718 348914 493954
rect 348294 493634 348914 493718
rect 348294 493398 348326 493634
rect 348562 493398 348646 493634
rect 348882 493398 348914 493634
rect 348294 457954 348914 493398
rect 348294 457718 348326 457954
rect 348562 457718 348646 457954
rect 348882 457718 348914 457954
rect 348294 457634 348914 457718
rect 348294 457398 348326 457634
rect 348562 457398 348646 457634
rect 348882 457398 348914 457634
rect 348294 421954 348914 457398
rect 348294 421718 348326 421954
rect 348562 421718 348646 421954
rect 348882 421718 348914 421954
rect 348294 421634 348914 421718
rect 348294 421398 348326 421634
rect 348562 421398 348646 421634
rect 348882 421398 348914 421634
rect 348294 385954 348914 421398
rect 348294 385718 348326 385954
rect 348562 385718 348646 385954
rect 348882 385718 348914 385954
rect 348294 385634 348914 385718
rect 348294 385398 348326 385634
rect 348562 385398 348646 385634
rect 348882 385398 348914 385634
rect 348294 349954 348914 385398
rect 348294 349718 348326 349954
rect 348562 349718 348646 349954
rect 348882 349718 348914 349954
rect 348294 349634 348914 349718
rect 348294 349398 348326 349634
rect 348562 349398 348646 349634
rect 348882 349398 348914 349634
rect 348294 313954 348914 349398
rect 348294 313718 348326 313954
rect 348562 313718 348646 313954
rect 348882 313718 348914 313954
rect 348294 313634 348914 313718
rect 348294 313398 348326 313634
rect 348562 313398 348646 313634
rect 348882 313398 348914 313634
rect 348294 277954 348914 313398
rect 348294 277718 348326 277954
rect 348562 277718 348646 277954
rect 348882 277718 348914 277954
rect 348294 277634 348914 277718
rect 348294 277398 348326 277634
rect 348562 277398 348646 277634
rect 348882 277398 348914 277634
rect 348294 241954 348914 277398
rect 348294 241718 348326 241954
rect 348562 241718 348646 241954
rect 348882 241718 348914 241954
rect 348294 241634 348914 241718
rect 348294 241398 348326 241634
rect 348562 241398 348646 241634
rect 348882 241398 348914 241634
rect 348294 205954 348914 241398
rect 348294 205718 348326 205954
rect 348562 205718 348646 205954
rect 348882 205718 348914 205954
rect 348294 205634 348914 205718
rect 348294 205398 348326 205634
rect 348562 205398 348646 205634
rect 348882 205398 348914 205634
rect 348294 169954 348914 205398
rect 348294 169718 348326 169954
rect 348562 169718 348646 169954
rect 348882 169718 348914 169954
rect 348294 169634 348914 169718
rect 348294 169398 348326 169634
rect 348562 169398 348646 169634
rect 348882 169398 348914 169634
rect 348294 133954 348914 169398
rect 348294 133718 348326 133954
rect 348562 133718 348646 133954
rect 348882 133718 348914 133954
rect 348294 133634 348914 133718
rect 348294 133398 348326 133634
rect 348562 133398 348646 133634
rect 348882 133398 348914 133634
rect 348294 97954 348914 133398
rect 348294 97718 348326 97954
rect 348562 97718 348646 97954
rect 348882 97718 348914 97954
rect 348294 97634 348914 97718
rect 348294 97398 348326 97634
rect 348562 97398 348646 97634
rect 348882 97398 348914 97634
rect 348294 61954 348914 97398
rect 348294 61718 348326 61954
rect 348562 61718 348646 61954
rect 348882 61718 348914 61954
rect 348294 61634 348914 61718
rect 348294 61398 348326 61634
rect 348562 61398 348646 61634
rect 348882 61398 348914 61634
rect 348294 25954 348914 61398
rect 348294 25718 348326 25954
rect 348562 25718 348646 25954
rect 348882 25718 348914 25954
rect 348294 25634 348914 25718
rect 348294 25398 348326 25634
rect 348562 25398 348646 25634
rect 348882 25398 348914 25634
rect 348294 -5146 348914 25398
rect 348294 -5382 348326 -5146
rect 348562 -5382 348646 -5146
rect 348882 -5382 348914 -5146
rect 348294 -5466 348914 -5382
rect 348294 -5702 348326 -5466
rect 348562 -5702 348646 -5466
rect 348882 -5702 348914 -5466
rect 348294 -7654 348914 -5702
rect 352794 710598 353414 711590
rect 352794 710362 352826 710598
rect 353062 710362 353146 710598
rect 353382 710362 353414 710598
rect 352794 710278 353414 710362
rect 352794 710042 352826 710278
rect 353062 710042 353146 710278
rect 353382 710042 353414 710278
rect 352794 678454 353414 710042
rect 352794 678218 352826 678454
rect 353062 678218 353146 678454
rect 353382 678218 353414 678454
rect 352794 678134 353414 678218
rect 352794 677898 352826 678134
rect 353062 677898 353146 678134
rect 353382 677898 353414 678134
rect 352794 642454 353414 677898
rect 352794 642218 352826 642454
rect 353062 642218 353146 642454
rect 353382 642218 353414 642454
rect 352794 642134 353414 642218
rect 352794 641898 352826 642134
rect 353062 641898 353146 642134
rect 353382 641898 353414 642134
rect 352794 606454 353414 641898
rect 352794 606218 352826 606454
rect 353062 606218 353146 606454
rect 353382 606218 353414 606454
rect 352794 606134 353414 606218
rect 352794 605898 352826 606134
rect 353062 605898 353146 606134
rect 353382 605898 353414 606134
rect 352794 570454 353414 605898
rect 352794 570218 352826 570454
rect 353062 570218 353146 570454
rect 353382 570218 353414 570454
rect 352794 570134 353414 570218
rect 352794 569898 352826 570134
rect 353062 569898 353146 570134
rect 353382 569898 353414 570134
rect 352794 534454 353414 569898
rect 352794 534218 352826 534454
rect 353062 534218 353146 534454
rect 353382 534218 353414 534454
rect 352794 534134 353414 534218
rect 352794 533898 352826 534134
rect 353062 533898 353146 534134
rect 353382 533898 353414 534134
rect 352794 498454 353414 533898
rect 352794 498218 352826 498454
rect 353062 498218 353146 498454
rect 353382 498218 353414 498454
rect 352794 498134 353414 498218
rect 352794 497898 352826 498134
rect 353062 497898 353146 498134
rect 353382 497898 353414 498134
rect 352794 462454 353414 497898
rect 352794 462218 352826 462454
rect 353062 462218 353146 462454
rect 353382 462218 353414 462454
rect 352794 462134 353414 462218
rect 352794 461898 352826 462134
rect 353062 461898 353146 462134
rect 353382 461898 353414 462134
rect 352794 426454 353414 461898
rect 352794 426218 352826 426454
rect 353062 426218 353146 426454
rect 353382 426218 353414 426454
rect 352794 426134 353414 426218
rect 352794 425898 352826 426134
rect 353062 425898 353146 426134
rect 353382 425898 353414 426134
rect 352794 390454 353414 425898
rect 352794 390218 352826 390454
rect 353062 390218 353146 390454
rect 353382 390218 353414 390454
rect 352794 390134 353414 390218
rect 352794 389898 352826 390134
rect 353062 389898 353146 390134
rect 353382 389898 353414 390134
rect 352794 354454 353414 389898
rect 352794 354218 352826 354454
rect 353062 354218 353146 354454
rect 353382 354218 353414 354454
rect 352794 354134 353414 354218
rect 352794 353898 352826 354134
rect 353062 353898 353146 354134
rect 353382 353898 353414 354134
rect 352794 318454 353414 353898
rect 352794 318218 352826 318454
rect 353062 318218 353146 318454
rect 353382 318218 353414 318454
rect 352794 318134 353414 318218
rect 352794 317898 352826 318134
rect 353062 317898 353146 318134
rect 353382 317898 353414 318134
rect 352794 282454 353414 317898
rect 352794 282218 352826 282454
rect 353062 282218 353146 282454
rect 353382 282218 353414 282454
rect 352794 282134 353414 282218
rect 352794 281898 352826 282134
rect 353062 281898 353146 282134
rect 353382 281898 353414 282134
rect 352794 246454 353414 281898
rect 352794 246218 352826 246454
rect 353062 246218 353146 246454
rect 353382 246218 353414 246454
rect 352794 246134 353414 246218
rect 352794 245898 352826 246134
rect 353062 245898 353146 246134
rect 353382 245898 353414 246134
rect 352794 210454 353414 245898
rect 352794 210218 352826 210454
rect 353062 210218 353146 210454
rect 353382 210218 353414 210454
rect 352794 210134 353414 210218
rect 352794 209898 352826 210134
rect 353062 209898 353146 210134
rect 353382 209898 353414 210134
rect 352794 174454 353414 209898
rect 352794 174218 352826 174454
rect 353062 174218 353146 174454
rect 353382 174218 353414 174454
rect 352794 174134 353414 174218
rect 352794 173898 352826 174134
rect 353062 173898 353146 174134
rect 353382 173898 353414 174134
rect 352794 138454 353414 173898
rect 352794 138218 352826 138454
rect 353062 138218 353146 138454
rect 353382 138218 353414 138454
rect 352794 138134 353414 138218
rect 352794 137898 352826 138134
rect 353062 137898 353146 138134
rect 353382 137898 353414 138134
rect 352794 102454 353414 137898
rect 352794 102218 352826 102454
rect 353062 102218 353146 102454
rect 353382 102218 353414 102454
rect 352794 102134 353414 102218
rect 352794 101898 352826 102134
rect 353062 101898 353146 102134
rect 353382 101898 353414 102134
rect 352794 66454 353414 101898
rect 352794 66218 352826 66454
rect 353062 66218 353146 66454
rect 353382 66218 353414 66454
rect 352794 66134 353414 66218
rect 352794 65898 352826 66134
rect 353062 65898 353146 66134
rect 353382 65898 353414 66134
rect 352794 30454 353414 65898
rect 352794 30218 352826 30454
rect 353062 30218 353146 30454
rect 353382 30218 353414 30454
rect 352794 30134 353414 30218
rect 352794 29898 352826 30134
rect 353062 29898 353146 30134
rect 353382 29898 353414 30134
rect 352794 -6106 353414 29898
rect 352794 -6342 352826 -6106
rect 353062 -6342 353146 -6106
rect 353382 -6342 353414 -6106
rect 352794 -6426 353414 -6342
rect 352794 -6662 352826 -6426
rect 353062 -6662 353146 -6426
rect 353382 -6662 353414 -6426
rect 352794 -7654 353414 -6662
rect 357294 711558 357914 711590
rect 357294 711322 357326 711558
rect 357562 711322 357646 711558
rect 357882 711322 357914 711558
rect 357294 711238 357914 711322
rect 357294 711002 357326 711238
rect 357562 711002 357646 711238
rect 357882 711002 357914 711238
rect 357294 682954 357914 711002
rect 357294 682718 357326 682954
rect 357562 682718 357646 682954
rect 357882 682718 357914 682954
rect 357294 682634 357914 682718
rect 357294 682398 357326 682634
rect 357562 682398 357646 682634
rect 357882 682398 357914 682634
rect 357294 646954 357914 682398
rect 357294 646718 357326 646954
rect 357562 646718 357646 646954
rect 357882 646718 357914 646954
rect 357294 646634 357914 646718
rect 357294 646398 357326 646634
rect 357562 646398 357646 646634
rect 357882 646398 357914 646634
rect 357294 610954 357914 646398
rect 357294 610718 357326 610954
rect 357562 610718 357646 610954
rect 357882 610718 357914 610954
rect 357294 610634 357914 610718
rect 357294 610398 357326 610634
rect 357562 610398 357646 610634
rect 357882 610398 357914 610634
rect 357294 574954 357914 610398
rect 357294 574718 357326 574954
rect 357562 574718 357646 574954
rect 357882 574718 357914 574954
rect 357294 574634 357914 574718
rect 357294 574398 357326 574634
rect 357562 574398 357646 574634
rect 357882 574398 357914 574634
rect 357294 538954 357914 574398
rect 357294 538718 357326 538954
rect 357562 538718 357646 538954
rect 357882 538718 357914 538954
rect 357294 538634 357914 538718
rect 357294 538398 357326 538634
rect 357562 538398 357646 538634
rect 357882 538398 357914 538634
rect 357294 502954 357914 538398
rect 357294 502718 357326 502954
rect 357562 502718 357646 502954
rect 357882 502718 357914 502954
rect 357294 502634 357914 502718
rect 357294 502398 357326 502634
rect 357562 502398 357646 502634
rect 357882 502398 357914 502634
rect 357294 466954 357914 502398
rect 357294 466718 357326 466954
rect 357562 466718 357646 466954
rect 357882 466718 357914 466954
rect 357294 466634 357914 466718
rect 357294 466398 357326 466634
rect 357562 466398 357646 466634
rect 357882 466398 357914 466634
rect 357294 430954 357914 466398
rect 357294 430718 357326 430954
rect 357562 430718 357646 430954
rect 357882 430718 357914 430954
rect 357294 430634 357914 430718
rect 357294 430398 357326 430634
rect 357562 430398 357646 430634
rect 357882 430398 357914 430634
rect 357294 394954 357914 430398
rect 357294 394718 357326 394954
rect 357562 394718 357646 394954
rect 357882 394718 357914 394954
rect 357294 394634 357914 394718
rect 357294 394398 357326 394634
rect 357562 394398 357646 394634
rect 357882 394398 357914 394634
rect 357294 358954 357914 394398
rect 357294 358718 357326 358954
rect 357562 358718 357646 358954
rect 357882 358718 357914 358954
rect 357294 358634 357914 358718
rect 357294 358398 357326 358634
rect 357562 358398 357646 358634
rect 357882 358398 357914 358634
rect 357294 322954 357914 358398
rect 357294 322718 357326 322954
rect 357562 322718 357646 322954
rect 357882 322718 357914 322954
rect 357294 322634 357914 322718
rect 357294 322398 357326 322634
rect 357562 322398 357646 322634
rect 357882 322398 357914 322634
rect 357294 286954 357914 322398
rect 357294 286718 357326 286954
rect 357562 286718 357646 286954
rect 357882 286718 357914 286954
rect 357294 286634 357914 286718
rect 357294 286398 357326 286634
rect 357562 286398 357646 286634
rect 357882 286398 357914 286634
rect 357294 250954 357914 286398
rect 357294 250718 357326 250954
rect 357562 250718 357646 250954
rect 357882 250718 357914 250954
rect 357294 250634 357914 250718
rect 357294 250398 357326 250634
rect 357562 250398 357646 250634
rect 357882 250398 357914 250634
rect 357294 214954 357914 250398
rect 357294 214718 357326 214954
rect 357562 214718 357646 214954
rect 357882 214718 357914 214954
rect 357294 214634 357914 214718
rect 357294 214398 357326 214634
rect 357562 214398 357646 214634
rect 357882 214398 357914 214634
rect 357294 178954 357914 214398
rect 357294 178718 357326 178954
rect 357562 178718 357646 178954
rect 357882 178718 357914 178954
rect 357294 178634 357914 178718
rect 357294 178398 357326 178634
rect 357562 178398 357646 178634
rect 357882 178398 357914 178634
rect 357294 142954 357914 178398
rect 357294 142718 357326 142954
rect 357562 142718 357646 142954
rect 357882 142718 357914 142954
rect 357294 142634 357914 142718
rect 357294 142398 357326 142634
rect 357562 142398 357646 142634
rect 357882 142398 357914 142634
rect 357294 106954 357914 142398
rect 357294 106718 357326 106954
rect 357562 106718 357646 106954
rect 357882 106718 357914 106954
rect 357294 106634 357914 106718
rect 357294 106398 357326 106634
rect 357562 106398 357646 106634
rect 357882 106398 357914 106634
rect 357294 70954 357914 106398
rect 357294 70718 357326 70954
rect 357562 70718 357646 70954
rect 357882 70718 357914 70954
rect 357294 70634 357914 70718
rect 357294 70398 357326 70634
rect 357562 70398 357646 70634
rect 357882 70398 357914 70634
rect 357294 34954 357914 70398
rect 357294 34718 357326 34954
rect 357562 34718 357646 34954
rect 357882 34718 357914 34954
rect 357294 34634 357914 34718
rect 357294 34398 357326 34634
rect 357562 34398 357646 34634
rect 357882 34398 357914 34634
rect 357294 -7066 357914 34398
rect 357294 -7302 357326 -7066
rect 357562 -7302 357646 -7066
rect 357882 -7302 357914 -7066
rect 357294 -7386 357914 -7302
rect 357294 -7622 357326 -7386
rect 357562 -7622 357646 -7386
rect 357882 -7622 357914 -7386
rect 357294 -7654 357914 -7622
rect 361794 704838 362414 711590
rect 361794 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 362414 704838
rect 361794 704518 362414 704602
rect 361794 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 362414 704518
rect 361794 687454 362414 704282
rect 361794 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 362414 687454
rect 361794 687134 362414 687218
rect 361794 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 362414 687134
rect 361794 651454 362414 686898
rect 361794 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 362414 651454
rect 361794 651134 362414 651218
rect 361794 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 362414 651134
rect 361794 615454 362414 650898
rect 361794 615218 361826 615454
rect 362062 615218 362146 615454
rect 362382 615218 362414 615454
rect 361794 615134 362414 615218
rect 361794 614898 361826 615134
rect 362062 614898 362146 615134
rect 362382 614898 362414 615134
rect 361794 579454 362414 614898
rect 361794 579218 361826 579454
rect 362062 579218 362146 579454
rect 362382 579218 362414 579454
rect 361794 579134 362414 579218
rect 361794 578898 361826 579134
rect 362062 578898 362146 579134
rect 362382 578898 362414 579134
rect 361794 543454 362414 578898
rect 361794 543218 361826 543454
rect 362062 543218 362146 543454
rect 362382 543218 362414 543454
rect 361794 543134 362414 543218
rect 361794 542898 361826 543134
rect 362062 542898 362146 543134
rect 362382 542898 362414 543134
rect 361794 507454 362414 542898
rect 361794 507218 361826 507454
rect 362062 507218 362146 507454
rect 362382 507218 362414 507454
rect 361794 507134 362414 507218
rect 361794 506898 361826 507134
rect 362062 506898 362146 507134
rect 362382 506898 362414 507134
rect 361794 471454 362414 506898
rect 361794 471218 361826 471454
rect 362062 471218 362146 471454
rect 362382 471218 362414 471454
rect 361794 471134 362414 471218
rect 361794 470898 361826 471134
rect 362062 470898 362146 471134
rect 362382 470898 362414 471134
rect 361794 435454 362414 470898
rect 361794 435218 361826 435454
rect 362062 435218 362146 435454
rect 362382 435218 362414 435454
rect 361794 435134 362414 435218
rect 361794 434898 361826 435134
rect 362062 434898 362146 435134
rect 362382 434898 362414 435134
rect 361794 399454 362414 434898
rect 361794 399218 361826 399454
rect 362062 399218 362146 399454
rect 362382 399218 362414 399454
rect 361794 399134 362414 399218
rect 361794 398898 361826 399134
rect 362062 398898 362146 399134
rect 362382 398898 362414 399134
rect 361794 363454 362414 398898
rect 361794 363218 361826 363454
rect 362062 363218 362146 363454
rect 362382 363218 362414 363454
rect 361794 363134 362414 363218
rect 361794 362898 361826 363134
rect 362062 362898 362146 363134
rect 362382 362898 362414 363134
rect 361794 327454 362414 362898
rect 361794 327218 361826 327454
rect 362062 327218 362146 327454
rect 362382 327218 362414 327454
rect 361794 327134 362414 327218
rect 361794 326898 361826 327134
rect 362062 326898 362146 327134
rect 362382 326898 362414 327134
rect 361794 291454 362414 326898
rect 361794 291218 361826 291454
rect 362062 291218 362146 291454
rect 362382 291218 362414 291454
rect 361794 291134 362414 291218
rect 361794 290898 361826 291134
rect 362062 290898 362146 291134
rect 362382 290898 362414 291134
rect 361794 255454 362414 290898
rect 361794 255218 361826 255454
rect 362062 255218 362146 255454
rect 362382 255218 362414 255454
rect 361794 255134 362414 255218
rect 361794 254898 361826 255134
rect 362062 254898 362146 255134
rect 362382 254898 362414 255134
rect 361794 219454 362414 254898
rect 361794 219218 361826 219454
rect 362062 219218 362146 219454
rect 362382 219218 362414 219454
rect 361794 219134 362414 219218
rect 361794 218898 361826 219134
rect 362062 218898 362146 219134
rect 362382 218898 362414 219134
rect 361794 183454 362414 218898
rect 361794 183218 361826 183454
rect 362062 183218 362146 183454
rect 362382 183218 362414 183454
rect 361794 183134 362414 183218
rect 361794 182898 361826 183134
rect 362062 182898 362146 183134
rect 362382 182898 362414 183134
rect 361794 147454 362414 182898
rect 361794 147218 361826 147454
rect 362062 147218 362146 147454
rect 362382 147218 362414 147454
rect 361794 147134 362414 147218
rect 361794 146898 361826 147134
rect 362062 146898 362146 147134
rect 362382 146898 362414 147134
rect 361794 111454 362414 146898
rect 361794 111218 361826 111454
rect 362062 111218 362146 111454
rect 362382 111218 362414 111454
rect 361794 111134 362414 111218
rect 361794 110898 361826 111134
rect 362062 110898 362146 111134
rect 362382 110898 362414 111134
rect 361794 75454 362414 110898
rect 361794 75218 361826 75454
rect 362062 75218 362146 75454
rect 362382 75218 362414 75454
rect 361794 75134 362414 75218
rect 361794 74898 361826 75134
rect 362062 74898 362146 75134
rect 362382 74898 362414 75134
rect 361794 39454 362414 74898
rect 361794 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 362414 39454
rect 361794 39134 362414 39218
rect 361794 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 362414 39134
rect 361794 3454 362414 38898
rect 361794 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 362414 3454
rect 361794 3134 362414 3218
rect 361794 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 362414 3134
rect 361794 -346 362414 2898
rect 361794 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 362414 -346
rect 361794 -666 362414 -582
rect 361794 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 362414 -666
rect 361794 -7654 362414 -902
rect 366294 705798 366914 711590
rect 366294 705562 366326 705798
rect 366562 705562 366646 705798
rect 366882 705562 366914 705798
rect 366294 705478 366914 705562
rect 366294 705242 366326 705478
rect 366562 705242 366646 705478
rect 366882 705242 366914 705478
rect 366294 691954 366914 705242
rect 366294 691718 366326 691954
rect 366562 691718 366646 691954
rect 366882 691718 366914 691954
rect 366294 691634 366914 691718
rect 366294 691398 366326 691634
rect 366562 691398 366646 691634
rect 366882 691398 366914 691634
rect 366294 655954 366914 691398
rect 366294 655718 366326 655954
rect 366562 655718 366646 655954
rect 366882 655718 366914 655954
rect 366294 655634 366914 655718
rect 366294 655398 366326 655634
rect 366562 655398 366646 655634
rect 366882 655398 366914 655634
rect 366294 619954 366914 655398
rect 366294 619718 366326 619954
rect 366562 619718 366646 619954
rect 366882 619718 366914 619954
rect 366294 619634 366914 619718
rect 366294 619398 366326 619634
rect 366562 619398 366646 619634
rect 366882 619398 366914 619634
rect 366294 583954 366914 619398
rect 366294 583718 366326 583954
rect 366562 583718 366646 583954
rect 366882 583718 366914 583954
rect 366294 583634 366914 583718
rect 366294 583398 366326 583634
rect 366562 583398 366646 583634
rect 366882 583398 366914 583634
rect 366294 547954 366914 583398
rect 366294 547718 366326 547954
rect 366562 547718 366646 547954
rect 366882 547718 366914 547954
rect 366294 547634 366914 547718
rect 366294 547398 366326 547634
rect 366562 547398 366646 547634
rect 366882 547398 366914 547634
rect 366294 511954 366914 547398
rect 366294 511718 366326 511954
rect 366562 511718 366646 511954
rect 366882 511718 366914 511954
rect 366294 511634 366914 511718
rect 366294 511398 366326 511634
rect 366562 511398 366646 511634
rect 366882 511398 366914 511634
rect 366294 475954 366914 511398
rect 366294 475718 366326 475954
rect 366562 475718 366646 475954
rect 366882 475718 366914 475954
rect 366294 475634 366914 475718
rect 366294 475398 366326 475634
rect 366562 475398 366646 475634
rect 366882 475398 366914 475634
rect 366294 439954 366914 475398
rect 366294 439718 366326 439954
rect 366562 439718 366646 439954
rect 366882 439718 366914 439954
rect 366294 439634 366914 439718
rect 366294 439398 366326 439634
rect 366562 439398 366646 439634
rect 366882 439398 366914 439634
rect 366294 403954 366914 439398
rect 366294 403718 366326 403954
rect 366562 403718 366646 403954
rect 366882 403718 366914 403954
rect 366294 403634 366914 403718
rect 366294 403398 366326 403634
rect 366562 403398 366646 403634
rect 366882 403398 366914 403634
rect 366294 367954 366914 403398
rect 366294 367718 366326 367954
rect 366562 367718 366646 367954
rect 366882 367718 366914 367954
rect 366294 367634 366914 367718
rect 366294 367398 366326 367634
rect 366562 367398 366646 367634
rect 366882 367398 366914 367634
rect 366294 331954 366914 367398
rect 366294 331718 366326 331954
rect 366562 331718 366646 331954
rect 366882 331718 366914 331954
rect 366294 331634 366914 331718
rect 366294 331398 366326 331634
rect 366562 331398 366646 331634
rect 366882 331398 366914 331634
rect 366294 295954 366914 331398
rect 366294 295718 366326 295954
rect 366562 295718 366646 295954
rect 366882 295718 366914 295954
rect 366294 295634 366914 295718
rect 366294 295398 366326 295634
rect 366562 295398 366646 295634
rect 366882 295398 366914 295634
rect 366294 259954 366914 295398
rect 366294 259718 366326 259954
rect 366562 259718 366646 259954
rect 366882 259718 366914 259954
rect 366294 259634 366914 259718
rect 366294 259398 366326 259634
rect 366562 259398 366646 259634
rect 366882 259398 366914 259634
rect 366294 223954 366914 259398
rect 366294 223718 366326 223954
rect 366562 223718 366646 223954
rect 366882 223718 366914 223954
rect 366294 223634 366914 223718
rect 366294 223398 366326 223634
rect 366562 223398 366646 223634
rect 366882 223398 366914 223634
rect 366294 187954 366914 223398
rect 366294 187718 366326 187954
rect 366562 187718 366646 187954
rect 366882 187718 366914 187954
rect 366294 187634 366914 187718
rect 366294 187398 366326 187634
rect 366562 187398 366646 187634
rect 366882 187398 366914 187634
rect 366294 151954 366914 187398
rect 366294 151718 366326 151954
rect 366562 151718 366646 151954
rect 366882 151718 366914 151954
rect 366294 151634 366914 151718
rect 366294 151398 366326 151634
rect 366562 151398 366646 151634
rect 366882 151398 366914 151634
rect 366294 115954 366914 151398
rect 366294 115718 366326 115954
rect 366562 115718 366646 115954
rect 366882 115718 366914 115954
rect 366294 115634 366914 115718
rect 366294 115398 366326 115634
rect 366562 115398 366646 115634
rect 366882 115398 366914 115634
rect 366294 79954 366914 115398
rect 366294 79718 366326 79954
rect 366562 79718 366646 79954
rect 366882 79718 366914 79954
rect 366294 79634 366914 79718
rect 366294 79398 366326 79634
rect 366562 79398 366646 79634
rect 366882 79398 366914 79634
rect 366294 43954 366914 79398
rect 366294 43718 366326 43954
rect 366562 43718 366646 43954
rect 366882 43718 366914 43954
rect 366294 43634 366914 43718
rect 366294 43398 366326 43634
rect 366562 43398 366646 43634
rect 366882 43398 366914 43634
rect 366294 7954 366914 43398
rect 366294 7718 366326 7954
rect 366562 7718 366646 7954
rect 366882 7718 366914 7954
rect 366294 7634 366914 7718
rect 366294 7398 366326 7634
rect 366562 7398 366646 7634
rect 366882 7398 366914 7634
rect 366294 -1306 366914 7398
rect 366294 -1542 366326 -1306
rect 366562 -1542 366646 -1306
rect 366882 -1542 366914 -1306
rect 366294 -1626 366914 -1542
rect 366294 -1862 366326 -1626
rect 366562 -1862 366646 -1626
rect 366882 -1862 366914 -1626
rect 366294 -7654 366914 -1862
rect 370794 706758 371414 711590
rect 370794 706522 370826 706758
rect 371062 706522 371146 706758
rect 371382 706522 371414 706758
rect 370794 706438 371414 706522
rect 370794 706202 370826 706438
rect 371062 706202 371146 706438
rect 371382 706202 371414 706438
rect 370794 696454 371414 706202
rect 370794 696218 370826 696454
rect 371062 696218 371146 696454
rect 371382 696218 371414 696454
rect 370794 696134 371414 696218
rect 370794 695898 370826 696134
rect 371062 695898 371146 696134
rect 371382 695898 371414 696134
rect 370794 660454 371414 695898
rect 370794 660218 370826 660454
rect 371062 660218 371146 660454
rect 371382 660218 371414 660454
rect 370794 660134 371414 660218
rect 370794 659898 370826 660134
rect 371062 659898 371146 660134
rect 371382 659898 371414 660134
rect 370794 624454 371414 659898
rect 370794 624218 370826 624454
rect 371062 624218 371146 624454
rect 371382 624218 371414 624454
rect 370794 624134 371414 624218
rect 370794 623898 370826 624134
rect 371062 623898 371146 624134
rect 371382 623898 371414 624134
rect 370794 588454 371414 623898
rect 370794 588218 370826 588454
rect 371062 588218 371146 588454
rect 371382 588218 371414 588454
rect 370794 588134 371414 588218
rect 370794 587898 370826 588134
rect 371062 587898 371146 588134
rect 371382 587898 371414 588134
rect 370794 552454 371414 587898
rect 370794 552218 370826 552454
rect 371062 552218 371146 552454
rect 371382 552218 371414 552454
rect 370794 552134 371414 552218
rect 370794 551898 370826 552134
rect 371062 551898 371146 552134
rect 371382 551898 371414 552134
rect 370794 516454 371414 551898
rect 370794 516218 370826 516454
rect 371062 516218 371146 516454
rect 371382 516218 371414 516454
rect 370794 516134 371414 516218
rect 370794 515898 370826 516134
rect 371062 515898 371146 516134
rect 371382 515898 371414 516134
rect 370794 480454 371414 515898
rect 370794 480218 370826 480454
rect 371062 480218 371146 480454
rect 371382 480218 371414 480454
rect 370794 480134 371414 480218
rect 370794 479898 370826 480134
rect 371062 479898 371146 480134
rect 371382 479898 371414 480134
rect 370794 444454 371414 479898
rect 370794 444218 370826 444454
rect 371062 444218 371146 444454
rect 371382 444218 371414 444454
rect 370794 444134 371414 444218
rect 370794 443898 370826 444134
rect 371062 443898 371146 444134
rect 371382 443898 371414 444134
rect 370794 408454 371414 443898
rect 370794 408218 370826 408454
rect 371062 408218 371146 408454
rect 371382 408218 371414 408454
rect 370794 408134 371414 408218
rect 370794 407898 370826 408134
rect 371062 407898 371146 408134
rect 371382 407898 371414 408134
rect 370794 372454 371414 407898
rect 370794 372218 370826 372454
rect 371062 372218 371146 372454
rect 371382 372218 371414 372454
rect 370794 372134 371414 372218
rect 370794 371898 370826 372134
rect 371062 371898 371146 372134
rect 371382 371898 371414 372134
rect 370794 336454 371414 371898
rect 370794 336218 370826 336454
rect 371062 336218 371146 336454
rect 371382 336218 371414 336454
rect 370794 336134 371414 336218
rect 370794 335898 370826 336134
rect 371062 335898 371146 336134
rect 371382 335898 371414 336134
rect 370794 300454 371414 335898
rect 370794 300218 370826 300454
rect 371062 300218 371146 300454
rect 371382 300218 371414 300454
rect 370794 300134 371414 300218
rect 370794 299898 370826 300134
rect 371062 299898 371146 300134
rect 371382 299898 371414 300134
rect 370794 264454 371414 299898
rect 370794 264218 370826 264454
rect 371062 264218 371146 264454
rect 371382 264218 371414 264454
rect 370794 264134 371414 264218
rect 370794 263898 370826 264134
rect 371062 263898 371146 264134
rect 371382 263898 371414 264134
rect 370794 228454 371414 263898
rect 370794 228218 370826 228454
rect 371062 228218 371146 228454
rect 371382 228218 371414 228454
rect 370794 228134 371414 228218
rect 370794 227898 370826 228134
rect 371062 227898 371146 228134
rect 371382 227898 371414 228134
rect 370794 192454 371414 227898
rect 370794 192218 370826 192454
rect 371062 192218 371146 192454
rect 371382 192218 371414 192454
rect 370794 192134 371414 192218
rect 370794 191898 370826 192134
rect 371062 191898 371146 192134
rect 371382 191898 371414 192134
rect 370794 156454 371414 191898
rect 370794 156218 370826 156454
rect 371062 156218 371146 156454
rect 371382 156218 371414 156454
rect 370794 156134 371414 156218
rect 370794 155898 370826 156134
rect 371062 155898 371146 156134
rect 371382 155898 371414 156134
rect 370794 120454 371414 155898
rect 370794 120218 370826 120454
rect 371062 120218 371146 120454
rect 371382 120218 371414 120454
rect 370794 120134 371414 120218
rect 370794 119898 370826 120134
rect 371062 119898 371146 120134
rect 371382 119898 371414 120134
rect 370794 84454 371414 119898
rect 370794 84218 370826 84454
rect 371062 84218 371146 84454
rect 371382 84218 371414 84454
rect 370794 84134 371414 84218
rect 370794 83898 370826 84134
rect 371062 83898 371146 84134
rect 371382 83898 371414 84134
rect 370794 48454 371414 83898
rect 370794 48218 370826 48454
rect 371062 48218 371146 48454
rect 371382 48218 371414 48454
rect 370794 48134 371414 48218
rect 370794 47898 370826 48134
rect 371062 47898 371146 48134
rect 371382 47898 371414 48134
rect 370794 12454 371414 47898
rect 370794 12218 370826 12454
rect 371062 12218 371146 12454
rect 371382 12218 371414 12454
rect 370794 12134 371414 12218
rect 370794 11898 370826 12134
rect 371062 11898 371146 12134
rect 371382 11898 371414 12134
rect 370794 -2266 371414 11898
rect 370794 -2502 370826 -2266
rect 371062 -2502 371146 -2266
rect 371382 -2502 371414 -2266
rect 370794 -2586 371414 -2502
rect 370794 -2822 370826 -2586
rect 371062 -2822 371146 -2586
rect 371382 -2822 371414 -2586
rect 370794 -7654 371414 -2822
rect 375294 707718 375914 711590
rect 375294 707482 375326 707718
rect 375562 707482 375646 707718
rect 375882 707482 375914 707718
rect 375294 707398 375914 707482
rect 375294 707162 375326 707398
rect 375562 707162 375646 707398
rect 375882 707162 375914 707398
rect 375294 700954 375914 707162
rect 375294 700718 375326 700954
rect 375562 700718 375646 700954
rect 375882 700718 375914 700954
rect 375294 700634 375914 700718
rect 375294 700398 375326 700634
rect 375562 700398 375646 700634
rect 375882 700398 375914 700634
rect 375294 664954 375914 700398
rect 375294 664718 375326 664954
rect 375562 664718 375646 664954
rect 375882 664718 375914 664954
rect 375294 664634 375914 664718
rect 375294 664398 375326 664634
rect 375562 664398 375646 664634
rect 375882 664398 375914 664634
rect 375294 628954 375914 664398
rect 375294 628718 375326 628954
rect 375562 628718 375646 628954
rect 375882 628718 375914 628954
rect 375294 628634 375914 628718
rect 375294 628398 375326 628634
rect 375562 628398 375646 628634
rect 375882 628398 375914 628634
rect 375294 592954 375914 628398
rect 375294 592718 375326 592954
rect 375562 592718 375646 592954
rect 375882 592718 375914 592954
rect 375294 592634 375914 592718
rect 375294 592398 375326 592634
rect 375562 592398 375646 592634
rect 375882 592398 375914 592634
rect 375294 556954 375914 592398
rect 375294 556718 375326 556954
rect 375562 556718 375646 556954
rect 375882 556718 375914 556954
rect 375294 556634 375914 556718
rect 375294 556398 375326 556634
rect 375562 556398 375646 556634
rect 375882 556398 375914 556634
rect 375294 520954 375914 556398
rect 375294 520718 375326 520954
rect 375562 520718 375646 520954
rect 375882 520718 375914 520954
rect 375294 520634 375914 520718
rect 375294 520398 375326 520634
rect 375562 520398 375646 520634
rect 375882 520398 375914 520634
rect 375294 484954 375914 520398
rect 375294 484718 375326 484954
rect 375562 484718 375646 484954
rect 375882 484718 375914 484954
rect 375294 484634 375914 484718
rect 375294 484398 375326 484634
rect 375562 484398 375646 484634
rect 375882 484398 375914 484634
rect 375294 448954 375914 484398
rect 375294 448718 375326 448954
rect 375562 448718 375646 448954
rect 375882 448718 375914 448954
rect 375294 448634 375914 448718
rect 375294 448398 375326 448634
rect 375562 448398 375646 448634
rect 375882 448398 375914 448634
rect 375294 412954 375914 448398
rect 375294 412718 375326 412954
rect 375562 412718 375646 412954
rect 375882 412718 375914 412954
rect 375294 412634 375914 412718
rect 375294 412398 375326 412634
rect 375562 412398 375646 412634
rect 375882 412398 375914 412634
rect 375294 376954 375914 412398
rect 375294 376718 375326 376954
rect 375562 376718 375646 376954
rect 375882 376718 375914 376954
rect 375294 376634 375914 376718
rect 375294 376398 375326 376634
rect 375562 376398 375646 376634
rect 375882 376398 375914 376634
rect 375294 340954 375914 376398
rect 375294 340718 375326 340954
rect 375562 340718 375646 340954
rect 375882 340718 375914 340954
rect 375294 340634 375914 340718
rect 375294 340398 375326 340634
rect 375562 340398 375646 340634
rect 375882 340398 375914 340634
rect 375294 304954 375914 340398
rect 375294 304718 375326 304954
rect 375562 304718 375646 304954
rect 375882 304718 375914 304954
rect 375294 304634 375914 304718
rect 375294 304398 375326 304634
rect 375562 304398 375646 304634
rect 375882 304398 375914 304634
rect 375294 268954 375914 304398
rect 375294 268718 375326 268954
rect 375562 268718 375646 268954
rect 375882 268718 375914 268954
rect 375294 268634 375914 268718
rect 375294 268398 375326 268634
rect 375562 268398 375646 268634
rect 375882 268398 375914 268634
rect 375294 232954 375914 268398
rect 375294 232718 375326 232954
rect 375562 232718 375646 232954
rect 375882 232718 375914 232954
rect 375294 232634 375914 232718
rect 375294 232398 375326 232634
rect 375562 232398 375646 232634
rect 375882 232398 375914 232634
rect 375294 196954 375914 232398
rect 375294 196718 375326 196954
rect 375562 196718 375646 196954
rect 375882 196718 375914 196954
rect 375294 196634 375914 196718
rect 375294 196398 375326 196634
rect 375562 196398 375646 196634
rect 375882 196398 375914 196634
rect 375294 160954 375914 196398
rect 375294 160718 375326 160954
rect 375562 160718 375646 160954
rect 375882 160718 375914 160954
rect 375294 160634 375914 160718
rect 375294 160398 375326 160634
rect 375562 160398 375646 160634
rect 375882 160398 375914 160634
rect 375294 124954 375914 160398
rect 375294 124718 375326 124954
rect 375562 124718 375646 124954
rect 375882 124718 375914 124954
rect 375294 124634 375914 124718
rect 375294 124398 375326 124634
rect 375562 124398 375646 124634
rect 375882 124398 375914 124634
rect 375294 88954 375914 124398
rect 375294 88718 375326 88954
rect 375562 88718 375646 88954
rect 375882 88718 375914 88954
rect 375294 88634 375914 88718
rect 375294 88398 375326 88634
rect 375562 88398 375646 88634
rect 375882 88398 375914 88634
rect 375294 52954 375914 88398
rect 375294 52718 375326 52954
rect 375562 52718 375646 52954
rect 375882 52718 375914 52954
rect 375294 52634 375914 52718
rect 375294 52398 375326 52634
rect 375562 52398 375646 52634
rect 375882 52398 375914 52634
rect 375294 16954 375914 52398
rect 375294 16718 375326 16954
rect 375562 16718 375646 16954
rect 375882 16718 375914 16954
rect 375294 16634 375914 16718
rect 375294 16398 375326 16634
rect 375562 16398 375646 16634
rect 375882 16398 375914 16634
rect 375294 -3226 375914 16398
rect 375294 -3462 375326 -3226
rect 375562 -3462 375646 -3226
rect 375882 -3462 375914 -3226
rect 375294 -3546 375914 -3462
rect 375294 -3782 375326 -3546
rect 375562 -3782 375646 -3546
rect 375882 -3782 375914 -3546
rect 375294 -7654 375914 -3782
rect 379794 708678 380414 711590
rect 379794 708442 379826 708678
rect 380062 708442 380146 708678
rect 380382 708442 380414 708678
rect 379794 708358 380414 708442
rect 379794 708122 379826 708358
rect 380062 708122 380146 708358
rect 380382 708122 380414 708358
rect 379794 669454 380414 708122
rect 379794 669218 379826 669454
rect 380062 669218 380146 669454
rect 380382 669218 380414 669454
rect 379794 669134 380414 669218
rect 379794 668898 379826 669134
rect 380062 668898 380146 669134
rect 380382 668898 380414 669134
rect 379794 633454 380414 668898
rect 379794 633218 379826 633454
rect 380062 633218 380146 633454
rect 380382 633218 380414 633454
rect 379794 633134 380414 633218
rect 379794 632898 379826 633134
rect 380062 632898 380146 633134
rect 380382 632898 380414 633134
rect 379794 597454 380414 632898
rect 379794 597218 379826 597454
rect 380062 597218 380146 597454
rect 380382 597218 380414 597454
rect 379794 597134 380414 597218
rect 379794 596898 379826 597134
rect 380062 596898 380146 597134
rect 380382 596898 380414 597134
rect 379794 561454 380414 596898
rect 379794 561218 379826 561454
rect 380062 561218 380146 561454
rect 380382 561218 380414 561454
rect 379794 561134 380414 561218
rect 379794 560898 379826 561134
rect 380062 560898 380146 561134
rect 380382 560898 380414 561134
rect 379794 525454 380414 560898
rect 379794 525218 379826 525454
rect 380062 525218 380146 525454
rect 380382 525218 380414 525454
rect 379794 525134 380414 525218
rect 379794 524898 379826 525134
rect 380062 524898 380146 525134
rect 380382 524898 380414 525134
rect 379794 489454 380414 524898
rect 379794 489218 379826 489454
rect 380062 489218 380146 489454
rect 380382 489218 380414 489454
rect 379794 489134 380414 489218
rect 379794 488898 379826 489134
rect 380062 488898 380146 489134
rect 380382 488898 380414 489134
rect 379794 453454 380414 488898
rect 379794 453218 379826 453454
rect 380062 453218 380146 453454
rect 380382 453218 380414 453454
rect 379794 453134 380414 453218
rect 379794 452898 379826 453134
rect 380062 452898 380146 453134
rect 380382 452898 380414 453134
rect 379794 417454 380414 452898
rect 379794 417218 379826 417454
rect 380062 417218 380146 417454
rect 380382 417218 380414 417454
rect 379794 417134 380414 417218
rect 379794 416898 379826 417134
rect 380062 416898 380146 417134
rect 380382 416898 380414 417134
rect 379794 381454 380414 416898
rect 379794 381218 379826 381454
rect 380062 381218 380146 381454
rect 380382 381218 380414 381454
rect 379794 381134 380414 381218
rect 379794 380898 379826 381134
rect 380062 380898 380146 381134
rect 380382 380898 380414 381134
rect 379794 345454 380414 380898
rect 379794 345218 379826 345454
rect 380062 345218 380146 345454
rect 380382 345218 380414 345454
rect 379794 345134 380414 345218
rect 379794 344898 379826 345134
rect 380062 344898 380146 345134
rect 380382 344898 380414 345134
rect 379794 309454 380414 344898
rect 379794 309218 379826 309454
rect 380062 309218 380146 309454
rect 380382 309218 380414 309454
rect 379794 309134 380414 309218
rect 379794 308898 379826 309134
rect 380062 308898 380146 309134
rect 380382 308898 380414 309134
rect 379794 273454 380414 308898
rect 379794 273218 379826 273454
rect 380062 273218 380146 273454
rect 380382 273218 380414 273454
rect 379794 273134 380414 273218
rect 379794 272898 379826 273134
rect 380062 272898 380146 273134
rect 380382 272898 380414 273134
rect 379794 237454 380414 272898
rect 379794 237218 379826 237454
rect 380062 237218 380146 237454
rect 380382 237218 380414 237454
rect 379794 237134 380414 237218
rect 379794 236898 379826 237134
rect 380062 236898 380146 237134
rect 380382 236898 380414 237134
rect 379794 201454 380414 236898
rect 379794 201218 379826 201454
rect 380062 201218 380146 201454
rect 380382 201218 380414 201454
rect 379794 201134 380414 201218
rect 379794 200898 379826 201134
rect 380062 200898 380146 201134
rect 380382 200898 380414 201134
rect 379794 165454 380414 200898
rect 379794 165218 379826 165454
rect 380062 165218 380146 165454
rect 380382 165218 380414 165454
rect 379794 165134 380414 165218
rect 379794 164898 379826 165134
rect 380062 164898 380146 165134
rect 380382 164898 380414 165134
rect 379794 129454 380414 164898
rect 379794 129218 379826 129454
rect 380062 129218 380146 129454
rect 380382 129218 380414 129454
rect 379794 129134 380414 129218
rect 379794 128898 379826 129134
rect 380062 128898 380146 129134
rect 380382 128898 380414 129134
rect 379794 93454 380414 128898
rect 379794 93218 379826 93454
rect 380062 93218 380146 93454
rect 380382 93218 380414 93454
rect 379794 93134 380414 93218
rect 379794 92898 379826 93134
rect 380062 92898 380146 93134
rect 380382 92898 380414 93134
rect 379794 57454 380414 92898
rect 379794 57218 379826 57454
rect 380062 57218 380146 57454
rect 380382 57218 380414 57454
rect 379794 57134 380414 57218
rect 379794 56898 379826 57134
rect 380062 56898 380146 57134
rect 380382 56898 380414 57134
rect 379794 21454 380414 56898
rect 379794 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 380414 21454
rect 379794 21134 380414 21218
rect 379794 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 380414 21134
rect 379794 -4186 380414 20898
rect 379794 -4422 379826 -4186
rect 380062 -4422 380146 -4186
rect 380382 -4422 380414 -4186
rect 379794 -4506 380414 -4422
rect 379794 -4742 379826 -4506
rect 380062 -4742 380146 -4506
rect 380382 -4742 380414 -4506
rect 379794 -7654 380414 -4742
rect 384294 709638 384914 711590
rect 384294 709402 384326 709638
rect 384562 709402 384646 709638
rect 384882 709402 384914 709638
rect 384294 709318 384914 709402
rect 384294 709082 384326 709318
rect 384562 709082 384646 709318
rect 384882 709082 384914 709318
rect 384294 673954 384914 709082
rect 384294 673718 384326 673954
rect 384562 673718 384646 673954
rect 384882 673718 384914 673954
rect 384294 673634 384914 673718
rect 384294 673398 384326 673634
rect 384562 673398 384646 673634
rect 384882 673398 384914 673634
rect 384294 637954 384914 673398
rect 384294 637718 384326 637954
rect 384562 637718 384646 637954
rect 384882 637718 384914 637954
rect 384294 637634 384914 637718
rect 384294 637398 384326 637634
rect 384562 637398 384646 637634
rect 384882 637398 384914 637634
rect 384294 601954 384914 637398
rect 384294 601718 384326 601954
rect 384562 601718 384646 601954
rect 384882 601718 384914 601954
rect 384294 601634 384914 601718
rect 384294 601398 384326 601634
rect 384562 601398 384646 601634
rect 384882 601398 384914 601634
rect 384294 565954 384914 601398
rect 384294 565718 384326 565954
rect 384562 565718 384646 565954
rect 384882 565718 384914 565954
rect 384294 565634 384914 565718
rect 384294 565398 384326 565634
rect 384562 565398 384646 565634
rect 384882 565398 384914 565634
rect 384294 529954 384914 565398
rect 384294 529718 384326 529954
rect 384562 529718 384646 529954
rect 384882 529718 384914 529954
rect 384294 529634 384914 529718
rect 384294 529398 384326 529634
rect 384562 529398 384646 529634
rect 384882 529398 384914 529634
rect 384294 493954 384914 529398
rect 384294 493718 384326 493954
rect 384562 493718 384646 493954
rect 384882 493718 384914 493954
rect 384294 493634 384914 493718
rect 384294 493398 384326 493634
rect 384562 493398 384646 493634
rect 384882 493398 384914 493634
rect 384294 457954 384914 493398
rect 384294 457718 384326 457954
rect 384562 457718 384646 457954
rect 384882 457718 384914 457954
rect 384294 457634 384914 457718
rect 384294 457398 384326 457634
rect 384562 457398 384646 457634
rect 384882 457398 384914 457634
rect 384294 421954 384914 457398
rect 384294 421718 384326 421954
rect 384562 421718 384646 421954
rect 384882 421718 384914 421954
rect 384294 421634 384914 421718
rect 384294 421398 384326 421634
rect 384562 421398 384646 421634
rect 384882 421398 384914 421634
rect 384294 385954 384914 421398
rect 384294 385718 384326 385954
rect 384562 385718 384646 385954
rect 384882 385718 384914 385954
rect 384294 385634 384914 385718
rect 384294 385398 384326 385634
rect 384562 385398 384646 385634
rect 384882 385398 384914 385634
rect 384294 349954 384914 385398
rect 384294 349718 384326 349954
rect 384562 349718 384646 349954
rect 384882 349718 384914 349954
rect 384294 349634 384914 349718
rect 384294 349398 384326 349634
rect 384562 349398 384646 349634
rect 384882 349398 384914 349634
rect 384294 313954 384914 349398
rect 384294 313718 384326 313954
rect 384562 313718 384646 313954
rect 384882 313718 384914 313954
rect 384294 313634 384914 313718
rect 384294 313398 384326 313634
rect 384562 313398 384646 313634
rect 384882 313398 384914 313634
rect 384294 277954 384914 313398
rect 384294 277718 384326 277954
rect 384562 277718 384646 277954
rect 384882 277718 384914 277954
rect 384294 277634 384914 277718
rect 384294 277398 384326 277634
rect 384562 277398 384646 277634
rect 384882 277398 384914 277634
rect 384294 241954 384914 277398
rect 384294 241718 384326 241954
rect 384562 241718 384646 241954
rect 384882 241718 384914 241954
rect 384294 241634 384914 241718
rect 384294 241398 384326 241634
rect 384562 241398 384646 241634
rect 384882 241398 384914 241634
rect 384294 205954 384914 241398
rect 384294 205718 384326 205954
rect 384562 205718 384646 205954
rect 384882 205718 384914 205954
rect 384294 205634 384914 205718
rect 384294 205398 384326 205634
rect 384562 205398 384646 205634
rect 384882 205398 384914 205634
rect 384294 169954 384914 205398
rect 384294 169718 384326 169954
rect 384562 169718 384646 169954
rect 384882 169718 384914 169954
rect 384294 169634 384914 169718
rect 384294 169398 384326 169634
rect 384562 169398 384646 169634
rect 384882 169398 384914 169634
rect 384294 133954 384914 169398
rect 384294 133718 384326 133954
rect 384562 133718 384646 133954
rect 384882 133718 384914 133954
rect 384294 133634 384914 133718
rect 384294 133398 384326 133634
rect 384562 133398 384646 133634
rect 384882 133398 384914 133634
rect 384294 97954 384914 133398
rect 384294 97718 384326 97954
rect 384562 97718 384646 97954
rect 384882 97718 384914 97954
rect 384294 97634 384914 97718
rect 384294 97398 384326 97634
rect 384562 97398 384646 97634
rect 384882 97398 384914 97634
rect 384294 61954 384914 97398
rect 384294 61718 384326 61954
rect 384562 61718 384646 61954
rect 384882 61718 384914 61954
rect 384294 61634 384914 61718
rect 384294 61398 384326 61634
rect 384562 61398 384646 61634
rect 384882 61398 384914 61634
rect 384294 25954 384914 61398
rect 384294 25718 384326 25954
rect 384562 25718 384646 25954
rect 384882 25718 384914 25954
rect 384294 25634 384914 25718
rect 384294 25398 384326 25634
rect 384562 25398 384646 25634
rect 384882 25398 384914 25634
rect 384294 -5146 384914 25398
rect 384294 -5382 384326 -5146
rect 384562 -5382 384646 -5146
rect 384882 -5382 384914 -5146
rect 384294 -5466 384914 -5382
rect 384294 -5702 384326 -5466
rect 384562 -5702 384646 -5466
rect 384882 -5702 384914 -5466
rect 384294 -7654 384914 -5702
rect 388794 710598 389414 711590
rect 388794 710362 388826 710598
rect 389062 710362 389146 710598
rect 389382 710362 389414 710598
rect 388794 710278 389414 710362
rect 388794 710042 388826 710278
rect 389062 710042 389146 710278
rect 389382 710042 389414 710278
rect 388794 678454 389414 710042
rect 388794 678218 388826 678454
rect 389062 678218 389146 678454
rect 389382 678218 389414 678454
rect 388794 678134 389414 678218
rect 388794 677898 388826 678134
rect 389062 677898 389146 678134
rect 389382 677898 389414 678134
rect 388794 642454 389414 677898
rect 388794 642218 388826 642454
rect 389062 642218 389146 642454
rect 389382 642218 389414 642454
rect 388794 642134 389414 642218
rect 388794 641898 388826 642134
rect 389062 641898 389146 642134
rect 389382 641898 389414 642134
rect 388794 606454 389414 641898
rect 388794 606218 388826 606454
rect 389062 606218 389146 606454
rect 389382 606218 389414 606454
rect 388794 606134 389414 606218
rect 388794 605898 388826 606134
rect 389062 605898 389146 606134
rect 389382 605898 389414 606134
rect 388794 570454 389414 605898
rect 388794 570218 388826 570454
rect 389062 570218 389146 570454
rect 389382 570218 389414 570454
rect 388794 570134 389414 570218
rect 388794 569898 388826 570134
rect 389062 569898 389146 570134
rect 389382 569898 389414 570134
rect 388794 534454 389414 569898
rect 388794 534218 388826 534454
rect 389062 534218 389146 534454
rect 389382 534218 389414 534454
rect 388794 534134 389414 534218
rect 388794 533898 388826 534134
rect 389062 533898 389146 534134
rect 389382 533898 389414 534134
rect 388794 498454 389414 533898
rect 388794 498218 388826 498454
rect 389062 498218 389146 498454
rect 389382 498218 389414 498454
rect 388794 498134 389414 498218
rect 388794 497898 388826 498134
rect 389062 497898 389146 498134
rect 389382 497898 389414 498134
rect 388794 462454 389414 497898
rect 388794 462218 388826 462454
rect 389062 462218 389146 462454
rect 389382 462218 389414 462454
rect 388794 462134 389414 462218
rect 388794 461898 388826 462134
rect 389062 461898 389146 462134
rect 389382 461898 389414 462134
rect 388794 426454 389414 461898
rect 388794 426218 388826 426454
rect 389062 426218 389146 426454
rect 389382 426218 389414 426454
rect 388794 426134 389414 426218
rect 388794 425898 388826 426134
rect 389062 425898 389146 426134
rect 389382 425898 389414 426134
rect 388794 390454 389414 425898
rect 388794 390218 388826 390454
rect 389062 390218 389146 390454
rect 389382 390218 389414 390454
rect 388794 390134 389414 390218
rect 388794 389898 388826 390134
rect 389062 389898 389146 390134
rect 389382 389898 389414 390134
rect 388794 354454 389414 389898
rect 388794 354218 388826 354454
rect 389062 354218 389146 354454
rect 389382 354218 389414 354454
rect 388794 354134 389414 354218
rect 388794 353898 388826 354134
rect 389062 353898 389146 354134
rect 389382 353898 389414 354134
rect 388794 318454 389414 353898
rect 388794 318218 388826 318454
rect 389062 318218 389146 318454
rect 389382 318218 389414 318454
rect 388794 318134 389414 318218
rect 388794 317898 388826 318134
rect 389062 317898 389146 318134
rect 389382 317898 389414 318134
rect 388794 282454 389414 317898
rect 388794 282218 388826 282454
rect 389062 282218 389146 282454
rect 389382 282218 389414 282454
rect 388794 282134 389414 282218
rect 388794 281898 388826 282134
rect 389062 281898 389146 282134
rect 389382 281898 389414 282134
rect 388794 246454 389414 281898
rect 388794 246218 388826 246454
rect 389062 246218 389146 246454
rect 389382 246218 389414 246454
rect 388794 246134 389414 246218
rect 388794 245898 388826 246134
rect 389062 245898 389146 246134
rect 389382 245898 389414 246134
rect 388794 210454 389414 245898
rect 388794 210218 388826 210454
rect 389062 210218 389146 210454
rect 389382 210218 389414 210454
rect 388794 210134 389414 210218
rect 388794 209898 388826 210134
rect 389062 209898 389146 210134
rect 389382 209898 389414 210134
rect 388794 174454 389414 209898
rect 388794 174218 388826 174454
rect 389062 174218 389146 174454
rect 389382 174218 389414 174454
rect 388794 174134 389414 174218
rect 388794 173898 388826 174134
rect 389062 173898 389146 174134
rect 389382 173898 389414 174134
rect 388794 138454 389414 173898
rect 388794 138218 388826 138454
rect 389062 138218 389146 138454
rect 389382 138218 389414 138454
rect 388794 138134 389414 138218
rect 388794 137898 388826 138134
rect 389062 137898 389146 138134
rect 389382 137898 389414 138134
rect 388794 102454 389414 137898
rect 388794 102218 388826 102454
rect 389062 102218 389146 102454
rect 389382 102218 389414 102454
rect 388794 102134 389414 102218
rect 388794 101898 388826 102134
rect 389062 101898 389146 102134
rect 389382 101898 389414 102134
rect 388794 66454 389414 101898
rect 388794 66218 388826 66454
rect 389062 66218 389146 66454
rect 389382 66218 389414 66454
rect 388794 66134 389414 66218
rect 388794 65898 388826 66134
rect 389062 65898 389146 66134
rect 389382 65898 389414 66134
rect 388794 30454 389414 65898
rect 388794 30218 388826 30454
rect 389062 30218 389146 30454
rect 389382 30218 389414 30454
rect 388794 30134 389414 30218
rect 388794 29898 388826 30134
rect 389062 29898 389146 30134
rect 389382 29898 389414 30134
rect 388794 -6106 389414 29898
rect 388794 -6342 388826 -6106
rect 389062 -6342 389146 -6106
rect 389382 -6342 389414 -6106
rect 388794 -6426 389414 -6342
rect 388794 -6662 388826 -6426
rect 389062 -6662 389146 -6426
rect 389382 -6662 389414 -6426
rect 388794 -7654 389414 -6662
rect 393294 711558 393914 711590
rect 393294 711322 393326 711558
rect 393562 711322 393646 711558
rect 393882 711322 393914 711558
rect 393294 711238 393914 711322
rect 393294 711002 393326 711238
rect 393562 711002 393646 711238
rect 393882 711002 393914 711238
rect 393294 682954 393914 711002
rect 393294 682718 393326 682954
rect 393562 682718 393646 682954
rect 393882 682718 393914 682954
rect 393294 682634 393914 682718
rect 393294 682398 393326 682634
rect 393562 682398 393646 682634
rect 393882 682398 393914 682634
rect 393294 646954 393914 682398
rect 393294 646718 393326 646954
rect 393562 646718 393646 646954
rect 393882 646718 393914 646954
rect 393294 646634 393914 646718
rect 393294 646398 393326 646634
rect 393562 646398 393646 646634
rect 393882 646398 393914 646634
rect 393294 610954 393914 646398
rect 393294 610718 393326 610954
rect 393562 610718 393646 610954
rect 393882 610718 393914 610954
rect 393294 610634 393914 610718
rect 393294 610398 393326 610634
rect 393562 610398 393646 610634
rect 393882 610398 393914 610634
rect 393294 574954 393914 610398
rect 393294 574718 393326 574954
rect 393562 574718 393646 574954
rect 393882 574718 393914 574954
rect 393294 574634 393914 574718
rect 393294 574398 393326 574634
rect 393562 574398 393646 574634
rect 393882 574398 393914 574634
rect 393294 538954 393914 574398
rect 393294 538718 393326 538954
rect 393562 538718 393646 538954
rect 393882 538718 393914 538954
rect 393294 538634 393914 538718
rect 393294 538398 393326 538634
rect 393562 538398 393646 538634
rect 393882 538398 393914 538634
rect 393294 502954 393914 538398
rect 393294 502718 393326 502954
rect 393562 502718 393646 502954
rect 393882 502718 393914 502954
rect 393294 502634 393914 502718
rect 393294 502398 393326 502634
rect 393562 502398 393646 502634
rect 393882 502398 393914 502634
rect 393294 466954 393914 502398
rect 393294 466718 393326 466954
rect 393562 466718 393646 466954
rect 393882 466718 393914 466954
rect 393294 466634 393914 466718
rect 393294 466398 393326 466634
rect 393562 466398 393646 466634
rect 393882 466398 393914 466634
rect 393294 430954 393914 466398
rect 393294 430718 393326 430954
rect 393562 430718 393646 430954
rect 393882 430718 393914 430954
rect 393294 430634 393914 430718
rect 393294 430398 393326 430634
rect 393562 430398 393646 430634
rect 393882 430398 393914 430634
rect 393294 394954 393914 430398
rect 393294 394718 393326 394954
rect 393562 394718 393646 394954
rect 393882 394718 393914 394954
rect 393294 394634 393914 394718
rect 393294 394398 393326 394634
rect 393562 394398 393646 394634
rect 393882 394398 393914 394634
rect 393294 358954 393914 394398
rect 393294 358718 393326 358954
rect 393562 358718 393646 358954
rect 393882 358718 393914 358954
rect 393294 358634 393914 358718
rect 393294 358398 393326 358634
rect 393562 358398 393646 358634
rect 393882 358398 393914 358634
rect 393294 322954 393914 358398
rect 393294 322718 393326 322954
rect 393562 322718 393646 322954
rect 393882 322718 393914 322954
rect 393294 322634 393914 322718
rect 393294 322398 393326 322634
rect 393562 322398 393646 322634
rect 393882 322398 393914 322634
rect 393294 286954 393914 322398
rect 393294 286718 393326 286954
rect 393562 286718 393646 286954
rect 393882 286718 393914 286954
rect 393294 286634 393914 286718
rect 393294 286398 393326 286634
rect 393562 286398 393646 286634
rect 393882 286398 393914 286634
rect 393294 250954 393914 286398
rect 393294 250718 393326 250954
rect 393562 250718 393646 250954
rect 393882 250718 393914 250954
rect 393294 250634 393914 250718
rect 393294 250398 393326 250634
rect 393562 250398 393646 250634
rect 393882 250398 393914 250634
rect 393294 214954 393914 250398
rect 393294 214718 393326 214954
rect 393562 214718 393646 214954
rect 393882 214718 393914 214954
rect 393294 214634 393914 214718
rect 393294 214398 393326 214634
rect 393562 214398 393646 214634
rect 393882 214398 393914 214634
rect 393294 178954 393914 214398
rect 393294 178718 393326 178954
rect 393562 178718 393646 178954
rect 393882 178718 393914 178954
rect 393294 178634 393914 178718
rect 393294 178398 393326 178634
rect 393562 178398 393646 178634
rect 393882 178398 393914 178634
rect 393294 142954 393914 178398
rect 393294 142718 393326 142954
rect 393562 142718 393646 142954
rect 393882 142718 393914 142954
rect 393294 142634 393914 142718
rect 393294 142398 393326 142634
rect 393562 142398 393646 142634
rect 393882 142398 393914 142634
rect 393294 106954 393914 142398
rect 393294 106718 393326 106954
rect 393562 106718 393646 106954
rect 393882 106718 393914 106954
rect 393294 106634 393914 106718
rect 393294 106398 393326 106634
rect 393562 106398 393646 106634
rect 393882 106398 393914 106634
rect 393294 70954 393914 106398
rect 393294 70718 393326 70954
rect 393562 70718 393646 70954
rect 393882 70718 393914 70954
rect 393294 70634 393914 70718
rect 393294 70398 393326 70634
rect 393562 70398 393646 70634
rect 393882 70398 393914 70634
rect 393294 34954 393914 70398
rect 393294 34718 393326 34954
rect 393562 34718 393646 34954
rect 393882 34718 393914 34954
rect 393294 34634 393914 34718
rect 393294 34398 393326 34634
rect 393562 34398 393646 34634
rect 393882 34398 393914 34634
rect 393294 -7066 393914 34398
rect 393294 -7302 393326 -7066
rect 393562 -7302 393646 -7066
rect 393882 -7302 393914 -7066
rect 393294 -7386 393914 -7302
rect 393294 -7622 393326 -7386
rect 393562 -7622 393646 -7386
rect 393882 -7622 393914 -7386
rect 393294 -7654 393914 -7622
rect 397794 704838 398414 711590
rect 397794 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 398414 704838
rect 397794 704518 398414 704602
rect 397794 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 398414 704518
rect 397794 687454 398414 704282
rect 397794 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 398414 687454
rect 397794 687134 398414 687218
rect 397794 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 398414 687134
rect 397794 651454 398414 686898
rect 397794 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 398414 651454
rect 397794 651134 398414 651218
rect 397794 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 398414 651134
rect 397794 615454 398414 650898
rect 397794 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 398414 615454
rect 397794 615134 398414 615218
rect 397794 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 398414 615134
rect 397794 579454 398414 614898
rect 397794 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 398414 579454
rect 397794 579134 398414 579218
rect 397794 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 398414 579134
rect 397794 543454 398414 578898
rect 397794 543218 397826 543454
rect 398062 543218 398146 543454
rect 398382 543218 398414 543454
rect 397794 543134 398414 543218
rect 397794 542898 397826 543134
rect 398062 542898 398146 543134
rect 398382 542898 398414 543134
rect 397794 507454 398414 542898
rect 397794 507218 397826 507454
rect 398062 507218 398146 507454
rect 398382 507218 398414 507454
rect 397794 507134 398414 507218
rect 397794 506898 397826 507134
rect 398062 506898 398146 507134
rect 398382 506898 398414 507134
rect 397794 471454 398414 506898
rect 397794 471218 397826 471454
rect 398062 471218 398146 471454
rect 398382 471218 398414 471454
rect 397794 471134 398414 471218
rect 397794 470898 397826 471134
rect 398062 470898 398146 471134
rect 398382 470898 398414 471134
rect 397794 435454 398414 470898
rect 397794 435218 397826 435454
rect 398062 435218 398146 435454
rect 398382 435218 398414 435454
rect 397794 435134 398414 435218
rect 397794 434898 397826 435134
rect 398062 434898 398146 435134
rect 398382 434898 398414 435134
rect 397794 399454 398414 434898
rect 397794 399218 397826 399454
rect 398062 399218 398146 399454
rect 398382 399218 398414 399454
rect 397794 399134 398414 399218
rect 397794 398898 397826 399134
rect 398062 398898 398146 399134
rect 398382 398898 398414 399134
rect 397794 363454 398414 398898
rect 397794 363218 397826 363454
rect 398062 363218 398146 363454
rect 398382 363218 398414 363454
rect 397794 363134 398414 363218
rect 397794 362898 397826 363134
rect 398062 362898 398146 363134
rect 398382 362898 398414 363134
rect 397794 327454 398414 362898
rect 397794 327218 397826 327454
rect 398062 327218 398146 327454
rect 398382 327218 398414 327454
rect 397794 327134 398414 327218
rect 397794 326898 397826 327134
rect 398062 326898 398146 327134
rect 398382 326898 398414 327134
rect 397794 291454 398414 326898
rect 397794 291218 397826 291454
rect 398062 291218 398146 291454
rect 398382 291218 398414 291454
rect 397794 291134 398414 291218
rect 397794 290898 397826 291134
rect 398062 290898 398146 291134
rect 398382 290898 398414 291134
rect 397794 255454 398414 290898
rect 397794 255218 397826 255454
rect 398062 255218 398146 255454
rect 398382 255218 398414 255454
rect 397794 255134 398414 255218
rect 397794 254898 397826 255134
rect 398062 254898 398146 255134
rect 398382 254898 398414 255134
rect 397794 219454 398414 254898
rect 397794 219218 397826 219454
rect 398062 219218 398146 219454
rect 398382 219218 398414 219454
rect 397794 219134 398414 219218
rect 397794 218898 397826 219134
rect 398062 218898 398146 219134
rect 398382 218898 398414 219134
rect 397794 183454 398414 218898
rect 397794 183218 397826 183454
rect 398062 183218 398146 183454
rect 398382 183218 398414 183454
rect 397794 183134 398414 183218
rect 397794 182898 397826 183134
rect 398062 182898 398146 183134
rect 398382 182898 398414 183134
rect 397794 147454 398414 182898
rect 397794 147218 397826 147454
rect 398062 147218 398146 147454
rect 398382 147218 398414 147454
rect 397794 147134 398414 147218
rect 397794 146898 397826 147134
rect 398062 146898 398146 147134
rect 398382 146898 398414 147134
rect 397794 111454 398414 146898
rect 397794 111218 397826 111454
rect 398062 111218 398146 111454
rect 398382 111218 398414 111454
rect 397794 111134 398414 111218
rect 397794 110898 397826 111134
rect 398062 110898 398146 111134
rect 398382 110898 398414 111134
rect 397794 75454 398414 110898
rect 397794 75218 397826 75454
rect 398062 75218 398146 75454
rect 398382 75218 398414 75454
rect 397794 75134 398414 75218
rect 397794 74898 397826 75134
rect 398062 74898 398146 75134
rect 398382 74898 398414 75134
rect 397794 39454 398414 74898
rect 397794 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 398414 39454
rect 397794 39134 398414 39218
rect 397794 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 398414 39134
rect 397794 3454 398414 38898
rect 397794 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 398414 3454
rect 397794 3134 398414 3218
rect 397794 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 398414 3134
rect 397794 -346 398414 2898
rect 397794 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 398414 -346
rect 397794 -666 398414 -582
rect 397794 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 398414 -666
rect 397794 -7654 398414 -902
rect 402294 705798 402914 711590
rect 402294 705562 402326 705798
rect 402562 705562 402646 705798
rect 402882 705562 402914 705798
rect 402294 705478 402914 705562
rect 402294 705242 402326 705478
rect 402562 705242 402646 705478
rect 402882 705242 402914 705478
rect 402294 691954 402914 705242
rect 402294 691718 402326 691954
rect 402562 691718 402646 691954
rect 402882 691718 402914 691954
rect 402294 691634 402914 691718
rect 402294 691398 402326 691634
rect 402562 691398 402646 691634
rect 402882 691398 402914 691634
rect 402294 655954 402914 691398
rect 402294 655718 402326 655954
rect 402562 655718 402646 655954
rect 402882 655718 402914 655954
rect 402294 655634 402914 655718
rect 402294 655398 402326 655634
rect 402562 655398 402646 655634
rect 402882 655398 402914 655634
rect 402294 619954 402914 655398
rect 402294 619718 402326 619954
rect 402562 619718 402646 619954
rect 402882 619718 402914 619954
rect 402294 619634 402914 619718
rect 402294 619398 402326 619634
rect 402562 619398 402646 619634
rect 402882 619398 402914 619634
rect 402294 583954 402914 619398
rect 402294 583718 402326 583954
rect 402562 583718 402646 583954
rect 402882 583718 402914 583954
rect 402294 583634 402914 583718
rect 402294 583398 402326 583634
rect 402562 583398 402646 583634
rect 402882 583398 402914 583634
rect 402294 547954 402914 583398
rect 402294 547718 402326 547954
rect 402562 547718 402646 547954
rect 402882 547718 402914 547954
rect 402294 547634 402914 547718
rect 402294 547398 402326 547634
rect 402562 547398 402646 547634
rect 402882 547398 402914 547634
rect 402294 511954 402914 547398
rect 402294 511718 402326 511954
rect 402562 511718 402646 511954
rect 402882 511718 402914 511954
rect 402294 511634 402914 511718
rect 402294 511398 402326 511634
rect 402562 511398 402646 511634
rect 402882 511398 402914 511634
rect 402294 475954 402914 511398
rect 402294 475718 402326 475954
rect 402562 475718 402646 475954
rect 402882 475718 402914 475954
rect 402294 475634 402914 475718
rect 402294 475398 402326 475634
rect 402562 475398 402646 475634
rect 402882 475398 402914 475634
rect 402294 439954 402914 475398
rect 402294 439718 402326 439954
rect 402562 439718 402646 439954
rect 402882 439718 402914 439954
rect 402294 439634 402914 439718
rect 402294 439398 402326 439634
rect 402562 439398 402646 439634
rect 402882 439398 402914 439634
rect 402294 403954 402914 439398
rect 402294 403718 402326 403954
rect 402562 403718 402646 403954
rect 402882 403718 402914 403954
rect 402294 403634 402914 403718
rect 402294 403398 402326 403634
rect 402562 403398 402646 403634
rect 402882 403398 402914 403634
rect 402294 367954 402914 403398
rect 402294 367718 402326 367954
rect 402562 367718 402646 367954
rect 402882 367718 402914 367954
rect 402294 367634 402914 367718
rect 402294 367398 402326 367634
rect 402562 367398 402646 367634
rect 402882 367398 402914 367634
rect 402294 331954 402914 367398
rect 402294 331718 402326 331954
rect 402562 331718 402646 331954
rect 402882 331718 402914 331954
rect 402294 331634 402914 331718
rect 402294 331398 402326 331634
rect 402562 331398 402646 331634
rect 402882 331398 402914 331634
rect 402294 295954 402914 331398
rect 402294 295718 402326 295954
rect 402562 295718 402646 295954
rect 402882 295718 402914 295954
rect 402294 295634 402914 295718
rect 402294 295398 402326 295634
rect 402562 295398 402646 295634
rect 402882 295398 402914 295634
rect 402294 259954 402914 295398
rect 402294 259718 402326 259954
rect 402562 259718 402646 259954
rect 402882 259718 402914 259954
rect 402294 259634 402914 259718
rect 402294 259398 402326 259634
rect 402562 259398 402646 259634
rect 402882 259398 402914 259634
rect 402294 223954 402914 259398
rect 402294 223718 402326 223954
rect 402562 223718 402646 223954
rect 402882 223718 402914 223954
rect 402294 223634 402914 223718
rect 402294 223398 402326 223634
rect 402562 223398 402646 223634
rect 402882 223398 402914 223634
rect 402294 187954 402914 223398
rect 402294 187718 402326 187954
rect 402562 187718 402646 187954
rect 402882 187718 402914 187954
rect 402294 187634 402914 187718
rect 402294 187398 402326 187634
rect 402562 187398 402646 187634
rect 402882 187398 402914 187634
rect 402294 151954 402914 187398
rect 402294 151718 402326 151954
rect 402562 151718 402646 151954
rect 402882 151718 402914 151954
rect 402294 151634 402914 151718
rect 402294 151398 402326 151634
rect 402562 151398 402646 151634
rect 402882 151398 402914 151634
rect 402294 115954 402914 151398
rect 402294 115718 402326 115954
rect 402562 115718 402646 115954
rect 402882 115718 402914 115954
rect 402294 115634 402914 115718
rect 402294 115398 402326 115634
rect 402562 115398 402646 115634
rect 402882 115398 402914 115634
rect 402294 79954 402914 115398
rect 402294 79718 402326 79954
rect 402562 79718 402646 79954
rect 402882 79718 402914 79954
rect 402294 79634 402914 79718
rect 402294 79398 402326 79634
rect 402562 79398 402646 79634
rect 402882 79398 402914 79634
rect 402294 43954 402914 79398
rect 402294 43718 402326 43954
rect 402562 43718 402646 43954
rect 402882 43718 402914 43954
rect 402294 43634 402914 43718
rect 402294 43398 402326 43634
rect 402562 43398 402646 43634
rect 402882 43398 402914 43634
rect 402294 7954 402914 43398
rect 402294 7718 402326 7954
rect 402562 7718 402646 7954
rect 402882 7718 402914 7954
rect 402294 7634 402914 7718
rect 402294 7398 402326 7634
rect 402562 7398 402646 7634
rect 402882 7398 402914 7634
rect 402294 -1306 402914 7398
rect 402294 -1542 402326 -1306
rect 402562 -1542 402646 -1306
rect 402882 -1542 402914 -1306
rect 402294 -1626 402914 -1542
rect 402294 -1862 402326 -1626
rect 402562 -1862 402646 -1626
rect 402882 -1862 402914 -1626
rect 402294 -7654 402914 -1862
rect 406794 706758 407414 711590
rect 406794 706522 406826 706758
rect 407062 706522 407146 706758
rect 407382 706522 407414 706758
rect 406794 706438 407414 706522
rect 406794 706202 406826 706438
rect 407062 706202 407146 706438
rect 407382 706202 407414 706438
rect 406794 696454 407414 706202
rect 406794 696218 406826 696454
rect 407062 696218 407146 696454
rect 407382 696218 407414 696454
rect 406794 696134 407414 696218
rect 406794 695898 406826 696134
rect 407062 695898 407146 696134
rect 407382 695898 407414 696134
rect 406794 660454 407414 695898
rect 406794 660218 406826 660454
rect 407062 660218 407146 660454
rect 407382 660218 407414 660454
rect 406794 660134 407414 660218
rect 406794 659898 406826 660134
rect 407062 659898 407146 660134
rect 407382 659898 407414 660134
rect 406794 624454 407414 659898
rect 406794 624218 406826 624454
rect 407062 624218 407146 624454
rect 407382 624218 407414 624454
rect 406794 624134 407414 624218
rect 406794 623898 406826 624134
rect 407062 623898 407146 624134
rect 407382 623898 407414 624134
rect 406794 588454 407414 623898
rect 406794 588218 406826 588454
rect 407062 588218 407146 588454
rect 407382 588218 407414 588454
rect 406794 588134 407414 588218
rect 406794 587898 406826 588134
rect 407062 587898 407146 588134
rect 407382 587898 407414 588134
rect 406794 552454 407414 587898
rect 406794 552218 406826 552454
rect 407062 552218 407146 552454
rect 407382 552218 407414 552454
rect 406794 552134 407414 552218
rect 406794 551898 406826 552134
rect 407062 551898 407146 552134
rect 407382 551898 407414 552134
rect 406794 516454 407414 551898
rect 406794 516218 406826 516454
rect 407062 516218 407146 516454
rect 407382 516218 407414 516454
rect 406794 516134 407414 516218
rect 406794 515898 406826 516134
rect 407062 515898 407146 516134
rect 407382 515898 407414 516134
rect 406794 480454 407414 515898
rect 406794 480218 406826 480454
rect 407062 480218 407146 480454
rect 407382 480218 407414 480454
rect 406794 480134 407414 480218
rect 406794 479898 406826 480134
rect 407062 479898 407146 480134
rect 407382 479898 407414 480134
rect 406794 444454 407414 479898
rect 406794 444218 406826 444454
rect 407062 444218 407146 444454
rect 407382 444218 407414 444454
rect 406794 444134 407414 444218
rect 406794 443898 406826 444134
rect 407062 443898 407146 444134
rect 407382 443898 407414 444134
rect 406794 408454 407414 443898
rect 406794 408218 406826 408454
rect 407062 408218 407146 408454
rect 407382 408218 407414 408454
rect 406794 408134 407414 408218
rect 406794 407898 406826 408134
rect 407062 407898 407146 408134
rect 407382 407898 407414 408134
rect 406794 372454 407414 407898
rect 406794 372218 406826 372454
rect 407062 372218 407146 372454
rect 407382 372218 407414 372454
rect 406794 372134 407414 372218
rect 406794 371898 406826 372134
rect 407062 371898 407146 372134
rect 407382 371898 407414 372134
rect 406794 336454 407414 371898
rect 406794 336218 406826 336454
rect 407062 336218 407146 336454
rect 407382 336218 407414 336454
rect 406794 336134 407414 336218
rect 406794 335898 406826 336134
rect 407062 335898 407146 336134
rect 407382 335898 407414 336134
rect 406794 300454 407414 335898
rect 406794 300218 406826 300454
rect 407062 300218 407146 300454
rect 407382 300218 407414 300454
rect 406794 300134 407414 300218
rect 406794 299898 406826 300134
rect 407062 299898 407146 300134
rect 407382 299898 407414 300134
rect 406794 264454 407414 299898
rect 406794 264218 406826 264454
rect 407062 264218 407146 264454
rect 407382 264218 407414 264454
rect 406794 264134 407414 264218
rect 406794 263898 406826 264134
rect 407062 263898 407146 264134
rect 407382 263898 407414 264134
rect 406794 228454 407414 263898
rect 406794 228218 406826 228454
rect 407062 228218 407146 228454
rect 407382 228218 407414 228454
rect 406794 228134 407414 228218
rect 406794 227898 406826 228134
rect 407062 227898 407146 228134
rect 407382 227898 407414 228134
rect 406794 192454 407414 227898
rect 406794 192218 406826 192454
rect 407062 192218 407146 192454
rect 407382 192218 407414 192454
rect 406794 192134 407414 192218
rect 406794 191898 406826 192134
rect 407062 191898 407146 192134
rect 407382 191898 407414 192134
rect 406794 156454 407414 191898
rect 406794 156218 406826 156454
rect 407062 156218 407146 156454
rect 407382 156218 407414 156454
rect 406794 156134 407414 156218
rect 406794 155898 406826 156134
rect 407062 155898 407146 156134
rect 407382 155898 407414 156134
rect 406794 120454 407414 155898
rect 406794 120218 406826 120454
rect 407062 120218 407146 120454
rect 407382 120218 407414 120454
rect 406794 120134 407414 120218
rect 406794 119898 406826 120134
rect 407062 119898 407146 120134
rect 407382 119898 407414 120134
rect 406794 84454 407414 119898
rect 406794 84218 406826 84454
rect 407062 84218 407146 84454
rect 407382 84218 407414 84454
rect 406794 84134 407414 84218
rect 406794 83898 406826 84134
rect 407062 83898 407146 84134
rect 407382 83898 407414 84134
rect 406794 48454 407414 83898
rect 406794 48218 406826 48454
rect 407062 48218 407146 48454
rect 407382 48218 407414 48454
rect 406794 48134 407414 48218
rect 406794 47898 406826 48134
rect 407062 47898 407146 48134
rect 407382 47898 407414 48134
rect 406794 12454 407414 47898
rect 406794 12218 406826 12454
rect 407062 12218 407146 12454
rect 407382 12218 407414 12454
rect 406794 12134 407414 12218
rect 406794 11898 406826 12134
rect 407062 11898 407146 12134
rect 407382 11898 407414 12134
rect 406794 -2266 407414 11898
rect 406794 -2502 406826 -2266
rect 407062 -2502 407146 -2266
rect 407382 -2502 407414 -2266
rect 406794 -2586 407414 -2502
rect 406794 -2822 406826 -2586
rect 407062 -2822 407146 -2586
rect 407382 -2822 407414 -2586
rect 406794 -7654 407414 -2822
rect 411294 707718 411914 711590
rect 411294 707482 411326 707718
rect 411562 707482 411646 707718
rect 411882 707482 411914 707718
rect 411294 707398 411914 707482
rect 411294 707162 411326 707398
rect 411562 707162 411646 707398
rect 411882 707162 411914 707398
rect 411294 700954 411914 707162
rect 411294 700718 411326 700954
rect 411562 700718 411646 700954
rect 411882 700718 411914 700954
rect 411294 700634 411914 700718
rect 411294 700398 411326 700634
rect 411562 700398 411646 700634
rect 411882 700398 411914 700634
rect 411294 664954 411914 700398
rect 411294 664718 411326 664954
rect 411562 664718 411646 664954
rect 411882 664718 411914 664954
rect 411294 664634 411914 664718
rect 411294 664398 411326 664634
rect 411562 664398 411646 664634
rect 411882 664398 411914 664634
rect 411294 628954 411914 664398
rect 411294 628718 411326 628954
rect 411562 628718 411646 628954
rect 411882 628718 411914 628954
rect 411294 628634 411914 628718
rect 411294 628398 411326 628634
rect 411562 628398 411646 628634
rect 411882 628398 411914 628634
rect 411294 592954 411914 628398
rect 411294 592718 411326 592954
rect 411562 592718 411646 592954
rect 411882 592718 411914 592954
rect 411294 592634 411914 592718
rect 411294 592398 411326 592634
rect 411562 592398 411646 592634
rect 411882 592398 411914 592634
rect 411294 556954 411914 592398
rect 411294 556718 411326 556954
rect 411562 556718 411646 556954
rect 411882 556718 411914 556954
rect 411294 556634 411914 556718
rect 411294 556398 411326 556634
rect 411562 556398 411646 556634
rect 411882 556398 411914 556634
rect 411294 520954 411914 556398
rect 411294 520718 411326 520954
rect 411562 520718 411646 520954
rect 411882 520718 411914 520954
rect 411294 520634 411914 520718
rect 411294 520398 411326 520634
rect 411562 520398 411646 520634
rect 411882 520398 411914 520634
rect 411294 484954 411914 520398
rect 411294 484718 411326 484954
rect 411562 484718 411646 484954
rect 411882 484718 411914 484954
rect 411294 484634 411914 484718
rect 411294 484398 411326 484634
rect 411562 484398 411646 484634
rect 411882 484398 411914 484634
rect 411294 448954 411914 484398
rect 411294 448718 411326 448954
rect 411562 448718 411646 448954
rect 411882 448718 411914 448954
rect 411294 448634 411914 448718
rect 411294 448398 411326 448634
rect 411562 448398 411646 448634
rect 411882 448398 411914 448634
rect 411294 412954 411914 448398
rect 411294 412718 411326 412954
rect 411562 412718 411646 412954
rect 411882 412718 411914 412954
rect 411294 412634 411914 412718
rect 411294 412398 411326 412634
rect 411562 412398 411646 412634
rect 411882 412398 411914 412634
rect 411294 376954 411914 412398
rect 411294 376718 411326 376954
rect 411562 376718 411646 376954
rect 411882 376718 411914 376954
rect 411294 376634 411914 376718
rect 411294 376398 411326 376634
rect 411562 376398 411646 376634
rect 411882 376398 411914 376634
rect 411294 340954 411914 376398
rect 411294 340718 411326 340954
rect 411562 340718 411646 340954
rect 411882 340718 411914 340954
rect 411294 340634 411914 340718
rect 411294 340398 411326 340634
rect 411562 340398 411646 340634
rect 411882 340398 411914 340634
rect 411294 304954 411914 340398
rect 411294 304718 411326 304954
rect 411562 304718 411646 304954
rect 411882 304718 411914 304954
rect 411294 304634 411914 304718
rect 411294 304398 411326 304634
rect 411562 304398 411646 304634
rect 411882 304398 411914 304634
rect 411294 268954 411914 304398
rect 411294 268718 411326 268954
rect 411562 268718 411646 268954
rect 411882 268718 411914 268954
rect 411294 268634 411914 268718
rect 411294 268398 411326 268634
rect 411562 268398 411646 268634
rect 411882 268398 411914 268634
rect 411294 232954 411914 268398
rect 411294 232718 411326 232954
rect 411562 232718 411646 232954
rect 411882 232718 411914 232954
rect 411294 232634 411914 232718
rect 411294 232398 411326 232634
rect 411562 232398 411646 232634
rect 411882 232398 411914 232634
rect 411294 196954 411914 232398
rect 411294 196718 411326 196954
rect 411562 196718 411646 196954
rect 411882 196718 411914 196954
rect 411294 196634 411914 196718
rect 411294 196398 411326 196634
rect 411562 196398 411646 196634
rect 411882 196398 411914 196634
rect 411294 160954 411914 196398
rect 411294 160718 411326 160954
rect 411562 160718 411646 160954
rect 411882 160718 411914 160954
rect 411294 160634 411914 160718
rect 411294 160398 411326 160634
rect 411562 160398 411646 160634
rect 411882 160398 411914 160634
rect 411294 124954 411914 160398
rect 411294 124718 411326 124954
rect 411562 124718 411646 124954
rect 411882 124718 411914 124954
rect 411294 124634 411914 124718
rect 411294 124398 411326 124634
rect 411562 124398 411646 124634
rect 411882 124398 411914 124634
rect 411294 88954 411914 124398
rect 411294 88718 411326 88954
rect 411562 88718 411646 88954
rect 411882 88718 411914 88954
rect 411294 88634 411914 88718
rect 411294 88398 411326 88634
rect 411562 88398 411646 88634
rect 411882 88398 411914 88634
rect 411294 52954 411914 88398
rect 411294 52718 411326 52954
rect 411562 52718 411646 52954
rect 411882 52718 411914 52954
rect 411294 52634 411914 52718
rect 411294 52398 411326 52634
rect 411562 52398 411646 52634
rect 411882 52398 411914 52634
rect 411294 16954 411914 52398
rect 411294 16718 411326 16954
rect 411562 16718 411646 16954
rect 411882 16718 411914 16954
rect 411294 16634 411914 16718
rect 411294 16398 411326 16634
rect 411562 16398 411646 16634
rect 411882 16398 411914 16634
rect 411294 -3226 411914 16398
rect 411294 -3462 411326 -3226
rect 411562 -3462 411646 -3226
rect 411882 -3462 411914 -3226
rect 411294 -3546 411914 -3462
rect 411294 -3782 411326 -3546
rect 411562 -3782 411646 -3546
rect 411882 -3782 411914 -3546
rect 411294 -7654 411914 -3782
rect 415794 708678 416414 711590
rect 415794 708442 415826 708678
rect 416062 708442 416146 708678
rect 416382 708442 416414 708678
rect 415794 708358 416414 708442
rect 415794 708122 415826 708358
rect 416062 708122 416146 708358
rect 416382 708122 416414 708358
rect 415794 669454 416414 708122
rect 415794 669218 415826 669454
rect 416062 669218 416146 669454
rect 416382 669218 416414 669454
rect 415794 669134 416414 669218
rect 415794 668898 415826 669134
rect 416062 668898 416146 669134
rect 416382 668898 416414 669134
rect 415794 633454 416414 668898
rect 415794 633218 415826 633454
rect 416062 633218 416146 633454
rect 416382 633218 416414 633454
rect 415794 633134 416414 633218
rect 415794 632898 415826 633134
rect 416062 632898 416146 633134
rect 416382 632898 416414 633134
rect 415794 597454 416414 632898
rect 415794 597218 415826 597454
rect 416062 597218 416146 597454
rect 416382 597218 416414 597454
rect 415794 597134 416414 597218
rect 415794 596898 415826 597134
rect 416062 596898 416146 597134
rect 416382 596898 416414 597134
rect 415794 561454 416414 596898
rect 415794 561218 415826 561454
rect 416062 561218 416146 561454
rect 416382 561218 416414 561454
rect 415794 561134 416414 561218
rect 415794 560898 415826 561134
rect 416062 560898 416146 561134
rect 416382 560898 416414 561134
rect 415794 525454 416414 560898
rect 415794 525218 415826 525454
rect 416062 525218 416146 525454
rect 416382 525218 416414 525454
rect 415794 525134 416414 525218
rect 415794 524898 415826 525134
rect 416062 524898 416146 525134
rect 416382 524898 416414 525134
rect 415794 489454 416414 524898
rect 415794 489218 415826 489454
rect 416062 489218 416146 489454
rect 416382 489218 416414 489454
rect 415794 489134 416414 489218
rect 415794 488898 415826 489134
rect 416062 488898 416146 489134
rect 416382 488898 416414 489134
rect 415794 453454 416414 488898
rect 415794 453218 415826 453454
rect 416062 453218 416146 453454
rect 416382 453218 416414 453454
rect 415794 453134 416414 453218
rect 415794 452898 415826 453134
rect 416062 452898 416146 453134
rect 416382 452898 416414 453134
rect 415794 417454 416414 452898
rect 415794 417218 415826 417454
rect 416062 417218 416146 417454
rect 416382 417218 416414 417454
rect 415794 417134 416414 417218
rect 415794 416898 415826 417134
rect 416062 416898 416146 417134
rect 416382 416898 416414 417134
rect 415794 381454 416414 416898
rect 415794 381218 415826 381454
rect 416062 381218 416146 381454
rect 416382 381218 416414 381454
rect 415794 381134 416414 381218
rect 415794 380898 415826 381134
rect 416062 380898 416146 381134
rect 416382 380898 416414 381134
rect 415794 345454 416414 380898
rect 415794 345218 415826 345454
rect 416062 345218 416146 345454
rect 416382 345218 416414 345454
rect 415794 345134 416414 345218
rect 415794 344898 415826 345134
rect 416062 344898 416146 345134
rect 416382 344898 416414 345134
rect 415794 309454 416414 344898
rect 415794 309218 415826 309454
rect 416062 309218 416146 309454
rect 416382 309218 416414 309454
rect 415794 309134 416414 309218
rect 415794 308898 415826 309134
rect 416062 308898 416146 309134
rect 416382 308898 416414 309134
rect 415794 273454 416414 308898
rect 415794 273218 415826 273454
rect 416062 273218 416146 273454
rect 416382 273218 416414 273454
rect 415794 273134 416414 273218
rect 415794 272898 415826 273134
rect 416062 272898 416146 273134
rect 416382 272898 416414 273134
rect 415794 237454 416414 272898
rect 415794 237218 415826 237454
rect 416062 237218 416146 237454
rect 416382 237218 416414 237454
rect 415794 237134 416414 237218
rect 415794 236898 415826 237134
rect 416062 236898 416146 237134
rect 416382 236898 416414 237134
rect 415794 201454 416414 236898
rect 415794 201218 415826 201454
rect 416062 201218 416146 201454
rect 416382 201218 416414 201454
rect 415794 201134 416414 201218
rect 415794 200898 415826 201134
rect 416062 200898 416146 201134
rect 416382 200898 416414 201134
rect 415794 165454 416414 200898
rect 415794 165218 415826 165454
rect 416062 165218 416146 165454
rect 416382 165218 416414 165454
rect 415794 165134 416414 165218
rect 415794 164898 415826 165134
rect 416062 164898 416146 165134
rect 416382 164898 416414 165134
rect 415794 129454 416414 164898
rect 415794 129218 415826 129454
rect 416062 129218 416146 129454
rect 416382 129218 416414 129454
rect 415794 129134 416414 129218
rect 415794 128898 415826 129134
rect 416062 128898 416146 129134
rect 416382 128898 416414 129134
rect 415794 93454 416414 128898
rect 415794 93218 415826 93454
rect 416062 93218 416146 93454
rect 416382 93218 416414 93454
rect 415794 93134 416414 93218
rect 415794 92898 415826 93134
rect 416062 92898 416146 93134
rect 416382 92898 416414 93134
rect 415794 57454 416414 92898
rect 415794 57218 415826 57454
rect 416062 57218 416146 57454
rect 416382 57218 416414 57454
rect 415794 57134 416414 57218
rect 415794 56898 415826 57134
rect 416062 56898 416146 57134
rect 416382 56898 416414 57134
rect 415794 21454 416414 56898
rect 415794 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 416414 21454
rect 415794 21134 416414 21218
rect 415794 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 416414 21134
rect 415794 -4186 416414 20898
rect 415794 -4422 415826 -4186
rect 416062 -4422 416146 -4186
rect 416382 -4422 416414 -4186
rect 415794 -4506 416414 -4422
rect 415794 -4742 415826 -4506
rect 416062 -4742 416146 -4506
rect 416382 -4742 416414 -4506
rect 415794 -7654 416414 -4742
rect 420294 709638 420914 711590
rect 420294 709402 420326 709638
rect 420562 709402 420646 709638
rect 420882 709402 420914 709638
rect 420294 709318 420914 709402
rect 420294 709082 420326 709318
rect 420562 709082 420646 709318
rect 420882 709082 420914 709318
rect 420294 673954 420914 709082
rect 420294 673718 420326 673954
rect 420562 673718 420646 673954
rect 420882 673718 420914 673954
rect 420294 673634 420914 673718
rect 420294 673398 420326 673634
rect 420562 673398 420646 673634
rect 420882 673398 420914 673634
rect 420294 637954 420914 673398
rect 420294 637718 420326 637954
rect 420562 637718 420646 637954
rect 420882 637718 420914 637954
rect 420294 637634 420914 637718
rect 420294 637398 420326 637634
rect 420562 637398 420646 637634
rect 420882 637398 420914 637634
rect 420294 601954 420914 637398
rect 420294 601718 420326 601954
rect 420562 601718 420646 601954
rect 420882 601718 420914 601954
rect 420294 601634 420914 601718
rect 420294 601398 420326 601634
rect 420562 601398 420646 601634
rect 420882 601398 420914 601634
rect 420294 565954 420914 601398
rect 420294 565718 420326 565954
rect 420562 565718 420646 565954
rect 420882 565718 420914 565954
rect 420294 565634 420914 565718
rect 420294 565398 420326 565634
rect 420562 565398 420646 565634
rect 420882 565398 420914 565634
rect 420294 529954 420914 565398
rect 420294 529718 420326 529954
rect 420562 529718 420646 529954
rect 420882 529718 420914 529954
rect 420294 529634 420914 529718
rect 420294 529398 420326 529634
rect 420562 529398 420646 529634
rect 420882 529398 420914 529634
rect 420294 493954 420914 529398
rect 420294 493718 420326 493954
rect 420562 493718 420646 493954
rect 420882 493718 420914 493954
rect 420294 493634 420914 493718
rect 420294 493398 420326 493634
rect 420562 493398 420646 493634
rect 420882 493398 420914 493634
rect 420294 457954 420914 493398
rect 420294 457718 420326 457954
rect 420562 457718 420646 457954
rect 420882 457718 420914 457954
rect 420294 457634 420914 457718
rect 420294 457398 420326 457634
rect 420562 457398 420646 457634
rect 420882 457398 420914 457634
rect 420294 421954 420914 457398
rect 420294 421718 420326 421954
rect 420562 421718 420646 421954
rect 420882 421718 420914 421954
rect 420294 421634 420914 421718
rect 420294 421398 420326 421634
rect 420562 421398 420646 421634
rect 420882 421398 420914 421634
rect 420294 385954 420914 421398
rect 420294 385718 420326 385954
rect 420562 385718 420646 385954
rect 420882 385718 420914 385954
rect 420294 385634 420914 385718
rect 420294 385398 420326 385634
rect 420562 385398 420646 385634
rect 420882 385398 420914 385634
rect 420294 349954 420914 385398
rect 420294 349718 420326 349954
rect 420562 349718 420646 349954
rect 420882 349718 420914 349954
rect 420294 349634 420914 349718
rect 420294 349398 420326 349634
rect 420562 349398 420646 349634
rect 420882 349398 420914 349634
rect 420294 313954 420914 349398
rect 420294 313718 420326 313954
rect 420562 313718 420646 313954
rect 420882 313718 420914 313954
rect 420294 313634 420914 313718
rect 420294 313398 420326 313634
rect 420562 313398 420646 313634
rect 420882 313398 420914 313634
rect 420294 277954 420914 313398
rect 420294 277718 420326 277954
rect 420562 277718 420646 277954
rect 420882 277718 420914 277954
rect 420294 277634 420914 277718
rect 420294 277398 420326 277634
rect 420562 277398 420646 277634
rect 420882 277398 420914 277634
rect 420294 241954 420914 277398
rect 420294 241718 420326 241954
rect 420562 241718 420646 241954
rect 420882 241718 420914 241954
rect 420294 241634 420914 241718
rect 420294 241398 420326 241634
rect 420562 241398 420646 241634
rect 420882 241398 420914 241634
rect 420294 205954 420914 241398
rect 420294 205718 420326 205954
rect 420562 205718 420646 205954
rect 420882 205718 420914 205954
rect 420294 205634 420914 205718
rect 420294 205398 420326 205634
rect 420562 205398 420646 205634
rect 420882 205398 420914 205634
rect 420294 169954 420914 205398
rect 420294 169718 420326 169954
rect 420562 169718 420646 169954
rect 420882 169718 420914 169954
rect 420294 169634 420914 169718
rect 420294 169398 420326 169634
rect 420562 169398 420646 169634
rect 420882 169398 420914 169634
rect 420294 133954 420914 169398
rect 420294 133718 420326 133954
rect 420562 133718 420646 133954
rect 420882 133718 420914 133954
rect 420294 133634 420914 133718
rect 420294 133398 420326 133634
rect 420562 133398 420646 133634
rect 420882 133398 420914 133634
rect 420294 97954 420914 133398
rect 420294 97718 420326 97954
rect 420562 97718 420646 97954
rect 420882 97718 420914 97954
rect 420294 97634 420914 97718
rect 420294 97398 420326 97634
rect 420562 97398 420646 97634
rect 420882 97398 420914 97634
rect 420294 61954 420914 97398
rect 420294 61718 420326 61954
rect 420562 61718 420646 61954
rect 420882 61718 420914 61954
rect 420294 61634 420914 61718
rect 420294 61398 420326 61634
rect 420562 61398 420646 61634
rect 420882 61398 420914 61634
rect 420294 25954 420914 61398
rect 420294 25718 420326 25954
rect 420562 25718 420646 25954
rect 420882 25718 420914 25954
rect 420294 25634 420914 25718
rect 420294 25398 420326 25634
rect 420562 25398 420646 25634
rect 420882 25398 420914 25634
rect 420294 -5146 420914 25398
rect 420294 -5382 420326 -5146
rect 420562 -5382 420646 -5146
rect 420882 -5382 420914 -5146
rect 420294 -5466 420914 -5382
rect 420294 -5702 420326 -5466
rect 420562 -5702 420646 -5466
rect 420882 -5702 420914 -5466
rect 420294 -7654 420914 -5702
rect 424794 710598 425414 711590
rect 424794 710362 424826 710598
rect 425062 710362 425146 710598
rect 425382 710362 425414 710598
rect 424794 710278 425414 710362
rect 424794 710042 424826 710278
rect 425062 710042 425146 710278
rect 425382 710042 425414 710278
rect 424794 678454 425414 710042
rect 424794 678218 424826 678454
rect 425062 678218 425146 678454
rect 425382 678218 425414 678454
rect 424794 678134 425414 678218
rect 424794 677898 424826 678134
rect 425062 677898 425146 678134
rect 425382 677898 425414 678134
rect 424794 642454 425414 677898
rect 424794 642218 424826 642454
rect 425062 642218 425146 642454
rect 425382 642218 425414 642454
rect 424794 642134 425414 642218
rect 424794 641898 424826 642134
rect 425062 641898 425146 642134
rect 425382 641898 425414 642134
rect 424794 606454 425414 641898
rect 424794 606218 424826 606454
rect 425062 606218 425146 606454
rect 425382 606218 425414 606454
rect 424794 606134 425414 606218
rect 424794 605898 424826 606134
rect 425062 605898 425146 606134
rect 425382 605898 425414 606134
rect 424794 570454 425414 605898
rect 424794 570218 424826 570454
rect 425062 570218 425146 570454
rect 425382 570218 425414 570454
rect 424794 570134 425414 570218
rect 424794 569898 424826 570134
rect 425062 569898 425146 570134
rect 425382 569898 425414 570134
rect 424794 534454 425414 569898
rect 424794 534218 424826 534454
rect 425062 534218 425146 534454
rect 425382 534218 425414 534454
rect 424794 534134 425414 534218
rect 424794 533898 424826 534134
rect 425062 533898 425146 534134
rect 425382 533898 425414 534134
rect 424794 498454 425414 533898
rect 424794 498218 424826 498454
rect 425062 498218 425146 498454
rect 425382 498218 425414 498454
rect 424794 498134 425414 498218
rect 424794 497898 424826 498134
rect 425062 497898 425146 498134
rect 425382 497898 425414 498134
rect 424794 462454 425414 497898
rect 424794 462218 424826 462454
rect 425062 462218 425146 462454
rect 425382 462218 425414 462454
rect 424794 462134 425414 462218
rect 424794 461898 424826 462134
rect 425062 461898 425146 462134
rect 425382 461898 425414 462134
rect 424794 426454 425414 461898
rect 424794 426218 424826 426454
rect 425062 426218 425146 426454
rect 425382 426218 425414 426454
rect 424794 426134 425414 426218
rect 424794 425898 424826 426134
rect 425062 425898 425146 426134
rect 425382 425898 425414 426134
rect 424794 390454 425414 425898
rect 424794 390218 424826 390454
rect 425062 390218 425146 390454
rect 425382 390218 425414 390454
rect 424794 390134 425414 390218
rect 424794 389898 424826 390134
rect 425062 389898 425146 390134
rect 425382 389898 425414 390134
rect 424794 354454 425414 389898
rect 424794 354218 424826 354454
rect 425062 354218 425146 354454
rect 425382 354218 425414 354454
rect 424794 354134 425414 354218
rect 424794 353898 424826 354134
rect 425062 353898 425146 354134
rect 425382 353898 425414 354134
rect 424794 318454 425414 353898
rect 424794 318218 424826 318454
rect 425062 318218 425146 318454
rect 425382 318218 425414 318454
rect 424794 318134 425414 318218
rect 424794 317898 424826 318134
rect 425062 317898 425146 318134
rect 425382 317898 425414 318134
rect 424794 282454 425414 317898
rect 424794 282218 424826 282454
rect 425062 282218 425146 282454
rect 425382 282218 425414 282454
rect 424794 282134 425414 282218
rect 424794 281898 424826 282134
rect 425062 281898 425146 282134
rect 425382 281898 425414 282134
rect 424794 246454 425414 281898
rect 424794 246218 424826 246454
rect 425062 246218 425146 246454
rect 425382 246218 425414 246454
rect 424794 246134 425414 246218
rect 424794 245898 424826 246134
rect 425062 245898 425146 246134
rect 425382 245898 425414 246134
rect 424794 210454 425414 245898
rect 424794 210218 424826 210454
rect 425062 210218 425146 210454
rect 425382 210218 425414 210454
rect 424794 210134 425414 210218
rect 424794 209898 424826 210134
rect 425062 209898 425146 210134
rect 425382 209898 425414 210134
rect 424794 174454 425414 209898
rect 424794 174218 424826 174454
rect 425062 174218 425146 174454
rect 425382 174218 425414 174454
rect 424794 174134 425414 174218
rect 424794 173898 424826 174134
rect 425062 173898 425146 174134
rect 425382 173898 425414 174134
rect 424794 138454 425414 173898
rect 424794 138218 424826 138454
rect 425062 138218 425146 138454
rect 425382 138218 425414 138454
rect 424794 138134 425414 138218
rect 424794 137898 424826 138134
rect 425062 137898 425146 138134
rect 425382 137898 425414 138134
rect 424794 102454 425414 137898
rect 424794 102218 424826 102454
rect 425062 102218 425146 102454
rect 425382 102218 425414 102454
rect 424794 102134 425414 102218
rect 424794 101898 424826 102134
rect 425062 101898 425146 102134
rect 425382 101898 425414 102134
rect 424794 66454 425414 101898
rect 424794 66218 424826 66454
rect 425062 66218 425146 66454
rect 425382 66218 425414 66454
rect 424794 66134 425414 66218
rect 424794 65898 424826 66134
rect 425062 65898 425146 66134
rect 425382 65898 425414 66134
rect 424794 30454 425414 65898
rect 424794 30218 424826 30454
rect 425062 30218 425146 30454
rect 425382 30218 425414 30454
rect 424794 30134 425414 30218
rect 424794 29898 424826 30134
rect 425062 29898 425146 30134
rect 425382 29898 425414 30134
rect 424794 -6106 425414 29898
rect 424794 -6342 424826 -6106
rect 425062 -6342 425146 -6106
rect 425382 -6342 425414 -6106
rect 424794 -6426 425414 -6342
rect 424794 -6662 424826 -6426
rect 425062 -6662 425146 -6426
rect 425382 -6662 425414 -6426
rect 424794 -7654 425414 -6662
rect 429294 711558 429914 711590
rect 429294 711322 429326 711558
rect 429562 711322 429646 711558
rect 429882 711322 429914 711558
rect 429294 711238 429914 711322
rect 429294 711002 429326 711238
rect 429562 711002 429646 711238
rect 429882 711002 429914 711238
rect 429294 682954 429914 711002
rect 429294 682718 429326 682954
rect 429562 682718 429646 682954
rect 429882 682718 429914 682954
rect 429294 682634 429914 682718
rect 429294 682398 429326 682634
rect 429562 682398 429646 682634
rect 429882 682398 429914 682634
rect 429294 646954 429914 682398
rect 429294 646718 429326 646954
rect 429562 646718 429646 646954
rect 429882 646718 429914 646954
rect 429294 646634 429914 646718
rect 429294 646398 429326 646634
rect 429562 646398 429646 646634
rect 429882 646398 429914 646634
rect 429294 610954 429914 646398
rect 429294 610718 429326 610954
rect 429562 610718 429646 610954
rect 429882 610718 429914 610954
rect 429294 610634 429914 610718
rect 429294 610398 429326 610634
rect 429562 610398 429646 610634
rect 429882 610398 429914 610634
rect 429294 574954 429914 610398
rect 429294 574718 429326 574954
rect 429562 574718 429646 574954
rect 429882 574718 429914 574954
rect 429294 574634 429914 574718
rect 429294 574398 429326 574634
rect 429562 574398 429646 574634
rect 429882 574398 429914 574634
rect 429294 538954 429914 574398
rect 429294 538718 429326 538954
rect 429562 538718 429646 538954
rect 429882 538718 429914 538954
rect 429294 538634 429914 538718
rect 429294 538398 429326 538634
rect 429562 538398 429646 538634
rect 429882 538398 429914 538634
rect 429294 502954 429914 538398
rect 429294 502718 429326 502954
rect 429562 502718 429646 502954
rect 429882 502718 429914 502954
rect 429294 502634 429914 502718
rect 429294 502398 429326 502634
rect 429562 502398 429646 502634
rect 429882 502398 429914 502634
rect 429294 466954 429914 502398
rect 429294 466718 429326 466954
rect 429562 466718 429646 466954
rect 429882 466718 429914 466954
rect 429294 466634 429914 466718
rect 429294 466398 429326 466634
rect 429562 466398 429646 466634
rect 429882 466398 429914 466634
rect 429294 430954 429914 466398
rect 429294 430718 429326 430954
rect 429562 430718 429646 430954
rect 429882 430718 429914 430954
rect 429294 430634 429914 430718
rect 429294 430398 429326 430634
rect 429562 430398 429646 430634
rect 429882 430398 429914 430634
rect 429294 394954 429914 430398
rect 429294 394718 429326 394954
rect 429562 394718 429646 394954
rect 429882 394718 429914 394954
rect 429294 394634 429914 394718
rect 429294 394398 429326 394634
rect 429562 394398 429646 394634
rect 429882 394398 429914 394634
rect 429294 358954 429914 394398
rect 429294 358718 429326 358954
rect 429562 358718 429646 358954
rect 429882 358718 429914 358954
rect 429294 358634 429914 358718
rect 429294 358398 429326 358634
rect 429562 358398 429646 358634
rect 429882 358398 429914 358634
rect 429294 322954 429914 358398
rect 429294 322718 429326 322954
rect 429562 322718 429646 322954
rect 429882 322718 429914 322954
rect 429294 322634 429914 322718
rect 429294 322398 429326 322634
rect 429562 322398 429646 322634
rect 429882 322398 429914 322634
rect 429294 286954 429914 322398
rect 429294 286718 429326 286954
rect 429562 286718 429646 286954
rect 429882 286718 429914 286954
rect 429294 286634 429914 286718
rect 429294 286398 429326 286634
rect 429562 286398 429646 286634
rect 429882 286398 429914 286634
rect 429294 250954 429914 286398
rect 429294 250718 429326 250954
rect 429562 250718 429646 250954
rect 429882 250718 429914 250954
rect 429294 250634 429914 250718
rect 429294 250398 429326 250634
rect 429562 250398 429646 250634
rect 429882 250398 429914 250634
rect 429294 214954 429914 250398
rect 429294 214718 429326 214954
rect 429562 214718 429646 214954
rect 429882 214718 429914 214954
rect 429294 214634 429914 214718
rect 429294 214398 429326 214634
rect 429562 214398 429646 214634
rect 429882 214398 429914 214634
rect 429294 178954 429914 214398
rect 429294 178718 429326 178954
rect 429562 178718 429646 178954
rect 429882 178718 429914 178954
rect 429294 178634 429914 178718
rect 429294 178398 429326 178634
rect 429562 178398 429646 178634
rect 429882 178398 429914 178634
rect 429294 142954 429914 178398
rect 429294 142718 429326 142954
rect 429562 142718 429646 142954
rect 429882 142718 429914 142954
rect 429294 142634 429914 142718
rect 429294 142398 429326 142634
rect 429562 142398 429646 142634
rect 429882 142398 429914 142634
rect 429294 106954 429914 142398
rect 429294 106718 429326 106954
rect 429562 106718 429646 106954
rect 429882 106718 429914 106954
rect 429294 106634 429914 106718
rect 429294 106398 429326 106634
rect 429562 106398 429646 106634
rect 429882 106398 429914 106634
rect 429294 70954 429914 106398
rect 429294 70718 429326 70954
rect 429562 70718 429646 70954
rect 429882 70718 429914 70954
rect 429294 70634 429914 70718
rect 429294 70398 429326 70634
rect 429562 70398 429646 70634
rect 429882 70398 429914 70634
rect 429294 34954 429914 70398
rect 429294 34718 429326 34954
rect 429562 34718 429646 34954
rect 429882 34718 429914 34954
rect 429294 34634 429914 34718
rect 429294 34398 429326 34634
rect 429562 34398 429646 34634
rect 429882 34398 429914 34634
rect 429294 -7066 429914 34398
rect 429294 -7302 429326 -7066
rect 429562 -7302 429646 -7066
rect 429882 -7302 429914 -7066
rect 429294 -7386 429914 -7302
rect 429294 -7622 429326 -7386
rect 429562 -7622 429646 -7386
rect 429882 -7622 429914 -7386
rect 429294 -7654 429914 -7622
rect 433794 704838 434414 711590
rect 433794 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 434414 704838
rect 433794 704518 434414 704602
rect 433794 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 434414 704518
rect 433794 687454 434414 704282
rect 433794 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 434414 687454
rect 433794 687134 434414 687218
rect 433794 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 434414 687134
rect 433794 651454 434414 686898
rect 433794 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 434414 651454
rect 433794 651134 434414 651218
rect 433794 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 434414 651134
rect 433794 615454 434414 650898
rect 433794 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 434414 615454
rect 433794 615134 434414 615218
rect 433794 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 434414 615134
rect 433794 579454 434414 614898
rect 433794 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 434414 579454
rect 433794 579134 434414 579218
rect 433794 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 434414 579134
rect 433794 543454 434414 578898
rect 433794 543218 433826 543454
rect 434062 543218 434146 543454
rect 434382 543218 434414 543454
rect 433794 543134 434414 543218
rect 433794 542898 433826 543134
rect 434062 542898 434146 543134
rect 434382 542898 434414 543134
rect 433794 507454 434414 542898
rect 433794 507218 433826 507454
rect 434062 507218 434146 507454
rect 434382 507218 434414 507454
rect 433794 507134 434414 507218
rect 433794 506898 433826 507134
rect 434062 506898 434146 507134
rect 434382 506898 434414 507134
rect 433794 471454 434414 506898
rect 433794 471218 433826 471454
rect 434062 471218 434146 471454
rect 434382 471218 434414 471454
rect 433794 471134 434414 471218
rect 433794 470898 433826 471134
rect 434062 470898 434146 471134
rect 434382 470898 434414 471134
rect 433794 435454 434414 470898
rect 433794 435218 433826 435454
rect 434062 435218 434146 435454
rect 434382 435218 434414 435454
rect 433794 435134 434414 435218
rect 433794 434898 433826 435134
rect 434062 434898 434146 435134
rect 434382 434898 434414 435134
rect 433794 399454 434414 434898
rect 433794 399218 433826 399454
rect 434062 399218 434146 399454
rect 434382 399218 434414 399454
rect 433794 399134 434414 399218
rect 433794 398898 433826 399134
rect 434062 398898 434146 399134
rect 434382 398898 434414 399134
rect 433794 363454 434414 398898
rect 433794 363218 433826 363454
rect 434062 363218 434146 363454
rect 434382 363218 434414 363454
rect 433794 363134 434414 363218
rect 433794 362898 433826 363134
rect 434062 362898 434146 363134
rect 434382 362898 434414 363134
rect 433794 327454 434414 362898
rect 433794 327218 433826 327454
rect 434062 327218 434146 327454
rect 434382 327218 434414 327454
rect 433794 327134 434414 327218
rect 433794 326898 433826 327134
rect 434062 326898 434146 327134
rect 434382 326898 434414 327134
rect 433794 291454 434414 326898
rect 433794 291218 433826 291454
rect 434062 291218 434146 291454
rect 434382 291218 434414 291454
rect 433794 291134 434414 291218
rect 433794 290898 433826 291134
rect 434062 290898 434146 291134
rect 434382 290898 434414 291134
rect 433794 255454 434414 290898
rect 433794 255218 433826 255454
rect 434062 255218 434146 255454
rect 434382 255218 434414 255454
rect 433794 255134 434414 255218
rect 433794 254898 433826 255134
rect 434062 254898 434146 255134
rect 434382 254898 434414 255134
rect 433794 219454 434414 254898
rect 433794 219218 433826 219454
rect 434062 219218 434146 219454
rect 434382 219218 434414 219454
rect 433794 219134 434414 219218
rect 433794 218898 433826 219134
rect 434062 218898 434146 219134
rect 434382 218898 434414 219134
rect 433794 183454 434414 218898
rect 433794 183218 433826 183454
rect 434062 183218 434146 183454
rect 434382 183218 434414 183454
rect 433794 183134 434414 183218
rect 433794 182898 433826 183134
rect 434062 182898 434146 183134
rect 434382 182898 434414 183134
rect 433794 147454 434414 182898
rect 433794 147218 433826 147454
rect 434062 147218 434146 147454
rect 434382 147218 434414 147454
rect 433794 147134 434414 147218
rect 433794 146898 433826 147134
rect 434062 146898 434146 147134
rect 434382 146898 434414 147134
rect 433794 111454 434414 146898
rect 433794 111218 433826 111454
rect 434062 111218 434146 111454
rect 434382 111218 434414 111454
rect 433794 111134 434414 111218
rect 433794 110898 433826 111134
rect 434062 110898 434146 111134
rect 434382 110898 434414 111134
rect 433794 75454 434414 110898
rect 433794 75218 433826 75454
rect 434062 75218 434146 75454
rect 434382 75218 434414 75454
rect 433794 75134 434414 75218
rect 433794 74898 433826 75134
rect 434062 74898 434146 75134
rect 434382 74898 434414 75134
rect 433794 39454 434414 74898
rect 433794 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 434414 39454
rect 433794 39134 434414 39218
rect 433794 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 434414 39134
rect 433794 3454 434414 38898
rect 433794 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 434414 3454
rect 433794 3134 434414 3218
rect 433794 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 434414 3134
rect 433794 -346 434414 2898
rect 433794 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 434414 -346
rect 433794 -666 434414 -582
rect 433794 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 434414 -666
rect 433794 -7654 434414 -902
rect 438294 705798 438914 711590
rect 438294 705562 438326 705798
rect 438562 705562 438646 705798
rect 438882 705562 438914 705798
rect 438294 705478 438914 705562
rect 438294 705242 438326 705478
rect 438562 705242 438646 705478
rect 438882 705242 438914 705478
rect 438294 691954 438914 705242
rect 438294 691718 438326 691954
rect 438562 691718 438646 691954
rect 438882 691718 438914 691954
rect 438294 691634 438914 691718
rect 438294 691398 438326 691634
rect 438562 691398 438646 691634
rect 438882 691398 438914 691634
rect 438294 655954 438914 691398
rect 438294 655718 438326 655954
rect 438562 655718 438646 655954
rect 438882 655718 438914 655954
rect 438294 655634 438914 655718
rect 438294 655398 438326 655634
rect 438562 655398 438646 655634
rect 438882 655398 438914 655634
rect 438294 619954 438914 655398
rect 438294 619718 438326 619954
rect 438562 619718 438646 619954
rect 438882 619718 438914 619954
rect 438294 619634 438914 619718
rect 438294 619398 438326 619634
rect 438562 619398 438646 619634
rect 438882 619398 438914 619634
rect 438294 583954 438914 619398
rect 438294 583718 438326 583954
rect 438562 583718 438646 583954
rect 438882 583718 438914 583954
rect 438294 583634 438914 583718
rect 438294 583398 438326 583634
rect 438562 583398 438646 583634
rect 438882 583398 438914 583634
rect 438294 547954 438914 583398
rect 438294 547718 438326 547954
rect 438562 547718 438646 547954
rect 438882 547718 438914 547954
rect 438294 547634 438914 547718
rect 438294 547398 438326 547634
rect 438562 547398 438646 547634
rect 438882 547398 438914 547634
rect 438294 511954 438914 547398
rect 438294 511718 438326 511954
rect 438562 511718 438646 511954
rect 438882 511718 438914 511954
rect 438294 511634 438914 511718
rect 438294 511398 438326 511634
rect 438562 511398 438646 511634
rect 438882 511398 438914 511634
rect 438294 475954 438914 511398
rect 438294 475718 438326 475954
rect 438562 475718 438646 475954
rect 438882 475718 438914 475954
rect 438294 475634 438914 475718
rect 438294 475398 438326 475634
rect 438562 475398 438646 475634
rect 438882 475398 438914 475634
rect 438294 439954 438914 475398
rect 438294 439718 438326 439954
rect 438562 439718 438646 439954
rect 438882 439718 438914 439954
rect 438294 439634 438914 439718
rect 438294 439398 438326 439634
rect 438562 439398 438646 439634
rect 438882 439398 438914 439634
rect 438294 403954 438914 439398
rect 438294 403718 438326 403954
rect 438562 403718 438646 403954
rect 438882 403718 438914 403954
rect 438294 403634 438914 403718
rect 438294 403398 438326 403634
rect 438562 403398 438646 403634
rect 438882 403398 438914 403634
rect 438294 367954 438914 403398
rect 438294 367718 438326 367954
rect 438562 367718 438646 367954
rect 438882 367718 438914 367954
rect 438294 367634 438914 367718
rect 438294 367398 438326 367634
rect 438562 367398 438646 367634
rect 438882 367398 438914 367634
rect 438294 331954 438914 367398
rect 438294 331718 438326 331954
rect 438562 331718 438646 331954
rect 438882 331718 438914 331954
rect 438294 331634 438914 331718
rect 438294 331398 438326 331634
rect 438562 331398 438646 331634
rect 438882 331398 438914 331634
rect 438294 295954 438914 331398
rect 438294 295718 438326 295954
rect 438562 295718 438646 295954
rect 438882 295718 438914 295954
rect 438294 295634 438914 295718
rect 438294 295398 438326 295634
rect 438562 295398 438646 295634
rect 438882 295398 438914 295634
rect 438294 259954 438914 295398
rect 438294 259718 438326 259954
rect 438562 259718 438646 259954
rect 438882 259718 438914 259954
rect 438294 259634 438914 259718
rect 438294 259398 438326 259634
rect 438562 259398 438646 259634
rect 438882 259398 438914 259634
rect 438294 223954 438914 259398
rect 438294 223718 438326 223954
rect 438562 223718 438646 223954
rect 438882 223718 438914 223954
rect 438294 223634 438914 223718
rect 438294 223398 438326 223634
rect 438562 223398 438646 223634
rect 438882 223398 438914 223634
rect 438294 187954 438914 223398
rect 438294 187718 438326 187954
rect 438562 187718 438646 187954
rect 438882 187718 438914 187954
rect 438294 187634 438914 187718
rect 438294 187398 438326 187634
rect 438562 187398 438646 187634
rect 438882 187398 438914 187634
rect 438294 151954 438914 187398
rect 438294 151718 438326 151954
rect 438562 151718 438646 151954
rect 438882 151718 438914 151954
rect 438294 151634 438914 151718
rect 438294 151398 438326 151634
rect 438562 151398 438646 151634
rect 438882 151398 438914 151634
rect 438294 115954 438914 151398
rect 438294 115718 438326 115954
rect 438562 115718 438646 115954
rect 438882 115718 438914 115954
rect 438294 115634 438914 115718
rect 438294 115398 438326 115634
rect 438562 115398 438646 115634
rect 438882 115398 438914 115634
rect 438294 79954 438914 115398
rect 438294 79718 438326 79954
rect 438562 79718 438646 79954
rect 438882 79718 438914 79954
rect 438294 79634 438914 79718
rect 438294 79398 438326 79634
rect 438562 79398 438646 79634
rect 438882 79398 438914 79634
rect 438294 43954 438914 79398
rect 438294 43718 438326 43954
rect 438562 43718 438646 43954
rect 438882 43718 438914 43954
rect 438294 43634 438914 43718
rect 438294 43398 438326 43634
rect 438562 43398 438646 43634
rect 438882 43398 438914 43634
rect 438294 7954 438914 43398
rect 438294 7718 438326 7954
rect 438562 7718 438646 7954
rect 438882 7718 438914 7954
rect 438294 7634 438914 7718
rect 438294 7398 438326 7634
rect 438562 7398 438646 7634
rect 438882 7398 438914 7634
rect 438294 -1306 438914 7398
rect 438294 -1542 438326 -1306
rect 438562 -1542 438646 -1306
rect 438882 -1542 438914 -1306
rect 438294 -1626 438914 -1542
rect 438294 -1862 438326 -1626
rect 438562 -1862 438646 -1626
rect 438882 -1862 438914 -1626
rect 438294 -7654 438914 -1862
rect 442794 706758 443414 711590
rect 442794 706522 442826 706758
rect 443062 706522 443146 706758
rect 443382 706522 443414 706758
rect 442794 706438 443414 706522
rect 442794 706202 442826 706438
rect 443062 706202 443146 706438
rect 443382 706202 443414 706438
rect 442794 696454 443414 706202
rect 442794 696218 442826 696454
rect 443062 696218 443146 696454
rect 443382 696218 443414 696454
rect 442794 696134 443414 696218
rect 442794 695898 442826 696134
rect 443062 695898 443146 696134
rect 443382 695898 443414 696134
rect 442794 660454 443414 695898
rect 442794 660218 442826 660454
rect 443062 660218 443146 660454
rect 443382 660218 443414 660454
rect 442794 660134 443414 660218
rect 442794 659898 442826 660134
rect 443062 659898 443146 660134
rect 443382 659898 443414 660134
rect 442794 624454 443414 659898
rect 442794 624218 442826 624454
rect 443062 624218 443146 624454
rect 443382 624218 443414 624454
rect 442794 624134 443414 624218
rect 442794 623898 442826 624134
rect 443062 623898 443146 624134
rect 443382 623898 443414 624134
rect 442794 588454 443414 623898
rect 442794 588218 442826 588454
rect 443062 588218 443146 588454
rect 443382 588218 443414 588454
rect 442794 588134 443414 588218
rect 442794 587898 442826 588134
rect 443062 587898 443146 588134
rect 443382 587898 443414 588134
rect 442794 552454 443414 587898
rect 442794 552218 442826 552454
rect 443062 552218 443146 552454
rect 443382 552218 443414 552454
rect 442794 552134 443414 552218
rect 442794 551898 442826 552134
rect 443062 551898 443146 552134
rect 443382 551898 443414 552134
rect 442794 516454 443414 551898
rect 442794 516218 442826 516454
rect 443062 516218 443146 516454
rect 443382 516218 443414 516454
rect 442794 516134 443414 516218
rect 442794 515898 442826 516134
rect 443062 515898 443146 516134
rect 443382 515898 443414 516134
rect 442794 480454 443414 515898
rect 442794 480218 442826 480454
rect 443062 480218 443146 480454
rect 443382 480218 443414 480454
rect 442794 480134 443414 480218
rect 442794 479898 442826 480134
rect 443062 479898 443146 480134
rect 443382 479898 443414 480134
rect 442794 444454 443414 479898
rect 442794 444218 442826 444454
rect 443062 444218 443146 444454
rect 443382 444218 443414 444454
rect 442794 444134 443414 444218
rect 442794 443898 442826 444134
rect 443062 443898 443146 444134
rect 443382 443898 443414 444134
rect 442794 408454 443414 443898
rect 442794 408218 442826 408454
rect 443062 408218 443146 408454
rect 443382 408218 443414 408454
rect 442794 408134 443414 408218
rect 442794 407898 442826 408134
rect 443062 407898 443146 408134
rect 443382 407898 443414 408134
rect 442794 372454 443414 407898
rect 442794 372218 442826 372454
rect 443062 372218 443146 372454
rect 443382 372218 443414 372454
rect 442794 372134 443414 372218
rect 442794 371898 442826 372134
rect 443062 371898 443146 372134
rect 443382 371898 443414 372134
rect 442794 336454 443414 371898
rect 442794 336218 442826 336454
rect 443062 336218 443146 336454
rect 443382 336218 443414 336454
rect 442794 336134 443414 336218
rect 442794 335898 442826 336134
rect 443062 335898 443146 336134
rect 443382 335898 443414 336134
rect 442794 300454 443414 335898
rect 442794 300218 442826 300454
rect 443062 300218 443146 300454
rect 443382 300218 443414 300454
rect 442794 300134 443414 300218
rect 442794 299898 442826 300134
rect 443062 299898 443146 300134
rect 443382 299898 443414 300134
rect 442794 264454 443414 299898
rect 442794 264218 442826 264454
rect 443062 264218 443146 264454
rect 443382 264218 443414 264454
rect 442794 264134 443414 264218
rect 442794 263898 442826 264134
rect 443062 263898 443146 264134
rect 443382 263898 443414 264134
rect 442794 228454 443414 263898
rect 442794 228218 442826 228454
rect 443062 228218 443146 228454
rect 443382 228218 443414 228454
rect 442794 228134 443414 228218
rect 442794 227898 442826 228134
rect 443062 227898 443146 228134
rect 443382 227898 443414 228134
rect 442794 192454 443414 227898
rect 442794 192218 442826 192454
rect 443062 192218 443146 192454
rect 443382 192218 443414 192454
rect 442794 192134 443414 192218
rect 442794 191898 442826 192134
rect 443062 191898 443146 192134
rect 443382 191898 443414 192134
rect 442794 156454 443414 191898
rect 442794 156218 442826 156454
rect 443062 156218 443146 156454
rect 443382 156218 443414 156454
rect 442794 156134 443414 156218
rect 442794 155898 442826 156134
rect 443062 155898 443146 156134
rect 443382 155898 443414 156134
rect 442794 120454 443414 155898
rect 442794 120218 442826 120454
rect 443062 120218 443146 120454
rect 443382 120218 443414 120454
rect 442794 120134 443414 120218
rect 442794 119898 442826 120134
rect 443062 119898 443146 120134
rect 443382 119898 443414 120134
rect 442794 84454 443414 119898
rect 442794 84218 442826 84454
rect 443062 84218 443146 84454
rect 443382 84218 443414 84454
rect 442794 84134 443414 84218
rect 442794 83898 442826 84134
rect 443062 83898 443146 84134
rect 443382 83898 443414 84134
rect 442794 48454 443414 83898
rect 442794 48218 442826 48454
rect 443062 48218 443146 48454
rect 443382 48218 443414 48454
rect 442794 48134 443414 48218
rect 442794 47898 442826 48134
rect 443062 47898 443146 48134
rect 443382 47898 443414 48134
rect 442794 12454 443414 47898
rect 442794 12218 442826 12454
rect 443062 12218 443146 12454
rect 443382 12218 443414 12454
rect 442794 12134 443414 12218
rect 442794 11898 442826 12134
rect 443062 11898 443146 12134
rect 443382 11898 443414 12134
rect 442794 -2266 443414 11898
rect 442794 -2502 442826 -2266
rect 443062 -2502 443146 -2266
rect 443382 -2502 443414 -2266
rect 442794 -2586 443414 -2502
rect 442794 -2822 442826 -2586
rect 443062 -2822 443146 -2586
rect 443382 -2822 443414 -2586
rect 442794 -7654 443414 -2822
rect 447294 707718 447914 711590
rect 447294 707482 447326 707718
rect 447562 707482 447646 707718
rect 447882 707482 447914 707718
rect 447294 707398 447914 707482
rect 447294 707162 447326 707398
rect 447562 707162 447646 707398
rect 447882 707162 447914 707398
rect 447294 700954 447914 707162
rect 447294 700718 447326 700954
rect 447562 700718 447646 700954
rect 447882 700718 447914 700954
rect 447294 700634 447914 700718
rect 447294 700398 447326 700634
rect 447562 700398 447646 700634
rect 447882 700398 447914 700634
rect 447294 664954 447914 700398
rect 447294 664718 447326 664954
rect 447562 664718 447646 664954
rect 447882 664718 447914 664954
rect 447294 664634 447914 664718
rect 447294 664398 447326 664634
rect 447562 664398 447646 664634
rect 447882 664398 447914 664634
rect 447294 628954 447914 664398
rect 447294 628718 447326 628954
rect 447562 628718 447646 628954
rect 447882 628718 447914 628954
rect 447294 628634 447914 628718
rect 447294 628398 447326 628634
rect 447562 628398 447646 628634
rect 447882 628398 447914 628634
rect 447294 592954 447914 628398
rect 447294 592718 447326 592954
rect 447562 592718 447646 592954
rect 447882 592718 447914 592954
rect 447294 592634 447914 592718
rect 447294 592398 447326 592634
rect 447562 592398 447646 592634
rect 447882 592398 447914 592634
rect 447294 556954 447914 592398
rect 447294 556718 447326 556954
rect 447562 556718 447646 556954
rect 447882 556718 447914 556954
rect 447294 556634 447914 556718
rect 447294 556398 447326 556634
rect 447562 556398 447646 556634
rect 447882 556398 447914 556634
rect 447294 520954 447914 556398
rect 447294 520718 447326 520954
rect 447562 520718 447646 520954
rect 447882 520718 447914 520954
rect 447294 520634 447914 520718
rect 447294 520398 447326 520634
rect 447562 520398 447646 520634
rect 447882 520398 447914 520634
rect 447294 484954 447914 520398
rect 447294 484718 447326 484954
rect 447562 484718 447646 484954
rect 447882 484718 447914 484954
rect 447294 484634 447914 484718
rect 447294 484398 447326 484634
rect 447562 484398 447646 484634
rect 447882 484398 447914 484634
rect 447294 448954 447914 484398
rect 447294 448718 447326 448954
rect 447562 448718 447646 448954
rect 447882 448718 447914 448954
rect 447294 448634 447914 448718
rect 447294 448398 447326 448634
rect 447562 448398 447646 448634
rect 447882 448398 447914 448634
rect 447294 412954 447914 448398
rect 447294 412718 447326 412954
rect 447562 412718 447646 412954
rect 447882 412718 447914 412954
rect 447294 412634 447914 412718
rect 447294 412398 447326 412634
rect 447562 412398 447646 412634
rect 447882 412398 447914 412634
rect 447294 376954 447914 412398
rect 447294 376718 447326 376954
rect 447562 376718 447646 376954
rect 447882 376718 447914 376954
rect 447294 376634 447914 376718
rect 447294 376398 447326 376634
rect 447562 376398 447646 376634
rect 447882 376398 447914 376634
rect 447294 340954 447914 376398
rect 447294 340718 447326 340954
rect 447562 340718 447646 340954
rect 447882 340718 447914 340954
rect 447294 340634 447914 340718
rect 447294 340398 447326 340634
rect 447562 340398 447646 340634
rect 447882 340398 447914 340634
rect 447294 304954 447914 340398
rect 447294 304718 447326 304954
rect 447562 304718 447646 304954
rect 447882 304718 447914 304954
rect 447294 304634 447914 304718
rect 447294 304398 447326 304634
rect 447562 304398 447646 304634
rect 447882 304398 447914 304634
rect 447294 268954 447914 304398
rect 447294 268718 447326 268954
rect 447562 268718 447646 268954
rect 447882 268718 447914 268954
rect 447294 268634 447914 268718
rect 447294 268398 447326 268634
rect 447562 268398 447646 268634
rect 447882 268398 447914 268634
rect 447294 232954 447914 268398
rect 447294 232718 447326 232954
rect 447562 232718 447646 232954
rect 447882 232718 447914 232954
rect 447294 232634 447914 232718
rect 447294 232398 447326 232634
rect 447562 232398 447646 232634
rect 447882 232398 447914 232634
rect 447294 196954 447914 232398
rect 447294 196718 447326 196954
rect 447562 196718 447646 196954
rect 447882 196718 447914 196954
rect 447294 196634 447914 196718
rect 447294 196398 447326 196634
rect 447562 196398 447646 196634
rect 447882 196398 447914 196634
rect 447294 160954 447914 196398
rect 447294 160718 447326 160954
rect 447562 160718 447646 160954
rect 447882 160718 447914 160954
rect 447294 160634 447914 160718
rect 447294 160398 447326 160634
rect 447562 160398 447646 160634
rect 447882 160398 447914 160634
rect 447294 124954 447914 160398
rect 447294 124718 447326 124954
rect 447562 124718 447646 124954
rect 447882 124718 447914 124954
rect 447294 124634 447914 124718
rect 447294 124398 447326 124634
rect 447562 124398 447646 124634
rect 447882 124398 447914 124634
rect 447294 88954 447914 124398
rect 447294 88718 447326 88954
rect 447562 88718 447646 88954
rect 447882 88718 447914 88954
rect 447294 88634 447914 88718
rect 447294 88398 447326 88634
rect 447562 88398 447646 88634
rect 447882 88398 447914 88634
rect 447294 52954 447914 88398
rect 447294 52718 447326 52954
rect 447562 52718 447646 52954
rect 447882 52718 447914 52954
rect 447294 52634 447914 52718
rect 447294 52398 447326 52634
rect 447562 52398 447646 52634
rect 447882 52398 447914 52634
rect 447294 16954 447914 52398
rect 447294 16718 447326 16954
rect 447562 16718 447646 16954
rect 447882 16718 447914 16954
rect 447294 16634 447914 16718
rect 447294 16398 447326 16634
rect 447562 16398 447646 16634
rect 447882 16398 447914 16634
rect 447294 -3226 447914 16398
rect 447294 -3462 447326 -3226
rect 447562 -3462 447646 -3226
rect 447882 -3462 447914 -3226
rect 447294 -3546 447914 -3462
rect 447294 -3782 447326 -3546
rect 447562 -3782 447646 -3546
rect 447882 -3782 447914 -3546
rect 447294 -7654 447914 -3782
rect 451794 708678 452414 711590
rect 451794 708442 451826 708678
rect 452062 708442 452146 708678
rect 452382 708442 452414 708678
rect 451794 708358 452414 708442
rect 451794 708122 451826 708358
rect 452062 708122 452146 708358
rect 452382 708122 452414 708358
rect 451794 669454 452414 708122
rect 451794 669218 451826 669454
rect 452062 669218 452146 669454
rect 452382 669218 452414 669454
rect 451794 669134 452414 669218
rect 451794 668898 451826 669134
rect 452062 668898 452146 669134
rect 452382 668898 452414 669134
rect 451794 633454 452414 668898
rect 451794 633218 451826 633454
rect 452062 633218 452146 633454
rect 452382 633218 452414 633454
rect 451794 633134 452414 633218
rect 451794 632898 451826 633134
rect 452062 632898 452146 633134
rect 452382 632898 452414 633134
rect 451794 597454 452414 632898
rect 451794 597218 451826 597454
rect 452062 597218 452146 597454
rect 452382 597218 452414 597454
rect 451794 597134 452414 597218
rect 451794 596898 451826 597134
rect 452062 596898 452146 597134
rect 452382 596898 452414 597134
rect 451794 561454 452414 596898
rect 451794 561218 451826 561454
rect 452062 561218 452146 561454
rect 452382 561218 452414 561454
rect 451794 561134 452414 561218
rect 451794 560898 451826 561134
rect 452062 560898 452146 561134
rect 452382 560898 452414 561134
rect 451794 525454 452414 560898
rect 451794 525218 451826 525454
rect 452062 525218 452146 525454
rect 452382 525218 452414 525454
rect 451794 525134 452414 525218
rect 451794 524898 451826 525134
rect 452062 524898 452146 525134
rect 452382 524898 452414 525134
rect 451794 489454 452414 524898
rect 451794 489218 451826 489454
rect 452062 489218 452146 489454
rect 452382 489218 452414 489454
rect 451794 489134 452414 489218
rect 451794 488898 451826 489134
rect 452062 488898 452146 489134
rect 452382 488898 452414 489134
rect 451794 453454 452414 488898
rect 451794 453218 451826 453454
rect 452062 453218 452146 453454
rect 452382 453218 452414 453454
rect 451794 453134 452414 453218
rect 451794 452898 451826 453134
rect 452062 452898 452146 453134
rect 452382 452898 452414 453134
rect 451794 417454 452414 452898
rect 451794 417218 451826 417454
rect 452062 417218 452146 417454
rect 452382 417218 452414 417454
rect 451794 417134 452414 417218
rect 451794 416898 451826 417134
rect 452062 416898 452146 417134
rect 452382 416898 452414 417134
rect 451794 381454 452414 416898
rect 451794 381218 451826 381454
rect 452062 381218 452146 381454
rect 452382 381218 452414 381454
rect 451794 381134 452414 381218
rect 451794 380898 451826 381134
rect 452062 380898 452146 381134
rect 452382 380898 452414 381134
rect 451794 345454 452414 380898
rect 451794 345218 451826 345454
rect 452062 345218 452146 345454
rect 452382 345218 452414 345454
rect 451794 345134 452414 345218
rect 451794 344898 451826 345134
rect 452062 344898 452146 345134
rect 452382 344898 452414 345134
rect 451794 309454 452414 344898
rect 451794 309218 451826 309454
rect 452062 309218 452146 309454
rect 452382 309218 452414 309454
rect 451794 309134 452414 309218
rect 451794 308898 451826 309134
rect 452062 308898 452146 309134
rect 452382 308898 452414 309134
rect 451794 273454 452414 308898
rect 451794 273218 451826 273454
rect 452062 273218 452146 273454
rect 452382 273218 452414 273454
rect 451794 273134 452414 273218
rect 451794 272898 451826 273134
rect 452062 272898 452146 273134
rect 452382 272898 452414 273134
rect 451794 237454 452414 272898
rect 451794 237218 451826 237454
rect 452062 237218 452146 237454
rect 452382 237218 452414 237454
rect 451794 237134 452414 237218
rect 451794 236898 451826 237134
rect 452062 236898 452146 237134
rect 452382 236898 452414 237134
rect 451794 201454 452414 236898
rect 451794 201218 451826 201454
rect 452062 201218 452146 201454
rect 452382 201218 452414 201454
rect 451794 201134 452414 201218
rect 451794 200898 451826 201134
rect 452062 200898 452146 201134
rect 452382 200898 452414 201134
rect 451794 165454 452414 200898
rect 451794 165218 451826 165454
rect 452062 165218 452146 165454
rect 452382 165218 452414 165454
rect 451794 165134 452414 165218
rect 451794 164898 451826 165134
rect 452062 164898 452146 165134
rect 452382 164898 452414 165134
rect 451794 129454 452414 164898
rect 451794 129218 451826 129454
rect 452062 129218 452146 129454
rect 452382 129218 452414 129454
rect 451794 129134 452414 129218
rect 451794 128898 451826 129134
rect 452062 128898 452146 129134
rect 452382 128898 452414 129134
rect 451794 93454 452414 128898
rect 451794 93218 451826 93454
rect 452062 93218 452146 93454
rect 452382 93218 452414 93454
rect 451794 93134 452414 93218
rect 451794 92898 451826 93134
rect 452062 92898 452146 93134
rect 452382 92898 452414 93134
rect 451794 57454 452414 92898
rect 451794 57218 451826 57454
rect 452062 57218 452146 57454
rect 452382 57218 452414 57454
rect 451794 57134 452414 57218
rect 451794 56898 451826 57134
rect 452062 56898 452146 57134
rect 452382 56898 452414 57134
rect 451794 21454 452414 56898
rect 451794 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 452414 21454
rect 451794 21134 452414 21218
rect 451794 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 452414 21134
rect 451794 -4186 452414 20898
rect 451794 -4422 451826 -4186
rect 452062 -4422 452146 -4186
rect 452382 -4422 452414 -4186
rect 451794 -4506 452414 -4422
rect 451794 -4742 451826 -4506
rect 452062 -4742 452146 -4506
rect 452382 -4742 452414 -4506
rect 451794 -7654 452414 -4742
rect 456294 709638 456914 711590
rect 456294 709402 456326 709638
rect 456562 709402 456646 709638
rect 456882 709402 456914 709638
rect 456294 709318 456914 709402
rect 456294 709082 456326 709318
rect 456562 709082 456646 709318
rect 456882 709082 456914 709318
rect 456294 673954 456914 709082
rect 456294 673718 456326 673954
rect 456562 673718 456646 673954
rect 456882 673718 456914 673954
rect 456294 673634 456914 673718
rect 456294 673398 456326 673634
rect 456562 673398 456646 673634
rect 456882 673398 456914 673634
rect 456294 637954 456914 673398
rect 456294 637718 456326 637954
rect 456562 637718 456646 637954
rect 456882 637718 456914 637954
rect 456294 637634 456914 637718
rect 456294 637398 456326 637634
rect 456562 637398 456646 637634
rect 456882 637398 456914 637634
rect 456294 601954 456914 637398
rect 456294 601718 456326 601954
rect 456562 601718 456646 601954
rect 456882 601718 456914 601954
rect 456294 601634 456914 601718
rect 456294 601398 456326 601634
rect 456562 601398 456646 601634
rect 456882 601398 456914 601634
rect 456294 565954 456914 601398
rect 456294 565718 456326 565954
rect 456562 565718 456646 565954
rect 456882 565718 456914 565954
rect 456294 565634 456914 565718
rect 456294 565398 456326 565634
rect 456562 565398 456646 565634
rect 456882 565398 456914 565634
rect 456294 529954 456914 565398
rect 456294 529718 456326 529954
rect 456562 529718 456646 529954
rect 456882 529718 456914 529954
rect 456294 529634 456914 529718
rect 456294 529398 456326 529634
rect 456562 529398 456646 529634
rect 456882 529398 456914 529634
rect 456294 493954 456914 529398
rect 456294 493718 456326 493954
rect 456562 493718 456646 493954
rect 456882 493718 456914 493954
rect 456294 493634 456914 493718
rect 456294 493398 456326 493634
rect 456562 493398 456646 493634
rect 456882 493398 456914 493634
rect 456294 457954 456914 493398
rect 456294 457718 456326 457954
rect 456562 457718 456646 457954
rect 456882 457718 456914 457954
rect 456294 457634 456914 457718
rect 456294 457398 456326 457634
rect 456562 457398 456646 457634
rect 456882 457398 456914 457634
rect 456294 421954 456914 457398
rect 456294 421718 456326 421954
rect 456562 421718 456646 421954
rect 456882 421718 456914 421954
rect 456294 421634 456914 421718
rect 456294 421398 456326 421634
rect 456562 421398 456646 421634
rect 456882 421398 456914 421634
rect 456294 385954 456914 421398
rect 456294 385718 456326 385954
rect 456562 385718 456646 385954
rect 456882 385718 456914 385954
rect 456294 385634 456914 385718
rect 456294 385398 456326 385634
rect 456562 385398 456646 385634
rect 456882 385398 456914 385634
rect 456294 349954 456914 385398
rect 456294 349718 456326 349954
rect 456562 349718 456646 349954
rect 456882 349718 456914 349954
rect 456294 349634 456914 349718
rect 456294 349398 456326 349634
rect 456562 349398 456646 349634
rect 456882 349398 456914 349634
rect 456294 313954 456914 349398
rect 456294 313718 456326 313954
rect 456562 313718 456646 313954
rect 456882 313718 456914 313954
rect 456294 313634 456914 313718
rect 456294 313398 456326 313634
rect 456562 313398 456646 313634
rect 456882 313398 456914 313634
rect 456294 277954 456914 313398
rect 456294 277718 456326 277954
rect 456562 277718 456646 277954
rect 456882 277718 456914 277954
rect 456294 277634 456914 277718
rect 456294 277398 456326 277634
rect 456562 277398 456646 277634
rect 456882 277398 456914 277634
rect 456294 241954 456914 277398
rect 456294 241718 456326 241954
rect 456562 241718 456646 241954
rect 456882 241718 456914 241954
rect 456294 241634 456914 241718
rect 456294 241398 456326 241634
rect 456562 241398 456646 241634
rect 456882 241398 456914 241634
rect 456294 205954 456914 241398
rect 456294 205718 456326 205954
rect 456562 205718 456646 205954
rect 456882 205718 456914 205954
rect 456294 205634 456914 205718
rect 456294 205398 456326 205634
rect 456562 205398 456646 205634
rect 456882 205398 456914 205634
rect 456294 169954 456914 205398
rect 456294 169718 456326 169954
rect 456562 169718 456646 169954
rect 456882 169718 456914 169954
rect 456294 169634 456914 169718
rect 456294 169398 456326 169634
rect 456562 169398 456646 169634
rect 456882 169398 456914 169634
rect 456294 133954 456914 169398
rect 456294 133718 456326 133954
rect 456562 133718 456646 133954
rect 456882 133718 456914 133954
rect 456294 133634 456914 133718
rect 456294 133398 456326 133634
rect 456562 133398 456646 133634
rect 456882 133398 456914 133634
rect 456294 97954 456914 133398
rect 456294 97718 456326 97954
rect 456562 97718 456646 97954
rect 456882 97718 456914 97954
rect 456294 97634 456914 97718
rect 456294 97398 456326 97634
rect 456562 97398 456646 97634
rect 456882 97398 456914 97634
rect 456294 61954 456914 97398
rect 456294 61718 456326 61954
rect 456562 61718 456646 61954
rect 456882 61718 456914 61954
rect 456294 61634 456914 61718
rect 456294 61398 456326 61634
rect 456562 61398 456646 61634
rect 456882 61398 456914 61634
rect 456294 25954 456914 61398
rect 456294 25718 456326 25954
rect 456562 25718 456646 25954
rect 456882 25718 456914 25954
rect 456294 25634 456914 25718
rect 456294 25398 456326 25634
rect 456562 25398 456646 25634
rect 456882 25398 456914 25634
rect 456294 -5146 456914 25398
rect 456294 -5382 456326 -5146
rect 456562 -5382 456646 -5146
rect 456882 -5382 456914 -5146
rect 456294 -5466 456914 -5382
rect 456294 -5702 456326 -5466
rect 456562 -5702 456646 -5466
rect 456882 -5702 456914 -5466
rect 456294 -7654 456914 -5702
rect 460794 710598 461414 711590
rect 460794 710362 460826 710598
rect 461062 710362 461146 710598
rect 461382 710362 461414 710598
rect 460794 710278 461414 710362
rect 460794 710042 460826 710278
rect 461062 710042 461146 710278
rect 461382 710042 461414 710278
rect 460794 678454 461414 710042
rect 460794 678218 460826 678454
rect 461062 678218 461146 678454
rect 461382 678218 461414 678454
rect 460794 678134 461414 678218
rect 460794 677898 460826 678134
rect 461062 677898 461146 678134
rect 461382 677898 461414 678134
rect 460794 642454 461414 677898
rect 460794 642218 460826 642454
rect 461062 642218 461146 642454
rect 461382 642218 461414 642454
rect 460794 642134 461414 642218
rect 460794 641898 460826 642134
rect 461062 641898 461146 642134
rect 461382 641898 461414 642134
rect 460794 606454 461414 641898
rect 460794 606218 460826 606454
rect 461062 606218 461146 606454
rect 461382 606218 461414 606454
rect 460794 606134 461414 606218
rect 460794 605898 460826 606134
rect 461062 605898 461146 606134
rect 461382 605898 461414 606134
rect 460794 570454 461414 605898
rect 460794 570218 460826 570454
rect 461062 570218 461146 570454
rect 461382 570218 461414 570454
rect 460794 570134 461414 570218
rect 460794 569898 460826 570134
rect 461062 569898 461146 570134
rect 461382 569898 461414 570134
rect 460794 534454 461414 569898
rect 460794 534218 460826 534454
rect 461062 534218 461146 534454
rect 461382 534218 461414 534454
rect 460794 534134 461414 534218
rect 460794 533898 460826 534134
rect 461062 533898 461146 534134
rect 461382 533898 461414 534134
rect 460794 498454 461414 533898
rect 460794 498218 460826 498454
rect 461062 498218 461146 498454
rect 461382 498218 461414 498454
rect 460794 498134 461414 498218
rect 460794 497898 460826 498134
rect 461062 497898 461146 498134
rect 461382 497898 461414 498134
rect 460794 462454 461414 497898
rect 460794 462218 460826 462454
rect 461062 462218 461146 462454
rect 461382 462218 461414 462454
rect 460794 462134 461414 462218
rect 460794 461898 460826 462134
rect 461062 461898 461146 462134
rect 461382 461898 461414 462134
rect 460794 426454 461414 461898
rect 460794 426218 460826 426454
rect 461062 426218 461146 426454
rect 461382 426218 461414 426454
rect 460794 426134 461414 426218
rect 460794 425898 460826 426134
rect 461062 425898 461146 426134
rect 461382 425898 461414 426134
rect 460794 390454 461414 425898
rect 460794 390218 460826 390454
rect 461062 390218 461146 390454
rect 461382 390218 461414 390454
rect 460794 390134 461414 390218
rect 460794 389898 460826 390134
rect 461062 389898 461146 390134
rect 461382 389898 461414 390134
rect 460794 354454 461414 389898
rect 460794 354218 460826 354454
rect 461062 354218 461146 354454
rect 461382 354218 461414 354454
rect 460794 354134 461414 354218
rect 460794 353898 460826 354134
rect 461062 353898 461146 354134
rect 461382 353898 461414 354134
rect 460794 318454 461414 353898
rect 460794 318218 460826 318454
rect 461062 318218 461146 318454
rect 461382 318218 461414 318454
rect 460794 318134 461414 318218
rect 460794 317898 460826 318134
rect 461062 317898 461146 318134
rect 461382 317898 461414 318134
rect 460794 282454 461414 317898
rect 460794 282218 460826 282454
rect 461062 282218 461146 282454
rect 461382 282218 461414 282454
rect 460794 282134 461414 282218
rect 460794 281898 460826 282134
rect 461062 281898 461146 282134
rect 461382 281898 461414 282134
rect 460794 246454 461414 281898
rect 460794 246218 460826 246454
rect 461062 246218 461146 246454
rect 461382 246218 461414 246454
rect 460794 246134 461414 246218
rect 460794 245898 460826 246134
rect 461062 245898 461146 246134
rect 461382 245898 461414 246134
rect 460794 210454 461414 245898
rect 460794 210218 460826 210454
rect 461062 210218 461146 210454
rect 461382 210218 461414 210454
rect 460794 210134 461414 210218
rect 460794 209898 460826 210134
rect 461062 209898 461146 210134
rect 461382 209898 461414 210134
rect 460794 174454 461414 209898
rect 460794 174218 460826 174454
rect 461062 174218 461146 174454
rect 461382 174218 461414 174454
rect 460794 174134 461414 174218
rect 460794 173898 460826 174134
rect 461062 173898 461146 174134
rect 461382 173898 461414 174134
rect 460794 138454 461414 173898
rect 460794 138218 460826 138454
rect 461062 138218 461146 138454
rect 461382 138218 461414 138454
rect 460794 138134 461414 138218
rect 460794 137898 460826 138134
rect 461062 137898 461146 138134
rect 461382 137898 461414 138134
rect 460794 102454 461414 137898
rect 460794 102218 460826 102454
rect 461062 102218 461146 102454
rect 461382 102218 461414 102454
rect 460794 102134 461414 102218
rect 460794 101898 460826 102134
rect 461062 101898 461146 102134
rect 461382 101898 461414 102134
rect 460794 66454 461414 101898
rect 460794 66218 460826 66454
rect 461062 66218 461146 66454
rect 461382 66218 461414 66454
rect 460794 66134 461414 66218
rect 460794 65898 460826 66134
rect 461062 65898 461146 66134
rect 461382 65898 461414 66134
rect 460794 30454 461414 65898
rect 460794 30218 460826 30454
rect 461062 30218 461146 30454
rect 461382 30218 461414 30454
rect 460794 30134 461414 30218
rect 460794 29898 460826 30134
rect 461062 29898 461146 30134
rect 461382 29898 461414 30134
rect 460794 -6106 461414 29898
rect 460794 -6342 460826 -6106
rect 461062 -6342 461146 -6106
rect 461382 -6342 461414 -6106
rect 460794 -6426 461414 -6342
rect 460794 -6662 460826 -6426
rect 461062 -6662 461146 -6426
rect 461382 -6662 461414 -6426
rect 460794 -7654 461414 -6662
rect 465294 711558 465914 711590
rect 465294 711322 465326 711558
rect 465562 711322 465646 711558
rect 465882 711322 465914 711558
rect 465294 711238 465914 711322
rect 465294 711002 465326 711238
rect 465562 711002 465646 711238
rect 465882 711002 465914 711238
rect 465294 682954 465914 711002
rect 465294 682718 465326 682954
rect 465562 682718 465646 682954
rect 465882 682718 465914 682954
rect 465294 682634 465914 682718
rect 465294 682398 465326 682634
rect 465562 682398 465646 682634
rect 465882 682398 465914 682634
rect 465294 646954 465914 682398
rect 465294 646718 465326 646954
rect 465562 646718 465646 646954
rect 465882 646718 465914 646954
rect 465294 646634 465914 646718
rect 465294 646398 465326 646634
rect 465562 646398 465646 646634
rect 465882 646398 465914 646634
rect 465294 610954 465914 646398
rect 465294 610718 465326 610954
rect 465562 610718 465646 610954
rect 465882 610718 465914 610954
rect 465294 610634 465914 610718
rect 465294 610398 465326 610634
rect 465562 610398 465646 610634
rect 465882 610398 465914 610634
rect 465294 574954 465914 610398
rect 465294 574718 465326 574954
rect 465562 574718 465646 574954
rect 465882 574718 465914 574954
rect 465294 574634 465914 574718
rect 465294 574398 465326 574634
rect 465562 574398 465646 574634
rect 465882 574398 465914 574634
rect 465294 538954 465914 574398
rect 465294 538718 465326 538954
rect 465562 538718 465646 538954
rect 465882 538718 465914 538954
rect 465294 538634 465914 538718
rect 465294 538398 465326 538634
rect 465562 538398 465646 538634
rect 465882 538398 465914 538634
rect 465294 502954 465914 538398
rect 465294 502718 465326 502954
rect 465562 502718 465646 502954
rect 465882 502718 465914 502954
rect 465294 502634 465914 502718
rect 465294 502398 465326 502634
rect 465562 502398 465646 502634
rect 465882 502398 465914 502634
rect 465294 466954 465914 502398
rect 465294 466718 465326 466954
rect 465562 466718 465646 466954
rect 465882 466718 465914 466954
rect 465294 466634 465914 466718
rect 465294 466398 465326 466634
rect 465562 466398 465646 466634
rect 465882 466398 465914 466634
rect 465294 430954 465914 466398
rect 465294 430718 465326 430954
rect 465562 430718 465646 430954
rect 465882 430718 465914 430954
rect 465294 430634 465914 430718
rect 465294 430398 465326 430634
rect 465562 430398 465646 430634
rect 465882 430398 465914 430634
rect 465294 394954 465914 430398
rect 465294 394718 465326 394954
rect 465562 394718 465646 394954
rect 465882 394718 465914 394954
rect 465294 394634 465914 394718
rect 465294 394398 465326 394634
rect 465562 394398 465646 394634
rect 465882 394398 465914 394634
rect 465294 358954 465914 394398
rect 465294 358718 465326 358954
rect 465562 358718 465646 358954
rect 465882 358718 465914 358954
rect 465294 358634 465914 358718
rect 465294 358398 465326 358634
rect 465562 358398 465646 358634
rect 465882 358398 465914 358634
rect 465294 322954 465914 358398
rect 465294 322718 465326 322954
rect 465562 322718 465646 322954
rect 465882 322718 465914 322954
rect 465294 322634 465914 322718
rect 465294 322398 465326 322634
rect 465562 322398 465646 322634
rect 465882 322398 465914 322634
rect 465294 286954 465914 322398
rect 465294 286718 465326 286954
rect 465562 286718 465646 286954
rect 465882 286718 465914 286954
rect 465294 286634 465914 286718
rect 465294 286398 465326 286634
rect 465562 286398 465646 286634
rect 465882 286398 465914 286634
rect 465294 250954 465914 286398
rect 465294 250718 465326 250954
rect 465562 250718 465646 250954
rect 465882 250718 465914 250954
rect 465294 250634 465914 250718
rect 465294 250398 465326 250634
rect 465562 250398 465646 250634
rect 465882 250398 465914 250634
rect 465294 214954 465914 250398
rect 465294 214718 465326 214954
rect 465562 214718 465646 214954
rect 465882 214718 465914 214954
rect 465294 214634 465914 214718
rect 465294 214398 465326 214634
rect 465562 214398 465646 214634
rect 465882 214398 465914 214634
rect 465294 178954 465914 214398
rect 465294 178718 465326 178954
rect 465562 178718 465646 178954
rect 465882 178718 465914 178954
rect 465294 178634 465914 178718
rect 465294 178398 465326 178634
rect 465562 178398 465646 178634
rect 465882 178398 465914 178634
rect 465294 142954 465914 178398
rect 465294 142718 465326 142954
rect 465562 142718 465646 142954
rect 465882 142718 465914 142954
rect 465294 142634 465914 142718
rect 465294 142398 465326 142634
rect 465562 142398 465646 142634
rect 465882 142398 465914 142634
rect 465294 106954 465914 142398
rect 465294 106718 465326 106954
rect 465562 106718 465646 106954
rect 465882 106718 465914 106954
rect 465294 106634 465914 106718
rect 465294 106398 465326 106634
rect 465562 106398 465646 106634
rect 465882 106398 465914 106634
rect 465294 70954 465914 106398
rect 465294 70718 465326 70954
rect 465562 70718 465646 70954
rect 465882 70718 465914 70954
rect 465294 70634 465914 70718
rect 465294 70398 465326 70634
rect 465562 70398 465646 70634
rect 465882 70398 465914 70634
rect 465294 34954 465914 70398
rect 465294 34718 465326 34954
rect 465562 34718 465646 34954
rect 465882 34718 465914 34954
rect 465294 34634 465914 34718
rect 465294 34398 465326 34634
rect 465562 34398 465646 34634
rect 465882 34398 465914 34634
rect 465294 -7066 465914 34398
rect 465294 -7302 465326 -7066
rect 465562 -7302 465646 -7066
rect 465882 -7302 465914 -7066
rect 465294 -7386 465914 -7302
rect 465294 -7622 465326 -7386
rect 465562 -7622 465646 -7386
rect 465882 -7622 465914 -7386
rect 465294 -7654 465914 -7622
rect 469794 704838 470414 711590
rect 469794 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 470414 704838
rect 469794 704518 470414 704602
rect 469794 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 470414 704518
rect 469794 687454 470414 704282
rect 469794 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 470414 687454
rect 469794 687134 470414 687218
rect 469794 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 470414 687134
rect 469794 651454 470414 686898
rect 469794 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 470414 651454
rect 469794 651134 470414 651218
rect 469794 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 470414 651134
rect 469794 615454 470414 650898
rect 469794 615218 469826 615454
rect 470062 615218 470146 615454
rect 470382 615218 470414 615454
rect 469794 615134 470414 615218
rect 469794 614898 469826 615134
rect 470062 614898 470146 615134
rect 470382 614898 470414 615134
rect 469794 579454 470414 614898
rect 469794 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 470414 579454
rect 469794 579134 470414 579218
rect 469794 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 470414 579134
rect 469794 543454 470414 578898
rect 469794 543218 469826 543454
rect 470062 543218 470146 543454
rect 470382 543218 470414 543454
rect 469794 543134 470414 543218
rect 469794 542898 469826 543134
rect 470062 542898 470146 543134
rect 470382 542898 470414 543134
rect 469794 507454 470414 542898
rect 469794 507218 469826 507454
rect 470062 507218 470146 507454
rect 470382 507218 470414 507454
rect 469794 507134 470414 507218
rect 469794 506898 469826 507134
rect 470062 506898 470146 507134
rect 470382 506898 470414 507134
rect 469794 471454 470414 506898
rect 469794 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 470414 471454
rect 469794 471134 470414 471218
rect 469794 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 470414 471134
rect 469794 435454 470414 470898
rect 469794 435218 469826 435454
rect 470062 435218 470146 435454
rect 470382 435218 470414 435454
rect 469794 435134 470414 435218
rect 469794 434898 469826 435134
rect 470062 434898 470146 435134
rect 470382 434898 470414 435134
rect 469794 399454 470414 434898
rect 469794 399218 469826 399454
rect 470062 399218 470146 399454
rect 470382 399218 470414 399454
rect 469794 399134 470414 399218
rect 469794 398898 469826 399134
rect 470062 398898 470146 399134
rect 470382 398898 470414 399134
rect 469794 363454 470414 398898
rect 469794 363218 469826 363454
rect 470062 363218 470146 363454
rect 470382 363218 470414 363454
rect 469794 363134 470414 363218
rect 469794 362898 469826 363134
rect 470062 362898 470146 363134
rect 470382 362898 470414 363134
rect 469794 327454 470414 362898
rect 469794 327218 469826 327454
rect 470062 327218 470146 327454
rect 470382 327218 470414 327454
rect 469794 327134 470414 327218
rect 469794 326898 469826 327134
rect 470062 326898 470146 327134
rect 470382 326898 470414 327134
rect 469794 291454 470414 326898
rect 469794 291218 469826 291454
rect 470062 291218 470146 291454
rect 470382 291218 470414 291454
rect 469794 291134 470414 291218
rect 469794 290898 469826 291134
rect 470062 290898 470146 291134
rect 470382 290898 470414 291134
rect 469794 255454 470414 290898
rect 469794 255218 469826 255454
rect 470062 255218 470146 255454
rect 470382 255218 470414 255454
rect 469794 255134 470414 255218
rect 469794 254898 469826 255134
rect 470062 254898 470146 255134
rect 470382 254898 470414 255134
rect 469794 219454 470414 254898
rect 469794 219218 469826 219454
rect 470062 219218 470146 219454
rect 470382 219218 470414 219454
rect 469794 219134 470414 219218
rect 469794 218898 469826 219134
rect 470062 218898 470146 219134
rect 470382 218898 470414 219134
rect 469794 183454 470414 218898
rect 469794 183218 469826 183454
rect 470062 183218 470146 183454
rect 470382 183218 470414 183454
rect 469794 183134 470414 183218
rect 469794 182898 469826 183134
rect 470062 182898 470146 183134
rect 470382 182898 470414 183134
rect 469794 147454 470414 182898
rect 469794 147218 469826 147454
rect 470062 147218 470146 147454
rect 470382 147218 470414 147454
rect 469794 147134 470414 147218
rect 469794 146898 469826 147134
rect 470062 146898 470146 147134
rect 470382 146898 470414 147134
rect 469794 111454 470414 146898
rect 469794 111218 469826 111454
rect 470062 111218 470146 111454
rect 470382 111218 470414 111454
rect 469794 111134 470414 111218
rect 469794 110898 469826 111134
rect 470062 110898 470146 111134
rect 470382 110898 470414 111134
rect 469794 75454 470414 110898
rect 469794 75218 469826 75454
rect 470062 75218 470146 75454
rect 470382 75218 470414 75454
rect 469794 75134 470414 75218
rect 469794 74898 469826 75134
rect 470062 74898 470146 75134
rect 470382 74898 470414 75134
rect 469794 39454 470414 74898
rect 469794 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 470414 39454
rect 469794 39134 470414 39218
rect 469794 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 470414 39134
rect 469794 3454 470414 38898
rect 469794 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 470414 3454
rect 469794 3134 470414 3218
rect 469794 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 470414 3134
rect 469794 -346 470414 2898
rect 469794 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 470414 -346
rect 469794 -666 470414 -582
rect 469794 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 470414 -666
rect 469794 -7654 470414 -902
rect 474294 705798 474914 711590
rect 474294 705562 474326 705798
rect 474562 705562 474646 705798
rect 474882 705562 474914 705798
rect 474294 705478 474914 705562
rect 474294 705242 474326 705478
rect 474562 705242 474646 705478
rect 474882 705242 474914 705478
rect 474294 691954 474914 705242
rect 474294 691718 474326 691954
rect 474562 691718 474646 691954
rect 474882 691718 474914 691954
rect 474294 691634 474914 691718
rect 474294 691398 474326 691634
rect 474562 691398 474646 691634
rect 474882 691398 474914 691634
rect 474294 655954 474914 691398
rect 474294 655718 474326 655954
rect 474562 655718 474646 655954
rect 474882 655718 474914 655954
rect 474294 655634 474914 655718
rect 474294 655398 474326 655634
rect 474562 655398 474646 655634
rect 474882 655398 474914 655634
rect 474294 619954 474914 655398
rect 474294 619718 474326 619954
rect 474562 619718 474646 619954
rect 474882 619718 474914 619954
rect 474294 619634 474914 619718
rect 474294 619398 474326 619634
rect 474562 619398 474646 619634
rect 474882 619398 474914 619634
rect 474294 583954 474914 619398
rect 474294 583718 474326 583954
rect 474562 583718 474646 583954
rect 474882 583718 474914 583954
rect 474294 583634 474914 583718
rect 474294 583398 474326 583634
rect 474562 583398 474646 583634
rect 474882 583398 474914 583634
rect 474294 547954 474914 583398
rect 474294 547718 474326 547954
rect 474562 547718 474646 547954
rect 474882 547718 474914 547954
rect 474294 547634 474914 547718
rect 474294 547398 474326 547634
rect 474562 547398 474646 547634
rect 474882 547398 474914 547634
rect 474294 511954 474914 547398
rect 474294 511718 474326 511954
rect 474562 511718 474646 511954
rect 474882 511718 474914 511954
rect 474294 511634 474914 511718
rect 474294 511398 474326 511634
rect 474562 511398 474646 511634
rect 474882 511398 474914 511634
rect 474294 475954 474914 511398
rect 474294 475718 474326 475954
rect 474562 475718 474646 475954
rect 474882 475718 474914 475954
rect 474294 475634 474914 475718
rect 474294 475398 474326 475634
rect 474562 475398 474646 475634
rect 474882 475398 474914 475634
rect 474294 439954 474914 475398
rect 474294 439718 474326 439954
rect 474562 439718 474646 439954
rect 474882 439718 474914 439954
rect 474294 439634 474914 439718
rect 474294 439398 474326 439634
rect 474562 439398 474646 439634
rect 474882 439398 474914 439634
rect 474294 403954 474914 439398
rect 474294 403718 474326 403954
rect 474562 403718 474646 403954
rect 474882 403718 474914 403954
rect 474294 403634 474914 403718
rect 474294 403398 474326 403634
rect 474562 403398 474646 403634
rect 474882 403398 474914 403634
rect 474294 367954 474914 403398
rect 474294 367718 474326 367954
rect 474562 367718 474646 367954
rect 474882 367718 474914 367954
rect 474294 367634 474914 367718
rect 474294 367398 474326 367634
rect 474562 367398 474646 367634
rect 474882 367398 474914 367634
rect 474294 331954 474914 367398
rect 474294 331718 474326 331954
rect 474562 331718 474646 331954
rect 474882 331718 474914 331954
rect 474294 331634 474914 331718
rect 474294 331398 474326 331634
rect 474562 331398 474646 331634
rect 474882 331398 474914 331634
rect 474294 295954 474914 331398
rect 474294 295718 474326 295954
rect 474562 295718 474646 295954
rect 474882 295718 474914 295954
rect 474294 295634 474914 295718
rect 474294 295398 474326 295634
rect 474562 295398 474646 295634
rect 474882 295398 474914 295634
rect 474294 259954 474914 295398
rect 474294 259718 474326 259954
rect 474562 259718 474646 259954
rect 474882 259718 474914 259954
rect 474294 259634 474914 259718
rect 474294 259398 474326 259634
rect 474562 259398 474646 259634
rect 474882 259398 474914 259634
rect 474294 223954 474914 259398
rect 474294 223718 474326 223954
rect 474562 223718 474646 223954
rect 474882 223718 474914 223954
rect 474294 223634 474914 223718
rect 474294 223398 474326 223634
rect 474562 223398 474646 223634
rect 474882 223398 474914 223634
rect 474294 187954 474914 223398
rect 474294 187718 474326 187954
rect 474562 187718 474646 187954
rect 474882 187718 474914 187954
rect 474294 187634 474914 187718
rect 474294 187398 474326 187634
rect 474562 187398 474646 187634
rect 474882 187398 474914 187634
rect 474294 151954 474914 187398
rect 474294 151718 474326 151954
rect 474562 151718 474646 151954
rect 474882 151718 474914 151954
rect 474294 151634 474914 151718
rect 474294 151398 474326 151634
rect 474562 151398 474646 151634
rect 474882 151398 474914 151634
rect 474294 115954 474914 151398
rect 474294 115718 474326 115954
rect 474562 115718 474646 115954
rect 474882 115718 474914 115954
rect 474294 115634 474914 115718
rect 474294 115398 474326 115634
rect 474562 115398 474646 115634
rect 474882 115398 474914 115634
rect 474294 79954 474914 115398
rect 474294 79718 474326 79954
rect 474562 79718 474646 79954
rect 474882 79718 474914 79954
rect 474294 79634 474914 79718
rect 474294 79398 474326 79634
rect 474562 79398 474646 79634
rect 474882 79398 474914 79634
rect 474294 43954 474914 79398
rect 474294 43718 474326 43954
rect 474562 43718 474646 43954
rect 474882 43718 474914 43954
rect 474294 43634 474914 43718
rect 474294 43398 474326 43634
rect 474562 43398 474646 43634
rect 474882 43398 474914 43634
rect 474294 7954 474914 43398
rect 474294 7718 474326 7954
rect 474562 7718 474646 7954
rect 474882 7718 474914 7954
rect 474294 7634 474914 7718
rect 474294 7398 474326 7634
rect 474562 7398 474646 7634
rect 474882 7398 474914 7634
rect 474294 -1306 474914 7398
rect 474294 -1542 474326 -1306
rect 474562 -1542 474646 -1306
rect 474882 -1542 474914 -1306
rect 474294 -1626 474914 -1542
rect 474294 -1862 474326 -1626
rect 474562 -1862 474646 -1626
rect 474882 -1862 474914 -1626
rect 474294 -7654 474914 -1862
rect 478794 706758 479414 711590
rect 478794 706522 478826 706758
rect 479062 706522 479146 706758
rect 479382 706522 479414 706758
rect 478794 706438 479414 706522
rect 478794 706202 478826 706438
rect 479062 706202 479146 706438
rect 479382 706202 479414 706438
rect 478794 696454 479414 706202
rect 478794 696218 478826 696454
rect 479062 696218 479146 696454
rect 479382 696218 479414 696454
rect 478794 696134 479414 696218
rect 478794 695898 478826 696134
rect 479062 695898 479146 696134
rect 479382 695898 479414 696134
rect 478794 660454 479414 695898
rect 478794 660218 478826 660454
rect 479062 660218 479146 660454
rect 479382 660218 479414 660454
rect 478794 660134 479414 660218
rect 478794 659898 478826 660134
rect 479062 659898 479146 660134
rect 479382 659898 479414 660134
rect 478794 624454 479414 659898
rect 478794 624218 478826 624454
rect 479062 624218 479146 624454
rect 479382 624218 479414 624454
rect 478794 624134 479414 624218
rect 478794 623898 478826 624134
rect 479062 623898 479146 624134
rect 479382 623898 479414 624134
rect 478794 588454 479414 623898
rect 478794 588218 478826 588454
rect 479062 588218 479146 588454
rect 479382 588218 479414 588454
rect 478794 588134 479414 588218
rect 478794 587898 478826 588134
rect 479062 587898 479146 588134
rect 479382 587898 479414 588134
rect 478794 552454 479414 587898
rect 478794 552218 478826 552454
rect 479062 552218 479146 552454
rect 479382 552218 479414 552454
rect 478794 552134 479414 552218
rect 478794 551898 478826 552134
rect 479062 551898 479146 552134
rect 479382 551898 479414 552134
rect 478794 516454 479414 551898
rect 478794 516218 478826 516454
rect 479062 516218 479146 516454
rect 479382 516218 479414 516454
rect 478794 516134 479414 516218
rect 478794 515898 478826 516134
rect 479062 515898 479146 516134
rect 479382 515898 479414 516134
rect 478794 480454 479414 515898
rect 478794 480218 478826 480454
rect 479062 480218 479146 480454
rect 479382 480218 479414 480454
rect 478794 480134 479414 480218
rect 478794 479898 478826 480134
rect 479062 479898 479146 480134
rect 479382 479898 479414 480134
rect 478794 444454 479414 479898
rect 478794 444218 478826 444454
rect 479062 444218 479146 444454
rect 479382 444218 479414 444454
rect 478794 444134 479414 444218
rect 478794 443898 478826 444134
rect 479062 443898 479146 444134
rect 479382 443898 479414 444134
rect 478794 408454 479414 443898
rect 478794 408218 478826 408454
rect 479062 408218 479146 408454
rect 479382 408218 479414 408454
rect 478794 408134 479414 408218
rect 478794 407898 478826 408134
rect 479062 407898 479146 408134
rect 479382 407898 479414 408134
rect 478794 372454 479414 407898
rect 478794 372218 478826 372454
rect 479062 372218 479146 372454
rect 479382 372218 479414 372454
rect 478794 372134 479414 372218
rect 478794 371898 478826 372134
rect 479062 371898 479146 372134
rect 479382 371898 479414 372134
rect 478794 336454 479414 371898
rect 478794 336218 478826 336454
rect 479062 336218 479146 336454
rect 479382 336218 479414 336454
rect 478794 336134 479414 336218
rect 478794 335898 478826 336134
rect 479062 335898 479146 336134
rect 479382 335898 479414 336134
rect 478794 300454 479414 335898
rect 478794 300218 478826 300454
rect 479062 300218 479146 300454
rect 479382 300218 479414 300454
rect 478794 300134 479414 300218
rect 478794 299898 478826 300134
rect 479062 299898 479146 300134
rect 479382 299898 479414 300134
rect 478794 264454 479414 299898
rect 478794 264218 478826 264454
rect 479062 264218 479146 264454
rect 479382 264218 479414 264454
rect 478794 264134 479414 264218
rect 478794 263898 478826 264134
rect 479062 263898 479146 264134
rect 479382 263898 479414 264134
rect 478794 228454 479414 263898
rect 478794 228218 478826 228454
rect 479062 228218 479146 228454
rect 479382 228218 479414 228454
rect 478794 228134 479414 228218
rect 478794 227898 478826 228134
rect 479062 227898 479146 228134
rect 479382 227898 479414 228134
rect 478794 192454 479414 227898
rect 478794 192218 478826 192454
rect 479062 192218 479146 192454
rect 479382 192218 479414 192454
rect 478794 192134 479414 192218
rect 478794 191898 478826 192134
rect 479062 191898 479146 192134
rect 479382 191898 479414 192134
rect 478794 156454 479414 191898
rect 478794 156218 478826 156454
rect 479062 156218 479146 156454
rect 479382 156218 479414 156454
rect 478794 156134 479414 156218
rect 478794 155898 478826 156134
rect 479062 155898 479146 156134
rect 479382 155898 479414 156134
rect 478794 120454 479414 155898
rect 478794 120218 478826 120454
rect 479062 120218 479146 120454
rect 479382 120218 479414 120454
rect 478794 120134 479414 120218
rect 478794 119898 478826 120134
rect 479062 119898 479146 120134
rect 479382 119898 479414 120134
rect 478794 84454 479414 119898
rect 478794 84218 478826 84454
rect 479062 84218 479146 84454
rect 479382 84218 479414 84454
rect 478794 84134 479414 84218
rect 478794 83898 478826 84134
rect 479062 83898 479146 84134
rect 479382 83898 479414 84134
rect 478794 48454 479414 83898
rect 478794 48218 478826 48454
rect 479062 48218 479146 48454
rect 479382 48218 479414 48454
rect 478794 48134 479414 48218
rect 478794 47898 478826 48134
rect 479062 47898 479146 48134
rect 479382 47898 479414 48134
rect 478794 12454 479414 47898
rect 478794 12218 478826 12454
rect 479062 12218 479146 12454
rect 479382 12218 479414 12454
rect 478794 12134 479414 12218
rect 478794 11898 478826 12134
rect 479062 11898 479146 12134
rect 479382 11898 479414 12134
rect 478794 -2266 479414 11898
rect 478794 -2502 478826 -2266
rect 479062 -2502 479146 -2266
rect 479382 -2502 479414 -2266
rect 478794 -2586 479414 -2502
rect 478794 -2822 478826 -2586
rect 479062 -2822 479146 -2586
rect 479382 -2822 479414 -2586
rect 478794 -7654 479414 -2822
rect 483294 707718 483914 711590
rect 483294 707482 483326 707718
rect 483562 707482 483646 707718
rect 483882 707482 483914 707718
rect 483294 707398 483914 707482
rect 483294 707162 483326 707398
rect 483562 707162 483646 707398
rect 483882 707162 483914 707398
rect 483294 700954 483914 707162
rect 483294 700718 483326 700954
rect 483562 700718 483646 700954
rect 483882 700718 483914 700954
rect 483294 700634 483914 700718
rect 483294 700398 483326 700634
rect 483562 700398 483646 700634
rect 483882 700398 483914 700634
rect 483294 664954 483914 700398
rect 483294 664718 483326 664954
rect 483562 664718 483646 664954
rect 483882 664718 483914 664954
rect 483294 664634 483914 664718
rect 483294 664398 483326 664634
rect 483562 664398 483646 664634
rect 483882 664398 483914 664634
rect 483294 628954 483914 664398
rect 483294 628718 483326 628954
rect 483562 628718 483646 628954
rect 483882 628718 483914 628954
rect 483294 628634 483914 628718
rect 483294 628398 483326 628634
rect 483562 628398 483646 628634
rect 483882 628398 483914 628634
rect 483294 592954 483914 628398
rect 483294 592718 483326 592954
rect 483562 592718 483646 592954
rect 483882 592718 483914 592954
rect 483294 592634 483914 592718
rect 483294 592398 483326 592634
rect 483562 592398 483646 592634
rect 483882 592398 483914 592634
rect 483294 556954 483914 592398
rect 483294 556718 483326 556954
rect 483562 556718 483646 556954
rect 483882 556718 483914 556954
rect 483294 556634 483914 556718
rect 483294 556398 483326 556634
rect 483562 556398 483646 556634
rect 483882 556398 483914 556634
rect 483294 520954 483914 556398
rect 483294 520718 483326 520954
rect 483562 520718 483646 520954
rect 483882 520718 483914 520954
rect 483294 520634 483914 520718
rect 483294 520398 483326 520634
rect 483562 520398 483646 520634
rect 483882 520398 483914 520634
rect 483294 484954 483914 520398
rect 483294 484718 483326 484954
rect 483562 484718 483646 484954
rect 483882 484718 483914 484954
rect 483294 484634 483914 484718
rect 483294 484398 483326 484634
rect 483562 484398 483646 484634
rect 483882 484398 483914 484634
rect 483294 448954 483914 484398
rect 483294 448718 483326 448954
rect 483562 448718 483646 448954
rect 483882 448718 483914 448954
rect 483294 448634 483914 448718
rect 483294 448398 483326 448634
rect 483562 448398 483646 448634
rect 483882 448398 483914 448634
rect 483294 412954 483914 448398
rect 483294 412718 483326 412954
rect 483562 412718 483646 412954
rect 483882 412718 483914 412954
rect 483294 412634 483914 412718
rect 483294 412398 483326 412634
rect 483562 412398 483646 412634
rect 483882 412398 483914 412634
rect 483294 376954 483914 412398
rect 483294 376718 483326 376954
rect 483562 376718 483646 376954
rect 483882 376718 483914 376954
rect 483294 376634 483914 376718
rect 483294 376398 483326 376634
rect 483562 376398 483646 376634
rect 483882 376398 483914 376634
rect 483294 340954 483914 376398
rect 483294 340718 483326 340954
rect 483562 340718 483646 340954
rect 483882 340718 483914 340954
rect 483294 340634 483914 340718
rect 483294 340398 483326 340634
rect 483562 340398 483646 340634
rect 483882 340398 483914 340634
rect 483294 304954 483914 340398
rect 483294 304718 483326 304954
rect 483562 304718 483646 304954
rect 483882 304718 483914 304954
rect 483294 304634 483914 304718
rect 483294 304398 483326 304634
rect 483562 304398 483646 304634
rect 483882 304398 483914 304634
rect 483294 268954 483914 304398
rect 483294 268718 483326 268954
rect 483562 268718 483646 268954
rect 483882 268718 483914 268954
rect 483294 268634 483914 268718
rect 483294 268398 483326 268634
rect 483562 268398 483646 268634
rect 483882 268398 483914 268634
rect 483294 232954 483914 268398
rect 483294 232718 483326 232954
rect 483562 232718 483646 232954
rect 483882 232718 483914 232954
rect 483294 232634 483914 232718
rect 483294 232398 483326 232634
rect 483562 232398 483646 232634
rect 483882 232398 483914 232634
rect 483294 196954 483914 232398
rect 483294 196718 483326 196954
rect 483562 196718 483646 196954
rect 483882 196718 483914 196954
rect 483294 196634 483914 196718
rect 483294 196398 483326 196634
rect 483562 196398 483646 196634
rect 483882 196398 483914 196634
rect 483294 160954 483914 196398
rect 483294 160718 483326 160954
rect 483562 160718 483646 160954
rect 483882 160718 483914 160954
rect 483294 160634 483914 160718
rect 483294 160398 483326 160634
rect 483562 160398 483646 160634
rect 483882 160398 483914 160634
rect 483294 124954 483914 160398
rect 483294 124718 483326 124954
rect 483562 124718 483646 124954
rect 483882 124718 483914 124954
rect 483294 124634 483914 124718
rect 483294 124398 483326 124634
rect 483562 124398 483646 124634
rect 483882 124398 483914 124634
rect 483294 88954 483914 124398
rect 483294 88718 483326 88954
rect 483562 88718 483646 88954
rect 483882 88718 483914 88954
rect 483294 88634 483914 88718
rect 483294 88398 483326 88634
rect 483562 88398 483646 88634
rect 483882 88398 483914 88634
rect 483294 52954 483914 88398
rect 483294 52718 483326 52954
rect 483562 52718 483646 52954
rect 483882 52718 483914 52954
rect 483294 52634 483914 52718
rect 483294 52398 483326 52634
rect 483562 52398 483646 52634
rect 483882 52398 483914 52634
rect 483294 16954 483914 52398
rect 483294 16718 483326 16954
rect 483562 16718 483646 16954
rect 483882 16718 483914 16954
rect 483294 16634 483914 16718
rect 483294 16398 483326 16634
rect 483562 16398 483646 16634
rect 483882 16398 483914 16634
rect 483294 -3226 483914 16398
rect 483294 -3462 483326 -3226
rect 483562 -3462 483646 -3226
rect 483882 -3462 483914 -3226
rect 483294 -3546 483914 -3462
rect 483294 -3782 483326 -3546
rect 483562 -3782 483646 -3546
rect 483882 -3782 483914 -3546
rect 483294 -7654 483914 -3782
rect 487794 708678 488414 711590
rect 487794 708442 487826 708678
rect 488062 708442 488146 708678
rect 488382 708442 488414 708678
rect 487794 708358 488414 708442
rect 487794 708122 487826 708358
rect 488062 708122 488146 708358
rect 488382 708122 488414 708358
rect 487794 669454 488414 708122
rect 487794 669218 487826 669454
rect 488062 669218 488146 669454
rect 488382 669218 488414 669454
rect 487794 669134 488414 669218
rect 487794 668898 487826 669134
rect 488062 668898 488146 669134
rect 488382 668898 488414 669134
rect 487794 633454 488414 668898
rect 487794 633218 487826 633454
rect 488062 633218 488146 633454
rect 488382 633218 488414 633454
rect 487794 633134 488414 633218
rect 487794 632898 487826 633134
rect 488062 632898 488146 633134
rect 488382 632898 488414 633134
rect 487794 597454 488414 632898
rect 487794 597218 487826 597454
rect 488062 597218 488146 597454
rect 488382 597218 488414 597454
rect 487794 597134 488414 597218
rect 487794 596898 487826 597134
rect 488062 596898 488146 597134
rect 488382 596898 488414 597134
rect 487794 561454 488414 596898
rect 487794 561218 487826 561454
rect 488062 561218 488146 561454
rect 488382 561218 488414 561454
rect 487794 561134 488414 561218
rect 487794 560898 487826 561134
rect 488062 560898 488146 561134
rect 488382 560898 488414 561134
rect 487794 525454 488414 560898
rect 487794 525218 487826 525454
rect 488062 525218 488146 525454
rect 488382 525218 488414 525454
rect 487794 525134 488414 525218
rect 487794 524898 487826 525134
rect 488062 524898 488146 525134
rect 488382 524898 488414 525134
rect 487794 489454 488414 524898
rect 487794 489218 487826 489454
rect 488062 489218 488146 489454
rect 488382 489218 488414 489454
rect 487794 489134 488414 489218
rect 487794 488898 487826 489134
rect 488062 488898 488146 489134
rect 488382 488898 488414 489134
rect 487794 453454 488414 488898
rect 487794 453218 487826 453454
rect 488062 453218 488146 453454
rect 488382 453218 488414 453454
rect 487794 453134 488414 453218
rect 487794 452898 487826 453134
rect 488062 452898 488146 453134
rect 488382 452898 488414 453134
rect 487794 417454 488414 452898
rect 487794 417218 487826 417454
rect 488062 417218 488146 417454
rect 488382 417218 488414 417454
rect 487794 417134 488414 417218
rect 487794 416898 487826 417134
rect 488062 416898 488146 417134
rect 488382 416898 488414 417134
rect 487794 381454 488414 416898
rect 487794 381218 487826 381454
rect 488062 381218 488146 381454
rect 488382 381218 488414 381454
rect 487794 381134 488414 381218
rect 487794 380898 487826 381134
rect 488062 380898 488146 381134
rect 488382 380898 488414 381134
rect 487794 345454 488414 380898
rect 487794 345218 487826 345454
rect 488062 345218 488146 345454
rect 488382 345218 488414 345454
rect 487794 345134 488414 345218
rect 487794 344898 487826 345134
rect 488062 344898 488146 345134
rect 488382 344898 488414 345134
rect 487794 309454 488414 344898
rect 487794 309218 487826 309454
rect 488062 309218 488146 309454
rect 488382 309218 488414 309454
rect 487794 309134 488414 309218
rect 487794 308898 487826 309134
rect 488062 308898 488146 309134
rect 488382 308898 488414 309134
rect 487794 273454 488414 308898
rect 487794 273218 487826 273454
rect 488062 273218 488146 273454
rect 488382 273218 488414 273454
rect 487794 273134 488414 273218
rect 487794 272898 487826 273134
rect 488062 272898 488146 273134
rect 488382 272898 488414 273134
rect 487794 237454 488414 272898
rect 487794 237218 487826 237454
rect 488062 237218 488146 237454
rect 488382 237218 488414 237454
rect 487794 237134 488414 237218
rect 487794 236898 487826 237134
rect 488062 236898 488146 237134
rect 488382 236898 488414 237134
rect 487794 201454 488414 236898
rect 487794 201218 487826 201454
rect 488062 201218 488146 201454
rect 488382 201218 488414 201454
rect 487794 201134 488414 201218
rect 487794 200898 487826 201134
rect 488062 200898 488146 201134
rect 488382 200898 488414 201134
rect 487794 165454 488414 200898
rect 487794 165218 487826 165454
rect 488062 165218 488146 165454
rect 488382 165218 488414 165454
rect 487794 165134 488414 165218
rect 487794 164898 487826 165134
rect 488062 164898 488146 165134
rect 488382 164898 488414 165134
rect 487794 129454 488414 164898
rect 487794 129218 487826 129454
rect 488062 129218 488146 129454
rect 488382 129218 488414 129454
rect 487794 129134 488414 129218
rect 487794 128898 487826 129134
rect 488062 128898 488146 129134
rect 488382 128898 488414 129134
rect 487794 93454 488414 128898
rect 487794 93218 487826 93454
rect 488062 93218 488146 93454
rect 488382 93218 488414 93454
rect 487794 93134 488414 93218
rect 487794 92898 487826 93134
rect 488062 92898 488146 93134
rect 488382 92898 488414 93134
rect 487794 57454 488414 92898
rect 487794 57218 487826 57454
rect 488062 57218 488146 57454
rect 488382 57218 488414 57454
rect 487794 57134 488414 57218
rect 487794 56898 487826 57134
rect 488062 56898 488146 57134
rect 488382 56898 488414 57134
rect 487794 21454 488414 56898
rect 487794 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 488414 21454
rect 487794 21134 488414 21218
rect 487794 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 488414 21134
rect 487794 -4186 488414 20898
rect 487794 -4422 487826 -4186
rect 488062 -4422 488146 -4186
rect 488382 -4422 488414 -4186
rect 487794 -4506 488414 -4422
rect 487794 -4742 487826 -4506
rect 488062 -4742 488146 -4506
rect 488382 -4742 488414 -4506
rect 487794 -7654 488414 -4742
rect 492294 709638 492914 711590
rect 492294 709402 492326 709638
rect 492562 709402 492646 709638
rect 492882 709402 492914 709638
rect 492294 709318 492914 709402
rect 492294 709082 492326 709318
rect 492562 709082 492646 709318
rect 492882 709082 492914 709318
rect 492294 673954 492914 709082
rect 492294 673718 492326 673954
rect 492562 673718 492646 673954
rect 492882 673718 492914 673954
rect 492294 673634 492914 673718
rect 492294 673398 492326 673634
rect 492562 673398 492646 673634
rect 492882 673398 492914 673634
rect 492294 637954 492914 673398
rect 492294 637718 492326 637954
rect 492562 637718 492646 637954
rect 492882 637718 492914 637954
rect 492294 637634 492914 637718
rect 492294 637398 492326 637634
rect 492562 637398 492646 637634
rect 492882 637398 492914 637634
rect 492294 601954 492914 637398
rect 492294 601718 492326 601954
rect 492562 601718 492646 601954
rect 492882 601718 492914 601954
rect 492294 601634 492914 601718
rect 492294 601398 492326 601634
rect 492562 601398 492646 601634
rect 492882 601398 492914 601634
rect 492294 565954 492914 601398
rect 492294 565718 492326 565954
rect 492562 565718 492646 565954
rect 492882 565718 492914 565954
rect 492294 565634 492914 565718
rect 492294 565398 492326 565634
rect 492562 565398 492646 565634
rect 492882 565398 492914 565634
rect 492294 529954 492914 565398
rect 492294 529718 492326 529954
rect 492562 529718 492646 529954
rect 492882 529718 492914 529954
rect 492294 529634 492914 529718
rect 492294 529398 492326 529634
rect 492562 529398 492646 529634
rect 492882 529398 492914 529634
rect 492294 493954 492914 529398
rect 492294 493718 492326 493954
rect 492562 493718 492646 493954
rect 492882 493718 492914 493954
rect 492294 493634 492914 493718
rect 492294 493398 492326 493634
rect 492562 493398 492646 493634
rect 492882 493398 492914 493634
rect 492294 457954 492914 493398
rect 492294 457718 492326 457954
rect 492562 457718 492646 457954
rect 492882 457718 492914 457954
rect 492294 457634 492914 457718
rect 492294 457398 492326 457634
rect 492562 457398 492646 457634
rect 492882 457398 492914 457634
rect 492294 421954 492914 457398
rect 492294 421718 492326 421954
rect 492562 421718 492646 421954
rect 492882 421718 492914 421954
rect 492294 421634 492914 421718
rect 492294 421398 492326 421634
rect 492562 421398 492646 421634
rect 492882 421398 492914 421634
rect 492294 385954 492914 421398
rect 492294 385718 492326 385954
rect 492562 385718 492646 385954
rect 492882 385718 492914 385954
rect 492294 385634 492914 385718
rect 492294 385398 492326 385634
rect 492562 385398 492646 385634
rect 492882 385398 492914 385634
rect 492294 349954 492914 385398
rect 492294 349718 492326 349954
rect 492562 349718 492646 349954
rect 492882 349718 492914 349954
rect 492294 349634 492914 349718
rect 492294 349398 492326 349634
rect 492562 349398 492646 349634
rect 492882 349398 492914 349634
rect 492294 313954 492914 349398
rect 492294 313718 492326 313954
rect 492562 313718 492646 313954
rect 492882 313718 492914 313954
rect 492294 313634 492914 313718
rect 492294 313398 492326 313634
rect 492562 313398 492646 313634
rect 492882 313398 492914 313634
rect 492294 277954 492914 313398
rect 492294 277718 492326 277954
rect 492562 277718 492646 277954
rect 492882 277718 492914 277954
rect 492294 277634 492914 277718
rect 492294 277398 492326 277634
rect 492562 277398 492646 277634
rect 492882 277398 492914 277634
rect 492294 241954 492914 277398
rect 492294 241718 492326 241954
rect 492562 241718 492646 241954
rect 492882 241718 492914 241954
rect 492294 241634 492914 241718
rect 492294 241398 492326 241634
rect 492562 241398 492646 241634
rect 492882 241398 492914 241634
rect 492294 205954 492914 241398
rect 492294 205718 492326 205954
rect 492562 205718 492646 205954
rect 492882 205718 492914 205954
rect 492294 205634 492914 205718
rect 492294 205398 492326 205634
rect 492562 205398 492646 205634
rect 492882 205398 492914 205634
rect 492294 169954 492914 205398
rect 492294 169718 492326 169954
rect 492562 169718 492646 169954
rect 492882 169718 492914 169954
rect 492294 169634 492914 169718
rect 492294 169398 492326 169634
rect 492562 169398 492646 169634
rect 492882 169398 492914 169634
rect 492294 133954 492914 169398
rect 492294 133718 492326 133954
rect 492562 133718 492646 133954
rect 492882 133718 492914 133954
rect 492294 133634 492914 133718
rect 492294 133398 492326 133634
rect 492562 133398 492646 133634
rect 492882 133398 492914 133634
rect 492294 97954 492914 133398
rect 492294 97718 492326 97954
rect 492562 97718 492646 97954
rect 492882 97718 492914 97954
rect 492294 97634 492914 97718
rect 492294 97398 492326 97634
rect 492562 97398 492646 97634
rect 492882 97398 492914 97634
rect 492294 61954 492914 97398
rect 492294 61718 492326 61954
rect 492562 61718 492646 61954
rect 492882 61718 492914 61954
rect 492294 61634 492914 61718
rect 492294 61398 492326 61634
rect 492562 61398 492646 61634
rect 492882 61398 492914 61634
rect 492294 25954 492914 61398
rect 492294 25718 492326 25954
rect 492562 25718 492646 25954
rect 492882 25718 492914 25954
rect 492294 25634 492914 25718
rect 492294 25398 492326 25634
rect 492562 25398 492646 25634
rect 492882 25398 492914 25634
rect 492294 -5146 492914 25398
rect 492294 -5382 492326 -5146
rect 492562 -5382 492646 -5146
rect 492882 -5382 492914 -5146
rect 492294 -5466 492914 -5382
rect 492294 -5702 492326 -5466
rect 492562 -5702 492646 -5466
rect 492882 -5702 492914 -5466
rect 492294 -7654 492914 -5702
rect 496794 710598 497414 711590
rect 496794 710362 496826 710598
rect 497062 710362 497146 710598
rect 497382 710362 497414 710598
rect 496794 710278 497414 710362
rect 496794 710042 496826 710278
rect 497062 710042 497146 710278
rect 497382 710042 497414 710278
rect 496794 678454 497414 710042
rect 496794 678218 496826 678454
rect 497062 678218 497146 678454
rect 497382 678218 497414 678454
rect 496794 678134 497414 678218
rect 496794 677898 496826 678134
rect 497062 677898 497146 678134
rect 497382 677898 497414 678134
rect 496794 642454 497414 677898
rect 496794 642218 496826 642454
rect 497062 642218 497146 642454
rect 497382 642218 497414 642454
rect 496794 642134 497414 642218
rect 496794 641898 496826 642134
rect 497062 641898 497146 642134
rect 497382 641898 497414 642134
rect 496794 606454 497414 641898
rect 496794 606218 496826 606454
rect 497062 606218 497146 606454
rect 497382 606218 497414 606454
rect 496794 606134 497414 606218
rect 496794 605898 496826 606134
rect 497062 605898 497146 606134
rect 497382 605898 497414 606134
rect 496794 570454 497414 605898
rect 496794 570218 496826 570454
rect 497062 570218 497146 570454
rect 497382 570218 497414 570454
rect 496794 570134 497414 570218
rect 496794 569898 496826 570134
rect 497062 569898 497146 570134
rect 497382 569898 497414 570134
rect 496794 534454 497414 569898
rect 496794 534218 496826 534454
rect 497062 534218 497146 534454
rect 497382 534218 497414 534454
rect 496794 534134 497414 534218
rect 496794 533898 496826 534134
rect 497062 533898 497146 534134
rect 497382 533898 497414 534134
rect 496794 498454 497414 533898
rect 496794 498218 496826 498454
rect 497062 498218 497146 498454
rect 497382 498218 497414 498454
rect 496794 498134 497414 498218
rect 496794 497898 496826 498134
rect 497062 497898 497146 498134
rect 497382 497898 497414 498134
rect 496794 462454 497414 497898
rect 496794 462218 496826 462454
rect 497062 462218 497146 462454
rect 497382 462218 497414 462454
rect 496794 462134 497414 462218
rect 496794 461898 496826 462134
rect 497062 461898 497146 462134
rect 497382 461898 497414 462134
rect 496794 426454 497414 461898
rect 496794 426218 496826 426454
rect 497062 426218 497146 426454
rect 497382 426218 497414 426454
rect 496794 426134 497414 426218
rect 496794 425898 496826 426134
rect 497062 425898 497146 426134
rect 497382 425898 497414 426134
rect 496794 390454 497414 425898
rect 496794 390218 496826 390454
rect 497062 390218 497146 390454
rect 497382 390218 497414 390454
rect 496794 390134 497414 390218
rect 496794 389898 496826 390134
rect 497062 389898 497146 390134
rect 497382 389898 497414 390134
rect 496794 354454 497414 389898
rect 496794 354218 496826 354454
rect 497062 354218 497146 354454
rect 497382 354218 497414 354454
rect 496794 354134 497414 354218
rect 496794 353898 496826 354134
rect 497062 353898 497146 354134
rect 497382 353898 497414 354134
rect 496794 318454 497414 353898
rect 496794 318218 496826 318454
rect 497062 318218 497146 318454
rect 497382 318218 497414 318454
rect 496794 318134 497414 318218
rect 496794 317898 496826 318134
rect 497062 317898 497146 318134
rect 497382 317898 497414 318134
rect 496794 282454 497414 317898
rect 496794 282218 496826 282454
rect 497062 282218 497146 282454
rect 497382 282218 497414 282454
rect 496794 282134 497414 282218
rect 496794 281898 496826 282134
rect 497062 281898 497146 282134
rect 497382 281898 497414 282134
rect 496794 246454 497414 281898
rect 496794 246218 496826 246454
rect 497062 246218 497146 246454
rect 497382 246218 497414 246454
rect 496794 246134 497414 246218
rect 496794 245898 496826 246134
rect 497062 245898 497146 246134
rect 497382 245898 497414 246134
rect 496794 210454 497414 245898
rect 496794 210218 496826 210454
rect 497062 210218 497146 210454
rect 497382 210218 497414 210454
rect 496794 210134 497414 210218
rect 496794 209898 496826 210134
rect 497062 209898 497146 210134
rect 497382 209898 497414 210134
rect 496794 174454 497414 209898
rect 496794 174218 496826 174454
rect 497062 174218 497146 174454
rect 497382 174218 497414 174454
rect 496794 174134 497414 174218
rect 496794 173898 496826 174134
rect 497062 173898 497146 174134
rect 497382 173898 497414 174134
rect 496794 138454 497414 173898
rect 496794 138218 496826 138454
rect 497062 138218 497146 138454
rect 497382 138218 497414 138454
rect 496794 138134 497414 138218
rect 496794 137898 496826 138134
rect 497062 137898 497146 138134
rect 497382 137898 497414 138134
rect 496794 102454 497414 137898
rect 496794 102218 496826 102454
rect 497062 102218 497146 102454
rect 497382 102218 497414 102454
rect 496794 102134 497414 102218
rect 496794 101898 496826 102134
rect 497062 101898 497146 102134
rect 497382 101898 497414 102134
rect 496794 66454 497414 101898
rect 496794 66218 496826 66454
rect 497062 66218 497146 66454
rect 497382 66218 497414 66454
rect 496794 66134 497414 66218
rect 496794 65898 496826 66134
rect 497062 65898 497146 66134
rect 497382 65898 497414 66134
rect 496794 30454 497414 65898
rect 496794 30218 496826 30454
rect 497062 30218 497146 30454
rect 497382 30218 497414 30454
rect 496794 30134 497414 30218
rect 496794 29898 496826 30134
rect 497062 29898 497146 30134
rect 497382 29898 497414 30134
rect 496794 -6106 497414 29898
rect 496794 -6342 496826 -6106
rect 497062 -6342 497146 -6106
rect 497382 -6342 497414 -6106
rect 496794 -6426 497414 -6342
rect 496794 -6662 496826 -6426
rect 497062 -6662 497146 -6426
rect 497382 -6662 497414 -6426
rect 496794 -7654 497414 -6662
rect 501294 711558 501914 711590
rect 501294 711322 501326 711558
rect 501562 711322 501646 711558
rect 501882 711322 501914 711558
rect 501294 711238 501914 711322
rect 501294 711002 501326 711238
rect 501562 711002 501646 711238
rect 501882 711002 501914 711238
rect 501294 682954 501914 711002
rect 501294 682718 501326 682954
rect 501562 682718 501646 682954
rect 501882 682718 501914 682954
rect 501294 682634 501914 682718
rect 501294 682398 501326 682634
rect 501562 682398 501646 682634
rect 501882 682398 501914 682634
rect 501294 646954 501914 682398
rect 501294 646718 501326 646954
rect 501562 646718 501646 646954
rect 501882 646718 501914 646954
rect 501294 646634 501914 646718
rect 501294 646398 501326 646634
rect 501562 646398 501646 646634
rect 501882 646398 501914 646634
rect 501294 610954 501914 646398
rect 501294 610718 501326 610954
rect 501562 610718 501646 610954
rect 501882 610718 501914 610954
rect 501294 610634 501914 610718
rect 501294 610398 501326 610634
rect 501562 610398 501646 610634
rect 501882 610398 501914 610634
rect 501294 574954 501914 610398
rect 501294 574718 501326 574954
rect 501562 574718 501646 574954
rect 501882 574718 501914 574954
rect 501294 574634 501914 574718
rect 501294 574398 501326 574634
rect 501562 574398 501646 574634
rect 501882 574398 501914 574634
rect 501294 538954 501914 574398
rect 501294 538718 501326 538954
rect 501562 538718 501646 538954
rect 501882 538718 501914 538954
rect 501294 538634 501914 538718
rect 501294 538398 501326 538634
rect 501562 538398 501646 538634
rect 501882 538398 501914 538634
rect 501294 502954 501914 538398
rect 501294 502718 501326 502954
rect 501562 502718 501646 502954
rect 501882 502718 501914 502954
rect 501294 502634 501914 502718
rect 501294 502398 501326 502634
rect 501562 502398 501646 502634
rect 501882 502398 501914 502634
rect 501294 466954 501914 502398
rect 501294 466718 501326 466954
rect 501562 466718 501646 466954
rect 501882 466718 501914 466954
rect 501294 466634 501914 466718
rect 501294 466398 501326 466634
rect 501562 466398 501646 466634
rect 501882 466398 501914 466634
rect 501294 430954 501914 466398
rect 501294 430718 501326 430954
rect 501562 430718 501646 430954
rect 501882 430718 501914 430954
rect 501294 430634 501914 430718
rect 501294 430398 501326 430634
rect 501562 430398 501646 430634
rect 501882 430398 501914 430634
rect 501294 394954 501914 430398
rect 501294 394718 501326 394954
rect 501562 394718 501646 394954
rect 501882 394718 501914 394954
rect 501294 394634 501914 394718
rect 501294 394398 501326 394634
rect 501562 394398 501646 394634
rect 501882 394398 501914 394634
rect 501294 358954 501914 394398
rect 501294 358718 501326 358954
rect 501562 358718 501646 358954
rect 501882 358718 501914 358954
rect 501294 358634 501914 358718
rect 501294 358398 501326 358634
rect 501562 358398 501646 358634
rect 501882 358398 501914 358634
rect 501294 322954 501914 358398
rect 501294 322718 501326 322954
rect 501562 322718 501646 322954
rect 501882 322718 501914 322954
rect 501294 322634 501914 322718
rect 501294 322398 501326 322634
rect 501562 322398 501646 322634
rect 501882 322398 501914 322634
rect 501294 286954 501914 322398
rect 501294 286718 501326 286954
rect 501562 286718 501646 286954
rect 501882 286718 501914 286954
rect 501294 286634 501914 286718
rect 501294 286398 501326 286634
rect 501562 286398 501646 286634
rect 501882 286398 501914 286634
rect 501294 250954 501914 286398
rect 501294 250718 501326 250954
rect 501562 250718 501646 250954
rect 501882 250718 501914 250954
rect 501294 250634 501914 250718
rect 501294 250398 501326 250634
rect 501562 250398 501646 250634
rect 501882 250398 501914 250634
rect 501294 214954 501914 250398
rect 501294 214718 501326 214954
rect 501562 214718 501646 214954
rect 501882 214718 501914 214954
rect 501294 214634 501914 214718
rect 501294 214398 501326 214634
rect 501562 214398 501646 214634
rect 501882 214398 501914 214634
rect 501294 178954 501914 214398
rect 501294 178718 501326 178954
rect 501562 178718 501646 178954
rect 501882 178718 501914 178954
rect 501294 178634 501914 178718
rect 501294 178398 501326 178634
rect 501562 178398 501646 178634
rect 501882 178398 501914 178634
rect 501294 142954 501914 178398
rect 501294 142718 501326 142954
rect 501562 142718 501646 142954
rect 501882 142718 501914 142954
rect 501294 142634 501914 142718
rect 501294 142398 501326 142634
rect 501562 142398 501646 142634
rect 501882 142398 501914 142634
rect 501294 106954 501914 142398
rect 501294 106718 501326 106954
rect 501562 106718 501646 106954
rect 501882 106718 501914 106954
rect 501294 106634 501914 106718
rect 501294 106398 501326 106634
rect 501562 106398 501646 106634
rect 501882 106398 501914 106634
rect 501294 70954 501914 106398
rect 501294 70718 501326 70954
rect 501562 70718 501646 70954
rect 501882 70718 501914 70954
rect 501294 70634 501914 70718
rect 501294 70398 501326 70634
rect 501562 70398 501646 70634
rect 501882 70398 501914 70634
rect 501294 34954 501914 70398
rect 501294 34718 501326 34954
rect 501562 34718 501646 34954
rect 501882 34718 501914 34954
rect 501294 34634 501914 34718
rect 501294 34398 501326 34634
rect 501562 34398 501646 34634
rect 501882 34398 501914 34634
rect 501294 -7066 501914 34398
rect 501294 -7302 501326 -7066
rect 501562 -7302 501646 -7066
rect 501882 -7302 501914 -7066
rect 501294 -7386 501914 -7302
rect 501294 -7622 501326 -7386
rect 501562 -7622 501646 -7386
rect 501882 -7622 501914 -7386
rect 501294 -7654 501914 -7622
rect 505794 704838 506414 711590
rect 505794 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 506414 704838
rect 505794 704518 506414 704602
rect 505794 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 506414 704518
rect 505794 687454 506414 704282
rect 505794 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 506414 687454
rect 505794 687134 506414 687218
rect 505794 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 506414 687134
rect 505794 651454 506414 686898
rect 505794 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 506414 651454
rect 505794 651134 506414 651218
rect 505794 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 506414 651134
rect 505794 615454 506414 650898
rect 505794 615218 505826 615454
rect 506062 615218 506146 615454
rect 506382 615218 506414 615454
rect 505794 615134 506414 615218
rect 505794 614898 505826 615134
rect 506062 614898 506146 615134
rect 506382 614898 506414 615134
rect 505794 579454 506414 614898
rect 505794 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 506414 579454
rect 505794 579134 506414 579218
rect 505794 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 506414 579134
rect 505794 543454 506414 578898
rect 505794 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 506414 543454
rect 505794 543134 506414 543218
rect 505794 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 506414 543134
rect 505794 507454 506414 542898
rect 505794 507218 505826 507454
rect 506062 507218 506146 507454
rect 506382 507218 506414 507454
rect 505794 507134 506414 507218
rect 505794 506898 505826 507134
rect 506062 506898 506146 507134
rect 506382 506898 506414 507134
rect 505794 471454 506414 506898
rect 505794 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 506414 471454
rect 505794 471134 506414 471218
rect 505794 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 506414 471134
rect 505794 435454 506414 470898
rect 505794 435218 505826 435454
rect 506062 435218 506146 435454
rect 506382 435218 506414 435454
rect 505794 435134 506414 435218
rect 505794 434898 505826 435134
rect 506062 434898 506146 435134
rect 506382 434898 506414 435134
rect 505794 399454 506414 434898
rect 505794 399218 505826 399454
rect 506062 399218 506146 399454
rect 506382 399218 506414 399454
rect 505794 399134 506414 399218
rect 505794 398898 505826 399134
rect 506062 398898 506146 399134
rect 506382 398898 506414 399134
rect 505794 363454 506414 398898
rect 505794 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 506414 363454
rect 505794 363134 506414 363218
rect 505794 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 506414 363134
rect 505794 327454 506414 362898
rect 505794 327218 505826 327454
rect 506062 327218 506146 327454
rect 506382 327218 506414 327454
rect 505794 327134 506414 327218
rect 505794 326898 505826 327134
rect 506062 326898 506146 327134
rect 506382 326898 506414 327134
rect 505794 291454 506414 326898
rect 505794 291218 505826 291454
rect 506062 291218 506146 291454
rect 506382 291218 506414 291454
rect 505794 291134 506414 291218
rect 505794 290898 505826 291134
rect 506062 290898 506146 291134
rect 506382 290898 506414 291134
rect 505794 255454 506414 290898
rect 505794 255218 505826 255454
rect 506062 255218 506146 255454
rect 506382 255218 506414 255454
rect 505794 255134 506414 255218
rect 505794 254898 505826 255134
rect 506062 254898 506146 255134
rect 506382 254898 506414 255134
rect 505794 219454 506414 254898
rect 505794 219218 505826 219454
rect 506062 219218 506146 219454
rect 506382 219218 506414 219454
rect 505794 219134 506414 219218
rect 505794 218898 505826 219134
rect 506062 218898 506146 219134
rect 506382 218898 506414 219134
rect 505794 183454 506414 218898
rect 505794 183218 505826 183454
rect 506062 183218 506146 183454
rect 506382 183218 506414 183454
rect 505794 183134 506414 183218
rect 505794 182898 505826 183134
rect 506062 182898 506146 183134
rect 506382 182898 506414 183134
rect 505794 147454 506414 182898
rect 505794 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 506414 147454
rect 505794 147134 506414 147218
rect 505794 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 506414 147134
rect 505794 111454 506414 146898
rect 505794 111218 505826 111454
rect 506062 111218 506146 111454
rect 506382 111218 506414 111454
rect 505794 111134 506414 111218
rect 505794 110898 505826 111134
rect 506062 110898 506146 111134
rect 506382 110898 506414 111134
rect 505794 75454 506414 110898
rect 505794 75218 505826 75454
rect 506062 75218 506146 75454
rect 506382 75218 506414 75454
rect 505794 75134 506414 75218
rect 505794 74898 505826 75134
rect 506062 74898 506146 75134
rect 506382 74898 506414 75134
rect 505794 39454 506414 74898
rect 505794 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 506414 39454
rect 505794 39134 506414 39218
rect 505794 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 506414 39134
rect 505794 3454 506414 38898
rect 505794 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 506414 3454
rect 505794 3134 506414 3218
rect 505794 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 506414 3134
rect 505794 -346 506414 2898
rect 505794 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 506414 -346
rect 505794 -666 506414 -582
rect 505794 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 506414 -666
rect 505794 -7654 506414 -902
rect 510294 705798 510914 711590
rect 510294 705562 510326 705798
rect 510562 705562 510646 705798
rect 510882 705562 510914 705798
rect 510294 705478 510914 705562
rect 510294 705242 510326 705478
rect 510562 705242 510646 705478
rect 510882 705242 510914 705478
rect 510294 691954 510914 705242
rect 510294 691718 510326 691954
rect 510562 691718 510646 691954
rect 510882 691718 510914 691954
rect 510294 691634 510914 691718
rect 510294 691398 510326 691634
rect 510562 691398 510646 691634
rect 510882 691398 510914 691634
rect 510294 655954 510914 691398
rect 510294 655718 510326 655954
rect 510562 655718 510646 655954
rect 510882 655718 510914 655954
rect 510294 655634 510914 655718
rect 510294 655398 510326 655634
rect 510562 655398 510646 655634
rect 510882 655398 510914 655634
rect 510294 619954 510914 655398
rect 510294 619718 510326 619954
rect 510562 619718 510646 619954
rect 510882 619718 510914 619954
rect 510294 619634 510914 619718
rect 510294 619398 510326 619634
rect 510562 619398 510646 619634
rect 510882 619398 510914 619634
rect 510294 583954 510914 619398
rect 510294 583718 510326 583954
rect 510562 583718 510646 583954
rect 510882 583718 510914 583954
rect 510294 583634 510914 583718
rect 510294 583398 510326 583634
rect 510562 583398 510646 583634
rect 510882 583398 510914 583634
rect 510294 547954 510914 583398
rect 510294 547718 510326 547954
rect 510562 547718 510646 547954
rect 510882 547718 510914 547954
rect 510294 547634 510914 547718
rect 510294 547398 510326 547634
rect 510562 547398 510646 547634
rect 510882 547398 510914 547634
rect 510294 511954 510914 547398
rect 510294 511718 510326 511954
rect 510562 511718 510646 511954
rect 510882 511718 510914 511954
rect 510294 511634 510914 511718
rect 510294 511398 510326 511634
rect 510562 511398 510646 511634
rect 510882 511398 510914 511634
rect 510294 475954 510914 511398
rect 510294 475718 510326 475954
rect 510562 475718 510646 475954
rect 510882 475718 510914 475954
rect 510294 475634 510914 475718
rect 510294 475398 510326 475634
rect 510562 475398 510646 475634
rect 510882 475398 510914 475634
rect 510294 439954 510914 475398
rect 510294 439718 510326 439954
rect 510562 439718 510646 439954
rect 510882 439718 510914 439954
rect 510294 439634 510914 439718
rect 510294 439398 510326 439634
rect 510562 439398 510646 439634
rect 510882 439398 510914 439634
rect 510294 403954 510914 439398
rect 510294 403718 510326 403954
rect 510562 403718 510646 403954
rect 510882 403718 510914 403954
rect 510294 403634 510914 403718
rect 510294 403398 510326 403634
rect 510562 403398 510646 403634
rect 510882 403398 510914 403634
rect 510294 367954 510914 403398
rect 510294 367718 510326 367954
rect 510562 367718 510646 367954
rect 510882 367718 510914 367954
rect 510294 367634 510914 367718
rect 510294 367398 510326 367634
rect 510562 367398 510646 367634
rect 510882 367398 510914 367634
rect 510294 331954 510914 367398
rect 510294 331718 510326 331954
rect 510562 331718 510646 331954
rect 510882 331718 510914 331954
rect 510294 331634 510914 331718
rect 510294 331398 510326 331634
rect 510562 331398 510646 331634
rect 510882 331398 510914 331634
rect 510294 295954 510914 331398
rect 510294 295718 510326 295954
rect 510562 295718 510646 295954
rect 510882 295718 510914 295954
rect 510294 295634 510914 295718
rect 510294 295398 510326 295634
rect 510562 295398 510646 295634
rect 510882 295398 510914 295634
rect 510294 259954 510914 295398
rect 510294 259718 510326 259954
rect 510562 259718 510646 259954
rect 510882 259718 510914 259954
rect 510294 259634 510914 259718
rect 510294 259398 510326 259634
rect 510562 259398 510646 259634
rect 510882 259398 510914 259634
rect 510294 223954 510914 259398
rect 510294 223718 510326 223954
rect 510562 223718 510646 223954
rect 510882 223718 510914 223954
rect 510294 223634 510914 223718
rect 510294 223398 510326 223634
rect 510562 223398 510646 223634
rect 510882 223398 510914 223634
rect 510294 187954 510914 223398
rect 510294 187718 510326 187954
rect 510562 187718 510646 187954
rect 510882 187718 510914 187954
rect 510294 187634 510914 187718
rect 510294 187398 510326 187634
rect 510562 187398 510646 187634
rect 510882 187398 510914 187634
rect 510294 151954 510914 187398
rect 510294 151718 510326 151954
rect 510562 151718 510646 151954
rect 510882 151718 510914 151954
rect 510294 151634 510914 151718
rect 510294 151398 510326 151634
rect 510562 151398 510646 151634
rect 510882 151398 510914 151634
rect 510294 115954 510914 151398
rect 510294 115718 510326 115954
rect 510562 115718 510646 115954
rect 510882 115718 510914 115954
rect 510294 115634 510914 115718
rect 510294 115398 510326 115634
rect 510562 115398 510646 115634
rect 510882 115398 510914 115634
rect 510294 79954 510914 115398
rect 510294 79718 510326 79954
rect 510562 79718 510646 79954
rect 510882 79718 510914 79954
rect 510294 79634 510914 79718
rect 510294 79398 510326 79634
rect 510562 79398 510646 79634
rect 510882 79398 510914 79634
rect 510294 43954 510914 79398
rect 510294 43718 510326 43954
rect 510562 43718 510646 43954
rect 510882 43718 510914 43954
rect 510294 43634 510914 43718
rect 510294 43398 510326 43634
rect 510562 43398 510646 43634
rect 510882 43398 510914 43634
rect 510294 7954 510914 43398
rect 510294 7718 510326 7954
rect 510562 7718 510646 7954
rect 510882 7718 510914 7954
rect 510294 7634 510914 7718
rect 510294 7398 510326 7634
rect 510562 7398 510646 7634
rect 510882 7398 510914 7634
rect 510294 -1306 510914 7398
rect 510294 -1542 510326 -1306
rect 510562 -1542 510646 -1306
rect 510882 -1542 510914 -1306
rect 510294 -1626 510914 -1542
rect 510294 -1862 510326 -1626
rect 510562 -1862 510646 -1626
rect 510882 -1862 510914 -1626
rect 510294 -7654 510914 -1862
rect 514794 706758 515414 711590
rect 514794 706522 514826 706758
rect 515062 706522 515146 706758
rect 515382 706522 515414 706758
rect 514794 706438 515414 706522
rect 514794 706202 514826 706438
rect 515062 706202 515146 706438
rect 515382 706202 515414 706438
rect 514794 696454 515414 706202
rect 514794 696218 514826 696454
rect 515062 696218 515146 696454
rect 515382 696218 515414 696454
rect 514794 696134 515414 696218
rect 514794 695898 514826 696134
rect 515062 695898 515146 696134
rect 515382 695898 515414 696134
rect 514794 660454 515414 695898
rect 514794 660218 514826 660454
rect 515062 660218 515146 660454
rect 515382 660218 515414 660454
rect 514794 660134 515414 660218
rect 514794 659898 514826 660134
rect 515062 659898 515146 660134
rect 515382 659898 515414 660134
rect 514794 624454 515414 659898
rect 514794 624218 514826 624454
rect 515062 624218 515146 624454
rect 515382 624218 515414 624454
rect 514794 624134 515414 624218
rect 514794 623898 514826 624134
rect 515062 623898 515146 624134
rect 515382 623898 515414 624134
rect 514794 588454 515414 623898
rect 514794 588218 514826 588454
rect 515062 588218 515146 588454
rect 515382 588218 515414 588454
rect 514794 588134 515414 588218
rect 514794 587898 514826 588134
rect 515062 587898 515146 588134
rect 515382 587898 515414 588134
rect 514794 552454 515414 587898
rect 514794 552218 514826 552454
rect 515062 552218 515146 552454
rect 515382 552218 515414 552454
rect 514794 552134 515414 552218
rect 514794 551898 514826 552134
rect 515062 551898 515146 552134
rect 515382 551898 515414 552134
rect 514794 516454 515414 551898
rect 514794 516218 514826 516454
rect 515062 516218 515146 516454
rect 515382 516218 515414 516454
rect 514794 516134 515414 516218
rect 514794 515898 514826 516134
rect 515062 515898 515146 516134
rect 515382 515898 515414 516134
rect 514794 480454 515414 515898
rect 514794 480218 514826 480454
rect 515062 480218 515146 480454
rect 515382 480218 515414 480454
rect 514794 480134 515414 480218
rect 514794 479898 514826 480134
rect 515062 479898 515146 480134
rect 515382 479898 515414 480134
rect 514794 444454 515414 479898
rect 514794 444218 514826 444454
rect 515062 444218 515146 444454
rect 515382 444218 515414 444454
rect 514794 444134 515414 444218
rect 514794 443898 514826 444134
rect 515062 443898 515146 444134
rect 515382 443898 515414 444134
rect 514794 408454 515414 443898
rect 514794 408218 514826 408454
rect 515062 408218 515146 408454
rect 515382 408218 515414 408454
rect 514794 408134 515414 408218
rect 514794 407898 514826 408134
rect 515062 407898 515146 408134
rect 515382 407898 515414 408134
rect 514794 372454 515414 407898
rect 514794 372218 514826 372454
rect 515062 372218 515146 372454
rect 515382 372218 515414 372454
rect 514794 372134 515414 372218
rect 514794 371898 514826 372134
rect 515062 371898 515146 372134
rect 515382 371898 515414 372134
rect 514794 336454 515414 371898
rect 514794 336218 514826 336454
rect 515062 336218 515146 336454
rect 515382 336218 515414 336454
rect 514794 336134 515414 336218
rect 514794 335898 514826 336134
rect 515062 335898 515146 336134
rect 515382 335898 515414 336134
rect 514794 300454 515414 335898
rect 514794 300218 514826 300454
rect 515062 300218 515146 300454
rect 515382 300218 515414 300454
rect 514794 300134 515414 300218
rect 514794 299898 514826 300134
rect 515062 299898 515146 300134
rect 515382 299898 515414 300134
rect 514794 264454 515414 299898
rect 514794 264218 514826 264454
rect 515062 264218 515146 264454
rect 515382 264218 515414 264454
rect 514794 264134 515414 264218
rect 514794 263898 514826 264134
rect 515062 263898 515146 264134
rect 515382 263898 515414 264134
rect 514794 228454 515414 263898
rect 514794 228218 514826 228454
rect 515062 228218 515146 228454
rect 515382 228218 515414 228454
rect 514794 228134 515414 228218
rect 514794 227898 514826 228134
rect 515062 227898 515146 228134
rect 515382 227898 515414 228134
rect 514794 192454 515414 227898
rect 514794 192218 514826 192454
rect 515062 192218 515146 192454
rect 515382 192218 515414 192454
rect 514794 192134 515414 192218
rect 514794 191898 514826 192134
rect 515062 191898 515146 192134
rect 515382 191898 515414 192134
rect 514794 156454 515414 191898
rect 514794 156218 514826 156454
rect 515062 156218 515146 156454
rect 515382 156218 515414 156454
rect 514794 156134 515414 156218
rect 514794 155898 514826 156134
rect 515062 155898 515146 156134
rect 515382 155898 515414 156134
rect 514794 120454 515414 155898
rect 514794 120218 514826 120454
rect 515062 120218 515146 120454
rect 515382 120218 515414 120454
rect 514794 120134 515414 120218
rect 514794 119898 514826 120134
rect 515062 119898 515146 120134
rect 515382 119898 515414 120134
rect 514794 84454 515414 119898
rect 514794 84218 514826 84454
rect 515062 84218 515146 84454
rect 515382 84218 515414 84454
rect 514794 84134 515414 84218
rect 514794 83898 514826 84134
rect 515062 83898 515146 84134
rect 515382 83898 515414 84134
rect 514794 48454 515414 83898
rect 514794 48218 514826 48454
rect 515062 48218 515146 48454
rect 515382 48218 515414 48454
rect 514794 48134 515414 48218
rect 514794 47898 514826 48134
rect 515062 47898 515146 48134
rect 515382 47898 515414 48134
rect 514794 12454 515414 47898
rect 514794 12218 514826 12454
rect 515062 12218 515146 12454
rect 515382 12218 515414 12454
rect 514794 12134 515414 12218
rect 514794 11898 514826 12134
rect 515062 11898 515146 12134
rect 515382 11898 515414 12134
rect 514794 -2266 515414 11898
rect 514794 -2502 514826 -2266
rect 515062 -2502 515146 -2266
rect 515382 -2502 515414 -2266
rect 514794 -2586 515414 -2502
rect 514794 -2822 514826 -2586
rect 515062 -2822 515146 -2586
rect 515382 -2822 515414 -2586
rect 514794 -7654 515414 -2822
rect 519294 707718 519914 711590
rect 519294 707482 519326 707718
rect 519562 707482 519646 707718
rect 519882 707482 519914 707718
rect 519294 707398 519914 707482
rect 519294 707162 519326 707398
rect 519562 707162 519646 707398
rect 519882 707162 519914 707398
rect 519294 700954 519914 707162
rect 519294 700718 519326 700954
rect 519562 700718 519646 700954
rect 519882 700718 519914 700954
rect 519294 700634 519914 700718
rect 519294 700398 519326 700634
rect 519562 700398 519646 700634
rect 519882 700398 519914 700634
rect 519294 664954 519914 700398
rect 519294 664718 519326 664954
rect 519562 664718 519646 664954
rect 519882 664718 519914 664954
rect 519294 664634 519914 664718
rect 519294 664398 519326 664634
rect 519562 664398 519646 664634
rect 519882 664398 519914 664634
rect 519294 628954 519914 664398
rect 519294 628718 519326 628954
rect 519562 628718 519646 628954
rect 519882 628718 519914 628954
rect 519294 628634 519914 628718
rect 519294 628398 519326 628634
rect 519562 628398 519646 628634
rect 519882 628398 519914 628634
rect 519294 592954 519914 628398
rect 519294 592718 519326 592954
rect 519562 592718 519646 592954
rect 519882 592718 519914 592954
rect 519294 592634 519914 592718
rect 519294 592398 519326 592634
rect 519562 592398 519646 592634
rect 519882 592398 519914 592634
rect 519294 556954 519914 592398
rect 519294 556718 519326 556954
rect 519562 556718 519646 556954
rect 519882 556718 519914 556954
rect 519294 556634 519914 556718
rect 519294 556398 519326 556634
rect 519562 556398 519646 556634
rect 519882 556398 519914 556634
rect 519294 520954 519914 556398
rect 519294 520718 519326 520954
rect 519562 520718 519646 520954
rect 519882 520718 519914 520954
rect 519294 520634 519914 520718
rect 519294 520398 519326 520634
rect 519562 520398 519646 520634
rect 519882 520398 519914 520634
rect 519294 484954 519914 520398
rect 519294 484718 519326 484954
rect 519562 484718 519646 484954
rect 519882 484718 519914 484954
rect 519294 484634 519914 484718
rect 519294 484398 519326 484634
rect 519562 484398 519646 484634
rect 519882 484398 519914 484634
rect 519294 448954 519914 484398
rect 519294 448718 519326 448954
rect 519562 448718 519646 448954
rect 519882 448718 519914 448954
rect 519294 448634 519914 448718
rect 519294 448398 519326 448634
rect 519562 448398 519646 448634
rect 519882 448398 519914 448634
rect 519294 412954 519914 448398
rect 519294 412718 519326 412954
rect 519562 412718 519646 412954
rect 519882 412718 519914 412954
rect 519294 412634 519914 412718
rect 519294 412398 519326 412634
rect 519562 412398 519646 412634
rect 519882 412398 519914 412634
rect 519294 376954 519914 412398
rect 519294 376718 519326 376954
rect 519562 376718 519646 376954
rect 519882 376718 519914 376954
rect 519294 376634 519914 376718
rect 519294 376398 519326 376634
rect 519562 376398 519646 376634
rect 519882 376398 519914 376634
rect 519294 340954 519914 376398
rect 519294 340718 519326 340954
rect 519562 340718 519646 340954
rect 519882 340718 519914 340954
rect 519294 340634 519914 340718
rect 519294 340398 519326 340634
rect 519562 340398 519646 340634
rect 519882 340398 519914 340634
rect 519294 304954 519914 340398
rect 519294 304718 519326 304954
rect 519562 304718 519646 304954
rect 519882 304718 519914 304954
rect 519294 304634 519914 304718
rect 519294 304398 519326 304634
rect 519562 304398 519646 304634
rect 519882 304398 519914 304634
rect 519294 268954 519914 304398
rect 519294 268718 519326 268954
rect 519562 268718 519646 268954
rect 519882 268718 519914 268954
rect 519294 268634 519914 268718
rect 519294 268398 519326 268634
rect 519562 268398 519646 268634
rect 519882 268398 519914 268634
rect 519294 232954 519914 268398
rect 519294 232718 519326 232954
rect 519562 232718 519646 232954
rect 519882 232718 519914 232954
rect 519294 232634 519914 232718
rect 519294 232398 519326 232634
rect 519562 232398 519646 232634
rect 519882 232398 519914 232634
rect 519294 196954 519914 232398
rect 519294 196718 519326 196954
rect 519562 196718 519646 196954
rect 519882 196718 519914 196954
rect 519294 196634 519914 196718
rect 519294 196398 519326 196634
rect 519562 196398 519646 196634
rect 519882 196398 519914 196634
rect 519294 160954 519914 196398
rect 519294 160718 519326 160954
rect 519562 160718 519646 160954
rect 519882 160718 519914 160954
rect 519294 160634 519914 160718
rect 519294 160398 519326 160634
rect 519562 160398 519646 160634
rect 519882 160398 519914 160634
rect 519294 124954 519914 160398
rect 519294 124718 519326 124954
rect 519562 124718 519646 124954
rect 519882 124718 519914 124954
rect 519294 124634 519914 124718
rect 519294 124398 519326 124634
rect 519562 124398 519646 124634
rect 519882 124398 519914 124634
rect 519294 88954 519914 124398
rect 519294 88718 519326 88954
rect 519562 88718 519646 88954
rect 519882 88718 519914 88954
rect 519294 88634 519914 88718
rect 519294 88398 519326 88634
rect 519562 88398 519646 88634
rect 519882 88398 519914 88634
rect 519294 52954 519914 88398
rect 519294 52718 519326 52954
rect 519562 52718 519646 52954
rect 519882 52718 519914 52954
rect 519294 52634 519914 52718
rect 519294 52398 519326 52634
rect 519562 52398 519646 52634
rect 519882 52398 519914 52634
rect 519294 16954 519914 52398
rect 519294 16718 519326 16954
rect 519562 16718 519646 16954
rect 519882 16718 519914 16954
rect 519294 16634 519914 16718
rect 519294 16398 519326 16634
rect 519562 16398 519646 16634
rect 519882 16398 519914 16634
rect 519294 -3226 519914 16398
rect 519294 -3462 519326 -3226
rect 519562 -3462 519646 -3226
rect 519882 -3462 519914 -3226
rect 519294 -3546 519914 -3462
rect 519294 -3782 519326 -3546
rect 519562 -3782 519646 -3546
rect 519882 -3782 519914 -3546
rect 519294 -7654 519914 -3782
rect 523794 708678 524414 711590
rect 523794 708442 523826 708678
rect 524062 708442 524146 708678
rect 524382 708442 524414 708678
rect 523794 708358 524414 708442
rect 523794 708122 523826 708358
rect 524062 708122 524146 708358
rect 524382 708122 524414 708358
rect 523794 669454 524414 708122
rect 523794 669218 523826 669454
rect 524062 669218 524146 669454
rect 524382 669218 524414 669454
rect 523794 669134 524414 669218
rect 523794 668898 523826 669134
rect 524062 668898 524146 669134
rect 524382 668898 524414 669134
rect 523794 633454 524414 668898
rect 523794 633218 523826 633454
rect 524062 633218 524146 633454
rect 524382 633218 524414 633454
rect 523794 633134 524414 633218
rect 523794 632898 523826 633134
rect 524062 632898 524146 633134
rect 524382 632898 524414 633134
rect 523794 597454 524414 632898
rect 523794 597218 523826 597454
rect 524062 597218 524146 597454
rect 524382 597218 524414 597454
rect 523794 597134 524414 597218
rect 523794 596898 523826 597134
rect 524062 596898 524146 597134
rect 524382 596898 524414 597134
rect 523794 561454 524414 596898
rect 523794 561218 523826 561454
rect 524062 561218 524146 561454
rect 524382 561218 524414 561454
rect 523794 561134 524414 561218
rect 523794 560898 523826 561134
rect 524062 560898 524146 561134
rect 524382 560898 524414 561134
rect 523794 525454 524414 560898
rect 523794 525218 523826 525454
rect 524062 525218 524146 525454
rect 524382 525218 524414 525454
rect 523794 525134 524414 525218
rect 523794 524898 523826 525134
rect 524062 524898 524146 525134
rect 524382 524898 524414 525134
rect 523794 489454 524414 524898
rect 523794 489218 523826 489454
rect 524062 489218 524146 489454
rect 524382 489218 524414 489454
rect 523794 489134 524414 489218
rect 523794 488898 523826 489134
rect 524062 488898 524146 489134
rect 524382 488898 524414 489134
rect 523794 453454 524414 488898
rect 523794 453218 523826 453454
rect 524062 453218 524146 453454
rect 524382 453218 524414 453454
rect 523794 453134 524414 453218
rect 523794 452898 523826 453134
rect 524062 452898 524146 453134
rect 524382 452898 524414 453134
rect 523794 417454 524414 452898
rect 523794 417218 523826 417454
rect 524062 417218 524146 417454
rect 524382 417218 524414 417454
rect 523794 417134 524414 417218
rect 523794 416898 523826 417134
rect 524062 416898 524146 417134
rect 524382 416898 524414 417134
rect 523794 381454 524414 416898
rect 523794 381218 523826 381454
rect 524062 381218 524146 381454
rect 524382 381218 524414 381454
rect 523794 381134 524414 381218
rect 523794 380898 523826 381134
rect 524062 380898 524146 381134
rect 524382 380898 524414 381134
rect 523794 345454 524414 380898
rect 523794 345218 523826 345454
rect 524062 345218 524146 345454
rect 524382 345218 524414 345454
rect 523794 345134 524414 345218
rect 523794 344898 523826 345134
rect 524062 344898 524146 345134
rect 524382 344898 524414 345134
rect 523794 309454 524414 344898
rect 523794 309218 523826 309454
rect 524062 309218 524146 309454
rect 524382 309218 524414 309454
rect 523794 309134 524414 309218
rect 523794 308898 523826 309134
rect 524062 308898 524146 309134
rect 524382 308898 524414 309134
rect 523794 273454 524414 308898
rect 523794 273218 523826 273454
rect 524062 273218 524146 273454
rect 524382 273218 524414 273454
rect 523794 273134 524414 273218
rect 523794 272898 523826 273134
rect 524062 272898 524146 273134
rect 524382 272898 524414 273134
rect 523794 237454 524414 272898
rect 523794 237218 523826 237454
rect 524062 237218 524146 237454
rect 524382 237218 524414 237454
rect 523794 237134 524414 237218
rect 523794 236898 523826 237134
rect 524062 236898 524146 237134
rect 524382 236898 524414 237134
rect 523794 201454 524414 236898
rect 523794 201218 523826 201454
rect 524062 201218 524146 201454
rect 524382 201218 524414 201454
rect 523794 201134 524414 201218
rect 523794 200898 523826 201134
rect 524062 200898 524146 201134
rect 524382 200898 524414 201134
rect 523794 165454 524414 200898
rect 523794 165218 523826 165454
rect 524062 165218 524146 165454
rect 524382 165218 524414 165454
rect 523794 165134 524414 165218
rect 523794 164898 523826 165134
rect 524062 164898 524146 165134
rect 524382 164898 524414 165134
rect 523794 129454 524414 164898
rect 523794 129218 523826 129454
rect 524062 129218 524146 129454
rect 524382 129218 524414 129454
rect 523794 129134 524414 129218
rect 523794 128898 523826 129134
rect 524062 128898 524146 129134
rect 524382 128898 524414 129134
rect 523794 93454 524414 128898
rect 523794 93218 523826 93454
rect 524062 93218 524146 93454
rect 524382 93218 524414 93454
rect 523794 93134 524414 93218
rect 523794 92898 523826 93134
rect 524062 92898 524146 93134
rect 524382 92898 524414 93134
rect 523794 57454 524414 92898
rect 523794 57218 523826 57454
rect 524062 57218 524146 57454
rect 524382 57218 524414 57454
rect 523794 57134 524414 57218
rect 523794 56898 523826 57134
rect 524062 56898 524146 57134
rect 524382 56898 524414 57134
rect 523794 21454 524414 56898
rect 523794 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 524414 21454
rect 523794 21134 524414 21218
rect 523794 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 524414 21134
rect 523794 -4186 524414 20898
rect 523794 -4422 523826 -4186
rect 524062 -4422 524146 -4186
rect 524382 -4422 524414 -4186
rect 523794 -4506 524414 -4422
rect 523794 -4742 523826 -4506
rect 524062 -4742 524146 -4506
rect 524382 -4742 524414 -4506
rect 523794 -7654 524414 -4742
rect 528294 709638 528914 711590
rect 528294 709402 528326 709638
rect 528562 709402 528646 709638
rect 528882 709402 528914 709638
rect 528294 709318 528914 709402
rect 528294 709082 528326 709318
rect 528562 709082 528646 709318
rect 528882 709082 528914 709318
rect 528294 673954 528914 709082
rect 528294 673718 528326 673954
rect 528562 673718 528646 673954
rect 528882 673718 528914 673954
rect 528294 673634 528914 673718
rect 528294 673398 528326 673634
rect 528562 673398 528646 673634
rect 528882 673398 528914 673634
rect 528294 637954 528914 673398
rect 528294 637718 528326 637954
rect 528562 637718 528646 637954
rect 528882 637718 528914 637954
rect 528294 637634 528914 637718
rect 528294 637398 528326 637634
rect 528562 637398 528646 637634
rect 528882 637398 528914 637634
rect 528294 601954 528914 637398
rect 528294 601718 528326 601954
rect 528562 601718 528646 601954
rect 528882 601718 528914 601954
rect 528294 601634 528914 601718
rect 528294 601398 528326 601634
rect 528562 601398 528646 601634
rect 528882 601398 528914 601634
rect 528294 565954 528914 601398
rect 528294 565718 528326 565954
rect 528562 565718 528646 565954
rect 528882 565718 528914 565954
rect 528294 565634 528914 565718
rect 528294 565398 528326 565634
rect 528562 565398 528646 565634
rect 528882 565398 528914 565634
rect 528294 529954 528914 565398
rect 528294 529718 528326 529954
rect 528562 529718 528646 529954
rect 528882 529718 528914 529954
rect 528294 529634 528914 529718
rect 528294 529398 528326 529634
rect 528562 529398 528646 529634
rect 528882 529398 528914 529634
rect 528294 493954 528914 529398
rect 528294 493718 528326 493954
rect 528562 493718 528646 493954
rect 528882 493718 528914 493954
rect 528294 493634 528914 493718
rect 528294 493398 528326 493634
rect 528562 493398 528646 493634
rect 528882 493398 528914 493634
rect 528294 457954 528914 493398
rect 528294 457718 528326 457954
rect 528562 457718 528646 457954
rect 528882 457718 528914 457954
rect 528294 457634 528914 457718
rect 528294 457398 528326 457634
rect 528562 457398 528646 457634
rect 528882 457398 528914 457634
rect 528294 421954 528914 457398
rect 528294 421718 528326 421954
rect 528562 421718 528646 421954
rect 528882 421718 528914 421954
rect 528294 421634 528914 421718
rect 528294 421398 528326 421634
rect 528562 421398 528646 421634
rect 528882 421398 528914 421634
rect 528294 385954 528914 421398
rect 528294 385718 528326 385954
rect 528562 385718 528646 385954
rect 528882 385718 528914 385954
rect 528294 385634 528914 385718
rect 528294 385398 528326 385634
rect 528562 385398 528646 385634
rect 528882 385398 528914 385634
rect 528294 349954 528914 385398
rect 528294 349718 528326 349954
rect 528562 349718 528646 349954
rect 528882 349718 528914 349954
rect 528294 349634 528914 349718
rect 528294 349398 528326 349634
rect 528562 349398 528646 349634
rect 528882 349398 528914 349634
rect 528294 313954 528914 349398
rect 528294 313718 528326 313954
rect 528562 313718 528646 313954
rect 528882 313718 528914 313954
rect 528294 313634 528914 313718
rect 528294 313398 528326 313634
rect 528562 313398 528646 313634
rect 528882 313398 528914 313634
rect 528294 277954 528914 313398
rect 528294 277718 528326 277954
rect 528562 277718 528646 277954
rect 528882 277718 528914 277954
rect 528294 277634 528914 277718
rect 528294 277398 528326 277634
rect 528562 277398 528646 277634
rect 528882 277398 528914 277634
rect 528294 241954 528914 277398
rect 528294 241718 528326 241954
rect 528562 241718 528646 241954
rect 528882 241718 528914 241954
rect 528294 241634 528914 241718
rect 528294 241398 528326 241634
rect 528562 241398 528646 241634
rect 528882 241398 528914 241634
rect 528294 205954 528914 241398
rect 528294 205718 528326 205954
rect 528562 205718 528646 205954
rect 528882 205718 528914 205954
rect 528294 205634 528914 205718
rect 528294 205398 528326 205634
rect 528562 205398 528646 205634
rect 528882 205398 528914 205634
rect 528294 169954 528914 205398
rect 528294 169718 528326 169954
rect 528562 169718 528646 169954
rect 528882 169718 528914 169954
rect 528294 169634 528914 169718
rect 528294 169398 528326 169634
rect 528562 169398 528646 169634
rect 528882 169398 528914 169634
rect 528294 133954 528914 169398
rect 528294 133718 528326 133954
rect 528562 133718 528646 133954
rect 528882 133718 528914 133954
rect 528294 133634 528914 133718
rect 528294 133398 528326 133634
rect 528562 133398 528646 133634
rect 528882 133398 528914 133634
rect 528294 97954 528914 133398
rect 528294 97718 528326 97954
rect 528562 97718 528646 97954
rect 528882 97718 528914 97954
rect 528294 97634 528914 97718
rect 528294 97398 528326 97634
rect 528562 97398 528646 97634
rect 528882 97398 528914 97634
rect 528294 61954 528914 97398
rect 528294 61718 528326 61954
rect 528562 61718 528646 61954
rect 528882 61718 528914 61954
rect 528294 61634 528914 61718
rect 528294 61398 528326 61634
rect 528562 61398 528646 61634
rect 528882 61398 528914 61634
rect 528294 25954 528914 61398
rect 528294 25718 528326 25954
rect 528562 25718 528646 25954
rect 528882 25718 528914 25954
rect 528294 25634 528914 25718
rect 528294 25398 528326 25634
rect 528562 25398 528646 25634
rect 528882 25398 528914 25634
rect 528294 -5146 528914 25398
rect 528294 -5382 528326 -5146
rect 528562 -5382 528646 -5146
rect 528882 -5382 528914 -5146
rect 528294 -5466 528914 -5382
rect 528294 -5702 528326 -5466
rect 528562 -5702 528646 -5466
rect 528882 -5702 528914 -5466
rect 528294 -7654 528914 -5702
rect 532794 710598 533414 711590
rect 532794 710362 532826 710598
rect 533062 710362 533146 710598
rect 533382 710362 533414 710598
rect 532794 710278 533414 710362
rect 532794 710042 532826 710278
rect 533062 710042 533146 710278
rect 533382 710042 533414 710278
rect 532794 678454 533414 710042
rect 532794 678218 532826 678454
rect 533062 678218 533146 678454
rect 533382 678218 533414 678454
rect 532794 678134 533414 678218
rect 532794 677898 532826 678134
rect 533062 677898 533146 678134
rect 533382 677898 533414 678134
rect 532794 642454 533414 677898
rect 532794 642218 532826 642454
rect 533062 642218 533146 642454
rect 533382 642218 533414 642454
rect 532794 642134 533414 642218
rect 532794 641898 532826 642134
rect 533062 641898 533146 642134
rect 533382 641898 533414 642134
rect 532794 606454 533414 641898
rect 532794 606218 532826 606454
rect 533062 606218 533146 606454
rect 533382 606218 533414 606454
rect 532794 606134 533414 606218
rect 532794 605898 532826 606134
rect 533062 605898 533146 606134
rect 533382 605898 533414 606134
rect 532794 570454 533414 605898
rect 532794 570218 532826 570454
rect 533062 570218 533146 570454
rect 533382 570218 533414 570454
rect 532794 570134 533414 570218
rect 532794 569898 532826 570134
rect 533062 569898 533146 570134
rect 533382 569898 533414 570134
rect 532794 534454 533414 569898
rect 532794 534218 532826 534454
rect 533062 534218 533146 534454
rect 533382 534218 533414 534454
rect 532794 534134 533414 534218
rect 532794 533898 532826 534134
rect 533062 533898 533146 534134
rect 533382 533898 533414 534134
rect 532794 498454 533414 533898
rect 532794 498218 532826 498454
rect 533062 498218 533146 498454
rect 533382 498218 533414 498454
rect 532794 498134 533414 498218
rect 532794 497898 532826 498134
rect 533062 497898 533146 498134
rect 533382 497898 533414 498134
rect 532794 462454 533414 497898
rect 532794 462218 532826 462454
rect 533062 462218 533146 462454
rect 533382 462218 533414 462454
rect 532794 462134 533414 462218
rect 532794 461898 532826 462134
rect 533062 461898 533146 462134
rect 533382 461898 533414 462134
rect 532794 426454 533414 461898
rect 532794 426218 532826 426454
rect 533062 426218 533146 426454
rect 533382 426218 533414 426454
rect 532794 426134 533414 426218
rect 532794 425898 532826 426134
rect 533062 425898 533146 426134
rect 533382 425898 533414 426134
rect 532794 390454 533414 425898
rect 532794 390218 532826 390454
rect 533062 390218 533146 390454
rect 533382 390218 533414 390454
rect 532794 390134 533414 390218
rect 532794 389898 532826 390134
rect 533062 389898 533146 390134
rect 533382 389898 533414 390134
rect 532794 354454 533414 389898
rect 532794 354218 532826 354454
rect 533062 354218 533146 354454
rect 533382 354218 533414 354454
rect 532794 354134 533414 354218
rect 532794 353898 532826 354134
rect 533062 353898 533146 354134
rect 533382 353898 533414 354134
rect 532794 318454 533414 353898
rect 532794 318218 532826 318454
rect 533062 318218 533146 318454
rect 533382 318218 533414 318454
rect 532794 318134 533414 318218
rect 532794 317898 532826 318134
rect 533062 317898 533146 318134
rect 533382 317898 533414 318134
rect 532794 282454 533414 317898
rect 532794 282218 532826 282454
rect 533062 282218 533146 282454
rect 533382 282218 533414 282454
rect 532794 282134 533414 282218
rect 532794 281898 532826 282134
rect 533062 281898 533146 282134
rect 533382 281898 533414 282134
rect 532794 246454 533414 281898
rect 532794 246218 532826 246454
rect 533062 246218 533146 246454
rect 533382 246218 533414 246454
rect 532794 246134 533414 246218
rect 532794 245898 532826 246134
rect 533062 245898 533146 246134
rect 533382 245898 533414 246134
rect 532794 210454 533414 245898
rect 532794 210218 532826 210454
rect 533062 210218 533146 210454
rect 533382 210218 533414 210454
rect 532794 210134 533414 210218
rect 532794 209898 532826 210134
rect 533062 209898 533146 210134
rect 533382 209898 533414 210134
rect 532794 174454 533414 209898
rect 532794 174218 532826 174454
rect 533062 174218 533146 174454
rect 533382 174218 533414 174454
rect 532794 174134 533414 174218
rect 532794 173898 532826 174134
rect 533062 173898 533146 174134
rect 533382 173898 533414 174134
rect 532794 138454 533414 173898
rect 532794 138218 532826 138454
rect 533062 138218 533146 138454
rect 533382 138218 533414 138454
rect 532794 138134 533414 138218
rect 532794 137898 532826 138134
rect 533062 137898 533146 138134
rect 533382 137898 533414 138134
rect 532794 102454 533414 137898
rect 532794 102218 532826 102454
rect 533062 102218 533146 102454
rect 533382 102218 533414 102454
rect 532794 102134 533414 102218
rect 532794 101898 532826 102134
rect 533062 101898 533146 102134
rect 533382 101898 533414 102134
rect 532794 66454 533414 101898
rect 532794 66218 532826 66454
rect 533062 66218 533146 66454
rect 533382 66218 533414 66454
rect 532794 66134 533414 66218
rect 532794 65898 532826 66134
rect 533062 65898 533146 66134
rect 533382 65898 533414 66134
rect 532794 30454 533414 65898
rect 532794 30218 532826 30454
rect 533062 30218 533146 30454
rect 533382 30218 533414 30454
rect 532794 30134 533414 30218
rect 532794 29898 532826 30134
rect 533062 29898 533146 30134
rect 533382 29898 533414 30134
rect 532794 -6106 533414 29898
rect 532794 -6342 532826 -6106
rect 533062 -6342 533146 -6106
rect 533382 -6342 533414 -6106
rect 532794 -6426 533414 -6342
rect 532794 -6662 532826 -6426
rect 533062 -6662 533146 -6426
rect 533382 -6662 533414 -6426
rect 532794 -7654 533414 -6662
rect 537294 711558 537914 711590
rect 537294 711322 537326 711558
rect 537562 711322 537646 711558
rect 537882 711322 537914 711558
rect 537294 711238 537914 711322
rect 537294 711002 537326 711238
rect 537562 711002 537646 711238
rect 537882 711002 537914 711238
rect 537294 682954 537914 711002
rect 537294 682718 537326 682954
rect 537562 682718 537646 682954
rect 537882 682718 537914 682954
rect 537294 682634 537914 682718
rect 537294 682398 537326 682634
rect 537562 682398 537646 682634
rect 537882 682398 537914 682634
rect 537294 646954 537914 682398
rect 537294 646718 537326 646954
rect 537562 646718 537646 646954
rect 537882 646718 537914 646954
rect 537294 646634 537914 646718
rect 537294 646398 537326 646634
rect 537562 646398 537646 646634
rect 537882 646398 537914 646634
rect 537294 610954 537914 646398
rect 537294 610718 537326 610954
rect 537562 610718 537646 610954
rect 537882 610718 537914 610954
rect 537294 610634 537914 610718
rect 537294 610398 537326 610634
rect 537562 610398 537646 610634
rect 537882 610398 537914 610634
rect 537294 574954 537914 610398
rect 537294 574718 537326 574954
rect 537562 574718 537646 574954
rect 537882 574718 537914 574954
rect 537294 574634 537914 574718
rect 537294 574398 537326 574634
rect 537562 574398 537646 574634
rect 537882 574398 537914 574634
rect 537294 538954 537914 574398
rect 537294 538718 537326 538954
rect 537562 538718 537646 538954
rect 537882 538718 537914 538954
rect 537294 538634 537914 538718
rect 537294 538398 537326 538634
rect 537562 538398 537646 538634
rect 537882 538398 537914 538634
rect 537294 502954 537914 538398
rect 537294 502718 537326 502954
rect 537562 502718 537646 502954
rect 537882 502718 537914 502954
rect 537294 502634 537914 502718
rect 537294 502398 537326 502634
rect 537562 502398 537646 502634
rect 537882 502398 537914 502634
rect 537294 466954 537914 502398
rect 537294 466718 537326 466954
rect 537562 466718 537646 466954
rect 537882 466718 537914 466954
rect 537294 466634 537914 466718
rect 537294 466398 537326 466634
rect 537562 466398 537646 466634
rect 537882 466398 537914 466634
rect 537294 430954 537914 466398
rect 537294 430718 537326 430954
rect 537562 430718 537646 430954
rect 537882 430718 537914 430954
rect 537294 430634 537914 430718
rect 537294 430398 537326 430634
rect 537562 430398 537646 430634
rect 537882 430398 537914 430634
rect 537294 394954 537914 430398
rect 537294 394718 537326 394954
rect 537562 394718 537646 394954
rect 537882 394718 537914 394954
rect 537294 394634 537914 394718
rect 537294 394398 537326 394634
rect 537562 394398 537646 394634
rect 537882 394398 537914 394634
rect 537294 358954 537914 394398
rect 537294 358718 537326 358954
rect 537562 358718 537646 358954
rect 537882 358718 537914 358954
rect 537294 358634 537914 358718
rect 537294 358398 537326 358634
rect 537562 358398 537646 358634
rect 537882 358398 537914 358634
rect 537294 322954 537914 358398
rect 537294 322718 537326 322954
rect 537562 322718 537646 322954
rect 537882 322718 537914 322954
rect 537294 322634 537914 322718
rect 537294 322398 537326 322634
rect 537562 322398 537646 322634
rect 537882 322398 537914 322634
rect 537294 286954 537914 322398
rect 537294 286718 537326 286954
rect 537562 286718 537646 286954
rect 537882 286718 537914 286954
rect 537294 286634 537914 286718
rect 537294 286398 537326 286634
rect 537562 286398 537646 286634
rect 537882 286398 537914 286634
rect 537294 250954 537914 286398
rect 537294 250718 537326 250954
rect 537562 250718 537646 250954
rect 537882 250718 537914 250954
rect 537294 250634 537914 250718
rect 537294 250398 537326 250634
rect 537562 250398 537646 250634
rect 537882 250398 537914 250634
rect 537294 214954 537914 250398
rect 537294 214718 537326 214954
rect 537562 214718 537646 214954
rect 537882 214718 537914 214954
rect 537294 214634 537914 214718
rect 537294 214398 537326 214634
rect 537562 214398 537646 214634
rect 537882 214398 537914 214634
rect 537294 178954 537914 214398
rect 537294 178718 537326 178954
rect 537562 178718 537646 178954
rect 537882 178718 537914 178954
rect 537294 178634 537914 178718
rect 537294 178398 537326 178634
rect 537562 178398 537646 178634
rect 537882 178398 537914 178634
rect 537294 142954 537914 178398
rect 537294 142718 537326 142954
rect 537562 142718 537646 142954
rect 537882 142718 537914 142954
rect 537294 142634 537914 142718
rect 537294 142398 537326 142634
rect 537562 142398 537646 142634
rect 537882 142398 537914 142634
rect 537294 106954 537914 142398
rect 537294 106718 537326 106954
rect 537562 106718 537646 106954
rect 537882 106718 537914 106954
rect 537294 106634 537914 106718
rect 537294 106398 537326 106634
rect 537562 106398 537646 106634
rect 537882 106398 537914 106634
rect 537294 70954 537914 106398
rect 537294 70718 537326 70954
rect 537562 70718 537646 70954
rect 537882 70718 537914 70954
rect 537294 70634 537914 70718
rect 537294 70398 537326 70634
rect 537562 70398 537646 70634
rect 537882 70398 537914 70634
rect 537294 34954 537914 70398
rect 537294 34718 537326 34954
rect 537562 34718 537646 34954
rect 537882 34718 537914 34954
rect 537294 34634 537914 34718
rect 537294 34398 537326 34634
rect 537562 34398 537646 34634
rect 537882 34398 537914 34634
rect 537294 -7066 537914 34398
rect 537294 -7302 537326 -7066
rect 537562 -7302 537646 -7066
rect 537882 -7302 537914 -7066
rect 537294 -7386 537914 -7302
rect 537294 -7622 537326 -7386
rect 537562 -7622 537646 -7386
rect 537882 -7622 537914 -7386
rect 537294 -7654 537914 -7622
rect 541794 704838 542414 711590
rect 541794 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 542414 704838
rect 541794 704518 542414 704602
rect 541794 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 542414 704518
rect 541794 687454 542414 704282
rect 541794 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 542414 687454
rect 541794 687134 542414 687218
rect 541794 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 542414 687134
rect 541794 651454 542414 686898
rect 541794 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 542414 651454
rect 541794 651134 542414 651218
rect 541794 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 542414 651134
rect 541794 615454 542414 650898
rect 541794 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 542414 615454
rect 541794 615134 542414 615218
rect 541794 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 542414 615134
rect 541794 579454 542414 614898
rect 541794 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 542414 579454
rect 541794 579134 542414 579218
rect 541794 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 542414 579134
rect 541794 543454 542414 578898
rect 541794 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 542414 543454
rect 541794 543134 542414 543218
rect 541794 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 542414 543134
rect 541794 507454 542414 542898
rect 541794 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 542414 507454
rect 541794 507134 542414 507218
rect 541794 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 542414 507134
rect 541794 471454 542414 506898
rect 541794 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 542414 471454
rect 541794 471134 542414 471218
rect 541794 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 542414 471134
rect 541794 435454 542414 470898
rect 541794 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 542414 435454
rect 541794 435134 542414 435218
rect 541794 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 542414 435134
rect 541794 399454 542414 434898
rect 541794 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 542414 399454
rect 541794 399134 542414 399218
rect 541794 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 542414 399134
rect 541794 363454 542414 398898
rect 541794 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 542414 363454
rect 541794 363134 542414 363218
rect 541794 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 542414 363134
rect 541794 327454 542414 362898
rect 541794 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 542414 327454
rect 541794 327134 542414 327218
rect 541794 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 542414 327134
rect 541794 291454 542414 326898
rect 541794 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 542414 291454
rect 541794 291134 542414 291218
rect 541794 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 542414 291134
rect 541794 255454 542414 290898
rect 541794 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 542414 255454
rect 541794 255134 542414 255218
rect 541794 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 542414 255134
rect 541794 219454 542414 254898
rect 541794 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 542414 219454
rect 541794 219134 542414 219218
rect 541794 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 542414 219134
rect 541794 183454 542414 218898
rect 541794 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 542414 183454
rect 541794 183134 542414 183218
rect 541794 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 542414 183134
rect 541794 147454 542414 182898
rect 541794 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 542414 147454
rect 541794 147134 542414 147218
rect 541794 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 542414 147134
rect 541794 111454 542414 146898
rect 541794 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 542414 111454
rect 541794 111134 542414 111218
rect 541794 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 542414 111134
rect 541794 75454 542414 110898
rect 541794 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 542414 75454
rect 541794 75134 542414 75218
rect 541794 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 542414 75134
rect 541794 39454 542414 74898
rect 541794 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 542414 39454
rect 541794 39134 542414 39218
rect 541794 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 542414 39134
rect 541794 3454 542414 38898
rect 541794 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 542414 3454
rect 541794 3134 542414 3218
rect 541794 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 542414 3134
rect 541794 -346 542414 2898
rect 541794 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 542414 -346
rect 541794 -666 542414 -582
rect 541794 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 542414 -666
rect 541794 -7654 542414 -902
rect 546294 705798 546914 711590
rect 546294 705562 546326 705798
rect 546562 705562 546646 705798
rect 546882 705562 546914 705798
rect 546294 705478 546914 705562
rect 546294 705242 546326 705478
rect 546562 705242 546646 705478
rect 546882 705242 546914 705478
rect 546294 691954 546914 705242
rect 546294 691718 546326 691954
rect 546562 691718 546646 691954
rect 546882 691718 546914 691954
rect 546294 691634 546914 691718
rect 546294 691398 546326 691634
rect 546562 691398 546646 691634
rect 546882 691398 546914 691634
rect 546294 655954 546914 691398
rect 546294 655718 546326 655954
rect 546562 655718 546646 655954
rect 546882 655718 546914 655954
rect 546294 655634 546914 655718
rect 546294 655398 546326 655634
rect 546562 655398 546646 655634
rect 546882 655398 546914 655634
rect 546294 619954 546914 655398
rect 546294 619718 546326 619954
rect 546562 619718 546646 619954
rect 546882 619718 546914 619954
rect 546294 619634 546914 619718
rect 546294 619398 546326 619634
rect 546562 619398 546646 619634
rect 546882 619398 546914 619634
rect 546294 583954 546914 619398
rect 546294 583718 546326 583954
rect 546562 583718 546646 583954
rect 546882 583718 546914 583954
rect 546294 583634 546914 583718
rect 546294 583398 546326 583634
rect 546562 583398 546646 583634
rect 546882 583398 546914 583634
rect 546294 547954 546914 583398
rect 546294 547718 546326 547954
rect 546562 547718 546646 547954
rect 546882 547718 546914 547954
rect 546294 547634 546914 547718
rect 546294 547398 546326 547634
rect 546562 547398 546646 547634
rect 546882 547398 546914 547634
rect 546294 511954 546914 547398
rect 546294 511718 546326 511954
rect 546562 511718 546646 511954
rect 546882 511718 546914 511954
rect 546294 511634 546914 511718
rect 546294 511398 546326 511634
rect 546562 511398 546646 511634
rect 546882 511398 546914 511634
rect 546294 475954 546914 511398
rect 546294 475718 546326 475954
rect 546562 475718 546646 475954
rect 546882 475718 546914 475954
rect 546294 475634 546914 475718
rect 546294 475398 546326 475634
rect 546562 475398 546646 475634
rect 546882 475398 546914 475634
rect 546294 439954 546914 475398
rect 546294 439718 546326 439954
rect 546562 439718 546646 439954
rect 546882 439718 546914 439954
rect 546294 439634 546914 439718
rect 546294 439398 546326 439634
rect 546562 439398 546646 439634
rect 546882 439398 546914 439634
rect 546294 403954 546914 439398
rect 546294 403718 546326 403954
rect 546562 403718 546646 403954
rect 546882 403718 546914 403954
rect 546294 403634 546914 403718
rect 546294 403398 546326 403634
rect 546562 403398 546646 403634
rect 546882 403398 546914 403634
rect 546294 367954 546914 403398
rect 546294 367718 546326 367954
rect 546562 367718 546646 367954
rect 546882 367718 546914 367954
rect 546294 367634 546914 367718
rect 546294 367398 546326 367634
rect 546562 367398 546646 367634
rect 546882 367398 546914 367634
rect 546294 331954 546914 367398
rect 546294 331718 546326 331954
rect 546562 331718 546646 331954
rect 546882 331718 546914 331954
rect 546294 331634 546914 331718
rect 546294 331398 546326 331634
rect 546562 331398 546646 331634
rect 546882 331398 546914 331634
rect 546294 295954 546914 331398
rect 546294 295718 546326 295954
rect 546562 295718 546646 295954
rect 546882 295718 546914 295954
rect 546294 295634 546914 295718
rect 546294 295398 546326 295634
rect 546562 295398 546646 295634
rect 546882 295398 546914 295634
rect 546294 259954 546914 295398
rect 546294 259718 546326 259954
rect 546562 259718 546646 259954
rect 546882 259718 546914 259954
rect 546294 259634 546914 259718
rect 546294 259398 546326 259634
rect 546562 259398 546646 259634
rect 546882 259398 546914 259634
rect 546294 223954 546914 259398
rect 546294 223718 546326 223954
rect 546562 223718 546646 223954
rect 546882 223718 546914 223954
rect 546294 223634 546914 223718
rect 546294 223398 546326 223634
rect 546562 223398 546646 223634
rect 546882 223398 546914 223634
rect 546294 187954 546914 223398
rect 546294 187718 546326 187954
rect 546562 187718 546646 187954
rect 546882 187718 546914 187954
rect 546294 187634 546914 187718
rect 546294 187398 546326 187634
rect 546562 187398 546646 187634
rect 546882 187398 546914 187634
rect 546294 151954 546914 187398
rect 546294 151718 546326 151954
rect 546562 151718 546646 151954
rect 546882 151718 546914 151954
rect 546294 151634 546914 151718
rect 546294 151398 546326 151634
rect 546562 151398 546646 151634
rect 546882 151398 546914 151634
rect 546294 115954 546914 151398
rect 546294 115718 546326 115954
rect 546562 115718 546646 115954
rect 546882 115718 546914 115954
rect 546294 115634 546914 115718
rect 546294 115398 546326 115634
rect 546562 115398 546646 115634
rect 546882 115398 546914 115634
rect 546294 79954 546914 115398
rect 546294 79718 546326 79954
rect 546562 79718 546646 79954
rect 546882 79718 546914 79954
rect 546294 79634 546914 79718
rect 546294 79398 546326 79634
rect 546562 79398 546646 79634
rect 546882 79398 546914 79634
rect 546294 43954 546914 79398
rect 546294 43718 546326 43954
rect 546562 43718 546646 43954
rect 546882 43718 546914 43954
rect 546294 43634 546914 43718
rect 546294 43398 546326 43634
rect 546562 43398 546646 43634
rect 546882 43398 546914 43634
rect 546294 7954 546914 43398
rect 546294 7718 546326 7954
rect 546562 7718 546646 7954
rect 546882 7718 546914 7954
rect 546294 7634 546914 7718
rect 546294 7398 546326 7634
rect 546562 7398 546646 7634
rect 546882 7398 546914 7634
rect 546294 -1306 546914 7398
rect 546294 -1542 546326 -1306
rect 546562 -1542 546646 -1306
rect 546882 -1542 546914 -1306
rect 546294 -1626 546914 -1542
rect 546294 -1862 546326 -1626
rect 546562 -1862 546646 -1626
rect 546882 -1862 546914 -1626
rect 546294 -7654 546914 -1862
rect 550794 706758 551414 711590
rect 550794 706522 550826 706758
rect 551062 706522 551146 706758
rect 551382 706522 551414 706758
rect 550794 706438 551414 706522
rect 550794 706202 550826 706438
rect 551062 706202 551146 706438
rect 551382 706202 551414 706438
rect 550794 696454 551414 706202
rect 550794 696218 550826 696454
rect 551062 696218 551146 696454
rect 551382 696218 551414 696454
rect 550794 696134 551414 696218
rect 550794 695898 550826 696134
rect 551062 695898 551146 696134
rect 551382 695898 551414 696134
rect 550794 660454 551414 695898
rect 550794 660218 550826 660454
rect 551062 660218 551146 660454
rect 551382 660218 551414 660454
rect 550794 660134 551414 660218
rect 550794 659898 550826 660134
rect 551062 659898 551146 660134
rect 551382 659898 551414 660134
rect 550794 624454 551414 659898
rect 550794 624218 550826 624454
rect 551062 624218 551146 624454
rect 551382 624218 551414 624454
rect 550794 624134 551414 624218
rect 550794 623898 550826 624134
rect 551062 623898 551146 624134
rect 551382 623898 551414 624134
rect 550794 588454 551414 623898
rect 550794 588218 550826 588454
rect 551062 588218 551146 588454
rect 551382 588218 551414 588454
rect 550794 588134 551414 588218
rect 550794 587898 550826 588134
rect 551062 587898 551146 588134
rect 551382 587898 551414 588134
rect 550794 552454 551414 587898
rect 550794 552218 550826 552454
rect 551062 552218 551146 552454
rect 551382 552218 551414 552454
rect 550794 552134 551414 552218
rect 550794 551898 550826 552134
rect 551062 551898 551146 552134
rect 551382 551898 551414 552134
rect 550794 516454 551414 551898
rect 550794 516218 550826 516454
rect 551062 516218 551146 516454
rect 551382 516218 551414 516454
rect 550794 516134 551414 516218
rect 550794 515898 550826 516134
rect 551062 515898 551146 516134
rect 551382 515898 551414 516134
rect 550794 480454 551414 515898
rect 550794 480218 550826 480454
rect 551062 480218 551146 480454
rect 551382 480218 551414 480454
rect 550794 480134 551414 480218
rect 550794 479898 550826 480134
rect 551062 479898 551146 480134
rect 551382 479898 551414 480134
rect 550794 444454 551414 479898
rect 550794 444218 550826 444454
rect 551062 444218 551146 444454
rect 551382 444218 551414 444454
rect 550794 444134 551414 444218
rect 550794 443898 550826 444134
rect 551062 443898 551146 444134
rect 551382 443898 551414 444134
rect 550794 408454 551414 443898
rect 550794 408218 550826 408454
rect 551062 408218 551146 408454
rect 551382 408218 551414 408454
rect 550794 408134 551414 408218
rect 550794 407898 550826 408134
rect 551062 407898 551146 408134
rect 551382 407898 551414 408134
rect 550794 372454 551414 407898
rect 550794 372218 550826 372454
rect 551062 372218 551146 372454
rect 551382 372218 551414 372454
rect 550794 372134 551414 372218
rect 550794 371898 550826 372134
rect 551062 371898 551146 372134
rect 551382 371898 551414 372134
rect 550794 336454 551414 371898
rect 550794 336218 550826 336454
rect 551062 336218 551146 336454
rect 551382 336218 551414 336454
rect 550794 336134 551414 336218
rect 550794 335898 550826 336134
rect 551062 335898 551146 336134
rect 551382 335898 551414 336134
rect 550794 300454 551414 335898
rect 550794 300218 550826 300454
rect 551062 300218 551146 300454
rect 551382 300218 551414 300454
rect 550794 300134 551414 300218
rect 550794 299898 550826 300134
rect 551062 299898 551146 300134
rect 551382 299898 551414 300134
rect 550794 264454 551414 299898
rect 550794 264218 550826 264454
rect 551062 264218 551146 264454
rect 551382 264218 551414 264454
rect 550794 264134 551414 264218
rect 550794 263898 550826 264134
rect 551062 263898 551146 264134
rect 551382 263898 551414 264134
rect 550794 228454 551414 263898
rect 550794 228218 550826 228454
rect 551062 228218 551146 228454
rect 551382 228218 551414 228454
rect 550794 228134 551414 228218
rect 550794 227898 550826 228134
rect 551062 227898 551146 228134
rect 551382 227898 551414 228134
rect 550794 192454 551414 227898
rect 550794 192218 550826 192454
rect 551062 192218 551146 192454
rect 551382 192218 551414 192454
rect 550794 192134 551414 192218
rect 550794 191898 550826 192134
rect 551062 191898 551146 192134
rect 551382 191898 551414 192134
rect 550794 156454 551414 191898
rect 550794 156218 550826 156454
rect 551062 156218 551146 156454
rect 551382 156218 551414 156454
rect 550794 156134 551414 156218
rect 550794 155898 550826 156134
rect 551062 155898 551146 156134
rect 551382 155898 551414 156134
rect 550794 120454 551414 155898
rect 550794 120218 550826 120454
rect 551062 120218 551146 120454
rect 551382 120218 551414 120454
rect 550794 120134 551414 120218
rect 550794 119898 550826 120134
rect 551062 119898 551146 120134
rect 551382 119898 551414 120134
rect 550794 84454 551414 119898
rect 550794 84218 550826 84454
rect 551062 84218 551146 84454
rect 551382 84218 551414 84454
rect 550794 84134 551414 84218
rect 550794 83898 550826 84134
rect 551062 83898 551146 84134
rect 551382 83898 551414 84134
rect 550794 48454 551414 83898
rect 550794 48218 550826 48454
rect 551062 48218 551146 48454
rect 551382 48218 551414 48454
rect 550794 48134 551414 48218
rect 550794 47898 550826 48134
rect 551062 47898 551146 48134
rect 551382 47898 551414 48134
rect 550794 12454 551414 47898
rect 550794 12218 550826 12454
rect 551062 12218 551146 12454
rect 551382 12218 551414 12454
rect 550794 12134 551414 12218
rect 550794 11898 550826 12134
rect 551062 11898 551146 12134
rect 551382 11898 551414 12134
rect 550794 -2266 551414 11898
rect 550794 -2502 550826 -2266
rect 551062 -2502 551146 -2266
rect 551382 -2502 551414 -2266
rect 550794 -2586 551414 -2502
rect 550794 -2822 550826 -2586
rect 551062 -2822 551146 -2586
rect 551382 -2822 551414 -2586
rect 550794 -7654 551414 -2822
rect 555294 707718 555914 711590
rect 555294 707482 555326 707718
rect 555562 707482 555646 707718
rect 555882 707482 555914 707718
rect 555294 707398 555914 707482
rect 555294 707162 555326 707398
rect 555562 707162 555646 707398
rect 555882 707162 555914 707398
rect 555294 700954 555914 707162
rect 555294 700718 555326 700954
rect 555562 700718 555646 700954
rect 555882 700718 555914 700954
rect 555294 700634 555914 700718
rect 555294 700398 555326 700634
rect 555562 700398 555646 700634
rect 555882 700398 555914 700634
rect 555294 664954 555914 700398
rect 555294 664718 555326 664954
rect 555562 664718 555646 664954
rect 555882 664718 555914 664954
rect 555294 664634 555914 664718
rect 555294 664398 555326 664634
rect 555562 664398 555646 664634
rect 555882 664398 555914 664634
rect 555294 628954 555914 664398
rect 555294 628718 555326 628954
rect 555562 628718 555646 628954
rect 555882 628718 555914 628954
rect 555294 628634 555914 628718
rect 555294 628398 555326 628634
rect 555562 628398 555646 628634
rect 555882 628398 555914 628634
rect 555294 592954 555914 628398
rect 555294 592718 555326 592954
rect 555562 592718 555646 592954
rect 555882 592718 555914 592954
rect 555294 592634 555914 592718
rect 555294 592398 555326 592634
rect 555562 592398 555646 592634
rect 555882 592398 555914 592634
rect 555294 556954 555914 592398
rect 555294 556718 555326 556954
rect 555562 556718 555646 556954
rect 555882 556718 555914 556954
rect 555294 556634 555914 556718
rect 555294 556398 555326 556634
rect 555562 556398 555646 556634
rect 555882 556398 555914 556634
rect 555294 520954 555914 556398
rect 555294 520718 555326 520954
rect 555562 520718 555646 520954
rect 555882 520718 555914 520954
rect 555294 520634 555914 520718
rect 555294 520398 555326 520634
rect 555562 520398 555646 520634
rect 555882 520398 555914 520634
rect 555294 484954 555914 520398
rect 555294 484718 555326 484954
rect 555562 484718 555646 484954
rect 555882 484718 555914 484954
rect 555294 484634 555914 484718
rect 555294 484398 555326 484634
rect 555562 484398 555646 484634
rect 555882 484398 555914 484634
rect 555294 448954 555914 484398
rect 555294 448718 555326 448954
rect 555562 448718 555646 448954
rect 555882 448718 555914 448954
rect 555294 448634 555914 448718
rect 555294 448398 555326 448634
rect 555562 448398 555646 448634
rect 555882 448398 555914 448634
rect 555294 412954 555914 448398
rect 555294 412718 555326 412954
rect 555562 412718 555646 412954
rect 555882 412718 555914 412954
rect 555294 412634 555914 412718
rect 555294 412398 555326 412634
rect 555562 412398 555646 412634
rect 555882 412398 555914 412634
rect 555294 376954 555914 412398
rect 555294 376718 555326 376954
rect 555562 376718 555646 376954
rect 555882 376718 555914 376954
rect 555294 376634 555914 376718
rect 555294 376398 555326 376634
rect 555562 376398 555646 376634
rect 555882 376398 555914 376634
rect 555294 340954 555914 376398
rect 555294 340718 555326 340954
rect 555562 340718 555646 340954
rect 555882 340718 555914 340954
rect 555294 340634 555914 340718
rect 555294 340398 555326 340634
rect 555562 340398 555646 340634
rect 555882 340398 555914 340634
rect 555294 304954 555914 340398
rect 555294 304718 555326 304954
rect 555562 304718 555646 304954
rect 555882 304718 555914 304954
rect 555294 304634 555914 304718
rect 555294 304398 555326 304634
rect 555562 304398 555646 304634
rect 555882 304398 555914 304634
rect 555294 268954 555914 304398
rect 555294 268718 555326 268954
rect 555562 268718 555646 268954
rect 555882 268718 555914 268954
rect 555294 268634 555914 268718
rect 555294 268398 555326 268634
rect 555562 268398 555646 268634
rect 555882 268398 555914 268634
rect 555294 232954 555914 268398
rect 555294 232718 555326 232954
rect 555562 232718 555646 232954
rect 555882 232718 555914 232954
rect 555294 232634 555914 232718
rect 555294 232398 555326 232634
rect 555562 232398 555646 232634
rect 555882 232398 555914 232634
rect 555294 196954 555914 232398
rect 555294 196718 555326 196954
rect 555562 196718 555646 196954
rect 555882 196718 555914 196954
rect 555294 196634 555914 196718
rect 555294 196398 555326 196634
rect 555562 196398 555646 196634
rect 555882 196398 555914 196634
rect 555294 160954 555914 196398
rect 555294 160718 555326 160954
rect 555562 160718 555646 160954
rect 555882 160718 555914 160954
rect 555294 160634 555914 160718
rect 555294 160398 555326 160634
rect 555562 160398 555646 160634
rect 555882 160398 555914 160634
rect 555294 124954 555914 160398
rect 555294 124718 555326 124954
rect 555562 124718 555646 124954
rect 555882 124718 555914 124954
rect 555294 124634 555914 124718
rect 555294 124398 555326 124634
rect 555562 124398 555646 124634
rect 555882 124398 555914 124634
rect 555294 88954 555914 124398
rect 555294 88718 555326 88954
rect 555562 88718 555646 88954
rect 555882 88718 555914 88954
rect 555294 88634 555914 88718
rect 555294 88398 555326 88634
rect 555562 88398 555646 88634
rect 555882 88398 555914 88634
rect 555294 52954 555914 88398
rect 555294 52718 555326 52954
rect 555562 52718 555646 52954
rect 555882 52718 555914 52954
rect 555294 52634 555914 52718
rect 555294 52398 555326 52634
rect 555562 52398 555646 52634
rect 555882 52398 555914 52634
rect 555294 16954 555914 52398
rect 555294 16718 555326 16954
rect 555562 16718 555646 16954
rect 555882 16718 555914 16954
rect 555294 16634 555914 16718
rect 555294 16398 555326 16634
rect 555562 16398 555646 16634
rect 555882 16398 555914 16634
rect 555294 -3226 555914 16398
rect 555294 -3462 555326 -3226
rect 555562 -3462 555646 -3226
rect 555882 -3462 555914 -3226
rect 555294 -3546 555914 -3462
rect 555294 -3782 555326 -3546
rect 555562 -3782 555646 -3546
rect 555882 -3782 555914 -3546
rect 555294 -7654 555914 -3782
rect 559794 708678 560414 711590
rect 559794 708442 559826 708678
rect 560062 708442 560146 708678
rect 560382 708442 560414 708678
rect 559794 708358 560414 708442
rect 559794 708122 559826 708358
rect 560062 708122 560146 708358
rect 560382 708122 560414 708358
rect 559794 669454 560414 708122
rect 559794 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 560414 669454
rect 559794 669134 560414 669218
rect 559794 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 560414 669134
rect 559794 633454 560414 668898
rect 559794 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 560414 633454
rect 559794 633134 560414 633218
rect 559794 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 560414 633134
rect 559794 597454 560414 632898
rect 559794 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 560414 597454
rect 559794 597134 560414 597218
rect 559794 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 560414 597134
rect 559794 561454 560414 596898
rect 559794 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 560414 561454
rect 559794 561134 560414 561218
rect 559794 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 560414 561134
rect 559794 525454 560414 560898
rect 559794 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 560414 525454
rect 559794 525134 560414 525218
rect 559794 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 560414 525134
rect 559794 489454 560414 524898
rect 559794 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 560414 489454
rect 559794 489134 560414 489218
rect 559794 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 560414 489134
rect 559794 453454 560414 488898
rect 559794 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 560414 453454
rect 559794 453134 560414 453218
rect 559794 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 560414 453134
rect 559794 417454 560414 452898
rect 559794 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 560414 417454
rect 559794 417134 560414 417218
rect 559794 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 560414 417134
rect 559794 381454 560414 416898
rect 559794 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 560414 381454
rect 559794 381134 560414 381218
rect 559794 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 560414 381134
rect 559794 345454 560414 380898
rect 559794 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 560414 345454
rect 559794 345134 560414 345218
rect 559794 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 560414 345134
rect 559794 309454 560414 344898
rect 559794 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 560414 309454
rect 559794 309134 560414 309218
rect 559794 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 560414 309134
rect 559794 273454 560414 308898
rect 559794 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 560414 273454
rect 559794 273134 560414 273218
rect 559794 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 560414 273134
rect 559794 237454 560414 272898
rect 559794 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 560414 237454
rect 559794 237134 560414 237218
rect 559794 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 560414 237134
rect 559794 201454 560414 236898
rect 559794 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 560414 201454
rect 559794 201134 560414 201218
rect 559794 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 560414 201134
rect 559794 165454 560414 200898
rect 559794 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 560414 165454
rect 559794 165134 560414 165218
rect 559794 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 560414 165134
rect 559794 129454 560414 164898
rect 559794 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 560414 129454
rect 559794 129134 560414 129218
rect 559794 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 560414 129134
rect 559794 93454 560414 128898
rect 559794 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 560414 93454
rect 559794 93134 560414 93218
rect 559794 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 560414 93134
rect 559794 57454 560414 92898
rect 559794 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 560414 57454
rect 559794 57134 560414 57218
rect 559794 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 560414 57134
rect 559794 21454 560414 56898
rect 559794 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 560414 21454
rect 559794 21134 560414 21218
rect 559794 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 560414 21134
rect 559794 -4186 560414 20898
rect 559794 -4422 559826 -4186
rect 560062 -4422 560146 -4186
rect 560382 -4422 560414 -4186
rect 559794 -4506 560414 -4422
rect 559794 -4742 559826 -4506
rect 560062 -4742 560146 -4506
rect 560382 -4742 560414 -4506
rect 559794 -7654 560414 -4742
rect 564294 709638 564914 711590
rect 564294 709402 564326 709638
rect 564562 709402 564646 709638
rect 564882 709402 564914 709638
rect 564294 709318 564914 709402
rect 564294 709082 564326 709318
rect 564562 709082 564646 709318
rect 564882 709082 564914 709318
rect 564294 673954 564914 709082
rect 564294 673718 564326 673954
rect 564562 673718 564646 673954
rect 564882 673718 564914 673954
rect 564294 673634 564914 673718
rect 564294 673398 564326 673634
rect 564562 673398 564646 673634
rect 564882 673398 564914 673634
rect 564294 637954 564914 673398
rect 564294 637718 564326 637954
rect 564562 637718 564646 637954
rect 564882 637718 564914 637954
rect 564294 637634 564914 637718
rect 564294 637398 564326 637634
rect 564562 637398 564646 637634
rect 564882 637398 564914 637634
rect 564294 601954 564914 637398
rect 564294 601718 564326 601954
rect 564562 601718 564646 601954
rect 564882 601718 564914 601954
rect 564294 601634 564914 601718
rect 564294 601398 564326 601634
rect 564562 601398 564646 601634
rect 564882 601398 564914 601634
rect 564294 565954 564914 601398
rect 564294 565718 564326 565954
rect 564562 565718 564646 565954
rect 564882 565718 564914 565954
rect 564294 565634 564914 565718
rect 564294 565398 564326 565634
rect 564562 565398 564646 565634
rect 564882 565398 564914 565634
rect 564294 529954 564914 565398
rect 564294 529718 564326 529954
rect 564562 529718 564646 529954
rect 564882 529718 564914 529954
rect 564294 529634 564914 529718
rect 564294 529398 564326 529634
rect 564562 529398 564646 529634
rect 564882 529398 564914 529634
rect 564294 493954 564914 529398
rect 564294 493718 564326 493954
rect 564562 493718 564646 493954
rect 564882 493718 564914 493954
rect 564294 493634 564914 493718
rect 564294 493398 564326 493634
rect 564562 493398 564646 493634
rect 564882 493398 564914 493634
rect 564294 457954 564914 493398
rect 564294 457718 564326 457954
rect 564562 457718 564646 457954
rect 564882 457718 564914 457954
rect 564294 457634 564914 457718
rect 564294 457398 564326 457634
rect 564562 457398 564646 457634
rect 564882 457398 564914 457634
rect 564294 421954 564914 457398
rect 564294 421718 564326 421954
rect 564562 421718 564646 421954
rect 564882 421718 564914 421954
rect 564294 421634 564914 421718
rect 564294 421398 564326 421634
rect 564562 421398 564646 421634
rect 564882 421398 564914 421634
rect 564294 385954 564914 421398
rect 564294 385718 564326 385954
rect 564562 385718 564646 385954
rect 564882 385718 564914 385954
rect 564294 385634 564914 385718
rect 564294 385398 564326 385634
rect 564562 385398 564646 385634
rect 564882 385398 564914 385634
rect 564294 349954 564914 385398
rect 564294 349718 564326 349954
rect 564562 349718 564646 349954
rect 564882 349718 564914 349954
rect 564294 349634 564914 349718
rect 564294 349398 564326 349634
rect 564562 349398 564646 349634
rect 564882 349398 564914 349634
rect 564294 313954 564914 349398
rect 564294 313718 564326 313954
rect 564562 313718 564646 313954
rect 564882 313718 564914 313954
rect 564294 313634 564914 313718
rect 564294 313398 564326 313634
rect 564562 313398 564646 313634
rect 564882 313398 564914 313634
rect 564294 277954 564914 313398
rect 564294 277718 564326 277954
rect 564562 277718 564646 277954
rect 564882 277718 564914 277954
rect 564294 277634 564914 277718
rect 564294 277398 564326 277634
rect 564562 277398 564646 277634
rect 564882 277398 564914 277634
rect 564294 241954 564914 277398
rect 564294 241718 564326 241954
rect 564562 241718 564646 241954
rect 564882 241718 564914 241954
rect 564294 241634 564914 241718
rect 564294 241398 564326 241634
rect 564562 241398 564646 241634
rect 564882 241398 564914 241634
rect 564294 205954 564914 241398
rect 564294 205718 564326 205954
rect 564562 205718 564646 205954
rect 564882 205718 564914 205954
rect 564294 205634 564914 205718
rect 564294 205398 564326 205634
rect 564562 205398 564646 205634
rect 564882 205398 564914 205634
rect 564294 169954 564914 205398
rect 564294 169718 564326 169954
rect 564562 169718 564646 169954
rect 564882 169718 564914 169954
rect 564294 169634 564914 169718
rect 564294 169398 564326 169634
rect 564562 169398 564646 169634
rect 564882 169398 564914 169634
rect 564294 133954 564914 169398
rect 564294 133718 564326 133954
rect 564562 133718 564646 133954
rect 564882 133718 564914 133954
rect 564294 133634 564914 133718
rect 564294 133398 564326 133634
rect 564562 133398 564646 133634
rect 564882 133398 564914 133634
rect 564294 97954 564914 133398
rect 564294 97718 564326 97954
rect 564562 97718 564646 97954
rect 564882 97718 564914 97954
rect 564294 97634 564914 97718
rect 564294 97398 564326 97634
rect 564562 97398 564646 97634
rect 564882 97398 564914 97634
rect 564294 61954 564914 97398
rect 564294 61718 564326 61954
rect 564562 61718 564646 61954
rect 564882 61718 564914 61954
rect 564294 61634 564914 61718
rect 564294 61398 564326 61634
rect 564562 61398 564646 61634
rect 564882 61398 564914 61634
rect 564294 25954 564914 61398
rect 564294 25718 564326 25954
rect 564562 25718 564646 25954
rect 564882 25718 564914 25954
rect 564294 25634 564914 25718
rect 564294 25398 564326 25634
rect 564562 25398 564646 25634
rect 564882 25398 564914 25634
rect 564294 -5146 564914 25398
rect 564294 -5382 564326 -5146
rect 564562 -5382 564646 -5146
rect 564882 -5382 564914 -5146
rect 564294 -5466 564914 -5382
rect 564294 -5702 564326 -5466
rect 564562 -5702 564646 -5466
rect 564882 -5702 564914 -5466
rect 564294 -7654 564914 -5702
rect 568794 710598 569414 711590
rect 568794 710362 568826 710598
rect 569062 710362 569146 710598
rect 569382 710362 569414 710598
rect 568794 710278 569414 710362
rect 568794 710042 568826 710278
rect 569062 710042 569146 710278
rect 569382 710042 569414 710278
rect 568794 678454 569414 710042
rect 568794 678218 568826 678454
rect 569062 678218 569146 678454
rect 569382 678218 569414 678454
rect 568794 678134 569414 678218
rect 568794 677898 568826 678134
rect 569062 677898 569146 678134
rect 569382 677898 569414 678134
rect 568794 642454 569414 677898
rect 568794 642218 568826 642454
rect 569062 642218 569146 642454
rect 569382 642218 569414 642454
rect 568794 642134 569414 642218
rect 568794 641898 568826 642134
rect 569062 641898 569146 642134
rect 569382 641898 569414 642134
rect 568794 606454 569414 641898
rect 568794 606218 568826 606454
rect 569062 606218 569146 606454
rect 569382 606218 569414 606454
rect 568794 606134 569414 606218
rect 568794 605898 568826 606134
rect 569062 605898 569146 606134
rect 569382 605898 569414 606134
rect 568794 570454 569414 605898
rect 568794 570218 568826 570454
rect 569062 570218 569146 570454
rect 569382 570218 569414 570454
rect 568794 570134 569414 570218
rect 568794 569898 568826 570134
rect 569062 569898 569146 570134
rect 569382 569898 569414 570134
rect 568794 534454 569414 569898
rect 568794 534218 568826 534454
rect 569062 534218 569146 534454
rect 569382 534218 569414 534454
rect 568794 534134 569414 534218
rect 568794 533898 568826 534134
rect 569062 533898 569146 534134
rect 569382 533898 569414 534134
rect 568794 498454 569414 533898
rect 568794 498218 568826 498454
rect 569062 498218 569146 498454
rect 569382 498218 569414 498454
rect 568794 498134 569414 498218
rect 568794 497898 568826 498134
rect 569062 497898 569146 498134
rect 569382 497898 569414 498134
rect 568794 462454 569414 497898
rect 568794 462218 568826 462454
rect 569062 462218 569146 462454
rect 569382 462218 569414 462454
rect 568794 462134 569414 462218
rect 568794 461898 568826 462134
rect 569062 461898 569146 462134
rect 569382 461898 569414 462134
rect 568794 426454 569414 461898
rect 568794 426218 568826 426454
rect 569062 426218 569146 426454
rect 569382 426218 569414 426454
rect 568794 426134 569414 426218
rect 568794 425898 568826 426134
rect 569062 425898 569146 426134
rect 569382 425898 569414 426134
rect 568794 390454 569414 425898
rect 568794 390218 568826 390454
rect 569062 390218 569146 390454
rect 569382 390218 569414 390454
rect 568794 390134 569414 390218
rect 568794 389898 568826 390134
rect 569062 389898 569146 390134
rect 569382 389898 569414 390134
rect 568794 354454 569414 389898
rect 568794 354218 568826 354454
rect 569062 354218 569146 354454
rect 569382 354218 569414 354454
rect 568794 354134 569414 354218
rect 568794 353898 568826 354134
rect 569062 353898 569146 354134
rect 569382 353898 569414 354134
rect 568794 318454 569414 353898
rect 568794 318218 568826 318454
rect 569062 318218 569146 318454
rect 569382 318218 569414 318454
rect 568794 318134 569414 318218
rect 568794 317898 568826 318134
rect 569062 317898 569146 318134
rect 569382 317898 569414 318134
rect 568794 282454 569414 317898
rect 568794 282218 568826 282454
rect 569062 282218 569146 282454
rect 569382 282218 569414 282454
rect 568794 282134 569414 282218
rect 568794 281898 568826 282134
rect 569062 281898 569146 282134
rect 569382 281898 569414 282134
rect 568794 246454 569414 281898
rect 568794 246218 568826 246454
rect 569062 246218 569146 246454
rect 569382 246218 569414 246454
rect 568794 246134 569414 246218
rect 568794 245898 568826 246134
rect 569062 245898 569146 246134
rect 569382 245898 569414 246134
rect 568794 210454 569414 245898
rect 568794 210218 568826 210454
rect 569062 210218 569146 210454
rect 569382 210218 569414 210454
rect 568794 210134 569414 210218
rect 568794 209898 568826 210134
rect 569062 209898 569146 210134
rect 569382 209898 569414 210134
rect 568794 174454 569414 209898
rect 568794 174218 568826 174454
rect 569062 174218 569146 174454
rect 569382 174218 569414 174454
rect 568794 174134 569414 174218
rect 568794 173898 568826 174134
rect 569062 173898 569146 174134
rect 569382 173898 569414 174134
rect 568794 138454 569414 173898
rect 568794 138218 568826 138454
rect 569062 138218 569146 138454
rect 569382 138218 569414 138454
rect 568794 138134 569414 138218
rect 568794 137898 568826 138134
rect 569062 137898 569146 138134
rect 569382 137898 569414 138134
rect 568794 102454 569414 137898
rect 568794 102218 568826 102454
rect 569062 102218 569146 102454
rect 569382 102218 569414 102454
rect 568794 102134 569414 102218
rect 568794 101898 568826 102134
rect 569062 101898 569146 102134
rect 569382 101898 569414 102134
rect 568794 66454 569414 101898
rect 568794 66218 568826 66454
rect 569062 66218 569146 66454
rect 569382 66218 569414 66454
rect 568794 66134 569414 66218
rect 568794 65898 568826 66134
rect 569062 65898 569146 66134
rect 569382 65898 569414 66134
rect 568794 30454 569414 65898
rect 568794 30218 568826 30454
rect 569062 30218 569146 30454
rect 569382 30218 569414 30454
rect 568794 30134 569414 30218
rect 568794 29898 568826 30134
rect 569062 29898 569146 30134
rect 569382 29898 569414 30134
rect 568794 -6106 569414 29898
rect 568794 -6342 568826 -6106
rect 569062 -6342 569146 -6106
rect 569382 -6342 569414 -6106
rect 568794 -6426 569414 -6342
rect 568794 -6662 568826 -6426
rect 569062 -6662 569146 -6426
rect 569382 -6662 569414 -6426
rect 568794 -7654 569414 -6662
rect 573294 711558 573914 711590
rect 573294 711322 573326 711558
rect 573562 711322 573646 711558
rect 573882 711322 573914 711558
rect 573294 711238 573914 711322
rect 573294 711002 573326 711238
rect 573562 711002 573646 711238
rect 573882 711002 573914 711238
rect 573294 682954 573914 711002
rect 573294 682718 573326 682954
rect 573562 682718 573646 682954
rect 573882 682718 573914 682954
rect 573294 682634 573914 682718
rect 573294 682398 573326 682634
rect 573562 682398 573646 682634
rect 573882 682398 573914 682634
rect 573294 646954 573914 682398
rect 573294 646718 573326 646954
rect 573562 646718 573646 646954
rect 573882 646718 573914 646954
rect 573294 646634 573914 646718
rect 573294 646398 573326 646634
rect 573562 646398 573646 646634
rect 573882 646398 573914 646634
rect 573294 610954 573914 646398
rect 573294 610718 573326 610954
rect 573562 610718 573646 610954
rect 573882 610718 573914 610954
rect 573294 610634 573914 610718
rect 573294 610398 573326 610634
rect 573562 610398 573646 610634
rect 573882 610398 573914 610634
rect 573294 574954 573914 610398
rect 573294 574718 573326 574954
rect 573562 574718 573646 574954
rect 573882 574718 573914 574954
rect 573294 574634 573914 574718
rect 573294 574398 573326 574634
rect 573562 574398 573646 574634
rect 573882 574398 573914 574634
rect 573294 538954 573914 574398
rect 573294 538718 573326 538954
rect 573562 538718 573646 538954
rect 573882 538718 573914 538954
rect 573294 538634 573914 538718
rect 573294 538398 573326 538634
rect 573562 538398 573646 538634
rect 573882 538398 573914 538634
rect 573294 502954 573914 538398
rect 573294 502718 573326 502954
rect 573562 502718 573646 502954
rect 573882 502718 573914 502954
rect 573294 502634 573914 502718
rect 573294 502398 573326 502634
rect 573562 502398 573646 502634
rect 573882 502398 573914 502634
rect 573294 466954 573914 502398
rect 573294 466718 573326 466954
rect 573562 466718 573646 466954
rect 573882 466718 573914 466954
rect 573294 466634 573914 466718
rect 573294 466398 573326 466634
rect 573562 466398 573646 466634
rect 573882 466398 573914 466634
rect 573294 430954 573914 466398
rect 573294 430718 573326 430954
rect 573562 430718 573646 430954
rect 573882 430718 573914 430954
rect 573294 430634 573914 430718
rect 573294 430398 573326 430634
rect 573562 430398 573646 430634
rect 573882 430398 573914 430634
rect 573294 394954 573914 430398
rect 573294 394718 573326 394954
rect 573562 394718 573646 394954
rect 573882 394718 573914 394954
rect 573294 394634 573914 394718
rect 573294 394398 573326 394634
rect 573562 394398 573646 394634
rect 573882 394398 573914 394634
rect 573294 358954 573914 394398
rect 573294 358718 573326 358954
rect 573562 358718 573646 358954
rect 573882 358718 573914 358954
rect 573294 358634 573914 358718
rect 573294 358398 573326 358634
rect 573562 358398 573646 358634
rect 573882 358398 573914 358634
rect 573294 322954 573914 358398
rect 573294 322718 573326 322954
rect 573562 322718 573646 322954
rect 573882 322718 573914 322954
rect 573294 322634 573914 322718
rect 573294 322398 573326 322634
rect 573562 322398 573646 322634
rect 573882 322398 573914 322634
rect 573294 286954 573914 322398
rect 573294 286718 573326 286954
rect 573562 286718 573646 286954
rect 573882 286718 573914 286954
rect 573294 286634 573914 286718
rect 573294 286398 573326 286634
rect 573562 286398 573646 286634
rect 573882 286398 573914 286634
rect 573294 250954 573914 286398
rect 573294 250718 573326 250954
rect 573562 250718 573646 250954
rect 573882 250718 573914 250954
rect 573294 250634 573914 250718
rect 573294 250398 573326 250634
rect 573562 250398 573646 250634
rect 573882 250398 573914 250634
rect 573294 214954 573914 250398
rect 573294 214718 573326 214954
rect 573562 214718 573646 214954
rect 573882 214718 573914 214954
rect 573294 214634 573914 214718
rect 573294 214398 573326 214634
rect 573562 214398 573646 214634
rect 573882 214398 573914 214634
rect 573294 178954 573914 214398
rect 573294 178718 573326 178954
rect 573562 178718 573646 178954
rect 573882 178718 573914 178954
rect 573294 178634 573914 178718
rect 573294 178398 573326 178634
rect 573562 178398 573646 178634
rect 573882 178398 573914 178634
rect 573294 142954 573914 178398
rect 573294 142718 573326 142954
rect 573562 142718 573646 142954
rect 573882 142718 573914 142954
rect 573294 142634 573914 142718
rect 573294 142398 573326 142634
rect 573562 142398 573646 142634
rect 573882 142398 573914 142634
rect 573294 106954 573914 142398
rect 573294 106718 573326 106954
rect 573562 106718 573646 106954
rect 573882 106718 573914 106954
rect 573294 106634 573914 106718
rect 573294 106398 573326 106634
rect 573562 106398 573646 106634
rect 573882 106398 573914 106634
rect 573294 70954 573914 106398
rect 573294 70718 573326 70954
rect 573562 70718 573646 70954
rect 573882 70718 573914 70954
rect 573294 70634 573914 70718
rect 573294 70398 573326 70634
rect 573562 70398 573646 70634
rect 573882 70398 573914 70634
rect 573294 34954 573914 70398
rect 573294 34718 573326 34954
rect 573562 34718 573646 34954
rect 573882 34718 573914 34954
rect 573294 34634 573914 34718
rect 573294 34398 573326 34634
rect 573562 34398 573646 34634
rect 573882 34398 573914 34634
rect 573294 -7066 573914 34398
rect 573294 -7302 573326 -7066
rect 573562 -7302 573646 -7066
rect 573882 -7302 573914 -7066
rect 573294 -7386 573914 -7302
rect 573294 -7622 573326 -7386
rect 573562 -7622 573646 -7386
rect 573882 -7622 573914 -7386
rect 573294 -7654 573914 -7622
rect 577794 704838 578414 711590
rect 577794 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 578414 704838
rect 577794 704518 578414 704602
rect 577794 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 578414 704518
rect 577794 687454 578414 704282
rect 577794 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 578414 687454
rect 577794 687134 578414 687218
rect 577794 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 578414 687134
rect 577794 651454 578414 686898
rect 577794 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 578414 651454
rect 577794 651134 578414 651218
rect 577794 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 578414 651134
rect 577794 615454 578414 650898
rect 577794 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 578414 615454
rect 577794 615134 578414 615218
rect 577794 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 578414 615134
rect 577794 579454 578414 614898
rect 577794 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 578414 579454
rect 577794 579134 578414 579218
rect 577794 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 578414 579134
rect 577794 543454 578414 578898
rect 577794 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 578414 543454
rect 577794 543134 578414 543218
rect 577794 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 578414 543134
rect 577794 507454 578414 542898
rect 577794 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 578414 507454
rect 577794 507134 578414 507218
rect 577794 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 578414 507134
rect 577794 471454 578414 506898
rect 577794 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 578414 471454
rect 577794 471134 578414 471218
rect 577794 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 578414 471134
rect 577794 435454 578414 470898
rect 577794 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 578414 435454
rect 577794 435134 578414 435218
rect 577794 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 578414 435134
rect 577794 399454 578414 434898
rect 577794 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 578414 399454
rect 577794 399134 578414 399218
rect 577794 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 578414 399134
rect 577794 363454 578414 398898
rect 577794 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 578414 363454
rect 577794 363134 578414 363218
rect 577794 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 578414 363134
rect 577794 327454 578414 362898
rect 577794 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 578414 327454
rect 577794 327134 578414 327218
rect 577794 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 578414 327134
rect 577794 291454 578414 326898
rect 577794 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 578414 291454
rect 577794 291134 578414 291218
rect 577794 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 578414 291134
rect 577794 255454 578414 290898
rect 577794 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 578414 255454
rect 577794 255134 578414 255218
rect 577794 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 578414 255134
rect 577794 219454 578414 254898
rect 577794 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 578414 219454
rect 577794 219134 578414 219218
rect 577794 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 578414 219134
rect 577794 183454 578414 218898
rect 577794 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 578414 183454
rect 577794 183134 578414 183218
rect 577794 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 578414 183134
rect 577794 147454 578414 182898
rect 577794 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 578414 147454
rect 577794 147134 578414 147218
rect 577794 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 578414 147134
rect 577794 111454 578414 146898
rect 577794 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 578414 111454
rect 577794 111134 578414 111218
rect 577794 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 578414 111134
rect 577794 75454 578414 110898
rect 577794 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 578414 75454
rect 577794 75134 578414 75218
rect 577794 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 578414 75134
rect 577794 39454 578414 74898
rect 577794 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 578414 39454
rect 577794 39134 578414 39218
rect 577794 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 578414 39134
rect 577794 3454 578414 38898
rect 577794 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 578414 3454
rect 577794 3134 578414 3218
rect 577794 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 578414 3134
rect 577794 -346 578414 2898
rect 577794 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 578414 -346
rect 577794 -666 578414 -582
rect 577794 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 578414 -666
rect 577794 -7654 578414 -902
rect 582294 705798 582914 711590
rect 592030 711558 592650 711590
rect 592030 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect 592030 711238 592650 711322
rect 592030 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect 591070 710598 591690 710630
rect 591070 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect 591070 710278 591690 710362
rect 591070 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect 590110 709638 590730 709670
rect 590110 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect 590110 709318 590730 709402
rect 590110 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect 589150 708678 589770 708710
rect 589150 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect 589150 708358 589770 708442
rect 589150 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect 588190 707718 588810 707750
rect 588190 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect 588190 707398 588810 707482
rect 588190 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect 587230 706758 587850 706790
rect 587230 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect 587230 706438 587850 706522
rect 587230 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect 582294 705562 582326 705798
rect 582562 705562 582646 705798
rect 582882 705562 582914 705798
rect 582294 705478 582914 705562
rect 582294 705242 582326 705478
rect 582562 705242 582646 705478
rect 582882 705242 582914 705478
rect 582294 691954 582914 705242
rect 586270 705798 586890 705830
rect 586270 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect 586270 705478 586890 705562
rect 586270 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect 582294 691718 582326 691954
rect 582562 691718 582646 691954
rect 582882 691718 582914 691954
rect 582294 691634 582914 691718
rect 582294 691398 582326 691634
rect 582562 691398 582646 691634
rect 582882 691398 582914 691634
rect 582294 655954 582914 691398
rect 582294 655718 582326 655954
rect 582562 655718 582646 655954
rect 582882 655718 582914 655954
rect 582294 655634 582914 655718
rect 582294 655398 582326 655634
rect 582562 655398 582646 655634
rect 582882 655398 582914 655634
rect 582294 619954 582914 655398
rect 582294 619718 582326 619954
rect 582562 619718 582646 619954
rect 582882 619718 582914 619954
rect 582294 619634 582914 619718
rect 582294 619398 582326 619634
rect 582562 619398 582646 619634
rect 582882 619398 582914 619634
rect 582294 583954 582914 619398
rect 582294 583718 582326 583954
rect 582562 583718 582646 583954
rect 582882 583718 582914 583954
rect 582294 583634 582914 583718
rect 582294 583398 582326 583634
rect 582562 583398 582646 583634
rect 582882 583398 582914 583634
rect 582294 547954 582914 583398
rect 582294 547718 582326 547954
rect 582562 547718 582646 547954
rect 582882 547718 582914 547954
rect 582294 547634 582914 547718
rect 582294 547398 582326 547634
rect 582562 547398 582646 547634
rect 582882 547398 582914 547634
rect 582294 511954 582914 547398
rect 582294 511718 582326 511954
rect 582562 511718 582646 511954
rect 582882 511718 582914 511954
rect 582294 511634 582914 511718
rect 582294 511398 582326 511634
rect 582562 511398 582646 511634
rect 582882 511398 582914 511634
rect 582294 475954 582914 511398
rect 582294 475718 582326 475954
rect 582562 475718 582646 475954
rect 582882 475718 582914 475954
rect 582294 475634 582914 475718
rect 582294 475398 582326 475634
rect 582562 475398 582646 475634
rect 582882 475398 582914 475634
rect 582294 439954 582914 475398
rect 582294 439718 582326 439954
rect 582562 439718 582646 439954
rect 582882 439718 582914 439954
rect 582294 439634 582914 439718
rect 582294 439398 582326 439634
rect 582562 439398 582646 439634
rect 582882 439398 582914 439634
rect 582294 403954 582914 439398
rect 582294 403718 582326 403954
rect 582562 403718 582646 403954
rect 582882 403718 582914 403954
rect 582294 403634 582914 403718
rect 582294 403398 582326 403634
rect 582562 403398 582646 403634
rect 582882 403398 582914 403634
rect 582294 367954 582914 403398
rect 582294 367718 582326 367954
rect 582562 367718 582646 367954
rect 582882 367718 582914 367954
rect 582294 367634 582914 367718
rect 582294 367398 582326 367634
rect 582562 367398 582646 367634
rect 582882 367398 582914 367634
rect 582294 331954 582914 367398
rect 582294 331718 582326 331954
rect 582562 331718 582646 331954
rect 582882 331718 582914 331954
rect 582294 331634 582914 331718
rect 582294 331398 582326 331634
rect 582562 331398 582646 331634
rect 582882 331398 582914 331634
rect 582294 295954 582914 331398
rect 582294 295718 582326 295954
rect 582562 295718 582646 295954
rect 582882 295718 582914 295954
rect 582294 295634 582914 295718
rect 582294 295398 582326 295634
rect 582562 295398 582646 295634
rect 582882 295398 582914 295634
rect 582294 259954 582914 295398
rect 582294 259718 582326 259954
rect 582562 259718 582646 259954
rect 582882 259718 582914 259954
rect 582294 259634 582914 259718
rect 582294 259398 582326 259634
rect 582562 259398 582646 259634
rect 582882 259398 582914 259634
rect 582294 223954 582914 259398
rect 582294 223718 582326 223954
rect 582562 223718 582646 223954
rect 582882 223718 582914 223954
rect 582294 223634 582914 223718
rect 582294 223398 582326 223634
rect 582562 223398 582646 223634
rect 582882 223398 582914 223634
rect 582294 187954 582914 223398
rect 582294 187718 582326 187954
rect 582562 187718 582646 187954
rect 582882 187718 582914 187954
rect 582294 187634 582914 187718
rect 582294 187398 582326 187634
rect 582562 187398 582646 187634
rect 582882 187398 582914 187634
rect 582294 151954 582914 187398
rect 582294 151718 582326 151954
rect 582562 151718 582646 151954
rect 582882 151718 582914 151954
rect 582294 151634 582914 151718
rect 582294 151398 582326 151634
rect 582562 151398 582646 151634
rect 582882 151398 582914 151634
rect 582294 115954 582914 151398
rect 582294 115718 582326 115954
rect 582562 115718 582646 115954
rect 582882 115718 582914 115954
rect 582294 115634 582914 115718
rect 582294 115398 582326 115634
rect 582562 115398 582646 115634
rect 582882 115398 582914 115634
rect 582294 79954 582914 115398
rect 582294 79718 582326 79954
rect 582562 79718 582646 79954
rect 582882 79718 582914 79954
rect 582294 79634 582914 79718
rect 582294 79398 582326 79634
rect 582562 79398 582646 79634
rect 582882 79398 582914 79634
rect 582294 43954 582914 79398
rect 582294 43718 582326 43954
rect 582562 43718 582646 43954
rect 582882 43718 582914 43954
rect 582294 43634 582914 43718
rect 582294 43398 582326 43634
rect 582562 43398 582646 43634
rect 582882 43398 582914 43634
rect 582294 7954 582914 43398
rect 582294 7718 582326 7954
rect 582562 7718 582646 7954
rect 582882 7718 582914 7954
rect 582294 7634 582914 7718
rect 582294 7398 582326 7634
rect 582562 7398 582646 7634
rect 582882 7398 582914 7634
rect 582294 -1306 582914 7398
rect 585310 704838 585930 704870
rect 585310 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect 585310 704518 585930 704602
rect 585310 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect 585310 687454 585930 704282
rect 585310 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 585930 687454
rect 585310 687134 585930 687218
rect 585310 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 585930 687134
rect 585310 651454 585930 686898
rect 585310 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 585930 651454
rect 585310 651134 585930 651218
rect 585310 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 585930 651134
rect 585310 615454 585930 650898
rect 585310 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 585930 615454
rect 585310 615134 585930 615218
rect 585310 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 585930 615134
rect 585310 579454 585930 614898
rect 585310 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 585930 579454
rect 585310 579134 585930 579218
rect 585310 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 585930 579134
rect 585310 543454 585930 578898
rect 585310 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 585930 543454
rect 585310 543134 585930 543218
rect 585310 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 585930 543134
rect 585310 507454 585930 542898
rect 585310 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 585930 507454
rect 585310 507134 585930 507218
rect 585310 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 585930 507134
rect 585310 471454 585930 506898
rect 585310 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 585930 471454
rect 585310 471134 585930 471218
rect 585310 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 585930 471134
rect 585310 435454 585930 470898
rect 585310 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 585930 435454
rect 585310 435134 585930 435218
rect 585310 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 585930 435134
rect 585310 399454 585930 434898
rect 585310 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 585930 399454
rect 585310 399134 585930 399218
rect 585310 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 585930 399134
rect 585310 363454 585930 398898
rect 585310 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 585930 363454
rect 585310 363134 585930 363218
rect 585310 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 585930 363134
rect 585310 327454 585930 362898
rect 585310 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 585930 327454
rect 585310 327134 585930 327218
rect 585310 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 585930 327134
rect 585310 291454 585930 326898
rect 585310 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 585930 291454
rect 585310 291134 585930 291218
rect 585310 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 585930 291134
rect 585310 255454 585930 290898
rect 585310 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 585930 255454
rect 585310 255134 585930 255218
rect 585310 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 585930 255134
rect 585310 219454 585930 254898
rect 585310 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 585930 219454
rect 585310 219134 585930 219218
rect 585310 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 585930 219134
rect 585310 183454 585930 218898
rect 585310 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 585930 183454
rect 585310 183134 585930 183218
rect 585310 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 585930 183134
rect 585310 147454 585930 182898
rect 585310 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 585930 147454
rect 585310 147134 585930 147218
rect 585310 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 585930 147134
rect 585310 111454 585930 146898
rect 585310 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 585930 111454
rect 585310 111134 585930 111218
rect 585310 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 585930 111134
rect 585310 75454 585930 110898
rect 585310 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 585930 75454
rect 585310 75134 585930 75218
rect 585310 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 585930 75134
rect 585310 39454 585930 74898
rect 585310 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 585930 39454
rect 585310 39134 585930 39218
rect 585310 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 585930 39134
rect 585310 3454 585930 38898
rect 585310 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 585930 3454
rect 585310 3134 585930 3218
rect 585310 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 585930 3134
rect 585310 -346 585930 2898
rect 585310 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect 585310 -666 585930 -582
rect 585310 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect 585310 -934 585930 -902
rect 586270 691954 586890 705242
rect 586270 691718 586302 691954
rect 586538 691718 586622 691954
rect 586858 691718 586890 691954
rect 586270 691634 586890 691718
rect 586270 691398 586302 691634
rect 586538 691398 586622 691634
rect 586858 691398 586890 691634
rect 586270 655954 586890 691398
rect 586270 655718 586302 655954
rect 586538 655718 586622 655954
rect 586858 655718 586890 655954
rect 586270 655634 586890 655718
rect 586270 655398 586302 655634
rect 586538 655398 586622 655634
rect 586858 655398 586890 655634
rect 586270 619954 586890 655398
rect 586270 619718 586302 619954
rect 586538 619718 586622 619954
rect 586858 619718 586890 619954
rect 586270 619634 586890 619718
rect 586270 619398 586302 619634
rect 586538 619398 586622 619634
rect 586858 619398 586890 619634
rect 586270 583954 586890 619398
rect 586270 583718 586302 583954
rect 586538 583718 586622 583954
rect 586858 583718 586890 583954
rect 586270 583634 586890 583718
rect 586270 583398 586302 583634
rect 586538 583398 586622 583634
rect 586858 583398 586890 583634
rect 586270 547954 586890 583398
rect 586270 547718 586302 547954
rect 586538 547718 586622 547954
rect 586858 547718 586890 547954
rect 586270 547634 586890 547718
rect 586270 547398 586302 547634
rect 586538 547398 586622 547634
rect 586858 547398 586890 547634
rect 586270 511954 586890 547398
rect 586270 511718 586302 511954
rect 586538 511718 586622 511954
rect 586858 511718 586890 511954
rect 586270 511634 586890 511718
rect 586270 511398 586302 511634
rect 586538 511398 586622 511634
rect 586858 511398 586890 511634
rect 586270 475954 586890 511398
rect 586270 475718 586302 475954
rect 586538 475718 586622 475954
rect 586858 475718 586890 475954
rect 586270 475634 586890 475718
rect 586270 475398 586302 475634
rect 586538 475398 586622 475634
rect 586858 475398 586890 475634
rect 586270 439954 586890 475398
rect 586270 439718 586302 439954
rect 586538 439718 586622 439954
rect 586858 439718 586890 439954
rect 586270 439634 586890 439718
rect 586270 439398 586302 439634
rect 586538 439398 586622 439634
rect 586858 439398 586890 439634
rect 586270 403954 586890 439398
rect 586270 403718 586302 403954
rect 586538 403718 586622 403954
rect 586858 403718 586890 403954
rect 586270 403634 586890 403718
rect 586270 403398 586302 403634
rect 586538 403398 586622 403634
rect 586858 403398 586890 403634
rect 586270 367954 586890 403398
rect 586270 367718 586302 367954
rect 586538 367718 586622 367954
rect 586858 367718 586890 367954
rect 586270 367634 586890 367718
rect 586270 367398 586302 367634
rect 586538 367398 586622 367634
rect 586858 367398 586890 367634
rect 586270 331954 586890 367398
rect 586270 331718 586302 331954
rect 586538 331718 586622 331954
rect 586858 331718 586890 331954
rect 586270 331634 586890 331718
rect 586270 331398 586302 331634
rect 586538 331398 586622 331634
rect 586858 331398 586890 331634
rect 586270 295954 586890 331398
rect 586270 295718 586302 295954
rect 586538 295718 586622 295954
rect 586858 295718 586890 295954
rect 586270 295634 586890 295718
rect 586270 295398 586302 295634
rect 586538 295398 586622 295634
rect 586858 295398 586890 295634
rect 586270 259954 586890 295398
rect 586270 259718 586302 259954
rect 586538 259718 586622 259954
rect 586858 259718 586890 259954
rect 586270 259634 586890 259718
rect 586270 259398 586302 259634
rect 586538 259398 586622 259634
rect 586858 259398 586890 259634
rect 586270 223954 586890 259398
rect 586270 223718 586302 223954
rect 586538 223718 586622 223954
rect 586858 223718 586890 223954
rect 586270 223634 586890 223718
rect 586270 223398 586302 223634
rect 586538 223398 586622 223634
rect 586858 223398 586890 223634
rect 586270 187954 586890 223398
rect 586270 187718 586302 187954
rect 586538 187718 586622 187954
rect 586858 187718 586890 187954
rect 586270 187634 586890 187718
rect 586270 187398 586302 187634
rect 586538 187398 586622 187634
rect 586858 187398 586890 187634
rect 586270 151954 586890 187398
rect 586270 151718 586302 151954
rect 586538 151718 586622 151954
rect 586858 151718 586890 151954
rect 586270 151634 586890 151718
rect 586270 151398 586302 151634
rect 586538 151398 586622 151634
rect 586858 151398 586890 151634
rect 586270 115954 586890 151398
rect 586270 115718 586302 115954
rect 586538 115718 586622 115954
rect 586858 115718 586890 115954
rect 586270 115634 586890 115718
rect 586270 115398 586302 115634
rect 586538 115398 586622 115634
rect 586858 115398 586890 115634
rect 586270 79954 586890 115398
rect 586270 79718 586302 79954
rect 586538 79718 586622 79954
rect 586858 79718 586890 79954
rect 586270 79634 586890 79718
rect 586270 79398 586302 79634
rect 586538 79398 586622 79634
rect 586858 79398 586890 79634
rect 586270 43954 586890 79398
rect 586270 43718 586302 43954
rect 586538 43718 586622 43954
rect 586858 43718 586890 43954
rect 586270 43634 586890 43718
rect 586270 43398 586302 43634
rect 586538 43398 586622 43634
rect 586858 43398 586890 43634
rect 586270 7954 586890 43398
rect 586270 7718 586302 7954
rect 586538 7718 586622 7954
rect 586858 7718 586890 7954
rect 586270 7634 586890 7718
rect 586270 7398 586302 7634
rect 586538 7398 586622 7634
rect 586858 7398 586890 7634
rect 582294 -1542 582326 -1306
rect 582562 -1542 582646 -1306
rect 582882 -1542 582914 -1306
rect 582294 -1626 582914 -1542
rect 582294 -1862 582326 -1626
rect 582562 -1862 582646 -1626
rect 582882 -1862 582914 -1626
rect 582294 -7654 582914 -1862
rect 586270 -1306 586890 7398
rect 586270 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect 586270 -1626 586890 -1542
rect 586270 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect 586270 -1894 586890 -1862
rect 587230 696454 587850 706202
rect 587230 696218 587262 696454
rect 587498 696218 587582 696454
rect 587818 696218 587850 696454
rect 587230 696134 587850 696218
rect 587230 695898 587262 696134
rect 587498 695898 587582 696134
rect 587818 695898 587850 696134
rect 587230 660454 587850 695898
rect 587230 660218 587262 660454
rect 587498 660218 587582 660454
rect 587818 660218 587850 660454
rect 587230 660134 587850 660218
rect 587230 659898 587262 660134
rect 587498 659898 587582 660134
rect 587818 659898 587850 660134
rect 587230 624454 587850 659898
rect 587230 624218 587262 624454
rect 587498 624218 587582 624454
rect 587818 624218 587850 624454
rect 587230 624134 587850 624218
rect 587230 623898 587262 624134
rect 587498 623898 587582 624134
rect 587818 623898 587850 624134
rect 587230 588454 587850 623898
rect 587230 588218 587262 588454
rect 587498 588218 587582 588454
rect 587818 588218 587850 588454
rect 587230 588134 587850 588218
rect 587230 587898 587262 588134
rect 587498 587898 587582 588134
rect 587818 587898 587850 588134
rect 587230 552454 587850 587898
rect 587230 552218 587262 552454
rect 587498 552218 587582 552454
rect 587818 552218 587850 552454
rect 587230 552134 587850 552218
rect 587230 551898 587262 552134
rect 587498 551898 587582 552134
rect 587818 551898 587850 552134
rect 587230 516454 587850 551898
rect 587230 516218 587262 516454
rect 587498 516218 587582 516454
rect 587818 516218 587850 516454
rect 587230 516134 587850 516218
rect 587230 515898 587262 516134
rect 587498 515898 587582 516134
rect 587818 515898 587850 516134
rect 587230 480454 587850 515898
rect 587230 480218 587262 480454
rect 587498 480218 587582 480454
rect 587818 480218 587850 480454
rect 587230 480134 587850 480218
rect 587230 479898 587262 480134
rect 587498 479898 587582 480134
rect 587818 479898 587850 480134
rect 587230 444454 587850 479898
rect 587230 444218 587262 444454
rect 587498 444218 587582 444454
rect 587818 444218 587850 444454
rect 587230 444134 587850 444218
rect 587230 443898 587262 444134
rect 587498 443898 587582 444134
rect 587818 443898 587850 444134
rect 587230 408454 587850 443898
rect 587230 408218 587262 408454
rect 587498 408218 587582 408454
rect 587818 408218 587850 408454
rect 587230 408134 587850 408218
rect 587230 407898 587262 408134
rect 587498 407898 587582 408134
rect 587818 407898 587850 408134
rect 587230 372454 587850 407898
rect 587230 372218 587262 372454
rect 587498 372218 587582 372454
rect 587818 372218 587850 372454
rect 587230 372134 587850 372218
rect 587230 371898 587262 372134
rect 587498 371898 587582 372134
rect 587818 371898 587850 372134
rect 587230 336454 587850 371898
rect 587230 336218 587262 336454
rect 587498 336218 587582 336454
rect 587818 336218 587850 336454
rect 587230 336134 587850 336218
rect 587230 335898 587262 336134
rect 587498 335898 587582 336134
rect 587818 335898 587850 336134
rect 587230 300454 587850 335898
rect 587230 300218 587262 300454
rect 587498 300218 587582 300454
rect 587818 300218 587850 300454
rect 587230 300134 587850 300218
rect 587230 299898 587262 300134
rect 587498 299898 587582 300134
rect 587818 299898 587850 300134
rect 587230 264454 587850 299898
rect 587230 264218 587262 264454
rect 587498 264218 587582 264454
rect 587818 264218 587850 264454
rect 587230 264134 587850 264218
rect 587230 263898 587262 264134
rect 587498 263898 587582 264134
rect 587818 263898 587850 264134
rect 587230 228454 587850 263898
rect 587230 228218 587262 228454
rect 587498 228218 587582 228454
rect 587818 228218 587850 228454
rect 587230 228134 587850 228218
rect 587230 227898 587262 228134
rect 587498 227898 587582 228134
rect 587818 227898 587850 228134
rect 587230 192454 587850 227898
rect 587230 192218 587262 192454
rect 587498 192218 587582 192454
rect 587818 192218 587850 192454
rect 587230 192134 587850 192218
rect 587230 191898 587262 192134
rect 587498 191898 587582 192134
rect 587818 191898 587850 192134
rect 587230 156454 587850 191898
rect 587230 156218 587262 156454
rect 587498 156218 587582 156454
rect 587818 156218 587850 156454
rect 587230 156134 587850 156218
rect 587230 155898 587262 156134
rect 587498 155898 587582 156134
rect 587818 155898 587850 156134
rect 587230 120454 587850 155898
rect 587230 120218 587262 120454
rect 587498 120218 587582 120454
rect 587818 120218 587850 120454
rect 587230 120134 587850 120218
rect 587230 119898 587262 120134
rect 587498 119898 587582 120134
rect 587818 119898 587850 120134
rect 587230 84454 587850 119898
rect 587230 84218 587262 84454
rect 587498 84218 587582 84454
rect 587818 84218 587850 84454
rect 587230 84134 587850 84218
rect 587230 83898 587262 84134
rect 587498 83898 587582 84134
rect 587818 83898 587850 84134
rect 587230 48454 587850 83898
rect 587230 48218 587262 48454
rect 587498 48218 587582 48454
rect 587818 48218 587850 48454
rect 587230 48134 587850 48218
rect 587230 47898 587262 48134
rect 587498 47898 587582 48134
rect 587818 47898 587850 48134
rect 587230 12454 587850 47898
rect 587230 12218 587262 12454
rect 587498 12218 587582 12454
rect 587818 12218 587850 12454
rect 587230 12134 587850 12218
rect 587230 11898 587262 12134
rect 587498 11898 587582 12134
rect 587818 11898 587850 12134
rect 587230 -2266 587850 11898
rect 587230 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect 587230 -2586 587850 -2502
rect 587230 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect 587230 -2854 587850 -2822
rect 588190 700954 588810 707162
rect 588190 700718 588222 700954
rect 588458 700718 588542 700954
rect 588778 700718 588810 700954
rect 588190 700634 588810 700718
rect 588190 700398 588222 700634
rect 588458 700398 588542 700634
rect 588778 700398 588810 700634
rect 588190 664954 588810 700398
rect 588190 664718 588222 664954
rect 588458 664718 588542 664954
rect 588778 664718 588810 664954
rect 588190 664634 588810 664718
rect 588190 664398 588222 664634
rect 588458 664398 588542 664634
rect 588778 664398 588810 664634
rect 588190 628954 588810 664398
rect 588190 628718 588222 628954
rect 588458 628718 588542 628954
rect 588778 628718 588810 628954
rect 588190 628634 588810 628718
rect 588190 628398 588222 628634
rect 588458 628398 588542 628634
rect 588778 628398 588810 628634
rect 588190 592954 588810 628398
rect 588190 592718 588222 592954
rect 588458 592718 588542 592954
rect 588778 592718 588810 592954
rect 588190 592634 588810 592718
rect 588190 592398 588222 592634
rect 588458 592398 588542 592634
rect 588778 592398 588810 592634
rect 588190 556954 588810 592398
rect 588190 556718 588222 556954
rect 588458 556718 588542 556954
rect 588778 556718 588810 556954
rect 588190 556634 588810 556718
rect 588190 556398 588222 556634
rect 588458 556398 588542 556634
rect 588778 556398 588810 556634
rect 588190 520954 588810 556398
rect 588190 520718 588222 520954
rect 588458 520718 588542 520954
rect 588778 520718 588810 520954
rect 588190 520634 588810 520718
rect 588190 520398 588222 520634
rect 588458 520398 588542 520634
rect 588778 520398 588810 520634
rect 588190 484954 588810 520398
rect 588190 484718 588222 484954
rect 588458 484718 588542 484954
rect 588778 484718 588810 484954
rect 588190 484634 588810 484718
rect 588190 484398 588222 484634
rect 588458 484398 588542 484634
rect 588778 484398 588810 484634
rect 588190 448954 588810 484398
rect 588190 448718 588222 448954
rect 588458 448718 588542 448954
rect 588778 448718 588810 448954
rect 588190 448634 588810 448718
rect 588190 448398 588222 448634
rect 588458 448398 588542 448634
rect 588778 448398 588810 448634
rect 588190 412954 588810 448398
rect 588190 412718 588222 412954
rect 588458 412718 588542 412954
rect 588778 412718 588810 412954
rect 588190 412634 588810 412718
rect 588190 412398 588222 412634
rect 588458 412398 588542 412634
rect 588778 412398 588810 412634
rect 588190 376954 588810 412398
rect 588190 376718 588222 376954
rect 588458 376718 588542 376954
rect 588778 376718 588810 376954
rect 588190 376634 588810 376718
rect 588190 376398 588222 376634
rect 588458 376398 588542 376634
rect 588778 376398 588810 376634
rect 588190 340954 588810 376398
rect 588190 340718 588222 340954
rect 588458 340718 588542 340954
rect 588778 340718 588810 340954
rect 588190 340634 588810 340718
rect 588190 340398 588222 340634
rect 588458 340398 588542 340634
rect 588778 340398 588810 340634
rect 588190 304954 588810 340398
rect 588190 304718 588222 304954
rect 588458 304718 588542 304954
rect 588778 304718 588810 304954
rect 588190 304634 588810 304718
rect 588190 304398 588222 304634
rect 588458 304398 588542 304634
rect 588778 304398 588810 304634
rect 588190 268954 588810 304398
rect 588190 268718 588222 268954
rect 588458 268718 588542 268954
rect 588778 268718 588810 268954
rect 588190 268634 588810 268718
rect 588190 268398 588222 268634
rect 588458 268398 588542 268634
rect 588778 268398 588810 268634
rect 588190 232954 588810 268398
rect 588190 232718 588222 232954
rect 588458 232718 588542 232954
rect 588778 232718 588810 232954
rect 588190 232634 588810 232718
rect 588190 232398 588222 232634
rect 588458 232398 588542 232634
rect 588778 232398 588810 232634
rect 588190 196954 588810 232398
rect 588190 196718 588222 196954
rect 588458 196718 588542 196954
rect 588778 196718 588810 196954
rect 588190 196634 588810 196718
rect 588190 196398 588222 196634
rect 588458 196398 588542 196634
rect 588778 196398 588810 196634
rect 588190 160954 588810 196398
rect 588190 160718 588222 160954
rect 588458 160718 588542 160954
rect 588778 160718 588810 160954
rect 588190 160634 588810 160718
rect 588190 160398 588222 160634
rect 588458 160398 588542 160634
rect 588778 160398 588810 160634
rect 588190 124954 588810 160398
rect 588190 124718 588222 124954
rect 588458 124718 588542 124954
rect 588778 124718 588810 124954
rect 588190 124634 588810 124718
rect 588190 124398 588222 124634
rect 588458 124398 588542 124634
rect 588778 124398 588810 124634
rect 588190 88954 588810 124398
rect 588190 88718 588222 88954
rect 588458 88718 588542 88954
rect 588778 88718 588810 88954
rect 588190 88634 588810 88718
rect 588190 88398 588222 88634
rect 588458 88398 588542 88634
rect 588778 88398 588810 88634
rect 588190 52954 588810 88398
rect 588190 52718 588222 52954
rect 588458 52718 588542 52954
rect 588778 52718 588810 52954
rect 588190 52634 588810 52718
rect 588190 52398 588222 52634
rect 588458 52398 588542 52634
rect 588778 52398 588810 52634
rect 588190 16954 588810 52398
rect 588190 16718 588222 16954
rect 588458 16718 588542 16954
rect 588778 16718 588810 16954
rect 588190 16634 588810 16718
rect 588190 16398 588222 16634
rect 588458 16398 588542 16634
rect 588778 16398 588810 16634
rect 588190 -3226 588810 16398
rect 588190 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect 588190 -3546 588810 -3462
rect 588190 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect 588190 -3814 588810 -3782
rect 589150 669454 589770 708122
rect 589150 669218 589182 669454
rect 589418 669218 589502 669454
rect 589738 669218 589770 669454
rect 589150 669134 589770 669218
rect 589150 668898 589182 669134
rect 589418 668898 589502 669134
rect 589738 668898 589770 669134
rect 589150 633454 589770 668898
rect 589150 633218 589182 633454
rect 589418 633218 589502 633454
rect 589738 633218 589770 633454
rect 589150 633134 589770 633218
rect 589150 632898 589182 633134
rect 589418 632898 589502 633134
rect 589738 632898 589770 633134
rect 589150 597454 589770 632898
rect 589150 597218 589182 597454
rect 589418 597218 589502 597454
rect 589738 597218 589770 597454
rect 589150 597134 589770 597218
rect 589150 596898 589182 597134
rect 589418 596898 589502 597134
rect 589738 596898 589770 597134
rect 589150 561454 589770 596898
rect 589150 561218 589182 561454
rect 589418 561218 589502 561454
rect 589738 561218 589770 561454
rect 589150 561134 589770 561218
rect 589150 560898 589182 561134
rect 589418 560898 589502 561134
rect 589738 560898 589770 561134
rect 589150 525454 589770 560898
rect 589150 525218 589182 525454
rect 589418 525218 589502 525454
rect 589738 525218 589770 525454
rect 589150 525134 589770 525218
rect 589150 524898 589182 525134
rect 589418 524898 589502 525134
rect 589738 524898 589770 525134
rect 589150 489454 589770 524898
rect 589150 489218 589182 489454
rect 589418 489218 589502 489454
rect 589738 489218 589770 489454
rect 589150 489134 589770 489218
rect 589150 488898 589182 489134
rect 589418 488898 589502 489134
rect 589738 488898 589770 489134
rect 589150 453454 589770 488898
rect 589150 453218 589182 453454
rect 589418 453218 589502 453454
rect 589738 453218 589770 453454
rect 589150 453134 589770 453218
rect 589150 452898 589182 453134
rect 589418 452898 589502 453134
rect 589738 452898 589770 453134
rect 589150 417454 589770 452898
rect 589150 417218 589182 417454
rect 589418 417218 589502 417454
rect 589738 417218 589770 417454
rect 589150 417134 589770 417218
rect 589150 416898 589182 417134
rect 589418 416898 589502 417134
rect 589738 416898 589770 417134
rect 589150 381454 589770 416898
rect 589150 381218 589182 381454
rect 589418 381218 589502 381454
rect 589738 381218 589770 381454
rect 589150 381134 589770 381218
rect 589150 380898 589182 381134
rect 589418 380898 589502 381134
rect 589738 380898 589770 381134
rect 589150 345454 589770 380898
rect 589150 345218 589182 345454
rect 589418 345218 589502 345454
rect 589738 345218 589770 345454
rect 589150 345134 589770 345218
rect 589150 344898 589182 345134
rect 589418 344898 589502 345134
rect 589738 344898 589770 345134
rect 589150 309454 589770 344898
rect 589150 309218 589182 309454
rect 589418 309218 589502 309454
rect 589738 309218 589770 309454
rect 589150 309134 589770 309218
rect 589150 308898 589182 309134
rect 589418 308898 589502 309134
rect 589738 308898 589770 309134
rect 589150 273454 589770 308898
rect 589150 273218 589182 273454
rect 589418 273218 589502 273454
rect 589738 273218 589770 273454
rect 589150 273134 589770 273218
rect 589150 272898 589182 273134
rect 589418 272898 589502 273134
rect 589738 272898 589770 273134
rect 589150 237454 589770 272898
rect 589150 237218 589182 237454
rect 589418 237218 589502 237454
rect 589738 237218 589770 237454
rect 589150 237134 589770 237218
rect 589150 236898 589182 237134
rect 589418 236898 589502 237134
rect 589738 236898 589770 237134
rect 589150 201454 589770 236898
rect 589150 201218 589182 201454
rect 589418 201218 589502 201454
rect 589738 201218 589770 201454
rect 589150 201134 589770 201218
rect 589150 200898 589182 201134
rect 589418 200898 589502 201134
rect 589738 200898 589770 201134
rect 589150 165454 589770 200898
rect 589150 165218 589182 165454
rect 589418 165218 589502 165454
rect 589738 165218 589770 165454
rect 589150 165134 589770 165218
rect 589150 164898 589182 165134
rect 589418 164898 589502 165134
rect 589738 164898 589770 165134
rect 589150 129454 589770 164898
rect 589150 129218 589182 129454
rect 589418 129218 589502 129454
rect 589738 129218 589770 129454
rect 589150 129134 589770 129218
rect 589150 128898 589182 129134
rect 589418 128898 589502 129134
rect 589738 128898 589770 129134
rect 589150 93454 589770 128898
rect 589150 93218 589182 93454
rect 589418 93218 589502 93454
rect 589738 93218 589770 93454
rect 589150 93134 589770 93218
rect 589150 92898 589182 93134
rect 589418 92898 589502 93134
rect 589738 92898 589770 93134
rect 589150 57454 589770 92898
rect 589150 57218 589182 57454
rect 589418 57218 589502 57454
rect 589738 57218 589770 57454
rect 589150 57134 589770 57218
rect 589150 56898 589182 57134
rect 589418 56898 589502 57134
rect 589738 56898 589770 57134
rect 589150 21454 589770 56898
rect 589150 21218 589182 21454
rect 589418 21218 589502 21454
rect 589738 21218 589770 21454
rect 589150 21134 589770 21218
rect 589150 20898 589182 21134
rect 589418 20898 589502 21134
rect 589738 20898 589770 21134
rect 589150 -4186 589770 20898
rect 589150 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect 589150 -4506 589770 -4422
rect 589150 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect 589150 -4774 589770 -4742
rect 590110 673954 590730 709082
rect 590110 673718 590142 673954
rect 590378 673718 590462 673954
rect 590698 673718 590730 673954
rect 590110 673634 590730 673718
rect 590110 673398 590142 673634
rect 590378 673398 590462 673634
rect 590698 673398 590730 673634
rect 590110 637954 590730 673398
rect 590110 637718 590142 637954
rect 590378 637718 590462 637954
rect 590698 637718 590730 637954
rect 590110 637634 590730 637718
rect 590110 637398 590142 637634
rect 590378 637398 590462 637634
rect 590698 637398 590730 637634
rect 590110 601954 590730 637398
rect 590110 601718 590142 601954
rect 590378 601718 590462 601954
rect 590698 601718 590730 601954
rect 590110 601634 590730 601718
rect 590110 601398 590142 601634
rect 590378 601398 590462 601634
rect 590698 601398 590730 601634
rect 590110 565954 590730 601398
rect 590110 565718 590142 565954
rect 590378 565718 590462 565954
rect 590698 565718 590730 565954
rect 590110 565634 590730 565718
rect 590110 565398 590142 565634
rect 590378 565398 590462 565634
rect 590698 565398 590730 565634
rect 590110 529954 590730 565398
rect 590110 529718 590142 529954
rect 590378 529718 590462 529954
rect 590698 529718 590730 529954
rect 590110 529634 590730 529718
rect 590110 529398 590142 529634
rect 590378 529398 590462 529634
rect 590698 529398 590730 529634
rect 590110 493954 590730 529398
rect 590110 493718 590142 493954
rect 590378 493718 590462 493954
rect 590698 493718 590730 493954
rect 590110 493634 590730 493718
rect 590110 493398 590142 493634
rect 590378 493398 590462 493634
rect 590698 493398 590730 493634
rect 590110 457954 590730 493398
rect 590110 457718 590142 457954
rect 590378 457718 590462 457954
rect 590698 457718 590730 457954
rect 590110 457634 590730 457718
rect 590110 457398 590142 457634
rect 590378 457398 590462 457634
rect 590698 457398 590730 457634
rect 590110 421954 590730 457398
rect 590110 421718 590142 421954
rect 590378 421718 590462 421954
rect 590698 421718 590730 421954
rect 590110 421634 590730 421718
rect 590110 421398 590142 421634
rect 590378 421398 590462 421634
rect 590698 421398 590730 421634
rect 590110 385954 590730 421398
rect 590110 385718 590142 385954
rect 590378 385718 590462 385954
rect 590698 385718 590730 385954
rect 590110 385634 590730 385718
rect 590110 385398 590142 385634
rect 590378 385398 590462 385634
rect 590698 385398 590730 385634
rect 590110 349954 590730 385398
rect 590110 349718 590142 349954
rect 590378 349718 590462 349954
rect 590698 349718 590730 349954
rect 590110 349634 590730 349718
rect 590110 349398 590142 349634
rect 590378 349398 590462 349634
rect 590698 349398 590730 349634
rect 590110 313954 590730 349398
rect 590110 313718 590142 313954
rect 590378 313718 590462 313954
rect 590698 313718 590730 313954
rect 590110 313634 590730 313718
rect 590110 313398 590142 313634
rect 590378 313398 590462 313634
rect 590698 313398 590730 313634
rect 590110 277954 590730 313398
rect 590110 277718 590142 277954
rect 590378 277718 590462 277954
rect 590698 277718 590730 277954
rect 590110 277634 590730 277718
rect 590110 277398 590142 277634
rect 590378 277398 590462 277634
rect 590698 277398 590730 277634
rect 590110 241954 590730 277398
rect 590110 241718 590142 241954
rect 590378 241718 590462 241954
rect 590698 241718 590730 241954
rect 590110 241634 590730 241718
rect 590110 241398 590142 241634
rect 590378 241398 590462 241634
rect 590698 241398 590730 241634
rect 590110 205954 590730 241398
rect 590110 205718 590142 205954
rect 590378 205718 590462 205954
rect 590698 205718 590730 205954
rect 590110 205634 590730 205718
rect 590110 205398 590142 205634
rect 590378 205398 590462 205634
rect 590698 205398 590730 205634
rect 590110 169954 590730 205398
rect 590110 169718 590142 169954
rect 590378 169718 590462 169954
rect 590698 169718 590730 169954
rect 590110 169634 590730 169718
rect 590110 169398 590142 169634
rect 590378 169398 590462 169634
rect 590698 169398 590730 169634
rect 590110 133954 590730 169398
rect 590110 133718 590142 133954
rect 590378 133718 590462 133954
rect 590698 133718 590730 133954
rect 590110 133634 590730 133718
rect 590110 133398 590142 133634
rect 590378 133398 590462 133634
rect 590698 133398 590730 133634
rect 590110 97954 590730 133398
rect 590110 97718 590142 97954
rect 590378 97718 590462 97954
rect 590698 97718 590730 97954
rect 590110 97634 590730 97718
rect 590110 97398 590142 97634
rect 590378 97398 590462 97634
rect 590698 97398 590730 97634
rect 590110 61954 590730 97398
rect 590110 61718 590142 61954
rect 590378 61718 590462 61954
rect 590698 61718 590730 61954
rect 590110 61634 590730 61718
rect 590110 61398 590142 61634
rect 590378 61398 590462 61634
rect 590698 61398 590730 61634
rect 590110 25954 590730 61398
rect 590110 25718 590142 25954
rect 590378 25718 590462 25954
rect 590698 25718 590730 25954
rect 590110 25634 590730 25718
rect 590110 25398 590142 25634
rect 590378 25398 590462 25634
rect 590698 25398 590730 25634
rect 590110 -5146 590730 25398
rect 590110 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect 590110 -5466 590730 -5382
rect 590110 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect 590110 -5734 590730 -5702
rect 591070 678454 591690 710042
rect 591070 678218 591102 678454
rect 591338 678218 591422 678454
rect 591658 678218 591690 678454
rect 591070 678134 591690 678218
rect 591070 677898 591102 678134
rect 591338 677898 591422 678134
rect 591658 677898 591690 678134
rect 591070 642454 591690 677898
rect 591070 642218 591102 642454
rect 591338 642218 591422 642454
rect 591658 642218 591690 642454
rect 591070 642134 591690 642218
rect 591070 641898 591102 642134
rect 591338 641898 591422 642134
rect 591658 641898 591690 642134
rect 591070 606454 591690 641898
rect 591070 606218 591102 606454
rect 591338 606218 591422 606454
rect 591658 606218 591690 606454
rect 591070 606134 591690 606218
rect 591070 605898 591102 606134
rect 591338 605898 591422 606134
rect 591658 605898 591690 606134
rect 591070 570454 591690 605898
rect 591070 570218 591102 570454
rect 591338 570218 591422 570454
rect 591658 570218 591690 570454
rect 591070 570134 591690 570218
rect 591070 569898 591102 570134
rect 591338 569898 591422 570134
rect 591658 569898 591690 570134
rect 591070 534454 591690 569898
rect 591070 534218 591102 534454
rect 591338 534218 591422 534454
rect 591658 534218 591690 534454
rect 591070 534134 591690 534218
rect 591070 533898 591102 534134
rect 591338 533898 591422 534134
rect 591658 533898 591690 534134
rect 591070 498454 591690 533898
rect 591070 498218 591102 498454
rect 591338 498218 591422 498454
rect 591658 498218 591690 498454
rect 591070 498134 591690 498218
rect 591070 497898 591102 498134
rect 591338 497898 591422 498134
rect 591658 497898 591690 498134
rect 591070 462454 591690 497898
rect 591070 462218 591102 462454
rect 591338 462218 591422 462454
rect 591658 462218 591690 462454
rect 591070 462134 591690 462218
rect 591070 461898 591102 462134
rect 591338 461898 591422 462134
rect 591658 461898 591690 462134
rect 591070 426454 591690 461898
rect 591070 426218 591102 426454
rect 591338 426218 591422 426454
rect 591658 426218 591690 426454
rect 591070 426134 591690 426218
rect 591070 425898 591102 426134
rect 591338 425898 591422 426134
rect 591658 425898 591690 426134
rect 591070 390454 591690 425898
rect 591070 390218 591102 390454
rect 591338 390218 591422 390454
rect 591658 390218 591690 390454
rect 591070 390134 591690 390218
rect 591070 389898 591102 390134
rect 591338 389898 591422 390134
rect 591658 389898 591690 390134
rect 591070 354454 591690 389898
rect 591070 354218 591102 354454
rect 591338 354218 591422 354454
rect 591658 354218 591690 354454
rect 591070 354134 591690 354218
rect 591070 353898 591102 354134
rect 591338 353898 591422 354134
rect 591658 353898 591690 354134
rect 591070 318454 591690 353898
rect 591070 318218 591102 318454
rect 591338 318218 591422 318454
rect 591658 318218 591690 318454
rect 591070 318134 591690 318218
rect 591070 317898 591102 318134
rect 591338 317898 591422 318134
rect 591658 317898 591690 318134
rect 591070 282454 591690 317898
rect 591070 282218 591102 282454
rect 591338 282218 591422 282454
rect 591658 282218 591690 282454
rect 591070 282134 591690 282218
rect 591070 281898 591102 282134
rect 591338 281898 591422 282134
rect 591658 281898 591690 282134
rect 591070 246454 591690 281898
rect 591070 246218 591102 246454
rect 591338 246218 591422 246454
rect 591658 246218 591690 246454
rect 591070 246134 591690 246218
rect 591070 245898 591102 246134
rect 591338 245898 591422 246134
rect 591658 245898 591690 246134
rect 591070 210454 591690 245898
rect 591070 210218 591102 210454
rect 591338 210218 591422 210454
rect 591658 210218 591690 210454
rect 591070 210134 591690 210218
rect 591070 209898 591102 210134
rect 591338 209898 591422 210134
rect 591658 209898 591690 210134
rect 591070 174454 591690 209898
rect 591070 174218 591102 174454
rect 591338 174218 591422 174454
rect 591658 174218 591690 174454
rect 591070 174134 591690 174218
rect 591070 173898 591102 174134
rect 591338 173898 591422 174134
rect 591658 173898 591690 174134
rect 591070 138454 591690 173898
rect 591070 138218 591102 138454
rect 591338 138218 591422 138454
rect 591658 138218 591690 138454
rect 591070 138134 591690 138218
rect 591070 137898 591102 138134
rect 591338 137898 591422 138134
rect 591658 137898 591690 138134
rect 591070 102454 591690 137898
rect 591070 102218 591102 102454
rect 591338 102218 591422 102454
rect 591658 102218 591690 102454
rect 591070 102134 591690 102218
rect 591070 101898 591102 102134
rect 591338 101898 591422 102134
rect 591658 101898 591690 102134
rect 591070 66454 591690 101898
rect 591070 66218 591102 66454
rect 591338 66218 591422 66454
rect 591658 66218 591690 66454
rect 591070 66134 591690 66218
rect 591070 65898 591102 66134
rect 591338 65898 591422 66134
rect 591658 65898 591690 66134
rect 591070 30454 591690 65898
rect 591070 30218 591102 30454
rect 591338 30218 591422 30454
rect 591658 30218 591690 30454
rect 591070 30134 591690 30218
rect 591070 29898 591102 30134
rect 591338 29898 591422 30134
rect 591658 29898 591690 30134
rect 591070 -6106 591690 29898
rect 591070 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect 591070 -6426 591690 -6342
rect 591070 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect 591070 -6694 591690 -6662
rect 592030 682954 592650 711002
rect 592030 682718 592062 682954
rect 592298 682718 592382 682954
rect 592618 682718 592650 682954
rect 592030 682634 592650 682718
rect 592030 682398 592062 682634
rect 592298 682398 592382 682634
rect 592618 682398 592650 682634
rect 592030 646954 592650 682398
rect 592030 646718 592062 646954
rect 592298 646718 592382 646954
rect 592618 646718 592650 646954
rect 592030 646634 592650 646718
rect 592030 646398 592062 646634
rect 592298 646398 592382 646634
rect 592618 646398 592650 646634
rect 592030 610954 592650 646398
rect 592030 610718 592062 610954
rect 592298 610718 592382 610954
rect 592618 610718 592650 610954
rect 592030 610634 592650 610718
rect 592030 610398 592062 610634
rect 592298 610398 592382 610634
rect 592618 610398 592650 610634
rect 592030 574954 592650 610398
rect 592030 574718 592062 574954
rect 592298 574718 592382 574954
rect 592618 574718 592650 574954
rect 592030 574634 592650 574718
rect 592030 574398 592062 574634
rect 592298 574398 592382 574634
rect 592618 574398 592650 574634
rect 592030 538954 592650 574398
rect 592030 538718 592062 538954
rect 592298 538718 592382 538954
rect 592618 538718 592650 538954
rect 592030 538634 592650 538718
rect 592030 538398 592062 538634
rect 592298 538398 592382 538634
rect 592618 538398 592650 538634
rect 592030 502954 592650 538398
rect 592030 502718 592062 502954
rect 592298 502718 592382 502954
rect 592618 502718 592650 502954
rect 592030 502634 592650 502718
rect 592030 502398 592062 502634
rect 592298 502398 592382 502634
rect 592618 502398 592650 502634
rect 592030 466954 592650 502398
rect 592030 466718 592062 466954
rect 592298 466718 592382 466954
rect 592618 466718 592650 466954
rect 592030 466634 592650 466718
rect 592030 466398 592062 466634
rect 592298 466398 592382 466634
rect 592618 466398 592650 466634
rect 592030 430954 592650 466398
rect 592030 430718 592062 430954
rect 592298 430718 592382 430954
rect 592618 430718 592650 430954
rect 592030 430634 592650 430718
rect 592030 430398 592062 430634
rect 592298 430398 592382 430634
rect 592618 430398 592650 430634
rect 592030 394954 592650 430398
rect 592030 394718 592062 394954
rect 592298 394718 592382 394954
rect 592618 394718 592650 394954
rect 592030 394634 592650 394718
rect 592030 394398 592062 394634
rect 592298 394398 592382 394634
rect 592618 394398 592650 394634
rect 592030 358954 592650 394398
rect 592030 358718 592062 358954
rect 592298 358718 592382 358954
rect 592618 358718 592650 358954
rect 592030 358634 592650 358718
rect 592030 358398 592062 358634
rect 592298 358398 592382 358634
rect 592618 358398 592650 358634
rect 592030 322954 592650 358398
rect 592030 322718 592062 322954
rect 592298 322718 592382 322954
rect 592618 322718 592650 322954
rect 592030 322634 592650 322718
rect 592030 322398 592062 322634
rect 592298 322398 592382 322634
rect 592618 322398 592650 322634
rect 592030 286954 592650 322398
rect 592030 286718 592062 286954
rect 592298 286718 592382 286954
rect 592618 286718 592650 286954
rect 592030 286634 592650 286718
rect 592030 286398 592062 286634
rect 592298 286398 592382 286634
rect 592618 286398 592650 286634
rect 592030 250954 592650 286398
rect 592030 250718 592062 250954
rect 592298 250718 592382 250954
rect 592618 250718 592650 250954
rect 592030 250634 592650 250718
rect 592030 250398 592062 250634
rect 592298 250398 592382 250634
rect 592618 250398 592650 250634
rect 592030 214954 592650 250398
rect 592030 214718 592062 214954
rect 592298 214718 592382 214954
rect 592618 214718 592650 214954
rect 592030 214634 592650 214718
rect 592030 214398 592062 214634
rect 592298 214398 592382 214634
rect 592618 214398 592650 214634
rect 592030 178954 592650 214398
rect 592030 178718 592062 178954
rect 592298 178718 592382 178954
rect 592618 178718 592650 178954
rect 592030 178634 592650 178718
rect 592030 178398 592062 178634
rect 592298 178398 592382 178634
rect 592618 178398 592650 178634
rect 592030 142954 592650 178398
rect 592030 142718 592062 142954
rect 592298 142718 592382 142954
rect 592618 142718 592650 142954
rect 592030 142634 592650 142718
rect 592030 142398 592062 142634
rect 592298 142398 592382 142634
rect 592618 142398 592650 142634
rect 592030 106954 592650 142398
rect 592030 106718 592062 106954
rect 592298 106718 592382 106954
rect 592618 106718 592650 106954
rect 592030 106634 592650 106718
rect 592030 106398 592062 106634
rect 592298 106398 592382 106634
rect 592618 106398 592650 106634
rect 592030 70954 592650 106398
rect 592030 70718 592062 70954
rect 592298 70718 592382 70954
rect 592618 70718 592650 70954
rect 592030 70634 592650 70718
rect 592030 70398 592062 70634
rect 592298 70398 592382 70634
rect 592618 70398 592650 70634
rect 592030 34954 592650 70398
rect 592030 34718 592062 34954
rect 592298 34718 592382 34954
rect 592618 34718 592650 34954
rect 592030 34634 592650 34718
rect 592030 34398 592062 34634
rect 592298 34398 592382 34634
rect 592618 34398 592650 34634
rect 592030 -7066 592650 34398
rect 592030 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect 592030 -7386 592650 -7302
rect 592030 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect 592030 -7654 592650 -7622
<< via4 >>
rect -8694 711322 -8458 711558
rect -8374 711322 -8138 711558
rect -8694 711002 -8458 711238
rect -8374 711002 -8138 711238
rect -8694 682718 -8458 682954
rect -8374 682718 -8138 682954
rect -8694 682398 -8458 682634
rect -8374 682398 -8138 682634
rect -8694 646718 -8458 646954
rect -8374 646718 -8138 646954
rect -8694 646398 -8458 646634
rect -8374 646398 -8138 646634
rect -8694 610718 -8458 610954
rect -8374 610718 -8138 610954
rect -8694 610398 -8458 610634
rect -8374 610398 -8138 610634
rect -8694 574718 -8458 574954
rect -8374 574718 -8138 574954
rect -8694 574398 -8458 574634
rect -8374 574398 -8138 574634
rect -8694 538718 -8458 538954
rect -8374 538718 -8138 538954
rect -8694 538398 -8458 538634
rect -8374 538398 -8138 538634
rect -8694 502718 -8458 502954
rect -8374 502718 -8138 502954
rect -8694 502398 -8458 502634
rect -8374 502398 -8138 502634
rect -8694 466718 -8458 466954
rect -8374 466718 -8138 466954
rect -8694 466398 -8458 466634
rect -8374 466398 -8138 466634
rect -8694 430718 -8458 430954
rect -8374 430718 -8138 430954
rect -8694 430398 -8458 430634
rect -8374 430398 -8138 430634
rect -8694 394718 -8458 394954
rect -8374 394718 -8138 394954
rect -8694 394398 -8458 394634
rect -8374 394398 -8138 394634
rect -8694 358718 -8458 358954
rect -8374 358718 -8138 358954
rect -8694 358398 -8458 358634
rect -8374 358398 -8138 358634
rect -8694 322718 -8458 322954
rect -8374 322718 -8138 322954
rect -8694 322398 -8458 322634
rect -8374 322398 -8138 322634
rect -8694 286718 -8458 286954
rect -8374 286718 -8138 286954
rect -8694 286398 -8458 286634
rect -8374 286398 -8138 286634
rect -8694 250718 -8458 250954
rect -8374 250718 -8138 250954
rect -8694 250398 -8458 250634
rect -8374 250398 -8138 250634
rect -8694 214718 -8458 214954
rect -8374 214718 -8138 214954
rect -8694 214398 -8458 214634
rect -8374 214398 -8138 214634
rect -8694 178718 -8458 178954
rect -8374 178718 -8138 178954
rect -8694 178398 -8458 178634
rect -8374 178398 -8138 178634
rect -8694 142718 -8458 142954
rect -8374 142718 -8138 142954
rect -8694 142398 -8458 142634
rect -8374 142398 -8138 142634
rect -8694 106718 -8458 106954
rect -8374 106718 -8138 106954
rect -8694 106398 -8458 106634
rect -8374 106398 -8138 106634
rect -8694 70718 -8458 70954
rect -8374 70718 -8138 70954
rect -8694 70398 -8458 70634
rect -8374 70398 -8138 70634
rect -8694 34718 -8458 34954
rect -8374 34718 -8138 34954
rect -8694 34398 -8458 34634
rect -8374 34398 -8138 34634
rect -7734 710362 -7498 710598
rect -7414 710362 -7178 710598
rect -7734 710042 -7498 710278
rect -7414 710042 -7178 710278
rect -7734 678218 -7498 678454
rect -7414 678218 -7178 678454
rect -7734 677898 -7498 678134
rect -7414 677898 -7178 678134
rect -7734 642218 -7498 642454
rect -7414 642218 -7178 642454
rect -7734 641898 -7498 642134
rect -7414 641898 -7178 642134
rect -7734 606218 -7498 606454
rect -7414 606218 -7178 606454
rect -7734 605898 -7498 606134
rect -7414 605898 -7178 606134
rect -7734 570218 -7498 570454
rect -7414 570218 -7178 570454
rect -7734 569898 -7498 570134
rect -7414 569898 -7178 570134
rect -7734 534218 -7498 534454
rect -7414 534218 -7178 534454
rect -7734 533898 -7498 534134
rect -7414 533898 -7178 534134
rect -7734 498218 -7498 498454
rect -7414 498218 -7178 498454
rect -7734 497898 -7498 498134
rect -7414 497898 -7178 498134
rect -7734 462218 -7498 462454
rect -7414 462218 -7178 462454
rect -7734 461898 -7498 462134
rect -7414 461898 -7178 462134
rect -7734 426218 -7498 426454
rect -7414 426218 -7178 426454
rect -7734 425898 -7498 426134
rect -7414 425898 -7178 426134
rect -7734 390218 -7498 390454
rect -7414 390218 -7178 390454
rect -7734 389898 -7498 390134
rect -7414 389898 -7178 390134
rect -7734 354218 -7498 354454
rect -7414 354218 -7178 354454
rect -7734 353898 -7498 354134
rect -7414 353898 -7178 354134
rect -7734 318218 -7498 318454
rect -7414 318218 -7178 318454
rect -7734 317898 -7498 318134
rect -7414 317898 -7178 318134
rect -7734 282218 -7498 282454
rect -7414 282218 -7178 282454
rect -7734 281898 -7498 282134
rect -7414 281898 -7178 282134
rect -7734 246218 -7498 246454
rect -7414 246218 -7178 246454
rect -7734 245898 -7498 246134
rect -7414 245898 -7178 246134
rect -7734 210218 -7498 210454
rect -7414 210218 -7178 210454
rect -7734 209898 -7498 210134
rect -7414 209898 -7178 210134
rect -7734 174218 -7498 174454
rect -7414 174218 -7178 174454
rect -7734 173898 -7498 174134
rect -7414 173898 -7178 174134
rect -7734 138218 -7498 138454
rect -7414 138218 -7178 138454
rect -7734 137898 -7498 138134
rect -7414 137898 -7178 138134
rect -7734 102218 -7498 102454
rect -7414 102218 -7178 102454
rect -7734 101898 -7498 102134
rect -7414 101898 -7178 102134
rect -7734 66218 -7498 66454
rect -7414 66218 -7178 66454
rect -7734 65898 -7498 66134
rect -7414 65898 -7178 66134
rect -7734 30218 -7498 30454
rect -7414 30218 -7178 30454
rect -7734 29898 -7498 30134
rect -7414 29898 -7178 30134
rect -6774 709402 -6538 709638
rect -6454 709402 -6218 709638
rect -6774 709082 -6538 709318
rect -6454 709082 -6218 709318
rect -6774 673718 -6538 673954
rect -6454 673718 -6218 673954
rect -6774 673398 -6538 673634
rect -6454 673398 -6218 673634
rect -6774 637718 -6538 637954
rect -6454 637718 -6218 637954
rect -6774 637398 -6538 637634
rect -6454 637398 -6218 637634
rect -6774 601718 -6538 601954
rect -6454 601718 -6218 601954
rect -6774 601398 -6538 601634
rect -6454 601398 -6218 601634
rect -6774 565718 -6538 565954
rect -6454 565718 -6218 565954
rect -6774 565398 -6538 565634
rect -6454 565398 -6218 565634
rect -6774 529718 -6538 529954
rect -6454 529718 -6218 529954
rect -6774 529398 -6538 529634
rect -6454 529398 -6218 529634
rect -6774 493718 -6538 493954
rect -6454 493718 -6218 493954
rect -6774 493398 -6538 493634
rect -6454 493398 -6218 493634
rect -6774 457718 -6538 457954
rect -6454 457718 -6218 457954
rect -6774 457398 -6538 457634
rect -6454 457398 -6218 457634
rect -6774 421718 -6538 421954
rect -6454 421718 -6218 421954
rect -6774 421398 -6538 421634
rect -6454 421398 -6218 421634
rect -6774 385718 -6538 385954
rect -6454 385718 -6218 385954
rect -6774 385398 -6538 385634
rect -6454 385398 -6218 385634
rect -6774 349718 -6538 349954
rect -6454 349718 -6218 349954
rect -6774 349398 -6538 349634
rect -6454 349398 -6218 349634
rect -6774 313718 -6538 313954
rect -6454 313718 -6218 313954
rect -6774 313398 -6538 313634
rect -6454 313398 -6218 313634
rect -6774 277718 -6538 277954
rect -6454 277718 -6218 277954
rect -6774 277398 -6538 277634
rect -6454 277398 -6218 277634
rect -6774 241718 -6538 241954
rect -6454 241718 -6218 241954
rect -6774 241398 -6538 241634
rect -6454 241398 -6218 241634
rect -6774 205718 -6538 205954
rect -6454 205718 -6218 205954
rect -6774 205398 -6538 205634
rect -6454 205398 -6218 205634
rect -6774 169718 -6538 169954
rect -6454 169718 -6218 169954
rect -6774 169398 -6538 169634
rect -6454 169398 -6218 169634
rect -6774 133718 -6538 133954
rect -6454 133718 -6218 133954
rect -6774 133398 -6538 133634
rect -6454 133398 -6218 133634
rect -6774 97718 -6538 97954
rect -6454 97718 -6218 97954
rect -6774 97398 -6538 97634
rect -6454 97398 -6218 97634
rect -6774 61718 -6538 61954
rect -6454 61718 -6218 61954
rect -6774 61398 -6538 61634
rect -6454 61398 -6218 61634
rect -6774 25718 -6538 25954
rect -6454 25718 -6218 25954
rect -6774 25398 -6538 25634
rect -6454 25398 -6218 25634
rect -5814 708442 -5578 708678
rect -5494 708442 -5258 708678
rect -5814 708122 -5578 708358
rect -5494 708122 -5258 708358
rect -5814 669218 -5578 669454
rect -5494 669218 -5258 669454
rect -5814 668898 -5578 669134
rect -5494 668898 -5258 669134
rect -5814 633218 -5578 633454
rect -5494 633218 -5258 633454
rect -5814 632898 -5578 633134
rect -5494 632898 -5258 633134
rect -5814 597218 -5578 597454
rect -5494 597218 -5258 597454
rect -5814 596898 -5578 597134
rect -5494 596898 -5258 597134
rect -5814 561218 -5578 561454
rect -5494 561218 -5258 561454
rect -5814 560898 -5578 561134
rect -5494 560898 -5258 561134
rect -5814 525218 -5578 525454
rect -5494 525218 -5258 525454
rect -5814 524898 -5578 525134
rect -5494 524898 -5258 525134
rect -5814 489218 -5578 489454
rect -5494 489218 -5258 489454
rect -5814 488898 -5578 489134
rect -5494 488898 -5258 489134
rect -5814 453218 -5578 453454
rect -5494 453218 -5258 453454
rect -5814 452898 -5578 453134
rect -5494 452898 -5258 453134
rect -5814 417218 -5578 417454
rect -5494 417218 -5258 417454
rect -5814 416898 -5578 417134
rect -5494 416898 -5258 417134
rect -5814 381218 -5578 381454
rect -5494 381218 -5258 381454
rect -5814 380898 -5578 381134
rect -5494 380898 -5258 381134
rect -5814 345218 -5578 345454
rect -5494 345218 -5258 345454
rect -5814 344898 -5578 345134
rect -5494 344898 -5258 345134
rect -5814 309218 -5578 309454
rect -5494 309218 -5258 309454
rect -5814 308898 -5578 309134
rect -5494 308898 -5258 309134
rect -5814 273218 -5578 273454
rect -5494 273218 -5258 273454
rect -5814 272898 -5578 273134
rect -5494 272898 -5258 273134
rect -5814 237218 -5578 237454
rect -5494 237218 -5258 237454
rect -5814 236898 -5578 237134
rect -5494 236898 -5258 237134
rect -5814 201218 -5578 201454
rect -5494 201218 -5258 201454
rect -5814 200898 -5578 201134
rect -5494 200898 -5258 201134
rect -5814 165218 -5578 165454
rect -5494 165218 -5258 165454
rect -5814 164898 -5578 165134
rect -5494 164898 -5258 165134
rect -5814 129218 -5578 129454
rect -5494 129218 -5258 129454
rect -5814 128898 -5578 129134
rect -5494 128898 -5258 129134
rect -5814 93218 -5578 93454
rect -5494 93218 -5258 93454
rect -5814 92898 -5578 93134
rect -5494 92898 -5258 93134
rect -5814 57218 -5578 57454
rect -5494 57218 -5258 57454
rect -5814 56898 -5578 57134
rect -5494 56898 -5258 57134
rect -5814 21218 -5578 21454
rect -5494 21218 -5258 21454
rect -5814 20898 -5578 21134
rect -5494 20898 -5258 21134
rect -4854 707482 -4618 707718
rect -4534 707482 -4298 707718
rect -4854 707162 -4618 707398
rect -4534 707162 -4298 707398
rect -4854 700718 -4618 700954
rect -4534 700718 -4298 700954
rect -4854 700398 -4618 700634
rect -4534 700398 -4298 700634
rect -4854 664718 -4618 664954
rect -4534 664718 -4298 664954
rect -4854 664398 -4618 664634
rect -4534 664398 -4298 664634
rect -4854 628718 -4618 628954
rect -4534 628718 -4298 628954
rect -4854 628398 -4618 628634
rect -4534 628398 -4298 628634
rect -4854 592718 -4618 592954
rect -4534 592718 -4298 592954
rect -4854 592398 -4618 592634
rect -4534 592398 -4298 592634
rect -4854 556718 -4618 556954
rect -4534 556718 -4298 556954
rect -4854 556398 -4618 556634
rect -4534 556398 -4298 556634
rect -4854 520718 -4618 520954
rect -4534 520718 -4298 520954
rect -4854 520398 -4618 520634
rect -4534 520398 -4298 520634
rect -4854 484718 -4618 484954
rect -4534 484718 -4298 484954
rect -4854 484398 -4618 484634
rect -4534 484398 -4298 484634
rect -4854 448718 -4618 448954
rect -4534 448718 -4298 448954
rect -4854 448398 -4618 448634
rect -4534 448398 -4298 448634
rect -4854 412718 -4618 412954
rect -4534 412718 -4298 412954
rect -4854 412398 -4618 412634
rect -4534 412398 -4298 412634
rect -4854 376718 -4618 376954
rect -4534 376718 -4298 376954
rect -4854 376398 -4618 376634
rect -4534 376398 -4298 376634
rect -4854 340718 -4618 340954
rect -4534 340718 -4298 340954
rect -4854 340398 -4618 340634
rect -4534 340398 -4298 340634
rect -4854 304718 -4618 304954
rect -4534 304718 -4298 304954
rect -4854 304398 -4618 304634
rect -4534 304398 -4298 304634
rect -4854 268718 -4618 268954
rect -4534 268718 -4298 268954
rect -4854 268398 -4618 268634
rect -4534 268398 -4298 268634
rect -4854 232718 -4618 232954
rect -4534 232718 -4298 232954
rect -4854 232398 -4618 232634
rect -4534 232398 -4298 232634
rect -4854 196718 -4618 196954
rect -4534 196718 -4298 196954
rect -4854 196398 -4618 196634
rect -4534 196398 -4298 196634
rect -4854 160718 -4618 160954
rect -4534 160718 -4298 160954
rect -4854 160398 -4618 160634
rect -4534 160398 -4298 160634
rect -4854 124718 -4618 124954
rect -4534 124718 -4298 124954
rect -4854 124398 -4618 124634
rect -4534 124398 -4298 124634
rect -4854 88718 -4618 88954
rect -4534 88718 -4298 88954
rect -4854 88398 -4618 88634
rect -4534 88398 -4298 88634
rect -4854 52718 -4618 52954
rect -4534 52718 -4298 52954
rect -4854 52398 -4618 52634
rect -4534 52398 -4298 52634
rect -4854 16718 -4618 16954
rect -4534 16718 -4298 16954
rect -4854 16398 -4618 16634
rect -4534 16398 -4298 16634
rect -3894 706522 -3658 706758
rect -3574 706522 -3338 706758
rect -3894 706202 -3658 706438
rect -3574 706202 -3338 706438
rect -3894 696218 -3658 696454
rect -3574 696218 -3338 696454
rect -3894 695898 -3658 696134
rect -3574 695898 -3338 696134
rect -3894 660218 -3658 660454
rect -3574 660218 -3338 660454
rect -3894 659898 -3658 660134
rect -3574 659898 -3338 660134
rect -3894 624218 -3658 624454
rect -3574 624218 -3338 624454
rect -3894 623898 -3658 624134
rect -3574 623898 -3338 624134
rect -3894 588218 -3658 588454
rect -3574 588218 -3338 588454
rect -3894 587898 -3658 588134
rect -3574 587898 -3338 588134
rect -3894 552218 -3658 552454
rect -3574 552218 -3338 552454
rect -3894 551898 -3658 552134
rect -3574 551898 -3338 552134
rect -3894 516218 -3658 516454
rect -3574 516218 -3338 516454
rect -3894 515898 -3658 516134
rect -3574 515898 -3338 516134
rect -3894 480218 -3658 480454
rect -3574 480218 -3338 480454
rect -3894 479898 -3658 480134
rect -3574 479898 -3338 480134
rect -3894 444218 -3658 444454
rect -3574 444218 -3338 444454
rect -3894 443898 -3658 444134
rect -3574 443898 -3338 444134
rect -3894 408218 -3658 408454
rect -3574 408218 -3338 408454
rect -3894 407898 -3658 408134
rect -3574 407898 -3338 408134
rect -3894 372218 -3658 372454
rect -3574 372218 -3338 372454
rect -3894 371898 -3658 372134
rect -3574 371898 -3338 372134
rect -3894 336218 -3658 336454
rect -3574 336218 -3338 336454
rect -3894 335898 -3658 336134
rect -3574 335898 -3338 336134
rect -3894 300218 -3658 300454
rect -3574 300218 -3338 300454
rect -3894 299898 -3658 300134
rect -3574 299898 -3338 300134
rect -3894 264218 -3658 264454
rect -3574 264218 -3338 264454
rect -3894 263898 -3658 264134
rect -3574 263898 -3338 264134
rect -3894 228218 -3658 228454
rect -3574 228218 -3338 228454
rect -3894 227898 -3658 228134
rect -3574 227898 -3338 228134
rect -3894 192218 -3658 192454
rect -3574 192218 -3338 192454
rect -3894 191898 -3658 192134
rect -3574 191898 -3338 192134
rect -3894 156218 -3658 156454
rect -3574 156218 -3338 156454
rect -3894 155898 -3658 156134
rect -3574 155898 -3338 156134
rect -3894 120218 -3658 120454
rect -3574 120218 -3338 120454
rect -3894 119898 -3658 120134
rect -3574 119898 -3338 120134
rect -3894 84218 -3658 84454
rect -3574 84218 -3338 84454
rect -3894 83898 -3658 84134
rect -3574 83898 -3338 84134
rect -3894 48218 -3658 48454
rect -3574 48218 -3338 48454
rect -3894 47898 -3658 48134
rect -3574 47898 -3338 48134
rect -3894 12218 -3658 12454
rect -3574 12218 -3338 12454
rect -3894 11898 -3658 12134
rect -3574 11898 -3338 12134
rect -2934 705562 -2698 705798
rect -2614 705562 -2378 705798
rect -2934 705242 -2698 705478
rect -2614 705242 -2378 705478
rect -2934 691718 -2698 691954
rect -2614 691718 -2378 691954
rect -2934 691398 -2698 691634
rect -2614 691398 -2378 691634
rect -2934 655718 -2698 655954
rect -2614 655718 -2378 655954
rect -2934 655398 -2698 655634
rect -2614 655398 -2378 655634
rect -2934 619718 -2698 619954
rect -2614 619718 -2378 619954
rect -2934 619398 -2698 619634
rect -2614 619398 -2378 619634
rect -2934 583718 -2698 583954
rect -2614 583718 -2378 583954
rect -2934 583398 -2698 583634
rect -2614 583398 -2378 583634
rect -2934 547718 -2698 547954
rect -2614 547718 -2378 547954
rect -2934 547398 -2698 547634
rect -2614 547398 -2378 547634
rect -2934 511718 -2698 511954
rect -2614 511718 -2378 511954
rect -2934 511398 -2698 511634
rect -2614 511398 -2378 511634
rect -2934 475718 -2698 475954
rect -2614 475718 -2378 475954
rect -2934 475398 -2698 475634
rect -2614 475398 -2378 475634
rect -2934 439718 -2698 439954
rect -2614 439718 -2378 439954
rect -2934 439398 -2698 439634
rect -2614 439398 -2378 439634
rect -2934 403718 -2698 403954
rect -2614 403718 -2378 403954
rect -2934 403398 -2698 403634
rect -2614 403398 -2378 403634
rect -2934 367718 -2698 367954
rect -2614 367718 -2378 367954
rect -2934 367398 -2698 367634
rect -2614 367398 -2378 367634
rect -2934 331718 -2698 331954
rect -2614 331718 -2378 331954
rect -2934 331398 -2698 331634
rect -2614 331398 -2378 331634
rect -2934 295718 -2698 295954
rect -2614 295718 -2378 295954
rect -2934 295398 -2698 295634
rect -2614 295398 -2378 295634
rect -2934 259718 -2698 259954
rect -2614 259718 -2378 259954
rect -2934 259398 -2698 259634
rect -2614 259398 -2378 259634
rect -2934 223718 -2698 223954
rect -2614 223718 -2378 223954
rect -2934 223398 -2698 223634
rect -2614 223398 -2378 223634
rect -2934 187718 -2698 187954
rect -2614 187718 -2378 187954
rect -2934 187398 -2698 187634
rect -2614 187398 -2378 187634
rect -2934 151718 -2698 151954
rect -2614 151718 -2378 151954
rect -2934 151398 -2698 151634
rect -2614 151398 -2378 151634
rect -2934 115718 -2698 115954
rect -2614 115718 -2378 115954
rect -2934 115398 -2698 115634
rect -2614 115398 -2378 115634
rect -2934 79718 -2698 79954
rect -2614 79718 -2378 79954
rect -2934 79398 -2698 79634
rect -2614 79398 -2378 79634
rect -2934 43718 -2698 43954
rect -2614 43718 -2378 43954
rect -2934 43398 -2698 43634
rect -2614 43398 -2378 43634
rect -2934 7718 -2698 7954
rect -2614 7718 -2378 7954
rect -2934 7398 -2698 7634
rect -2614 7398 -2378 7634
rect -1974 704602 -1738 704838
rect -1654 704602 -1418 704838
rect -1974 704282 -1738 704518
rect -1654 704282 -1418 704518
rect -1974 687218 -1738 687454
rect -1654 687218 -1418 687454
rect -1974 686898 -1738 687134
rect -1654 686898 -1418 687134
rect -1974 651218 -1738 651454
rect -1654 651218 -1418 651454
rect -1974 650898 -1738 651134
rect -1654 650898 -1418 651134
rect -1974 615218 -1738 615454
rect -1654 615218 -1418 615454
rect -1974 614898 -1738 615134
rect -1654 614898 -1418 615134
rect -1974 579218 -1738 579454
rect -1654 579218 -1418 579454
rect -1974 578898 -1738 579134
rect -1654 578898 -1418 579134
rect -1974 543218 -1738 543454
rect -1654 543218 -1418 543454
rect -1974 542898 -1738 543134
rect -1654 542898 -1418 543134
rect -1974 507218 -1738 507454
rect -1654 507218 -1418 507454
rect -1974 506898 -1738 507134
rect -1654 506898 -1418 507134
rect -1974 471218 -1738 471454
rect -1654 471218 -1418 471454
rect -1974 470898 -1738 471134
rect -1654 470898 -1418 471134
rect -1974 435218 -1738 435454
rect -1654 435218 -1418 435454
rect -1974 434898 -1738 435134
rect -1654 434898 -1418 435134
rect -1974 399218 -1738 399454
rect -1654 399218 -1418 399454
rect -1974 398898 -1738 399134
rect -1654 398898 -1418 399134
rect -1974 363218 -1738 363454
rect -1654 363218 -1418 363454
rect -1974 362898 -1738 363134
rect -1654 362898 -1418 363134
rect -1974 327218 -1738 327454
rect -1654 327218 -1418 327454
rect -1974 326898 -1738 327134
rect -1654 326898 -1418 327134
rect -1974 291218 -1738 291454
rect -1654 291218 -1418 291454
rect -1974 290898 -1738 291134
rect -1654 290898 -1418 291134
rect -1974 255218 -1738 255454
rect -1654 255218 -1418 255454
rect -1974 254898 -1738 255134
rect -1654 254898 -1418 255134
rect -1974 219218 -1738 219454
rect -1654 219218 -1418 219454
rect -1974 218898 -1738 219134
rect -1654 218898 -1418 219134
rect -1974 183218 -1738 183454
rect -1654 183218 -1418 183454
rect -1974 182898 -1738 183134
rect -1654 182898 -1418 183134
rect -1974 147218 -1738 147454
rect -1654 147218 -1418 147454
rect -1974 146898 -1738 147134
rect -1654 146898 -1418 147134
rect -1974 111218 -1738 111454
rect -1654 111218 -1418 111454
rect -1974 110898 -1738 111134
rect -1654 110898 -1418 111134
rect -1974 75218 -1738 75454
rect -1654 75218 -1418 75454
rect -1974 74898 -1738 75134
rect -1654 74898 -1418 75134
rect -1974 39218 -1738 39454
rect -1654 39218 -1418 39454
rect -1974 38898 -1738 39134
rect -1654 38898 -1418 39134
rect -1974 3218 -1738 3454
rect -1654 3218 -1418 3454
rect -1974 2898 -1738 3134
rect -1654 2898 -1418 3134
rect -1974 -582 -1738 -346
rect -1654 -582 -1418 -346
rect -1974 -902 -1738 -666
rect -1654 -902 -1418 -666
rect 1826 704602 2062 704838
rect 2146 704602 2382 704838
rect 1826 704282 2062 704518
rect 2146 704282 2382 704518
rect 1826 687218 2062 687454
rect 2146 687218 2382 687454
rect 1826 686898 2062 687134
rect 2146 686898 2382 687134
rect 1826 651218 2062 651454
rect 2146 651218 2382 651454
rect 1826 650898 2062 651134
rect 2146 650898 2382 651134
rect 1826 615218 2062 615454
rect 2146 615218 2382 615454
rect 1826 614898 2062 615134
rect 2146 614898 2382 615134
rect 1826 579218 2062 579454
rect 2146 579218 2382 579454
rect 1826 578898 2062 579134
rect 2146 578898 2382 579134
rect 1826 543218 2062 543454
rect 2146 543218 2382 543454
rect 1826 542898 2062 543134
rect 2146 542898 2382 543134
rect 1826 507218 2062 507454
rect 2146 507218 2382 507454
rect 1826 506898 2062 507134
rect 2146 506898 2382 507134
rect 1826 471218 2062 471454
rect 2146 471218 2382 471454
rect 1826 470898 2062 471134
rect 2146 470898 2382 471134
rect 1826 435218 2062 435454
rect 2146 435218 2382 435454
rect 1826 434898 2062 435134
rect 2146 434898 2382 435134
rect 1826 399218 2062 399454
rect 2146 399218 2382 399454
rect 1826 398898 2062 399134
rect 2146 398898 2382 399134
rect 1826 363218 2062 363454
rect 2146 363218 2382 363454
rect 1826 362898 2062 363134
rect 2146 362898 2382 363134
rect 1826 327218 2062 327454
rect 2146 327218 2382 327454
rect 1826 326898 2062 327134
rect 2146 326898 2382 327134
rect 1826 291218 2062 291454
rect 2146 291218 2382 291454
rect 1826 290898 2062 291134
rect 2146 290898 2382 291134
rect 1826 255218 2062 255454
rect 2146 255218 2382 255454
rect 1826 254898 2062 255134
rect 2146 254898 2382 255134
rect 1826 219218 2062 219454
rect 2146 219218 2382 219454
rect 1826 218898 2062 219134
rect 2146 218898 2382 219134
rect 1826 183218 2062 183454
rect 2146 183218 2382 183454
rect 1826 182898 2062 183134
rect 2146 182898 2382 183134
rect 1826 147218 2062 147454
rect 2146 147218 2382 147454
rect 1826 146898 2062 147134
rect 2146 146898 2382 147134
rect 1826 111218 2062 111454
rect 2146 111218 2382 111454
rect 1826 110898 2062 111134
rect 2146 110898 2382 111134
rect 1826 75218 2062 75454
rect 2146 75218 2382 75454
rect 1826 74898 2062 75134
rect 2146 74898 2382 75134
rect 1826 39218 2062 39454
rect 2146 39218 2382 39454
rect 1826 38898 2062 39134
rect 2146 38898 2382 39134
rect 1826 3218 2062 3454
rect 2146 3218 2382 3454
rect 1826 2898 2062 3134
rect 2146 2898 2382 3134
rect 1826 -582 2062 -346
rect 2146 -582 2382 -346
rect 1826 -902 2062 -666
rect 2146 -902 2382 -666
rect -2934 -1542 -2698 -1306
rect -2614 -1542 -2378 -1306
rect -2934 -1862 -2698 -1626
rect -2614 -1862 -2378 -1626
rect -3894 -2502 -3658 -2266
rect -3574 -2502 -3338 -2266
rect -3894 -2822 -3658 -2586
rect -3574 -2822 -3338 -2586
rect -4854 -3462 -4618 -3226
rect -4534 -3462 -4298 -3226
rect -4854 -3782 -4618 -3546
rect -4534 -3782 -4298 -3546
rect -5814 -4422 -5578 -4186
rect -5494 -4422 -5258 -4186
rect -5814 -4742 -5578 -4506
rect -5494 -4742 -5258 -4506
rect -6774 -5382 -6538 -5146
rect -6454 -5382 -6218 -5146
rect -6774 -5702 -6538 -5466
rect -6454 -5702 -6218 -5466
rect -7734 -6342 -7498 -6106
rect -7414 -6342 -7178 -6106
rect -7734 -6662 -7498 -6426
rect -7414 -6662 -7178 -6426
rect -8694 -7302 -8458 -7066
rect -8374 -7302 -8138 -7066
rect -8694 -7622 -8458 -7386
rect -8374 -7622 -8138 -7386
rect 6326 705562 6562 705798
rect 6646 705562 6882 705798
rect 6326 705242 6562 705478
rect 6646 705242 6882 705478
rect 6326 691718 6562 691954
rect 6646 691718 6882 691954
rect 6326 691398 6562 691634
rect 6646 691398 6882 691634
rect 6326 655718 6562 655954
rect 6646 655718 6882 655954
rect 6326 655398 6562 655634
rect 6646 655398 6882 655634
rect 6326 619718 6562 619954
rect 6646 619718 6882 619954
rect 6326 619398 6562 619634
rect 6646 619398 6882 619634
rect 6326 583718 6562 583954
rect 6646 583718 6882 583954
rect 6326 583398 6562 583634
rect 6646 583398 6882 583634
rect 6326 547718 6562 547954
rect 6646 547718 6882 547954
rect 6326 547398 6562 547634
rect 6646 547398 6882 547634
rect 6326 511718 6562 511954
rect 6646 511718 6882 511954
rect 6326 511398 6562 511634
rect 6646 511398 6882 511634
rect 6326 475718 6562 475954
rect 6646 475718 6882 475954
rect 6326 475398 6562 475634
rect 6646 475398 6882 475634
rect 6326 439718 6562 439954
rect 6646 439718 6882 439954
rect 6326 439398 6562 439634
rect 6646 439398 6882 439634
rect 6326 403718 6562 403954
rect 6646 403718 6882 403954
rect 6326 403398 6562 403634
rect 6646 403398 6882 403634
rect 6326 367718 6562 367954
rect 6646 367718 6882 367954
rect 6326 367398 6562 367634
rect 6646 367398 6882 367634
rect 6326 331718 6562 331954
rect 6646 331718 6882 331954
rect 6326 331398 6562 331634
rect 6646 331398 6882 331634
rect 6326 295718 6562 295954
rect 6646 295718 6882 295954
rect 6326 295398 6562 295634
rect 6646 295398 6882 295634
rect 6326 259718 6562 259954
rect 6646 259718 6882 259954
rect 6326 259398 6562 259634
rect 6646 259398 6882 259634
rect 6326 223718 6562 223954
rect 6646 223718 6882 223954
rect 6326 223398 6562 223634
rect 6646 223398 6882 223634
rect 6326 187718 6562 187954
rect 6646 187718 6882 187954
rect 6326 187398 6562 187634
rect 6646 187398 6882 187634
rect 6326 151718 6562 151954
rect 6646 151718 6882 151954
rect 6326 151398 6562 151634
rect 6646 151398 6882 151634
rect 6326 115718 6562 115954
rect 6646 115718 6882 115954
rect 6326 115398 6562 115634
rect 6646 115398 6882 115634
rect 6326 79718 6562 79954
rect 6646 79718 6882 79954
rect 6326 79398 6562 79634
rect 6646 79398 6882 79634
rect 6326 43718 6562 43954
rect 6646 43718 6882 43954
rect 6326 43398 6562 43634
rect 6646 43398 6882 43634
rect 6326 7718 6562 7954
rect 6646 7718 6882 7954
rect 6326 7398 6562 7634
rect 6646 7398 6882 7634
rect 6326 -1542 6562 -1306
rect 6646 -1542 6882 -1306
rect 6326 -1862 6562 -1626
rect 6646 -1862 6882 -1626
rect 10826 706522 11062 706758
rect 11146 706522 11382 706758
rect 10826 706202 11062 706438
rect 11146 706202 11382 706438
rect 10826 696218 11062 696454
rect 11146 696218 11382 696454
rect 10826 695898 11062 696134
rect 11146 695898 11382 696134
rect 10826 660218 11062 660454
rect 11146 660218 11382 660454
rect 10826 659898 11062 660134
rect 11146 659898 11382 660134
rect 10826 624218 11062 624454
rect 11146 624218 11382 624454
rect 10826 623898 11062 624134
rect 11146 623898 11382 624134
rect 10826 588218 11062 588454
rect 11146 588218 11382 588454
rect 10826 587898 11062 588134
rect 11146 587898 11382 588134
rect 10826 552218 11062 552454
rect 11146 552218 11382 552454
rect 10826 551898 11062 552134
rect 11146 551898 11382 552134
rect 10826 516218 11062 516454
rect 11146 516218 11382 516454
rect 10826 515898 11062 516134
rect 11146 515898 11382 516134
rect 10826 480218 11062 480454
rect 11146 480218 11382 480454
rect 10826 479898 11062 480134
rect 11146 479898 11382 480134
rect 10826 444218 11062 444454
rect 11146 444218 11382 444454
rect 10826 443898 11062 444134
rect 11146 443898 11382 444134
rect 10826 408218 11062 408454
rect 11146 408218 11382 408454
rect 10826 407898 11062 408134
rect 11146 407898 11382 408134
rect 10826 372218 11062 372454
rect 11146 372218 11382 372454
rect 10826 371898 11062 372134
rect 11146 371898 11382 372134
rect 10826 336218 11062 336454
rect 11146 336218 11382 336454
rect 10826 335898 11062 336134
rect 11146 335898 11382 336134
rect 10826 300218 11062 300454
rect 11146 300218 11382 300454
rect 10826 299898 11062 300134
rect 11146 299898 11382 300134
rect 10826 264218 11062 264454
rect 11146 264218 11382 264454
rect 10826 263898 11062 264134
rect 11146 263898 11382 264134
rect 10826 228218 11062 228454
rect 11146 228218 11382 228454
rect 10826 227898 11062 228134
rect 11146 227898 11382 228134
rect 10826 192218 11062 192454
rect 11146 192218 11382 192454
rect 10826 191898 11062 192134
rect 11146 191898 11382 192134
rect 10826 156218 11062 156454
rect 11146 156218 11382 156454
rect 10826 155898 11062 156134
rect 11146 155898 11382 156134
rect 10826 120218 11062 120454
rect 11146 120218 11382 120454
rect 10826 119898 11062 120134
rect 11146 119898 11382 120134
rect 10826 84218 11062 84454
rect 11146 84218 11382 84454
rect 10826 83898 11062 84134
rect 11146 83898 11382 84134
rect 10826 48218 11062 48454
rect 11146 48218 11382 48454
rect 10826 47898 11062 48134
rect 11146 47898 11382 48134
rect 10826 12218 11062 12454
rect 11146 12218 11382 12454
rect 10826 11898 11062 12134
rect 11146 11898 11382 12134
rect 10826 -2502 11062 -2266
rect 11146 -2502 11382 -2266
rect 10826 -2822 11062 -2586
rect 11146 -2822 11382 -2586
rect 15326 707482 15562 707718
rect 15646 707482 15882 707718
rect 15326 707162 15562 707398
rect 15646 707162 15882 707398
rect 15326 700718 15562 700954
rect 15646 700718 15882 700954
rect 15326 700398 15562 700634
rect 15646 700398 15882 700634
rect 15326 664718 15562 664954
rect 15646 664718 15882 664954
rect 15326 664398 15562 664634
rect 15646 664398 15882 664634
rect 15326 628718 15562 628954
rect 15646 628718 15882 628954
rect 15326 628398 15562 628634
rect 15646 628398 15882 628634
rect 15326 592718 15562 592954
rect 15646 592718 15882 592954
rect 15326 592398 15562 592634
rect 15646 592398 15882 592634
rect 15326 556718 15562 556954
rect 15646 556718 15882 556954
rect 15326 556398 15562 556634
rect 15646 556398 15882 556634
rect 15326 520718 15562 520954
rect 15646 520718 15882 520954
rect 15326 520398 15562 520634
rect 15646 520398 15882 520634
rect 15326 484718 15562 484954
rect 15646 484718 15882 484954
rect 15326 484398 15562 484634
rect 15646 484398 15882 484634
rect 15326 448718 15562 448954
rect 15646 448718 15882 448954
rect 15326 448398 15562 448634
rect 15646 448398 15882 448634
rect 15326 412718 15562 412954
rect 15646 412718 15882 412954
rect 15326 412398 15562 412634
rect 15646 412398 15882 412634
rect 15326 376718 15562 376954
rect 15646 376718 15882 376954
rect 15326 376398 15562 376634
rect 15646 376398 15882 376634
rect 15326 340718 15562 340954
rect 15646 340718 15882 340954
rect 15326 340398 15562 340634
rect 15646 340398 15882 340634
rect 15326 304718 15562 304954
rect 15646 304718 15882 304954
rect 15326 304398 15562 304634
rect 15646 304398 15882 304634
rect 15326 268718 15562 268954
rect 15646 268718 15882 268954
rect 15326 268398 15562 268634
rect 15646 268398 15882 268634
rect 15326 232718 15562 232954
rect 15646 232718 15882 232954
rect 15326 232398 15562 232634
rect 15646 232398 15882 232634
rect 15326 196718 15562 196954
rect 15646 196718 15882 196954
rect 15326 196398 15562 196634
rect 15646 196398 15882 196634
rect 15326 160718 15562 160954
rect 15646 160718 15882 160954
rect 15326 160398 15562 160634
rect 15646 160398 15882 160634
rect 15326 124718 15562 124954
rect 15646 124718 15882 124954
rect 15326 124398 15562 124634
rect 15646 124398 15882 124634
rect 15326 88718 15562 88954
rect 15646 88718 15882 88954
rect 15326 88398 15562 88634
rect 15646 88398 15882 88634
rect 15326 52718 15562 52954
rect 15646 52718 15882 52954
rect 15326 52398 15562 52634
rect 15646 52398 15882 52634
rect 15326 16718 15562 16954
rect 15646 16718 15882 16954
rect 15326 16398 15562 16634
rect 15646 16398 15882 16634
rect 15326 -3462 15562 -3226
rect 15646 -3462 15882 -3226
rect 15326 -3782 15562 -3546
rect 15646 -3782 15882 -3546
rect 19826 708442 20062 708678
rect 20146 708442 20382 708678
rect 19826 708122 20062 708358
rect 20146 708122 20382 708358
rect 19826 669218 20062 669454
rect 20146 669218 20382 669454
rect 19826 668898 20062 669134
rect 20146 668898 20382 669134
rect 19826 633218 20062 633454
rect 20146 633218 20382 633454
rect 19826 632898 20062 633134
rect 20146 632898 20382 633134
rect 19826 597218 20062 597454
rect 20146 597218 20382 597454
rect 19826 596898 20062 597134
rect 20146 596898 20382 597134
rect 19826 561218 20062 561454
rect 20146 561218 20382 561454
rect 19826 560898 20062 561134
rect 20146 560898 20382 561134
rect 19826 525218 20062 525454
rect 20146 525218 20382 525454
rect 19826 524898 20062 525134
rect 20146 524898 20382 525134
rect 19826 489218 20062 489454
rect 20146 489218 20382 489454
rect 19826 488898 20062 489134
rect 20146 488898 20382 489134
rect 19826 453218 20062 453454
rect 20146 453218 20382 453454
rect 19826 452898 20062 453134
rect 20146 452898 20382 453134
rect 19826 417218 20062 417454
rect 20146 417218 20382 417454
rect 19826 416898 20062 417134
rect 20146 416898 20382 417134
rect 19826 381218 20062 381454
rect 20146 381218 20382 381454
rect 19826 380898 20062 381134
rect 20146 380898 20382 381134
rect 19826 345218 20062 345454
rect 20146 345218 20382 345454
rect 19826 344898 20062 345134
rect 20146 344898 20382 345134
rect 19826 309218 20062 309454
rect 20146 309218 20382 309454
rect 19826 308898 20062 309134
rect 20146 308898 20382 309134
rect 19826 273218 20062 273454
rect 20146 273218 20382 273454
rect 19826 272898 20062 273134
rect 20146 272898 20382 273134
rect 19826 237218 20062 237454
rect 20146 237218 20382 237454
rect 19826 236898 20062 237134
rect 20146 236898 20382 237134
rect 19826 201218 20062 201454
rect 20146 201218 20382 201454
rect 19826 200898 20062 201134
rect 20146 200898 20382 201134
rect 19826 165218 20062 165454
rect 20146 165218 20382 165454
rect 19826 164898 20062 165134
rect 20146 164898 20382 165134
rect 19826 129218 20062 129454
rect 20146 129218 20382 129454
rect 19826 128898 20062 129134
rect 20146 128898 20382 129134
rect 19826 93218 20062 93454
rect 20146 93218 20382 93454
rect 19826 92898 20062 93134
rect 20146 92898 20382 93134
rect 19826 57218 20062 57454
rect 20146 57218 20382 57454
rect 19826 56898 20062 57134
rect 20146 56898 20382 57134
rect 19826 21218 20062 21454
rect 20146 21218 20382 21454
rect 19826 20898 20062 21134
rect 20146 20898 20382 21134
rect 19826 -4422 20062 -4186
rect 20146 -4422 20382 -4186
rect 19826 -4742 20062 -4506
rect 20146 -4742 20382 -4506
rect 24326 709402 24562 709638
rect 24646 709402 24882 709638
rect 24326 709082 24562 709318
rect 24646 709082 24882 709318
rect 24326 673718 24562 673954
rect 24646 673718 24882 673954
rect 24326 673398 24562 673634
rect 24646 673398 24882 673634
rect 24326 637718 24562 637954
rect 24646 637718 24882 637954
rect 24326 637398 24562 637634
rect 24646 637398 24882 637634
rect 24326 601718 24562 601954
rect 24646 601718 24882 601954
rect 24326 601398 24562 601634
rect 24646 601398 24882 601634
rect 24326 565718 24562 565954
rect 24646 565718 24882 565954
rect 24326 565398 24562 565634
rect 24646 565398 24882 565634
rect 24326 529718 24562 529954
rect 24646 529718 24882 529954
rect 24326 529398 24562 529634
rect 24646 529398 24882 529634
rect 24326 493718 24562 493954
rect 24646 493718 24882 493954
rect 24326 493398 24562 493634
rect 24646 493398 24882 493634
rect 24326 457718 24562 457954
rect 24646 457718 24882 457954
rect 24326 457398 24562 457634
rect 24646 457398 24882 457634
rect 24326 421718 24562 421954
rect 24646 421718 24882 421954
rect 24326 421398 24562 421634
rect 24646 421398 24882 421634
rect 24326 385718 24562 385954
rect 24646 385718 24882 385954
rect 24326 385398 24562 385634
rect 24646 385398 24882 385634
rect 24326 349718 24562 349954
rect 24646 349718 24882 349954
rect 24326 349398 24562 349634
rect 24646 349398 24882 349634
rect 24326 313718 24562 313954
rect 24646 313718 24882 313954
rect 24326 313398 24562 313634
rect 24646 313398 24882 313634
rect 24326 277718 24562 277954
rect 24646 277718 24882 277954
rect 24326 277398 24562 277634
rect 24646 277398 24882 277634
rect 24326 241718 24562 241954
rect 24646 241718 24882 241954
rect 24326 241398 24562 241634
rect 24646 241398 24882 241634
rect 24326 205718 24562 205954
rect 24646 205718 24882 205954
rect 24326 205398 24562 205634
rect 24646 205398 24882 205634
rect 24326 169718 24562 169954
rect 24646 169718 24882 169954
rect 24326 169398 24562 169634
rect 24646 169398 24882 169634
rect 24326 133718 24562 133954
rect 24646 133718 24882 133954
rect 24326 133398 24562 133634
rect 24646 133398 24882 133634
rect 24326 97718 24562 97954
rect 24646 97718 24882 97954
rect 24326 97398 24562 97634
rect 24646 97398 24882 97634
rect 24326 61718 24562 61954
rect 24646 61718 24882 61954
rect 24326 61398 24562 61634
rect 24646 61398 24882 61634
rect 24326 25718 24562 25954
rect 24646 25718 24882 25954
rect 24326 25398 24562 25634
rect 24646 25398 24882 25634
rect 24326 -5382 24562 -5146
rect 24646 -5382 24882 -5146
rect 24326 -5702 24562 -5466
rect 24646 -5702 24882 -5466
rect 28826 710362 29062 710598
rect 29146 710362 29382 710598
rect 28826 710042 29062 710278
rect 29146 710042 29382 710278
rect 28826 678218 29062 678454
rect 29146 678218 29382 678454
rect 28826 677898 29062 678134
rect 29146 677898 29382 678134
rect 28826 642218 29062 642454
rect 29146 642218 29382 642454
rect 28826 641898 29062 642134
rect 29146 641898 29382 642134
rect 28826 606218 29062 606454
rect 29146 606218 29382 606454
rect 28826 605898 29062 606134
rect 29146 605898 29382 606134
rect 28826 570218 29062 570454
rect 29146 570218 29382 570454
rect 28826 569898 29062 570134
rect 29146 569898 29382 570134
rect 28826 534218 29062 534454
rect 29146 534218 29382 534454
rect 28826 533898 29062 534134
rect 29146 533898 29382 534134
rect 28826 498218 29062 498454
rect 29146 498218 29382 498454
rect 28826 497898 29062 498134
rect 29146 497898 29382 498134
rect 28826 462218 29062 462454
rect 29146 462218 29382 462454
rect 28826 461898 29062 462134
rect 29146 461898 29382 462134
rect 28826 426218 29062 426454
rect 29146 426218 29382 426454
rect 28826 425898 29062 426134
rect 29146 425898 29382 426134
rect 28826 390218 29062 390454
rect 29146 390218 29382 390454
rect 28826 389898 29062 390134
rect 29146 389898 29382 390134
rect 28826 354218 29062 354454
rect 29146 354218 29382 354454
rect 28826 353898 29062 354134
rect 29146 353898 29382 354134
rect 28826 318218 29062 318454
rect 29146 318218 29382 318454
rect 28826 317898 29062 318134
rect 29146 317898 29382 318134
rect 28826 282218 29062 282454
rect 29146 282218 29382 282454
rect 28826 281898 29062 282134
rect 29146 281898 29382 282134
rect 28826 246218 29062 246454
rect 29146 246218 29382 246454
rect 28826 245898 29062 246134
rect 29146 245898 29382 246134
rect 28826 210218 29062 210454
rect 29146 210218 29382 210454
rect 28826 209898 29062 210134
rect 29146 209898 29382 210134
rect 28826 174218 29062 174454
rect 29146 174218 29382 174454
rect 28826 173898 29062 174134
rect 29146 173898 29382 174134
rect 28826 138218 29062 138454
rect 29146 138218 29382 138454
rect 28826 137898 29062 138134
rect 29146 137898 29382 138134
rect 28826 102218 29062 102454
rect 29146 102218 29382 102454
rect 28826 101898 29062 102134
rect 29146 101898 29382 102134
rect 28826 66218 29062 66454
rect 29146 66218 29382 66454
rect 28826 65898 29062 66134
rect 29146 65898 29382 66134
rect 28826 30218 29062 30454
rect 29146 30218 29382 30454
rect 28826 29898 29062 30134
rect 29146 29898 29382 30134
rect 28826 -6342 29062 -6106
rect 29146 -6342 29382 -6106
rect 28826 -6662 29062 -6426
rect 29146 -6662 29382 -6426
rect 33326 711322 33562 711558
rect 33646 711322 33882 711558
rect 33326 711002 33562 711238
rect 33646 711002 33882 711238
rect 33326 682718 33562 682954
rect 33646 682718 33882 682954
rect 33326 682398 33562 682634
rect 33646 682398 33882 682634
rect 33326 646718 33562 646954
rect 33646 646718 33882 646954
rect 33326 646398 33562 646634
rect 33646 646398 33882 646634
rect 33326 610718 33562 610954
rect 33646 610718 33882 610954
rect 33326 610398 33562 610634
rect 33646 610398 33882 610634
rect 33326 574718 33562 574954
rect 33646 574718 33882 574954
rect 33326 574398 33562 574634
rect 33646 574398 33882 574634
rect 33326 538718 33562 538954
rect 33646 538718 33882 538954
rect 33326 538398 33562 538634
rect 33646 538398 33882 538634
rect 33326 502718 33562 502954
rect 33646 502718 33882 502954
rect 33326 502398 33562 502634
rect 33646 502398 33882 502634
rect 33326 466718 33562 466954
rect 33646 466718 33882 466954
rect 33326 466398 33562 466634
rect 33646 466398 33882 466634
rect 33326 430718 33562 430954
rect 33646 430718 33882 430954
rect 33326 430398 33562 430634
rect 33646 430398 33882 430634
rect 33326 394718 33562 394954
rect 33646 394718 33882 394954
rect 33326 394398 33562 394634
rect 33646 394398 33882 394634
rect 33326 358718 33562 358954
rect 33646 358718 33882 358954
rect 33326 358398 33562 358634
rect 33646 358398 33882 358634
rect 33326 322718 33562 322954
rect 33646 322718 33882 322954
rect 33326 322398 33562 322634
rect 33646 322398 33882 322634
rect 33326 286718 33562 286954
rect 33646 286718 33882 286954
rect 33326 286398 33562 286634
rect 33646 286398 33882 286634
rect 33326 250718 33562 250954
rect 33646 250718 33882 250954
rect 33326 250398 33562 250634
rect 33646 250398 33882 250634
rect 33326 214718 33562 214954
rect 33646 214718 33882 214954
rect 33326 214398 33562 214634
rect 33646 214398 33882 214634
rect 33326 178718 33562 178954
rect 33646 178718 33882 178954
rect 33326 178398 33562 178634
rect 33646 178398 33882 178634
rect 33326 142718 33562 142954
rect 33646 142718 33882 142954
rect 33326 142398 33562 142634
rect 33646 142398 33882 142634
rect 33326 106718 33562 106954
rect 33646 106718 33882 106954
rect 33326 106398 33562 106634
rect 33646 106398 33882 106634
rect 33326 70718 33562 70954
rect 33646 70718 33882 70954
rect 33326 70398 33562 70634
rect 33646 70398 33882 70634
rect 33326 34718 33562 34954
rect 33646 34718 33882 34954
rect 33326 34398 33562 34634
rect 33646 34398 33882 34634
rect 33326 -7302 33562 -7066
rect 33646 -7302 33882 -7066
rect 33326 -7622 33562 -7386
rect 33646 -7622 33882 -7386
rect 37826 704602 38062 704838
rect 38146 704602 38382 704838
rect 37826 704282 38062 704518
rect 38146 704282 38382 704518
rect 37826 687218 38062 687454
rect 38146 687218 38382 687454
rect 37826 686898 38062 687134
rect 38146 686898 38382 687134
rect 37826 651218 38062 651454
rect 38146 651218 38382 651454
rect 37826 650898 38062 651134
rect 38146 650898 38382 651134
rect 37826 615218 38062 615454
rect 38146 615218 38382 615454
rect 37826 614898 38062 615134
rect 38146 614898 38382 615134
rect 37826 579218 38062 579454
rect 38146 579218 38382 579454
rect 37826 578898 38062 579134
rect 38146 578898 38382 579134
rect 37826 543218 38062 543454
rect 38146 543218 38382 543454
rect 37826 542898 38062 543134
rect 38146 542898 38382 543134
rect 37826 507218 38062 507454
rect 38146 507218 38382 507454
rect 37826 506898 38062 507134
rect 38146 506898 38382 507134
rect 37826 471218 38062 471454
rect 38146 471218 38382 471454
rect 37826 470898 38062 471134
rect 38146 470898 38382 471134
rect 37826 435218 38062 435454
rect 38146 435218 38382 435454
rect 37826 434898 38062 435134
rect 38146 434898 38382 435134
rect 37826 399218 38062 399454
rect 38146 399218 38382 399454
rect 37826 398898 38062 399134
rect 38146 398898 38382 399134
rect 37826 363218 38062 363454
rect 38146 363218 38382 363454
rect 37826 362898 38062 363134
rect 38146 362898 38382 363134
rect 37826 327218 38062 327454
rect 38146 327218 38382 327454
rect 37826 326898 38062 327134
rect 38146 326898 38382 327134
rect 37826 291218 38062 291454
rect 38146 291218 38382 291454
rect 37826 290898 38062 291134
rect 38146 290898 38382 291134
rect 37826 255218 38062 255454
rect 38146 255218 38382 255454
rect 37826 254898 38062 255134
rect 38146 254898 38382 255134
rect 37826 219218 38062 219454
rect 38146 219218 38382 219454
rect 37826 218898 38062 219134
rect 38146 218898 38382 219134
rect 37826 183218 38062 183454
rect 38146 183218 38382 183454
rect 37826 182898 38062 183134
rect 38146 182898 38382 183134
rect 37826 147218 38062 147454
rect 38146 147218 38382 147454
rect 37826 146898 38062 147134
rect 38146 146898 38382 147134
rect 37826 111218 38062 111454
rect 38146 111218 38382 111454
rect 37826 110898 38062 111134
rect 38146 110898 38382 111134
rect 37826 75218 38062 75454
rect 38146 75218 38382 75454
rect 37826 74898 38062 75134
rect 38146 74898 38382 75134
rect 37826 39218 38062 39454
rect 38146 39218 38382 39454
rect 37826 38898 38062 39134
rect 38146 38898 38382 39134
rect 37826 3218 38062 3454
rect 38146 3218 38382 3454
rect 37826 2898 38062 3134
rect 38146 2898 38382 3134
rect 37826 -582 38062 -346
rect 38146 -582 38382 -346
rect 37826 -902 38062 -666
rect 38146 -902 38382 -666
rect 42326 705562 42562 705798
rect 42646 705562 42882 705798
rect 42326 705242 42562 705478
rect 42646 705242 42882 705478
rect 42326 691718 42562 691954
rect 42646 691718 42882 691954
rect 42326 691398 42562 691634
rect 42646 691398 42882 691634
rect 42326 655718 42562 655954
rect 42646 655718 42882 655954
rect 42326 655398 42562 655634
rect 42646 655398 42882 655634
rect 42326 619718 42562 619954
rect 42646 619718 42882 619954
rect 42326 619398 42562 619634
rect 42646 619398 42882 619634
rect 42326 583718 42562 583954
rect 42646 583718 42882 583954
rect 42326 583398 42562 583634
rect 42646 583398 42882 583634
rect 42326 547718 42562 547954
rect 42646 547718 42882 547954
rect 42326 547398 42562 547634
rect 42646 547398 42882 547634
rect 42326 511718 42562 511954
rect 42646 511718 42882 511954
rect 42326 511398 42562 511634
rect 42646 511398 42882 511634
rect 42326 475718 42562 475954
rect 42646 475718 42882 475954
rect 42326 475398 42562 475634
rect 42646 475398 42882 475634
rect 42326 439718 42562 439954
rect 42646 439718 42882 439954
rect 42326 439398 42562 439634
rect 42646 439398 42882 439634
rect 42326 403718 42562 403954
rect 42646 403718 42882 403954
rect 42326 403398 42562 403634
rect 42646 403398 42882 403634
rect 42326 367718 42562 367954
rect 42646 367718 42882 367954
rect 42326 367398 42562 367634
rect 42646 367398 42882 367634
rect 42326 331718 42562 331954
rect 42646 331718 42882 331954
rect 42326 331398 42562 331634
rect 42646 331398 42882 331634
rect 42326 295718 42562 295954
rect 42646 295718 42882 295954
rect 42326 295398 42562 295634
rect 42646 295398 42882 295634
rect 42326 259718 42562 259954
rect 42646 259718 42882 259954
rect 42326 259398 42562 259634
rect 42646 259398 42882 259634
rect 42326 223718 42562 223954
rect 42646 223718 42882 223954
rect 42326 223398 42562 223634
rect 42646 223398 42882 223634
rect 42326 187718 42562 187954
rect 42646 187718 42882 187954
rect 42326 187398 42562 187634
rect 42646 187398 42882 187634
rect 42326 151718 42562 151954
rect 42646 151718 42882 151954
rect 42326 151398 42562 151634
rect 42646 151398 42882 151634
rect 42326 115718 42562 115954
rect 42646 115718 42882 115954
rect 42326 115398 42562 115634
rect 42646 115398 42882 115634
rect 42326 79718 42562 79954
rect 42646 79718 42882 79954
rect 42326 79398 42562 79634
rect 42646 79398 42882 79634
rect 42326 43718 42562 43954
rect 42646 43718 42882 43954
rect 42326 43398 42562 43634
rect 42646 43398 42882 43634
rect 42326 7718 42562 7954
rect 42646 7718 42882 7954
rect 42326 7398 42562 7634
rect 42646 7398 42882 7634
rect 42326 -1542 42562 -1306
rect 42646 -1542 42882 -1306
rect 42326 -1862 42562 -1626
rect 42646 -1862 42882 -1626
rect 46826 706522 47062 706758
rect 47146 706522 47382 706758
rect 46826 706202 47062 706438
rect 47146 706202 47382 706438
rect 46826 696218 47062 696454
rect 47146 696218 47382 696454
rect 46826 695898 47062 696134
rect 47146 695898 47382 696134
rect 46826 660218 47062 660454
rect 47146 660218 47382 660454
rect 46826 659898 47062 660134
rect 47146 659898 47382 660134
rect 46826 624218 47062 624454
rect 47146 624218 47382 624454
rect 46826 623898 47062 624134
rect 47146 623898 47382 624134
rect 46826 588218 47062 588454
rect 47146 588218 47382 588454
rect 46826 587898 47062 588134
rect 47146 587898 47382 588134
rect 46826 552218 47062 552454
rect 47146 552218 47382 552454
rect 46826 551898 47062 552134
rect 47146 551898 47382 552134
rect 46826 516218 47062 516454
rect 47146 516218 47382 516454
rect 46826 515898 47062 516134
rect 47146 515898 47382 516134
rect 46826 480218 47062 480454
rect 47146 480218 47382 480454
rect 46826 479898 47062 480134
rect 47146 479898 47382 480134
rect 46826 444218 47062 444454
rect 47146 444218 47382 444454
rect 46826 443898 47062 444134
rect 47146 443898 47382 444134
rect 46826 408218 47062 408454
rect 47146 408218 47382 408454
rect 46826 407898 47062 408134
rect 47146 407898 47382 408134
rect 46826 372218 47062 372454
rect 47146 372218 47382 372454
rect 46826 371898 47062 372134
rect 47146 371898 47382 372134
rect 46826 336218 47062 336454
rect 47146 336218 47382 336454
rect 46826 335898 47062 336134
rect 47146 335898 47382 336134
rect 46826 300218 47062 300454
rect 47146 300218 47382 300454
rect 46826 299898 47062 300134
rect 47146 299898 47382 300134
rect 46826 264218 47062 264454
rect 47146 264218 47382 264454
rect 46826 263898 47062 264134
rect 47146 263898 47382 264134
rect 46826 228218 47062 228454
rect 47146 228218 47382 228454
rect 46826 227898 47062 228134
rect 47146 227898 47382 228134
rect 46826 192218 47062 192454
rect 47146 192218 47382 192454
rect 46826 191898 47062 192134
rect 47146 191898 47382 192134
rect 46826 156218 47062 156454
rect 47146 156218 47382 156454
rect 46826 155898 47062 156134
rect 47146 155898 47382 156134
rect 46826 120218 47062 120454
rect 47146 120218 47382 120454
rect 46826 119898 47062 120134
rect 47146 119898 47382 120134
rect 46826 84218 47062 84454
rect 47146 84218 47382 84454
rect 46826 83898 47062 84134
rect 47146 83898 47382 84134
rect 46826 48218 47062 48454
rect 47146 48218 47382 48454
rect 46826 47898 47062 48134
rect 47146 47898 47382 48134
rect 46826 12218 47062 12454
rect 47146 12218 47382 12454
rect 46826 11898 47062 12134
rect 47146 11898 47382 12134
rect 46826 -2502 47062 -2266
rect 47146 -2502 47382 -2266
rect 46826 -2822 47062 -2586
rect 47146 -2822 47382 -2586
rect 51326 707482 51562 707718
rect 51646 707482 51882 707718
rect 51326 707162 51562 707398
rect 51646 707162 51882 707398
rect 51326 700718 51562 700954
rect 51646 700718 51882 700954
rect 51326 700398 51562 700634
rect 51646 700398 51882 700634
rect 51326 664718 51562 664954
rect 51646 664718 51882 664954
rect 51326 664398 51562 664634
rect 51646 664398 51882 664634
rect 51326 628718 51562 628954
rect 51646 628718 51882 628954
rect 51326 628398 51562 628634
rect 51646 628398 51882 628634
rect 51326 592718 51562 592954
rect 51646 592718 51882 592954
rect 51326 592398 51562 592634
rect 51646 592398 51882 592634
rect 51326 556718 51562 556954
rect 51646 556718 51882 556954
rect 51326 556398 51562 556634
rect 51646 556398 51882 556634
rect 51326 520718 51562 520954
rect 51646 520718 51882 520954
rect 51326 520398 51562 520634
rect 51646 520398 51882 520634
rect 51326 484718 51562 484954
rect 51646 484718 51882 484954
rect 51326 484398 51562 484634
rect 51646 484398 51882 484634
rect 51326 448718 51562 448954
rect 51646 448718 51882 448954
rect 51326 448398 51562 448634
rect 51646 448398 51882 448634
rect 51326 412718 51562 412954
rect 51646 412718 51882 412954
rect 51326 412398 51562 412634
rect 51646 412398 51882 412634
rect 51326 376718 51562 376954
rect 51646 376718 51882 376954
rect 51326 376398 51562 376634
rect 51646 376398 51882 376634
rect 51326 340718 51562 340954
rect 51646 340718 51882 340954
rect 51326 340398 51562 340634
rect 51646 340398 51882 340634
rect 51326 304718 51562 304954
rect 51646 304718 51882 304954
rect 51326 304398 51562 304634
rect 51646 304398 51882 304634
rect 51326 268718 51562 268954
rect 51646 268718 51882 268954
rect 51326 268398 51562 268634
rect 51646 268398 51882 268634
rect 51326 232718 51562 232954
rect 51646 232718 51882 232954
rect 51326 232398 51562 232634
rect 51646 232398 51882 232634
rect 51326 196718 51562 196954
rect 51646 196718 51882 196954
rect 51326 196398 51562 196634
rect 51646 196398 51882 196634
rect 51326 160718 51562 160954
rect 51646 160718 51882 160954
rect 51326 160398 51562 160634
rect 51646 160398 51882 160634
rect 51326 124718 51562 124954
rect 51646 124718 51882 124954
rect 51326 124398 51562 124634
rect 51646 124398 51882 124634
rect 51326 88718 51562 88954
rect 51646 88718 51882 88954
rect 51326 88398 51562 88634
rect 51646 88398 51882 88634
rect 51326 52718 51562 52954
rect 51646 52718 51882 52954
rect 51326 52398 51562 52634
rect 51646 52398 51882 52634
rect 51326 16718 51562 16954
rect 51646 16718 51882 16954
rect 51326 16398 51562 16634
rect 51646 16398 51882 16634
rect 51326 -3462 51562 -3226
rect 51646 -3462 51882 -3226
rect 51326 -3782 51562 -3546
rect 51646 -3782 51882 -3546
rect 55826 708442 56062 708678
rect 56146 708442 56382 708678
rect 55826 708122 56062 708358
rect 56146 708122 56382 708358
rect 55826 669218 56062 669454
rect 56146 669218 56382 669454
rect 55826 668898 56062 669134
rect 56146 668898 56382 669134
rect 55826 633218 56062 633454
rect 56146 633218 56382 633454
rect 55826 632898 56062 633134
rect 56146 632898 56382 633134
rect 55826 597218 56062 597454
rect 56146 597218 56382 597454
rect 55826 596898 56062 597134
rect 56146 596898 56382 597134
rect 55826 561218 56062 561454
rect 56146 561218 56382 561454
rect 55826 560898 56062 561134
rect 56146 560898 56382 561134
rect 55826 525218 56062 525454
rect 56146 525218 56382 525454
rect 55826 524898 56062 525134
rect 56146 524898 56382 525134
rect 55826 489218 56062 489454
rect 56146 489218 56382 489454
rect 55826 488898 56062 489134
rect 56146 488898 56382 489134
rect 55826 453218 56062 453454
rect 56146 453218 56382 453454
rect 55826 452898 56062 453134
rect 56146 452898 56382 453134
rect 55826 417218 56062 417454
rect 56146 417218 56382 417454
rect 55826 416898 56062 417134
rect 56146 416898 56382 417134
rect 55826 381218 56062 381454
rect 56146 381218 56382 381454
rect 55826 380898 56062 381134
rect 56146 380898 56382 381134
rect 55826 345218 56062 345454
rect 56146 345218 56382 345454
rect 55826 344898 56062 345134
rect 56146 344898 56382 345134
rect 55826 309218 56062 309454
rect 56146 309218 56382 309454
rect 55826 308898 56062 309134
rect 56146 308898 56382 309134
rect 55826 273218 56062 273454
rect 56146 273218 56382 273454
rect 55826 272898 56062 273134
rect 56146 272898 56382 273134
rect 55826 237218 56062 237454
rect 56146 237218 56382 237454
rect 55826 236898 56062 237134
rect 56146 236898 56382 237134
rect 55826 201218 56062 201454
rect 56146 201218 56382 201454
rect 55826 200898 56062 201134
rect 56146 200898 56382 201134
rect 55826 165218 56062 165454
rect 56146 165218 56382 165454
rect 55826 164898 56062 165134
rect 56146 164898 56382 165134
rect 55826 129218 56062 129454
rect 56146 129218 56382 129454
rect 55826 128898 56062 129134
rect 56146 128898 56382 129134
rect 55826 93218 56062 93454
rect 56146 93218 56382 93454
rect 55826 92898 56062 93134
rect 56146 92898 56382 93134
rect 55826 57218 56062 57454
rect 56146 57218 56382 57454
rect 55826 56898 56062 57134
rect 56146 56898 56382 57134
rect 55826 21218 56062 21454
rect 56146 21218 56382 21454
rect 55826 20898 56062 21134
rect 56146 20898 56382 21134
rect 55826 -4422 56062 -4186
rect 56146 -4422 56382 -4186
rect 55826 -4742 56062 -4506
rect 56146 -4742 56382 -4506
rect 60326 709402 60562 709638
rect 60646 709402 60882 709638
rect 60326 709082 60562 709318
rect 60646 709082 60882 709318
rect 60326 673718 60562 673954
rect 60646 673718 60882 673954
rect 60326 673398 60562 673634
rect 60646 673398 60882 673634
rect 60326 637718 60562 637954
rect 60646 637718 60882 637954
rect 60326 637398 60562 637634
rect 60646 637398 60882 637634
rect 60326 601718 60562 601954
rect 60646 601718 60882 601954
rect 60326 601398 60562 601634
rect 60646 601398 60882 601634
rect 60326 565718 60562 565954
rect 60646 565718 60882 565954
rect 60326 565398 60562 565634
rect 60646 565398 60882 565634
rect 60326 529718 60562 529954
rect 60646 529718 60882 529954
rect 60326 529398 60562 529634
rect 60646 529398 60882 529634
rect 60326 493718 60562 493954
rect 60646 493718 60882 493954
rect 60326 493398 60562 493634
rect 60646 493398 60882 493634
rect 60326 457718 60562 457954
rect 60646 457718 60882 457954
rect 60326 457398 60562 457634
rect 60646 457398 60882 457634
rect 60326 421718 60562 421954
rect 60646 421718 60882 421954
rect 60326 421398 60562 421634
rect 60646 421398 60882 421634
rect 60326 385718 60562 385954
rect 60646 385718 60882 385954
rect 60326 385398 60562 385634
rect 60646 385398 60882 385634
rect 60326 349718 60562 349954
rect 60646 349718 60882 349954
rect 60326 349398 60562 349634
rect 60646 349398 60882 349634
rect 60326 313718 60562 313954
rect 60646 313718 60882 313954
rect 60326 313398 60562 313634
rect 60646 313398 60882 313634
rect 60326 277718 60562 277954
rect 60646 277718 60882 277954
rect 60326 277398 60562 277634
rect 60646 277398 60882 277634
rect 60326 241718 60562 241954
rect 60646 241718 60882 241954
rect 60326 241398 60562 241634
rect 60646 241398 60882 241634
rect 60326 205718 60562 205954
rect 60646 205718 60882 205954
rect 60326 205398 60562 205634
rect 60646 205398 60882 205634
rect 60326 169718 60562 169954
rect 60646 169718 60882 169954
rect 60326 169398 60562 169634
rect 60646 169398 60882 169634
rect 60326 133718 60562 133954
rect 60646 133718 60882 133954
rect 60326 133398 60562 133634
rect 60646 133398 60882 133634
rect 60326 97718 60562 97954
rect 60646 97718 60882 97954
rect 60326 97398 60562 97634
rect 60646 97398 60882 97634
rect 60326 61718 60562 61954
rect 60646 61718 60882 61954
rect 60326 61398 60562 61634
rect 60646 61398 60882 61634
rect 60326 25718 60562 25954
rect 60646 25718 60882 25954
rect 60326 25398 60562 25634
rect 60646 25398 60882 25634
rect 60326 -5382 60562 -5146
rect 60646 -5382 60882 -5146
rect 60326 -5702 60562 -5466
rect 60646 -5702 60882 -5466
rect 64826 710362 65062 710598
rect 65146 710362 65382 710598
rect 64826 710042 65062 710278
rect 65146 710042 65382 710278
rect 64826 678218 65062 678454
rect 65146 678218 65382 678454
rect 64826 677898 65062 678134
rect 65146 677898 65382 678134
rect 64826 642218 65062 642454
rect 65146 642218 65382 642454
rect 64826 641898 65062 642134
rect 65146 641898 65382 642134
rect 64826 606218 65062 606454
rect 65146 606218 65382 606454
rect 64826 605898 65062 606134
rect 65146 605898 65382 606134
rect 64826 570218 65062 570454
rect 65146 570218 65382 570454
rect 64826 569898 65062 570134
rect 65146 569898 65382 570134
rect 64826 534218 65062 534454
rect 65146 534218 65382 534454
rect 64826 533898 65062 534134
rect 65146 533898 65382 534134
rect 64826 498218 65062 498454
rect 65146 498218 65382 498454
rect 64826 497898 65062 498134
rect 65146 497898 65382 498134
rect 64826 462218 65062 462454
rect 65146 462218 65382 462454
rect 64826 461898 65062 462134
rect 65146 461898 65382 462134
rect 64826 426218 65062 426454
rect 65146 426218 65382 426454
rect 64826 425898 65062 426134
rect 65146 425898 65382 426134
rect 64826 390218 65062 390454
rect 65146 390218 65382 390454
rect 64826 389898 65062 390134
rect 65146 389898 65382 390134
rect 64826 354218 65062 354454
rect 65146 354218 65382 354454
rect 64826 353898 65062 354134
rect 65146 353898 65382 354134
rect 64826 318218 65062 318454
rect 65146 318218 65382 318454
rect 64826 317898 65062 318134
rect 65146 317898 65382 318134
rect 64826 282218 65062 282454
rect 65146 282218 65382 282454
rect 64826 281898 65062 282134
rect 65146 281898 65382 282134
rect 64826 246218 65062 246454
rect 65146 246218 65382 246454
rect 64826 245898 65062 246134
rect 65146 245898 65382 246134
rect 64826 210218 65062 210454
rect 65146 210218 65382 210454
rect 64826 209898 65062 210134
rect 65146 209898 65382 210134
rect 64826 174218 65062 174454
rect 65146 174218 65382 174454
rect 64826 173898 65062 174134
rect 65146 173898 65382 174134
rect 64826 138218 65062 138454
rect 65146 138218 65382 138454
rect 64826 137898 65062 138134
rect 65146 137898 65382 138134
rect 64826 102218 65062 102454
rect 65146 102218 65382 102454
rect 64826 101898 65062 102134
rect 65146 101898 65382 102134
rect 64826 66218 65062 66454
rect 65146 66218 65382 66454
rect 64826 65898 65062 66134
rect 65146 65898 65382 66134
rect 64826 30218 65062 30454
rect 65146 30218 65382 30454
rect 64826 29898 65062 30134
rect 65146 29898 65382 30134
rect 64826 -6342 65062 -6106
rect 65146 -6342 65382 -6106
rect 64826 -6662 65062 -6426
rect 65146 -6662 65382 -6426
rect 69326 711322 69562 711558
rect 69646 711322 69882 711558
rect 69326 711002 69562 711238
rect 69646 711002 69882 711238
rect 69326 682718 69562 682954
rect 69646 682718 69882 682954
rect 69326 682398 69562 682634
rect 69646 682398 69882 682634
rect 69326 646718 69562 646954
rect 69646 646718 69882 646954
rect 69326 646398 69562 646634
rect 69646 646398 69882 646634
rect 69326 610718 69562 610954
rect 69646 610718 69882 610954
rect 69326 610398 69562 610634
rect 69646 610398 69882 610634
rect 69326 574718 69562 574954
rect 69646 574718 69882 574954
rect 69326 574398 69562 574634
rect 69646 574398 69882 574634
rect 69326 538718 69562 538954
rect 69646 538718 69882 538954
rect 69326 538398 69562 538634
rect 69646 538398 69882 538634
rect 69326 502718 69562 502954
rect 69646 502718 69882 502954
rect 69326 502398 69562 502634
rect 69646 502398 69882 502634
rect 69326 466718 69562 466954
rect 69646 466718 69882 466954
rect 69326 466398 69562 466634
rect 69646 466398 69882 466634
rect 69326 430718 69562 430954
rect 69646 430718 69882 430954
rect 69326 430398 69562 430634
rect 69646 430398 69882 430634
rect 69326 394718 69562 394954
rect 69646 394718 69882 394954
rect 69326 394398 69562 394634
rect 69646 394398 69882 394634
rect 69326 358718 69562 358954
rect 69646 358718 69882 358954
rect 69326 358398 69562 358634
rect 69646 358398 69882 358634
rect 69326 322718 69562 322954
rect 69646 322718 69882 322954
rect 69326 322398 69562 322634
rect 69646 322398 69882 322634
rect 69326 286718 69562 286954
rect 69646 286718 69882 286954
rect 69326 286398 69562 286634
rect 69646 286398 69882 286634
rect 69326 250718 69562 250954
rect 69646 250718 69882 250954
rect 69326 250398 69562 250634
rect 69646 250398 69882 250634
rect 69326 214718 69562 214954
rect 69646 214718 69882 214954
rect 69326 214398 69562 214634
rect 69646 214398 69882 214634
rect 69326 178718 69562 178954
rect 69646 178718 69882 178954
rect 69326 178398 69562 178634
rect 69646 178398 69882 178634
rect 69326 142718 69562 142954
rect 69646 142718 69882 142954
rect 69326 142398 69562 142634
rect 69646 142398 69882 142634
rect 69326 106718 69562 106954
rect 69646 106718 69882 106954
rect 69326 106398 69562 106634
rect 69646 106398 69882 106634
rect 69326 70718 69562 70954
rect 69646 70718 69882 70954
rect 69326 70398 69562 70634
rect 69646 70398 69882 70634
rect 69326 34718 69562 34954
rect 69646 34718 69882 34954
rect 69326 34398 69562 34634
rect 69646 34398 69882 34634
rect 69326 -7302 69562 -7066
rect 69646 -7302 69882 -7066
rect 69326 -7622 69562 -7386
rect 69646 -7622 69882 -7386
rect 73826 704602 74062 704838
rect 74146 704602 74382 704838
rect 73826 704282 74062 704518
rect 74146 704282 74382 704518
rect 73826 687218 74062 687454
rect 74146 687218 74382 687454
rect 73826 686898 74062 687134
rect 74146 686898 74382 687134
rect 73826 651218 74062 651454
rect 74146 651218 74382 651454
rect 73826 650898 74062 651134
rect 74146 650898 74382 651134
rect 73826 615218 74062 615454
rect 74146 615218 74382 615454
rect 73826 614898 74062 615134
rect 74146 614898 74382 615134
rect 73826 579218 74062 579454
rect 74146 579218 74382 579454
rect 73826 578898 74062 579134
rect 74146 578898 74382 579134
rect 73826 543218 74062 543454
rect 74146 543218 74382 543454
rect 73826 542898 74062 543134
rect 74146 542898 74382 543134
rect 73826 507218 74062 507454
rect 74146 507218 74382 507454
rect 73826 506898 74062 507134
rect 74146 506898 74382 507134
rect 73826 471218 74062 471454
rect 74146 471218 74382 471454
rect 73826 470898 74062 471134
rect 74146 470898 74382 471134
rect 73826 435218 74062 435454
rect 74146 435218 74382 435454
rect 73826 434898 74062 435134
rect 74146 434898 74382 435134
rect 73826 399218 74062 399454
rect 74146 399218 74382 399454
rect 73826 398898 74062 399134
rect 74146 398898 74382 399134
rect 73826 363218 74062 363454
rect 74146 363218 74382 363454
rect 73826 362898 74062 363134
rect 74146 362898 74382 363134
rect 73826 327218 74062 327454
rect 74146 327218 74382 327454
rect 73826 326898 74062 327134
rect 74146 326898 74382 327134
rect 73826 291218 74062 291454
rect 74146 291218 74382 291454
rect 73826 290898 74062 291134
rect 74146 290898 74382 291134
rect 73826 255218 74062 255454
rect 74146 255218 74382 255454
rect 73826 254898 74062 255134
rect 74146 254898 74382 255134
rect 73826 219218 74062 219454
rect 74146 219218 74382 219454
rect 73826 218898 74062 219134
rect 74146 218898 74382 219134
rect 73826 183218 74062 183454
rect 74146 183218 74382 183454
rect 73826 182898 74062 183134
rect 74146 182898 74382 183134
rect 73826 147218 74062 147454
rect 74146 147218 74382 147454
rect 73826 146898 74062 147134
rect 74146 146898 74382 147134
rect 73826 111218 74062 111454
rect 74146 111218 74382 111454
rect 73826 110898 74062 111134
rect 74146 110898 74382 111134
rect 73826 75218 74062 75454
rect 74146 75218 74382 75454
rect 73826 74898 74062 75134
rect 74146 74898 74382 75134
rect 73826 39218 74062 39454
rect 74146 39218 74382 39454
rect 73826 38898 74062 39134
rect 74146 38898 74382 39134
rect 73826 3218 74062 3454
rect 74146 3218 74382 3454
rect 73826 2898 74062 3134
rect 74146 2898 74382 3134
rect 73826 -582 74062 -346
rect 74146 -582 74382 -346
rect 73826 -902 74062 -666
rect 74146 -902 74382 -666
rect 78326 705562 78562 705798
rect 78646 705562 78882 705798
rect 78326 705242 78562 705478
rect 78646 705242 78882 705478
rect 78326 691718 78562 691954
rect 78646 691718 78882 691954
rect 78326 691398 78562 691634
rect 78646 691398 78882 691634
rect 78326 655718 78562 655954
rect 78646 655718 78882 655954
rect 78326 655398 78562 655634
rect 78646 655398 78882 655634
rect 78326 619718 78562 619954
rect 78646 619718 78882 619954
rect 78326 619398 78562 619634
rect 78646 619398 78882 619634
rect 78326 583718 78562 583954
rect 78646 583718 78882 583954
rect 78326 583398 78562 583634
rect 78646 583398 78882 583634
rect 78326 547718 78562 547954
rect 78646 547718 78882 547954
rect 78326 547398 78562 547634
rect 78646 547398 78882 547634
rect 78326 511718 78562 511954
rect 78646 511718 78882 511954
rect 78326 511398 78562 511634
rect 78646 511398 78882 511634
rect 78326 475718 78562 475954
rect 78646 475718 78882 475954
rect 78326 475398 78562 475634
rect 78646 475398 78882 475634
rect 78326 439718 78562 439954
rect 78646 439718 78882 439954
rect 78326 439398 78562 439634
rect 78646 439398 78882 439634
rect 78326 403718 78562 403954
rect 78646 403718 78882 403954
rect 78326 403398 78562 403634
rect 78646 403398 78882 403634
rect 78326 367718 78562 367954
rect 78646 367718 78882 367954
rect 78326 367398 78562 367634
rect 78646 367398 78882 367634
rect 78326 331718 78562 331954
rect 78646 331718 78882 331954
rect 78326 331398 78562 331634
rect 78646 331398 78882 331634
rect 78326 295718 78562 295954
rect 78646 295718 78882 295954
rect 78326 295398 78562 295634
rect 78646 295398 78882 295634
rect 78326 259718 78562 259954
rect 78646 259718 78882 259954
rect 78326 259398 78562 259634
rect 78646 259398 78882 259634
rect 78326 223718 78562 223954
rect 78646 223718 78882 223954
rect 78326 223398 78562 223634
rect 78646 223398 78882 223634
rect 78326 187718 78562 187954
rect 78646 187718 78882 187954
rect 78326 187398 78562 187634
rect 78646 187398 78882 187634
rect 78326 151718 78562 151954
rect 78646 151718 78882 151954
rect 78326 151398 78562 151634
rect 78646 151398 78882 151634
rect 78326 115718 78562 115954
rect 78646 115718 78882 115954
rect 78326 115398 78562 115634
rect 78646 115398 78882 115634
rect 78326 79718 78562 79954
rect 78646 79718 78882 79954
rect 78326 79398 78562 79634
rect 78646 79398 78882 79634
rect 78326 43718 78562 43954
rect 78646 43718 78882 43954
rect 78326 43398 78562 43634
rect 78646 43398 78882 43634
rect 78326 7718 78562 7954
rect 78646 7718 78882 7954
rect 78326 7398 78562 7634
rect 78646 7398 78882 7634
rect 78326 -1542 78562 -1306
rect 78646 -1542 78882 -1306
rect 78326 -1862 78562 -1626
rect 78646 -1862 78882 -1626
rect 82826 706522 83062 706758
rect 83146 706522 83382 706758
rect 82826 706202 83062 706438
rect 83146 706202 83382 706438
rect 82826 696218 83062 696454
rect 83146 696218 83382 696454
rect 82826 695898 83062 696134
rect 83146 695898 83382 696134
rect 82826 660218 83062 660454
rect 83146 660218 83382 660454
rect 82826 659898 83062 660134
rect 83146 659898 83382 660134
rect 82826 624218 83062 624454
rect 83146 624218 83382 624454
rect 82826 623898 83062 624134
rect 83146 623898 83382 624134
rect 82826 588218 83062 588454
rect 83146 588218 83382 588454
rect 82826 587898 83062 588134
rect 83146 587898 83382 588134
rect 82826 552218 83062 552454
rect 83146 552218 83382 552454
rect 82826 551898 83062 552134
rect 83146 551898 83382 552134
rect 82826 516218 83062 516454
rect 83146 516218 83382 516454
rect 82826 515898 83062 516134
rect 83146 515898 83382 516134
rect 82826 480218 83062 480454
rect 83146 480218 83382 480454
rect 82826 479898 83062 480134
rect 83146 479898 83382 480134
rect 82826 444218 83062 444454
rect 83146 444218 83382 444454
rect 82826 443898 83062 444134
rect 83146 443898 83382 444134
rect 82826 408218 83062 408454
rect 83146 408218 83382 408454
rect 82826 407898 83062 408134
rect 83146 407898 83382 408134
rect 82826 372218 83062 372454
rect 83146 372218 83382 372454
rect 82826 371898 83062 372134
rect 83146 371898 83382 372134
rect 82826 336218 83062 336454
rect 83146 336218 83382 336454
rect 82826 335898 83062 336134
rect 83146 335898 83382 336134
rect 82826 300218 83062 300454
rect 83146 300218 83382 300454
rect 82826 299898 83062 300134
rect 83146 299898 83382 300134
rect 82826 264218 83062 264454
rect 83146 264218 83382 264454
rect 82826 263898 83062 264134
rect 83146 263898 83382 264134
rect 82826 228218 83062 228454
rect 83146 228218 83382 228454
rect 82826 227898 83062 228134
rect 83146 227898 83382 228134
rect 82826 192218 83062 192454
rect 83146 192218 83382 192454
rect 82826 191898 83062 192134
rect 83146 191898 83382 192134
rect 82826 156218 83062 156454
rect 83146 156218 83382 156454
rect 82826 155898 83062 156134
rect 83146 155898 83382 156134
rect 82826 120218 83062 120454
rect 83146 120218 83382 120454
rect 82826 119898 83062 120134
rect 83146 119898 83382 120134
rect 82826 84218 83062 84454
rect 83146 84218 83382 84454
rect 82826 83898 83062 84134
rect 83146 83898 83382 84134
rect 82826 48218 83062 48454
rect 83146 48218 83382 48454
rect 82826 47898 83062 48134
rect 83146 47898 83382 48134
rect 82826 12218 83062 12454
rect 83146 12218 83382 12454
rect 82826 11898 83062 12134
rect 83146 11898 83382 12134
rect 82826 -2502 83062 -2266
rect 83146 -2502 83382 -2266
rect 82826 -2822 83062 -2586
rect 83146 -2822 83382 -2586
rect 87326 707482 87562 707718
rect 87646 707482 87882 707718
rect 87326 707162 87562 707398
rect 87646 707162 87882 707398
rect 87326 700718 87562 700954
rect 87646 700718 87882 700954
rect 87326 700398 87562 700634
rect 87646 700398 87882 700634
rect 87326 664718 87562 664954
rect 87646 664718 87882 664954
rect 87326 664398 87562 664634
rect 87646 664398 87882 664634
rect 87326 628718 87562 628954
rect 87646 628718 87882 628954
rect 87326 628398 87562 628634
rect 87646 628398 87882 628634
rect 87326 592718 87562 592954
rect 87646 592718 87882 592954
rect 87326 592398 87562 592634
rect 87646 592398 87882 592634
rect 87326 556718 87562 556954
rect 87646 556718 87882 556954
rect 87326 556398 87562 556634
rect 87646 556398 87882 556634
rect 87326 520718 87562 520954
rect 87646 520718 87882 520954
rect 87326 520398 87562 520634
rect 87646 520398 87882 520634
rect 87326 484718 87562 484954
rect 87646 484718 87882 484954
rect 87326 484398 87562 484634
rect 87646 484398 87882 484634
rect 87326 448718 87562 448954
rect 87646 448718 87882 448954
rect 87326 448398 87562 448634
rect 87646 448398 87882 448634
rect 87326 412718 87562 412954
rect 87646 412718 87882 412954
rect 87326 412398 87562 412634
rect 87646 412398 87882 412634
rect 87326 376718 87562 376954
rect 87646 376718 87882 376954
rect 87326 376398 87562 376634
rect 87646 376398 87882 376634
rect 87326 340718 87562 340954
rect 87646 340718 87882 340954
rect 87326 340398 87562 340634
rect 87646 340398 87882 340634
rect 87326 304718 87562 304954
rect 87646 304718 87882 304954
rect 87326 304398 87562 304634
rect 87646 304398 87882 304634
rect 87326 268718 87562 268954
rect 87646 268718 87882 268954
rect 87326 268398 87562 268634
rect 87646 268398 87882 268634
rect 87326 232718 87562 232954
rect 87646 232718 87882 232954
rect 87326 232398 87562 232634
rect 87646 232398 87882 232634
rect 87326 196718 87562 196954
rect 87646 196718 87882 196954
rect 87326 196398 87562 196634
rect 87646 196398 87882 196634
rect 87326 160718 87562 160954
rect 87646 160718 87882 160954
rect 87326 160398 87562 160634
rect 87646 160398 87882 160634
rect 87326 124718 87562 124954
rect 87646 124718 87882 124954
rect 87326 124398 87562 124634
rect 87646 124398 87882 124634
rect 87326 88718 87562 88954
rect 87646 88718 87882 88954
rect 87326 88398 87562 88634
rect 87646 88398 87882 88634
rect 87326 52718 87562 52954
rect 87646 52718 87882 52954
rect 87326 52398 87562 52634
rect 87646 52398 87882 52634
rect 87326 16718 87562 16954
rect 87646 16718 87882 16954
rect 87326 16398 87562 16634
rect 87646 16398 87882 16634
rect 87326 -3462 87562 -3226
rect 87646 -3462 87882 -3226
rect 87326 -3782 87562 -3546
rect 87646 -3782 87882 -3546
rect 91826 708442 92062 708678
rect 92146 708442 92382 708678
rect 91826 708122 92062 708358
rect 92146 708122 92382 708358
rect 91826 669218 92062 669454
rect 92146 669218 92382 669454
rect 91826 668898 92062 669134
rect 92146 668898 92382 669134
rect 91826 633218 92062 633454
rect 92146 633218 92382 633454
rect 91826 632898 92062 633134
rect 92146 632898 92382 633134
rect 91826 597218 92062 597454
rect 92146 597218 92382 597454
rect 91826 596898 92062 597134
rect 92146 596898 92382 597134
rect 91826 561218 92062 561454
rect 92146 561218 92382 561454
rect 91826 560898 92062 561134
rect 92146 560898 92382 561134
rect 91826 525218 92062 525454
rect 92146 525218 92382 525454
rect 91826 524898 92062 525134
rect 92146 524898 92382 525134
rect 91826 489218 92062 489454
rect 92146 489218 92382 489454
rect 91826 488898 92062 489134
rect 92146 488898 92382 489134
rect 91826 453218 92062 453454
rect 92146 453218 92382 453454
rect 91826 452898 92062 453134
rect 92146 452898 92382 453134
rect 91826 417218 92062 417454
rect 92146 417218 92382 417454
rect 91826 416898 92062 417134
rect 92146 416898 92382 417134
rect 91826 381218 92062 381454
rect 92146 381218 92382 381454
rect 91826 380898 92062 381134
rect 92146 380898 92382 381134
rect 91826 345218 92062 345454
rect 92146 345218 92382 345454
rect 91826 344898 92062 345134
rect 92146 344898 92382 345134
rect 91826 309218 92062 309454
rect 92146 309218 92382 309454
rect 91826 308898 92062 309134
rect 92146 308898 92382 309134
rect 91826 273218 92062 273454
rect 92146 273218 92382 273454
rect 91826 272898 92062 273134
rect 92146 272898 92382 273134
rect 91826 237218 92062 237454
rect 92146 237218 92382 237454
rect 91826 236898 92062 237134
rect 92146 236898 92382 237134
rect 91826 201218 92062 201454
rect 92146 201218 92382 201454
rect 91826 200898 92062 201134
rect 92146 200898 92382 201134
rect 91826 165218 92062 165454
rect 92146 165218 92382 165454
rect 91826 164898 92062 165134
rect 92146 164898 92382 165134
rect 91826 129218 92062 129454
rect 92146 129218 92382 129454
rect 91826 128898 92062 129134
rect 92146 128898 92382 129134
rect 91826 93218 92062 93454
rect 92146 93218 92382 93454
rect 91826 92898 92062 93134
rect 92146 92898 92382 93134
rect 91826 57218 92062 57454
rect 92146 57218 92382 57454
rect 91826 56898 92062 57134
rect 92146 56898 92382 57134
rect 91826 21218 92062 21454
rect 92146 21218 92382 21454
rect 91826 20898 92062 21134
rect 92146 20898 92382 21134
rect 91826 -4422 92062 -4186
rect 92146 -4422 92382 -4186
rect 91826 -4742 92062 -4506
rect 92146 -4742 92382 -4506
rect 96326 709402 96562 709638
rect 96646 709402 96882 709638
rect 96326 709082 96562 709318
rect 96646 709082 96882 709318
rect 96326 673718 96562 673954
rect 96646 673718 96882 673954
rect 96326 673398 96562 673634
rect 96646 673398 96882 673634
rect 96326 637718 96562 637954
rect 96646 637718 96882 637954
rect 96326 637398 96562 637634
rect 96646 637398 96882 637634
rect 96326 601718 96562 601954
rect 96646 601718 96882 601954
rect 96326 601398 96562 601634
rect 96646 601398 96882 601634
rect 96326 565718 96562 565954
rect 96646 565718 96882 565954
rect 96326 565398 96562 565634
rect 96646 565398 96882 565634
rect 96326 529718 96562 529954
rect 96646 529718 96882 529954
rect 96326 529398 96562 529634
rect 96646 529398 96882 529634
rect 96326 493718 96562 493954
rect 96646 493718 96882 493954
rect 96326 493398 96562 493634
rect 96646 493398 96882 493634
rect 96326 457718 96562 457954
rect 96646 457718 96882 457954
rect 96326 457398 96562 457634
rect 96646 457398 96882 457634
rect 96326 421718 96562 421954
rect 96646 421718 96882 421954
rect 96326 421398 96562 421634
rect 96646 421398 96882 421634
rect 96326 385718 96562 385954
rect 96646 385718 96882 385954
rect 96326 385398 96562 385634
rect 96646 385398 96882 385634
rect 96326 349718 96562 349954
rect 96646 349718 96882 349954
rect 96326 349398 96562 349634
rect 96646 349398 96882 349634
rect 96326 313718 96562 313954
rect 96646 313718 96882 313954
rect 96326 313398 96562 313634
rect 96646 313398 96882 313634
rect 96326 277718 96562 277954
rect 96646 277718 96882 277954
rect 96326 277398 96562 277634
rect 96646 277398 96882 277634
rect 96326 241718 96562 241954
rect 96646 241718 96882 241954
rect 96326 241398 96562 241634
rect 96646 241398 96882 241634
rect 96326 205718 96562 205954
rect 96646 205718 96882 205954
rect 96326 205398 96562 205634
rect 96646 205398 96882 205634
rect 100826 710362 101062 710598
rect 101146 710362 101382 710598
rect 100826 710042 101062 710278
rect 101146 710042 101382 710278
rect 100826 678218 101062 678454
rect 101146 678218 101382 678454
rect 100826 677898 101062 678134
rect 101146 677898 101382 678134
rect 100826 642218 101062 642454
rect 101146 642218 101382 642454
rect 100826 641898 101062 642134
rect 101146 641898 101382 642134
rect 100826 606218 101062 606454
rect 101146 606218 101382 606454
rect 100826 605898 101062 606134
rect 101146 605898 101382 606134
rect 100826 570218 101062 570454
rect 101146 570218 101382 570454
rect 100826 569898 101062 570134
rect 101146 569898 101382 570134
rect 100826 534218 101062 534454
rect 101146 534218 101382 534454
rect 100826 533898 101062 534134
rect 101146 533898 101382 534134
rect 100826 498218 101062 498454
rect 101146 498218 101382 498454
rect 100826 497898 101062 498134
rect 101146 497898 101382 498134
rect 100826 462218 101062 462454
rect 101146 462218 101382 462454
rect 100826 461898 101062 462134
rect 101146 461898 101382 462134
rect 100826 426218 101062 426454
rect 101146 426218 101382 426454
rect 100826 425898 101062 426134
rect 101146 425898 101382 426134
rect 100826 390218 101062 390454
rect 101146 390218 101382 390454
rect 100826 389898 101062 390134
rect 101146 389898 101382 390134
rect 100826 354218 101062 354454
rect 101146 354218 101382 354454
rect 100826 353898 101062 354134
rect 101146 353898 101382 354134
rect 100826 318218 101062 318454
rect 101146 318218 101382 318454
rect 100826 317898 101062 318134
rect 101146 317898 101382 318134
rect 100826 282218 101062 282454
rect 101146 282218 101382 282454
rect 100826 281898 101062 282134
rect 101146 281898 101382 282134
rect 100826 246218 101062 246454
rect 101146 246218 101382 246454
rect 100826 245898 101062 246134
rect 101146 245898 101382 246134
rect 100826 210218 101062 210454
rect 101146 210218 101382 210454
rect 100826 209898 101062 210134
rect 101146 209898 101382 210134
rect 96326 169718 96562 169954
rect 96646 169718 96882 169954
rect 96326 169398 96562 169634
rect 96646 169398 96882 169634
rect 96326 133718 96562 133954
rect 96646 133718 96882 133954
rect 96326 133398 96562 133634
rect 96646 133398 96882 133634
rect 96326 97718 96562 97954
rect 96646 97718 96882 97954
rect 96326 97398 96562 97634
rect 96646 97398 96882 97634
rect 96326 61718 96562 61954
rect 96646 61718 96882 61954
rect 96326 61398 96562 61634
rect 96646 61398 96882 61634
rect 105326 711322 105562 711558
rect 105646 711322 105882 711558
rect 105326 711002 105562 711238
rect 105646 711002 105882 711238
rect 105326 682718 105562 682954
rect 105646 682718 105882 682954
rect 105326 682398 105562 682634
rect 105646 682398 105882 682634
rect 105326 646718 105562 646954
rect 105646 646718 105882 646954
rect 105326 646398 105562 646634
rect 105646 646398 105882 646634
rect 105326 610718 105562 610954
rect 105646 610718 105882 610954
rect 105326 610398 105562 610634
rect 105646 610398 105882 610634
rect 105326 574718 105562 574954
rect 105646 574718 105882 574954
rect 105326 574398 105562 574634
rect 105646 574398 105882 574634
rect 105326 538718 105562 538954
rect 105646 538718 105882 538954
rect 105326 538398 105562 538634
rect 105646 538398 105882 538634
rect 105326 502718 105562 502954
rect 105646 502718 105882 502954
rect 105326 502398 105562 502634
rect 105646 502398 105882 502634
rect 105326 466718 105562 466954
rect 105646 466718 105882 466954
rect 105326 466398 105562 466634
rect 105646 466398 105882 466634
rect 105326 430718 105562 430954
rect 105646 430718 105882 430954
rect 105326 430398 105562 430634
rect 105646 430398 105882 430634
rect 105326 394718 105562 394954
rect 105646 394718 105882 394954
rect 105326 394398 105562 394634
rect 105646 394398 105882 394634
rect 105326 358718 105562 358954
rect 105646 358718 105882 358954
rect 105326 358398 105562 358634
rect 105646 358398 105882 358634
rect 105326 322718 105562 322954
rect 105646 322718 105882 322954
rect 105326 322398 105562 322634
rect 105646 322398 105882 322634
rect 105326 286718 105562 286954
rect 105646 286718 105882 286954
rect 105326 286398 105562 286634
rect 105646 286398 105882 286634
rect 109826 704602 110062 704838
rect 110146 704602 110382 704838
rect 109826 704282 110062 704518
rect 110146 704282 110382 704518
rect 109826 687218 110062 687454
rect 110146 687218 110382 687454
rect 109826 686898 110062 687134
rect 110146 686898 110382 687134
rect 109826 651218 110062 651454
rect 110146 651218 110382 651454
rect 109826 650898 110062 651134
rect 110146 650898 110382 651134
rect 109826 615218 110062 615454
rect 110146 615218 110382 615454
rect 109826 614898 110062 615134
rect 110146 614898 110382 615134
rect 109826 579218 110062 579454
rect 110146 579218 110382 579454
rect 109826 578898 110062 579134
rect 110146 578898 110382 579134
rect 109826 543218 110062 543454
rect 110146 543218 110382 543454
rect 109826 542898 110062 543134
rect 110146 542898 110382 543134
rect 109826 507218 110062 507454
rect 110146 507218 110382 507454
rect 109826 506898 110062 507134
rect 110146 506898 110382 507134
rect 109826 471218 110062 471454
rect 110146 471218 110382 471454
rect 109826 470898 110062 471134
rect 110146 470898 110382 471134
rect 109826 435218 110062 435454
rect 110146 435218 110382 435454
rect 109826 434898 110062 435134
rect 110146 434898 110382 435134
rect 109826 399218 110062 399454
rect 110146 399218 110382 399454
rect 109826 398898 110062 399134
rect 110146 398898 110382 399134
rect 109826 363218 110062 363454
rect 110146 363218 110382 363454
rect 109826 362898 110062 363134
rect 110146 362898 110382 363134
rect 109826 327218 110062 327454
rect 110146 327218 110382 327454
rect 109826 326898 110062 327134
rect 110146 326898 110382 327134
rect 109826 291218 110062 291454
rect 110146 291218 110382 291454
rect 109826 290898 110062 291134
rect 110146 290898 110382 291134
rect 105326 250718 105562 250954
rect 105646 250718 105882 250954
rect 105326 250398 105562 250634
rect 105646 250398 105882 250634
rect 105326 214718 105562 214954
rect 105646 214718 105882 214954
rect 105326 214398 105562 214634
rect 105646 214398 105882 214634
rect 100826 174218 101062 174454
rect 101146 174218 101382 174454
rect 100826 173898 101062 174134
rect 101146 173898 101382 174134
rect 100826 138218 101062 138454
rect 101146 138218 101382 138454
rect 100826 137898 101062 138134
rect 101146 137898 101382 138134
rect 100826 102218 101062 102454
rect 101146 102218 101382 102454
rect 100826 101898 101062 102134
rect 101146 101898 101382 102134
rect 100826 66218 101062 66454
rect 101146 66218 101382 66454
rect 100826 65898 101062 66134
rect 101146 65898 101382 66134
rect 96326 25718 96562 25954
rect 96646 25718 96882 25954
rect 96326 25398 96562 25634
rect 96646 25398 96882 25634
rect 96326 -5382 96562 -5146
rect 96646 -5382 96882 -5146
rect 96326 -5702 96562 -5466
rect 96646 -5702 96882 -5466
rect 105326 178718 105562 178954
rect 105646 178718 105882 178954
rect 105326 178398 105562 178634
rect 105646 178398 105882 178634
rect 105326 142718 105562 142954
rect 105646 142718 105882 142954
rect 105326 142398 105562 142634
rect 105646 142398 105882 142634
rect 105326 106718 105562 106954
rect 105646 106718 105882 106954
rect 105326 106398 105562 106634
rect 105646 106398 105882 106634
rect 105326 70718 105562 70954
rect 105646 70718 105882 70954
rect 105326 70398 105562 70634
rect 105646 70398 105882 70634
rect 100826 30218 101062 30454
rect 101146 30218 101382 30454
rect 100826 29898 101062 30134
rect 101146 29898 101382 30134
rect 100826 -6342 101062 -6106
rect 101146 -6342 101382 -6106
rect 100826 -6662 101062 -6426
rect 101146 -6662 101382 -6426
rect 114326 705562 114562 705798
rect 114646 705562 114882 705798
rect 114326 705242 114562 705478
rect 114646 705242 114882 705478
rect 114326 691718 114562 691954
rect 114646 691718 114882 691954
rect 114326 691398 114562 691634
rect 114646 691398 114882 691634
rect 114326 655718 114562 655954
rect 114646 655718 114882 655954
rect 114326 655398 114562 655634
rect 114646 655398 114882 655634
rect 114326 619718 114562 619954
rect 114646 619718 114882 619954
rect 114326 619398 114562 619634
rect 114646 619398 114882 619634
rect 114326 583718 114562 583954
rect 114646 583718 114882 583954
rect 114326 583398 114562 583634
rect 114646 583398 114882 583634
rect 114326 547718 114562 547954
rect 114646 547718 114882 547954
rect 114326 547398 114562 547634
rect 114646 547398 114882 547634
rect 114326 511718 114562 511954
rect 114646 511718 114882 511954
rect 114326 511398 114562 511634
rect 114646 511398 114882 511634
rect 114326 475718 114562 475954
rect 114646 475718 114882 475954
rect 114326 475398 114562 475634
rect 114646 475398 114882 475634
rect 114326 439718 114562 439954
rect 114646 439718 114882 439954
rect 114326 439398 114562 439634
rect 114646 439398 114882 439634
rect 114326 403718 114562 403954
rect 114646 403718 114882 403954
rect 114326 403398 114562 403634
rect 114646 403398 114882 403634
rect 114326 367718 114562 367954
rect 114646 367718 114882 367954
rect 114326 367398 114562 367634
rect 114646 367398 114882 367634
rect 114326 331718 114562 331954
rect 114646 331718 114882 331954
rect 114326 331398 114562 331634
rect 114646 331398 114882 331634
rect 114326 295718 114562 295954
rect 114646 295718 114882 295954
rect 114326 295398 114562 295634
rect 114646 295398 114882 295634
rect 109826 255218 110062 255454
rect 110146 255218 110382 255454
rect 109826 254898 110062 255134
rect 110146 254898 110382 255134
rect 109826 219218 110062 219454
rect 110146 219218 110382 219454
rect 109826 218898 110062 219134
rect 110146 218898 110382 219134
rect 109826 183218 110062 183454
rect 110146 183218 110382 183454
rect 109826 182898 110062 183134
rect 110146 182898 110382 183134
rect 109826 147218 110062 147454
rect 110146 147218 110382 147454
rect 109826 146898 110062 147134
rect 110146 146898 110382 147134
rect 109826 111218 110062 111454
rect 110146 111218 110382 111454
rect 109826 110898 110062 111134
rect 110146 110898 110382 111134
rect 109826 75218 110062 75454
rect 110146 75218 110382 75454
rect 109826 74898 110062 75134
rect 110146 74898 110382 75134
rect 105326 34718 105562 34954
rect 105646 34718 105882 34954
rect 105326 34398 105562 34634
rect 105646 34398 105882 34634
rect 105326 -7302 105562 -7066
rect 105646 -7302 105882 -7066
rect 105326 -7622 105562 -7386
rect 105646 -7622 105882 -7386
rect 118826 706522 119062 706758
rect 119146 706522 119382 706758
rect 118826 706202 119062 706438
rect 119146 706202 119382 706438
rect 118826 696218 119062 696454
rect 119146 696218 119382 696454
rect 118826 695898 119062 696134
rect 119146 695898 119382 696134
rect 118826 660218 119062 660454
rect 119146 660218 119382 660454
rect 118826 659898 119062 660134
rect 119146 659898 119382 660134
rect 118826 624218 119062 624454
rect 119146 624218 119382 624454
rect 118826 623898 119062 624134
rect 119146 623898 119382 624134
rect 118826 588218 119062 588454
rect 119146 588218 119382 588454
rect 118826 587898 119062 588134
rect 119146 587898 119382 588134
rect 118826 552218 119062 552454
rect 119146 552218 119382 552454
rect 118826 551898 119062 552134
rect 119146 551898 119382 552134
rect 118826 516218 119062 516454
rect 119146 516218 119382 516454
rect 118826 515898 119062 516134
rect 119146 515898 119382 516134
rect 118826 480218 119062 480454
rect 119146 480218 119382 480454
rect 118826 479898 119062 480134
rect 119146 479898 119382 480134
rect 118826 444218 119062 444454
rect 119146 444218 119382 444454
rect 118826 443898 119062 444134
rect 119146 443898 119382 444134
rect 118826 408218 119062 408454
rect 119146 408218 119382 408454
rect 118826 407898 119062 408134
rect 119146 407898 119382 408134
rect 118826 372218 119062 372454
rect 119146 372218 119382 372454
rect 118826 371898 119062 372134
rect 119146 371898 119382 372134
rect 118826 336218 119062 336454
rect 119146 336218 119382 336454
rect 118826 335898 119062 336134
rect 119146 335898 119382 336134
rect 118826 300218 119062 300454
rect 119146 300218 119382 300454
rect 118826 299898 119062 300134
rect 119146 299898 119382 300134
rect 118826 264218 119062 264454
rect 119146 264218 119382 264454
rect 118826 263898 119062 264134
rect 119146 263898 119382 264134
rect 114326 259718 114562 259954
rect 114646 259718 114882 259954
rect 114326 259398 114562 259634
rect 114646 259398 114882 259634
rect 114326 223718 114562 223954
rect 114646 223718 114882 223954
rect 114326 223398 114562 223634
rect 114646 223398 114882 223634
rect 114326 187718 114562 187954
rect 114646 187718 114882 187954
rect 114326 187398 114562 187634
rect 114646 187398 114882 187634
rect 114326 151718 114562 151954
rect 114646 151718 114882 151954
rect 114326 151398 114562 151634
rect 114646 151398 114882 151634
rect 114326 115718 114562 115954
rect 114646 115718 114882 115954
rect 114326 115398 114562 115634
rect 114646 115398 114882 115634
rect 114326 79718 114562 79954
rect 114646 79718 114882 79954
rect 114326 79398 114562 79634
rect 114646 79398 114882 79634
rect 109826 39218 110062 39454
rect 110146 39218 110382 39454
rect 109826 38898 110062 39134
rect 110146 38898 110382 39134
rect 109826 3218 110062 3454
rect 110146 3218 110382 3454
rect 109826 2898 110062 3134
rect 110146 2898 110382 3134
rect 109826 -582 110062 -346
rect 110146 -582 110382 -346
rect 109826 -902 110062 -666
rect 110146 -902 110382 -666
rect 123326 707482 123562 707718
rect 123646 707482 123882 707718
rect 123326 707162 123562 707398
rect 123646 707162 123882 707398
rect 123326 700718 123562 700954
rect 123646 700718 123882 700954
rect 123326 700398 123562 700634
rect 123646 700398 123882 700634
rect 123326 664718 123562 664954
rect 123646 664718 123882 664954
rect 123326 664398 123562 664634
rect 123646 664398 123882 664634
rect 123326 628718 123562 628954
rect 123646 628718 123882 628954
rect 123326 628398 123562 628634
rect 123646 628398 123882 628634
rect 123326 592718 123562 592954
rect 123646 592718 123882 592954
rect 123326 592398 123562 592634
rect 123646 592398 123882 592634
rect 123326 556718 123562 556954
rect 123646 556718 123882 556954
rect 123326 556398 123562 556634
rect 123646 556398 123882 556634
rect 123326 520718 123562 520954
rect 123646 520718 123882 520954
rect 123326 520398 123562 520634
rect 123646 520398 123882 520634
rect 123326 484718 123562 484954
rect 123646 484718 123882 484954
rect 123326 484398 123562 484634
rect 123646 484398 123882 484634
rect 123326 448718 123562 448954
rect 123646 448718 123882 448954
rect 123326 448398 123562 448634
rect 123646 448398 123882 448634
rect 123326 412718 123562 412954
rect 123646 412718 123882 412954
rect 123326 412398 123562 412634
rect 123646 412398 123882 412634
rect 123326 376718 123562 376954
rect 123646 376718 123882 376954
rect 123326 376398 123562 376634
rect 123646 376398 123882 376634
rect 123326 340718 123562 340954
rect 123646 340718 123882 340954
rect 123326 340398 123562 340634
rect 123646 340398 123882 340634
rect 123326 304718 123562 304954
rect 123646 304718 123882 304954
rect 123326 304398 123562 304634
rect 123646 304398 123882 304634
rect 123326 268718 123562 268954
rect 123646 268718 123882 268954
rect 123326 268398 123562 268634
rect 123646 268398 123882 268634
rect 127826 708442 128062 708678
rect 128146 708442 128382 708678
rect 127826 708122 128062 708358
rect 128146 708122 128382 708358
rect 127826 669218 128062 669454
rect 128146 669218 128382 669454
rect 127826 668898 128062 669134
rect 128146 668898 128382 669134
rect 127826 633218 128062 633454
rect 128146 633218 128382 633454
rect 127826 632898 128062 633134
rect 128146 632898 128382 633134
rect 127826 597218 128062 597454
rect 128146 597218 128382 597454
rect 127826 596898 128062 597134
rect 128146 596898 128382 597134
rect 127826 561218 128062 561454
rect 128146 561218 128382 561454
rect 127826 560898 128062 561134
rect 128146 560898 128382 561134
rect 127826 525218 128062 525454
rect 128146 525218 128382 525454
rect 127826 524898 128062 525134
rect 128146 524898 128382 525134
rect 127826 489218 128062 489454
rect 128146 489218 128382 489454
rect 127826 488898 128062 489134
rect 128146 488898 128382 489134
rect 127826 453218 128062 453454
rect 128146 453218 128382 453454
rect 127826 452898 128062 453134
rect 128146 452898 128382 453134
rect 127826 417218 128062 417454
rect 128146 417218 128382 417454
rect 127826 416898 128062 417134
rect 128146 416898 128382 417134
rect 127826 381218 128062 381454
rect 128146 381218 128382 381454
rect 127826 380898 128062 381134
rect 128146 380898 128382 381134
rect 127826 345218 128062 345454
rect 128146 345218 128382 345454
rect 127826 344898 128062 345134
rect 128146 344898 128382 345134
rect 127826 309218 128062 309454
rect 128146 309218 128382 309454
rect 127826 308898 128062 309134
rect 128146 308898 128382 309134
rect 127826 273218 128062 273454
rect 128146 273218 128382 273454
rect 127826 272898 128062 273134
rect 128146 272898 128382 273134
rect 132326 709402 132562 709638
rect 132646 709402 132882 709638
rect 132326 709082 132562 709318
rect 132646 709082 132882 709318
rect 132326 673718 132562 673954
rect 132646 673718 132882 673954
rect 132326 673398 132562 673634
rect 132646 673398 132882 673634
rect 132326 637718 132562 637954
rect 132646 637718 132882 637954
rect 132326 637398 132562 637634
rect 132646 637398 132882 637634
rect 132326 601718 132562 601954
rect 132646 601718 132882 601954
rect 132326 601398 132562 601634
rect 132646 601398 132882 601634
rect 132326 565718 132562 565954
rect 132646 565718 132882 565954
rect 132326 565398 132562 565634
rect 132646 565398 132882 565634
rect 132326 529718 132562 529954
rect 132646 529718 132882 529954
rect 132326 529398 132562 529634
rect 132646 529398 132882 529634
rect 132326 493718 132562 493954
rect 132646 493718 132882 493954
rect 132326 493398 132562 493634
rect 132646 493398 132882 493634
rect 132326 457718 132562 457954
rect 132646 457718 132882 457954
rect 132326 457398 132562 457634
rect 132646 457398 132882 457634
rect 132326 421718 132562 421954
rect 132646 421718 132882 421954
rect 132326 421398 132562 421634
rect 132646 421398 132882 421634
rect 132326 385718 132562 385954
rect 132646 385718 132882 385954
rect 132326 385398 132562 385634
rect 132646 385398 132882 385634
rect 132326 349718 132562 349954
rect 132646 349718 132882 349954
rect 132326 349398 132562 349634
rect 132646 349398 132882 349634
rect 132326 313718 132562 313954
rect 132646 313718 132882 313954
rect 132326 313398 132562 313634
rect 132646 313398 132882 313634
rect 132326 277718 132562 277954
rect 132646 277718 132882 277954
rect 132326 277398 132562 277634
rect 132646 277398 132882 277634
rect 136826 710362 137062 710598
rect 137146 710362 137382 710598
rect 136826 710042 137062 710278
rect 137146 710042 137382 710278
rect 136826 678218 137062 678454
rect 137146 678218 137382 678454
rect 136826 677898 137062 678134
rect 137146 677898 137382 678134
rect 136826 642218 137062 642454
rect 137146 642218 137382 642454
rect 136826 641898 137062 642134
rect 137146 641898 137382 642134
rect 136826 606218 137062 606454
rect 137146 606218 137382 606454
rect 136826 605898 137062 606134
rect 137146 605898 137382 606134
rect 136826 570218 137062 570454
rect 137146 570218 137382 570454
rect 136826 569898 137062 570134
rect 137146 569898 137382 570134
rect 136826 534218 137062 534454
rect 137146 534218 137382 534454
rect 136826 533898 137062 534134
rect 137146 533898 137382 534134
rect 136826 498218 137062 498454
rect 137146 498218 137382 498454
rect 136826 497898 137062 498134
rect 137146 497898 137382 498134
rect 136826 462218 137062 462454
rect 137146 462218 137382 462454
rect 136826 461898 137062 462134
rect 137146 461898 137382 462134
rect 136826 426218 137062 426454
rect 137146 426218 137382 426454
rect 136826 425898 137062 426134
rect 137146 425898 137382 426134
rect 136826 390218 137062 390454
rect 137146 390218 137382 390454
rect 136826 389898 137062 390134
rect 137146 389898 137382 390134
rect 136826 354218 137062 354454
rect 137146 354218 137382 354454
rect 136826 353898 137062 354134
rect 137146 353898 137382 354134
rect 136826 318218 137062 318454
rect 137146 318218 137382 318454
rect 136826 317898 137062 318134
rect 137146 317898 137382 318134
rect 136826 282218 137062 282454
rect 137146 282218 137382 282454
rect 136826 281898 137062 282134
rect 137146 281898 137382 282134
rect 141326 711322 141562 711558
rect 141646 711322 141882 711558
rect 141326 711002 141562 711238
rect 141646 711002 141882 711238
rect 141326 682718 141562 682954
rect 141646 682718 141882 682954
rect 141326 682398 141562 682634
rect 141646 682398 141882 682634
rect 141326 646718 141562 646954
rect 141646 646718 141882 646954
rect 141326 646398 141562 646634
rect 141646 646398 141882 646634
rect 141326 610718 141562 610954
rect 141646 610718 141882 610954
rect 141326 610398 141562 610634
rect 141646 610398 141882 610634
rect 141326 574718 141562 574954
rect 141646 574718 141882 574954
rect 141326 574398 141562 574634
rect 141646 574398 141882 574634
rect 141326 538718 141562 538954
rect 141646 538718 141882 538954
rect 141326 538398 141562 538634
rect 141646 538398 141882 538634
rect 141326 502718 141562 502954
rect 141646 502718 141882 502954
rect 141326 502398 141562 502634
rect 141646 502398 141882 502634
rect 141326 466718 141562 466954
rect 141646 466718 141882 466954
rect 141326 466398 141562 466634
rect 141646 466398 141882 466634
rect 141326 430718 141562 430954
rect 141646 430718 141882 430954
rect 141326 430398 141562 430634
rect 141646 430398 141882 430634
rect 141326 394718 141562 394954
rect 141646 394718 141882 394954
rect 141326 394398 141562 394634
rect 141646 394398 141882 394634
rect 141326 358718 141562 358954
rect 141646 358718 141882 358954
rect 141326 358398 141562 358634
rect 141646 358398 141882 358634
rect 141326 322718 141562 322954
rect 141646 322718 141882 322954
rect 141326 322398 141562 322634
rect 141646 322398 141882 322634
rect 141326 286718 141562 286954
rect 141646 286718 141882 286954
rect 141326 286398 141562 286634
rect 141646 286398 141882 286634
rect 145826 704602 146062 704838
rect 146146 704602 146382 704838
rect 145826 704282 146062 704518
rect 146146 704282 146382 704518
rect 145826 687218 146062 687454
rect 146146 687218 146382 687454
rect 145826 686898 146062 687134
rect 146146 686898 146382 687134
rect 145826 651218 146062 651454
rect 146146 651218 146382 651454
rect 145826 650898 146062 651134
rect 146146 650898 146382 651134
rect 145826 615218 146062 615454
rect 146146 615218 146382 615454
rect 145826 614898 146062 615134
rect 146146 614898 146382 615134
rect 145826 579218 146062 579454
rect 146146 579218 146382 579454
rect 145826 578898 146062 579134
rect 146146 578898 146382 579134
rect 145826 543218 146062 543454
rect 146146 543218 146382 543454
rect 145826 542898 146062 543134
rect 146146 542898 146382 543134
rect 145826 507218 146062 507454
rect 146146 507218 146382 507454
rect 145826 506898 146062 507134
rect 146146 506898 146382 507134
rect 145826 471218 146062 471454
rect 146146 471218 146382 471454
rect 145826 470898 146062 471134
rect 146146 470898 146382 471134
rect 145826 435218 146062 435454
rect 146146 435218 146382 435454
rect 145826 434898 146062 435134
rect 146146 434898 146382 435134
rect 145826 399218 146062 399454
rect 146146 399218 146382 399454
rect 145826 398898 146062 399134
rect 146146 398898 146382 399134
rect 145826 363218 146062 363454
rect 146146 363218 146382 363454
rect 145826 362898 146062 363134
rect 146146 362898 146382 363134
rect 145826 327218 146062 327454
rect 146146 327218 146382 327454
rect 145826 326898 146062 327134
rect 146146 326898 146382 327134
rect 145826 291218 146062 291454
rect 146146 291218 146382 291454
rect 145826 290898 146062 291134
rect 146146 290898 146382 291134
rect 150326 705562 150562 705798
rect 150646 705562 150882 705798
rect 150326 705242 150562 705478
rect 150646 705242 150882 705478
rect 150326 691718 150562 691954
rect 150646 691718 150882 691954
rect 150326 691398 150562 691634
rect 150646 691398 150882 691634
rect 150326 655718 150562 655954
rect 150646 655718 150882 655954
rect 150326 655398 150562 655634
rect 150646 655398 150882 655634
rect 150326 619718 150562 619954
rect 150646 619718 150882 619954
rect 150326 619398 150562 619634
rect 150646 619398 150882 619634
rect 150326 583718 150562 583954
rect 150646 583718 150882 583954
rect 150326 583398 150562 583634
rect 150646 583398 150882 583634
rect 150326 547718 150562 547954
rect 150646 547718 150882 547954
rect 150326 547398 150562 547634
rect 150646 547398 150882 547634
rect 150326 511718 150562 511954
rect 150646 511718 150882 511954
rect 150326 511398 150562 511634
rect 150646 511398 150882 511634
rect 150326 475718 150562 475954
rect 150646 475718 150882 475954
rect 150326 475398 150562 475634
rect 150646 475398 150882 475634
rect 150326 439718 150562 439954
rect 150646 439718 150882 439954
rect 150326 439398 150562 439634
rect 150646 439398 150882 439634
rect 150326 403718 150562 403954
rect 150646 403718 150882 403954
rect 150326 403398 150562 403634
rect 150646 403398 150882 403634
rect 150326 367718 150562 367954
rect 150646 367718 150882 367954
rect 150326 367398 150562 367634
rect 150646 367398 150882 367634
rect 150326 331718 150562 331954
rect 150646 331718 150882 331954
rect 150326 331398 150562 331634
rect 150646 331398 150882 331634
rect 150326 295718 150562 295954
rect 150646 295718 150882 295954
rect 150326 295398 150562 295634
rect 150646 295398 150882 295634
rect 154826 706522 155062 706758
rect 155146 706522 155382 706758
rect 154826 706202 155062 706438
rect 155146 706202 155382 706438
rect 154826 696218 155062 696454
rect 155146 696218 155382 696454
rect 154826 695898 155062 696134
rect 155146 695898 155382 696134
rect 154826 660218 155062 660454
rect 155146 660218 155382 660454
rect 154826 659898 155062 660134
rect 155146 659898 155382 660134
rect 154826 624218 155062 624454
rect 155146 624218 155382 624454
rect 154826 623898 155062 624134
rect 155146 623898 155382 624134
rect 154826 588218 155062 588454
rect 155146 588218 155382 588454
rect 154826 587898 155062 588134
rect 155146 587898 155382 588134
rect 154826 552218 155062 552454
rect 155146 552218 155382 552454
rect 154826 551898 155062 552134
rect 155146 551898 155382 552134
rect 154826 516218 155062 516454
rect 155146 516218 155382 516454
rect 154826 515898 155062 516134
rect 155146 515898 155382 516134
rect 154826 480218 155062 480454
rect 155146 480218 155382 480454
rect 154826 479898 155062 480134
rect 155146 479898 155382 480134
rect 154826 444218 155062 444454
rect 155146 444218 155382 444454
rect 154826 443898 155062 444134
rect 155146 443898 155382 444134
rect 154826 408218 155062 408454
rect 155146 408218 155382 408454
rect 154826 407898 155062 408134
rect 155146 407898 155382 408134
rect 154826 372218 155062 372454
rect 155146 372218 155382 372454
rect 154826 371898 155062 372134
rect 155146 371898 155382 372134
rect 154826 336218 155062 336454
rect 155146 336218 155382 336454
rect 154826 335898 155062 336134
rect 155146 335898 155382 336134
rect 154826 300218 155062 300454
rect 155146 300218 155382 300454
rect 154826 299898 155062 300134
rect 155146 299898 155382 300134
rect 154826 264218 155062 264454
rect 155146 264218 155382 264454
rect 154826 263898 155062 264134
rect 155146 263898 155382 264134
rect 159326 707482 159562 707718
rect 159646 707482 159882 707718
rect 159326 707162 159562 707398
rect 159646 707162 159882 707398
rect 159326 700718 159562 700954
rect 159646 700718 159882 700954
rect 159326 700398 159562 700634
rect 159646 700398 159882 700634
rect 159326 664718 159562 664954
rect 159646 664718 159882 664954
rect 159326 664398 159562 664634
rect 159646 664398 159882 664634
rect 159326 628718 159562 628954
rect 159646 628718 159882 628954
rect 159326 628398 159562 628634
rect 159646 628398 159882 628634
rect 159326 592718 159562 592954
rect 159646 592718 159882 592954
rect 159326 592398 159562 592634
rect 159646 592398 159882 592634
rect 159326 556718 159562 556954
rect 159646 556718 159882 556954
rect 159326 556398 159562 556634
rect 159646 556398 159882 556634
rect 159326 520718 159562 520954
rect 159646 520718 159882 520954
rect 159326 520398 159562 520634
rect 159646 520398 159882 520634
rect 159326 484718 159562 484954
rect 159646 484718 159882 484954
rect 159326 484398 159562 484634
rect 159646 484398 159882 484634
rect 159326 448718 159562 448954
rect 159646 448718 159882 448954
rect 159326 448398 159562 448634
rect 159646 448398 159882 448634
rect 159326 412718 159562 412954
rect 159646 412718 159882 412954
rect 159326 412398 159562 412634
rect 159646 412398 159882 412634
rect 159326 376718 159562 376954
rect 159646 376718 159882 376954
rect 159326 376398 159562 376634
rect 159646 376398 159882 376634
rect 159326 340718 159562 340954
rect 159646 340718 159882 340954
rect 159326 340398 159562 340634
rect 159646 340398 159882 340634
rect 159326 304718 159562 304954
rect 159646 304718 159882 304954
rect 159326 304398 159562 304634
rect 159646 304398 159882 304634
rect 159326 268718 159562 268954
rect 159646 268718 159882 268954
rect 159326 268398 159562 268634
rect 159646 268398 159882 268634
rect 163826 708442 164062 708678
rect 164146 708442 164382 708678
rect 163826 708122 164062 708358
rect 164146 708122 164382 708358
rect 163826 669218 164062 669454
rect 164146 669218 164382 669454
rect 163826 668898 164062 669134
rect 164146 668898 164382 669134
rect 163826 633218 164062 633454
rect 164146 633218 164382 633454
rect 163826 632898 164062 633134
rect 164146 632898 164382 633134
rect 163826 597218 164062 597454
rect 164146 597218 164382 597454
rect 163826 596898 164062 597134
rect 164146 596898 164382 597134
rect 163826 561218 164062 561454
rect 164146 561218 164382 561454
rect 163826 560898 164062 561134
rect 164146 560898 164382 561134
rect 163826 525218 164062 525454
rect 164146 525218 164382 525454
rect 163826 524898 164062 525134
rect 164146 524898 164382 525134
rect 163826 489218 164062 489454
rect 164146 489218 164382 489454
rect 163826 488898 164062 489134
rect 164146 488898 164382 489134
rect 163826 453218 164062 453454
rect 164146 453218 164382 453454
rect 163826 452898 164062 453134
rect 164146 452898 164382 453134
rect 163826 417218 164062 417454
rect 164146 417218 164382 417454
rect 163826 416898 164062 417134
rect 164146 416898 164382 417134
rect 163826 381218 164062 381454
rect 164146 381218 164382 381454
rect 163826 380898 164062 381134
rect 164146 380898 164382 381134
rect 163826 345218 164062 345454
rect 164146 345218 164382 345454
rect 163826 344898 164062 345134
rect 164146 344898 164382 345134
rect 163826 309218 164062 309454
rect 164146 309218 164382 309454
rect 163826 308898 164062 309134
rect 164146 308898 164382 309134
rect 163826 273218 164062 273454
rect 164146 273218 164382 273454
rect 163826 272898 164062 273134
rect 164146 272898 164382 273134
rect 168326 709402 168562 709638
rect 168646 709402 168882 709638
rect 168326 709082 168562 709318
rect 168646 709082 168882 709318
rect 168326 673718 168562 673954
rect 168646 673718 168882 673954
rect 168326 673398 168562 673634
rect 168646 673398 168882 673634
rect 168326 637718 168562 637954
rect 168646 637718 168882 637954
rect 168326 637398 168562 637634
rect 168646 637398 168882 637634
rect 168326 601718 168562 601954
rect 168646 601718 168882 601954
rect 168326 601398 168562 601634
rect 168646 601398 168882 601634
rect 168326 565718 168562 565954
rect 168646 565718 168882 565954
rect 168326 565398 168562 565634
rect 168646 565398 168882 565634
rect 168326 529718 168562 529954
rect 168646 529718 168882 529954
rect 168326 529398 168562 529634
rect 168646 529398 168882 529634
rect 168326 493718 168562 493954
rect 168646 493718 168882 493954
rect 168326 493398 168562 493634
rect 168646 493398 168882 493634
rect 168326 457718 168562 457954
rect 168646 457718 168882 457954
rect 168326 457398 168562 457634
rect 168646 457398 168882 457634
rect 168326 421718 168562 421954
rect 168646 421718 168882 421954
rect 168326 421398 168562 421634
rect 168646 421398 168882 421634
rect 168326 385718 168562 385954
rect 168646 385718 168882 385954
rect 168326 385398 168562 385634
rect 168646 385398 168882 385634
rect 168326 349718 168562 349954
rect 168646 349718 168882 349954
rect 168326 349398 168562 349634
rect 168646 349398 168882 349634
rect 168326 313718 168562 313954
rect 168646 313718 168882 313954
rect 168326 313398 168562 313634
rect 168646 313398 168882 313634
rect 168326 277718 168562 277954
rect 168646 277718 168882 277954
rect 168326 277398 168562 277634
rect 168646 277398 168882 277634
rect 172826 710362 173062 710598
rect 173146 710362 173382 710598
rect 172826 710042 173062 710278
rect 173146 710042 173382 710278
rect 172826 678218 173062 678454
rect 173146 678218 173382 678454
rect 172826 677898 173062 678134
rect 173146 677898 173382 678134
rect 172826 642218 173062 642454
rect 173146 642218 173382 642454
rect 172826 641898 173062 642134
rect 173146 641898 173382 642134
rect 172826 606218 173062 606454
rect 173146 606218 173382 606454
rect 172826 605898 173062 606134
rect 173146 605898 173382 606134
rect 172826 570218 173062 570454
rect 173146 570218 173382 570454
rect 172826 569898 173062 570134
rect 173146 569898 173382 570134
rect 172826 534218 173062 534454
rect 173146 534218 173382 534454
rect 172826 533898 173062 534134
rect 173146 533898 173382 534134
rect 172826 498218 173062 498454
rect 173146 498218 173382 498454
rect 172826 497898 173062 498134
rect 173146 497898 173382 498134
rect 172826 462218 173062 462454
rect 173146 462218 173382 462454
rect 172826 461898 173062 462134
rect 173146 461898 173382 462134
rect 172826 426218 173062 426454
rect 173146 426218 173382 426454
rect 172826 425898 173062 426134
rect 173146 425898 173382 426134
rect 172826 390218 173062 390454
rect 173146 390218 173382 390454
rect 172826 389898 173062 390134
rect 173146 389898 173382 390134
rect 172826 354218 173062 354454
rect 173146 354218 173382 354454
rect 172826 353898 173062 354134
rect 173146 353898 173382 354134
rect 172826 318218 173062 318454
rect 173146 318218 173382 318454
rect 172826 317898 173062 318134
rect 173146 317898 173382 318134
rect 172826 282218 173062 282454
rect 173146 282218 173382 282454
rect 172826 281898 173062 282134
rect 173146 281898 173382 282134
rect 177326 711322 177562 711558
rect 177646 711322 177882 711558
rect 177326 711002 177562 711238
rect 177646 711002 177882 711238
rect 177326 682718 177562 682954
rect 177646 682718 177882 682954
rect 177326 682398 177562 682634
rect 177646 682398 177882 682634
rect 177326 646718 177562 646954
rect 177646 646718 177882 646954
rect 177326 646398 177562 646634
rect 177646 646398 177882 646634
rect 177326 610718 177562 610954
rect 177646 610718 177882 610954
rect 177326 610398 177562 610634
rect 177646 610398 177882 610634
rect 177326 574718 177562 574954
rect 177646 574718 177882 574954
rect 177326 574398 177562 574634
rect 177646 574398 177882 574634
rect 177326 538718 177562 538954
rect 177646 538718 177882 538954
rect 177326 538398 177562 538634
rect 177646 538398 177882 538634
rect 177326 502718 177562 502954
rect 177646 502718 177882 502954
rect 177326 502398 177562 502634
rect 177646 502398 177882 502634
rect 177326 466718 177562 466954
rect 177646 466718 177882 466954
rect 177326 466398 177562 466634
rect 177646 466398 177882 466634
rect 177326 430718 177562 430954
rect 177646 430718 177882 430954
rect 177326 430398 177562 430634
rect 177646 430398 177882 430634
rect 177326 394718 177562 394954
rect 177646 394718 177882 394954
rect 177326 394398 177562 394634
rect 177646 394398 177882 394634
rect 177326 358718 177562 358954
rect 177646 358718 177882 358954
rect 177326 358398 177562 358634
rect 177646 358398 177882 358634
rect 177326 322718 177562 322954
rect 177646 322718 177882 322954
rect 177326 322398 177562 322634
rect 177646 322398 177882 322634
rect 177326 286718 177562 286954
rect 177646 286718 177882 286954
rect 177326 286398 177562 286634
rect 177646 286398 177882 286634
rect 181826 704602 182062 704838
rect 182146 704602 182382 704838
rect 181826 704282 182062 704518
rect 182146 704282 182382 704518
rect 181826 687218 182062 687454
rect 182146 687218 182382 687454
rect 181826 686898 182062 687134
rect 182146 686898 182382 687134
rect 181826 651218 182062 651454
rect 182146 651218 182382 651454
rect 181826 650898 182062 651134
rect 182146 650898 182382 651134
rect 181826 615218 182062 615454
rect 182146 615218 182382 615454
rect 181826 614898 182062 615134
rect 182146 614898 182382 615134
rect 181826 579218 182062 579454
rect 182146 579218 182382 579454
rect 181826 578898 182062 579134
rect 182146 578898 182382 579134
rect 181826 543218 182062 543454
rect 182146 543218 182382 543454
rect 181826 542898 182062 543134
rect 182146 542898 182382 543134
rect 181826 507218 182062 507454
rect 182146 507218 182382 507454
rect 181826 506898 182062 507134
rect 182146 506898 182382 507134
rect 181826 471218 182062 471454
rect 182146 471218 182382 471454
rect 181826 470898 182062 471134
rect 182146 470898 182382 471134
rect 181826 435218 182062 435454
rect 182146 435218 182382 435454
rect 181826 434898 182062 435134
rect 182146 434898 182382 435134
rect 181826 399218 182062 399454
rect 182146 399218 182382 399454
rect 181826 398898 182062 399134
rect 182146 398898 182382 399134
rect 181826 363218 182062 363454
rect 182146 363218 182382 363454
rect 181826 362898 182062 363134
rect 182146 362898 182382 363134
rect 181826 327218 182062 327454
rect 182146 327218 182382 327454
rect 181826 326898 182062 327134
rect 182146 326898 182382 327134
rect 181826 291218 182062 291454
rect 182146 291218 182382 291454
rect 181826 290898 182062 291134
rect 182146 290898 182382 291134
rect 186326 705562 186562 705798
rect 186646 705562 186882 705798
rect 186326 705242 186562 705478
rect 186646 705242 186882 705478
rect 186326 691718 186562 691954
rect 186646 691718 186882 691954
rect 186326 691398 186562 691634
rect 186646 691398 186882 691634
rect 186326 655718 186562 655954
rect 186646 655718 186882 655954
rect 186326 655398 186562 655634
rect 186646 655398 186882 655634
rect 186326 619718 186562 619954
rect 186646 619718 186882 619954
rect 186326 619398 186562 619634
rect 186646 619398 186882 619634
rect 186326 583718 186562 583954
rect 186646 583718 186882 583954
rect 186326 583398 186562 583634
rect 186646 583398 186882 583634
rect 186326 547718 186562 547954
rect 186646 547718 186882 547954
rect 186326 547398 186562 547634
rect 186646 547398 186882 547634
rect 186326 511718 186562 511954
rect 186646 511718 186882 511954
rect 186326 511398 186562 511634
rect 186646 511398 186882 511634
rect 186326 475718 186562 475954
rect 186646 475718 186882 475954
rect 186326 475398 186562 475634
rect 186646 475398 186882 475634
rect 186326 439718 186562 439954
rect 186646 439718 186882 439954
rect 186326 439398 186562 439634
rect 186646 439398 186882 439634
rect 186326 403718 186562 403954
rect 186646 403718 186882 403954
rect 186326 403398 186562 403634
rect 186646 403398 186882 403634
rect 186326 367718 186562 367954
rect 186646 367718 186882 367954
rect 186326 367398 186562 367634
rect 186646 367398 186882 367634
rect 186326 331718 186562 331954
rect 186646 331718 186882 331954
rect 186326 331398 186562 331634
rect 186646 331398 186882 331634
rect 186326 295718 186562 295954
rect 186646 295718 186882 295954
rect 186326 295398 186562 295634
rect 186646 295398 186882 295634
rect 190826 706522 191062 706758
rect 191146 706522 191382 706758
rect 190826 706202 191062 706438
rect 191146 706202 191382 706438
rect 190826 696218 191062 696454
rect 191146 696218 191382 696454
rect 190826 695898 191062 696134
rect 191146 695898 191382 696134
rect 190826 660218 191062 660454
rect 191146 660218 191382 660454
rect 190826 659898 191062 660134
rect 191146 659898 191382 660134
rect 190826 624218 191062 624454
rect 191146 624218 191382 624454
rect 190826 623898 191062 624134
rect 191146 623898 191382 624134
rect 190826 588218 191062 588454
rect 191146 588218 191382 588454
rect 190826 587898 191062 588134
rect 191146 587898 191382 588134
rect 190826 552218 191062 552454
rect 191146 552218 191382 552454
rect 190826 551898 191062 552134
rect 191146 551898 191382 552134
rect 190826 516218 191062 516454
rect 191146 516218 191382 516454
rect 190826 515898 191062 516134
rect 191146 515898 191382 516134
rect 190826 480218 191062 480454
rect 191146 480218 191382 480454
rect 190826 479898 191062 480134
rect 191146 479898 191382 480134
rect 190826 444218 191062 444454
rect 191146 444218 191382 444454
rect 190826 443898 191062 444134
rect 191146 443898 191382 444134
rect 190826 408218 191062 408454
rect 191146 408218 191382 408454
rect 190826 407898 191062 408134
rect 191146 407898 191382 408134
rect 190826 372218 191062 372454
rect 191146 372218 191382 372454
rect 190826 371898 191062 372134
rect 191146 371898 191382 372134
rect 190826 336218 191062 336454
rect 191146 336218 191382 336454
rect 190826 335898 191062 336134
rect 191146 335898 191382 336134
rect 190826 300218 191062 300454
rect 191146 300218 191382 300454
rect 190826 299898 191062 300134
rect 191146 299898 191382 300134
rect 118826 192218 119062 192454
rect 119146 192218 119382 192454
rect 118826 191898 119062 192134
rect 119146 191898 119382 192134
rect 118826 156218 119062 156454
rect 119146 156218 119382 156454
rect 118826 155898 119062 156134
rect 119146 155898 119382 156134
rect 118826 48218 119062 48454
rect 119146 48218 119382 48454
rect 118826 47898 119062 48134
rect 119146 47898 119382 48134
rect 114326 43718 114562 43954
rect 114646 43718 114882 43954
rect 114326 43398 114562 43634
rect 114646 43398 114882 43634
rect 114326 7718 114562 7954
rect 114646 7718 114882 7954
rect 114326 7398 114562 7634
rect 114646 7398 114882 7634
rect 114326 -1542 114562 -1306
rect 114646 -1542 114882 -1306
rect 114326 -1862 114562 -1626
rect 114646 -1862 114882 -1626
rect 123326 196718 123562 196954
rect 123646 196718 123882 196954
rect 123326 196398 123562 196634
rect 123646 196398 123882 196634
rect 123326 160718 123562 160954
rect 123646 160718 123882 160954
rect 123326 160398 123562 160634
rect 123646 160398 123882 160634
rect 124250 255218 124486 255454
rect 124250 254898 124486 255134
rect 154970 255218 155206 255454
rect 154970 254898 155206 255134
rect 185690 255218 185926 255454
rect 185690 254898 185926 255134
rect 139610 223718 139846 223954
rect 139610 223398 139846 223634
rect 170330 223718 170566 223954
rect 170330 223398 170566 223634
rect 124250 219218 124486 219454
rect 124250 218898 124486 219134
rect 154970 219218 155206 219454
rect 154970 218898 155206 219134
rect 185690 219218 185926 219454
rect 185690 218898 185926 219134
rect 141326 178718 141562 178954
rect 141646 178718 141882 178954
rect 141326 178398 141562 178634
rect 141646 178398 141882 178634
rect 145826 183218 146062 183454
rect 146146 183218 146382 183454
rect 145826 182898 146062 183134
rect 146146 182898 146382 183134
rect 145826 147218 146062 147454
rect 146146 147218 146382 147454
rect 145826 146898 146062 147134
rect 146146 146898 146382 147134
rect 141326 142718 141562 142954
rect 141646 142718 141882 142954
rect 141326 142398 141562 142634
rect 141646 142398 141882 142634
rect 150326 187718 150562 187954
rect 150646 187718 150882 187954
rect 150326 187398 150562 187634
rect 150646 187398 150882 187634
rect 154826 192218 155062 192454
rect 155146 192218 155382 192454
rect 154826 191898 155062 192134
rect 155146 191898 155382 192134
rect 150326 151718 150562 151954
rect 150646 151718 150882 151954
rect 150326 151398 150562 151634
rect 150646 151398 150882 151634
rect 154826 156218 155062 156454
rect 155146 156218 155382 156454
rect 154826 155898 155062 156134
rect 155146 155898 155382 156134
rect 159326 196718 159562 196954
rect 159646 196718 159882 196954
rect 159326 196398 159562 196634
rect 159646 196398 159882 196634
rect 159326 160718 159562 160954
rect 159646 160718 159882 160954
rect 159326 160398 159562 160634
rect 159646 160398 159882 160634
rect 177326 178718 177562 178954
rect 177646 178718 177882 178954
rect 177326 178398 177562 178634
rect 177646 178398 177882 178634
rect 177326 142718 177562 142954
rect 177646 142718 177882 142954
rect 177326 142398 177562 142634
rect 177646 142398 177882 142634
rect 181826 183218 182062 183454
rect 182146 183218 182382 183454
rect 181826 182898 182062 183134
rect 182146 182898 182382 183134
rect 181826 147218 182062 147454
rect 182146 147218 182382 147454
rect 181826 146898 182062 147134
rect 182146 146898 182382 147134
rect 186326 187718 186562 187954
rect 186646 187718 186882 187954
rect 186326 187398 186562 187634
rect 186646 187398 186882 187634
rect 186326 151718 186562 151954
rect 186646 151718 186882 151954
rect 186326 151398 186562 151634
rect 186646 151398 186882 151634
rect 139610 115718 139846 115954
rect 139610 115398 139846 115634
rect 170330 115718 170566 115954
rect 170330 115398 170566 115634
rect 124250 111218 124486 111454
rect 124250 110898 124486 111134
rect 154970 111218 155206 111454
rect 154970 110898 155206 111134
rect 185690 111218 185926 111454
rect 185690 110898 185926 111134
rect 123326 52718 123562 52954
rect 123646 52718 123882 52954
rect 123326 52398 123562 52634
rect 123646 52398 123882 52634
rect 118826 12218 119062 12454
rect 119146 12218 119382 12454
rect 118826 11898 119062 12134
rect 119146 11898 119382 12134
rect 118826 -2502 119062 -2266
rect 119146 -2502 119382 -2266
rect 118826 -2822 119062 -2586
rect 119146 -2822 119382 -2586
rect 123326 16718 123562 16954
rect 123646 16718 123882 16954
rect 123326 16398 123562 16634
rect 123646 16398 123882 16634
rect 123326 -3462 123562 -3226
rect 123646 -3462 123882 -3226
rect 123326 -3782 123562 -3546
rect 123646 -3782 123882 -3546
rect 127826 57218 128062 57454
rect 128146 57218 128382 57454
rect 127826 56898 128062 57134
rect 128146 56898 128382 57134
rect 127826 21218 128062 21454
rect 128146 21218 128382 21454
rect 127826 20898 128062 21134
rect 128146 20898 128382 21134
rect 127826 -4422 128062 -4186
rect 128146 -4422 128382 -4186
rect 127826 -4742 128062 -4506
rect 128146 -4742 128382 -4506
rect 132326 61718 132562 61954
rect 132646 61718 132882 61954
rect 132326 61398 132562 61634
rect 132646 61398 132882 61634
rect 136826 66218 137062 66454
rect 137146 66218 137382 66454
rect 136826 65898 137062 66134
rect 137146 65898 137382 66134
rect 132326 25718 132562 25954
rect 132646 25718 132882 25954
rect 132326 25398 132562 25634
rect 132646 25398 132882 25634
rect 132326 -5382 132562 -5146
rect 132646 -5382 132882 -5146
rect 132326 -5702 132562 -5466
rect 132646 -5702 132882 -5466
rect 141326 70718 141562 70954
rect 141646 70718 141882 70954
rect 141326 70398 141562 70634
rect 141646 70398 141882 70634
rect 136826 30218 137062 30454
rect 137146 30218 137382 30454
rect 136826 29898 137062 30134
rect 137146 29898 137382 30134
rect 136826 -6342 137062 -6106
rect 137146 -6342 137382 -6106
rect 136826 -6662 137062 -6426
rect 137146 -6662 137382 -6426
rect 141326 34718 141562 34954
rect 141646 34718 141882 34954
rect 141326 34398 141562 34634
rect 141646 34398 141882 34634
rect 145826 75218 146062 75454
rect 146146 75218 146382 75454
rect 145826 74898 146062 75134
rect 146146 74898 146382 75134
rect 145826 39218 146062 39454
rect 146146 39218 146382 39454
rect 145826 38898 146062 39134
rect 146146 38898 146382 39134
rect 141326 -7302 141562 -7066
rect 141646 -7302 141882 -7066
rect 141326 -7622 141562 -7386
rect 141646 -7622 141882 -7386
rect 150326 43718 150562 43954
rect 150646 43718 150882 43954
rect 150326 43398 150562 43634
rect 150646 43398 150882 43634
rect 145826 3218 146062 3454
rect 146146 3218 146382 3454
rect 145826 2898 146062 3134
rect 146146 2898 146382 3134
rect 145826 -582 146062 -346
rect 146146 -582 146382 -346
rect 145826 -902 146062 -666
rect 146146 -902 146382 -666
rect 154826 48218 155062 48454
rect 155146 48218 155382 48454
rect 154826 47898 155062 48134
rect 155146 47898 155382 48134
rect 150326 7718 150562 7954
rect 150646 7718 150882 7954
rect 150326 7398 150562 7634
rect 150646 7398 150882 7634
rect 150326 -1542 150562 -1306
rect 150646 -1542 150882 -1306
rect 150326 -1862 150562 -1626
rect 150646 -1862 150882 -1626
rect 159326 52718 159562 52954
rect 159646 52718 159882 52954
rect 159326 52398 159562 52634
rect 159646 52398 159882 52634
rect 154826 12218 155062 12454
rect 155146 12218 155382 12454
rect 154826 11898 155062 12134
rect 155146 11898 155382 12134
rect 154826 -2502 155062 -2266
rect 155146 -2502 155382 -2266
rect 154826 -2822 155062 -2586
rect 155146 -2822 155382 -2586
rect 163826 57218 164062 57454
rect 164146 57218 164382 57454
rect 163826 56898 164062 57134
rect 164146 56898 164382 57134
rect 159326 16718 159562 16954
rect 159646 16718 159882 16954
rect 159326 16398 159562 16634
rect 159646 16398 159882 16634
rect 159326 -3462 159562 -3226
rect 159646 -3462 159882 -3226
rect 159326 -3782 159562 -3546
rect 159646 -3782 159882 -3546
rect 168326 61718 168562 61954
rect 168646 61718 168882 61954
rect 168326 61398 168562 61634
rect 168646 61398 168882 61634
rect 163826 21218 164062 21454
rect 164146 21218 164382 21454
rect 163826 20898 164062 21134
rect 164146 20898 164382 21134
rect 163826 -4422 164062 -4186
rect 164146 -4422 164382 -4186
rect 163826 -4742 164062 -4506
rect 164146 -4742 164382 -4506
rect 172826 66218 173062 66454
rect 173146 66218 173382 66454
rect 172826 65898 173062 66134
rect 173146 65898 173382 66134
rect 168326 25718 168562 25954
rect 168646 25718 168882 25954
rect 168326 25398 168562 25634
rect 168646 25398 168882 25634
rect 168326 -5382 168562 -5146
rect 168646 -5382 168882 -5146
rect 168326 -5702 168562 -5466
rect 168646 -5702 168882 -5466
rect 177326 70718 177562 70954
rect 177646 70718 177882 70954
rect 177326 70398 177562 70634
rect 177646 70398 177882 70634
rect 172826 30218 173062 30454
rect 173146 30218 173382 30454
rect 172826 29898 173062 30134
rect 173146 29898 173382 30134
rect 172826 -6342 173062 -6106
rect 173146 -6342 173382 -6106
rect 172826 -6662 173062 -6426
rect 173146 -6662 173382 -6426
rect 177326 34718 177562 34954
rect 177646 34718 177882 34954
rect 177326 34398 177562 34634
rect 177646 34398 177882 34634
rect 177326 -7302 177562 -7066
rect 177646 -7302 177882 -7066
rect 177326 -7622 177562 -7386
rect 177646 -7622 177882 -7386
rect 181826 75218 182062 75454
rect 182146 75218 182382 75454
rect 181826 74898 182062 75134
rect 182146 74898 182382 75134
rect 181826 39218 182062 39454
rect 182146 39218 182382 39454
rect 181826 38898 182062 39134
rect 182146 38898 182382 39134
rect 181826 3218 182062 3454
rect 182146 3218 182382 3454
rect 181826 2898 182062 3134
rect 182146 2898 182382 3134
rect 181826 -582 182062 -346
rect 182146 -582 182382 -346
rect 181826 -902 182062 -666
rect 182146 -902 182382 -666
rect 195326 707482 195562 707718
rect 195646 707482 195882 707718
rect 195326 707162 195562 707398
rect 195646 707162 195882 707398
rect 195326 700718 195562 700954
rect 195646 700718 195882 700954
rect 195326 700398 195562 700634
rect 195646 700398 195882 700634
rect 195326 664718 195562 664954
rect 195646 664718 195882 664954
rect 195326 664398 195562 664634
rect 195646 664398 195882 664634
rect 195326 628718 195562 628954
rect 195646 628718 195882 628954
rect 195326 628398 195562 628634
rect 195646 628398 195882 628634
rect 195326 592718 195562 592954
rect 195646 592718 195882 592954
rect 195326 592398 195562 592634
rect 195646 592398 195882 592634
rect 195326 556718 195562 556954
rect 195646 556718 195882 556954
rect 195326 556398 195562 556634
rect 195646 556398 195882 556634
rect 195326 520718 195562 520954
rect 195646 520718 195882 520954
rect 195326 520398 195562 520634
rect 195646 520398 195882 520634
rect 195326 484718 195562 484954
rect 195646 484718 195882 484954
rect 195326 484398 195562 484634
rect 195646 484398 195882 484634
rect 195326 448718 195562 448954
rect 195646 448718 195882 448954
rect 195326 448398 195562 448634
rect 195646 448398 195882 448634
rect 195326 412718 195562 412954
rect 195646 412718 195882 412954
rect 195326 412398 195562 412634
rect 195646 412398 195882 412634
rect 195326 376718 195562 376954
rect 195646 376718 195882 376954
rect 195326 376398 195562 376634
rect 195646 376398 195882 376634
rect 195326 340718 195562 340954
rect 195646 340718 195882 340954
rect 195326 340398 195562 340634
rect 195646 340398 195882 340634
rect 195326 304718 195562 304954
rect 195646 304718 195882 304954
rect 195326 304398 195562 304634
rect 195646 304398 195882 304634
rect 195326 268718 195562 268954
rect 195646 268718 195882 268954
rect 195326 268398 195562 268634
rect 195646 268398 195882 268634
rect 190826 264218 191062 264454
rect 191146 264218 191382 264454
rect 190826 263898 191062 264134
rect 191146 263898 191382 264134
rect 190826 192218 191062 192454
rect 191146 192218 191382 192454
rect 190826 191898 191062 192134
rect 191146 191898 191382 192134
rect 190826 156218 191062 156454
rect 191146 156218 191382 156454
rect 190826 155898 191062 156134
rect 191146 155898 191382 156134
rect 186326 43718 186562 43954
rect 186646 43718 186882 43954
rect 186326 43398 186562 43634
rect 186646 43398 186882 43634
rect 186326 7718 186562 7954
rect 186646 7718 186882 7954
rect 186326 7398 186562 7634
rect 186646 7398 186882 7634
rect 186326 -1542 186562 -1306
rect 186646 -1542 186882 -1306
rect 186326 -1862 186562 -1626
rect 186646 -1862 186882 -1626
rect 199826 708442 200062 708678
rect 200146 708442 200382 708678
rect 199826 708122 200062 708358
rect 200146 708122 200382 708358
rect 199826 669218 200062 669454
rect 200146 669218 200382 669454
rect 199826 668898 200062 669134
rect 200146 668898 200382 669134
rect 199826 633218 200062 633454
rect 200146 633218 200382 633454
rect 199826 632898 200062 633134
rect 200146 632898 200382 633134
rect 199826 597218 200062 597454
rect 200146 597218 200382 597454
rect 199826 596898 200062 597134
rect 200146 596898 200382 597134
rect 199826 561218 200062 561454
rect 200146 561218 200382 561454
rect 199826 560898 200062 561134
rect 200146 560898 200382 561134
rect 199826 525218 200062 525454
rect 200146 525218 200382 525454
rect 199826 524898 200062 525134
rect 200146 524898 200382 525134
rect 199826 489218 200062 489454
rect 200146 489218 200382 489454
rect 199826 488898 200062 489134
rect 200146 488898 200382 489134
rect 199826 453218 200062 453454
rect 200146 453218 200382 453454
rect 199826 452898 200062 453134
rect 200146 452898 200382 453134
rect 199826 417218 200062 417454
rect 200146 417218 200382 417454
rect 199826 416898 200062 417134
rect 200146 416898 200382 417134
rect 199826 381218 200062 381454
rect 200146 381218 200382 381454
rect 199826 380898 200062 381134
rect 200146 380898 200382 381134
rect 199826 345218 200062 345454
rect 200146 345218 200382 345454
rect 199826 344898 200062 345134
rect 200146 344898 200382 345134
rect 199826 309218 200062 309454
rect 200146 309218 200382 309454
rect 199826 308898 200062 309134
rect 200146 308898 200382 309134
rect 199826 273218 200062 273454
rect 200146 273218 200382 273454
rect 199826 272898 200062 273134
rect 200146 272898 200382 273134
rect 195326 232718 195562 232954
rect 195646 232718 195882 232954
rect 195326 232398 195562 232634
rect 195646 232398 195882 232634
rect 195326 196718 195562 196954
rect 195646 196718 195882 196954
rect 195326 196398 195562 196634
rect 195646 196398 195882 196634
rect 195326 160718 195562 160954
rect 195646 160718 195882 160954
rect 195326 160398 195562 160634
rect 195646 160398 195882 160634
rect 195326 124718 195562 124954
rect 195646 124718 195882 124954
rect 195326 124398 195562 124634
rect 195646 124398 195882 124634
rect 195326 88718 195562 88954
rect 195646 88718 195882 88954
rect 195326 88398 195562 88634
rect 195646 88398 195882 88634
rect 199826 237218 200062 237454
rect 200146 237218 200382 237454
rect 199826 236898 200062 237134
rect 200146 236898 200382 237134
rect 199826 201218 200062 201454
rect 200146 201218 200382 201454
rect 199826 200898 200062 201134
rect 200146 200898 200382 201134
rect 195326 52718 195562 52954
rect 195646 52718 195882 52954
rect 195326 52398 195562 52634
rect 195646 52398 195882 52634
rect 190826 48218 191062 48454
rect 191146 48218 191382 48454
rect 190826 47898 191062 48134
rect 191146 47898 191382 48134
rect 190826 12218 191062 12454
rect 191146 12218 191382 12454
rect 190826 11898 191062 12134
rect 191146 11898 191382 12134
rect 190826 -2502 191062 -2266
rect 191146 -2502 191382 -2266
rect 190826 -2822 191062 -2586
rect 191146 -2822 191382 -2586
rect 204326 709402 204562 709638
rect 204646 709402 204882 709638
rect 204326 709082 204562 709318
rect 204646 709082 204882 709318
rect 204326 673718 204562 673954
rect 204646 673718 204882 673954
rect 204326 673398 204562 673634
rect 204646 673398 204882 673634
rect 204326 637718 204562 637954
rect 204646 637718 204882 637954
rect 204326 637398 204562 637634
rect 204646 637398 204882 637634
rect 204326 601718 204562 601954
rect 204646 601718 204882 601954
rect 204326 601398 204562 601634
rect 204646 601398 204882 601634
rect 204326 565718 204562 565954
rect 204646 565718 204882 565954
rect 204326 565398 204562 565634
rect 204646 565398 204882 565634
rect 204326 529718 204562 529954
rect 204646 529718 204882 529954
rect 204326 529398 204562 529634
rect 204646 529398 204882 529634
rect 204326 493718 204562 493954
rect 204646 493718 204882 493954
rect 204326 493398 204562 493634
rect 204646 493398 204882 493634
rect 204326 457718 204562 457954
rect 204646 457718 204882 457954
rect 204326 457398 204562 457634
rect 204646 457398 204882 457634
rect 204326 421718 204562 421954
rect 204646 421718 204882 421954
rect 204326 421398 204562 421634
rect 204646 421398 204882 421634
rect 204326 385718 204562 385954
rect 204646 385718 204882 385954
rect 204326 385398 204562 385634
rect 204646 385398 204882 385634
rect 204326 349718 204562 349954
rect 204646 349718 204882 349954
rect 204326 349398 204562 349634
rect 204646 349398 204882 349634
rect 204326 313718 204562 313954
rect 204646 313718 204882 313954
rect 204326 313398 204562 313634
rect 204646 313398 204882 313634
rect 204326 277718 204562 277954
rect 204646 277718 204882 277954
rect 204326 277398 204562 277634
rect 204646 277398 204882 277634
rect 204326 241718 204562 241954
rect 204646 241718 204882 241954
rect 204326 241398 204562 241634
rect 204646 241398 204882 241634
rect 204326 205718 204562 205954
rect 204646 205718 204882 205954
rect 204326 205398 204562 205634
rect 204646 205398 204882 205634
rect 199826 165218 200062 165454
rect 200146 165218 200382 165454
rect 199826 164898 200062 165134
rect 200146 164898 200382 165134
rect 199826 129218 200062 129454
rect 200146 129218 200382 129454
rect 199826 128898 200062 129134
rect 200146 128898 200382 129134
rect 199826 93218 200062 93454
rect 200146 93218 200382 93454
rect 199826 92898 200062 93134
rect 200146 92898 200382 93134
rect 199826 57218 200062 57454
rect 200146 57218 200382 57454
rect 199826 56898 200062 57134
rect 200146 56898 200382 57134
rect 195326 16718 195562 16954
rect 195646 16718 195882 16954
rect 195326 16398 195562 16634
rect 195646 16398 195882 16634
rect 195326 -3462 195562 -3226
rect 195646 -3462 195882 -3226
rect 195326 -3782 195562 -3546
rect 195646 -3782 195882 -3546
rect 208826 710362 209062 710598
rect 209146 710362 209382 710598
rect 208826 710042 209062 710278
rect 209146 710042 209382 710278
rect 208826 678218 209062 678454
rect 209146 678218 209382 678454
rect 208826 677898 209062 678134
rect 209146 677898 209382 678134
rect 208826 642218 209062 642454
rect 209146 642218 209382 642454
rect 208826 641898 209062 642134
rect 209146 641898 209382 642134
rect 208826 606218 209062 606454
rect 209146 606218 209382 606454
rect 208826 605898 209062 606134
rect 209146 605898 209382 606134
rect 208826 570218 209062 570454
rect 209146 570218 209382 570454
rect 208826 569898 209062 570134
rect 209146 569898 209382 570134
rect 208826 534218 209062 534454
rect 209146 534218 209382 534454
rect 208826 533898 209062 534134
rect 209146 533898 209382 534134
rect 208826 498218 209062 498454
rect 209146 498218 209382 498454
rect 208826 497898 209062 498134
rect 209146 497898 209382 498134
rect 208826 462218 209062 462454
rect 209146 462218 209382 462454
rect 208826 461898 209062 462134
rect 209146 461898 209382 462134
rect 208826 426218 209062 426454
rect 209146 426218 209382 426454
rect 208826 425898 209062 426134
rect 209146 425898 209382 426134
rect 208826 390218 209062 390454
rect 209146 390218 209382 390454
rect 208826 389898 209062 390134
rect 209146 389898 209382 390134
rect 208826 354218 209062 354454
rect 209146 354218 209382 354454
rect 208826 353898 209062 354134
rect 209146 353898 209382 354134
rect 208826 318218 209062 318454
rect 209146 318218 209382 318454
rect 208826 317898 209062 318134
rect 209146 317898 209382 318134
rect 208826 282218 209062 282454
rect 209146 282218 209382 282454
rect 208826 281898 209062 282134
rect 209146 281898 209382 282134
rect 208826 246218 209062 246454
rect 209146 246218 209382 246454
rect 208826 245898 209062 246134
rect 209146 245898 209382 246134
rect 208826 210218 209062 210454
rect 209146 210218 209382 210454
rect 208826 209898 209062 210134
rect 209146 209898 209382 210134
rect 204326 169718 204562 169954
rect 204646 169718 204882 169954
rect 204326 169398 204562 169634
rect 204646 169398 204882 169634
rect 204326 133718 204562 133954
rect 204646 133718 204882 133954
rect 204326 133398 204562 133634
rect 204646 133398 204882 133634
rect 204326 97718 204562 97954
rect 204646 97718 204882 97954
rect 204326 97398 204562 97634
rect 204646 97398 204882 97634
rect 213326 711322 213562 711558
rect 213646 711322 213882 711558
rect 213326 711002 213562 711238
rect 213646 711002 213882 711238
rect 213326 682718 213562 682954
rect 213646 682718 213882 682954
rect 213326 682398 213562 682634
rect 213646 682398 213882 682634
rect 213326 646718 213562 646954
rect 213646 646718 213882 646954
rect 213326 646398 213562 646634
rect 213646 646398 213882 646634
rect 213326 610718 213562 610954
rect 213646 610718 213882 610954
rect 213326 610398 213562 610634
rect 213646 610398 213882 610634
rect 213326 574718 213562 574954
rect 213646 574718 213882 574954
rect 213326 574398 213562 574634
rect 213646 574398 213882 574634
rect 213326 538718 213562 538954
rect 213646 538718 213882 538954
rect 213326 538398 213562 538634
rect 213646 538398 213882 538634
rect 213326 502718 213562 502954
rect 213646 502718 213882 502954
rect 213326 502398 213562 502634
rect 213646 502398 213882 502634
rect 213326 466718 213562 466954
rect 213646 466718 213882 466954
rect 213326 466398 213562 466634
rect 213646 466398 213882 466634
rect 213326 430718 213562 430954
rect 213646 430718 213882 430954
rect 213326 430398 213562 430634
rect 213646 430398 213882 430634
rect 213326 394718 213562 394954
rect 213646 394718 213882 394954
rect 213326 394398 213562 394634
rect 213646 394398 213882 394634
rect 213326 358718 213562 358954
rect 213646 358718 213882 358954
rect 213326 358398 213562 358634
rect 213646 358398 213882 358634
rect 213326 322718 213562 322954
rect 213646 322718 213882 322954
rect 213326 322398 213562 322634
rect 213646 322398 213882 322634
rect 213326 286718 213562 286954
rect 213646 286718 213882 286954
rect 213326 286398 213562 286634
rect 213646 286398 213882 286634
rect 213326 250718 213562 250954
rect 213646 250718 213882 250954
rect 213326 250398 213562 250634
rect 213646 250398 213882 250634
rect 213326 214718 213562 214954
rect 213646 214718 213882 214954
rect 213326 214398 213562 214634
rect 213646 214398 213882 214634
rect 208826 174218 209062 174454
rect 209146 174218 209382 174454
rect 208826 173898 209062 174134
rect 209146 173898 209382 174134
rect 204326 61718 204562 61954
rect 204646 61718 204882 61954
rect 204326 61398 204562 61634
rect 204646 61398 204882 61634
rect 199826 21218 200062 21454
rect 200146 21218 200382 21454
rect 199826 20898 200062 21134
rect 200146 20898 200382 21134
rect 199826 -4422 200062 -4186
rect 200146 -4422 200382 -4186
rect 199826 -4742 200062 -4506
rect 200146 -4742 200382 -4506
rect 208826 138218 209062 138454
rect 209146 138218 209382 138454
rect 208826 137898 209062 138134
rect 209146 137898 209382 138134
rect 208826 102218 209062 102454
rect 209146 102218 209382 102454
rect 208826 101898 209062 102134
rect 209146 101898 209382 102134
rect 208826 66218 209062 66454
rect 209146 66218 209382 66454
rect 208826 65898 209062 66134
rect 209146 65898 209382 66134
rect 204326 25718 204562 25954
rect 204646 25718 204882 25954
rect 204326 25398 204562 25634
rect 204646 25398 204882 25634
rect 204326 -5382 204562 -5146
rect 204646 -5382 204882 -5146
rect 204326 -5702 204562 -5466
rect 204646 -5702 204882 -5466
rect 213326 178718 213562 178954
rect 213646 178718 213882 178954
rect 213326 178398 213562 178634
rect 213646 178398 213882 178634
rect 213326 142718 213562 142954
rect 213646 142718 213882 142954
rect 213326 142398 213562 142634
rect 213646 142398 213882 142634
rect 213326 106718 213562 106954
rect 213646 106718 213882 106954
rect 213326 106398 213562 106634
rect 213646 106398 213882 106634
rect 213326 70718 213562 70954
rect 213646 70718 213882 70954
rect 213326 70398 213562 70634
rect 213646 70398 213882 70634
rect 208826 30218 209062 30454
rect 209146 30218 209382 30454
rect 208826 29898 209062 30134
rect 209146 29898 209382 30134
rect 208826 -6342 209062 -6106
rect 209146 -6342 209382 -6106
rect 208826 -6662 209062 -6426
rect 209146 -6662 209382 -6426
rect 213326 34718 213562 34954
rect 213646 34718 213882 34954
rect 213326 34398 213562 34634
rect 213646 34398 213882 34634
rect 213326 -7302 213562 -7066
rect 213646 -7302 213882 -7066
rect 213326 -7622 213562 -7386
rect 213646 -7622 213882 -7386
rect 217826 704602 218062 704838
rect 218146 704602 218382 704838
rect 217826 704282 218062 704518
rect 218146 704282 218382 704518
rect 217826 687218 218062 687454
rect 218146 687218 218382 687454
rect 217826 686898 218062 687134
rect 218146 686898 218382 687134
rect 217826 651218 218062 651454
rect 218146 651218 218382 651454
rect 217826 650898 218062 651134
rect 218146 650898 218382 651134
rect 217826 615218 218062 615454
rect 218146 615218 218382 615454
rect 217826 614898 218062 615134
rect 218146 614898 218382 615134
rect 217826 579218 218062 579454
rect 218146 579218 218382 579454
rect 217826 578898 218062 579134
rect 218146 578898 218382 579134
rect 217826 543218 218062 543454
rect 218146 543218 218382 543454
rect 217826 542898 218062 543134
rect 218146 542898 218382 543134
rect 217826 507218 218062 507454
rect 218146 507218 218382 507454
rect 217826 506898 218062 507134
rect 218146 506898 218382 507134
rect 217826 471218 218062 471454
rect 218146 471218 218382 471454
rect 217826 470898 218062 471134
rect 218146 470898 218382 471134
rect 217826 435218 218062 435454
rect 218146 435218 218382 435454
rect 217826 434898 218062 435134
rect 218146 434898 218382 435134
rect 217826 399218 218062 399454
rect 218146 399218 218382 399454
rect 217826 398898 218062 399134
rect 218146 398898 218382 399134
rect 217826 363218 218062 363454
rect 218146 363218 218382 363454
rect 217826 362898 218062 363134
rect 218146 362898 218382 363134
rect 217826 327218 218062 327454
rect 218146 327218 218382 327454
rect 217826 326898 218062 327134
rect 218146 326898 218382 327134
rect 217826 291218 218062 291454
rect 218146 291218 218382 291454
rect 217826 290898 218062 291134
rect 218146 290898 218382 291134
rect 217826 255218 218062 255454
rect 218146 255218 218382 255454
rect 217826 254898 218062 255134
rect 218146 254898 218382 255134
rect 217826 219218 218062 219454
rect 218146 219218 218382 219454
rect 217826 218898 218062 219134
rect 218146 218898 218382 219134
rect 217826 183218 218062 183454
rect 218146 183218 218382 183454
rect 217826 182898 218062 183134
rect 218146 182898 218382 183134
rect 217826 147218 218062 147454
rect 218146 147218 218382 147454
rect 217826 146898 218062 147134
rect 218146 146898 218382 147134
rect 217826 111218 218062 111454
rect 218146 111218 218382 111454
rect 217826 110898 218062 111134
rect 218146 110898 218382 111134
rect 217826 75218 218062 75454
rect 218146 75218 218382 75454
rect 217826 74898 218062 75134
rect 218146 74898 218382 75134
rect 217826 39218 218062 39454
rect 218146 39218 218382 39454
rect 217826 38898 218062 39134
rect 218146 38898 218382 39134
rect 217826 3218 218062 3454
rect 218146 3218 218382 3454
rect 217826 2898 218062 3134
rect 218146 2898 218382 3134
rect 217826 -582 218062 -346
rect 218146 -582 218382 -346
rect 217826 -902 218062 -666
rect 218146 -902 218382 -666
rect 222326 705562 222562 705798
rect 222646 705562 222882 705798
rect 222326 705242 222562 705478
rect 222646 705242 222882 705478
rect 222326 691718 222562 691954
rect 222646 691718 222882 691954
rect 222326 691398 222562 691634
rect 222646 691398 222882 691634
rect 222326 655718 222562 655954
rect 222646 655718 222882 655954
rect 222326 655398 222562 655634
rect 222646 655398 222882 655634
rect 222326 619718 222562 619954
rect 222646 619718 222882 619954
rect 222326 619398 222562 619634
rect 222646 619398 222882 619634
rect 222326 583718 222562 583954
rect 222646 583718 222882 583954
rect 222326 583398 222562 583634
rect 222646 583398 222882 583634
rect 222326 547718 222562 547954
rect 222646 547718 222882 547954
rect 222326 547398 222562 547634
rect 222646 547398 222882 547634
rect 222326 511718 222562 511954
rect 222646 511718 222882 511954
rect 222326 511398 222562 511634
rect 222646 511398 222882 511634
rect 222326 475718 222562 475954
rect 222646 475718 222882 475954
rect 222326 475398 222562 475634
rect 222646 475398 222882 475634
rect 222326 439718 222562 439954
rect 222646 439718 222882 439954
rect 222326 439398 222562 439634
rect 222646 439398 222882 439634
rect 222326 403718 222562 403954
rect 222646 403718 222882 403954
rect 222326 403398 222562 403634
rect 222646 403398 222882 403634
rect 222326 367718 222562 367954
rect 222646 367718 222882 367954
rect 222326 367398 222562 367634
rect 222646 367398 222882 367634
rect 222326 331718 222562 331954
rect 222646 331718 222882 331954
rect 222326 331398 222562 331634
rect 222646 331398 222882 331634
rect 222326 295718 222562 295954
rect 222646 295718 222882 295954
rect 222326 295398 222562 295634
rect 222646 295398 222882 295634
rect 222326 259718 222562 259954
rect 222646 259718 222882 259954
rect 222326 259398 222562 259634
rect 222646 259398 222882 259634
rect 222326 223718 222562 223954
rect 222646 223718 222882 223954
rect 222326 223398 222562 223634
rect 222646 223398 222882 223634
rect 222326 187718 222562 187954
rect 222646 187718 222882 187954
rect 222326 187398 222562 187634
rect 222646 187398 222882 187634
rect 222326 151718 222562 151954
rect 222646 151718 222882 151954
rect 222326 151398 222562 151634
rect 222646 151398 222882 151634
rect 222326 115718 222562 115954
rect 222646 115718 222882 115954
rect 222326 115398 222562 115634
rect 222646 115398 222882 115634
rect 222326 79718 222562 79954
rect 222646 79718 222882 79954
rect 222326 79398 222562 79634
rect 222646 79398 222882 79634
rect 222326 43718 222562 43954
rect 222646 43718 222882 43954
rect 222326 43398 222562 43634
rect 222646 43398 222882 43634
rect 222326 7718 222562 7954
rect 222646 7718 222882 7954
rect 222326 7398 222562 7634
rect 222646 7398 222882 7634
rect 222326 -1542 222562 -1306
rect 222646 -1542 222882 -1306
rect 222326 -1862 222562 -1626
rect 222646 -1862 222882 -1626
rect 226826 706522 227062 706758
rect 227146 706522 227382 706758
rect 226826 706202 227062 706438
rect 227146 706202 227382 706438
rect 226826 696218 227062 696454
rect 227146 696218 227382 696454
rect 226826 695898 227062 696134
rect 227146 695898 227382 696134
rect 226826 660218 227062 660454
rect 227146 660218 227382 660454
rect 226826 659898 227062 660134
rect 227146 659898 227382 660134
rect 226826 624218 227062 624454
rect 227146 624218 227382 624454
rect 226826 623898 227062 624134
rect 227146 623898 227382 624134
rect 226826 588218 227062 588454
rect 227146 588218 227382 588454
rect 226826 587898 227062 588134
rect 227146 587898 227382 588134
rect 226826 552218 227062 552454
rect 227146 552218 227382 552454
rect 226826 551898 227062 552134
rect 227146 551898 227382 552134
rect 226826 516218 227062 516454
rect 227146 516218 227382 516454
rect 226826 515898 227062 516134
rect 227146 515898 227382 516134
rect 226826 480218 227062 480454
rect 227146 480218 227382 480454
rect 226826 479898 227062 480134
rect 227146 479898 227382 480134
rect 226826 444218 227062 444454
rect 227146 444218 227382 444454
rect 226826 443898 227062 444134
rect 227146 443898 227382 444134
rect 226826 408218 227062 408454
rect 227146 408218 227382 408454
rect 226826 407898 227062 408134
rect 227146 407898 227382 408134
rect 226826 372218 227062 372454
rect 227146 372218 227382 372454
rect 226826 371898 227062 372134
rect 227146 371898 227382 372134
rect 226826 336218 227062 336454
rect 227146 336218 227382 336454
rect 226826 335898 227062 336134
rect 227146 335898 227382 336134
rect 226826 300218 227062 300454
rect 227146 300218 227382 300454
rect 226826 299898 227062 300134
rect 227146 299898 227382 300134
rect 226826 264218 227062 264454
rect 227146 264218 227382 264454
rect 226826 263898 227062 264134
rect 227146 263898 227382 264134
rect 226826 228218 227062 228454
rect 227146 228218 227382 228454
rect 226826 227898 227062 228134
rect 227146 227898 227382 228134
rect 226826 192218 227062 192454
rect 227146 192218 227382 192454
rect 226826 191898 227062 192134
rect 227146 191898 227382 192134
rect 226826 156218 227062 156454
rect 227146 156218 227382 156454
rect 226826 155898 227062 156134
rect 227146 155898 227382 156134
rect 226826 120218 227062 120454
rect 227146 120218 227382 120454
rect 226826 119898 227062 120134
rect 227146 119898 227382 120134
rect 226826 84218 227062 84454
rect 227146 84218 227382 84454
rect 226826 83898 227062 84134
rect 227146 83898 227382 84134
rect 226826 48218 227062 48454
rect 227146 48218 227382 48454
rect 226826 47898 227062 48134
rect 227146 47898 227382 48134
rect 226826 12218 227062 12454
rect 227146 12218 227382 12454
rect 226826 11898 227062 12134
rect 227146 11898 227382 12134
rect 226826 -2502 227062 -2266
rect 227146 -2502 227382 -2266
rect 226826 -2822 227062 -2586
rect 227146 -2822 227382 -2586
rect 231326 707482 231562 707718
rect 231646 707482 231882 707718
rect 231326 707162 231562 707398
rect 231646 707162 231882 707398
rect 231326 700718 231562 700954
rect 231646 700718 231882 700954
rect 231326 700398 231562 700634
rect 231646 700398 231882 700634
rect 231326 664718 231562 664954
rect 231646 664718 231882 664954
rect 231326 664398 231562 664634
rect 231646 664398 231882 664634
rect 231326 628718 231562 628954
rect 231646 628718 231882 628954
rect 231326 628398 231562 628634
rect 231646 628398 231882 628634
rect 231326 592718 231562 592954
rect 231646 592718 231882 592954
rect 231326 592398 231562 592634
rect 231646 592398 231882 592634
rect 231326 556718 231562 556954
rect 231646 556718 231882 556954
rect 231326 556398 231562 556634
rect 231646 556398 231882 556634
rect 231326 520718 231562 520954
rect 231646 520718 231882 520954
rect 231326 520398 231562 520634
rect 231646 520398 231882 520634
rect 231326 484718 231562 484954
rect 231646 484718 231882 484954
rect 231326 484398 231562 484634
rect 231646 484398 231882 484634
rect 231326 448718 231562 448954
rect 231646 448718 231882 448954
rect 231326 448398 231562 448634
rect 231646 448398 231882 448634
rect 231326 412718 231562 412954
rect 231646 412718 231882 412954
rect 231326 412398 231562 412634
rect 231646 412398 231882 412634
rect 231326 376718 231562 376954
rect 231646 376718 231882 376954
rect 231326 376398 231562 376634
rect 231646 376398 231882 376634
rect 231326 340718 231562 340954
rect 231646 340718 231882 340954
rect 231326 340398 231562 340634
rect 231646 340398 231882 340634
rect 231326 304718 231562 304954
rect 231646 304718 231882 304954
rect 231326 304398 231562 304634
rect 231646 304398 231882 304634
rect 231326 268718 231562 268954
rect 231646 268718 231882 268954
rect 231326 268398 231562 268634
rect 231646 268398 231882 268634
rect 231326 232718 231562 232954
rect 231646 232718 231882 232954
rect 231326 232398 231562 232634
rect 231646 232398 231882 232634
rect 231326 196718 231562 196954
rect 231646 196718 231882 196954
rect 231326 196398 231562 196634
rect 231646 196398 231882 196634
rect 231326 160718 231562 160954
rect 231646 160718 231882 160954
rect 231326 160398 231562 160634
rect 231646 160398 231882 160634
rect 231326 124718 231562 124954
rect 231646 124718 231882 124954
rect 231326 124398 231562 124634
rect 231646 124398 231882 124634
rect 231326 88718 231562 88954
rect 231646 88718 231882 88954
rect 231326 88398 231562 88634
rect 231646 88398 231882 88634
rect 231326 52718 231562 52954
rect 231646 52718 231882 52954
rect 231326 52398 231562 52634
rect 231646 52398 231882 52634
rect 231326 16718 231562 16954
rect 231646 16718 231882 16954
rect 231326 16398 231562 16634
rect 231646 16398 231882 16634
rect 231326 -3462 231562 -3226
rect 231646 -3462 231882 -3226
rect 231326 -3782 231562 -3546
rect 231646 -3782 231882 -3546
rect 235826 708442 236062 708678
rect 236146 708442 236382 708678
rect 235826 708122 236062 708358
rect 236146 708122 236382 708358
rect 235826 669218 236062 669454
rect 236146 669218 236382 669454
rect 235826 668898 236062 669134
rect 236146 668898 236382 669134
rect 235826 633218 236062 633454
rect 236146 633218 236382 633454
rect 235826 632898 236062 633134
rect 236146 632898 236382 633134
rect 235826 597218 236062 597454
rect 236146 597218 236382 597454
rect 235826 596898 236062 597134
rect 236146 596898 236382 597134
rect 235826 561218 236062 561454
rect 236146 561218 236382 561454
rect 235826 560898 236062 561134
rect 236146 560898 236382 561134
rect 235826 525218 236062 525454
rect 236146 525218 236382 525454
rect 235826 524898 236062 525134
rect 236146 524898 236382 525134
rect 235826 489218 236062 489454
rect 236146 489218 236382 489454
rect 235826 488898 236062 489134
rect 236146 488898 236382 489134
rect 235826 453218 236062 453454
rect 236146 453218 236382 453454
rect 235826 452898 236062 453134
rect 236146 452898 236382 453134
rect 235826 417218 236062 417454
rect 236146 417218 236382 417454
rect 235826 416898 236062 417134
rect 236146 416898 236382 417134
rect 235826 381218 236062 381454
rect 236146 381218 236382 381454
rect 235826 380898 236062 381134
rect 236146 380898 236382 381134
rect 235826 345218 236062 345454
rect 236146 345218 236382 345454
rect 235826 344898 236062 345134
rect 236146 344898 236382 345134
rect 235826 309218 236062 309454
rect 236146 309218 236382 309454
rect 235826 308898 236062 309134
rect 236146 308898 236382 309134
rect 235826 273218 236062 273454
rect 236146 273218 236382 273454
rect 235826 272898 236062 273134
rect 236146 272898 236382 273134
rect 235826 237218 236062 237454
rect 236146 237218 236382 237454
rect 235826 236898 236062 237134
rect 236146 236898 236382 237134
rect 235826 201218 236062 201454
rect 236146 201218 236382 201454
rect 235826 200898 236062 201134
rect 236146 200898 236382 201134
rect 235826 165218 236062 165454
rect 236146 165218 236382 165454
rect 235826 164898 236062 165134
rect 236146 164898 236382 165134
rect 235826 129218 236062 129454
rect 236146 129218 236382 129454
rect 235826 128898 236062 129134
rect 236146 128898 236382 129134
rect 235826 93218 236062 93454
rect 236146 93218 236382 93454
rect 235826 92898 236062 93134
rect 236146 92898 236382 93134
rect 235826 57218 236062 57454
rect 236146 57218 236382 57454
rect 235826 56898 236062 57134
rect 236146 56898 236382 57134
rect 235826 21218 236062 21454
rect 236146 21218 236382 21454
rect 235826 20898 236062 21134
rect 236146 20898 236382 21134
rect 235826 -4422 236062 -4186
rect 236146 -4422 236382 -4186
rect 235826 -4742 236062 -4506
rect 236146 -4742 236382 -4506
rect 240326 709402 240562 709638
rect 240646 709402 240882 709638
rect 240326 709082 240562 709318
rect 240646 709082 240882 709318
rect 240326 673718 240562 673954
rect 240646 673718 240882 673954
rect 240326 673398 240562 673634
rect 240646 673398 240882 673634
rect 240326 637718 240562 637954
rect 240646 637718 240882 637954
rect 240326 637398 240562 637634
rect 240646 637398 240882 637634
rect 240326 601718 240562 601954
rect 240646 601718 240882 601954
rect 240326 601398 240562 601634
rect 240646 601398 240882 601634
rect 240326 565718 240562 565954
rect 240646 565718 240882 565954
rect 240326 565398 240562 565634
rect 240646 565398 240882 565634
rect 240326 529718 240562 529954
rect 240646 529718 240882 529954
rect 240326 529398 240562 529634
rect 240646 529398 240882 529634
rect 240326 493718 240562 493954
rect 240646 493718 240882 493954
rect 240326 493398 240562 493634
rect 240646 493398 240882 493634
rect 240326 457718 240562 457954
rect 240646 457718 240882 457954
rect 240326 457398 240562 457634
rect 240646 457398 240882 457634
rect 240326 421718 240562 421954
rect 240646 421718 240882 421954
rect 240326 421398 240562 421634
rect 240646 421398 240882 421634
rect 240326 385718 240562 385954
rect 240646 385718 240882 385954
rect 240326 385398 240562 385634
rect 240646 385398 240882 385634
rect 240326 349718 240562 349954
rect 240646 349718 240882 349954
rect 240326 349398 240562 349634
rect 240646 349398 240882 349634
rect 240326 313718 240562 313954
rect 240646 313718 240882 313954
rect 240326 313398 240562 313634
rect 240646 313398 240882 313634
rect 240326 277718 240562 277954
rect 240646 277718 240882 277954
rect 240326 277398 240562 277634
rect 240646 277398 240882 277634
rect 240326 241718 240562 241954
rect 240646 241718 240882 241954
rect 240326 241398 240562 241634
rect 240646 241398 240882 241634
rect 240326 205718 240562 205954
rect 240646 205718 240882 205954
rect 240326 205398 240562 205634
rect 240646 205398 240882 205634
rect 240326 169718 240562 169954
rect 240646 169718 240882 169954
rect 240326 169398 240562 169634
rect 240646 169398 240882 169634
rect 240326 133718 240562 133954
rect 240646 133718 240882 133954
rect 240326 133398 240562 133634
rect 240646 133398 240882 133634
rect 240326 97718 240562 97954
rect 240646 97718 240882 97954
rect 240326 97398 240562 97634
rect 240646 97398 240882 97634
rect 240326 61718 240562 61954
rect 240646 61718 240882 61954
rect 240326 61398 240562 61634
rect 240646 61398 240882 61634
rect 240326 25718 240562 25954
rect 240646 25718 240882 25954
rect 240326 25398 240562 25634
rect 240646 25398 240882 25634
rect 240326 -5382 240562 -5146
rect 240646 -5382 240882 -5146
rect 240326 -5702 240562 -5466
rect 240646 -5702 240882 -5466
rect 244826 710362 245062 710598
rect 245146 710362 245382 710598
rect 244826 710042 245062 710278
rect 245146 710042 245382 710278
rect 244826 678218 245062 678454
rect 245146 678218 245382 678454
rect 244826 677898 245062 678134
rect 245146 677898 245382 678134
rect 244826 642218 245062 642454
rect 245146 642218 245382 642454
rect 244826 641898 245062 642134
rect 245146 641898 245382 642134
rect 244826 606218 245062 606454
rect 245146 606218 245382 606454
rect 244826 605898 245062 606134
rect 245146 605898 245382 606134
rect 244826 570218 245062 570454
rect 245146 570218 245382 570454
rect 244826 569898 245062 570134
rect 245146 569898 245382 570134
rect 244826 534218 245062 534454
rect 245146 534218 245382 534454
rect 244826 533898 245062 534134
rect 245146 533898 245382 534134
rect 244826 498218 245062 498454
rect 245146 498218 245382 498454
rect 244826 497898 245062 498134
rect 245146 497898 245382 498134
rect 244826 462218 245062 462454
rect 245146 462218 245382 462454
rect 244826 461898 245062 462134
rect 245146 461898 245382 462134
rect 244826 426218 245062 426454
rect 245146 426218 245382 426454
rect 244826 425898 245062 426134
rect 245146 425898 245382 426134
rect 244826 390218 245062 390454
rect 245146 390218 245382 390454
rect 244826 389898 245062 390134
rect 245146 389898 245382 390134
rect 244826 354218 245062 354454
rect 245146 354218 245382 354454
rect 244826 353898 245062 354134
rect 245146 353898 245382 354134
rect 244826 318218 245062 318454
rect 245146 318218 245382 318454
rect 244826 317898 245062 318134
rect 245146 317898 245382 318134
rect 244826 282218 245062 282454
rect 245146 282218 245382 282454
rect 244826 281898 245062 282134
rect 245146 281898 245382 282134
rect 244826 246218 245062 246454
rect 245146 246218 245382 246454
rect 244826 245898 245062 246134
rect 245146 245898 245382 246134
rect 244826 210218 245062 210454
rect 245146 210218 245382 210454
rect 244826 209898 245062 210134
rect 245146 209898 245382 210134
rect 244826 174218 245062 174454
rect 245146 174218 245382 174454
rect 244826 173898 245062 174134
rect 245146 173898 245382 174134
rect 244826 138218 245062 138454
rect 245146 138218 245382 138454
rect 244826 137898 245062 138134
rect 245146 137898 245382 138134
rect 244826 102218 245062 102454
rect 245146 102218 245382 102454
rect 244826 101898 245062 102134
rect 245146 101898 245382 102134
rect 244826 66218 245062 66454
rect 245146 66218 245382 66454
rect 244826 65898 245062 66134
rect 245146 65898 245382 66134
rect 244826 30218 245062 30454
rect 245146 30218 245382 30454
rect 244826 29898 245062 30134
rect 245146 29898 245382 30134
rect 244826 -6342 245062 -6106
rect 245146 -6342 245382 -6106
rect 244826 -6662 245062 -6426
rect 245146 -6662 245382 -6426
rect 249326 711322 249562 711558
rect 249646 711322 249882 711558
rect 249326 711002 249562 711238
rect 249646 711002 249882 711238
rect 249326 682718 249562 682954
rect 249646 682718 249882 682954
rect 249326 682398 249562 682634
rect 249646 682398 249882 682634
rect 249326 646718 249562 646954
rect 249646 646718 249882 646954
rect 249326 646398 249562 646634
rect 249646 646398 249882 646634
rect 249326 610718 249562 610954
rect 249646 610718 249882 610954
rect 249326 610398 249562 610634
rect 249646 610398 249882 610634
rect 249326 574718 249562 574954
rect 249646 574718 249882 574954
rect 249326 574398 249562 574634
rect 249646 574398 249882 574634
rect 249326 538718 249562 538954
rect 249646 538718 249882 538954
rect 249326 538398 249562 538634
rect 249646 538398 249882 538634
rect 249326 502718 249562 502954
rect 249646 502718 249882 502954
rect 249326 502398 249562 502634
rect 249646 502398 249882 502634
rect 249326 466718 249562 466954
rect 249646 466718 249882 466954
rect 249326 466398 249562 466634
rect 249646 466398 249882 466634
rect 249326 430718 249562 430954
rect 249646 430718 249882 430954
rect 249326 430398 249562 430634
rect 249646 430398 249882 430634
rect 249326 394718 249562 394954
rect 249646 394718 249882 394954
rect 249326 394398 249562 394634
rect 249646 394398 249882 394634
rect 249326 358718 249562 358954
rect 249646 358718 249882 358954
rect 249326 358398 249562 358634
rect 249646 358398 249882 358634
rect 249326 322718 249562 322954
rect 249646 322718 249882 322954
rect 249326 322398 249562 322634
rect 249646 322398 249882 322634
rect 249326 286718 249562 286954
rect 249646 286718 249882 286954
rect 249326 286398 249562 286634
rect 249646 286398 249882 286634
rect 249326 250718 249562 250954
rect 249646 250718 249882 250954
rect 249326 250398 249562 250634
rect 249646 250398 249882 250634
rect 249326 214718 249562 214954
rect 249646 214718 249882 214954
rect 249326 214398 249562 214634
rect 249646 214398 249882 214634
rect 249326 178718 249562 178954
rect 249646 178718 249882 178954
rect 249326 178398 249562 178634
rect 249646 178398 249882 178634
rect 249326 142718 249562 142954
rect 249646 142718 249882 142954
rect 249326 142398 249562 142634
rect 249646 142398 249882 142634
rect 249326 106718 249562 106954
rect 249646 106718 249882 106954
rect 249326 106398 249562 106634
rect 249646 106398 249882 106634
rect 249326 70718 249562 70954
rect 249646 70718 249882 70954
rect 249326 70398 249562 70634
rect 249646 70398 249882 70634
rect 249326 34718 249562 34954
rect 249646 34718 249882 34954
rect 249326 34398 249562 34634
rect 249646 34398 249882 34634
rect 249326 -7302 249562 -7066
rect 249646 -7302 249882 -7066
rect 249326 -7622 249562 -7386
rect 249646 -7622 249882 -7386
rect 253826 704602 254062 704838
rect 254146 704602 254382 704838
rect 253826 704282 254062 704518
rect 254146 704282 254382 704518
rect 253826 687218 254062 687454
rect 254146 687218 254382 687454
rect 253826 686898 254062 687134
rect 254146 686898 254382 687134
rect 253826 651218 254062 651454
rect 254146 651218 254382 651454
rect 253826 650898 254062 651134
rect 254146 650898 254382 651134
rect 253826 615218 254062 615454
rect 254146 615218 254382 615454
rect 253826 614898 254062 615134
rect 254146 614898 254382 615134
rect 253826 579218 254062 579454
rect 254146 579218 254382 579454
rect 253826 578898 254062 579134
rect 254146 578898 254382 579134
rect 253826 543218 254062 543454
rect 254146 543218 254382 543454
rect 253826 542898 254062 543134
rect 254146 542898 254382 543134
rect 253826 507218 254062 507454
rect 254146 507218 254382 507454
rect 253826 506898 254062 507134
rect 254146 506898 254382 507134
rect 253826 471218 254062 471454
rect 254146 471218 254382 471454
rect 253826 470898 254062 471134
rect 254146 470898 254382 471134
rect 253826 435218 254062 435454
rect 254146 435218 254382 435454
rect 253826 434898 254062 435134
rect 254146 434898 254382 435134
rect 253826 399218 254062 399454
rect 254146 399218 254382 399454
rect 253826 398898 254062 399134
rect 254146 398898 254382 399134
rect 253826 363218 254062 363454
rect 254146 363218 254382 363454
rect 253826 362898 254062 363134
rect 254146 362898 254382 363134
rect 253826 327218 254062 327454
rect 254146 327218 254382 327454
rect 253826 326898 254062 327134
rect 254146 326898 254382 327134
rect 253826 291218 254062 291454
rect 254146 291218 254382 291454
rect 253826 290898 254062 291134
rect 254146 290898 254382 291134
rect 253826 255218 254062 255454
rect 254146 255218 254382 255454
rect 253826 254898 254062 255134
rect 254146 254898 254382 255134
rect 253826 219218 254062 219454
rect 254146 219218 254382 219454
rect 253826 218898 254062 219134
rect 254146 218898 254382 219134
rect 253826 183218 254062 183454
rect 254146 183218 254382 183454
rect 253826 182898 254062 183134
rect 254146 182898 254382 183134
rect 253826 147218 254062 147454
rect 254146 147218 254382 147454
rect 253826 146898 254062 147134
rect 254146 146898 254382 147134
rect 253826 111218 254062 111454
rect 254146 111218 254382 111454
rect 253826 110898 254062 111134
rect 254146 110898 254382 111134
rect 253826 75218 254062 75454
rect 254146 75218 254382 75454
rect 253826 74898 254062 75134
rect 254146 74898 254382 75134
rect 253826 39218 254062 39454
rect 254146 39218 254382 39454
rect 253826 38898 254062 39134
rect 254146 38898 254382 39134
rect 253826 3218 254062 3454
rect 254146 3218 254382 3454
rect 253826 2898 254062 3134
rect 254146 2898 254382 3134
rect 253826 -582 254062 -346
rect 254146 -582 254382 -346
rect 253826 -902 254062 -666
rect 254146 -902 254382 -666
rect 258326 705562 258562 705798
rect 258646 705562 258882 705798
rect 258326 705242 258562 705478
rect 258646 705242 258882 705478
rect 258326 691718 258562 691954
rect 258646 691718 258882 691954
rect 258326 691398 258562 691634
rect 258646 691398 258882 691634
rect 258326 655718 258562 655954
rect 258646 655718 258882 655954
rect 258326 655398 258562 655634
rect 258646 655398 258882 655634
rect 258326 619718 258562 619954
rect 258646 619718 258882 619954
rect 258326 619398 258562 619634
rect 258646 619398 258882 619634
rect 258326 583718 258562 583954
rect 258646 583718 258882 583954
rect 258326 583398 258562 583634
rect 258646 583398 258882 583634
rect 258326 547718 258562 547954
rect 258646 547718 258882 547954
rect 258326 547398 258562 547634
rect 258646 547398 258882 547634
rect 258326 511718 258562 511954
rect 258646 511718 258882 511954
rect 258326 511398 258562 511634
rect 258646 511398 258882 511634
rect 258326 475718 258562 475954
rect 258646 475718 258882 475954
rect 258326 475398 258562 475634
rect 258646 475398 258882 475634
rect 258326 439718 258562 439954
rect 258646 439718 258882 439954
rect 258326 439398 258562 439634
rect 258646 439398 258882 439634
rect 258326 403718 258562 403954
rect 258646 403718 258882 403954
rect 258326 403398 258562 403634
rect 258646 403398 258882 403634
rect 258326 367718 258562 367954
rect 258646 367718 258882 367954
rect 258326 367398 258562 367634
rect 258646 367398 258882 367634
rect 258326 331718 258562 331954
rect 258646 331718 258882 331954
rect 258326 331398 258562 331634
rect 258646 331398 258882 331634
rect 258326 295718 258562 295954
rect 258646 295718 258882 295954
rect 258326 295398 258562 295634
rect 258646 295398 258882 295634
rect 258326 259718 258562 259954
rect 258646 259718 258882 259954
rect 258326 259398 258562 259634
rect 258646 259398 258882 259634
rect 258326 223718 258562 223954
rect 258646 223718 258882 223954
rect 258326 223398 258562 223634
rect 258646 223398 258882 223634
rect 258326 187718 258562 187954
rect 258646 187718 258882 187954
rect 258326 187398 258562 187634
rect 258646 187398 258882 187634
rect 258326 151718 258562 151954
rect 258646 151718 258882 151954
rect 258326 151398 258562 151634
rect 258646 151398 258882 151634
rect 258326 115718 258562 115954
rect 258646 115718 258882 115954
rect 258326 115398 258562 115634
rect 258646 115398 258882 115634
rect 258326 79718 258562 79954
rect 258646 79718 258882 79954
rect 258326 79398 258562 79634
rect 258646 79398 258882 79634
rect 258326 43718 258562 43954
rect 258646 43718 258882 43954
rect 258326 43398 258562 43634
rect 258646 43398 258882 43634
rect 258326 7718 258562 7954
rect 258646 7718 258882 7954
rect 258326 7398 258562 7634
rect 258646 7398 258882 7634
rect 258326 -1542 258562 -1306
rect 258646 -1542 258882 -1306
rect 258326 -1862 258562 -1626
rect 258646 -1862 258882 -1626
rect 262826 706522 263062 706758
rect 263146 706522 263382 706758
rect 262826 706202 263062 706438
rect 263146 706202 263382 706438
rect 262826 696218 263062 696454
rect 263146 696218 263382 696454
rect 262826 695898 263062 696134
rect 263146 695898 263382 696134
rect 262826 660218 263062 660454
rect 263146 660218 263382 660454
rect 262826 659898 263062 660134
rect 263146 659898 263382 660134
rect 262826 624218 263062 624454
rect 263146 624218 263382 624454
rect 262826 623898 263062 624134
rect 263146 623898 263382 624134
rect 262826 588218 263062 588454
rect 263146 588218 263382 588454
rect 262826 587898 263062 588134
rect 263146 587898 263382 588134
rect 262826 552218 263062 552454
rect 263146 552218 263382 552454
rect 262826 551898 263062 552134
rect 263146 551898 263382 552134
rect 262826 516218 263062 516454
rect 263146 516218 263382 516454
rect 262826 515898 263062 516134
rect 263146 515898 263382 516134
rect 262826 480218 263062 480454
rect 263146 480218 263382 480454
rect 262826 479898 263062 480134
rect 263146 479898 263382 480134
rect 262826 444218 263062 444454
rect 263146 444218 263382 444454
rect 262826 443898 263062 444134
rect 263146 443898 263382 444134
rect 262826 408218 263062 408454
rect 263146 408218 263382 408454
rect 262826 407898 263062 408134
rect 263146 407898 263382 408134
rect 262826 372218 263062 372454
rect 263146 372218 263382 372454
rect 262826 371898 263062 372134
rect 263146 371898 263382 372134
rect 262826 336218 263062 336454
rect 263146 336218 263382 336454
rect 262826 335898 263062 336134
rect 263146 335898 263382 336134
rect 262826 300218 263062 300454
rect 263146 300218 263382 300454
rect 262826 299898 263062 300134
rect 263146 299898 263382 300134
rect 262826 264218 263062 264454
rect 263146 264218 263382 264454
rect 262826 263898 263062 264134
rect 263146 263898 263382 264134
rect 262826 228218 263062 228454
rect 263146 228218 263382 228454
rect 262826 227898 263062 228134
rect 263146 227898 263382 228134
rect 262826 192218 263062 192454
rect 263146 192218 263382 192454
rect 262826 191898 263062 192134
rect 263146 191898 263382 192134
rect 262826 156218 263062 156454
rect 263146 156218 263382 156454
rect 262826 155898 263062 156134
rect 263146 155898 263382 156134
rect 262826 120218 263062 120454
rect 263146 120218 263382 120454
rect 262826 119898 263062 120134
rect 263146 119898 263382 120134
rect 262826 84218 263062 84454
rect 263146 84218 263382 84454
rect 262826 83898 263062 84134
rect 263146 83898 263382 84134
rect 262826 48218 263062 48454
rect 263146 48218 263382 48454
rect 262826 47898 263062 48134
rect 263146 47898 263382 48134
rect 262826 12218 263062 12454
rect 263146 12218 263382 12454
rect 262826 11898 263062 12134
rect 263146 11898 263382 12134
rect 262826 -2502 263062 -2266
rect 263146 -2502 263382 -2266
rect 262826 -2822 263062 -2586
rect 263146 -2822 263382 -2586
rect 267326 707482 267562 707718
rect 267646 707482 267882 707718
rect 267326 707162 267562 707398
rect 267646 707162 267882 707398
rect 267326 700718 267562 700954
rect 267646 700718 267882 700954
rect 267326 700398 267562 700634
rect 267646 700398 267882 700634
rect 267326 664718 267562 664954
rect 267646 664718 267882 664954
rect 267326 664398 267562 664634
rect 267646 664398 267882 664634
rect 267326 628718 267562 628954
rect 267646 628718 267882 628954
rect 267326 628398 267562 628634
rect 267646 628398 267882 628634
rect 267326 592718 267562 592954
rect 267646 592718 267882 592954
rect 267326 592398 267562 592634
rect 267646 592398 267882 592634
rect 267326 556718 267562 556954
rect 267646 556718 267882 556954
rect 267326 556398 267562 556634
rect 267646 556398 267882 556634
rect 267326 520718 267562 520954
rect 267646 520718 267882 520954
rect 267326 520398 267562 520634
rect 267646 520398 267882 520634
rect 267326 484718 267562 484954
rect 267646 484718 267882 484954
rect 267326 484398 267562 484634
rect 267646 484398 267882 484634
rect 267326 448718 267562 448954
rect 267646 448718 267882 448954
rect 267326 448398 267562 448634
rect 267646 448398 267882 448634
rect 267326 412718 267562 412954
rect 267646 412718 267882 412954
rect 267326 412398 267562 412634
rect 267646 412398 267882 412634
rect 267326 376718 267562 376954
rect 267646 376718 267882 376954
rect 267326 376398 267562 376634
rect 267646 376398 267882 376634
rect 267326 340718 267562 340954
rect 267646 340718 267882 340954
rect 267326 340398 267562 340634
rect 267646 340398 267882 340634
rect 267326 304718 267562 304954
rect 267646 304718 267882 304954
rect 267326 304398 267562 304634
rect 267646 304398 267882 304634
rect 267326 268718 267562 268954
rect 267646 268718 267882 268954
rect 267326 268398 267562 268634
rect 267646 268398 267882 268634
rect 267326 232718 267562 232954
rect 267646 232718 267882 232954
rect 267326 232398 267562 232634
rect 267646 232398 267882 232634
rect 267326 196718 267562 196954
rect 267646 196718 267882 196954
rect 267326 196398 267562 196634
rect 267646 196398 267882 196634
rect 267326 160718 267562 160954
rect 267646 160718 267882 160954
rect 267326 160398 267562 160634
rect 267646 160398 267882 160634
rect 267326 124718 267562 124954
rect 267646 124718 267882 124954
rect 267326 124398 267562 124634
rect 267646 124398 267882 124634
rect 267326 88718 267562 88954
rect 267646 88718 267882 88954
rect 267326 88398 267562 88634
rect 267646 88398 267882 88634
rect 267326 52718 267562 52954
rect 267646 52718 267882 52954
rect 267326 52398 267562 52634
rect 267646 52398 267882 52634
rect 267326 16718 267562 16954
rect 267646 16718 267882 16954
rect 267326 16398 267562 16634
rect 267646 16398 267882 16634
rect 267326 -3462 267562 -3226
rect 267646 -3462 267882 -3226
rect 267326 -3782 267562 -3546
rect 267646 -3782 267882 -3546
rect 271826 708442 272062 708678
rect 272146 708442 272382 708678
rect 271826 708122 272062 708358
rect 272146 708122 272382 708358
rect 271826 669218 272062 669454
rect 272146 669218 272382 669454
rect 271826 668898 272062 669134
rect 272146 668898 272382 669134
rect 271826 633218 272062 633454
rect 272146 633218 272382 633454
rect 271826 632898 272062 633134
rect 272146 632898 272382 633134
rect 271826 597218 272062 597454
rect 272146 597218 272382 597454
rect 271826 596898 272062 597134
rect 272146 596898 272382 597134
rect 271826 561218 272062 561454
rect 272146 561218 272382 561454
rect 271826 560898 272062 561134
rect 272146 560898 272382 561134
rect 271826 525218 272062 525454
rect 272146 525218 272382 525454
rect 271826 524898 272062 525134
rect 272146 524898 272382 525134
rect 271826 489218 272062 489454
rect 272146 489218 272382 489454
rect 271826 488898 272062 489134
rect 272146 488898 272382 489134
rect 271826 453218 272062 453454
rect 272146 453218 272382 453454
rect 271826 452898 272062 453134
rect 272146 452898 272382 453134
rect 271826 417218 272062 417454
rect 272146 417218 272382 417454
rect 271826 416898 272062 417134
rect 272146 416898 272382 417134
rect 271826 381218 272062 381454
rect 272146 381218 272382 381454
rect 271826 380898 272062 381134
rect 272146 380898 272382 381134
rect 271826 345218 272062 345454
rect 272146 345218 272382 345454
rect 271826 344898 272062 345134
rect 272146 344898 272382 345134
rect 271826 309218 272062 309454
rect 272146 309218 272382 309454
rect 271826 308898 272062 309134
rect 272146 308898 272382 309134
rect 271826 273218 272062 273454
rect 272146 273218 272382 273454
rect 271826 272898 272062 273134
rect 272146 272898 272382 273134
rect 271826 237218 272062 237454
rect 272146 237218 272382 237454
rect 271826 236898 272062 237134
rect 272146 236898 272382 237134
rect 271826 201218 272062 201454
rect 272146 201218 272382 201454
rect 271826 200898 272062 201134
rect 272146 200898 272382 201134
rect 271826 165218 272062 165454
rect 272146 165218 272382 165454
rect 271826 164898 272062 165134
rect 272146 164898 272382 165134
rect 271826 129218 272062 129454
rect 272146 129218 272382 129454
rect 271826 128898 272062 129134
rect 272146 128898 272382 129134
rect 271826 93218 272062 93454
rect 272146 93218 272382 93454
rect 271826 92898 272062 93134
rect 272146 92898 272382 93134
rect 271826 57218 272062 57454
rect 272146 57218 272382 57454
rect 271826 56898 272062 57134
rect 272146 56898 272382 57134
rect 271826 21218 272062 21454
rect 272146 21218 272382 21454
rect 271826 20898 272062 21134
rect 272146 20898 272382 21134
rect 271826 -4422 272062 -4186
rect 272146 -4422 272382 -4186
rect 271826 -4742 272062 -4506
rect 272146 -4742 272382 -4506
rect 276326 709402 276562 709638
rect 276646 709402 276882 709638
rect 276326 709082 276562 709318
rect 276646 709082 276882 709318
rect 276326 673718 276562 673954
rect 276646 673718 276882 673954
rect 276326 673398 276562 673634
rect 276646 673398 276882 673634
rect 276326 637718 276562 637954
rect 276646 637718 276882 637954
rect 276326 637398 276562 637634
rect 276646 637398 276882 637634
rect 276326 601718 276562 601954
rect 276646 601718 276882 601954
rect 276326 601398 276562 601634
rect 276646 601398 276882 601634
rect 276326 565718 276562 565954
rect 276646 565718 276882 565954
rect 276326 565398 276562 565634
rect 276646 565398 276882 565634
rect 276326 529718 276562 529954
rect 276646 529718 276882 529954
rect 276326 529398 276562 529634
rect 276646 529398 276882 529634
rect 276326 493718 276562 493954
rect 276646 493718 276882 493954
rect 276326 493398 276562 493634
rect 276646 493398 276882 493634
rect 276326 457718 276562 457954
rect 276646 457718 276882 457954
rect 276326 457398 276562 457634
rect 276646 457398 276882 457634
rect 276326 421718 276562 421954
rect 276646 421718 276882 421954
rect 276326 421398 276562 421634
rect 276646 421398 276882 421634
rect 276326 385718 276562 385954
rect 276646 385718 276882 385954
rect 276326 385398 276562 385634
rect 276646 385398 276882 385634
rect 276326 349718 276562 349954
rect 276646 349718 276882 349954
rect 276326 349398 276562 349634
rect 276646 349398 276882 349634
rect 276326 313718 276562 313954
rect 276646 313718 276882 313954
rect 276326 313398 276562 313634
rect 276646 313398 276882 313634
rect 276326 277718 276562 277954
rect 276646 277718 276882 277954
rect 276326 277398 276562 277634
rect 276646 277398 276882 277634
rect 276326 241718 276562 241954
rect 276646 241718 276882 241954
rect 276326 241398 276562 241634
rect 276646 241398 276882 241634
rect 276326 205718 276562 205954
rect 276646 205718 276882 205954
rect 276326 205398 276562 205634
rect 276646 205398 276882 205634
rect 276326 169718 276562 169954
rect 276646 169718 276882 169954
rect 276326 169398 276562 169634
rect 276646 169398 276882 169634
rect 276326 133718 276562 133954
rect 276646 133718 276882 133954
rect 276326 133398 276562 133634
rect 276646 133398 276882 133634
rect 276326 97718 276562 97954
rect 276646 97718 276882 97954
rect 276326 97398 276562 97634
rect 276646 97398 276882 97634
rect 276326 61718 276562 61954
rect 276646 61718 276882 61954
rect 276326 61398 276562 61634
rect 276646 61398 276882 61634
rect 276326 25718 276562 25954
rect 276646 25718 276882 25954
rect 276326 25398 276562 25634
rect 276646 25398 276882 25634
rect 276326 -5382 276562 -5146
rect 276646 -5382 276882 -5146
rect 276326 -5702 276562 -5466
rect 276646 -5702 276882 -5466
rect 280826 710362 281062 710598
rect 281146 710362 281382 710598
rect 280826 710042 281062 710278
rect 281146 710042 281382 710278
rect 280826 678218 281062 678454
rect 281146 678218 281382 678454
rect 280826 677898 281062 678134
rect 281146 677898 281382 678134
rect 280826 642218 281062 642454
rect 281146 642218 281382 642454
rect 280826 641898 281062 642134
rect 281146 641898 281382 642134
rect 280826 606218 281062 606454
rect 281146 606218 281382 606454
rect 280826 605898 281062 606134
rect 281146 605898 281382 606134
rect 280826 570218 281062 570454
rect 281146 570218 281382 570454
rect 280826 569898 281062 570134
rect 281146 569898 281382 570134
rect 280826 534218 281062 534454
rect 281146 534218 281382 534454
rect 280826 533898 281062 534134
rect 281146 533898 281382 534134
rect 280826 498218 281062 498454
rect 281146 498218 281382 498454
rect 280826 497898 281062 498134
rect 281146 497898 281382 498134
rect 280826 462218 281062 462454
rect 281146 462218 281382 462454
rect 280826 461898 281062 462134
rect 281146 461898 281382 462134
rect 280826 426218 281062 426454
rect 281146 426218 281382 426454
rect 280826 425898 281062 426134
rect 281146 425898 281382 426134
rect 280826 390218 281062 390454
rect 281146 390218 281382 390454
rect 280826 389898 281062 390134
rect 281146 389898 281382 390134
rect 280826 354218 281062 354454
rect 281146 354218 281382 354454
rect 280826 353898 281062 354134
rect 281146 353898 281382 354134
rect 280826 318218 281062 318454
rect 281146 318218 281382 318454
rect 280826 317898 281062 318134
rect 281146 317898 281382 318134
rect 280826 282218 281062 282454
rect 281146 282218 281382 282454
rect 280826 281898 281062 282134
rect 281146 281898 281382 282134
rect 280826 246218 281062 246454
rect 281146 246218 281382 246454
rect 280826 245898 281062 246134
rect 281146 245898 281382 246134
rect 280826 210218 281062 210454
rect 281146 210218 281382 210454
rect 280826 209898 281062 210134
rect 281146 209898 281382 210134
rect 280826 174218 281062 174454
rect 281146 174218 281382 174454
rect 280826 173898 281062 174134
rect 281146 173898 281382 174134
rect 280826 138218 281062 138454
rect 281146 138218 281382 138454
rect 280826 137898 281062 138134
rect 281146 137898 281382 138134
rect 280826 102218 281062 102454
rect 281146 102218 281382 102454
rect 280826 101898 281062 102134
rect 281146 101898 281382 102134
rect 280826 66218 281062 66454
rect 281146 66218 281382 66454
rect 280826 65898 281062 66134
rect 281146 65898 281382 66134
rect 280826 30218 281062 30454
rect 281146 30218 281382 30454
rect 280826 29898 281062 30134
rect 281146 29898 281382 30134
rect 280826 -6342 281062 -6106
rect 281146 -6342 281382 -6106
rect 280826 -6662 281062 -6426
rect 281146 -6662 281382 -6426
rect 285326 711322 285562 711558
rect 285646 711322 285882 711558
rect 285326 711002 285562 711238
rect 285646 711002 285882 711238
rect 285326 682718 285562 682954
rect 285646 682718 285882 682954
rect 285326 682398 285562 682634
rect 285646 682398 285882 682634
rect 285326 646718 285562 646954
rect 285646 646718 285882 646954
rect 285326 646398 285562 646634
rect 285646 646398 285882 646634
rect 285326 610718 285562 610954
rect 285646 610718 285882 610954
rect 285326 610398 285562 610634
rect 285646 610398 285882 610634
rect 285326 574718 285562 574954
rect 285646 574718 285882 574954
rect 285326 574398 285562 574634
rect 285646 574398 285882 574634
rect 285326 538718 285562 538954
rect 285646 538718 285882 538954
rect 285326 538398 285562 538634
rect 285646 538398 285882 538634
rect 285326 502718 285562 502954
rect 285646 502718 285882 502954
rect 285326 502398 285562 502634
rect 285646 502398 285882 502634
rect 285326 466718 285562 466954
rect 285646 466718 285882 466954
rect 285326 466398 285562 466634
rect 285646 466398 285882 466634
rect 285326 430718 285562 430954
rect 285646 430718 285882 430954
rect 285326 430398 285562 430634
rect 285646 430398 285882 430634
rect 285326 394718 285562 394954
rect 285646 394718 285882 394954
rect 285326 394398 285562 394634
rect 285646 394398 285882 394634
rect 285326 358718 285562 358954
rect 285646 358718 285882 358954
rect 285326 358398 285562 358634
rect 285646 358398 285882 358634
rect 285326 322718 285562 322954
rect 285646 322718 285882 322954
rect 285326 322398 285562 322634
rect 285646 322398 285882 322634
rect 285326 286718 285562 286954
rect 285646 286718 285882 286954
rect 285326 286398 285562 286634
rect 285646 286398 285882 286634
rect 285326 250718 285562 250954
rect 285646 250718 285882 250954
rect 285326 250398 285562 250634
rect 285646 250398 285882 250634
rect 285326 214718 285562 214954
rect 285646 214718 285882 214954
rect 285326 214398 285562 214634
rect 285646 214398 285882 214634
rect 285326 178718 285562 178954
rect 285646 178718 285882 178954
rect 285326 178398 285562 178634
rect 285646 178398 285882 178634
rect 285326 142718 285562 142954
rect 285646 142718 285882 142954
rect 285326 142398 285562 142634
rect 285646 142398 285882 142634
rect 285326 106718 285562 106954
rect 285646 106718 285882 106954
rect 285326 106398 285562 106634
rect 285646 106398 285882 106634
rect 285326 70718 285562 70954
rect 285646 70718 285882 70954
rect 285326 70398 285562 70634
rect 285646 70398 285882 70634
rect 285326 34718 285562 34954
rect 285646 34718 285882 34954
rect 285326 34398 285562 34634
rect 285646 34398 285882 34634
rect 285326 -7302 285562 -7066
rect 285646 -7302 285882 -7066
rect 285326 -7622 285562 -7386
rect 285646 -7622 285882 -7386
rect 289826 704602 290062 704838
rect 290146 704602 290382 704838
rect 289826 704282 290062 704518
rect 290146 704282 290382 704518
rect 289826 687218 290062 687454
rect 290146 687218 290382 687454
rect 289826 686898 290062 687134
rect 290146 686898 290382 687134
rect 289826 651218 290062 651454
rect 290146 651218 290382 651454
rect 289826 650898 290062 651134
rect 290146 650898 290382 651134
rect 289826 615218 290062 615454
rect 290146 615218 290382 615454
rect 289826 614898 290062 615134
rect 290146 614898 290382 615134
rect 289826 579218 290062 579454
rect 290146 579218 290382 579454
rect 289826 578898 290062 579134
rect 290146 578898 290382 579134
rect 289826 543218 290062 543454
rect 290146 543218 290382 543454
rect 289826 542898 290062 543134
rect 290146 542898 290382 543134
rect 289826 507218 290062 507454
rect 290146 507218 290382 507454
rect 289826 506898 290062 507134
rect 290146 506898 290382 507134
rect 289826 471218 290062 471454
rect 290146 471218 290382 471454
rect 289826 470898 290062 471134
rect 290146 470898 290382 471134
rect 289826 435218 290062 435454
rect 290146 435218 290382 435454
rect 289826 434898 290062 435134
rect 290146 434898 290382 435134
rect 289826 399218 290062 399454
rect 290146 399218 290382 399454
rect 289826 398898 290062 399134
rect 290146 398898 290382 399134
rect 289826 363218 290062 363454
rect 290146 363218 290382 363454
rect 289826 362898 290062 363134
rect 290146 362898 290382 363134
rect 289826 327218 290062 327454
rect 290146 327218 290382 327454
rect 289826 326898 290062 327134
rect 290146 326898 290382 327134
rect 289826 291218 290062 291454
rect 290146 291218 290382 291454
rect 289826 290898 290062 291134
rect 290146 290898 290382 291134
rect 289826 255218 290062 255454
rect 290146 255218 290382 255454
rect 289826 254898 290062 255134
rect 290146 254898 290382 255134
rect 289826 219218 290062 219454
rect 290146 219218 290382 219454
rect 289826 218898 290062 219134
rect 290146 218898 290382 219134
rect 289826 183218 290062 183454
rect 290146 183218 290382 183454
rect 289826 182898 290062 183134
rect 290146 182898 290382 183134
rect 289826 147218 290062 147454
rect 290146 147218 290382 147454
rect 289826 146898 290062 147134
rect 290146 146898 290382 147134
rect 289826 111218 290062 111454
rect 290146 111218 290382 111454
rect 289826 110898 290062 111134
rect 290146 110898 290382 111134
rect 289826 75218 290062 75454
rect 290146 75218 290382 75454
rect 289826 74898 290062 75134
rect 290146 74898 290382 75134
rect 289826 39218 290062 39454
rect 290146 39218 290382 39454
rect 289826 38898 290062 39134
rect 290146 38898 290382 39134
rect 289826 3218 290062 3454
rect 290146 3218 290382 3454
rect 289826 2898 290062 3134
rect 290146 2898 290382 3134
rect 289826 -582 290062 -346
rect 290146 -582 290382 -346
rect 289826 -902 290062 -666
rect 290146 -902 290382 -666
rect 294326 705562 294562 705798
rect 294646 705562 294882 705798
rect 294326 705242 294562 705478
rect 294646 705242 294882 705478
rect 294326 691718 294562 691954
rect 294646 691718 294882 691954
rect 294326 691398 294562 691634
rect 294646 691398 294882 691634
rect 294326 655718 294562 655954
rect 294646 655718 294882 655954
rect 294326 655398 294562 655634
rect 294646 655398 294882 655634
rect 294326 619718 294562 619954
rect 294646 619718 294882 619954
rect 294326 619398 294562 619634
rect 294646 619398 294882 619634
rect 294326 583718 294562 583954
rect 294646 583718 294882 583954
rect 294326 583398 294562 583634
rect 294646 583398 294882 583634
rect 294326 547718 294562 547954
rect 294646 547718 294882 547954
rect 294326 547398 294562 547634
rect 294646 547398 294882 547634
rect 294326 511718 294562 511954
rect 294646 511718 294882 511954
rect 294326 511398 294562 511634
rect 294646 511398 294882 511634
rect 294326 475718 294562 475954
rect 294646 475718 294882 475954
rect 294326 475398 294562 475634
rect 294646 475398 294882 475634
rect 294326 439718 294562 439954
rect 294646 439718 294882 439954
rect 294326 439398 294562 439634
rect 294646 439398 294882 439634
rect 294326 403718 294562 403954
rect 294646 403718 294882 403954
rect 294326 403398 294562 403634
rect 294646 403398 294882 403634
rect 294326 367718 294562 367954
rect 294646 367718 294882 367954
rect 294326 367398 294562 367634
rect 294646 367398 294882 367634
rect 294326 331718 294562 331954
rect 294646 331718 294882 331954
rect 294326 331398 294562 331634
rect 294646 331398 294882 331634
rect 294326 295718 294562 295954
rect 294646 295718 294882 295954
rect 294326 295398 294562 295634
rect 294646 295398 294882 295634
rect 294326 259718 294562 259954
rect 294646 259718 294882 259954
rect 294326 259398 294562 259634
rect 294646 259398 294882 259634
rect 294326 223718 294562 223954
rect 294646 223718 294882 223954
rect 294326 223398 294562 223634
rect 294646 223398 294882 223634
rect 294326 187718 294562 187954
rect 294646 187718 294882 187954
rect 294326 187398 294562 187634
rect 294646 187398 294882 187634
rect 294326 151718 294562 151954
rect 294646 151718 294882 151954
rect 294326 151398 294562 151634
rect 294646 151398 294882 151634
rect 294326 115718 294562 115954
rect 294646 115718 294882 115954
rect 294326 115398 294562 115634
rect 294646 115398 294882 115634
rect 294326 79718 294562 79954
rect 294646 79718 294882 79954
rect 294326 79398 294562 79634
rect 294646 79398 294882 79634
rect 294326 43718 294562 43954
rect 294646 43718 294882 43954
rect 294326 43398 294562 43634
rect 294646 43398 294882 43634
rect 294326 7718 294562 7954
rect 294646 7718 294882 7954
rect 294326 7398 294562 7634
rect 294646 7398 294882 7634
rect 294326 -1542 294562 -1306
rect 294646 -1542 294882 -1306
rect 294326 -1862 294562 -1626
rect 294646 -1862 294882 -1626
rect 298826 706522 299062 706758
rect 299146 706522 299382 706758
rect 298826 706202 299062 706438
rect 299146 706202 299382 706438
rect 298826 696218 299062 696454
rect 299146 696218 299382 696454
rect 298826 695898 299062 696134
rect 299146 695898 299382 696134
rect 298826 660218 299062 660454
rect 299146 660218 299382 660454
rect 298826 659898 299062 660134
rect 299146 659898 299382 660134
rect 298826 624218 299062 624454
rect 299146 624218 299382 624454
rect 298826 623898 299062 624134
rect 299146 623898 299382 624134
rect 298826 588218 299062 588454
rect 299146 588218 299382 588454
rect 298826 587898 299062 588134
rect 299146 587898 299382 588134
rect 298826 552218 299062 552454
rect 299146 552218 299382 552454
rect 298826 551898 299062 552134
rect 299146 551898 299382 552134
rect 298826 516218 299062 516454
rect 299146 516218 299382 516454
rect 298826 515898 299062 516134
rect 299146 515898 299382 516134
rect 298826 480218 299062 480454
rect 299146 480218 299382 480454
rect 298826 479898 299062 480134
rect 299146 479898 299382 480134
rect 298826 444218 299062 444454
rect 299146 444218 299382 444454
rect 298826 443898 299062 444134
rect 299146 443898 299382 444134
rect 298826 408218 299062 408454
rect 299146 408218 299382 408454
rect 298826 407898 299062 408134
rect 299146 407898 299382 408134
rect 298826 372218 299062 372454
rect 299146 372218 299382 372454
rect 298826 371898 299062 372134
rect 299146 371898 299382 372134
rect 298826 336218 299062 336454
rect 299146 336218 299382 336454
rect 298826 335898 299062 336134
rect 299146 335898 299382 336134
rect 298826 300218 299062 300454
rect 299146 300218 299382 300454
rect 298826 299898 299062 300134
rect 299146 299898 299382 300134
rect 298826 264218 299062 264454
rect 299146 264218 299382 264454
rect 298826 263898 299062 264134
rect 299146 263898 299382 264134
rect 298826 228218 299062 228454
rect 299146 228218 299382 228454
rect 298826 227898 299062 228134
rect 299146 227898 299382 228134
rect 298826 192218 299062 192454
rect 299146 192218 299382 192454
rect 298826 191898 299062 192134
rect 299146 191898 299382 192134
rect 298826 156218 299062 156454
rect 299146 156218 299382 156454
rect 298826 155898 299062 156134
rect 299146 155898 299382 156134
rect 298826 120218 299062 120454
rect 299146 120218 299382 120454
rect 298826 119898 299062 120134
rect 299146 119898 299382 120134
rect 298826 84218 299062 84454
rect 299146 84218 299382 84454
rect 298826 83898 299062 84134
rect 299146 83898 299382 84134
rect 298826 48218 299062 48454
rect 299146 48218 299382 48454
rect 298826 47898 299062 48134
rect 299146 47898 299382 48134
rect 298826 12218 299062 12454
rect 299146 12218 299382 12454
rect 298826 11898 299062 12134
rect 299146 11898 299382 12134
rect 298826 -2502 299062 -2266
rect 299146 -2502 299382 -2266
rect 298826 -2822 299062 -2586
rect 299146 -2822 299382 -2586
rect 303326 707482 303562 707718
rect 303646 707482 303882 707718
rect 303326 707162 303562 707398
rect 303646 707162 303882 707398
rect 303326 700718 303562 700954
rect 303646 700718 303882 700954
rect 303326 700398 303562 700634
rect 303646 700398 303882 700634
rect 303326 664718 303562 664954
rect 303646 664718 303882 664954
rect 303326 664398 303562 664634
rect 303646 664398 303882 664634
rect 303326 628718 303562 628954
rect 303646 628718 303882 628954
rect 303326 628398 303562 628634
rect 303646 628398 303882 628634
rect 303326 592718 303562 592954
rect 303646 592718 303882 592954
rect 303326 592398 303562 592634
rect 303646 592398 303882 592634
rect 303326 556718 303562 556954
rect 303646 556718 303882 556954
rect 303326 556398 303562 556634
rect 303646 556398 303882 556634
rect 303326 520718 303562 520954
rect 303646 520718 303882 520954
rect 303326 520398 303562 520634
rect 303646 520398 303882 520634
rect 303326 484718 303562 484954
rect 303646 484718 303882 484954
rect 303326 484398 303562 484634
rect 303646 484398 303882 484634
rect 303326 448718 303562 448954
rect 303646 448718 303882 448954
rect 303326 448398 303562 448634
rect 303646 448398 303882 448634
rect 303326 412718 303562 412954
rect 303646 412718 303882 412954
rect 303326 412398 303562 412634
rect 303646 412398 303882 412634
rect 303326 376718 303562 376954
rect 303646 376718 303882 376954
rect 303326 376398 303562 376634
rect 303646 376398 303882 376634
rect 303326 340718 303562 340954
rect 303646 340718 303882 340954
rect 303326 340398 303562 340634
rect 303646 340398 303882 340634
rect 303326 304718 303562 304954
rect 303646 304718 303882 304954
rect 303326 304398 303562 304634
rect 303646 304398 303882 304634
rect 303326 268718 303562 268954
rect 303646 268718 303882 268954
rect 303326 268398 303562 268634
rect 303646 268398 303882 268634
rect 303326 232718 303562 232954
rect 303646 232718 303882 232954
rect 303326 232398 303562 232634
rect 303646 232398 303882 232634
rect 303326 196718 303562 196954
rect 303646 196718 303882 196954
rect 303326 196398 303562 196634
rect 303646 196398 303882 196634
rect 303326 160718 303562 160954
rect 303646 160718 303882 160954
rect 303326 160398 303562 160634
rect 303646 160398 303882 160634
rect 303326 124718 303562 124954
rect 303646 124718 303882 124954
rect 303326 124398 303562 124634
rect 303646 124398 303882 124634
rect 303326 88718 303562 88954
rect 303646 88718 303882 88954
rect 303326 88398 303562 88634
rect 303646 88398 303882 88634
rect 303326 52718 303562 52954
rect 303646 52718 303882 52954
rect 303326 52398 303562 52634
rect 303646 52398 303882 52634
rect 303326 16718 303562 16954
rect 303646 16718 303882 16954
rect 303326 16398 303562 16634
rect 303646 16398 303882 16634
rect 303326 -3462 303562 -3226
rect 303646 -3462 303882 -3226
rect 303326 -3782 303562 -3546
rect 303646 -3782 303882 -3546
rect 307826 708442 308062 708678
rect 308146 708442 308382 708678
rect 307826 708122 308062 708358
rect 308146 708122 308382 708358
rect 307826 669218 308062 669454
rect 308146 669218 308382 669454
rect 307826 668898 308062 669134
rect 308146 668898 308382 669134
rect 307826 633218 308062 633454
rect 308146 633218 308382 633454
rect 307826 632898 308062 633134
rect 308146 632898 308382 633134
rect 307826 597218 308062 597454
rect 308146 597218 308382 597454
rect 307826 596898 308062 597134
rect 308146 596898 308382 597134
rect 307826 561218 308062 561454
rect 308146 561218 308382 561454
rect 307826 560898 308062 561134
rect 308146 560898 308382 561134
rect 307826 525218 308062 525454
rect 308146 525218 308382 525454
rect 307826 524898 308062 525134
rect 308146 524898 308382 525134
rect 307826 489218 308062 489454
rect 308146 489218 308382 489454
rect 307826 488898 308062 489134
rect 308146 488898 308382 489134
rect 307826 453218 308062 453454
rect 308146 453218 308382 453454
rect 307826 452898 308062 453134
rect 308146 452898 308382 453134
rect 307826 417218 308062 417454
rect 308146 417218 308382 417454
rect 307826 416898 308062 417134
rect 308146 416898 308382 417134
rect 307826 381218 308062 381454
rect 308146 381218 308382 381454
rect 307826 380898 308062 381134
rect 308146 380898 308382 381134
rect 307826 345218 308062 345454
rect 308146 345218 308382 345454
rect 307826 344898 308062 345134
rect 308146 344898 308382 345134
rect 307826 309218 308062 309454
rect 308146 309218 308382 309454
rect 307826 308898 308062 309134
rect 308146 308898 308382 309134
rect 307826 273218 308062 273454
rect 308146 273218 308382 273454
rect 307826 272898 308062 273134
rect 308146 272898 308382 273134
rect 307826 237218 308062 237454
rect 308146 237218 308382 237454
rect 307826 236898 308062 237134
rect 308146 236898 308382 237134
rect 307826 201218 308062 201454
rect 308146 201218 308382 201454
rect 307826 200898 308062 201134
rect 308146 200898 308382 201134
rect 307826 165218 308062 165454
rect 308146 165218 308382 165454
rect 307826 164898 308062 165134
rect 308146 164898 308382 165134
rect 307826 129218 308062 129454
rect 308146 129218 308382 129454
rect 307826 128898 308062 129134
rect 308146 128898 308382 129134
rect 307826 93218 308062 93454
rect 308146 93218 308382 93454
rect 307826 92898 308062 93134
rect 308146 92898 308382 93134
rect 307826 57218 308062 57454
rect 308146 57218 308382 57454
rect 307826 56898 308062 57134
rect 308146 56898 308382 57134
rect 307826 21218 308062 21454
rect 308146 21218 308382 21454
rect 307826 20898 308062 21134
rect 308146 20898 308382 21134
rect 307826 -4422 308062 -4186
rect 308146 -4422 308382 -4186
rect 307826 -4742 308062 -4506
rect 308146 -4742 308382 -4506
rect 312326 709402 312562 709638
rect 312646 709402 312882 709638
rect 312326 709082 312562 709318
rect 312646 709082 312882 709318
rect 312326 673718 312562 673954
rect 312646 673718 312882 673954
rect 312326 673398 312562 673634
rect 312646 673398 312882 673634
rect 312326 637718 312562 637954
rect 312646 637718 312882 637954
rect 312326 637398 312562 637634
rect 312646 637398 312882 637634
rect 312326 601718 312562 601954
rect 312646 601718 312882 601954
rect 312326 601398 312562 601634
rect 312646 601398 312882 601634
rect 312326 565718 312562 565954
rect 312646 565718 312882 565954
rect 312326 565398 312562 565634
rect 312646 565398 312882 565634
rect 312326 529718 312562 529954
rect 312646 529718 312882 529954
rect 312326 529398 312562 529634
rect 312646 529398 312882 529634
rect 312326 493718 312562 493954
rect 312646 493718 312882 493954
rect 312326 493398 312562 493634
rect 312646 493398 312882 493634
rect 312326 457718 312562 457954
rect 312646 457718 312882 457954
rect 312326 457398 312562 457634
rect 312646 457398 312882 457634
rect 312326 421718 312562 421954
rect 312646 421718 312882 421954
rect 312326 421398 312562 421634
rect 312646 421398 312882 421634
rect 312326 385718 312562 385954
rect 312646 385718 312882 385954
rect 312326 385398 312562 385634
rect 312646 385398 312882 385634
rect 312326 349718 312562 349954
rect 312646 349718 312882 349954
rect 312326 349398 312562 349634
rect 312646 349398 312882 349634
rect 312326 313718 312562 313954
rect 312646 313718 312882 313954
rect 312326 313398 312562 313634
rect 312646 313398 312882 313634
rect 312326 277718 312562 277954
rect 312646 277718 312882 277954
rect 312326 277398 312562 277634
rect 312646 277398 312882 277634
rect 312326 241718 312562 241954
rect 312646 241718 312882 241954
rect 312326 241398 312562 241634
rect 312646 241398 312882 241634
rect 312326 205718 312562 205954
rect 312646 205718 312882 205954
rect 312326 205398 312562 205634
rect 312646 205398 312882 205634
rect 312326 169718 312562 169954
rect 312646 169718 312882 169954
rect 312326 169398 312562 169634
rect 312646 169398 312882 169634
rect 312326 133718 312562 133954
rect 312646 133718 312882 133954
rect 312326 133398 312562 133634
rect 312646 133398 312882 133634
rect 312326 97718 312562 97954
rect 312646 97718 312882 97954
rect 312326 97398 312562 97634
rect 312646 97398 312882 97634
rect 312326 61718 312562 61954
rect 312646 61718 312882 61954
rect 312326 61398 312562 61634
rect 312646 61398 312882 61634
rect 312326 25718 312562 25954
rect 312646 25718 312882 25954
rect 312326 25398 312562 25634
rect 312646 25398 312882 25634
rect 312326 -5382 312562 -5146
rect 312646 -5382 312882 -5146
rect 312326 -5702 312562 -5466
rect 312646 -5702 312882 -5466
rect 316826 710362 317062 710598
rect 317146 710362 317382 710598
rect 316826 710042 317062 710278
rect 317146 710042 317382 710278
rect 316826 678218 317062 678454
rect 317146 678218 317382 678454
rect 316826 677898 317062 678134
rect 317146 677898 317382 678134
rect 316826 642218 317062 642454
rect 317146 642218 317382 642454
rect 316826 641898 317062 642134
rect 317146 641898 317382 642134
rect 316826 606218 317062 606454
rect 317146 606218 317382 606454
rect 316826 605898 317062 606134
rect 317146 605898 317382 606134
rect 316826 570218 317062 570454
rect 317146 570218 317382 570454
rect 316826 569898 317062 570134
rect 317146 569898 317382 570134
rect 316826 534218 317062 534454
rect 317146 534218 317382 534454
rect 316826 533898 317062 534134
rect 317146 533898 317382 534134
rect 316826 498218 317062 498454
rect 317146 498218 317382 498454
rect 316826 497898 317062 498134
rect 317146 497898 317382 498134
rect 316826 462218 317062 462454
rect 317146 462218 317382 462454
rect 316826 461898 317062 462134
rect 317146 461898 317382 462134
rect 316826 426218 317062 426454
rect 317146 426218 317382 426454
rect 316826 425898 317062 426134
rect 317146 425898 317382 426134
rect 316826 390218 317062 390454
rect 317146 390218 317382 390454
rect 316826 389898 317062 390134
rect 317146 389898 317382 390134
rect 316826 354218 317062 354454
rect 317146 354218 317382 354454
rect 316826 353898 317062 354134
rect 317146 353898 317382 354134
rect 316826 318218 317062 318454
rect 317146 318218 317382 318454
rect 316826 317898 317062 318134
rect 317146 317898 317382 318134
rect 316826 282218 317062 282454
rect 317146 282218 317382 282454
rect 316826 281898 317062 282134
rect 317146 281898 317382 282134
rect 316826 246218 317062 246454
rect 317146 246218 317382 246454
rect 316826 245898 317062 246134
rect 317146 245898 317382 246134
rect 316826 210218 317062 210454
rect 317146 210218 317382 210454
rect 316826 209898 317062 210134
rect 317146 209898 317382 210134
rect 316826 174218 317062 174454
rect 317146 174218 317382 174454
rect 316826 173898 317062 174134
rect 317146 173898 317382 174134
rect 316826 138218 317062 138454
rect 317146 138218 317382 138454
rect 316826 137898 317062 138134
rect 317146 137898 317382 138134
rect 316826 102218 317062 102454
rect 317146 102218 317382 102454
rect 316826 101898 317062 102134
rect 317146 101898 317382 102134
rect 316826 66218 317062 66454
rect 317146 66218 317382 66454
rect 316826 65898 317062 66134
rect 317146 65898 317382 66134
rect 316826 30218 317062 30454
rect 317146 30218 317382 30454
rect 316826 29898 317062 30134
rect 317146 29898 317382 30134
rect 316826 -6342 317062 -6106
rect 317146 -6342 317382 -6106
rect 316826 -6662 317062 -6426
rect 317146 -6662 317382 -6426
rect 321326 711322 321562 711558
rect 321646 711322 321882 711558
rect 321326 711002 321562 711238
rect 321646 711002 321882 711238
rect 321326 682718 321562 682954
rect 321646 682718 321882 682954
rect 321326 682398 321562 682634
rect 321646 682398 321882 682634
rect 321326 646718 321562 646954
rect 321646 646718 321882 646954
rect 321326 646398 321562 646634
rect 321646 646398 321882 646634
rect 321326 610718 321562 610954
rect 321646 610718 321882 610954
rect 321326 610398 321562 610634
rect 321646 610398 321882 610634
rect 321326 574718 321562 574954
rect 321646 574718 321882 574954
rect 321326 574398 321562 574634
rect 321646 574398 321882 574634
rect 321326 538718 321562 538954
rect 321646 538718 321882 538954
rect 321326 538398 321562 538634
rect 321646 538398 321882 538634
rect 321326 502718 321562 502954
rect 321646 502718 321882 502954
rect 321326 502398 321562 502634
rect 321646 502398 321882 502634
rect 321326 466718 321562 466954
rect 321646 466718 321882 466954
rect 321326 466398 321562 466634
rect 321646 466398 321882 466634
rect 321326 430718 321562 430954
rect 321646 430718 321882 430954
rect 321326 430398 321562 430634
rect 321646 430398 321882 430634
rect 321326 394718 321562 394954
rect 321646 394718 321882 394954
rect 321326 394398 321562 394634
rect 321646 394398 321882 394634
rect 321326 358718 321562 358954
rect 321646 358718 321882 358954
rect 321326 358398 321562 358634
rect 321646 358398 321882 358634
rect 321326 322718 321562 322954
rect 321646 322718 321882 322954
rect 321326 322398 321562 322634
rect 321646 322398 321882 322634
rect 321326 286718 321562 286954
rect 321646 286718 321882 286954
rect 321326 286398 321562 286634
rect 321646 286398 321882 286634
rect 321326 250718 321562 250954
rect 321646 250718 321882 250954
rect 321326 250398 321562 250634
rect 321646 250398 321882 250634
rect 321326 214718 321562 214954
rect 321646 214718 321882 214954
rect 321326 214398 321562 214634
rect 321646 214398 321882 214634
rect 321326 178718 321562 178954
rect 321646 178718 321882 178954
rect 321326 178398 321562 178634
rect 321646 178398 321882 178634
rect 321326 142718 321562 142954
rect 321646 142718 321882 142954
rect 321326 142398 321562 142634
rect 321646 142398 321882 142634
rect 321326 106718 321562 106954
rect 321646 106718 321882 106954
rect 321326 106398 321562 106634
rect 321646 106398 321882 106634
rect 321326 70718 321562 70954
rect 321646 70718 321882 70954
rect 321326 70398 321562 70634
rect 321646 70398 321882 70634
rect 321326 34718 321562 34954
rect 321646 34718 321882 34954
rect 321326 34398 321562 34634
rect 321646 34398 321882 34634
rect 321326 -7302 321562 -7066
rect 321646 -7302 321882 -7066
rect 321326 -7622 321562 -7386
rect 321646 -7622 321882 -7386
rect 325826 704602 326062 704838
rect 326146 704602 326382 704838
rect 325826 704282 326062 704518
rect 326146 704282 326382 704518
rect 325826 687218 326062 687454
rect 326146 687218 326382 687454
rect 325826 686898 326062 687134
rect 326146 686898 326382 687134
rect 325826 651218 326062 651454
rect 326146 651218 326382 651454
rect 325826 650898 326062 651134
rect 326146 650898 326382 651134
rect 325826 615218 326062 615454
rect 326146 615218 326382 615454
rect 325826 614898 326062 615134
rect 326146 614898 326382 615134
rect 325826 579218 326062 579454
rect 326146 579218 326382 579454
rect 325826 578898 326062 579134
rect 326146 578898 326382 579134
rect 325826 543218 326062 543454
rect 326146 543218 326382 543454
rect 325826 542898 326062 543134
rect 326146 542898 326382 543134
rect 325826 507218 326062 507454
rect 326146 507218 326382 507454
rect 325826 506898 326062 507134
rect 326146 506898 326382 507134
rect 325826 471218 326062 471454
rect 326146 471218 326382 471454
rect 325826 470898 326062 471134
rect 326146 470898 326382 471134
rect 325826 435218 326062 435454
rect 326146 435218 326382 435454
rect 325826 434898 326062 435134
rect 326146 434898 326382 435134
rect 325826 399218 326062 399454
rect 326146 399218 326382 399454
rect 325826 398898 326062 399134
rect 326146 398898 326382 399134
rect 325826 363218 326062 363454
rect 326146 363218 326382 363454
rect 325826 362898 326062 363134
rect 326146 362898 326382 363134
rect 325826 327218 326062 327454
rect 326146 327218 326382 327454
rect 325826 326898 326062 327134
rect 326146 326898 326382 327134
rect 325826 291218 326062 291454
rect 326146 291218 326382 291454
rect 325826 290898 326062 291134
rect 326146 290898 326382 291134
rect 325826 255218 326062 255454
rect 326146 255218 326382 255454
rect 325826 254898 326062 255134
rect 326146 254898 326382 255134
rect 325826 219218 326062 219454
rect 326146 219218 326382 219454
rect 325826 218898 326062 219134
rect 326146 218898 326382 219134
rect 325826 183218 326062 183454
rect 326146 183218 326382 183454
rect 325826 182898 326062 183134
rect 326146 182898 326382 183134
rect 325826 147218 326062 147454
rect 326146 147218 326382 147454
rect 325826 146898 326062 147134
rect 326146 146898 326382 147134
rect 325826 111218 326062 111454
rect 326146 111218 326382 111454
rect 325826 110898 326062 111134
rect 326146 110898 326382 111134
rect 325826 75218 326062 75454
rect 326146 75218 326382 75454
rect 325826 74898 326062 75134
rect 326146 74898 326382 75134
rect 325826 39218 326062 39454
rect 326146 39218 326382 39454
rect 325826 38898 326062 39134
rect 326146 38898 326382 39134
rect 325826 3218 326062 3454
rect 326146 3218 326382 3454
rect 325826 2898 326062 3134
rect 326146 2898 326382 3134
rect 325826 -582 326062 -346
rect 326146 -582 326382 -346
rect 325826 -902 326062 -666
rect 326146 -902 326382 -666
rect 330326 705562 330562 705798
rect 330646 705562 330882 705798
rect 330326 705242 330562 705478
rect 330646 705242 330882 705478
rect 330326 691718 330562 691954
rect 330646 691718 330882 691954
rect 330326 691398 330562 691634
rect 330646 691398 330882 691634
rect 330326 655718 330562 655954
rect 330646 655718 330882 655954
rect 330326 655398 330562 655634
rect 330646 655398 330882 655634
rect 330326 619718 330562 619954
rect 330646 619718 330882 619954
rect 330326 619398 330562 619634
rect 330646 619398 330882 619634
rect 330326 583718 330562 583954
rect 330646 583718 330882 583954
rect 330326 583398 330562 583634
rect 330646 583398 330882 583634
rect 330326 547718 330562 547954
rect 330646 547718 330882 547954
rect 330326 547398 330562 547634
rect 330646 547398 330882 547634
rect 330326 511718 330562 511954
rect 330646 511718 330882 511954
rect 330326 511398 330562 511634
rect 330646 511398 330882 511634
rect 330326 475718 330562 475954
rect 330646 475718 330882 475954
rect 330326 475398 330562 475634
rect 330646 475398 330882 475634
rect 330326 439718 330562 439954
rect 330646 439718 330882 439954
rect 330326 439398 330562 439634
rect 330646 439398 330882 439634
rect 330326 403718 330562 403954
rect 330646 403718 330882 403954
rect 330326 403398 330562 403634
rect 330646 403398 330882 403634
rect 330326 367718 330562 367954
rect 330646 367718 330882 367954
rect 330326 367398 330562 367634
rect 330646 367398 330882 367634
rect 330326 331718 330562 331954
rect 330646 331718 330882 331954
rect 330326 331398 330562 331634
rect 330646 331398 330882 331634
rect 330326 295718 330562 295954
rect 330646 295718 330882 295954
rect 330326 295398 330562 295634
rect 330646 295398 330882 295634
rect 330326 259718 330562 259954
rect 330646 259718 330882 259954
rect 330326 259398 330562 259634
rect 330646 259398 330882 259634
rect 330326 223718 330562 223954
rect 330646 223718 330882 223954
rect 330326 223398 330562 223634
rect 330646 223398 330882 223634
rect 330326 187718 330562 187954
rect 330646 187718 330882 187954
rect 330326 187398 330562 187634
rect 330646 187398 330882 187634
rect 330326 151718 330562 151954
rect 330646 151718 330882 151954
rect 330326 151398 330562 151634
rect 330646 151398 330882 151634
rect 330326 115718 330562 115954
rect 330646 115718 330882 115954
rect 330326 115398 330562 115634
rect 330646 115398 330882 115634
rect 330326 79718 330562 79954
rect 330646 79718 330882 79954
rect 330326 79398 330562 79634
rect 330646 79398 330882 79634
rect 330326 43718 330562 43954
rect 330646 43718 330882 43954
rect 330326 43398 330562 43634
rect 330646 43398 330882 43634
rect 330326 7718 330562 7954
rect 330646 7718 330882 7954
rect 330326 7398 330562 7634
rect 330646 7398 330882 7634
rect 330326 -1542 330562 -1306
rect 330646 -1542 330882 -1306
rect 330326 -1862 330562 -1626
rect 330646 -1862 330882 -1626
rect 334826 706522 335062 706758
rect 335146 706522 335382 706758
rect 334826 706202 335062 706438
rect 335146 706202 335382 706438
rect 334826 696218 335062 696454
rect 335146 696218 335382 696454
rect 334826 695898 335062 696134
rect 335146 695898 335382 696134
rect 334826 660218 335062 660454
rect 335146 660218 335382 660454
rect 334826 659898 335062 660134
rect 335146 659898 335382 660134
rect 334826 624218 335062 624454
rect 335146 624218 335382 624454
rect 334826 623898 335062 624134
rect 335146 623898 335382 624134
rect 334826 588218 335062 588454
rect 335146 588218 335382 588454
rect 334826 587898 335062 588134
rect 335146 587898 335382 588134
rect 334826 552218 335062 552454
rect 335146 552218 335382 552454
rect 334826 551898 335062 552134
rect 335146 551898 335382 552134
rect 334826 516218 335062 516454
rect 335146 516218 335382 516454
rect 334826 515898 335062 516134
rect 335146 515898 335382 516134
rect 334826 480218 335062 480454
rect 335146 480218 335382 480454
rect 334826 479898 335062 480134
rect 335146 479898 335382 480134
rect 334826 444218 335062 444454
rect 335146 444218 335382 444454
rect 334826 443898 335062 444134
rect 335146 443898 335382 444134
rect 334826 408218 335062 408454
rect 335146 408218 335382 408454
rect 334826 407898 335062 408134
rect 335146 407898 335382 408134
rect 334826 372218 335062 372454
rect 335146 372218 335382 372454
rect 334826 371898 335062 372134
rect 335146 371898 335382 372134
rect 334826 336218 335062 336454
rect 335146 336218 335382 336454
rect 334826 335898 335062 336134
rect 335146 335898 335382 336134
rect 334826 300218 335062 300454
rect 335146 300218 335382 300454
rect 334826 299898 335062 300134
rect 335146 299898 335382 300134
rect 334826 264218 335062 264454
rect 335146 264218 335382 264454
rect 334826 263898 335062 264134
rect 335146 263898 335382 264134
rect 334826 228218 335062 228454
rect 335146 228218 335382 228454
rect 334826 227898 335062 228134
rect 335146 227898 335382 228134
rect 334826 192218 335062 192454
rect 335146 192218 335382 192454
rect 334826 191898 335062 192134
rect 335146 191898 335382 192134
rect 334826 156218 335062 156454
rect 335146 156218 335382 156454
rect 334826 155898 335062 156134
rect 335146 155898 335382 156134
rect 334826 120218 335062 120454
rect 335146 120218 335382 120454
rect 334826 119898 335062 120134
rect 335146 119898 335382 120134
rect 334826 84218 335062 84454
rect 335146 84218 335382 84454
rect 334826 83898 335062 84134
rect 335146 83898 335382 84134
rect 334826 48218 335062 48454
rect 335146 48218 335382 48454
rect 334826 47898 335062 48134
rect 335146 47898 335382 48134
rect 334826 12218 335062 12454
rect 335146 12218 335382 12454
rect 334826 11898 335062 12134
rect 335146 11898 335382 12134
rect 334826 -2502 335062 -2266
rect 335146 -2502 335382 -2266
rect 334826 -2822 335062 -2586
rect 335146 -2822 335382 -2586
rect 339326 707482 339562 707718
rect 339646 707482 339882 707718
rect 339326 707162 339562 707398
rect 339646 707162 339882 707398
rect 339326 700718 339562 700954
rect 339646 700718 339882 700954
rect 339326 700398 339562 700634
rect 339646 700398 339882 700634
rect 339326 664718 339562 664954
rect 339646 664718 339882 664954
rect 339326 664398 339562 664634
rect 339646 664398 339882 664634
rect 339326 628718 339562 628954
rect 339646 628718 339882 628954
rect 339326 628398 339562 628634
rect 339646 628398 339882 628634
rect 339326 592718 339562 592954
rect 339646 592718 339882 592954
rect 339326 592398 339562 592634
rect 339646 592398 339882 592634
rect 339326 556718 339562 556954
rect 339646 556718 339882 556954
rect 339326 556398 339562 556634
rect 339646 556398 339882 556634
rect 339326 520718 339562 520954
rect 339646 520718 339882 520954
rect 339326 520398 339562 520634
rect 339646 520398 339882 520634
rect 339326 484718 339562 484954
rect 339646 484718 339882 484954
rect 339326 484398 339562 484634
rect 339646 484398 339882 484634
rect 339326 448718 339562 448954
rect 339646 448718 339882 448954
rect 339326 448398 339562 448634
rect 339646 448398 339882 448634
rect 339326 412718 339562 412954
rect 339646 412718 339882 412954
rect 339326 412398 339562 412634
rect 339646 412398 339882 412634
rect 339326 376718 339562 376954
rect 339646 376718 339882 376954
rect 339326 376398 339562 376634
rect 339646 376398 339882 376634
rect 339326 340718 339562 340954
rect 339646 340718 339882 340954
rect 339326 340398 339562 340634
rect 339646 340398 339882 340634
rect 339326 304718 339562 304954
rect 339646 304718 339882 304954
rect 339326 304398 339562 304634
rect 339646 304398 339882 304634
rect 339326 268718 339562 268954
rect 339646 268718 339882 268954
rect 339326 268398 339562 268634
rect 339646 268398 339882 268634
rect 339326 232718 339562 232954
rect 339646 232718 339882 232954
rect 339326 232398 339562 232634
rect 339646 232398 339882 232634
rect 339326 196718 339562 196954
rect 339646 196718 339882 196954
rect 339326 196398 339562 196634
rect 339646 196398 339882 196634
rect 339326 160718 339562 160954
rect 339646 160718 339882 160954
rect 339326 160398 339562 160634
rect 339646 160398 339882 160634
rect 339326 124718 339562 124954
rect 339646 124718 339882 124954
rect 339326 124398 339562 124634
rect 339646 124398 339882 124634
rect 339326 88718 339562 88954
rect 339646 88718 339882 88954
rect 339326 88398 339562 88634
rect 339646 88398 339882 88634
rect 339326 52718 339562 52954
rect 339646 52718 339882 52954
rect 339326 52398 339562 52634
rect 339646 52398 339882 52634
rect 339326 16718 339562 16954
rect 339646 16718 339882 16954
rect 339326 16398 339562 16634
rect 339646 16398 339882 16634
rect 339326 -3462 339562 -3226
rect 339646 -3462 339882 -3226
rect 339326 -3782 339562 -3546
rect 339646 -3782 339882 -3546
rect 343826 708442 344062 708678
rect 344146 708442 344382 708678
rect 343826 708122 344062 708358
rect 344146 708122 344382 708358
rect 343826 669218 344062 669454
rect 344146 669218 344382 669454
rect 343826 668898 344062 669134
rect 344146 668898 344382 669134
rect 343826 633218 344062 633454
rect 344146 633218 344382 633454
rect 343826 632898 344062 633134
rect 344146 632898 344382 633134
rect 343826 597218 344062 597454
rect 344146 597218 344382 597454
rect 343826 596898 344062 597134
rect 344146 596898 344382 597134
rect 343826 561218 344062 561454
rect 344146 561218 344382 561454
rect 343826 560898 344062 561134
rect 344146 560898 344382 561134
rect 343826 525218 344062 525454
rect 344146 525218 344382 525454
rect 343826 524898 344062 525134
rect 344146 524898 344382 525134
rect 343826 489218 344062 489454
rect 344146 489218 344382 489454
rect 343826 488898 344062 489134
rect 344146 488898 344382 489134
rect 343826 453218 344062 453454
rect 344146 453218 344382 453454
rect 343826 452898 344062 453134
rect 344146 452898 344382 453134
rect 343826 417218 344062 417454
rect 344146 417218 344382 417454
rect 343826 416898 344062 417134
rect 344146 416898 344382 417134
rect 343826 381218 344062 381454
rect 344146 381218 344382 381454
rect 343826 380898 344062 381134
rect 344146 380898 344382 381134
rect 343826 345218 344062 345454
rect 344146 345218 344382 345454
rect 343826 344898 344062 345134
rect 344146 344898 344382 345134
rect 343826 309218 344062 309454
rect 344146 309218 344382 309454
rect 343826 308898 344062 309134
rect 344146 308898 344382 309134
rect 343826 273218 344062 273454
rect 344146 273218 344382 273454
rect 343826 272898 344062 273134
rect 344146 272898 344382 273134
rect 343826 237218 344062 237454
rect 344146 237218 344382 237454
rect 343826 236898 344062 237134
rect 344146 236898 344382 237134
rect 343826 201218 344062 201454
rect 344146 201218 344382 201454
rect 343826 200898 344062 201134
rect 344146 200898 344382 201134
rect 343826 165218 344062 165454
rect 344146 165218 344382 165454
rect 343826 164898 344062 165134
rect 344146 164898 344382 165134
rect 343826 129218 344062 129454
rect 344146 129218 344382 129454
rect 343826 128898 344062 129134
rect 344146 128898 344382 129134
rect 343826 93218 344062 93454
rect 344146 93218 344382 93454
rect 343826 92898 344062 93134
rect 344146 92898 344382 93134
rect 343826 57218 344062 57454
rect 344146 57218 344382 57454
rect 343826 56898 344062 57134
rect 344146 56898 344382 57134
rect 343826 21218 344062 21454
rect 344146 21218 344382 21454
rect 343826 20898 344062 21134
rect 344146 20898 344382 21134
rect 343826 -4422 344062 -4186
rect 344146 -4422 344382 -4186
rect 343826 -4742 344062 -4506
rect 344146 -4742 344382 -4506
rect 348326 709402 348562 709638
rect 348646 709402 348882 709638
rect 348326 709082 348562 709318
rect 348646 709082 348882 709318
rect 348326 673718 348562 673954
rect 348646 673718 348882 673954
rect 348326 673398 348562 673634
rect 348646 673398 348882 673634
rect 348326 637718 348562 637954
rect 348646 637718 348882 637954
rect 348326 637398 348562 637634
rect 348646 637398 348882 637634
rect 348326 601718 348562 601954
rect 348646 601718 348882 601954
rect 348326 601398 348562 601634
rect 348646 601398 348882 601634
rect 348326 565718 348562 565954
rect 348646 565718 348882 565954
rect 348326 565398 348562 565634
rect 348646 565398 348882 565634
rect 348326 529718 348562 529954
rect 348646 529718 348882 529954
rect 348326 529398 348562 529634
rect 348646 529398 348882 529634
rect 348326 493718 348562 493954
rect 348646 493718 348882 493954
rect 348326 493398 348562 493634
rect 348646 493398 348882 493634
rect 348326 457718 348562 457954
rect 348646 457718 348882 457954
rect 348326 457398 348562 457634
rect 348646 457398 348882 457634
rect 348326 421718 348562 421954
rect 348646 421718 348882 421954
rect 348326 421398 348562 421634
rect 348646 421398 348882 421634
rect 348326 385718 348562 385954
rect 348646 385718 348882 385954
rect 348326 385398 348562 385634
rect 348646 385398 348882 385634
rect 348326 349718 348562 349954
rect 348646 349718 348882 349954
rect 348326 349398 348562 349634
rect 348646 349398 348882 349634
rect 348326 313718 348562 313954
rect 348646 313718 348882 313954
rect 348326 313398 348562 313634
rect 348646 313398 348882 313634
rect 348326 277718 348562 277954
rect 348646 277718 348882 277954
rect 348326 277398 348562 277634
rect 348646 277398 348882 277634
rect 348326 241718 348562 241954
rect 348646 241718 348882 241954
rect 348326 241398 348562 241634
rect 348646 241398 348882 241634
rect 348326 205718 348562 205954
rect 348646 205718 348882 205954
rect 348326 205398 348562 205634
rect 348646 205398 348882 205634
rect 348326 169718 348562 169954
rect 348646 169718 348882 169954
rect 348326 169398 348562 169634
rect 348646 169398 348882 169634
rect 348326 133718 348562 133954
rect 348646 133718 348882 133954
rect 348326 133398 348562 133634
rect 348646 133398 348882 133634
rect 348326 97718 348562 97954
rect 348646 97718 348882 97954
rect 348326 97398 348562 97634
rect 348646 97398 348882 97634
rect 348326 61718 348562 61954
rect 348646 61718 348882 61954
rect 348326 61398 348562 61634
rect 348646 61398 348882 61634
rect 348326 25718 348562 25954
rect 348646 25718 348882 25954
rect 348326 25398 348562 25634
rect 348646 25398 348882 25634
rect 348326 -5382 348562 -5146
rect 348646 -5382 348882 -5146
rect 348326 -5702 348562 -5466
rect 348646 -5702 348882 -5466
rect 352826 710362 353062 710598
rect 353146 710362 353382 710598
rect 352826 710042 353062 710278
rect 353146 710042 353382 710278
rect 352826 678218 353062 678454
rect 353146 678218 353382 678454
rect 352826 677898 353062 678134
rect 353146 677898 353382 678134
rect 352826 642218 353062 642454
rect 353146 642218 353382 642454
rect 352826 641898 353062 642134
rect 353146 641898 353382 642134
rect 352826 606218 353062 606454
rect 353146 606218 353382 606454
rect 352826 605898 353062 606134
rect 353146 605898 353382 606134
rect 352826 570218 353062 570454
rect 353146 570218 353382 570454
rect 352826 569898 353062 570134
rect 353146 569898 353382 570134
rect 352826 534218 353062 534454
rect 353146 534218 353382 534454
rect 352826 533898 353062 534134
rect 353146 533898 353382 534134
rect 352826 498218 353062 498454
rect 353146 498218 353382 498454
rect 352826 497898 353062 498134
rect 353146 497898 353382 498134
rect 352826 462218 353062 462454
rect 353146 462218 353382 462454
rect 352826 461898 353062 462134
rect 353146 461898 353382 462134
rect 352826 426218 353062 426454
rect 353146 426218 353382 426454
rect 352826 425898 353062 426134
rect 353146 425898 353382 426134
rect 352826 390218 353062 390454
rect 353146 390218 353382 390454
rect 352826 389898 353062 390134
rect 353146 389898 353382 390134
rect 352826 354218 353062 354454
rect 353146 354218 353382 354454
rect 352826 353898 353062 354134
rect 353146 353898 353382 354134
rect 352826 318218 353062 318454
rect 353146 318218 353382 318454
rect 352826 317898 353062 318134
rect 353146 317898 353382 318134
rect 352826 282218 353062 282454
rect 353146 282218 353382 282454
rect 352826 281898 353062 282134
rect 353146 281898 353382 282134
rect 352826 246218 353062 246454
rect 353146 246218 353382 246454
rect 352826 245898 353062 246134
rect 353146 245898 353382 246134
rect 352826 210218 353062 210454
rect 353146 210218 353382 210454
rect 352826 209898 353062 210134
rect 353146 209898 353382 210134
rect 352826 174218 353062 174454
rect 353146 174218 353382 174454
rect 352826 173898 353062 174134
rect 353146 173898 353382 174134
rect 352826 138218 353062 138454
rect 353146 138218 353382 138454
rect 352826 137898 353062 138134
rect 353146 137898 353382 138134
rect 352826 102218 353062 102454
rect 353146 102218 353382 102454
rect 352826 101898 353062 102134
rect 353146 101898 353382 102134
rect 352826 66218 353062 66454
rect 353146 66218 353382 66454
rect 352826 65898 353062 66134
rect 353146 65898 353382 66134
rect 352826 30218 353062 30454
rect 353146 30218 353382 30454
rect 352826 29898 353062 30134
rect 353146 29898 353382 30134
rect 352826 -6342 353062 -6106
rect 353146 -6342 353382 -6106
rect 352826 -6662 353062 -6426
rect 353146 -6662 353382 -6426
rect 357326 711322 357562 711558
rect 357646 711322 357882 711558
rect 357326 711002 357562 711238
rect 357646 711002 357882 711238
rect 357326 682718 357562 682954
rect 357646 682718 357882 682954
rect 357326 682398 357562 682634
rect 357646 682398 357882 682634
rect 357326 646718 357562 646954
rect 357646 646718 357882 646954
rect 357326 646398 357562 646634
rect 357646 646398 357882 646634
rect 357326 610718 357562 610954
rect 357646 610718 357882 610954
rect 357326 610398 357562 610634
rect 357646 610398 357882 610634
rect 357326 574718 357562 574954
rect 357646 574718 357882 574954
rect 357326 574398 357562 574634
rect 357646 574398 357882 574634
rect 357326 538718 357562 538954
rect 357646 538718 357882 538954
rect 357326 538398 357562 538634
rect 357646 538398 357882 538634
rect 357326 502718 357562 502954
rect 357646 502718 357882 502954
rect 357326 502398 357562 502634
rect 357646 502398 357882 502634
rect 357326 466718 357562 466954
rect 357646 466718 357882 466954
rect 357326 466398 357562 466634
rect 357646 466398 357882 466634
rect 357326 430718 357562 430954
rect 357646 430718 357882 430954
rect 357326 430398 357562 430634
rect 357646 430398 357882 430634
rect 357326 394718 357562 394954
rect 357646 394718 357882 394954
rect 357326 394398 357562 394634
rect 357646 394398 357882 394634
rect 357326 358718 357562 358954
rect 357646 358718 357882 358954
rect 357326 358398 357562 358634
rect 357646 358398 357882 358634
rect 357326 322718 357562 322954
rect 357646 322718 357882 322954
rect 357326 322398 357562 322634
rect 357646 322398 357882 322634
rect 357326 286718 357562 286954
rect 357646 286718 357882 286954
rect 357326 286398 357562 286634
rect 357646 286398 357882 286634
rect 357326 250718 357562 250954
rect 357646 250718 357882 250954
rect 357326 250398 357562 250634
rect 357646 250398 357882 250634
rect 357326 214718 357562 214954
rect 357646 214718 357882 214954
rect 357326 214398 357562 214634
rect 357646 214398 357882 214634
rect 357326 178718 357562 178954
rect 357646 178718 357882 178954
rect 357326 178398 357562 178634
rect 357646 178398 357882 178634
rect 357326 142718 357562 142954
rect 357646 142718 357882 142954
rect 357326 142398 357562 142634
rect 357646 142398 357882 142634
rect 357326 106718 357562 106954
rect 357646 106718 357882 106954
rect 357326 106398 357562 106634
rect 357646 106398 357882 106634
rect 357326 70718 357562 70954
rect 357646 70718 357882 70954
rect 357326 70398 357562 70634
rect 357646 70398 357882 70634
rect 357326 34718 357562 34954
rect 357646 34718 357882 34954
rect 357326 34398 357562 34634
rect 357646 34398 357882 34634
rect 357326 -7302 357562 -7066
rect 357646 -7302 357882 -7066
rect 357326 -7622 357562 -7386
rect 357646 -7622 357882 -7386
rect 361826 704602 362062 704838
rect 362146 704602 362382 704838
rect 361826 704282 362062 704518
rect 362146 704282 362382 704518
rect 361826 687218 362062 687454
rect 362146 687218 362382 687454
rect 361826 686898 362062 687134
rect 362146 686898 362382 687134
rect 361826 651218 362062 651454
rect 362146 651218 362382 651454
rect 361826 650898 362062 651134
rect 362146 650898 362382 651134
rect 361826 615218 362062 615454
rect 362146 615218 362382 615454
rect 361826 614898 362062 615134
rect 362146 614898 362382 615134
rect 361826 579218 362062 579454
rect 362146 579218 362382 579454
rect 361826 578898 362062 579134
rect 362146 578898 362382 579134
rect 361826 543218 362062 543454
rect 362146 543218 362382 543454
rect 361826 542898 362062 543134
rect 362146 542898 362382 543134
rect 361826 507218 362062 507454
rect 362146 507218 362382 507454
rect 361826 506898 362062 507134
rect 362146 506898 362382 507134
rect 361826 471218 362062 471454
rect 362146 471218 362382 471454
rect 361826 470898 362062 471134
rect 362146 470898 362382 471134
rect 361826 435218 362062 435454
rect 362146 435218 362382 435454
rect 361826 434898 362062 435134
rect 362146 434898 362382 435134
rect 361826 399218 362062 399454
rect 362146 399218 362382 399454
rect 361826 398898 362062 399134
rect 362146 398898 362382 399134
rect 361826 363218 362062 363454
rect 362146 363218 362382 363454
rect 361826 362898 362062 363134
rect 362146 362898 362382 363134
rect 361826 327218 362062 327454
rect 362146 327218 362382 327454
rect 361826 326898 362062 327134
rect 362146 326898 362382 327134
rect 361826 291218 362062 291454
rect 362146 291218 362382 291454
rect 361826 290898 362062 291134
rect 362146 290898 362382 291134
rect 361826 255218 362062 255454
rect 362146 255218 362382 255454
rect 361826 254898 362062 255134
rect 362146 254898 362382 255134
rect 361826 219218 362062 219454
rect 362146 219218 362382 219454
rect 361826 218898 362062 219134
rect 362146 218898 362382 219134
rect 361826 183218 362062 183454
rect 362146 183218 362382 183454
rect 361826 182898 362062 183134
rect 362146 182898 362382 183134
rect 361826 147218 362062 147454
rect 362146 147218 362382 147454
rect 361826 146898 362062 147134
rect 362146 146898 362382 147134
rect 361826 111218 362062 111454
rect 362146 111218 362382 111454
rect 361826 110898 362062 111134
rect 362146 110898 362382 111134
rect 361826 75218 362062 75454
rect 362146 75218 362382 75454
rect 361826 74898 362062 75134
rect 362146 74898 362382 75134
rect 361826 39218 362062 39454
rect 362146 39218 362382 39454
rect 361826 38898 362062 39134
rect 362146 38898 362382 39134
rect 361826 3218 362062 3454
rect 362146 3218 362382 3454
rect 361826 2898 362062 3134
rect 362146 2898 362382 3134
rect 361826 -582 362062 -346
rect 362146 -582 362382 -346
rect 361826 -902 362062 -666
rect 362146 -902 362382 -666
rect 366326 705562 366562 705798
rect 366646 705562 366882 705798
rect 366326 705242 366562 705478
rect 366646 705242 366882 705478
rect 366326 691718 366562 691954
rect 366646 691718 366882 691954
rect 366326 691398 366562 691634
rect 366646 691398 366882 691634
rect 366326 655718 366562 655954
rect 366646 655718 366882 655954
rect 366326 655398 366562 655634
rect 366646 655398 366882 655634
rect 366326 619718 366562 619954
rect 366646 619718 366882 619954
rect 366326 619398 366562 619634
rect 366646 619398 366882 619634
rect 366326 583718 366562 583954
rect 366646 583718 366882 583954
rect 366326 583398 366562 583634
rect 366646 583398 366882 583634
rect 366326 547718 366562 547954
rect 366646 547718 366882 547954
rect 366326 547398 366562 547634
rect 366646 547398 366882 547634
rect 366326 511718 366562 511954
rect 366646 511718 366882 511954
rect 366326 511398 366562 511634
rect 366646 511398 366882 511634
rect 366326 475718 366562 475954
rect 366646 475718 366882 475954
rect 366326 475398 366562 475634
rect 366646 475398 366882 475634
rect 366326 439718 366562 439954
rect 366646 439718 366882 439954
rect 366326 439398 366562 439634
rect 366646 439398 366882 439634
rect 366326 403718 366562 403954
rect 366646 403718 366882 403954
rect 366326 403398 366562 403634
rect 366646 403398 366882 403634
rect 366326 367718 366562 367954
rect 366646 367718 366882 367954
rect 366326 367398 366562 367634
rect 366646 367398 366882 367634
rect 366326 331718 366562 331954
rect 366646 331718 366882 331954
rect 366326 331398 366562 331634
rect 366646 331398 366882 331634
rect 366326 295718 366562 295954
rect 366646 295718 366882 295954
rect 366326 295398 366562 295634
rect 366646 295398 366882 295634
rect 366326 259718 366562 259954
rect 366646 259718 366882 259954
rect 366326 259398 366562 259634
rect 366646 259398 366882 259634
rect 366326 223718 366562 223954
rect 366646 223718 366882 223954
rect 366326 223398 366562 223634
rect 366646 223398 366882 223634
rect 366326 187718 366562 187954
rect 366646 187718 366882 187954
rect 366326 187398 366562 187634
rect 366646 187398 366882 187634
rect 366326 151718 366562 151954
rect 366646 151718 366882 151954
rect 366326 151398 366562 151634
rect 366646 151398 366882 151634
rect 366326 115718 366562 115954
rect 366646 115718 366882 115954
rect 366326 115398 366562 115634
rect 366646 115398 366882 115634
rect 366326 79718 366562 79954
rect 366646 79718 366882 79954
rect 366326 79398 366562 79634
rect 366646 79398 366882 79634
rect 366326 43718 366562 43954
rect 366646 43718 366882 43954
rect 366326 43398 366562 43634
rect 366646 43398 366882 43634
rect 366326 7718 366562 7954
rect 366646 7718 366882 7954
rect 366326 7398 366562 7634
rect 366646 7398 366882 7634
rect 366326 -1542 366562 -1306
rect 366646 -1542 366882 -1306
rect 366326 -1862 366562 -1626
rect 366646 -1862 366882 -1626
rect 370826 706522 371062 706758
rect 371146 706522 371382 706758
rect 370826 706202 371062 706438
rect 371146 706202 371382 706438
rect 370826 696218 371062 696454
rect 371146 696218 371382 696454
rect 370826 695898 371062 696134
rect 371146 695898 371382 696134
rect 370826 660218 371062 660454
rect 371146 660218 371382 660454
rect 370826 659898 371062 660134
rect 371146 659898 371382 660134
rect 370826 624218 371062 624454
rect 371146 624218 371382 624454
rect 370826 623898 371062 624134
rect 371146 623898 371382 624134
rect 370826 588218 371062 588454
rect 371146 588218 371382 588454
rect 370826 587898 371062 588134
rect 371146 587898 371382 588134
rect 370826 552218 371062 552454
rect 371146 552218 371382 552454
rect 370826 551898 371062 552134
rect 371146 551898 371382 552134
rect 370826 516218 371062 516454
rect 371146 516218 371382 516454
rect 370826 515898 371062 516134
rect 371146 515898 371382 516134
rect 370826 480218 371062 480454
rect 371146 480218 371382 480454
rect 370826 479898 371062 480134
rect 371146 479898 371382 480134
rect 370826 444218 371062 444454
rect 371146 444218 371382 444454
rect 370826 443898 371062 444134
rect 371146 443898 371382 444134
rect 370826 408218 371062 408454
rect 371146 408218 371382 408454
rect 370826 407898 371062 408134
rect 371146 407898 371382 408134
rect 370826 372218 371062 372454
rect 371146 372218 371382 372454
rect 370826 371898 371062 372134
rect 371146 371898 371382 372134
rect 370826 336218 371062 336454
rect 371146 336218 371382 336454
rect 370826 335898 371062 336134
rect 371146 335898 371382 336134
rect 370826 300218 371062 300454
rect 371146 300218 371382 300454
rect 370826 299898 371062 300134
rect 371146 299898 371382 300134
rect 370826 264218 371062 264454
rect 371146 264218 371382 264454
rect 370826 263898 371062 264134
rect 371146 263898 371382 264134
rect 370826 228218 371062 228454
rect 371146 228218 371382 228454
rect 370826 227898 371062 228134
rect 371146 227898 371382 228134
rect 370826 192218 371062 192454
rect 371146 192218 371382 192454
rect 370826 191898 371062 192134
rect 371146 191898 371382 192134
rect 370826 156218 371062 156454
rect 371146 156218 371382 156454
rect 370826 155898 371062 156134
rect 371146 155898 371382 156134
rect 370826 120218 371062 120454
rect 371146 120218 371382 120454
rect 370826 119898 371062 120134
rect 371146 119898 371382 120134
rect 370826 84218 371062 84454
rect 371146 84218 371382 84454
rect 370826 83898 371062 84134
rect 371146 83898 371382 84134
rect 370826 48218 371062 48454
rect 371146 48218 371382 48454
rect 370826 47898 371062 48134
rect 371146 47898 371382 48134
rect 370826 12218 371062 12454
rect 371146 12218 371382 12454
rect 370826 11898 371062 12134
rect 371146 11898 371382 12134
rect 370826 -2502 371062 -2266
rect 371146 -2502 371382 -2266
rect 370826 -2822 371062 -2586
rect 371146 -2822 371382 -2586
rect 375326 707482 375562 707718
rect 375646 707482 375882 707718
rect 375326 707162 375562 707398
rect 375646 707162 375882 707398
rect 375326 700718 375562 700954
rect 375646 700718 375882 700954
rect 375326 700398 375562 700634
rect 375646 700398 375882 700634
rect 375326 664718 375562 664954
rect 375646 664718 375882 664954
rect 375326 664398 375562 664634
rect 375646 664398 375882 664634
rect 375326 628718 375562 628954
rect 375646 628718 375882 628954
rect 375326 628398 375562 628634
rect 375646 628398 375882 628634
rect 375326 592718 375562 592954
rect 375646 592718 375882 592954
rect 375326 592398 375562 592634
rect 375646 592398 375882 592634
rect 375326 556718 375562 556954
rect 375646 556718 375882 556954
rect 375326 556398 375562 556634
rect 375646 556398 375882 556634
rect 375326 520718 375562 520954
rect 375646 520718 375882 520954
rect 375326 520398 375562 520634
rect 375646 520398 375882 520634
rect 375326 484718 375562 484954
rect 375646 484718 375882 484954
rect 375326 484398 375562 484634
rect 375646 484398 375882 484634
rect 375326 448718 375562 448954
rect 375646 448718 375882 448954
rect 375326 448398 375562 448634
rect 375646 448398 375882 448634
rect 375326 412718 375562 412954
rect 375646 412718 375882 412954
rect 375326 412398 375562 412634
rect 375646 412398 375882 412634
rect 375326 376718 375562 376954
rect 375646 376718 375882 376954
rect 375326 376398 375562 376634
rect 375646 376398 375882 376634
rect 375326 340718 375562 340954
rect 375646 340718 375882 340954
rect 375326 340398 375562 340634
rect 375646 340398 375882 340634
rect 375326 304718 375562 304954
rect 375646 304718 375882 304954
rect 375326 304398 375562 304634
rect 375646 304398 375882 304634
rect 375326 268718 375562 268954
rect 375646 268718 375882 268954
rect 375326 268398 375562 268634
rect 375646 268398 375882 268634
rect 375326 232718 375562 232954
rect 375646 232718 375882 232954
rect 375326 232398 375562 232634
rect 375646 232398 375882 232634
rect 375326 196718 375562 196954
rect 375646 196718 375882 196954
rect 375326 196398 375562 196634
rect 375646 196398 375882 196634
rect 375326 160718 375562 160954
rect 375646 160718 375882 160954
rect 375326 160398 375562 160634
rect 375646 160398 375882 160634
rect 375326 124718 375562 124954
rect 375646 124718 375882 124954
rect 375326 124398 375562 124634
rect 375646 124398 375882 124634
rect 375326 88718 375562 88954
rect 375646 88718 375882 88954
rect 375326 88398 375562 88634
rect 375646 88398 375882 88634
rect 375326 52718 375562 52954
rect 375646 52718 375882 52954
rect 375326 52398 375562 52634
rect 375646 52398 375882 52634
rect 375326 16718 375562 16954
rect 375646 16718 375882 16954
rect 375326 16398 375562 16634
rect 375646 16398 375882 16634
rect 375326 -3462 375562 -3226
rect 375646 -3462 375882 -3226
rect 375326 -3782 375562 -3546
rect 375646 -3782 375882 -3546
rect 379826 708442 380062 708678
rect 380146 708442 380382 708678
rect 379826 708122 380062 708358
rect 380146 708122 380382 708358
rect 379826 669218 380062 669454
rect 380146 669218 380382 669454
rect 379826 668898 380062 669134
rect 380146 668898 380382 669134
rect 379826 633218 380062 633454
rect 380146 633218 380382 633454
rect 379826 632898 380062 633134
rect 380146 632898 380382 633134
rect 379826 597218 380062 597454
rect 380146 597218 380382 597454
rect 379826 596898 380062 597134
rect 380146 596898 380382 597134
rect 379826 561218 380062 561454
rect 380146 561218 380382 561454
rect 379826 560898 380062 561134
rect 380146 560898 380382 561134
rect 379826 525218 380062 525454
rect 380146 525218 380382 525454
rect 379826 524898 380062 525134
rect 380146 524898 380382 525134
rect 379826 489218 380062 489454
rect 380146 489218 380382 489454
rect 379826 488898 380062 489134
rect 380146 488898 380382 489134
rect 379826 453218 380062 453454
rect 380146 453218 380382 453454
rect 379826 452898 380062 453134
rect 380146 452898 380382 453134
rect 379826 417218 380062 417454
rect 380146 417218 380382 417454
rect 379826 416898 380062 417134
rect 380146 416898 380382 417134
rect 379826 381218 380062 381454
rect 380146 381218 380382 381454
rect 379826 380898 380062 381134
rect 380146 380898 380382 381134
rect 379826 345218 380062 345454
rect 380146 345218 380382 345454
rect 379826 344898 380062 345134
rect 380146 344898 380382 345134
rect 379826 309218 380062 309454
rect 380146 309218 380382 309454
rect 379826 308898 380062 309134
rect 380146 308898 380382 309134
rect 379826 273218 380062 273454
rect 380146 273218 380382 273454
rect 379826 272898 380062 273134
rect 380146 272898 380382 273134
rect 379826 237218 380062 237454
rect 380146 237218 380382 237454
rect 379826 236898 380062 237134
rect 380146 236898 380382 237134
rect 379826 201218 380062 201454
rect 380146 201218 380382 201454
rect 379826 200898 380062 201134
rect 380146 200898 380382 201134
rect 379826 165218 380062 165454
rect 380146 165218 380382 165454
rect 379826 164898 380062 165134
rect 380146 164898 380382 165134
rect 379826 129218 380062 129454
rect 380146 129218 380382 129454
rect 379826 128898 380062 129134
rect 380146 128898 380382 129134
rect 379826 93218 380062 93454
rect 380146 93218 380382 93454
rect 379826 92898 380062 93134
rect 380146 92898 380382 93134
rect 379826 57218 380062 57454
rect 380146 57218 380382 57454
rect 379826 56898 380062 57134
rect 380146 56898 380382 57134
rect 379826 21218 380062 21454
rect 380146 21218 380382 21454
rect 379826 20898 380062 21134
rect 380146 20898 380382 21134
rect 379826 -4422 380062 -4186
rect 380146 -4422 380382 -4186
rect 379826 -4742 380062 -4506
rect 380146 -4742 380382 -4506
rect 384326 709402 384562 709638
rect 384646 709402 384882 709638
rect 384326 709082 384562 709318
rect 384646 709082 384882 709318
rect 384326 673718 384562 673954
rect 384646 673718 384882 673954
rect 384326 673398 384562 673634
rect 384646 673398 384882 673634
rect 384326 637718 384562 637954
rect 384646 637718 384882 637954
rect 384326 637398 384562 637634
rect 384646 637398 384882 637634
rect 384326 601718 384562 601954
rect 384646 601718 384882 601954
rect 384326 601398 384562 601634
rect 384646 601398 384882 601634
rect 384326 565718 384562 565954
rect 384646 565718 384882 565954
rect 384326 565398 384562 565634
rect 384646 565398 384882 565634
rect 384326 529718 384562 529954
rect 384646 529718 384882 529954
rect 384326 529398 384562 529634
rect 384646 529398 384882 529634
rect 384326 493718 384562 493954
rect 384646 493718 384882 493954
rect 384326 493398 384562 493634
rect 384646 493398 384882 493634
rect 384326 457718 384562 457954
rect 384646 457718 384882 457954
rect 384326 457398 384562 457634
rect 384646 457398 384882 457634
rect 384326 421718 384562 421954
rect 384646 421718 384882 421954
rect 384326 421398 384562 421634
rect 384646 421398 384882 421634
rect 384326 385718 384562 385954
rect 384646 385718 384882 385954
rect 384326 385398 384562 385634
rect 384646 385398 384882 385634
rect 384326 349718 384562 349954
rect 384646 349718 384882 349954
rect 384326 349398 384562 349634
rect 384646 349398 384882 349634
rect 384326 313718 384562 313954
rect 384646 313718 384882 313954
rect 384326 313398 384562 313634
rect 384646 313398 384882 313634
rect 384326 277718 384562 277954
rect 384646 277718 384882 277954
rect 384326 277398 384562 277634
rect 384646 277398 384882 277634
rect 384326 241718 384562 241954
rect 384646 241718 384882 241954
rect 384326 241398 384562 241634
rect 384646 241398 384882 241634
rect 384326 205718 384562 205954
rect 384646 205718 384882 205954
rect 384326 205398 384562 205634
rect 384646 205398 384882 205634
rect 384326 169718 384562 169954
rect 384646 169718 384882 169954
rect 384326 169398 384562 169634
rect 384646 169398 384882 169634
rect 384326 133718 384562 133954
rect 384646 133718 384882 133954
rect 384326 133398 384562 133634
rect 384646 133398 384882 133634
rect 384326 97718 384562 97954
rect 384646 97718 384882 97954
rect 384326 97398 384562 97634
rect 384646 97398 384882 97634
rect 384326 61718 384562 61954
rect 384646 61718 384882 61954
rect 384326 61398 384562 61634
rect 384646 61398 384882 61634
rect 384326 25718 384562 25954
rect 384646 25718 384882 25954
rect 384326 25398 384562 25634
rect 384646 25398 384882 25634
rect 384326 -5382 384562 -5146
rect 384646 -5382 384882 -5146
rect 384326 -5702 384562 -5466
rect 384646 -5702 384882 -5466
rect 388826 710362 389062 710598
rect 389146 710362 389382 710598
rect 388826 710042 389062 710278
rect 389146 710042 389382 710278
rect 388826 678218 389062 678454
rect 389146 678218 389382 678454
rect 388826 677898 389062 678134
rect 389146 677898 389382 678134
rect 388826 642218 389062 642454
rect 389146 642218 389382 642454
rect 388826 641898 389062 642134
rect 389146 641898 389382 642134
rect 388826 606218 389062 606454
rect 389146 606218 389382 606454
rect 388826 605898 389062 606134
rect 389146 605898 389382 606134
rect 388826 570218 389062 570454
rect 389146 570218 389382 570454
rect 388826 569898 389062 570134
rect 389146 569898 389382 570134
rect 388826 534218 389062 534454
rect 389146 534218 389382 534454
rect 388826 533898 389062 534134
rect 389146 533898 389382 534134
rect 388826 498218 389062 498454
rect 389146 498218 389382 498454
rect 388826 497898 389062 498134
rect 389146 497898 389382 498134
rect 388826 462218 389062 462454
rect 389146 462218 389382 462454
rect 388826 461898 389062 462134
rect 389146 461898 389382 462134
rect 388826 426218 389062 426454
rect 389146 426218 389382 426454
rect 388826 425898 389062 426134
rect 389146 425898 389382 426134
rect 388826 390218 389062 390454
rect 389146 390218 389382 390454
rect 388826 389898 389062 390134
rect 389146 389898 389382 390134
rect 388826 354218 389062 354454
rect 389146 354218 389382 354454
rect 388826 353898 389062 354134
rect 389146 353898 389382 354134
rect 388826 318218 389062 318454
rect 389146 318218 389382 318454
rect 388826 317898 389062 318134
rect 389146 317898 389382 318134
rect 388826 282218 389062 282454
rect 389146 282218 389382 282454
rect 388826 281898 389062 282134
rect 389146 281898 389382 282134
rect 388826 246218 389062 246454
rect 389146 246218 389382 246454
rect 388826 245898 389062 246134
rect 389146 245898 389382 246134
rect 388826 210218 389062 210454
rect 389146 210218 389382 210454
rect 388826 209898 389062 210134
rect 389146 209898 389382 210134
rect 388826 174218 389062 174454
rect 389146 174218 389382 174454
rect 388826 173898 389062 174134
rect 389146 173898 389382 174134
rect 388826 138218 389062 138454
rect 389146 138218 389382 138454
rect 388826 137898 389062 138134
rect 389146 137898 389382 138134
rect 388826 102218 389062 102454
rect 389146 102218 389382 102454
rect 388826 101898 389062 102134
rect 389146 101898 389382 102134
rect 388826 66218 389062 66454
rect 389146 66218 389382 66454
rect 388826 65898 389062 66134
rect 389146 65898 389382 66134
rect 388826 30218 389062 30454
rect 389146 30218 389382 30454
rect 388826 29898 389062 30134
rect 389146 29898 389382 30134
rect 388826 -6342 389062 -6106
rect 389146 -6342 389382 -6106
rect 388826 -6662 389062 -6426
rect 389146 -6662 389382 -6426
rect 393326 711322 393562 711558
rect 393646 711322 393882 711558
rect 393326 711002 393562 711238
rect 393646 711002 393882 711238
rect 393326 682718 393562 682954
rect 393646 682718 393882 682954
rect 393326 682398 393562 682634
rect 393646 682398 393882 682634
rect 393326 646718 393562 646954
rect 393646 646718 393882 646954
rect 393326 646398 393562 646634
rect 393646 646398 393882 646634
rect 393326 610718 393562 610954
rect 393646 610718 393882 610954
rect 393326 610398 393562 610634
rect 393646 610398 393882 610634
rect 393326 574718 393562 574954
rect 393646 574718 393882 574954
rect 393326 574398 393562 574634
rect 393646 574398 393882 574634
rect 393326 538718 393562 538954
rect 393646 538718 393882 538954
rect 393326 538398 393562 538634
rect 393646 538398 393882 538634
rect 393326 502718 393562 502954
rect 393646 502718 393882 502954
rect 393326 502398 393562 502634
rect 393646 502398 393882 502634
rect 393326 466718 393562 466954
rect 393646 466718 393882 466954
rect 393326 466398 393562 466634
rect 393646 466398 393882 466634
rect 393326 430718 393562 430954
rect 393646 430718 393882 430954
rect 393326 430398 393562 430634
rect 393646 430398 393882 430634
rect 393326 394718 393562 394954
rect 393646 394718 393882 394954
rect 393326 394398 393562 394634
rect 393646 394398 393882 394634
rect 393326 358718 393562 358954
rect 393646 358718 393882 358954
rect 393326 358398 393562 358634
rect 393646 358398 393882 358634
rect 393326 322718 393562 322954
rect 393646 322718 393882 322954
rect 393326 322398 393562 322634
rect 393646 322398 393882 322634
rect 393326 286718 393562 286954
rect 393646 286718 393882 286954
rect 393326 286398 393562 286634
rect 393646 286398 393882 286634
rect 393326 250718 393562 250954
rect 393646 250718 393882 250954
rect 393326 250398 393562 250634
rect 393646 250398 393882 250634
rect 393326 214718 393562 214954
rect 393646 214718 393882 214954
rect 393326 214398 393562 214634
rect 393646 214398 393882 214634
rect 393326 178718 393562 178954
rect 393646 178718 393882 178954
rect 393326 178398 393562 178634
rect 393646 178398 393882 178634
rect 393326 142718 393562 142954
rect 393646 142718 393882 142954
rect 393326 142398 393562 142634
rect 393646 142398 393882 142634
rect 393326 106718 393562 106954
rect 393646 106718 393882 106954
rect 393326 106398 393562 106634
rect 393646 106398 393882 106634
rect 393326 70718 393562 70954
rect 393646 70718 393882 70954
rect 393326 70398 393562 70634
rect 393646 70398 393882 70634
rect 393326 34718 393562 34954
rect 393646 34718 393882 34954
rect 393326 34398 393562 34634
rect 393646 34398 393882 34634
rect 393326 -7302 393562 -7066
rect 393646 -7302 393882 -7066
rect 393326 -7622 393562 -7386
rect 393646 -7622 393882 -7386
rect 397826 704602 398062 704838
rect 398146 704602 398382 704838
rect 397826 704282 398062 704518
rect 398146 704282 398382 704518
rect 397826 687218 398062 687454
rect 398146 687218 398382 687454
rect 397826 686898 398062 687134
rect 398146 686898 398382 687134
rect 397826 651218 398062 651454
rect 398146 651218 398382 651454
rect 397826 650898 398062 651134
rect 398146 650898 398382 651134
rect 397826 615218 398062 615454
rect 398146 615218 398382 615454
rect 397826 614898 398062 615134
rect 398146 614898 398382 615134
rect 397826 579218 398062 579454
rect 398146 579218 398382 579454
rect 397826 578898 398062 579134
rect 398146 578898 398382 579134
rect 397826 543218 398062 543454
rect 398146 543218 398382 543454
rect 397826 542898 398062 543134
rect 398146 542898 398382 543134
rect 397826 507218 398062 507454
rect 398146 507218 398382 507454
rect 397826 506898 398062 507134
rect 398146 506898 398382 507134
rect 397826 471218 398062 471454
rect 398146 471218 398382 471454
rect 397826 470898 398062 471134
rect 398146 470898 398382 471134
rect 397826 435218 398062 435454
rect 398146 435218 398382 435454
rect 397826 434898 398062 435134
rect 398146 434898 398382 435134
rect 397826 399218 398062 399454
rect 398146 399218 398382 399454
rect 397826 398898 398062 399134
rect 398146 398898 398382 399134
rect 397826 363218 398062 363454
rect 398146 363218 398382 363454
rect 397826 362898 398062 363134
rect 398146 362898 398382 363134
rect 397826 327218 398062 327454
rect 398146 327218 398382 327454
rect 397826 326898 398062 327134
rect 398146 326898 398382 327134
rect 397826 291218 398062 291454
rect 398146 291218 398382 291454
rect 397826 290898 398062 291134
rect 398146 290898 398382 291134
rect 397826 255218 398062 255454
rect 398146 255218 398382 255454
rect 397826 254898 398062 255134
rect 398146 254898 398382 255134
rect 397826 219218 398062 219454
rect 398146 219218 398382 219454
rect 397826 218898 398062 219134
rect 398146 218898 398382 219134
rect 397826 183218 398062 183454
rect 398146 183218 398382 183454
rect 397826 182898 398062 183134
rect 398146 182898 398382 183134
rect 397826 147218 398062 147454
rect 398146 147218 398382 147454
rect 397826 146898 398062 147134
rect 398146 146898 398382 147134
rect 397826 111218 398062 111454
rect 398146 111218 398382 111454
rect 397826 110898 398062 111134
rect 398146 110898 398382 111134
rect 397826 75218 398062 75454
rect 398146 75218 398382 75454
rect 397826 74898 398062 75134
rect 398146 74898 398382 75134
rect 397826 39218 398062 39454
rect 398146 39218 398382 39454
rect 397826 38898 398062 39134
rect 398146 38898 398382 39134
rect 397826 3218 398062 3454
rect 398146 3218 398382 3454
rect 397826 2898 398062 3134
rect 398146 2898 398382 3134
rect 397826 -582 398062 -346
rect 398146 -582 398382 -346
rect 397826 -902 398062 -666
rect 398146 -902 398382 -666
rect 402326 705562 402562 705798
rect 402646 705562 402882 705798
rect 402326 705242 402562 705478
rect 402646 705242 402882 705478
rect 402326 691718 402562 691954
rect 402646 691718 402882 691954
rect 402326 691398 402562 691634
rect 402646 691398 402882 691634
rect 402326 655718 402562 655954
rect 402646 655718 402882 655954
rect 402326 655398 402562 655634
rect 402646 655398 402882 655634
rect 402326 619718 402562 619954
rect 402646 619718 402882 619954
rect 402326 619398 402562 619634
rect 402646 619398 402882 619634
rect 402326 583718 402562 583954
rect 402646 583718 402882 583954
rect 402326 583398 402562 583634
rect 402646 583398 402882 583634
rect 402326 547718 402562 547954
rect 402646 547718 402882 547954
rect 402326 547398 402562 547634
rect 402646 547398 402882 547634
rect 402326 511718 402562 511954
rect 402646 511718 402882 511954
rect 402326 511398 402562 511634
rect 402646 511398 402882 511634
rect 402326 475718 402562 475954
rect 402646 475718 402882 475954
rect 402326 475398 402562 475634
rect 402646 475398 402882 475634
rect 402326 439718 402562 439954
rect 402646 439718 402882 439954
rect 402326 439398 402562 439634
rect 402646 439398 402882 439634
rect 402326 403718 402562 403954
rect 402646 403718 402882 403954
rect 402326 403398 402562 403634
rect 402646 403398 402882 403634
rect 402326 367718 402562 367954
rect 402646 367718 402882 367954
rect 402326 367398 402562 367634
rect 402646 367398 402882 367634
rect 402326 331718 402562 331954
rect 402646 331718 402882 331954
rect 402326 331398 402562 331634
rect 402646 331398 402882 331634
rect 402326 295718 402562 295954
rect 402646 295718 402882 295954
rect 402326 295398 402562 295634
rect 402646 295398 402882 295634
rect 402326 259718 402562 259954
rect 402646 259718 402882 259954
rect 402326 259398 402562 259634
rect 402646 259398 402882 259634
rect 402326 223718 402562 223954
rect 402646 223718 402882 223954
rect 402326 223398 402562 223634
rect 402646 223398 402882 223634
rect 402326 187718 402562 187954
rect 402646 187718 402882 187954
rect 402326 187398 402562 187634
rect 402646 187398 402882 187634
rect 402326 151718 402562 151954
rect 402646 151718 402882 151954
rect 402326 151398 402562 151634
rect 402646 151398 402882 151634
rect 402326 115718 402562 115954
rect 402646 115718 402882 115954
rect 402326 115398 402562 115634
rect 402646 115398 402882 115634
rect 402326 79718 402562 79954
rect 402646 79718 402882 79954
rect 402326 79398 402562 79634
rect 402646 79398 402882 79634
rect 402326 43718 402562 43954
rect 402646 43718 402882 43954
rect 402326 43398 402562 43634
rect 402646 43398 402882 43634
rect 402326 7718 402562 7954
rect 402646 7718 402882 7954
rect 402326 7398 402562 7634
rect 402646 7398 402882 7634
rect 402326 -1542 402562 -1306
rect 402646 -1542 402882 -1306
rect 402326 -1862 402562 -1626
rect 402646 -1862 402882 -1626
rect 406826 706522 407062 706758
rect 407146 706522 407382 706758
rect 406826 706202 407062 706438
rect 407146 706202 407382 706438
rect 406826 696218 407062 696454
rect 407146 696218 407382 696454
rect 406826 695898 407062 696134
rect 407146 695898 407382 696134
rect 406826 660218 407062 660454
rect 407146 660218 407382 660454
rect 406826 659898 407062 660134
rect 407146 659898 407382 660134
rect 406826 624218 407062 624454
rect 407146 624218 407382 624454
rect 406826 623898 407062 624134
rect 407146 623898 407382 624134
rect 406826 588218 407062 588454
rect 407146 588218 407382 588454
rect 406826 587898 407062 588134
rect 407146 587898 407382 588134
rect 406826 552218 407062 552454
rect 407146 552218 407382 552454
rect 406826 551898 407062 552134
rect 407146 551898 407382 552134
rect 406826 516218 407062 516454
rect 407146 516218 407382 516454
rect 406826 515898 407062 516134
rect 407146 515898 407382 516134
rect 406826 480218 407062 480454
rect 407146 480218 407382 480454
rect 406826 479898 407062 480134
rect 407146 479898 407382 480134
rect 406826 444218 407062 444454
rect 407146 444218 407382 444454
rect 406826 443898 407062 444134
rect 407146 443898 407382 444134
rect 406826 408218 407062 408454
rect 407146 408218 407382 408454
rect 406826 407898 407062 408134
rect 407146 407898 407382 408134
rect 406826 372218 407062 372454
rect 407146 372218 407382 372454
rect 406826 371898 407062 372134
rect 407146 371898 407382 372134
rect 406826 336218 407062 336454
rect 407146 336218 407382 336454
rect 406826 335898 407062 336134
rect 407146 335898 407382 336134
rect 406826 300218 407062 300454
rect 407146 300218 407382 300454
rect 406826 299898 407062 300134
rect 407146 299898 407382 300134
rect 406826 264218 407062 264454
rect 407146 264218 407382 264454
rect 406826 263898 407062 264134
rect 407146 263898 407382 264134
rect 406826 228218 407062 228454
rect 407146 228218 407382 228454
rect 406826 227898 407062 228134
rect 407146 227898 407382 228134
rect 406826 192218 407062 192454
rect 407146 192218 407382 192454
rect 406826 191898 407062 192134
rect 407146 191898 407382 192134
rect 406826 156218 407062 156454
rect 407146 156218 407382 156454
rect 406826 155898 407062 156134
rect 407146 155898 407382 156134
rect 406826 120218 407062 120454
rect 407146 120218 407382 120454
rect 406826 119898 407062 120134
rect 407146 119898 407382 120134
rect 406826 84218 407062 84454
rect 407146 84218 407382 84454
rect 406826 83898 407062 84134
rect 407146 83898 407382 84134
rect 406826 48218 407062 48454
rect 407146 48218 407382 48454
rect 406826 47898 407062 48134
rect 407146 47898 407382 48134
rect 406826 12218 407062 12454
rect 407146 12218 407382 12454
rect 406826 11898 407062 12134
rect 407146 11898 407382 12134
rect 406826 -2502 407062 -2266
rect 407146 -2502 407382 -2266
rect 406826 -2822 407062 -2586
rect 407146 -2822 407382 -2586
rect 411326 707482 411562 707718
rect 411646 707482 411882 707718
rect 411326 707162 411562 707398
rect 411646 707162 411882 707398
rect 411326 700718 411562 700954
rect 411646 700718 411882 700954
rect 411326 700398 411562 700634
rect 411646 700398 411882 700634
rect 411326 664718 411562 664954
rect 411646 664718 411882 664954
rect 411326 664398 411562 664634
rect 411646 664398 411882 664634
rect 411326 628718 411562 628954
rect 411646 628718 411882 628954
rect 411326 628398 411562 628634
rect 411646 628398 411882 628634
rect 411326 592718 411562 592954
rect 411646 592718 411882 592954
rect 411326 592398 411562 592634
rect 411646 592398 411882 592634
rect 411326 556718 411562 556954
rect 411646 556718 411882 556954
rect 411326 556398 411562 556634
rect 411646 556398 411882 556634
rect 411326 520718 411562 520954
rect 411646 520718 411882 520954
rect 411326 520398 411562 520634
rect 411646 520398 411882 520634
rect 411326 484718 411562 484954
rect 411646 484718 411882 484954
rect 411326 484398 411562 484634
rect 411646 484398 411882 484634
rect 411326 448718 411562 448954
rect 411646 448718 411882 448954
rect 411326 448398 411562 448634
rect 411646 448398 411882 448634
rect 411326 412718 411562 412954
rect 411646 412718 411882 412954
rect 411326 412398 411562 412634
rect 411646 412398 411882 412634
rect 411326 376718 411562 376954
rect 411646 376718 411882 376954
rect 411326 376398 411562 376634
rect 411646 376398 411882 376634
rect 411326 340718 411562 340954
rect 411646 340718 411882 340954
rect 411326 340398 411562 340634
rect 411646 340398 411882 340634
rect 411326 304718 411562 304954
rect 411646 304718 411882 304954
rect 411326 304398 411562 304634
rect 411646 304398 411882 304634
rect 411326 268718 411562 268954
rect 411646 268718 411882 268954
rect 411326 268398 411562 268634
rect 411646 268398 411882 268634
rect 411326 232718 411562 232954
rect 411646 232718 411882 232954
rect 411326 232398 411562 232634
rect 411646 232398 411882 232634
rect 411326 196718 411562 196954
rect 411646 196718 411882 196954
rect 411326 196398 411562 196634
rect 411646 196398 411882 196634
rect 411326 160718 411562 160954
rect 411646 160718 411882 160954
rect 411326 160398 411562 160634
rect 411646 160398 411882 160634
rect 411326 124718 411562 124954
rect 411646 124718 411882 124954
rect 411326 124398 411562 124634
rect 411646 124398 411882 124634
rect 411326 88718 411562 88954
rect 411646 88718 411882 88954
rect 411326 88398 411562 88634
rect 411646 88398 411882 88634
rect 411326 52718 411562 52954
rect 411646 52718 411882 52954
rect 411326 52398 411562 52634
rect 411646 52398 411882 52634
rect 411326 16718 411562 16954
rect 411646 16718 411882 16954
rect 411326 16398 411562 16634
rect 411646 16398 411882 16634
rect 411326 -3462 411562 -3226
rect 411646 -3462 411882 -3226
rect 411326 -3782 411562 -3546
rect 411646 -3782 411882 -3546
rect 415826 708442 416062 708678
rect 416146 708442 416382 708678
rect 415826 708122 416062 708358
rect 416146 708122 416382 708358
rect 415826 669218 416062 669454
rect 416146 669218 416382 669454
rect 415826 668898 416062 669134
rect 416146 668898 416382 669134
rect 415826 633218 416062 633454
rect 416146 633218 416382 633454
rect 415826 632898 416062 633134
rect 416146 632898 416382 633134
rect 415826 597218 416062 597454
rect 416146 597218 416382 597454
rect 415826 596898 416062 597134
rect 416146 596898 416382 597134
rect 415826 561218 416062 561454
rect 416146 561218 416382 561454
rect 415826 560898 416062 561134
rect 416146 560898 416382 561134
rect 415826 525218 416062 525454
rect 416146 525218 416382 525454
rect 415826 524898 416062 525134
rect 416146 524898 416382 525134
rect 415826 489218 416062 489454
rect 416146 489218 416382 489454
rect 415826 488898 416062 489134
rect 416146 488898 416382 489134
rect 415826 453218 416062 453454
rect 416146 453218 416382 453454
rect 415826 452898 416062 453134
rect 416146 452898 416382 453134
rect 415826 417218 416062 417454
rect 416146 417218 416382 417454
rect 415826 416898 416062 417134
rect 416146 416898 416382 417134
rect 415826 381218 416062 381454
rect 416146 381218 416382 381454
rect 415826 380898 416062 381134
rect 416146 380898 416382 381134
rect 415826 345218 416062 345454
rect 416146 345218 416382 345454
rect 415826 344898 416062 345134
rect 416146 344898 416382 345134
rect 415826 309218 416062 309454
rect 416146 309218 416382 309454
rect 415826 308898 416062 309134
rect 416146 308898 416382 309134
rect 415826 273218 416062 273454
rect 416146 273218 416382 273454
rect 415826 272898 416062 273134
rect 416146 272898 416382 273134
rect 415826 237218 416062 237454
rect 416146 237218 416382 237454
rect 415826 236898 416062 237134
rect 416146 236898 416382 237134
rect 415826 201218 416062 201454
rect 416146 201218 416382 201454
rect 415826 200898 416062 201134
rect 416146 200898 416382 201134
rect 415826 165218 416062 165454
rect 416146 165218 416382 165454
rect 415826 164898 416062 165134
rect 416146 164898 416382 165134
rect 415826 129218 416062 129454
rect 416146 129218 416382 129454
rect 415826 128898 416062 129134
rect 416146 128898 416382 129134
rect 415826 93218 416062 93454
rect 416146 93218 416382 93454
rect 415826 92898 416062 93134
rect 416146 92898 416382 93134
rect 415826 57218 416062 57454
rect 416146 57218 416382 57454
rect 415826 56898 416062 57134
rect 416146 56898 416382 57134
rect 415826 21218 416062 21454
rect 416146 21218 416382 21454
rect 415826 20898 416062 21134
rect 416146 20898 416382 21134
rect 415826 -4422 416062 -4186
rect 416146 -4422 416382 -4186
rect 415826 -4742 416062 -4506
rect 416146 -4742 416382 -4506
rect 420326 709402 420562 709638
rect 420646 709402 420882 709638
rect 420326 709082 420562 709318
rect 420646 709082 420882 709318
rect 420326 673718 420562 673954
rect 420646 673718 420882 673954
rect 420326 673398 420562 673634
rect 420646 673398 420882 673634
rect 420326 637718 420562 637954
rect 420646 637718 420882 637954
rect 420326 637398 420562 637634
rect 420646 637398 420882 637634
rect 420326 601718 420562 601954
rect 420646 601718 420882 601954
rect 420326 601398 420562 601634
rect 420646 601398 420882 601634
rect 420326 565718 420562 565954
rect 420646 565718 420882 565954
rect 420326 565398 420562 565634
rect 420646 565398 420882 565634
rect 420326 529718 420562 529954
rect 420646 529718 420882 529954
rect 420326 529398 420562 529634
rect 420646 529398 420882 529634
rect 420326 493718 420562 493954
rect 420646 493718 420882 493954
rect 420326 493398 420562 493634
rect 420646 493398 420882 493634
rect 420326 457718 420562 457954
rect 420646 457718 420882 457954
rect 420326 457398 420562 457634
rect 420646 457398 420882 457634
rect 420326 421718 420562 421954
rect 420646 421718 420882 421954
rect 420326 421398 420562 421634
rect 420646 421398 420882 421634
rect 420326 385718 420562 385954
rect 420646 385718 420882 385954
rect 420326 385398 420562 385634
rect 420646 385398 420882 385634
rect 420326 349718 420562 349954
rect 420646 349718 420882 349954
rect 420326 349398 420562 349634
rect 420646 349398 420882 349634
rect 420326 313718 420562 313954
rect 420646 313718 420882 313954
rect 420326 313398 420562 313634
rect 420646 313398 420882 313634
rect 420326 277718 420562 277954
rect 420646 277718 420882 277954
rect 420326 277398 420562 277634
rect 420646 277398 420882 277634
rect 420326 241718 420562 241954
rect 420646 241718 420882 241954
rect 420326 241398 420562 241634
rect 420646 241398 420882 241634
rect 420326 205718 420562 205954
rect 420646 205718 420882 205954
rect 420326 205398 420562 205634
rect 420646 205398 420882 205634
rect 420326 169718 420562 169954
rect 420646 169718 420882 169954
rect 420326 169398 420562 169634
rect 420646 169398 420882 169634
rect 420326 133718 420562 133954
rect 420646 133718 420882 133954
rect 420326 133398 420562 133634
rect 420646 133398 420882 133634
rect 420326 97718 420562 97954
rect 420646 97718 420882 97954
rect 420326 97398 420562 97634
rect 420646 97398 420882 97634
rect 420326 61718 420562 61954
rect 420646 61718 420882 61954
rect 420326 61398 420562 61634
rect 420646 61398 420882 61634
rect 420326 25718 420562 25954
rect 420646 25718 420882 25954
rect 420326 25398 420562 25634
rect 420646 25398 420882 25634
rect 420326 -5382 420562 -5146
rect 420646 -5382 420882 -5146
rect 420326 -5702 420562 -5466
rect 420646 -5702 420882 -5466
rect 424826 710362 425062 710598
rect 425146 710362 425382 710598
rect 424826 710042 425062 710278
rect 425146 710042 425382 710278
rect 424826 678218 425062 678454
rect 425146 678218 425382 678454
rect 424826 677898 425062 678134
rect 425146 677898 425382 678134
rect 424826 642218 425062 642454
rect 425146 642218 425382 642454
rect 424826 641898 425062 642134
rect 425146 641898 425382 642134
rect 424826 606218 425062 606454
rect 425146 606218 425382 606454
rect 424826 605898 425062 606134
rect 425146 605898 425382 606134
rect 424826 570218 425062 570454
rect 425146 570218 425382 570454
rect 424826 569898 425062 570134
rect 425146 569898 425382 570134
rect 424826 534218 425062 534454
rect 425146 534218 425382 534454
rect 424826 533898 425062 534134
rect 425146 533898 425382 534134
rect 424826 498218 425062 498454
rect 425146 498218 425382 498454
rect 424826 497898 425062 498134
rect 425146 497898 425382 498134
rect 424826 462218 425062 462454
rect 425146 462218 425382 462454
rect 424826 461898 425062 462134
rect 425146 461898 425382 462134
rect 424826 426218 425062 426454
rect 425146 426218 425382 426454
rect 424826 425898 425062 426134
rect 425146 425898 425382 426134
rect 424826 390218 425062 390454
rect 425146 390218 425382 390454
rect 424826 389898 425062 390134
rect 425146 389898 425382 390134
rect 424826 354218 425062 354454
rect 425146 354218 425382 354454
rect 424826 353898 425062 354134
rect 425146 353898 425382 354134
rect 424826 318218 425062 318454
rect 425146 318218 425382 318454
rect 424826 317898 425062 318134
rect 425146 317898 425382 318134
rect 424826 282218 425062 282454
rect 425146 282218 425382 282454
rect 424826 281898 425062 282134
rect 425146 281898 425382 282134
rect 424826 246218 425062 246454
rect 425146 246218 425382 246454
rect 424826 245898 425062 246134
rect 425146 245898 425382 246134
rect 424826 210218 425062 210454
rect 425146 210218 425382 210454
rect 424826 209898 425062 210134
rect 425146 209898 425382 210134
rect 424826 174218 425062 174454
rect 425146 174218 425382 174454
rect 424826 173898 425062 174134
rect 425146 173898 425382 174134
rect 424826 138218 425062 138454
rect 425146 138218 425382 138454
rect 424826 137898 425062 138134
rect 425146 137898 425382 138134
rect 424826 102218 425062 102454
rect 425146 102218 425382 102454
rect 424826 101898 425062 102134
rect 425146 101898 425382 102134
rect 424826 66218 425062 66454
rect 425146 66218 425382 66454
rect 424826 65898 425062 66134
rect 425146 65898 425382 66134
rect 424826 30218 425062 30454
rect 425146 30218 425382 30454
rect 424826 29898 425062 30134
rect 425146 29898 425382 30134
rect 424826 -6342 425062 -6106
rect 425146 -6342 425382 -6106
rect 424826 -6662 425062 -6426
rect 425146 -6662 425382 -6426
rect 429326 711322 429562 711558
rect 429646 711322 429882 711558
rect 429326 711002 429562 711238
rect 429646 711002 429882 711238
rect 429326 682718 429562 682954
rect 429646 682718 429882 682954
rect 429326 682398 429562 682634
rect 429646 682398 429882 682634
rect 429326 646718 429562 646954
rect 429646 646718 429882 646954
rect 429326 646398 429562 646634
rect 429646 646398 429882 646634
rect 429326 610718 429562 610954
rect 429646 610718 429882 610954
rect 429326 610398 429562 610634
rect 429646 610398 429882 610634
rect 429326 574718 429562 574954
rect 429646 574718 429882 574954
rect 429326 574398 429562 574634
rect 429646 574398 429882 574634
rect 429326 538718 429562 538954
rect 429646 538718 429882 538954
rect 429326 538398 429562 538634
rect 429646 538398 429882 538634
rect 429326 502718 429562 502954
rect 429646 502718 429882 502954
rect 429326 502398 429562 502634
rect 429646 502398 429882 502634
rect 429326 466718 429562 466954
rect 429646 466718 429882 466954
rect 429326 466398 429562 466634
rect 429646 466398 429882 466634
rect 429326 430718 429562 430954
rect 429646 430718 429882 430954
rect 429326 430398 429562 430634
rect 429646 430398 429882 430634
rect 429326 394718 429562 394954
rect 429646 394718 429882 394954
rect 429326 394398 429562 394634
rect 429646 394398 429882 394634
rect 429326 358718 429562 358954
rect 429646 358718 429882 358954
rect 429326 358398 429562 358634
rect 429646 358398 429882 358634
rect 429326 322718 429562 322954
rect 429646 322718 429882 322954
rect 429326 322398 429562 322634
rect 429646 322398 429882 322634
rect 429326 286718 429562 286954
rect 429646 286718 429882 286954
rect 429326 286398 429562 286634
rect 429646 286398 429882 286634
rect 429326 250718 429562 250954
rect 429646 250718 429882 250954
rect 429326 250398 429562 250634
rect 429646 250398 429882 250634
rect 429326 214718 429562 214954
rect 429646 214718 429882 214954
rect 429326 214398 429562 214634
rect 429646 214398 429882 214634
rect 429326 178718 429562 178954
rect 429646 178718 429882 178954
rect 429326 178398 429562 178634
rect 429646 178398 429882 178634
rect 429326 142718 429562 142954
rect 429646 142718 429882 142954
rect 429326 142398 429562 142634
rect 429646 142398 429882 142634
rect 429326 106718 429562 106954
rect 429646 106718 429882 106954
rect 429326 106398 429562 106634
rect 429646 106398 429882 106634
rect 429326 70718 429562 70954
rect 429646 70718 429882 70954
rect 429326 70398 429562 70634
rect 429646 70398 429882 70634
rect 429326 34718 429562 34954
rect 429646 34718 429882 34954
rect 429326 34398 429562 34634
rect 429646 34398 429882 34634
rect 429326 -7302 429562 -7066
rect 429646 -7302 429882 -7066
rect 429326 -7622 429562 -7386
rect 429646 -7622 429882 -7386
rect 433826 704602 434062 704838
rect 434146 704602 434382 704838
rect 433826 704282 434062 704518
rect 434146 704282 434382 704518
rect 433826 687218 434062 687454
rect 434146 687218 434382 687454
rect 433826 686898 434062 687134
rect 434146 686898 434382 687134
rect 433826 651218 434062 651454
rect 434146 651218 434382 651454
rect 433826 650898 434062 651134
rect 434146 650898 434382 651134
rect 433826 615218 434062 615454
rect 434146 615218 434382 615454
rect 433826 614898 434062 615134
rect 434146 614898 434382 615134
rect 433826 579218 434062 579454
rect 434146 579218 434382 579454
rect 433826 578898 434062 579134
rect 434146 578898 434382 579134
rect 433826 543218 434062 543454
rect 434146 543218 434382 543454
rect 433826 542898 434062 543134
rect 434146 542898 434382 543134
rect 433826 507218 434062 507454
rect 434146 507218 434382 507454
rect 433826 506898 434062 507134
rect 434146 506898 434382 507134
rect 433826 471218 434062 471454
rect 434146 471218 434382 471454
rect 433826 470898 434062 471134
rect 434146 470898 434382 471134
rect 433826 435218 434062 435454
rect 434146 435218 434382 435454
rect 433826 434898 434062 435134
rect 434146 434898 434382 435134
rect 433826 399218 434062 399454
rect 434146 399218 434382 399454
rect 433826 398898 434062 399134
rect 434146 398898 434382 399134
rect 433826 363218 434062 363454
rect 434146 363218 434382 363454
rect 433826 362898 434062 363134
rect 434146 362898 434382 363134
rect 433826 327218 434062 327454
rect 434146 327218 434382 327454
rect 433826 326898 434062 327134
rect 434146 326898 434382 327134
rect 433826 291218 434062 291454
rect 434146 291218 434382 291454
rect 433826 290898 434062 291134
rect 434146 290898 434382 291134
rect 433826 255218 434062 255454
rect 434146 255218 434382 255454
rect 433826 254898 434062 255134
rect 434146 254898 434382 255134
rect 433826 219218 434062 219454
rect 434146 219218 434382 219454
rect 433826 218898 434062 219134
rect 434146 218898 434382 219134
rect 433826 183218 434062 183454
rect 434146 183218 434382 183454
rect 433826 182898 434062 183134
rect 434146 182898 434382 183134
rect 433826 147218 434062 147454
rect 434146 147218 434382 147454
rect 433826 146898 434062 147134
rect 434146 146898 434382 147134
rect 433826 111218 434062 111454
rect 434146 111218 434382 111454
rect 433826 110898 434062 111134
rect 434146 110898 434382 111134
rect 433826 75218 434062 75454
rect 434146 75218 434382 75454
rect 433826 74898 434062 75134
rect 434146 74898 434382 75134
rect 433826 39218 434062 39454
rect 434146 39218 434382 39454
rect 433826 38898 434062 39134
rect 434146 38898 434382 39134
rect 433826 3218 434062 3454
rect 434146 3218 434382 3454
rect 433826 2898 434062 3134
rect 434146 2898 434382 3134
rect 433826 -582 434062 -346
rect 434146 -582 434382 -346
rect 433826 -902 434062 -666
rect 434146 -902 434382 -666
rect 438326 705562 438562 705798
rect 438646 705562 438882 705798
rect 438326 705242 438562 705478
rect 438646 705242 438882 705478
rect 438326 691718 438562 691954
rect 438646 691718 438882 691954
rect 438326 691398 438562 691634
rect 438646 691398 438882 691634
rect 438326 655718 438562 655954
rect 438646 655718 438882 655954
rect 438326 655398 438562 655634
rect 438646 655398 438882 655634
rect 438326 619718 438562 619954
rect 438646 619718 438882 619954
rect 438326 619398 438562 619634
rect 438646 619398 438882 619634
rect 438326 583718 438562 583954
rect 438646 583718 438882 583954
rect 438326 583398 438562 583634
rect 438646 583398 438882 583634
rect 438326 547718 438562 547954
rect 438646 547718 438882 547954
rect 438326 547398 438562 547634
rect 438646 547398 438882 547634
rect 438326 511718 438562 511954
rect 438646 511718 438882 511954
rect 438326 511398 438562 511634
rect 438646 511398 438882 511634
rect 438326 475718 438562 475954
rect 438646 475718 438882 475954
rect 438326 475398 438562 475634
rect 438646 475398 438882 475634
rect 438326 439718 438562 439954
rect 438646 439718 438882 439954
rect 438326 439398 438562 439634
rect 438646 439398 438882 439634
rect 438326 403718 438562 403954
rect 438646 403718 438882 403954
rect 438326 403398 438562 403634
rect 438646 403398 438882 403634
rect 438326 367718 438562 367954
rect 438646 367718 438882 367954
rect 438326 367398 438562 367634
rect 438646 367398 438882 367634
rect 438326 331718 438562 331954
rect 438646 331718 438882 331954
rect 438326 331398 438562 331634
rect 438646 331398 438882 331634
rect 438326 295718 438562 295954
rect 438646 295718 438882 295954
rect 438326 295398 438562 295634
rect 438646 295398 438882 295634
rect 438326 259718 438562 259954
rect 438646 259718 438882 259954
rect 438326 259398 438562 259634
rect 438646 259398 438882 259634
rect 438326 223718 438562 223954
rect 438646 223718 438882 223954
rect 438326 223398 438562 223634
rect 438646 223398 438882 223634
rect 438326 187718 438562 187954
rect 438646 187718 438882 187954
rect 438326 187398 438562 187634
rect 438646 187398 438882 187634
rect 438326 151718 438562 151954
rect 438646 151718 438882 151954
rect 438326 151398 438562 151634
rect 438646 151398 438882 151634
rect 438326 115718 438562 115954
rect 438646 115718 438882 115954
rect 438326 115398 438562 115634
rect 438646 115398 438882 115634
rect 438326 79718 438562 79954
rect 438646 79718 438882 79954
rect 438326 79398 438562 79634
rect 438646 79398 438882 79634
rect 438326 43718 438562 43954
rect 438646 43718 438882 43954
rect 438326 43398 438562 43634
rect 438646 43398 438882 43634
rect 438326 7718 438562 7954
rect 438646 7718 438882 7954
rect 438326 7398 438562 7634
rect 438646 7398 438882 7634
rect 438326 -1542 438562 -1306
rect 438646 -1542 438882 -1306
rect 438326 -1862 438562 -1626
rect 438646 -1862 438882 -1626
rect 442826 706522 443062 706758
rect 443146 706522 443382 706758
rect 442826 706202 443062 706438
rect 443146 706202 443382 706438
rect 442826 696218 443062 696454
rect 443146 696218 443382 696454
rect 442826 695898 443062 696134
rect 443146 695898 443382 696134
rect 442826 660218 443062 660454
rect 443146 660218 443382 660454
rect 442826 659898 443062 660134
rect 443146 659898 443382 660134
rect 442826 624218 443062 624454
rect 443146 624218 443382 624454
rect 442826 623898 443062 624134
rect 443146 623898 443382 624134
rect 442826 588218 443062 588454
rect 443146 588218 443382 588454
rect 442826 587898 443062 588134
rect 443146 587898 443382 588134
rect 442826 552218 443062 552454
rect 443146 552218 443382 552454
rect 442826 551898 443062 552134
rect 443146 551898 443382 552134
rect 442826 516218 443062 516454
rect 443146 516218 443382 516454
rect 442826 515898 443062 516134
rect 443146 515898 443382 516134
rect 442826 480218 443062 480454
rect 443146 480218 443382 480454
rect 442826 479898 443062 480134
rect 443146 479898 443382 480134
rect 442826 444218 443062 444454
rect 443146 444218 443382 444454
rect 442826 443898 443062 444134
rect 443146 443898 443382 444134
rect 442826 408218 443062 408454
rect 443146 408218 443382 408454
rect 442826 407898 443062 408134
rect 443146 407898 443382 408134
rect 442826 372218 443062 372454
rect 443146 372218 443382 372454
rect 442826 371898 443062 372134
rect 443146 371898 443382 372134
rect 442826 336218 443062 336454
rect 443146 336218 443382 336454
rect 442826 335898 443062 336134
rect 443146 335898 443382 336134
rect 442826 300218 443062 300454
rect 443146 300218 443382 300454
rect 442826 299898 443062 300134
rect 443146 299898 443382 300134
rect 442826 264218 443062 264454
rect 443146 264218 443382 264454
rect 442826 263898 443062 264134
rect 443146 263898 443382 264134
rect 442826 228218 443062 228454
rect 443146 228218 443382 228454
rect 442826 227898 443062 228134
rect 443146 227898 443382 228134
rect 442826 192218 443062 192454
rect 443146 192218 443382 192454
rect 442826 191898 443062 192134
rect 443146 191898 443382 192134
rect 442826 156218 443062 156454
rect 443146 156218 443382 156454
rect 442826 155898 443062 156134
rect 443146 155898 443382 156134
rect 442826 120218 443062 120454
rect 443146 120218 443382 120454
rect 442826 119898 443062 120134
rect 443146 119898 443382 120134
rect 442826 84218 443062 84454
rect 443146 84218 443382 84454
rect 442826 83898 443062 84134
rect 443146 83898 443382 84134
rect 442826 48218 443062 48454
rect 443146 48218 443382 48454
rect 442826 47898 443062 48134
rect 443146 47898 443382 48134
rect 442826 12218 443062 12454
rect 443146 12218 443382 12454
rect 442826 11898 443062 12134
rect 443146 11898 443382 12134
rect 442826 -2502 443062 -2266
rect 443146 -2502 443382 -2266
rect 442826 -2822 443062 -2586
rect 443146 -2822 443382 -2586
rect 447326 707482 447562 707718
rect 447646 707482 447882 707718
rect 447326 707162 447562 707398
rect 447646 707162 447882 707398
rect 447326 700718 447562 700954
rect 447646 700718 447882 700954
rect 447326 700398 447562 700634
rect 447646 700398 447882 700634
rect 447326 664718 447562 664954
rect 447646 664718 447882 664954
rect 447326 664398 447562 664634
rect 447646 664398 447882 664634
rect 447326 628718 447562 628954
rect 447646 628718 447882 628954
rect 447326 628398 447562 628634
rect 447646 628398 447882 628634
rect 447326 592718 447562 592954
rect 447646 592718 447882 592954
rect 447326 592398 447562 592634
rect 447646 592398 447882 592634
rect 447326 556718 447562 556954
rect 447646 556718 447882 556954
rect 447326 556398 447562 556634
rect 447646 556398 447882 556634
rect 447326 520718 447562 520954
rect 447646 520718 447882 520954
rect 447326 520398 447562 520634
rect 447646 520398 447882 520634
rect 447326 484718 447562 484954
rect 447646 484718 447882 484954
rect 447326 484398 447562 484634
rect 447646 484398 447882 484634
rect 447326 448718 447562 448954
rect 447646 448718 447882 448954
rect 447326 448398 447562 448634
rect 447646 448398 447882 448634
rect 447326 412718 447562 412954
rect 447646 412718 447882 412954
rect 447326 412398 447562 412634
rect 447646 412398 447882 412634
rect 447326 376718 447562 376954
rect 447646 376718 447882 376954
rect 447326 376398 447562 376634
rect 447646 376398 447882 376634
rect 447326 340718 447562 340954
rect 447646 340718 447882 340954
rect 447326 340398 447562 340634
rect 447646 340398 447882 340634
rect 447326 304718 447562 304954
rect 447646 304718 447882 304954
rect 447326 304398 447562 304634
rect 447646 304398 447882 304634
rect 447326 268718 447562 268954
rect 447646 268718 447882 268954
rect 447326 268398 447562 268634
rect 447646 268398 447882 268634
rect 447326 232718 447562 232954
rect 447646 232718 447882 232954
rect 447326 232398 447562 232634
rect 447646 232398 447882 232634
rect 447326 196718 447562 196954
rect 447646 196718 447882 196954
rect 447326 196398 447562 196634
rect 447646 196398 447882 196634
rect 447326 160718 447562 160954
rect 447646 160718 447882 160954
rect 447326 160398 447562 160634
rect 447646 160398 447882 160634
rect 447326 124718 447562 124954
rect 447646 124718 447882 124954
rect 447326 124398 447562 124634
rect 447646 124398 447882 124634
rect 447326 88718 447562 88954
rect 447646 88718 447882 88954
rect 447326 88398 447562 88634
rect 447646 88398 447882 88634
rect 447326 52718 447562 52954
rect 447646 52718 447882 52954
rect 447326 52398 447562 52634
rect 447646 52398 447882 52634
rect 447326 16718 447562 16954
rect 447646 16718 447882 16954
rect 447326 16398 447562 16634
rect 447646 16398 447882 16634
rect 447326 -3462 447562 -3226
rect 447646 -3462 447882 -3226
rect 447326 -3782 447562 -3546
rect 447646 -3782 447882 -3546
rect 451826 708442 452062 708678
rect 452146 708442 452382 708678
rect 451826 708122 452062 708358
rect 452146 708122 452382 708358
rect 451826 669218 452062 669454
rect 452146 669218 452382 669454
rect 451826 668898 452062 669134
rect 452146 668898 452382 669134
rect 451826 633218 452062 633454
rect 452146 633218 452382 633454
rect 451826 632898 452062 633134
rect 452146 632898 452382 633134
rect 451826 597218 452062 597454
rect 452146 597218 452382 597454
rect 451826 596898 452062 597134
rect 452146 596898 452382 597134
rect 451826 561218 452062 561454
rect 452146 561218 452382 561454
rect 451826 560898 452062 561134
rect 452146 560898 452382 561134
rect 451826 525218 452062 525454
rect 452146 525218 452382 525454
rect 451826 524898 452062 525134
rect 452146 524898 452382 525134
rect 451826 489218 452062 489454
rect 452146 489218 452382 489454
rect 451826 488898 452062 489134
rect 452146 488898 452382 489134
rect 451826 453218 452062 453454
rect 452146 453218 452382 453454
rect 451826 452898 452062 453134
rect 452146 452898 452382 453134
rect 451826 417218 452062 417454
rect 452146 417218 452382 417454
rect 451826 416898 452062 417134
rect 452146 416898 452382 417134
rect 451826 381218 452062 381454
rect 452146 381218 452382 381454
rect 451826 380898 452062 381134
rect 452146 380898 452382 381134
rect 451826 345218 452062 345454
rect 452146 345218 452382 345454
rect 451826 344898 452062 345134
rect 452146 344898 452382 345134
rect 451826 309218 452062 309454
rect 452146 309218 452382 309454
rect 451826 308898 452062 309134
rect 452146 308898 452382 309134
rect 451826 273218 452062 273454
rect 452146 273218 452382 273454
rect 451826 272898 452062 273134
rect 452146 272898 452382 273134
rect 451826 237218 452062 237454
rect 452146 237218 452382 237454
rect 451826 236898 452062 237134
rect 452146 236898 452382 237134
rect 451826 201218 452062 201454
rect 452146 201218 452382 201454
rect 451826 200898 452062 201134
rect 452146 200898 452382 201134
rect 451826 165218 452062 165454
rect 452146 165218 452382 165454
rect 451826 164898 452062 165134
rect 452146 164898 452382 165134
rect 451826 129218 452062 129454
rect 452146 129218 452382 129454
rect 451826 128898 452062 129134
rect 452146 128898 452382 129134
rect 451826 93218 452062 93454
rect 452146 93218 452382 93454
rect 451826 92898 452062 93134
rect 452146 92898 452382 93134
rect 451826 57218 452062 57454
rect 452146 57218 452382 57454
rect 451826 56898 452062 57134
rect 452146 56898 452382 57134
rect 451826 21218 452062 21454
rect 452146 21218 452382 21454
rect 451826 20898 452062 21134
rect 452146 20898 452382 21134
rect 451826 -4422 452062 -4186
rect 452146 -4422 452382 -4186
rect 451826 -4742 452062 -4506
rect 452146 -4742 452382 -4506
rect 456326 709402 456562 709638
rect 456646 709402 456882 709638
rect 456326 709082 456562 709318
rect 456646 709082 456882 709318
rect 456326 673718 456562 673954
rect 456646 673718 456882 673954
rect 456326 673398 456562 673634
rect 456646 673398 456882 673634
rect 456326 637718 456562 637954
rect 456646 637718 456882 637954
rect 456326 637398 456562 637634
rect 456646 637398 456882 637634
rect 456326 601718 456562 601954
rect 456646 601718 456882 601954
rect 456326 601398 456562 601634
rect 456646 601398 456882 601634
rect 456326 565718 456562 565954
rect 456646 565718 456882 565954
rect 456326 565398 456562 565634
rect 456646 565398 456882 565634
rect 456326 529718 456562 529954
rect 456646 529718 456882 529954
rect 456326 529398 456562 529634
rect 456646 529398 456882 529634
rect 456326 493718 456562 493954
rect 456646 493718 456882 493954
rect 456326 493398 456562 493634
rect 456646 493398 456882 493634
rect 456326 457718 456562 457954
rect 456646 457718 456882 457954
rect 456326 457398 456562 457634
rect 456646 457398 456882 457634
rect 456326 421718 456562 421954
rect 456646 421718 456882 421954
rect 456326 421398 456562 421634
rect 456646 421398 456882 421634
rect 456326 385718 456562 385954
rect 456646 385718 456882 385954
rect 456326 385398 456562 385634
rect 456646 385398 456882 385634
rect 456326 349718 456562 349954
rect 456646 349718 456882 349954
rect 456326 349398 456562 349634
rect 456646 349398 456882 349634
rect 456326 313718 456562 313954
rect 456646 313718 456882 313954
rect 456326 313398 456562 313634
rect 456646 313398 456882 313634
rect 456326 277718 456562 277954
rect 456646 277718 456882 277954
rect 456326 277398 456562 277634
rect 456646 277398 456882 277634
rect 456326 241718 456562 241954
rect 456646 241718 456882 241954
rect 456326 241398 456562 241634
rect 456646 241398 456882 241634
rect 456326 205718 456562 205954
rect 456646 205718 456882 205954
rect 456326 205398 456562 205634
rect 456646 205398 456882 205634
rect 456326 169718 456562 169954
rect 456646 169718 456882 169954
rect 456326 169398 456562 169634
rect 456646 169398 456882 169634
rect 456326 133718 456562 133954
rect 456646 133718 456882 133954
rect 456326 133398 456562 133634
rect 456646 133398 456882 133634
rect 456326 97718 456562 97954
rect 456646 97718 456882 97954
rect 456326 97398 456562 97634
rect 456646 97398 456882 97634
rect 456326 61718 456562 61954
rect 456646 61718 456882 61954
rect 456326 61398 456562 61634
rect 456646 61398 456882 61634
rect 456326 25718 456562 25954
rect 456646 25718 456882 25954
rect 456326 25398 456562 25634
rect 456646 25398 456882 25634
rect 456326 -5382 456562 -5146
rect 456646 -5382 456882 -5146
rect 456326 -5702 456562 -5466
rect 456646 -5702 456882 -5466
rect 460826 710362 461062 710598
rect 461146 710362 461382 710598
rect 460826 710042 461062 710278
rect 461146 710042 461382 710278
rect 460826 678218 461062 678454
rect 461146 678218 461382 678454
rect 460826 677898 461062 678134
rect 461146 677898 461382 678134
rect 460826 642218 461062 642454
rect 461146 642218 461382 642454
rect 460826 641898 461062 642134
rect 461146 641898 461382 642134
rect 460826 606218 461062 606454
rect 461146 606218 461382 606454
rect 460826 605898 461062 606134
rect 461146 605898 461382 606134
rect 460826 570218 461062 570454
rect 461146 570218 461382 570454
rect 460826 569898 461062 570134
rect 461146 569898 461382 570134
rect 460826 534218 461062 534454
rect 461146 534218 461382 534454
rect 460826 533898 461062 534134
rect 461146 533898 461382 534134
rect 460826 498218 461062 498454
rect 461146 498218 461382 498454
rect 460826 497898 461062 498134
rect 461146 497898 461382 498134
rect 460826 462218 461062 462454
rect 461146 462218 461382 462454
rect 460826 461898 461062 462134
rect 461146 461898 461382 462134
rect 460826 426218 461062 426454
rect 461146 426218 461382 426454
rect 460826 425898 461062 426134
rect 461146 425898 461382 426134
rect 460826 390218 461062 390454
rect 461146 390218 461382 390454
rect 460826 389898 461062 390134
rect 461146 389898 461382 390134
rect 460826 354218 461062 354454
rect 461146 354218 461382 354454
rect 460826 353898 461062 354134
rect 461146 353898 461382 354134
rect 460826 318218 461062 318454
rect 461146 318218 461382 318454
rect 460826 317898 461062 318134
rect 461146 317898 461382 318134
rect 460826 282218 461062 282454
rect 461146 282218 461382 282454
rect 460826 281898 461062 282134
rect 461146 281898 461382 282134
rect 460826 246218 461062 246454
rect 461146 246218 461382 246454
rect 460826 245898 461062 246134
rect 461146 245898 461382 246134
rect 460826 210218 461062 210454
rect 461146 210218 461382 210454
rect 460826 209898 461062 210134
rect 461146 209898 461382 210134
rect 460826 174218 461062 174454
rect 461146 174218 461382 174454
rect 460826 173898 461062 174134
rect 461146 173898 461382 174134
rect 460826 138218 461062 138454
rect 461146 138218 461382 138454
rect 460826 137898 461062 138134
rect 461146 137898 461382 138134
rect 460826 102218 461062 102454
rect 461146 102218 461382 102454
rect 460826 101898 461062 102134
rect 461146 101898 461382 102134
rect 460826 66218 461062 66454
rect 461146 66218 461382 66454
rect 460826 65898 461062 66134
rect 461146 65898 461382 66134
rect 460826 30218 461062 30454
rect 461146 30218 461382 30454
rect 460826 29898 461062 30134
rect 461146 29898 461382 30134
rect 460826 -6342 461062 -6106
rect 461146 -6342 461382 -6106
rect 460826 -6662 461062 -6426
rect 461146 -6662 461382 -6426
rect 465326 711322 465562 711558
rect 465646 711322 465882 711558
rect 465326 711002 465562 711238
rect 465646 711002 465882 711238
rect 465326 682718 465562 682954
rect 465646 682718 465882 682954
rect 465326 682398 465562 682634
rect 465646 682398 465882 682634
rect 465326 646718 465562 646954
rect 465646 646718 465882 646954
rect 465326 646398 465562 646634
rect 465646 646398 465882 646634
rect 465326 610718 465562 610954
rect 465646 610718 465882 610954
rect 465326 610398 465562 610634
rect 465646 610398 465882 610634
rect 465326 574718 465562 574954
rect 465646 574718 465882 574954
rect 465326 574398 465562 574634
rect 465646 574398 465882 574634
rect 465326 538718 465562 538954
rect 465646 538718 465882 538954
rect 465326 538398 465562 538634
rect 465646 538398 465882 538634
rect 465326 502718 465562 502954
rect 465646 502718 465882 502954
rect 465326 502398 465562 502634
rect 465646 502398 465882 502634
rect 465326 466718 465562 466954
rect 465646 466718 465882 466954
rect 465326 466398 465562 466634
rect 465646 466398 465882 466634
rect 465326 430718 465562 430954
rect 465646 430718 465882 430954
rect 465326 430398 465562 430634
rect 465646 430398 465882 430634
rect 465326 394718 465562 394954
rect 465646 394718 465882 394954
rect 465326 394398 465562 394634
rect 465646 394398 465882 394634
rect 465326 358718 465562 358954
rect 465646 358718 465882 358954
rect 465326 358398 465562 358634
rect 465646 358398 465882 358634
rect 465326 322718 465562 322954
rect 465646 322718 465882 322954
rect 465326 322398 465562 322634
rect 465646 322398 465882 322634
rect 465326 286718 465562 286954
rect 465646 286718 465882 286954
rect 465326 286398 465562 286634
rect 465646 286398 465882 286634
rect 465326 250718 465562 250954
rect 465646 250718 465882 250954
rect 465326 250398 465562 250634
rect 465646 250398 465882 250634
rect 465326 214718 465562 214954
rect 465646 214718 465882 214954
rect 465326 214398 465562 214634
rect 465646 214398 465882 214634
rect 465326 178718 465562 178954
rect 465646 178718 465882 178954
rect 465326 178398 465562 178634
rect 465646 178398 465882 178634
rect 465326 142718 465562 142954
rect 465646 142718 465882 142954
rect 465326 142398 465562 142634
rect 465646 142398 465882 142634
rect 465326 106718 465562 106954
rect 465646 106718 465882 106954
rect 465326 106398 465562 106634
rect 465646 106398 465882 106634
rect 465326 70718 465562 70954
rect 465646 70718 465882 70954
rect 465326 70398 465562 70634
rect 465646 70398 465882 70634
rect 465326 34718 465562 34954
rect 465646 34718 465882 34954
rect 465326 34398 465562 34634
rect 465646 34398 465882 34634
rect 465326 -7302 465562 -7066
rect 465646 -7302 465882 -7066
rect 465326 -7622 465562 -7386
rect 465646 -7622 465882 -7386
rect 469826 704602 470062 704838
rect 470146 704602 470382 704838
rect 469826 704282 470062 704518
rect 470146 704282 470382 704518
rect 469826 687218 470062 687454
rect 470146 687218 470382 687454
rect 469826 686898 470062 687134
rect 470146 686898 470382 687134
rect 469826 651218 470062 651454
rect 470146 651218 470382 651454
rect 469826 650898 470062 651134
rect 470146 650898 470382 651134
rect 469826 615218 470062 615454
rect 470146 615218 470382 615454
rect 469826 614898 470062 615134
rect 470146 614898 470382 615134
rect 469826 579218 470062 579454
rect 470146 579218 470382 579454
rect 469826 578898 470062 579134
rect 470146 578898 470382 579134
rect 469826 543218 470062 543454
rect 470146 543218 470382 543454
rect 469826 542898 470062 543134
rect 470146 542898 470382 543134
rect 469826 507218 470062 507454
rect 470146 507218 470382 507454
rect 469826 506898 470062 507134
rect 470146 506898 470382 507134
rect 469826 471218 470062 471454
rect 470146 471218 470382 471454
rect 469826 470898 470062 471134
rect 470146 470898 470382 471134
rect 469826 435218 470062 435454
rect 470146 435218 470382 435454
rect 469826 434898 470062 435134
rect 470146 434898 470382 435134
rect 469826 399218 470062 399454
rect 470146 399218 470382 399454
rect 469826 398898 470062 399134
rect 470146 398898 470382 399134
rect 469826 363218 470062 363454
rect 470146 363218 470382 363454
rect 469826 362898 470062 363134
rect 470146 362898 470382 363134
rect 469826 327218 470062 327454
rect 470146 327218 470382 327454
rect 469826 326898 470062 327134
rect 470146 326898 470382 327134
rect 469826 291218 470062 291454
rect 470146 291218 470382 291454
rect 469826 290898 470062 291134
rect 470146 290898 470382 291134
rect 469826 255218 470062 255454
rect 470146 255218 470382 255454
rect 469826 254898 470062 255134
rect 470146 254898 470382 255134
rect 469826 219218 470062 219454
rect 470146 219218 470382 219454
rect 469826 218898 470062 219134
rect 470146 218898 470382 219134
rect 469826 183218 470062 183454
rect 470146 183218 470382 183454
rect 469826 182898 470062 183134
rect 470146 182898 470382 183134
rect 469826 147218 470062 147454
rect 470146 147218 470382 147454
rect 469826 146898 470062 147134
rect 470146 146898 470382 147134
rect 469826 111218 470062 111454
rect 470146 111218 470382 111454
rect 469826 110898 470062 111134
rect 470146 110898 470382 111134
rect 469826 75218 470062 75454
rect 470146 75218 470382 75454
rect 469826 74898 470062 75134
rect 470146 74898 470382 75134
rect 469826 39218 470062 39454
rect 470146 39218 470382 39454
rect 469826 38898 470062 39134
rect 470146 38898 470382 39134
rect 469826 3218 470062 3454
rect 470146 3218 470382 3454
rect 469826 2898 470062 3134
rect 470146 2898 470382 3134
rect 469826 -582 470062 -346
rect 470146 -582 470382 -346
rect 469826 -902 470062 -666
rect 470146 -902 470382 -666
rect 474326 705562 474562 705798
rect 474646 705562 474882 705798
rect 474326 705242 474562 705478
rect 474646 705242 474882 705478
rect 474326 691718 474562 691954
rect 474646 691718 474882 691954
rect 474326 691398 474562 691634
rect 474646 691398 474882 691634
rect 474326 655718 474562 655954
rect 474646 655718 474882 655954
rect 474326 655398 474562 655634
rect 474646 655398 474882 655634
rect 474326 619718 474562 619954
rect 474646 619718 474882 619954
rect 474326 619398 474562 619634
rect 474646 619398 474882 619634
rect 474326 583718 474562 583954
rect 474646 583718 474882 583954
rect 474326 583398 474562 583634
rect 474646 583398 474882 583634
rect 474326 547718 474562 547954
rect 474646 547718 474882 547954
rect 474326 547398 474562 547634
rect 474646 547398 474882 547634
rect 474326 511718 474562 511954
rect 474646 511718 474882 511954
rect 474326 511398 474562 511634
rect 474646 511398 474882 511634
rect 474326 475718 474562 475954
rect 474646 475718 474882 475954
rect 474326 475398 474562 475634
rect 474646 475398 474882 475634
rect 474326 439718 474562 439954
rect 474646 439718 474882 439954
rect 474326 439398 474562 439634
rect 474646 439398 474882 439634
rect 474326 403718 474562 403954
rect 474646 403718 474882 403954
rect 474326 403398 474562 403634
rect 474646 403398 474882 403634
rect 474326 367718 474562 367954
rect 474646 367718 474882 367954
rect 474326 367398 474562 367634
rect 474646 367398 474882 367634
rect 474326 331718 474562 331954
rect 474646 331718 474882 331954
rect 474326 331398 474562 331634
rect 474646 331398 474882 331634
rect 474326 295718 474562 295954
rect 474646 295718 474882 295954
rect 474326 295398 474562 295634
rect 474646 295398 474882 295634
rect 474326 259718 474562 259954
rect 474646 259718 474882 259954
rect 474326 259398 474562 259634
rect 474646 259398 474882 259634
rect 474326 223718 474562 223954
rect 474646 223718 474882 223954
rect 474326 223398 474562 223634
rect 474646 223398 474882 223634
rect 474326 187718 474562 187954
rect 474646 187718 474882 187954
rect 474326 187398 474562 187634
rect 474646 187398 474882 187634
rect 474326 151718 474562 151954
rect 474646 151718 474882 151954
rect 474326 151398 474562 151634
rect 474646 151398 474882 151634
rect 474326 115718 474562 115954
rect 474646 115718 474882 115954
rect 474326 115398 474562 115634
rect 474646 115398 474882 115634
rect 474326 79718 474562 79954
rect 474646 79718 474882 79954
rect 474326 79398 474562 79634
rect 474646 79398 474882 79634
rect 474326 43718 474562 43954
rect 474646 43718 474882 43954
rect 474326 43398 474562 43634
rect 474646 43398 474882 43634
rect 474326 7718 474562 7954
rect 474646 7718 474882 7954
rect 474326 7398 474562 7634
rect 474646 7398 474882 7634
rect 474326 -1542 474562 -1306
rect 474646 -1542 474882 -1306
rect 474326 -1862 474562 -1626
rect 474646 -1862 474882 -1626
rect 478826 706522 479062 706758
rect 479146 706522 479382 706758
rect 478826 706202 479062 706438
rect 479146 706202 479382 706438
rect 478826 696218 479062 696454
rect 479146 696218 479382 696454
rect 478826 695898 479062 696134
rect 479146 695898 479382 696134
rect 478826 660218 479062 660454
rect 479146 660218 479382 660454
rect 478826 659898 479062 660134
rect 479146 659898 479382 660134
rect 478826 624218 479062 624454
rect 479146 624218 479382 624454
rect 478826 623898 479062 624134
rect 479146 623898 479382 624134
rect 478826 588218 479062 588454
rect 479146 588218 479382 588454
rect 478826 587898 479062 588134
rect 479146 587898 479382 588134
rect 478826 552218 479062 552454
rect 479146 552218 479382 552454
rect 478826 551898 479062 552134
rect 479146 551898 479382 552134
rect 478826 516218 479062 516454
rect 479146 516218 479382 516454
rect 478826 515898 479062 516134
rect 479146 515898 479382 516134
rect 478826 480218 479062 480454
rect 479146 480218 479382 480454
rect 478826 479898 479062 480134
rect 479146 479898 479382 480134
rect 478826 444218 479062 444454
rect 479146 444218 479382 444454
rect 478826 443898 479062 444134
rect 479146 443898 479382 444134
rect 478826 408218 479062 408454
rect 479146 408218 479382 408454
rect 478826 407898 479062 408134
rect 479146 407898 479382 408134
rect 478826 372218 479062 372454
rect 479146 372218 479382 372454
rect 478826 371898 479062 372134
rect 479146 371898 479382 372134
rect 478826 336218 479062 336454
rect 479146 336218 479382 336454
rect 478826 335898 479062 336134
rect 479146 335898 479382 336134
rect 478826 300218 479062 300454
rect 479146 300218 479382 300454
rect 478826 299898 479062 300134
rect 479146 299898 479382 300134
rect 478826 264218 479062 264454
rect 479146 264218 479382 264454
rect 478826 263898 479062 264134
rect 479146 263898 479382 264134
rect 478826 228218 479062 228454
rect 479146 228218 479382 228454
rect 478826 227898 479062 228134
rect 479146 227898 479382 228134
rect 478826 192218 479062 192454
rect 479146 192218 479382 192454
rect 478826 191898 479062 192134
rect 479146 191898 479382 192134
rect 478826 156218 479062 156454
rect 479146 156218 479382 156454
rect 478826 155898 479062 156134
rect 479146 155898 479382 156134
rect 478826 120218 479062 120454
rect 479146 120218 479382 120454
rect 478826 119898 479062 120134
rect 479146 119898 479382 120134
rect 478826 84218 479062 84454
rect 479146 84218 479382 84454
rect 478826 83898 479062 84134
rect 479146 83898 479382 84134
rect 478826 48218 479062 48454
rect 479146 48218 479382 48454
rect 478826 47898 479062 48134
rect 479146 47898 479382 48134
rect 478826 12218 479062 12454
rect 479146 12218 479382 12454
rect 478826 11898 479062 12134
rect 479146 11898 479382 12134
rect 478826 -2502 479062 -2266
rect 479146 -2502 479382 -2266
rect 478826 -2822 479062 -2586
rect 479146 -2822 479382 -2586
rect 483326 707482 483562 707718
rect 483646 707482 483882 707718
rect 483326 707162 483562 707398
rect 483646 707162 483882 707398
rect 483326 700718 483562 700954
rect 483646 700718 483882 700954
rect 483326 700398 483562 700634
rect 483646 700398 483882 700634
rect 483326 664718 483562 664954
rect 483646 664718 483882 664954
rect 483326 664398 483562 664634
rect 483646 664398 483882 664634
rect 483326 628718 483562 628954
rect 483646 628718 483882 628954
rect 483326 628398 483562 628634
rect 483646 628398 483882 628634
rect 483326 592718 483562 592954
rect 483646 592718 483882 592954
rect 483326 592398 483562 592634
rect 483646 592398 483882 592634
rect 483326 556718 483562 556954
rect 483646 556718 483882 556954
rect 483326 556398 483562 556634
rect 483646 556398 483882 556634
rect 483326 520718 483562 520954
rect 483646 520718 483882 520954
rect 483326 520398 483562 520634
rect 483646 520398 483882 520634
rect 483326 484718 483562 484954
rect 483646 484718 483882 484954
rect 483326 484398 483562 484634
rect 483646 484398 483882 484634
rect 483326 448718 483562 448954
rect 483646 448718 483882 448954
rect 483326 448398 483562 448634
rect 483646 448398 483882 448634
rect 483326 412718 483562 412954
rect 483646 412718 483882 412954
rect 483326 412398 483562 412634
rect 483646 412398 483882 412634
rect 483326 376718 483562 376954
rect 483646 376718 483882 376954
rect 483326 376398 483562 376634
rect 483646 376398 483882 376634
rect 483326 340718 483562 340954
rect 483646 340718 483882 340954
rect 483326 340398 483562 340634
rect 483646 340398 483882 340634
rect 483326 304718 483562 304954
rect 483646 304718 483882 304954
rect 483326 304398 483562 304634
rect 483646 304398 483882 304634
rect 483326 268718 483562 268954
rect 483646 268718 483882 268954
rect 483326 268398 483562 268634
rect 483646 268398 483882 268634
rect 483326 232718 483562 232954
rect 483646 232718 483882 232954
rect 483326 232398 483562 232634
rect 483646 232398 483882 232634
rect 483326 196718 483562 196954
rect 483646 196718 483882 196954
rect 483326 196398 483562 196634
rect 483646 196398 483882 196634
rect 483326 160718 483562 160954
rect 483646 160718 483882 160954
rect 483326 160398 483562 160634
rect 483646 160398 483882 160634
rect 483326 124718 483562 124954
rect 483646 124718 483882 124954
rect 483326 124398 483562 124634
rect 483646 124398 483882 124634
rect 483326 88718 483562 88954
rect 483646 88718 483882 88954
rect 483326 88398 483562 88634
rect 483646 88398 483882 88634
rect 483326 52718 483562 52954
rect 483646 52718 483882 52954
rect 483326 52398 483562 52634
rect 483646 52398 483882 52634
rect 483326 16718 483562 16954
rect 483646 16718 483882 16954
rect 483326 16398 483562 16634
rect 483646 16398 483882 16634
rect 483326 -3462 483562 -3226
rect 483646 -3462 483882 -3226
rect 483326 -3782 483562 -3546
rect 483646 -3782 483882 -3546
rect 487826 708442 488062 708678
rect 488146 708442 488382 708678
rect 487826 708122 488062 708358
rect 488146 708122 488382 708358
rect 487826 669218 488062 669454
rect 488146 669218 488382 669454
rect 487826 668898 488062 669134
rect 488146 668898 488382 669134
rect 487826 633218 488062 633454
rect 488146 633218 488382 633454
rect 487826 632898 488062 633134
rect 488146 632898 488382 633134
rect 487826 597218 488062 597454
rect 488146 597218 488382 597454
rect 487826 596898 488062 597134
rect 488146 596898 488382 597134
rect 487826 561218 488062 561454
rect 488146 561218 488382 561454
rect 487826 560898 488062 561134
rect 488146 560898 488382 561134
rect 487826 525218 488062 525454
rect 488146 525218 488382 525454
rect 487826 524898 488062 525134
rect 488146 524898 488382 525134
rect 487826 489218 488062 489454
rect 488146 489218 488382 489454
rect 487826 488898 488062 489134
rect 488146 488898 488382 489134
rect 487826 453218 488062 453454
rect 488146 453218 488382 453454
rect 487826 452898 488062 453134
rect 488146 452898 488382 453134
rect 487826 417218 488062 417454
rect 488146 417218 488382 417454
rect 487826 416898 488062 417134
rect 488146 416898 488382 417134
rect 487826 381218 488062 381454
rect 488146 381218 488382 381454
rect 487826 380898 488062 381134
rect 488146 380898 488382 381134
rect 487826 345218 488062 345454
rect 488146 345218 488382 345454
rect 487826 344898 488062 345134
rect 488146 344898 488382 345134
rect 487826 309218 488062 309454
rect 488146 309218 488382 309454
rect 487826 308898 488062 309134
rect 488146 308898 488382 309134
rect 487826 273218 488062 273454
rect 488146 273218 488382 273454
rect 487826 272898 488062 273134
rect 488146 272898 488382 273134
rect 487826 237218 488062 237454
rect 488146 237218 488382 237454
rect 487826 236898 488062 237134
rect 488146 236898 488382 237134
rect 487826 201218 488062 201454
rect 488146 201218 488382 201454
rect 487826 200898 488062 201134
rect 488146 200898 488382 201134
rect 487826 165218 488062 165454
rect 488146 165218 488382 165454
rect 487826 164898 488062 165134
rect 488146 164898 488382 165134
rect 487826 129218 488062 129454
rect 488146 129218 488382 129454
rect 487826 128898 488062 129134
rect 488146 128898 488382 129134
rect 487826 93218 488062 93454
rect 488146 93218 488382 93454
rect 487826 92898 488062 93134
rect 488146 92898 488382 93134
rect 487826 57218 488062 57454
rect 488146 57218 488382 57454
rect 487826 56898 488062 57134
rect 488146 56898 488382 57134
rect 487826 21218 488062 21454
rect 488146 21218 488382 21454
rect 487826 20898 488062 21134
rect 488146 20898 488382 21134
rect 487826 -4422 488062 -4186
rect 488146 -4422 488382 -4186
rect 487826 -4742 488062 -4506
rect 488146 -4742 488382 -4506
rect 492326 709402 492562 709638
rect 492646 709402 492882 709638
rect 492326 709082 492562 709318
rect 492646 709082 492882 709318
rect 492326 673718 492562 673954
rect 492646 673718 492882 673954
rect 492326 673398 492562 673634
rect 492646 673398 492882 673634
rect 492326 637718 492562 637954
rect 492646 637718 492882 637954
rect 492326 637398 492562 637634
rect 492646 637398 492882 637634
rect 492326 601718 492562 601954
rect 492646 601718 492882 601954
rect 492326 601398 492562 601634
rect 492646 601398 492882 601634
rect 492326 565718 492562 565954
rect 492646 565718 492882 565954
rect 492326 565398 492562 565634
rect 492646 565398 492882 565634
rect 492326 529718 492562 529954
rect 492646 529718 492882 529954
rect 492326 529398 492562 529634
rect 492646 529398 492882 529634
rect 492326 493718 492562 493954
rect 492646 493718 492882 493954
rect 492326 493398 492562 493634
rect 492646 493398 492882 493634
rect 492326 457718 492562 457954
rect 492646 457718 492882 457954
rect 492326 457398 492562 457634
rect 492646 457398 492882 457634
rect 492326 421718 492562 421954
rect 492646 421718 492882 421954
rect 492326 421398 492562 421634
rect 492646 421398 492882 421634
rect 492326 385718 492562 385954
rect 492646 385718 492882 385954
rect 492326 385398 492562 385634
rect 492646 385398 492882 385634
rect 492326 349718 492562 349954
rect 492646 349718 492882 349954
rect 492326 349398 492562 349634
rect 492646 349398 492882 349634
rect 492326 313718 492562 313954
rect 492646 313718 492882 313954
rect 492326 313398 492562 313634
rect 492646 313398 492882 313634
rect 492326 277718 492562 277954
rect 492646 277718 492882 277954
rect 492326 277398 492562 277634
rect 492646 277398 492882 277634
rect 492326 241718 492562 241954
rect 492646 241718 492882 241954
rect 492326 241398 492562 241634
rect 492646 241398 492882 241634
rect 492326 205718 492562 205954
rect 492646 205718 492882 205954
rect 492326 205398 492562 205634
rect 492646 205398 492882 205634
rect 492326 169718 492562 169954
rect 492646 169718 492882 169954
rect 492326 169398 492562 169634
rect 492646 169398 492882 169634
rect 492326 133718 492562 133954
rect 492646 133718 492882 133954
rect 492326 133398 492562 133634
rect 492646 133398 492882 133634
rect 492326 97718 492562 97954
rect 492646 97718 492882 97954
rect 492326 97398 492562 97634
rect 492646 97398 492882 97634
rect 492326 61718 492562 61954
rect 492646 61718 492882 61954
rect 492326 61398 492562 61634
rect 492646 61398 492882 61634
rect 492326 25718 492562 25954
rect 492646 25718 492882 25954
rect 492326 25398 492562 25634
rect 492646 25398 492882 25634
rect 492326 -5382 492562 -5146
rect 492646 -5382 492882 -5146
rect 492326 -5702 492562 -5466
rect 492646 -5702 492882 -5466
rect 496826 710362 497062 710598
rect 497146 710362 497382 710598
rect 496826 710042 497062 710278
rect 497146 710042 497382 710278
rect 496826 678218 497062 678454
rect 497146 678218 497382 678454
rect 496826 677898 497062 678134
rect 497146 677898 497382 678134
rect 496826 642218 497062 642454
rect 497146 642218 497382 642454
rect 496826 641898 497062 642134
rect 497146 641898 497382 642134
rect 496826 606218 497062 606454
rect 497146 606218 497382 606454
rect 496826 605898 497062 606134
rect 497146 605898 497382 606134
rect 496826 570218 497062 570454
rect 497146 570218 497382 570454
rect 496826 569898 497062 570134
rect 497146 569898 497382 570134
rect 496826 534218 497062 534454
rect 497146 534218 497382 534454
rect 496826 533898 497062 534134
rect 497146 533898 497382 534134
rect 496826 498218 497062 498454
rect 497146 498218 497382 498454
rect 496826 497898 497062 498134
rect 497146 497898 497382 498134
rect 496826 462218 497062 462454
rect 497146 462218 497382 462454
rect 496826 461898 497062 462134
rect 497146 461898 497382 462134
rect 496826 426218 497062 426454
rect 497146 426218 497382 426454
rect 496826 425898 497062 426134
rect 497146 425898 497382 426134
rect 496826 390218 497062 390454
rect 497146 390218 497382 390454
rect 496826 389898 497062 390134
rect 497146 389898 497382 390134
rect 496826 354218 497062 354454
rect 497146 354218 497382 354454
rect 496826 353898 497062 354134
rect 497146 353898 497382 354134
rect 496826 318218 497062 318454
rect 497146 318218 497382 318454
rect 496826 317898 497062 318134
rect 497146 317898 497382 318134
rect 496826 282218 497062 282454
rect 497146 282218 497382 282454
rect 496826 281898 497062 282134
rect 497146 281898 497382 282134
rect 496826 246218 497062 246454
rect 497146 246218 497382 246454
rect 496826 245898 497062 246134
rect 497146 245898 497382 246134
rect 496826 210218 497062 210454
rect 497146 210218 497382 210454
rect 496826 209898 497062 210134
rect 497146 209898 497382 210134
rect 496826 174218 497062 174454
rect 497146 174218 497382 174454
rect 496826 173898 497062 174134
rect 497146 173898 497382 174134
rect 496826 138218 497062 138454
rect 497146 138218 497382 138454
rect 496826 137898 497062 138134
rect 497146 137898 497382 138134
rect 496826 102218 497062 102454
rect 497146 102218 497382 102454
rect 496826 101898 497062 102134
rect 497146 101898 497382 102134
rect 496826 66218 497062 66454
rect 497146 66218 497382 66454
rect 496826 65898 497062 66134
rect 497146 65898 497382 66134
rect 496826 30218 497062 30454
rect 497146 30218 497382 30454
rect 496826 29898 497062 30134
rect 497146 29898 497382 30134
rect 496826 -6342 497062 -6106
rect 497146 -6342 497382 -6106
rect 496826 -6662 497062 -6426
rect 497146 -6662 497382 -6426
rect 501326 711322 501562 711558
rect 501646 711322 501882 711558
rect 501326 711002 501562 711238
rect 501646 711002 501882 711238
rect 501326 682718 501562 682954
rect 501646 682718 501882 682954
rect 501326 682398 501562 682634
rect 501646 682398 501882 682634
rect 501326 646718 501562 646954
rect 501646 646718 501882 646954
rect 501326 646398 501562 646634
rect 501646 646398 501882 646634
rect 501326 610718 501562 610954
rect 501646 610718 501882 610954
rect 501326 610398 501562 610634
rect 501646 610398 501882 610634
rect 501326 574718 501562 574954
rect 501646 574718 501882 574954
rect 501326 574398 501562 574634
rect 501646 574398 501882 574634
rect 501326 538718 501562 538954
rect 501646 538718 501882 538954
rect 501326 538398 501562 538634
rect 501646 538398 501882 538634
rect 501326 502718 501562 502954
rect 501646 502718 501882 502954
rect 501326 502398 501562 502634
rect 501646 502398 501882 502634
rect 501326 466718 501562 466954
rect 501646 466718 501882 466954
rect 501326 466398 501562 466634
rect 501646 466398 501882 466634
rect 501326 430718 501562 430954
rect 501646 430718 501882 430954
rect 501326 430398 501562 430634
rect 501646 430398 501882 430634
rect 501326 394718 501562 394954
rect 501646 394718 501882 394954
rect 501326 394398 501562 394634
rect 501646 394398 501882 394634
rect 501326 358718 501562 358954
rect 501646 358718 501882 358954
rect 501326 358398 501562 358634
rect 501646 358398 501882 358634
rect 501326 322718 501562 322954
rect 501646 322718 501882 322954
rect 501326 322398 501562 322634
rect 501646 322398 501882 322634
rect 501326 286718 501562 286954
rect 501646 286718 501882 286954
rect 501326 286398 501562 286634
rect 501646 286398 501882 286634
rect 501326 250718 501562 250954
rect 501646 250718 501882 250954
rect 501326 250398 501562 250634
rect 501646 250398 501882 250634
rect 501326 214718 501562 214954
rect 501646 214718 501882 214954
rect 501326 214398 501562 214634
rect 501646 214398 501882 214634
rect 501326 178718 501562 178954
rect 501646 178718 501882 178954
rect 501326 178398 501562 178634
rect 501646 178398 501882 178634
rect 501326 142718 501562 142954
rect 501646 142718 501882 142954
rect 501326 142398 501562 142634
rect 501646 142398 501882 142634
rect 501326 106718 501562 106954
rect 501646 106718 501882 106954
rect 501326 106398 501562 106634
rect 501646 106398 501882 106634
rect 501326 70718 501562 70954
rect 501646 70718 501882 70954
rect 501326 70398 501562 70634
rect 501646 70398 501882 70634
rect 501326 34718 501562 34954
rect 501646 34718 501882 34954
rect 501326 34398 501562 34634
rect 501646 34398 501882 34634
rect 501326 -7302 501562 -7066
rect 501646 -7302 501882 -7066
rect 501326 -7622 501562 -7386
rect 501646 -7622 501882 -7386
rect 505826 704602 506062 704838
rect 506146 704602 506382 704838
rect 505826 704282 506062 704518
rect 506146 704282 506382 704518
rect 505826 687218 506062 687454
rect 506146 687218 506382 687454
rect 505826 686898 506062 687134
rect 506146 686898 506382 687134
rect 505826 651218 506062 651454
rect 506146 651218 506382 651454
rect 505826 650898 506062 651134
rect 506146 650898 506382 651134
rect 505826 615218 506062 615454
rect 506146 615218 506382 615454
rect 505826 614898 506062 615134
rect 506146 614898 506382 615134
rect 505826 579218 506062 579454
rect 506146 579218 506382 579454
rect 505826 578898 506062 579134
rect 506146 578898 506382 579134
rect 505826 543218 506062 543454
rect 506146 543218 506382 543454
rect 505826 542898 506062 543134
rect 506146 542898 506382 543134
rect 505826 507218 506062 507454
rect 506146 507218 506382 507454
rect 505826 506898 506062 507134
rect 506146 506898 506382 507134
rect 505826 471218 506062 471454
rect 506146 471218 506382 471454
rect 505826 470898 506062 471134
rect 506146 470898 506382 471134
rect 505826 435218 506062 435454
rect 506146 435218 506382 435454
rect 505826 434898 506062 435134
rect 506146 434898 506382 435134
rect 505826 399218 506062 399454
rect 506146 399218 506382 399454
rect 505826 398898 506062 399134
rect 506146 398898 506382 399134
rect 505826 363218 506062 363454
rect 506146 363218 506382 363454
rect 505826 362898 506062 363134
rect 506146 362898 506382 363134
rect 505826 327218 506062 327454
rect 506146 327218 506382 327454
rect 505826 326898 506062 327134
rect 506146 326898 506382 327134
rect 505826 291218 506062 291454
rect 506146 291218 506382 291454
rect 505826 290898 506062 291134
rect 506146 290898 506382 291134
rect 505826 255218 506062 255454
rect 506146 255218 506382 255454
rect 505826 254898 506062 255134
rect 506146 254898 506382 255134
rect 505826 219218 506062 219454
rect 506146 219218 506382 219454
rect 505826 218898 506062 219134
rect 506146 218898 506382 219134
rect 505826 183218 506062 183454
rect 506146 183218 506382 183454
rect 505826 182898 506062 183134
rect 506146 182898 506382 183134
rect 505826 147218 506062 147454
rect 506146 147218 506382 147454
rect 505826 146898 506062 147134
rect 506146 146898 506382 147134
rect 505826 111218 506062 111454
rect 506146 111218 506382 111454
rect 505826 110898 506062 111134
rect 506146 110898 506382 111134
rect 505826 75218 506062 75454
rect 506146 75218 506382 75454
rect 505826 74898 506062 75134
rect 506146 74898 506382 75134
rect 505826 39218 506062 39454
rect 506146 39218 506382 39454
rect 505826 38898 506062 39134
rect 506146 38898 506382 39134
rect 505826 3218 506062 3454
rect 506146 3218 506382 3454
rect 505826 2898 506062 3134
rect 506146 2898 506382 3134
rect 505826 -582 506062 -346
rect 506146 -582 506382 -346
rect 505826 -902 506062 -666
rect 506146 -902 506382 -666
rect 510326 705562 510562 705798
rect 510646 705562 510882 705798
rect 510326 705242 510562 705478
rect 510646 705242 510882 705478
rect 510326 691718 510562 691954
rect 510646 691718 510882 691954
rect 510326 691398 510562 691634
rect 510646 691398 510882 691634
rect 510326 655718 510562 655954
rect 510646 655718 510882 655954
rect 510326 655398 510562 655634
rect 510646 655398 510882 655634
rect 510326 619718 510562 619954
rect 510646 619718 510882 619954
rect 510326 619398 510562 619634
rect 510646 619398 510882 619634
rect 510326 583718 510562 583954
rect 510646 583718 510882 583954
rect 510326 583398 510562 583634
rect 510646 583398 510882 583634
rect 510326 547718 510562 547954
rect 510646 547718 510882 547954
rect 510326 547398 510562 547634
rect 510646 547398 510882 547634
rect 510326 511718 510562 511954
rect 510646 511718 510882 511954
rect 510326 511398 510562 511634
rect 510646 511398 510882 511634
rect 510326 475718 510562 475954
rect 510646 475718 510882 475954
rect 510326 475398 510562 475634
rect 510646 475398 510882 475634
rect 510326 439718 510562 439954
rect 510646 439718 510882 439954
rect 510326 439398 510562 439634
rect 510646 439398 510882 439634
rect 510326 403718 510562 403954
rect 510646 403718 510882 403954
rect 510326 403398 510562 403634
rect 510646 403398 510882 403634
rect 510326 367718 510562 367954
rect 510646 367718 510882 367954
rect 510326 367398 510562 367634
rect 510646 367398 510882 367634
rect 510326 331718 510562 331954
rect 510646 331718 510882 331954
rect 510326 331398 510562 331634
rect 510646 331398 510882 331634
rect 510326 295718 510562 295954
rect 510646 295718 510882 295954
rect 510326 295398 510562 295634
rect 510646 295398 510882 295634
rect 510326 259718 510562 259954
rect 510646 259718 510882 259954
rect 510326 259398 510562 259634
rect 510646 259398 510882 259634
rect 510326 223718 510562 223954
rect 510646 223718 510882 223954
rect 510326 223398 510562 223634
rect 510646 223398 510882 223634
rect 510326 187718 510562 187954
rect 510646 187718 510882 187954
rect 510326 187398 510562 187634
rect 510646 187398 510882 187634
rect 510326 151718 510562 151954
rect 510646 151718 510882 151954
rect 510326 151398 510562 151634
rect 510646 151398 510882 151634
rect 510326 115718 510562 115954
rect 510646 115718 510882 115954
rect 510326 115398 510562 115634
rect 510646 115398 510882 115634
rect 510326 79718 510562 79954
rect 510646 79718 510882 79954
rect 510326 79398 510562 79634
rect 510646 79398 510882 79634
rect 510326 43718 510562 43954
rect 510646 43718 510882 43954
rect 510326 43398 510562 43634
rect 510646 43398 510882 43634
rect 510326 7718 510562 7954
rect 510646 7718 510882 7954
rect 510326 7398 510562 7634
rect 510646 7398 510882 7634
rect 510326 -1542 510562 -1306
rect 510646 -1542 510882 -1306
rect 510326 -1862 510562 -1626
rect 510646 -1862 510882 -1626
rect 514826 706522 515062 706758
rect 515146 706522 515382 706758
rect 514826 706202 515062 706438
rect 515146 706202 515382 706438
rect 514826 696218 515062 696454
rect 515146 696218 515382 696454
rect 514826 695898 515062 696134
rect 515146 695898 515382 696134
rect 514826 660218 515062 660454
rect 515146 660218 515382 660454
rect 514826 659898 515062 660134
rect 515146 659898 515382 660134
rect 514826 624218 515062 624454
rect 515146 624218 515382 624454
rect 514826 623898 515062 624134
rect 515146 623898 515382 624134
rect 514826 588218 515062 588454
rect 515146 588218 515382 588454
rect 514826 587898 515062 588134
rect 515146 587898 515382 588134
rect 514826 552218 515062 552454
rect 515146 552218 515382 552454
rect 514826 551898 515062 552134
rect 515146 551898 515382 552134
rect 514826 516218 515062 516454
rect 515146 516218 515382 516454
rect 514826 515898 515062 516134
rect 515146 515898 515382 516134
rect 514826 480218 515062 480454
rect 515146 480218 515382 480454
rect 514826 479898 515062 480134
rect 515146 479898 515382 480134
rect 514826 444218 515062 444454
rect 515146 444218 515382 444454
rect 514826 443898 515062 444134
rect 515146 443898 515382 444134
rect 514826 408218 515062 408454
rect 515146 408218 515382 408454
rect 514826 407898 515062 408134
rect 515146 407898 515382 408134
rect 514826 372218 515062 372454
rect 515146 372218 515382 372454
rect 514826 371898 515062 372134
rect 515146 371898 515382 372134
rect 514826 336218 515062 336454
rect 515146 336218 515382 336454
rect 514826 335898 515062 336134
rect 515146 335898 515382 336134
rect 514826 300218 515062 300454
rect 515146 300218 515382 300454
rect 514826 299898 515062 300134
rect 515146 299898 515382 300134
rect 514826 264218 515062 264454
rect 515146 264218 515382 264454
rect 514826 263898 515062 264134
rect 515146 263898 515382 264134
rect 514826 228218 515062 228454
rect 515146 228218 515382 228454
rect 514826 227898 515062 228134
rect 515146 227898 515382 228134
rect 514826 192218 515062 192454
rect 515146 192218 515382 192454
rect 514826 191898 515062 192134
rect 515146 191898 515382 192134
rect 514826 156218 515062 156454
rect 515146 156218 515382 156454
rect 514826 155898 515062 156134
rect 515146 155898 515382 156134
rect 514826 120218 515062 120454
rect 515146 120218 515382 120454
rect 514826 119898 515062 120134
rect 515146 119898 515382 120134
rect 514826 84218 515062 84454
rect 515146 84218 515382 84454
rect 514826 83898 515062 84134
rect 515146 83898 515382 84134
rect 514826 48218 515062 48454
rect 515146 48218 515382 48454
rect 514826 47898 515062 48134
rect 515146 47898 515382 48134
rect 514826 12218 515062 12454
rect 515146 12218 515382 12454
rect 514826 11898 515062 12134
rect 515146 11898 515382 12134
rect 514826 -2502 515062 -2266
rect 515146 -2502 515382 -2266
rect 514826 -2822 515062 -2586
rect 515146 -2822 515382 -2586
rect 519326 707482 519562 707718
rect 519646 707482 519882 707718
rect 519326 707162 519562 707398
rect 519646 707162 519882 707398
rect 519326 700718 519562 700954
rect 519646 700718 519882 700954
rect 519326 700398 519562 700634
rect 519646 700398 519882 700634
rect 519326 664718 519562 664954
rect 519646 664718 519882 664954
rect 519326 664398 519562 664634
rect 519646 664398 519882 664634
rect 519326 628718 519562 628954
rect 519646 628718 519882 628954
rect 519326 628398 519562 628634
rect 519646 628398 519882 628634
rect 519326 592718 519562 592954
rect 519646 592718 519882 592954
rect 519326 592398 519562 592634
rect 519646 592398 519882 592634
rect 519326 556718 519562 556954
rect 519646 556718 519882 556954
rect 519326 556398 519562 556634
rect 519646 556398 519882 556634
rect 519326 520718 519562 520954
rect 519646 520718 519882 520954
rect 519326 520398 519562 520634
rect 519646 520398 519882 520634
rect 519326 484718 519562 484954
rect 519646 484718 519882 484954
rect 519326 484398 519562 484634
rect 519646 484398 519882 484634
rect 519326 448718 519562 448954
rect 519646 448718 519882 448954
rect 519326 448398 519562 448634
rect 519646 448398 519882 448634
rect 519326 412718 519562 412954
rect 519646 412718 519882 412954
rect 519326 412398 519562 412634
rect 519646 412398 519882 412634
rect 519326 376718 519562 376954
rect 519646 376718 519882 376954
rect 519326 376398 519562 376634
rect 519646 376398 519882 376634
rect 519326 340718 519562 340954
rect 519646 340718 519882 340954
rect 519326 340398 519562 340634
rect 519646 340398 519882 340634
rect 519326 304718 519562 304954
rect 519646 304718 519882 304954
rect 519326 304398 519562 304634
rect 519646 304398 519882 304634
rect 519326 268718 519562 268954
rect 519646 268718 519882 268954
rect 519326 268398 519562 268634
rect 519646 268398 519882 268634
rect 519326 232718 519562 232954
rect 519646 232718 519882 232954
rect 519326 232398 519562 232634
rect 519646 232398 519882 232634
rect 519326 196718 519562 196954
rect 519646 196718 519882 196954
rect 519326 196398 519562 196634
rect 519646 196398 519882 196634
rect 519326 160718 519562 160954
rect 519646 160718 519882 160954
rect 519326 160398 519562 160634
rect 519646 160398 519882 160634
rect 519326 124718 519562 124954
rect 519646 124718 519882 124954
rect 519326 124398 519562 124634
rect 519646 124398 519882 124634
rect 519326 88718 519562 88954
rect 519646 88718 519882 88954
rect 519326 88398 519562 88634
rect 519646 88398 519882 88634
rect 519326 52718 519562 52954
rect 519646 52718 519882 52954
rect 519326 52398 519562 52634
rect 519646 52398 519882 52634
rect 519326 16718 519562 16954
rect 519646 16718 519882 16954
rect 519326 16398 519562 16634
rect 519646 16398 519882 16634
rect 519326 -3462 519562 -3226
rect 519646 -3462 519882 -3226
rect 519326 -3782 519562 -3546
rect 519646 -3782 519882 -3546
rect 523826 708442 524062 708678
rect 524146 708442 524382 708678
rect 523826 708122 524062 708358
rect 524146 708122 524382 708358
rect 523826 669218 524062 669454
rect 524146 669218 524382 669454
rect 523826 668898 524062 669134
rect 524146 668898 524382 669134
rect 523826 633218 524062 633454
rect 524146 633218 524382 633454
rect 523826 632898 524062 633134
rect 524146 632898 524382 633134
rect 523826 597218 524062 597454
rect 524146 597218 524382 597454
rect 523826 596898 524062 597134
rect 524146 596898 524382 597134
rect 523826 561218 524062 561454
rect 524146 561218 524382 561454
rect 523826 560898 524062 561134
rect 524146 560898 524382 561134
rect 523826 525218 524062 525454
rect 524146 525218 524382 525454
rect 523826 524898 524062 525134
rect 524146 524898 524382 525134
rect 523826 489218 524062 489454
rect 524146 489218 524382 489454
rect 523826 488898 524062 489134
rect 524146 488898 524382 489134
rect 523826 453218 524062 453454
rect 524146 453218 524382 453454
rect 523826 452898 524062 453134
rect 524146 452898 524382 453134
rect 523826 417218 524062 417454
rect 524146 417218 524382 417454
rect 523826 416898 524062 417134
rect 524146 416898 524382 417134
rect 523826 381218 524062 381454
rect 524146 381218 524382 381454
rect 523826 380898 524062 381134
rect 524146 380898 524382 381134
rect 523826 345218 524062 345454
rect 524146 345218 524382 345454
rect 523826 344898 524062 345134
rect 524146 344898 524382 345134
rect 523826 309218 524062 309454
rect 524146 309218 524382 309454
rect 523826 308898 524062 309134
rect 524146 308898 524382 309134
rect 523826 273218 524062 273454
rect 524146 273218 524382 273454
rect 523826 272898 524062 273134
rect 524146 272898 524382 273134
rect 523826 237218 524062 237454
rect 524146 237218 524382 237454
rect 523826 236898 524062 237134
rect 524146 236898 524382 237134
rect 523826 201218 524062 201454
rect 524146 201218 524382 201454
rect 523826 200898 524062 201134
rect 524146 200898 524382 201134
rect 523826 165218 524062 165454
rect 524146 165218 524382 165454
rect 523826 164898 524062 165134
rect 524146 164898 524382 165134
rect 523826 129218 524062 129454
rect 524146 129218 524382 129454
rect 523826 128898 524062 129134
rect 524146 128898 524382 129134
rect 523826 93218 524062 93454
rect 524146 93218 524382 93454
rect 523826 92898 524062 93134
rect 524146 92898 524382 93134
rect 523826 57218 524062 57454
rect 524146 57218 524382 57454
rect 523826 56898 524062 57134
rect 524146 56898 524382 57134
rect 523826 21218 524062 21454
rect 524146 21218 524382 21454
rect 523826 20898 524062 21134
rect 524146 20898 524382 21134
rect 523826 -4422 524062 -4186
rect 524146 -4422 524382 -4186
rect 523826 -4742 524062 -4506
rect 524146 -4742 524382 -4506
rect 528326 709402 528562 709638
rect 528646 709402 528882 709638
rect 528326 709082 528562 709318
rect 528646 709082 528882 709318
rect 528326 673718 528562 673954
rect 528646 673718 528882 673954
rect 528326 673398 528562 673634
rect 528646 673398 528882 673634
rect 528326 637718 528562 637954
rect 528646 637718 528882 637954
rect 528326 637398 528562 637634
rect 528646 637398 528882 637634
rect 528326 601718 528562 601954
rect 528646 601718 528882 601954
rect 528326 601398 528562 601634
rect 528646 601398 528882 601634
rect 528326 565718 528562 565954
rect 528646 565718 528882 565954
rect 528326 565398 528562 565634
rect 528646 565398 528882 565634
rect 528326 529718 528562 529954
rect 528646 529718 528882 529954
rect 528326 529398 528562 529634
rect 528646 529398 528882 529634
rect 528326 493718 528562 493954
rect 528646 493718 528882 493954
rect 528326 493398 528562 493634
rect 528646 493398 528882 493634
rect 528326 457718 528562 457954
rect 528646 457718 528882 457954
rect 528326 457398 528562 457634
rect 528646 457398 528882 457634
rect 528326 421718 528562 421954
rect 528646 421718 528882 421954
rect 528326 421398 528562 421634
rect 528646 421398 528882 421634
rect 528326 385718 528562 385954
rect 528646 385718 528882 385954
rect 528326 385398 528562 385634
rect 528646 385398 528882 385634
rect 528326 349718 528562 349954
rect 528646 349718 528882 349954
rect 528326 349398 528562 349634
rect 528646 349398 528882 349634
rect 528326 313718 528562 313954
rect 528646 313718 528882 313954
rect 528326 313398 528562 313634
rect 528646 313398 528882 313634
rect 528326 277718 528562 277954
rect 528646 277718 528882 277954
rect 528326 277398 528562 277634
rect 528646 277398 528882 277634
rect 528326 241718 528562 241954
rect 528646 241718 528882 241954
rect 528326 241398 528562 241634
rect 528646 241398 528882 241634
rect 528326 205718 528562 205954
rect 528646 205718 528882 205954
rect 528326 205398 528562 205634
rect 528646 205398 528882 205634
rect 528326 169718 528562 169954
rect 528646 169718 528882 169954
rect 528326 169398 528562 169634
rect 528646 169398 528882 169634
rect 528326 133718 528562 133954
rect 528646 133718 528882 133954
rect 528326 133398 528562 133634
rect 528646 133398 528882 133634
rect 528326 97718 528562 97954
rect 528646 97718 528882 97954
rect 528326 97398 528562 97634
rect 528646 97398 528882 97634
rect 528326 61718 528562 61954
rect 528646 61718 528882 61954
rect 528326 61398 528562 61634
rect 528646 61398 528882 61634
rect 528326 25718 528562 25954
rect 528646 25718 528882 25954
rect 528326 25398 528562 25634
rect 528646 25398 528882 25634
rect 528326 -5382 528562 -5146
rect 528646 -5382 528882 -5146
rect 528326 -5702 528562 -5466
rect 528646 -5702 528882 -5466
rect 532826 710362 533062 710598
rect 533146 710362 533382 710598
rect 532826 710042 533062 710278
rect 533146 710042 533382 710278
rect 532826 678218 533062 678454
rect 533146 678218 533382 678454
rect 532826 677898 533062 678134
rect 533146 677898 533382 678134
rect 532826 642218 533062 642454
rect 533146 642218 533382 642454
rect 532826 641898 533062 642134
rect 533146 641898 533382 642134
rect 532826 606218 533062 606454
rect 533146 606218 533382 606454
rect 532826 605898 533062 606134
rect 533146 605898 533382 606134
rect 532826 570218 533062 570454
rect 533146 570218 533382 570454
rect 532826 569898 533062 570134
rect 533146 569898 533382 570134
rect 532826 534218 533062 534454
rect 533146 534218 533382 534454
rect 532826 533898 533062 534134
rect 533146 533898 533382 534134
rect 532826 498218 533062 498454
rect 533146 498218 533382 498454
rect 532826 497898 533062 498134
rect 533146 497898 533382 498134
rect 532826 462218 533062 462454
rect 533146 462218 533382 462454
rect 532826 461898 533062 462134
rect 533146 461898 533382 462134
rect 532826 426218 533062 426454
rect 533146 426218 533382 426454
rect 532826 425898 533062 426134
rect 533146 425898 533382 426134
rect 532826 390218 533062 390454
rect 533146 390218 533382 390454
rect 532826 389898 533062 390134
rect 533146 389898 533382 390134
rect 532826 354218 533062 354454
rect 533146 354218 533382 354454
rect 532826 353898 533062 354134
rect 533146 353898 533382 354134
rect 532826 318218 533062 318454
rect 533146 318218 533382 318454
rect 532826 317898 533062 318134
rect 533146 317898 533382 318134
rect 532826 282218 533062 282454
rect 533146 282218 533382 282454
rect 532826 281898 533062 282134
rect 533146 281898 533382 282134
rect 532826 246218 533062 246454
rect 533146 246218 533382 246454
rect 532826 245898 533062 246134
rect 533146 245898 533382 246134
rect 532826 210218 533062 210454
rect 533146 210218 533382 210454
rect 532826 209898 533062 210134
rect 533146 209898 533382 210134
rect 532826 174218 533062 174454
rect 533146 174218 533382 174454
rect 532826 173898 533062 174134
rect 533146 173898 533382 174134
rect 532826 138218 533062 138454
rect 533146 138218 533382 138454
rect 532826 137898 533062 138134
rect 533146 137898 533382 138134
rect 532826 102218 533062 102454
rect 533146 102218 533382 102454
rect 532826 101898 533062 102134
rect 533146 101898 533382 102134
rect 532826 66218 533062 66454
rect 533146 66218 533382 66454
rect 532826 65898 533062 66134
rect 533146 65898 533382 66134
rect 532826 30218 533062 30454
rect 533146 30218 533382 30454
rect 532826 29898 533062 30134
rect 533146 29898 533382 30134
rect 532826 -6342 533062 -6106
rect 533146 -6342 533382 -6106
rect 532826 -6662 533062 -6426
rect 533146 -6662 533382 -6426
rect 537326 711322 537562 711558
rect 537646 711322 537882 711558
rect 537326 711002 537562 711238
rect 537646 711002 537882 711238
rect 537326 682718 537562 682954
rect 537646 682718 537882 682954
rect 537326 682398 537562 682634
rect 537646 682398 537882 682634
rect 537326 646718 537562 646954
rect 537646 646718 537882 646954
rect 537326 646398 537562 646634
rect 537646 646398 537882 646634
rect 537326 610718 537562 610954
rect 537646 610718 537882 610954
rect 537326 610398 537562 610634
rect 537646 610398 537882 610634
rect 537326 574718 537562 574954
rect 537646 574718 537882 574954
rect 537326 574398 537562 574634
rect 537646 574398 537882 574634
rect 537326 538718 537562 538954
rect 537646 538718 537882 538954
rect 537326 538398 537562 538634
rect 537646 538398 537882 538634
rect 537326 502718 537562 502954
rect 537646 502718 537882 502954
rect 537326 502398 537562 502634
rect 537646 502398 537882 502634
rect 537326 466718 537562 466954
rect 537646 466718 537882 466954
rect 537326 466398 537562 466634
rect 537646 466398 537882 466634
rect 537326 430718 537562 430954
rect 537646 430718 537882 430954
rect 537326 430398 537562 430634
rect 537646 430398 537882 430634
rect 537326 394718 537562 394954
rect 537646 394718 537882 394954
rect 537326 394398 537562 394634
rect 537646 394398 537882 394634
rect 537326 358718 537562 358954
rect 537646 358718 537882 358954
rect 537326 358398 537562 358634
rect 537646 358398 537882 358634
rect 537326 322718 537562 322954
rect 537646 322718 537882 322954
rect 537326 322398 537562 322634
rect 537646 322398 537882 322634
rect 537326 286718 537562 286954
rect 537646 286718 537882 286954
rect 537326 286398 537562 286634
rect 537646 286398 537882 286634
rect 537326 250718 537562 250954
rect 537646 250718 537882 250954
rect 537326 250398 537562 250634
rect 537646 250398 537882 250634
rect 537326 214718 537562 214954
rect 537646 214718 537882 214954
rect 537326 214398 537562 214634
rect 537646 214398 537882 214634
rect 537326 178718 537562 178954
rect 537646 178718 537882 178954
rect 537326 178398 537562 178634
rect 537646 178398 537882 178634
rect 537326 142718 537562 142954
rect 537646 142718 537882 142954
rect 537326 142398 537562 142634
rect 537646 142398 537882 142634
rect 537326 106718 537562 106954
rect 537646 106718 537882 106954
rect 537326 106398 537562 106634
rect 537646 106398 537882 106634
rect 537326 70718 537562 70954
rect 537646 70718 537882 70954
rect 537326 70398 537562 70634
rect 537646 70398 537882 70634
rect 537326 34718 537562 34954
rect 537646 34718 537882 34954
rect 537326 34398 537562 34634
rect 537646 34398 537882 34634
rect 537326 -7302 537562 -7066
rect 537646 -7302 537882 -7066
rect 537326 -7622 537562 -7386
rect 537646 -7622 537882 -7386
rect 541826 704602 542062 704838
rect 542146 704602 542382 704838
rect 541826 704282 542062 704518
rect 542146 704282 542382 704518
rect 541826 687218 542062 687454
rect 542146 687218 542382 687454
rect 541826 686898 542062 687134
rect 542146 686898 542382 687134
rect 541826 651218 542062 651454
rect 542146 651218 542382 651454
rect 541826 650898 542062 651134
rect 542146 650898 542382 651134
rect 541826 615218 542062 615454
rect 542146 615218 542382 615454
rect 541826 614898 542062 615134
rect 542146 614898 542382 615134
rect 541826 579218 542062 579454
rect 542146 579218 542382 579454
rect 541826 578898 542062 579134
rect 542146 578898 542382 579134
rect 541826 543218 542062 543454
rect 542146 543218 542382 543454
rect 541826 542898 542062 543134
rect 542146 542898 542382 543134
rect 541826 507218 542062 507454
rect 542146 507218 542382 507454
rect 541826 506898 542062 507134
rect 542146 506898 542382 507134
rect 541826 471218 542062 471454
rect 542146 471218 542382 471454
rect 541826 470898 542062 471134
rect 542146 470898 542382 471134
rect 541826 435218 542062 435454
rect 542146 435218 542382 435454
rect 541826 434898 542062 435134
rect 542146 434898 542382 435134
rect 541826 399218 542062 399454
rect 542146 399218 542382 399454
rect 541826 398898 542062 399134
rect 542146 398898 542382 399134
rect 541826 363218 542062 363454
rect 542146 363218 542382 363454
rect 541826 362898 542062 363134
rect 542146 362898 542382 363134
rect 541826 327218 542062 327454
rect 542146 327218 542382 327454
rect 541826 326898 542062 327134
rect 542146 326898 542382 327134
rect 541826 291218 542062 291454
rect 542146 291218 542382 291454
rect 541826 290898 542062 291134
rect 542146 290898 542382 291134
rect 541826 255218 542062 255454
rect 542146 255218 542382 255454
rect 541826 254898 542062 255134
rect 542146 254898 542382 255134
rect 541826 219218 542062 219454
rect 542146 219218 542382 219454
rect 541826 218898 542062 219134
rect 542146 218898 542382 219134
rect 541826 183218 542062 183454
rect 542146 183218 542382 183454
rect 541826 182898 542062 183134
rect 542146 182898 542382 183134
rect 541826 147218 542062 147454
rect 542146 147218 542382 147454
rect 541826 146898 542062 147134
rect 542146 146898 542382 147134
rect 541826 111218 542062 111454
rect 542146 111218 542382 111454
rect 541826 110898 542062 111134
rect 542146 110898 542382 111134
rect 541826 75218 542062 75454
rect 542146 75218 542382 75454
rect 541826 74898 542062 75134
rect 542146 74898 542382 75134
rect 541826 39218 542062 39454
rect 542146 39218 542382 39454
rect 541826 38898 542062 39134
rect 542146 38898 542382 39134
rect 541826 3218 542062 3454
rect 542146 3218 542382 3454
rect 541826 2898 542062 3134
rect 542146 2898 542382 3134
rect 541826 -582 542062 -346
rect 542146 -582 542382 -346
rect 541826 -902 542062 -666
rect 542146 -902 542382 -666
rect 546326 705562 546562 705798
rect 546646 705562 546882 705798
rect 546326 705242 546562 705478
rect 546646 705242 546882 705478
rect 546326 691718 546562 691954
rect 546646 691718 546882 691954
rect 546326 691398 546562 691634
rect 546646 691398 546882 691634
rect 546326 655718 546562 655954
rect 546646 655718 546882 655954
rect 546326 655398 546562 655634
rect 546646 655398 546882 655634
rect 546326 619718 546562 619954
rect 546646 619718 546882 619954
rect 546326 619398 546562 619634
rect 546646 619398 546882 619634
rect 546326 583718 546562 583954
rect 546646 583718 546882 583954
rect 546326 583398 546562 583634
rect 546646 583398 546882 583634
rect 546326 547718 546562 547954
rect 546646 547718 546882 547954
rect 546326 547398 546562 547634
rect 546646 547398 546882 547634
rect 546326 511718 546562 511954
rect 546646 511718 546882 511954
rect 546326 511398 546562 511634
rect 546646 511398 546882 511634
rect 546326 475718 546562 475954
rect 546646 475718 546882 475954
rect 546326 475398 546562 475634
rect 546646 475398 546882 475634
rect 546326 439718 546562 439954
rect 546646 439718 546882 439954
rect 546326 439398 546562 439634
rect 546646 439398 546882 439634
rect 546326 403718 546562 403954
rect 546646 403718 546882 403954
rect 546326 403398 546562 403634
rect 546646 403398 546882 403634
rect 546326 367718 546562 367954
rect 546646 367718 546882 367954
rect 546326 367398 546562 367634
rect 546646 367398 546882 367634
rect 546326 331718 546562 331954
rect 546646 331718 546882 331954
rect 546326 331398 546562 331634
rect 546646 331398 546882 331634
rect 546326 295718 546562 295954
rect 546646 295718 546882 295954
rect 546326 295398 546562 295634
rect 546646 295398 546882 295634
rect 546326 259718 546562 259954
rect 546646 259718 546882 259954
rect 546326 259398 546562 259634
rect 546646 259398 546882 259634
rect 546326 223718 546562 223954
rect 546646 223718 546882 223954
rect 546326 223398 546562 223634
rect 546646 223398 546882 223634
rect 546326 187718 546562 187954
rect 546646 187718 546882 187954
rect 546326 187398 546562 187634
rect 546646 187398 546882 187634
rect 546326 151718 546562 151954
rect 546646 151718 546882 151954
rect 546326 151398 546562 151634
rect 546646 151398 546882 151634
rect 546326 115718 546562 115954
rect 546646 115718 546882 115954
rect 546326 115398 546562 115634
rect 546646 115398 546882 115634
rect 546326 79718 546562 79954
rect 546646 79718 546882 79954
rect 546326 79398 546562 79634
rect 546646 79398 546882 79634
rect 546326 43718 546562 43954
rect 546646 43718 546882 43954
rect 546326 43398 546562 43634
rect 546646 43398 546882 43634
rect 546326 7718 546562 7954
rect 546646 7718 546882 7954
rect 546326 7398 546562 7634
rect 546646 7398 546882 7634
rect 546326 -1542 546562 -1306
rect 546646 -1542 546882 -1306
rect 546326 -1862 546562 -1626
rect 546646 -1862 546882 -1626
rect 550826 706522 551062 706758
rect 551146 706522 551382 706758
rect 550826 706202 551062 706438
rect 551146 706202 551382 706438
rect 550826 696218 551062 696454
rect 551146 696218 551382 696454
rect 550826 695898 551062 696134
rect 551146 695898 551382 696134
rect 550826 660218 551062 660454
rect 551146 660218 551382 660454
rect 550826 659898 551062 660134
rect 551146 659898 551382 660134
rect 550826 624218 551062 624454
rect 551146 624218 551382 624454
rect 550826 623898 551062 624134
rect 551146 623898 551382 624134
rect 550826 588218 551062 588454
rect 551146 588218 551382 588454
rect 550826 587898 551062 588134
rect 551146 587898 551382 588134
rect 550826 552218 551062 552454
rect 551146 552218 551382 552454
rect 550826 551898 551062 552134
rect 551146 551898 551382 552134
rect 550826 516218 551062 516454
rect 551146 516218 551382 516454
rect 550826 515898 551062 516134
rect 551146 515898 551382 516134
rect 550826 480218 551062 480454
rect 551146 480218 551382 480454
rect 550826 479898 551062 480134
rect 551146 479898 551382 480134
rect 550826 444218 551062 444454
rect 551146 444218 551382 444454
rect 550826 443898 551062 444134
rect 551146 443898 551382 444134
rect 550826 408218 551062 408454
rect 551146 408218 551382 408454
rect 550826 407898 551062 408134
rect 551146 407898 551382 408134
rect 550826 372218 551062 372454
rect 551146 372218 551382 372454
rect 550826 371898 551062 372134
rect 551146 371898 551382 372134
rect 550826 336218 551062 336454
rect 551146 336218 551382 336454
rect 550826 335898 551062 336134
rect 551146 335898 551382 336134
rect 550826 300218 551062 300454
rect 551146 300218 551382 300454
rect 550826 299898 551062 300134
rect 551146 299898 551382 300134
rect 550826 264218 551062 264454
rect 551146 264218 551382 264454
rect 550826 263898 551062 264134
rect 551146 263898 551382 264134
rect 550826 228218 551062 228454
rect 551146 228218 551382 228454
rect 550826 227898 551062 228134
rect 551146 227898 551382 228134
rect 550826 192218 551062 192454
rect 551146 192218 551382 192454
rect 550826 191898 551062 192134
rect 551146 191898 551382 192134
rect 550826 156218 551062 156454
rect 551146 156218 551382 156454
rect 550826 155898 551062 156134
rect 551146 155898 551382 156134
rect 550826 120218 551062 120454
rect 551146 120218 551382 120454
rect 550826 119898 551062 120134
rect 551146 119898 551382 120134
rect 550826 84218 551062 84454
rect 551146 84218 551382 84454
rect 550826 83898 551062 84134
rect 551146 83898 551382 84134
rect 550826 48218 551062 48454
rect 551146 48218 551382 48454
rect 550826 47898 551062 48134
rect 551146 47898 551382 48134
rect 550826 12218 551062 12454
rect 551146 12218 551382 12454
rect 550826 11898 551062 12134
rect 551146 11898 551382 12134
rect 550826 -2502 551062 -2266
rect 551146 -2502 551382 -2266
rect 550826 -2822 551062 -2586
rect 551146 -2822 551382 -2586
rect 555326 707482 555562 707718
rect 555646 707482 555882 707718
rect 555326 707162 555562 707398
rect 555646 707162 555882 707398
rect 555326 700718 555562 700954
rect 555646 700718 555882 700954
rect 555326 700398 555562 700634
rect 555646 700398 555882 700634
rect 555326 664718 555562 664954
rect 555646 664718 555882 664954
rect 555326 664398 555562 664634
rect 555646 664398 555882 664634
rect 555326 628718 555562 628954
rect 555646 628718 555882 628954
rect 555326 628398 555562 628634
rect 555646 628398 555882 628634
rect 555326 592718 555562 592954
rect 555646 592718 555882 592954
rect 555326 592398 555562 592634
rect 555646 592398 555882 592634
rect 555326 556718 555562 556954
rect 555646 556718 555882 556954
rect 555326 556398 555562 556634
rect 555646 556398 555882 556634
rect 555326 520718 555562 520954
rect 555646 520718 555882 520954
rect 555326 520398 555562 520634
rect 555646 520398 555882 520634
rect 555326 484718 555562 484954
rect 555646 484718 555882 484954
rect 555326 484398 555562 484634
rect 555646 484398 555882 484634
rect 555326 448718 555562 448954
rect 555646 448718 555882 448954
rect 555326 448398 555562 448634
rect 555646 448398 555882 448634
rect 555326 412718 555562 412954
rect 555646 412718 555882 412954
rect 555326 412398 555562 412634
rect 555646 412398 555882 412634
rect 555326 376718 555562 376954
rect 555646 376718 555882 376954
rect 555326 376398 555562 376634
rect 555646 376398 555882 376634
rect 555326 340718 555562 340954
rect 555646 340718 555882 340954
rect 555326 340398 555562 340634
rect 555646 340398 555882 340634
rect 555326 304718 555562 304954
rect 555646 304718 555882 304954
rect 555326 304398 555562 304634
rect 555646 304398 555882 304634
rect 555326 268718 555562 268954
rect 555646 268718 555882 268954
rect 555326 268398 555562 268634
rect 555646 268398 555882 268634
rect 555326 232718 555562 232954
rect 555646 232718 555882 232954
rect 555326 232398 555562 232634
rect 555646 232398 555882 232634
rect 555326 196718 555562 196954
rect 555646 196718 555882 196954
rect 555326 196398 555562 196634
rect 555646 196398 555882 196634
rect 555326 160718 555562 160954
rect 555646 160718 555882 160954
rect 555326 160398 555562 160634
rect 555646 160398 555882 160634
rect 555326 124718 555562 124954
rect 555646 124718 555882 124954
rect 555326 124398 555562 124634
rect 555646 124398 555882 124634
rect 555326 88718 555562 88954
rect 555646 88718 555882 88954
rect 555326 88398 555562 88634
rect 555646 88398 555882 88634
rect 555326 52718 555562 52954
rect 555646 52718 555882 52954
rect 555326 52398 555562 52634
rect 555646 52398 555882 52634
rect 555326 16718 555562 16954
rect 555646 16718 555882 16954
rect 555326 16398 555562 16634
rect 555646 16398 555882 16634
rect 555326 -3462 555562 -3226
rect 555646 -3462 555882 -3226
rect 555326 -3782 555562 -3546
rect 555646 -3782 555882 -3546
rect 559826 708442 560062 708678
rect 560146 708442 560382 708678
rect 559826 708122 560062 708358
rect 560146 708122 560382 708358
rect 559826 669218 560062 669454
rect 560146 669218 560382 669454
rect 559826 668898 560062 669134
rect 560146 668898 560382 669134
rect 559826 633218 560062 633454
rect 560146 633218 560382 633454
rect 559826 632898 560062 633134
rect 560146 632898 560382 633134
rect 559826 597218 560062 597454
rect 560146 597218 560382 597454
rect 559826 596898 560062 597134
rect 560146 596898 560382 597134
rect 559826 561218 560062 561454
rect 560146 561218 560382 561454
rect 559826 560898 560062 561134
rect 560146 560898 560382 561134
rect 559826 525218 560062 525454
rect 560146 525218 560382 525454
rect 559826 524898 560062 525134
rect 560146 524898 560382 525134
rect 559826 489218 560062 489454
rect 560146 489218 560382 489454
rect 559826 488898 560062 489134
rect 560146 488898 560382 489134
rect 559826 453218 560062 453454
rect 560146 453218 560382 453454
rect 559826 452898 560062 453134
rect 560146 452898 560382 453134
rect 559826 417218 560062 417454
rect 560146 417218 560382 417454
rect 559826 416898 560062 417134
rect 560146 416898 560382 417134
rect 559826 381218 560062 381454
rect 560146 381218 560382 381454
rect 559826 380898 560062 381134
rect 560146 380898 560382 381134
rect 559826 345218 560062 345454
rect 560146 345218 560382 345454
rect 559826 344898 560062 345134
rect 560146 344898 560382 345134
rect 559826 309218 560062 309454
rect 560146 309218 560382 309454
rect 559826 308898 560062 309134
rect 560146 308898 560382 309134
rect 559826 273218 560062 273454
rect 560146 273218 560382 273454
rect 559826 272898 560062 273134
rect 560146 272898 560382 273134
rect 559826 237218 560062 237454
rect 560146 237218 560382 237454
rect 559826 236898 560062 237134
rect 560146 236898 560382 237134
rect 559826 201218 560062 201454
rect 560146 201218 560382 201454
rect 559826 200898 560062 201134
rect 560146 200898 560382 201134
rect 559826 165218 560062 165454
rect 560146 165218 560382 165454
rect 559826 164898 560062 165134
rect 560146 164898 560382 165134
rect 559826 129218 560062 129454
rect 560146 129218 560382 129454
rect 559826 128898 560062 129134
rect 560146 128898 560382 129134
rect 559826 93218 560062 93454
rect 560146 93218 560382 93454
rect 559826 92898 560062 93134
rect 560146 92898 560382 93134
rect 559826 57218 560062 57454
rect 560146 57218 560382 57454
rect 559826 56898 560062 57134
rect 560146 56898 560382 57134
rect 559826 21218 560062 21454
rect 560146 21218 560382 21454
rect 559826 20898 560062 21134
rect 560146 20898 560382 21134
rect 559826 -4422 560062 -4186
rect 560146 -4422 560382 -4186
rect 559826 -4742 560062 -4506
rect 560146 -4742 560382 -4506
rect 564326 709402 564562 709638
rect 564646 709402 564882 709638
rect 564326 709082 564562 709318
rect 564646 709082 564882 709318
rect 564326 673718 564562 673954
rect 564646 673718 564882 673954
rect 564326 673398 564562 673634
rect 564646 673398 564882 673634
rect 564326 637718 564562 637954
rect 564646 637718 564882 637954
rect 564326 637398 564562 637634
rect 564646 637398 564882 637634
rect 564326 601718 564562 601954
rect 564646 601718 564882 601954
rect 564326 601398 564562 601634
rect 564646 601398 564882 601634
rect 564326 565718 564562 565954
rect 564646 565718 564882 565954
rect 564326 565398 564562 565634
rect 564646 565398 564882 565634
rect 564326 529718 564562 529954
rect 564646 529718 564882 529954
rect 564326 529398 564562 529634
rect 564646 529398 564882 529634
rect 564326 493718 564562 493954
rect 564646 493718 564882 493954
rect 564326 493398 564562 493634
rect 564646 493398 564882 493634
rect 564326 457718 564562 457954
rect 564646 457718 564882 457954
rect 564326 457398 564562 457634
rect 564646 457398 564882 457634
rect 564326 421718 564562 421954
rect 564646 421718 564882 421954
rect 564326 421398 564562 421634
rect 564646 421398 564882 421634
rect 564326 385718 564562 385954
rect 564646 385718 564882 385954
rect 564326 385398 564562 385634
rect 564646 385398 564882 385634
rect 564326 349718 564562 349954
rect 564646 349718 564882 349954
rect 564326 349398 564562 349634
rect 564646 349398 564882 349634
rect 564326 313718 564562 313954
rect 564646 313718 564882 313954
rect 564326 313398 564562 313634
rect 564646 313398 564882 313634
rect 564326 277718 564562 277954
rect 564646 277718 564882 277954
rect 564326 277398 564562 277634
rect 564646 277398 564882 277634
rect 564326 241718 564562 241954
rect 564646 241718 564882 241954
rect 564326 241398 564562 241634
rect 564646 241398 564882 241634
rect 564326 205718 564562 205954
rect 564646 205718 564882 205954
rect 564326 205398 564562 205634
rect 564646 205398 564882 205634
rect 564326 169718 564562 169954
rect 564646 169718 564882 169954
rect 564326 169398 564562 169634
rect 564646 169398 564882 169634
rect 564326 133718 564562 133954
rect 564646 133718 564882 133954
rect 564326 133398 564562 133634
rect 564646 133398 564882 133634
rect 564326 97718 564562 97954
rect 564646 97718 564882 97954
rect 564326 97398 564562 97634
rect 564646 97398 564882 97634
rect 564326 61718 564562 61954
rect 564646 61718 564882 61954
rect 564326 61398 564562 61634
rect 564646 61398 564882 61634
rect 564326 25718 564562 25954
rect 564646 25718 564882 25954
rect 564326 25398 564562 25634
rect 564646 25398 564882 25634
rect 564326 -5382 564562 -5146
rect 564646 -5382 564882 -5146
rect 564326 -5702 564562 -5466
rect 564646 -5702 564882 -5466
rect 568826 710362 569062 710598
rect 569146 710362 569382 710598
rect 568826 710042 569062 710278
rect 569146 710042 569382 710278
rect 568826 678218 569062 678454
rect 569146 678218 569382 678454
rect 568826 677898 569062 678134
rect 569146 677898 569382 678134
rect 568826 642218 569062 642454
rect 569146 642218 569382 642454
rect 568826 641898 569062 642134
rect 569146 641898 569382 642134
rect 568826 606218 569062 606454
rect 569146 606218 569382 606454
rect 568826 605898 569062 606134
rect 569146 605898 569382 606134
rect 568826 570218 569062 570454
rect 569146 570218 569382 570454
rect 568826 569898 569062 570134
rect 569146 569898 569382 570134
rect 568826 534218 569062 534454
rect 569146 534218 569382 534454
rect 568826 533898 569062 534134
rect 569146 533898 569382 534134
rect 568826 498218 569062 498454
rect 569146 498218 569382 498454
rect 568826 497898 569062 498134
rect 569146 497898 569382 498134
rect 568826 462218 569062 462454
rect 569146 462218 569382 462454
rect 568826 461898 569062 462134
rect 569146 461898 569382 462134
rect 568826 426218 569062 426454
rect 569146 426218 569382 426454
rect 568826 425898 569062 426134
rect 569146 425898 569382 426134
rect 568826 390218 569062 390454
rect 569146 390218 569382 390454
rect 568826 389898 569062 390134
rect 569146 389898 569382 390134
rect 568826 354218 569062 354454
rect 569146 354218 569382 354454
rect 568826 353898 569062 354134
rect 569146 353898 569382 354134
rect 568826 318218 569062 318454
rect 569146 318218 569382 318454
rect 568826 317898 569062 318134
rect 569146 317898 569382 318134
rect 568826 282218 569062 282454
rect 569146 282218 569382 282454
rect 568826 281898 569062 282134
rect 569146 281898 569382 282134
rect 568826 246218 569062 246454
rect 569146 246218 569382 246454
rect 568826 245898 569062 246134
rect 569146 245898 569382 246134
rect 568826 210218 569062 210454
rect 569146 210218 569382 210454
rect 568826 209898 569062 210134
rect 569146 209898 569382 210134
rect 568826 174218 569062 174454
rect 569146 174218 569382 174454
rect 568826 173898 569062 174134
rect 569146 173898 569382 174134
rect 568826 138218 569062 138454
rect 569146 138218 569382 138454
rect 568826 137898 569062 138134
rect 569146 137898 569382 138134
rect 568826 102218 569062 102454
rect 569146 102218 569382 102454
rect 568826 101898 569062 102134
rect 569146 101898 569382 102134
rect 568826 66218 569062 66454
rect 569146 66218 569382 66454
rect 568826 65898 569062 66134
rect 569146 65898 569382 66134
rect 568826 30218 569062 30454
rect 569146 30218 569382 30454
rect 568826 29898 569062 30134
rect 569146 29898 569382 30134
rect 568826 -6342 569062 -6106
rect 569146 -6342 569382 -6106
rect 568826 -6662 569062 -6426
rect 569146 -6662 569382 -6426
rect 573326 711322 573562 711558
rect 573646 711322 573882 711558
rect 573326 711002 573562 711238
rect 573646 711002 573882 711238
rect 573326 682718 573562 682954
rect 573646 682718 573882 682954
rect 573326 682398 573562 682634
rect 573646 682398 573882 682634
rect 573326 646718 573562 646954
rect 573646 646718 573882 646954
rect 573326 646398 573562 646634
rect 573646 646398 573882 646634
rect 573326 610718 573562 610954
rect 573646 610718 573882 610954
rect 573326 610398 573562 610634
rect 573646 610398 573882 610634
rect 573326 574718 573562 574954
rect 573646 574718 573882 574954
rect 573326 574398 573562 574634
rect 573646 574398 573882 574634
rect 573326 538718 573562 538954
rect 573646 538718 573882 538954
rect 573326 538398 573562 538634
rect 573646 538398 573882 538634
rect 573326 502718 573562 502954
rect 573646 502718 573882 502954
rect 573326 502398 573562 502634
rect 573646 502398 573882 502634
rect 573326 466718 573562 466954
rect 573646 466718 573882 466954
rect 573326 466398 573562 466634
rect 573646 466398 573882 466634
rect 573326 430718 573562 430954
rect 573646 430718 573882 430954
rect 573326 430398 573562 430634
rect 573646 430398 573882 430634
rect 573326 394718 573562 394954
rect 573646 394718 573882 394954
rect 573326 394398 573562 394634
rect 573646 394398 573882 394634
rect 573326 358718 573562 358954
rect 573646 358718 573882 358954
rect 573326 358398 573562 358634
rect 573646 358398 573882 358634
rect 573326 322718 573562 322954
rect 573646 322718 573882 322954
rect 573326 322398 573562 322634
rect 573646 322398 573882 322634
rect 573326 286718 573562 286954
rect 573646 286718 573882 286954
rect 573326 286398 573562 286634
rect 573646 286398 573882 286634
rect 573326 250718 573562 250954
rect 573646 250718 573882 250954
rect 573326 250398 573562 250634
rect 573646 250398 573882 250634
rect 573326 214718 573562 214954
rect 573646 214718 573882 214954
rect 573326 214398 573562 214634
rect 573646 214398 573882 214634
rect 573326 178718 573562 178954
rect 573646 178718 573882 178954
rect 573326 178398 573562 178634
rect 573646 178398 573882 178634
rect 573326 142718 573562 142954
rect 573646 142718 573882 142954
rect 573326 142398 573562 142634
rect 573646 142398 573882 142634
rect 573326 106718 573562 106954
rect 573646 106718 573882 106954
rect 573326 106398 573562 106634
rect 573646 106398 573882 106634
rect 573326 70718 573562 70954
rect 573646 70718 573882 70954
rect 573326 70398 573562 70634
rect 573646 70398 573882 70634
rect 573326 34718 573562 34954
rect 573646 34718 573882 34954
rect 573326 34398 573562 34634
rect 573646 34398 573882 34634
rect 573326 -7302 573562 -7066
rect 573646 -7302 573882 -7066
rect 573326 -7622 573562 -7386
rect 573646 -7622 573882 -7386
rect 577826 704602 578062 704838
rect 578146 704602 578382 704838
rect 577826 704282 578062 704518
rect 578146 704282 578382 704518
rect 577826 687218 578062 687454
rect 578146 687218 578382 687454
rect 577826 686898 578062 687134
rect 578146 686898 578382 687134
rect 577826 651218 578062 651454
rect 578146 651218 578382 651454
rect 577826 650898 578062 651134
rect 578146 650898 578382 651134
rect 577826 615218 578062 615454
rect 578146 615218 578382 615454
rect 577826 614898 578062 615134
rect 578146 614898 578382 615134
rect 577826 579218 578062 579454
rect 578146 579218 578382 579454
rect 577826 578898 578062 579134
rect 578146 578898 578382 579134
rect 577826 543218 578062 543454
rect 578146 543218 578382 543454
rect 577826 542898 578062 543134
rect 578146 542898 578382 543134
rect 577826 507218 578062 507454
rect 578146 507218 578382 507454
rect 577826 506898 578062 507134
rect 578146 506898 578382 507134
rect 577826 471218 578062 471454
rect 578146 471218 578382 471454
rect 577826 470898 578062 471134
rect 578146 470898 578382 471134
rect 577826 435218 578062 435454
rect 578146 435218 578382 435454
rect 577826 434898 578062 435134
rect 578146 434898 578382 435134
rect 577826 399218 578062 399454
rect 578146 399218 578382 399454
rect 577826 398898 578062 399134
rect 578146 398898 578382 399134
rect 577826 363218 578062 363454
rect 578146 363218 578382 363454
rect 577826 362898 578062 363134
rect 578146 362898 578382 363134
rect 577826 327218 578062 327454
rect 578146 327218 578382 327454
rect 577826 326898 578062 327134
rect 578146 326898 578382 327134
rect 577826 291218 578062 291454
rect 578146 291218 578382 291454
rect 577826 290898 578062 291134
rect 578146 290898 578382 291134
rect 577826 255218 578062 255454
rect 578146 255218 578382 255454
rect 577826 254898 578062 255134
rect 578146 254898 578382 255134
rect 577826 219218 578062 219454
rect 578146 219218 578382 219454
rect 577826 218898 578062 219134
rect 578146 218898 578382 219134
rect 577826 183218 578062 183454
rect 578146 183218 578382 183454
rect 577826 182898 578062 183134
rect 578146 182898 578382 183134
rect 577826 147218 578062 147454
rect 578146 147218 578382 147454
rect 577826 146898 578062 147134
rect 578146 146898 578382 147134
rect 577826 111218 578062 111454
rect 578146 111218 578382 111454
rect 577826 110898 578062 111134
rect 578146 110898 578382 111134
rect 577826 75218 578062 75454
rect 578146 75218 578382 75454
rect 577826 74898 578062 75134
rect 578146 74898 578382 75134
rect 577826 39218 578062 39454
rect 578146 39218 578382 39454
rect 577826 38898 578062 39134
rect 578146 38898 578382 39134
rect 577826 3218 578062 3454
rect 578146 3218 578382 3454
rect 577826 2898 578062 3134
rect 578146 2898 578382 3134
rect 577826 -582 578062 -346
rect 578146 -582 578382 -346
rect 577826 -902 578062 -666
rect 578146 -902 578382 -666
rect 592062 711322 592298 711558
rect 592382 711322 592618 711558
rect 592062 711002 592298 711238
rect 592382 711002 592618 711238
rect 591102 710362 591338 710598
rect 591422 710362 591658 710598
rect 591102 710042 591338 710278
rect 591422 710042 591658 710278
rect 590142 709402 590378 709638
rect 590462 709402 590698 709638
rect 590142 709082 590378 709318
rect 590462 709082 590698 709318
rect 589182 708442 589418 708678
rect 589502 708442 589738 708678
rect 589182 708122 589418 708358
rect 589502 708122 589738 708358
rect 588222 707482 588458 707718
rect 588542 707482 588778 707718
rect 588222 707162 588458 707398
rect 588542 707162 588778 707398
rect 587262 706522 587498 706758
rect 587582 706522 587818 706758
rect 587262 706202 587498 706438
rect 587582 706202 587818 706438
rect 582326 705562 582562 705798
rect 582646 705562 582882 705798
rect 582326 705242 582562 705478
rect 582646 705242 582882 705478
rect 586302 705562 586538 705798
rect 586622 705562 586858 705798
rect 586302 705242 586538 705478
rect 586622 705242 586858 705478
rect 582326 691718 582562 691954
rect 582646 691718 582882 691954
rect 582326 691398 582562 691634
rect 582646 691398 582882 691634
rect 582326 655718 582562 655954
rect 582646 655718 582882 655954
rect 582326 655398 582562 655634
rect 582646 655398 582882 655634
rect 582326 619718 582562 619954
rect 582646 619718 582882 619954
rect 582326 619398 582562 619634
rect 582646 619398 582882 619634
rect 582326 583718 582562 583954
rect 582646 583718 582882 583954
rect 582326 583398 582562 583634
rect 582646 583398 582882 583634
rect 582326 547718 582562 547954
rect 582646 547718 582882 547954
rect 582326 547398 582562 547634
rect 582646 547398 582882 547634
rect 582326 511718 582562 511954
rect 582646 511718 582882 511954
rect 582326 511398 582562 511634
rect 582646 511398 582882 511634
rect 582326 475718 582562 475954
rect 582646 475718 582882 475954
rect 582326 475398 582562 475634
rect 582646 475398 582882 475634
rect 582326 439718 582562 439954
rect 582646 439718 582882 439954
rect 582326 439398 582562 439634
rect 582646 439398 582882 439634
rect 582326 403718 582562 403954
rect 582646 403718 582882 403954
rect 582326 403398 582562 403634
rect 582646 403398 582882 403634
rect 582326 367718 582562 367954
rect 582646 367718 582882 367954
rect 582326 367398 582562 367634
rect 582646 367398 582882 367634
rect 582326 331718 582562 331954
rect 582646 331718 582882 331954
rect 582326 331398 582562 331634
rect 582646 331398 582882 331634
rect 582326 295718 582562 295954
rect 582646 295718 582882 295954
rect 582326 295398 582562 295634
rect 582646 295398 582882 295634
rect 582326 259718 582562 259954
rect 582646 259718 582882 259954
rect 582326 259398 582562 259634
rect 582646 259398 582882 259634
rect 582326 223718 582562 223954
rect 582646 223718 582882 223954
rect 582326 223398 582562 223634
rect 582646 223398 582882 223634
rect 582326 187718 582562 187954
rect 582646 187718 582882 187954
rect 582326 187398 582562 187634
rect 582646 187398 582882 187634
rect 582326 151718 582562 151954
rect 582646 151718 582882 151954
rect 582326 151398 582562 151634
rect 582646 151398 582882 151634
rect 582326 115718 582562 115954
rect 582646 115718 582882 115954
rect 582326 115398 582562 115634
rect 582646 115398 582882 115634
rect 582326 79718 582562 79954
rect 582646 79718 582882 79954
rect 582326 79398 582562 79634
rect 582646 79398 582882 79634
rect 582326 43718 582562 43954
rect 582646 43718 582882 43954
rect 582326 43398 582562 43634
rect 582646 43398 582882 43634
rect 582326 7718 582562 7954
rect 582646 7718 582882 7954
rect 582326 7398 582562 7634
rect 582646 7398 582882 7634
rect 585342 704602 585578 704838
rect 585662 704602 585898 704838
rect 585342 704282 585578 704518
rect 585662 704282 585898 704518
rect 585342 687218 585578 687454
rect 585662 687218 585898 687454
rect 585342 686898 585578 687134
rect 585662 686898 585898 687134
rect 585342 651218 585578 651454
rect 585662 651218 585898 651454
rect 585342 650898 585578 651134
rect 585662 650898 585898 651134
rect 585342 615218 585578 615454
rect 585662 615218 585898 615454
rect 585342 614898 585578 615134
rect 585662 614898 585898 615134
rect 585342 579218 585578 579454
rect 585662 579218 585898 579454
rect 585342 578898 585578 579134
rect 585662 578898 585898 579134
rect 585342 543218 585578 543454
rect 585662 543218 585898 543454
rect 585342 542898 585578 543134
rect 585662 542898 585898 543134
rect 585342 507218 585578 507454
rect 585662 507218 585898 507454
rect 585342 506898 585578 507134
rect 585662 506898 585898 507134
rect 585342 471218 585578 471454
rect 585662 471218 585898 471454
rect 585342 470898 585578 471134
rect 585662 470898 585898 471134
rect 585342 435218 585578 435454
rect 585662 435218 585898 435454
rect 585342 434898 585578 435134
rect 585662 434898 585898 435134
rect 585342 399218 585578 399454
rect 585662 399218 585898 399454
rect 585342 398898 585578 399134
rect 585662 398898 585898 399134
rect 585342 363218 585578 363454
rect 585662 363218 585898 363454
rect 585342 362898 585578 363134
rect 585662 362898 585898 363134
rect 585342 327218 585578 327454
rect 585662 327218 585898 327454
rect 585342 326898 585578 327134
rect 585662 326898 585898 327134
rect 585342 291218 585578 291454
rect 585662 291218 585898 291454
rect 585342 290898 585578 291134
rect 585662 290898 585898 291134
rect 585342 255218 585578 255454
rect 585662 255218 585898 255454
rect 585342 254898 585578 255134
rect 585662 254898 585898 255134
rect 585342 219218 585578 219454
rect 585662 219218 585898 219454
rect 585342 218898 585578 219134
rect 585662 218898 585898 219134
rect 585342 183218 585578 183454
rect 585662 183218 585898 183454
rect 585342 182898 585578 183134
rect 585662 182898 585898 183134
rect 585342 147218 585578 147454
rect 585662 147218 585898 147454
rect 585342 146898 585578 147134
rect 585662 146898 585898 147134
rect 585342 111218 585578 111454
rect 585662 111218 585898 111454
rect 585342 110898 585578 111134
rect 585662 110898 585898 111134
rect 585342 75218 585578 75454
rect 585662 75218 585898 75454
rect 585342 74898 585578 75134
rect 585662 74898 585898 75134
rect 585342 39218 585578 39454
rect 585662 39218 585898 39454
rect 585342 38898 585578 39134
rect 585662 38898 585898 39134
rect 585342 3218 585578 3454
rect 585662 3218 585898 3454
rect 585342 2898 585578 3134
rect 585662 2898 585898 3134
rect 585342 -582 585578 -346
rect 585662 -582 585898 -346
rect 585342 -902 585578 -666
rect 585662 -902 585898 -666
rect 586302 691718 586538 691954
rect 586622 691718 586858 691954
rect 586302 691398 586538 691634
rect 586622 691398 586858 691634
rect 586302 655718 586538 655954
rect 586622 655718 586858 655954
rect 586302 655398 586538 655634
rect 586622 655398 586858 655634
rect 586302 619718 586538 619954
rect 586622 619718 586858 619954
rect 586302 619398 586538 619634
rect 586622 619398 586858 619634
rect 586302 583718 586538 583954
rect 586622 583718 586858 583954
rect 586302 583398 586538 583634
rect 586622 583398 586858 583634
rect 586302 547718 586538 547954
rect 586622 547718 586858 547954
rect 586302 547398 586538 547634
rect 586622 547398 586858 547634
rect 586302 511718 586538 511954
rect 586622 511718 586858 511954
rect 586302 511398 586538 511634
rect 586622 511398 586858 511634
rect 586302 475718 586538 475954
rect 586622 475718 586858 475954
rect 586302 475398 586538 475634
rect 586622 475398 586858 475634
rect 586302 439718 586538 439954
rect 586622 439718 586858 439954
rect 586302 439398 586538 439634
rect 586622 439398 586858 439634
rect 586302 403718 586538 403954
rect 586622 403718 586858 403954
rect 586302 403398 586538 403634
rect 586622 403398 586858 403634
rect 586302 367718 586538 367954
rect 586622 367718 586858 367954
rect 586302 367398 586538 367634
rect 586622 367398 586858 367634
rect 586302 331718 586538 331954
rect 586622 331718 586858 331954
rect 586302 331398 586538 331634
rect 586622 331398 586858 331634
rect 586302 295718 586538 295954
rect 586622 295718 586858 295954
rect 586302 295398 586538 295634
rect 586622 295398 586858 295634
rect 586302 259718 586538 259954
rect 586622 259718 586858 259954
rect 586302 259398 586538 259634
rect 586622 259398 586858 259634
rect 586302 223718 586538 223954
rect 586622 223718 586858 223954
rect 586302 223398 586538 223634
rect 586622 223398 586858 223634
rect 586302 187718 586538 187954
rect 586622 187718 586858 187954
rect 586302 187398 586538 187634
rect 586622 187398 586858 187634
rect 586302 151718 586538 151954
rect 586622 151718 586858 151954
rect 586302 151398 586538 151634
rect 586622 151398 586858 151634
rect 586302 115718 586538 115954
rect 586622 115718 586858 115954
rect 586302 115398 586538 115634
rect 586622 115398 586858 115634
rect 586302 79718 586538 79954
rect 586622 79718 586858 79954
rect 586302 79398 586538 79634
rect 586622 79398 586858 79634
rect 586302 43718 586538 43954
rect 586622 43718 586858 43954
rect 586302 43398 586538 43634
rect 586622 43398 586858 43634
rect 586302 7718 586538 7954
rect 586622 7718 586858 7954
rect 586302 7398 586538 7634
rect 586622 7398 586858 7634
rect 582326 -1542 582562 -1306
rect 582646 -1542 582882 -1306
rect 582326 -1862 582562 -1626
rect 582646 -1862 582882 -1626
rect 586302 -1542 586538 -1306
rect 586622 -1542 586858 -1306
rect 586302 -1862 586538 -1626
rect 586622 -1862 586858 -1626
rect 587262 696218 587498 696454
rect 587582 696218 587818 696454
rect 587262 695898 587498 696134
rect 587582 695898 587818 696134
rect 587262 660218 587498 660454
rect 587582 660218 587818 660454
rect 587262 659898 587498 660134
rect 587582 659898 587818 660134
rect 587262 624218 587498 624454
rect 587582 624218 587818 624454
rect 587262 623898 587498 624134
rect 587582 623898 587818 624134
rect 587262 588218 587498 588454
rect 587582 588218 587818 588454
rect 587262 587898 587498 588134
rect 587582 587898 587818 588134
rect 587262 552218 587498 552454
rect 587582 552218 587818 552454
rect 587262 551898 587498 552134
rect 587582 551898 587818 552134
rect 587262 516218 587498 516454
rect 587582 516218 587818 516454
rect 587262 515898 587498 516134
rect 587582 515898 587818 516134
rect 587262 480218 587498 480454
rect 587582 480218 587818 480454
rect 587262 479898 587498 480134
rect 587582 479898 587818 480134
rect 587262 444218 587498 444454
rect 587582 444218 587818 444454
rect 587262 443898 587498 444134
rect 587582 443898 587818 444134
rect 587262 408218 587498 408454
rect 587582 408218 587818 408454
rect 587262 407898 587498 408134
rect 587582 407898 587818 408134
rect 587262 372218 587498 372454
rect 587582 372218 587818 372454
rect 587262 371898 587498 372134
rect 587582 371898 587818 372134
rect 587262 336218 587498 336454
rect 587582 336218 587818 336454
rect 587262 335898 587498 336134
rect 587582 335898 587818 336134
rect 587262 300218 587498 300454
rect 587582 300218 587818 300454
rect 587262 299898 587498 300134
rect 587582 299898 587818 300134
rect 587262 264218 587498 264454
rect 587582 264218 587818 264454
rect 587262 263898 587498 264134
rect 587582 263898 587818 264134
rect 587262 228218 587498 228454
rect 587582 228218 587818 228454
rect 587262 227898 587498 228134
rect 587582 227898 587818 228134
rect 587262 192218 587498 192454
rect 587582 192218 587818 192454
rect 587262 191898 587498 192134
rect 587582 191898 587818 192134
rect 587262 156218 587498 156454
rect 587582 156218 587818 156454
rect 587262 155898 587498 156134
rect 587582 155898 587818 156134
rect 587262 120218 587498 120454
rect 587582 120218 587818 120454
rect 587262 119898 587498 120134
rect 587582 119898 587818 120134
rect 587262 84218 587498 84454
rect 587582 84218 587818 84454
rect 587262 83898 587498 84134
rect 587582 83898 587818 84134
rect 587262 48218 587498 48454
rect 587582 48218 587818 48454
rect 587262 47898 587498 48134
rect 587582 47898 587818 48134
rect 587262 12218 587498 12454
rect 587582 12218 587818 12454
rect 587262 11898 587498 12134
rect 587582 11898 587818 12134
rect 587262 -2502 587498 -2266
rect 587582 -2502 587818 -2266
rect 587262 -2822 587498 -2586
rect 587582 -2822 587818 -2586
rect 588222 700718 588458 700954
rect 588542 700718 588778 700954
rect 588222 700398 588458 700634
rect 588542 700398 588778 700634
rect 588222 664718 588458 664954
rect 588542 664718 588778 664954
rect 588222 664398 588458 664634
rect 588542 664398 588778 664634
rect 588222 628718 588458 628954
rect 588542 628718 588778 628954
rect 588222 628398 588458 628634
rect 588542 628398 588778 628634
rect 588222 592718 588458 592954
rect 588542 592718 588778 592954
rect 588222 592398 588458 592634
rect 588542 592398 588778 592634
rect 588222 556718 588458 556954
rect 588542 556718 588778 556954
rect 588222 556398 588458 556634
rect 588542 556398 588778 556634
rect 588222 520718 588458 520954
rect 588542 520718 588778 520954
rect 588222 520398 588458 520634
rect 588542 520398 588778 520634
rect 588222 484718 588458 484954
rect 588542 484718 588778 484954
rect 588222 484398 588458 484634
rect 588542 484398 588778 484634
rect 588222 448718 588458 448954
rect 588542 448718 588778 448954
rect 588222 448398 588458 448634
rect 588542 448398 588778 448634
rect 588222 412718 588458 412954
rect 588542 412718 588778 412954
rect 588222 412398 588458 412634
rect 588542 412398 588778 412634
rect 588222 376718 588458 376954
rect 588542 376718 588778 376954
rect 588222 376398 588458 376634
rect 588542 376398 588778 376634
rect 588222 340718 588458 340954
rect 588542 340718 588778 340954
rect 588222 340398 588458 340634
rect 588542 340398 588778 340634
rect 588222 304718 588458 304954
rect 588542 304718 588778 304954
rect 588222 304398 588458 304634
rect 588542 304398 588778 304634
rect 588222 268718 588458 268954
rect 588542 268718 588778 268954
rect 588222 268398 588458 268634
rect 588542 268398 588778 268634
rect 588222 232718 588458 232954
rect 588542 232718 588778 232954
rect 588222 232398 588458 232634
rect 588542 232398 588778 232634
rect 588222 196718 588458 196954
rect 588542 196718 588778 196954
rect 588222 196398 588458 196634
rect 588542 196398 588778 196634
rect 588222 160718 588458 160954
rect 588542 160718 588778 160954
rect 588222 160398 588458 160634
rect 588542 160398 588778 160634
rect 588222 124718 588458 124954
rect 588542 124718 588778 124954
rect 588222 124398 588458 124634
rect 588542 124398 588778 124634
rect 588222 88718 588458 88954
rect 588542 88718 588778 88954
rect 588222 88398 588458 88634
rect 588542 88398 588778 88634
rect 588222 52718 588458 52954
rect 588542 52718 588778 52954
rect 588222 52398 588458 52634
rect 588542 52398 588778 52634
rect 588222 16718 588458 16954
rect 588542 16718 588778 16954
rect 588222 16398 588458 16634
rect 588542 16398 588778 16634
rect 588222 -3462 588458 -3226
rect 588542 -3462 588778 -3226
rect 588222 -3782 588458 -3546
rect 588542 -3782 588778 -3546
rect 589182 669218 589418 669454
rect 589502 669218 589738 669454
rect 589182 668898 589418 669134
rect 589502 668898 589738 669134
rect 589182 633218 589418 633454
rect 589502 633218 589738 633454
rect 589182 632898 589418 633134
rect 589502 632898 589738 633134
rect 589182 597218 589418 597454
rect 589502 597218 589738 597454
rect 589182 596898 589418 597134
rect 589502 596898 589738 597134
rect 589182 561218 589418 561454
rect 589502 561218 589738 561454
rect 589182 560898 589418 561134
rect 589502 560898 589738 561134
rect 589182 525218 589418 525454
rect 589502 525218 589738 525454
rect 589182 524898 589418 525134
rect 589502 524898 589738 525134
rect 589182 489218 589418 489454
rect 589502 489218 589738 489454
rect 589182 488898 589418 489134
rect 589502 488898 589738 489134
rect 589182 453218 589418 453454
rect 589502 453218 589738 453454
rect 589182 452898 589418 453134
rect 589502 452898 589738 453134
rect 589182 417218 589418 417454
rect 589502 417218 589738 417454
rect 589182 416898 589418 417134
rect 589502 416898 589738 417134
rect 589182 381218 589418 381454
rect 589502 381218 589738 381454
rect 589182 380898 589418 381134
rect 589502 380898 589738 381134
rect 589182 345218 589418 345454
rect 589502 345218 589738 345454
rect 589182 344898 589418 345134
rect 589502 344898 589738 345134
rect 589182 309218 589418 309454
rect 589502 309218 589738 309454
rect 589182 308898 589418 309134
rect 589502 308898 589738 309134
rect 589182 273218 589418 273454
rect 589502 273218 589738 273454
rect 589182 272898 589418 273134
rect 589502 272898 589738 273134
rect 589182 237218 589418 237454
rect 589502 237218 589738 237454
rect 589182 236898 589418 237134
rect 589502 236898 589738 237134
rect 589182 201218 589418 201454
rect 589502 201218 589738 201454
rect 589182 200898 589418 201134
rect 589502 200898 589738 201134
rect 589182 165218 589418 165454
rect 589502 165218 589738 165454
rect 589182 164898 589418 165134
rect 589502 164898 589738 165134
rect 589182 129218 589418 129454
rect 589502 129218 589738 129454
rect 589182 128898 589418 129134
rect 589502 128898 589738 129134
rect 589182 93218 589418 93454
rect 589502 93218 589738 93454
rect 589182 92898 589418 93134
rect 589502 92898 589738 93134
rect 589182 57218 589418 57454
rect 589502 57218 589738 57454
rect 589182 56898 589418 57134
rect 589502 56898 589738 57134
rect 589182 21218 589418 21454
rect 589502 21218 589738 21454
rect 589182 20898 589418 21134
rect 589502 20898 589738 21134
rect 589182 -4422 589418 -4186
rect 589502 -4422 589738 -4186
rect 589182 -4742 589418 -4506
rect 589502 -4742 589738 -4506
rect 590142 673718 590378 673954
rect 590462 673718 590698 673954
rect 590142 673398 590378 673634
rect 590462 673398 590698 673634
rect 590142 637718 590378 637954
rect 590462 637718 590698 637954
rect 590142 637398 590378 637634
rect 590462 637398 590698 637634
rect 590142 601718 590378 601954
rect 590462 601718 590698 601954
rect 590142 601398 590378 601634
rect 590462 601398 590698 601634
rect 590142 565718 590378 565954
rect 590462 565718 590698 565954
rect 590142 565398 590378 565634
rect 590462 565398 590698 565634
rect 590142 529718 590378 529954
rect 590462 529718 590698 529954
rect 590142 529398 590378 529634
rect 590462 529398 590698 529634
rect 590142 493718 590378 493954
rect 590462 493718 590698 493954
rect 590142 493398 590378 493634
rect 590462 493398 590698 493634
rect 590142 457718 590378 457954
rect 590462 457718 590698 457954
rect 590142 457398 590378 457634
rect 590462 457398 590698 457634
rect 590142 421718 590378 421954
rect 590462 421718 590698 421954
rect 590142 421398 590378 421634
rect 590462 421398 590698 421634
rect 590142 385718 590378 385954
rect 590462 385718 590698 385954
rect 590142 385398 590378 385634
rect 590462 385398 590698 385634
rect 590142 349718 590378 349954
rect 590462 349718 590698 349954
rect 590142 349398 590378 349634
rect 590462 349398 590698 349634
rect 590142 313718 590378 313954
rect 590462 313718 590698 313954
rect 590142 313398 590378 313634
rect 590462 313398 590698 313634
rect 590142 277718 590378 277954
rect 590462 277718 590698 277954
rect 590142 277398 590378 277634
rect 590462 277398 590698 277634
rect 590142 241718 590378 241954
rect 590462 241718 590698 241954
rect 590142 241398 590378 241634
rect 590462 241398 590698 241634
rect 590142 205718 590378 205954
rect 590462 205718 590698 205954
rect 590142 205398 590378 205634
rect 590462 205398 590698 205634
rect 590142 169718 590378 169954
rect 590462 169718 590698 169954
rect 590142 169398 590378 169634
rect 590462 169398 590698 169634
rect 590142 133718 590378 133954
rect 590462 133718 590698 133954
rect 590142 133398 590378 133634
rect 590462 133398 590698 133634
rect 590142 97718 590378 97954
rect 590462 97718 590698 97954
rect 590142 97398 590378 97634
rect 590462 97398 590698 97634
rect 590142 61718 590378 61954
rect 590462 61718 590698 61954
rect 590142 61398 590378 61634
rect 590462 61398 590698 61634
rect 590142 25718 590378 25954
rect 590462 25718 590698 25954
rect 590142 25398 590378 25634
rect 590462 25398 590698 25634
rect 590142 -5382 590378 -5146
rect 590462 -5382 590698 -5146
rect 590142 -5702 590378 -5466
rect 590462 -5702 590698 -5466
rect 591102 678218 591338 678454
rect 591422 678218 591658 678454
rect 591102 677898 591338 678134
rect 591422 677898 591658 678134
rect 591102 642218 591338 642454
rect 591422 642218 591658 642454
rect 591102 641898 591338 642134
rect 591422 641898 591658 642134
rect 591102 606218 591338 606454
rect 591422 606218 591658 606454
rect 591102 605898 591338 606134
rect 591422 605898 591658 606134
rect 591102 570218 591338 570454
rect 591422 570218 591658 570454
rect 591102 569898 591338 570134
rect 591422 569898 591658 570134
rect 591102 534218 591338 534454
rect 591422 534218 591658 534454
rect 591102 533898 591338 534134
rect 591422 533898 591658 534134
rect 591102 498218 591338 498454
rect 591422 498218 591658 498454
rect 591102 497898 591338 498134
rect 591422 497898 591658 498134
rect 591102 462218 591338 462454
rect 591422 462218 591658 462454
rect 591102 461898 591338 462134
rect 591422 461898 591658 462134
rect 591102 426218 591338 426454
rect 591422 426218 591658 426454
rect 591102 425898 591338 426134
rect 591422 425898 591658 426134
rect 591102 390218 591338 390454
rect 591422 390218 591658 390454
rect 591102 389898 591338 390134
rect 591422 389898 591658 390134
rect 591102 354218 591338 354454
rect 591422 354218 591658 354454
rect 591102 353898 591338 354134
rect 591422 353898 591658 354134
rect 591102 318218 591338 318454
rect 591422 318218 591658 318454
rect 591102 317898 591338 318134
rect 591422 317898 591658 318134
rect 591102 282218 591338 282454
rect 591422 282218 591658 282454
rect 591102 281898 591338 282134
rect 591422 281898 591658 282134
rect 591102 246218 591338 246454
rect 591422 246218 591658 246454
rect 591102 245898 591338 246134
rect 591422 245898 591658 246134
rect 591102 210218 591338 210454
rect 591422 210218 591658 210454
rect 591102 209898 591338 210134
rect 591422 209898 591658 210134
rect 591102 174218 591338 174454
rect 591422 174218 591658 174454
rect 591102 173898 591338 174134
rect 591422 173898 591658 174134
rect 591102 138218 591338 138454
rect 591422 138218 591658 138454
rect 591102 137898 591338 138134
rect 591422 137898 591658 138134
rect 591102 102218 591338 102454
rect 591422 102218 591658 102454
rect 591102 101898 591338 102134
rect 591422 101898 591658 102134
rect 591102 66218 591338 66454
rect 591422 66218 591658 66454
rect 591102 65898 591338 66134
rect 591422 65898 591658 66134
rect 591102 30218 591338 30454
rect 591422 30218 591658 30454
rect 591102 29898 591338 30134
rect 591422 29898 591658 30134
rect 591102 -6342 591338 -6106
rect 591422 -6342 591658 -6106
rect 591102 -6662 591338 -6426
rect 591422 -6662 591658 -6426
rect 592062 682718 592298 682954
rect 592382 682718 592618 682954
rect 592062 682398 592298 682634
rect 592382 682398 592618 682634
rect 592062 646718 592298 646954
rect 592382 646718 592618 646954
rect 592062 646398 592298 646634
rect 592382 646398 592618 646634
rect 592062 610718 592298 610954
rect 592382 610718 592618 610954
rect 592062 610398 592298 610634
rect 592382 610398 592618 610634
rect 592062 574718 592298 574954
rect 592382 574718 592618 574954
rect 592062 574398 592298 574634
rect 592382 574398 592618 574634
rect 592062 538718 592298 538954
rect 592382 538718 592618 538954
rect 592062 538398 592298 538634
rect 592382 538398 592618 538634
rect 592062 502718 592298 502954
rect 592382 502718 592618 502954
rect 592062 502398 592298 502634
rect 592382 502398 592618 502634
rect 592062 466718 592298 466954
rect 592382 466718 592618 466954
rect 592062 466398 592298 466634
rect 592382 466398 592618 466634
rect 592062 430718 592298 430954
rect 592382 430718 592618 430954
rect 592062 430398 592298 430634
rect 592382 430398 592618 430634
rect 592062 394718 592298 394954
rect 592382 394718 592618 394954
rect 592062 394398 592298 394634
rect 592382 394398 592618 394634
rect 592062 358718 592298 358954
rect 592382 358718 592618 358954
rect 592062 358398 592298 358634
rect 592382 358398 592618 358634
rect 592062 322718 592298 322954
rect 592382 322718 592618 322954
rect 592062 322398 592298 322634
rect 592382 322398 592618 322634
rect 592062 286718 592298 286954
rect 592382 286718 592618 286954
rect 592062 286398 592298 286634
rect 592382 286398 592618 286634
rect 592062 250718 592298 250954
rect 592382 250718 592618 250954
rect 592062 250398 592298 250634
rect 592382 250398 592618 250634
rect 592062 214718 592298 214954
rect 592382 214718 592618 214954
rect 592062 214398 592298 214634
rect 592382 214398 592618 214634
rect 592062 178718 592298 178954
rect 592382 178718 592618 178954
rect 592062 178398 592298 178634
rect 592382 178398 592618 178634
rect 592062 142718 592298 142954
rect 592382 142718 592618 142954
rect 592062 142398 592298 142634
rect 592382 142398 592618 142634
rect 592062 106718 592298 106954
rect 592382 106718 592618 106954
rect 592062 106398 592298 106634
rect 592382 106398 592618 106634
rect 592062 70718 592298 70954
rect 592382 70718 592618 70954
rect 592062 70398 592298 70634
rect 592382 70398 592618 70634
rect 592062 34718 592298 34954
rect 592382 34718 592618 34954
rect 592062 34398 592298 34634
rect 592382 34398 592618 34634
rect 592062 -7302 592298 -7066
rect 592382 -7302 592618 -7066
rect 592062 -7622 592298 -7386
rect 592382 -7622 592618 -7386
<< metal5 >>
rect -8726 711558 592650 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 33326 711558
rect 33562 711322 33646 711558
rect 33882 711322 69326 711558
rect 69562 711322 69646 711558
rect 69882 711322 105326 711558
rect 105562 711322 105646 711558
rect 105882 711322 141326 711558
rect 141562 711322 141646 711558
rect 141882 711322 177326 711558
rect 177562 711322 177646 711558
rect 177882 711322 213326 711558
rect 213562 711322 213646 711558
rect 213882 711322 249326 711558
rect 249562 711322 249646 711558
rect 249882 711322 285326 711558
rect 285562 711322 285646 711558
rect 285882 711322 321326 711558
rect 321562 711322 321646 711558
rect 321882 711322 357326 711558
rect 357562 711322 357646 711558
rect 357882 711322 393326 711558
rect 393562 711322 393646 711558
rect 393882 711322 429326 711558
rect 429562 711322 429646 711558
rect 429882 711322 465326 711558
rect 465562 711322 465646 711558
rect 465882 711322 501326 711558
rect 501562 711322 501646 711558
rect 501882 711322 537326 711558
rect 537562 711322 537646 711558
rect 537882 711322 573326 711558
rect 573562 711322 573646 711558
rect 573882 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect -8726 711238 592650 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 33326 711238
rect 33562 711002 33646 711238
rect 33882 711002 69326 711238
rect 69562 711002 69646 711238
rect 69882 711002 105326 711238
rect 105562 711002 105646 711238
rect 105882 711002 141326 711238
rect 141562 711002 141646 711238
rect 141882 711002 177326 711238
rect 177562 711002 177646 711238
rect 177882 711002 213326 711238
rect 213562 711002 213646 711238
rect 213882 711002 249326 711238
rect 249562 711002 249646 711238
rect 249882 711002 285326 711238
rect 285562 711002 285646 711238
rect 285882 711002 321326 711238
rect 321562 711002 321646 711238
rect 321882 711002 357326 711238
rect 357562 711002 357646 711238
rect 357882 711002 393326 711238
rect 393562 711002 393646 711238
rect 393882 711002 429326 711238
rect 429562 711002 429646 711238
rect 429882 711002 465326 711238
rect 465562 711002 465646 711238
rect 465882 711002 501326 711238
rect 501562 711002 501646 711238
rect 501882 711002 537326 711238
rect 537562 711002 537646 711238
rect 537882 711002 573326 711238
rect 573562 711002 573646 711238
rect 573882 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect -8726 710970 592650 711002
rect -7766 710598 591690 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 28826 710598
rect 29062 710362 29146 710598
rect 29382 710362 64826 710598
rect 65062 710362 65146 710598
rect 65382 710362 100826 710598
rect 101062 710362 101146 710598
rect 101382 710362 136826 710598
rect 137062 710362 137146 710598
rect 137382 710362 172826 710598
rect 173062 710362 173146 710598
rect 173382 710362 208826 710598
rect 209062 710362 209146 710598
rect 209382 710362 244826 710598
rect 245062 710362 245146 710598
rect 245382 710362 280826 710598
rect 281062 710362 281146 710598
rect 281382 710362 316826 710598
rect 317062 710362 317146 710598
rect 317382 710362 352826 710598
rect 353062 710362 353146 710598
rect 353382 710362 388826 710598
rect 389062 710362 389146 710598
rect 389382 710362 424826 710598
rect 425062 710362 425146 710598
rect 425382 710362 460826 710598
rect 461062 710362 461146 710598
rect 461382 710362 496826 710598
rect 497062 710362 497146 710598
rect 497382 710362 532826 710598
rect 533062 710362 533146 710598
rect 533382 710362 568826 710598
rect 569062 710362 569146 710598
rect 569382 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect -7766 710278 591690 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 28826 710278
rect 29062 710042 29146 710278
rect 29382 710042 64826 710278
rect 65062 710042 65146 710278
rect 65382 710042 100826 710278
rect 101062 710042 101146 710278
rect 101382 710042 136826 710278
rect 137062 710042 137146 710278
rect 137382 710042 172826 710278
rect 173062 710042 173146 710278
rect 173382 710042 208826 710278
rect 209062 710042 209146 710278
rect 209382 710042 244826 710278
rect 245062 710042 245146 710278
rect 245382 710042 280826 710278
rect 281062 710042 281146 710278
rect 281382 710042 316826 710278
rect 317062 710042 317146 710278
rect 317382 710042 352826 710278
rect 353062 710042 353146 710278
rect 353382 710042 388826 710278
rect 389062 710042 389146 710278
rect 389382 710042 424826 710278
rect 425062 710042 425146 710278
rect 425382 710042 460826 710278
rect 461062 710042 461146 710278
rect 461382 710042 496826 710278
rect 497062 710042 497146 710278
rect 497382 710042 532826 710278
rect 533062 710042 533146 710278
rect 533382 710042 568826 710278
rect 569062 710042 569146 710278
rect 569382 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect -7766 710010 591690 710042
rect -6806 709638 590730 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 24326 709638
rect 24562 709402 24646 709638
rect 24882 709402 60326 709638
rect 60562 709402 60646 709638
rect 60882 709402 96326 709638
rect 96562 709402 96646 709638
rect 96882 709402 132326 709638
rect 132562 709402 132646 709638
rect 132882 709402 168326 709638
rect 168562 709402 168646 709638
rect 168882 709402 204326 709638
rect 204562 709402 204646 709638
rect 204882 709402 240326 709638
rect 240562 709402 240646 709638
rect 240882 709402 276326 709638
rect 276562 709402 276646 709638
rect 276882 709402 312326 709638
rect 312562 709402 312646 709638
rect 312882 709402 348326 709638
rect 348562 709402 348646 709638
rect 348882 709402 384326 709638
rect 384562 709402 384646 709638
rect 384882 709402 420326 709638
rect 420562 709402 420646 709638
rect 420882 709402 456326 709638
rect 456562 709402 456646 709638
rect 456882 709402 492326 709638
rect 492562 709402 492646 709638
rect 492882 709402 528326 709638
rect 528562 709402 528646 709638
rect 528882 709402 564326 709638
rect 564562 709402 564646 709638
rect 564882 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect -6806 709318 590730 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 24326 709318
rect 24562 709082 24646 709318
rect 24882 709082 60326 709318
rect 60562 709082 60646 709318
rect 60882 709082 96326 709318
rect 96562 709082 96646 709318
rect 96882 709082 132326 709318
rect 132562 709082 132646 709318
rect 132882 709082 168326 709318
rect 168562 709082 168646 709318
rect 168882 709082 204326 709318
rect 204562 709082 204646 709318
rect 204882 709082 240326 709318
rect 240562 709082 240646 709318
rect 240882 709082 276326 709318
rect 276562 709082 276646 709318
rect 276882 709082 312326 709318
rect 312562 709082 312646 709318
rect 312882 709082 348326 709318
rect 348562 709082 348646 709318
rect 348882 709082 384326 709318
rect 384562 709082 384646 709318
rect 384882 709082 420326 709318
rect 420562 709082 420646 709318
rect 420882 709082 456326 709318
rect 456562 709082 456646 709318
rect 456882 709082 492326 709318
rect 492562 709082 492646 709318
rect 492882 709082 528326 709318
rect 528562 709082 528646 709318
rect 528882 709082 564326 709318
rect 564562 709082 564646 709318
rect 564882 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect -6806 709050 590730 709082
rect -5846 708678 589770 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 19826 708678
rect 20062 708442 20146 708678
rect 20382 708442 55826 708678
rect 56062 708442 56146 708678
rect 56382 708442 91826 708678
rect 92062 708442 92146 708678
rect 92382 708442 127826 708678
rect 128062 708442 128146 708678
rect 128382 708442 163826 708678
rect 164062 708442 164146 708678
rect 164382 708442 199826 708678
rect 200062 708442 200146 708678
rect 200382 708442 235826 708678
rect 236062 708442 236146 708678
rect 236382 708442 271826 708678
rect 272062 708442 272146 708678
rect 272382 708442 307826 708678
rect 308062 708442 308146 708678
rect 308382 708442 343826 708678
rect 344062 708442 344146 708678
rect 344382 708442 379826 708678
rect 380062 708442 380146 708678
rect 380382 708442 415826 708678
rect 416062 708442 416146 708678
rect 416382 708442 451826 708678
rect 452062 708442 452146 708678
rect 452382 708442 487826 708678
rect 488062 708442 488146 708678
rect 488382 708442 523826 708678
rect 524062 708442 524146 708678
rect 524382 708442 559826 708678
rect 560062 708442 560146 708678
rect 560382 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect -5846 708358 589770 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 19826 708358
rect 20062 708122 20146 708358
rect 20382 708122 55826 708358
rect 56062 708122 56146 708358
rect 56382 708122 91826 708358
rect 92062 708122 92146 708358
rect 92382 708122 127826 708358
rect 128062 708122 128146 708358
rect 128382 708122 163826 708358
rect 164062 708122 164146 708358
rect 164382 708122 199826 708358
rect 200062 708122 200146 708358
rect 200382 708122 235826 708358
rect 236062 708122 236146 708358
rect 236382 708122 271826 708358
rect 272062 708122 272146 708358
rect 272382 708122 307826 708358
rect 308062 708122 308146 708358
rect 308382 708122 343826 708358
rect 344062 708122 344146 708358
rect 344382 708122 379826 708358
rect 380062 708122 380146 708358
rect 380382 708122 415826 708358
rect 416062 708122 416146 708358
rect 416382 708122 451826 708358
rect 452062 708122 452146 708358
rect 452382 708122 487826 708358
rect 488062 708122 488146 708358
rect 488382 708122 523826 708358
rect 524062 708122 524146 708358
rect 524382 708122 559826 708358
rect 560062 708122 560146 708358
rect 560382 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect -5846 708090 589770 708122
rect -4886 707718 588810 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 15326 707718
rect 15562 707482 15646 707718
rect 15882 707482 51326 707718
rect 51562 707482 51646 707718
rect 51882 707482 87326 707718
rect 87562 707482 87646 707718
rect 87882 707482 123326 707718
rect 123562 707482 123646 707718
rect 123882 707482 159326 707718
rect 159562 707482 159646 707718
rect 159882 707482 195326 707718
rect 195562 707482 195646 707718
rect 195882 707482 231326 707718
rect 231562 707482 231646 707718
rect 231882 707482 267326 707718
rect 267562 707482 267646 707718
rect 267882 707482 303326 707718
rect 303562 707482 303646 707718
rect 303882 707482 339326 707718
rect 339562 707482 339646 707718
rect 339882 707482 375326 707718
rect 375562 707482 375646 707718
rect 375882 707482 411326 707718
rect 411562 707482 411646 707718
rect 411882 707482 447326 707718
rect 447562 707482 447646 707718
rect 447882 707482 483326 707718
rect 483562 707482 483646 707718
rect 483882 707482 519326 707718
rect 519562 707482 519646 707718
rect 519882 707482 555326 707718
rect 555562 707482 555646 707718
rect 555882 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect -4886 707398 588810 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 15326 707398
rect 15562 707162 15646 707398
rect 15882 707162 51326 707398
rect 51562 707162 51646 707398
rect 51882 707162 87326 707398
rect 87562 707162 87646 707398
rect 87882 707162 123326 707398
rect 123562 707162 123646 707398
rect 123882 707162 159326 707398
rect 159562 707162 159646 707398
rect 159882 707162 195326 707398
rect 195562 707162 195646 707398
rect 195882 707162 231326 707398
rect 231562 707162 231646 707398
rect 231882 707162 267326 707398
rect 267562 707162 267646 707398
rect 267882 707162 303326 707398
rect 303562 707162 303646 707398
rect 303882 707162 339326 707398
rect 339562 707162 339646 707398
rect 339882 707162 375326 707398
rect 375562 707162 375646 707398
rect 375882 707162 411326 707398
rect 411562 707162 411646 707398
rect 411882 707162 447326 707398
rect 447562 707162 447646 707398
rect 447882 707162 483326 707398
rect 483562 707162 483646 707398
rect 483882 707162 519326 707398
rect 519562 707162 519646 707398
rect 519882 707162 555326 707398
rect 555562 707162 555646 707398
rect 555882 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect -4886 707130 588810 707162
rect -3926 706758 587850 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 10826 706758
rect 11062 706522 11146 706758
rect 11382 706522 46826 706758
rect 47062 706522 47146 706758
rect 47382 706522 82826 706758
rect 83062 706522 83146 706758
rect 83382 706522 118826 706758
rect 119062 706522 119146 706758
rect 119382 706522 154826 706758
rect 155062 706522 155146 706758
rect 155382 706522 190826 706758
rect 191062 706522 191146 706758
rect 191382 706522 226826 706758
rect 227062 706522 227146 706758
rect 227382 706522 262826 706758
rect 263062 706522 263146 706758
rect 263382 706522 298826 706758
rect 299062 706522 299146 706758
rect 299382 706522 334826 706758
rect 335062 706522 335146 706758
rect 335382 706522 370826 706758
rect 371062 706522 371146 706758
rect 371382 706522 406826 706758
rect 407062 706522 407146 706758
rect 407382 706522 442826 706758
rect 443062 706522 443146 706758
rect 443382 706522 478826 706758
rect 479062 706522 479146 706758
rect 479382 706522 514826 706758
rect 515062 706522 515146 706758
rect 515382 706522 550826 706758
rect 551062 706522 551146 706758
rect 551382 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect -3926 706438 587850 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 10826 706438
rect 11062 706202 11146 706438
rect 11382 706202 46826 706438
rect 47062 706202 47146 706438
rect 47382 706202 82826 706438
rect 83062 706202 83146 706438
rect 83382 706202 118826 706438
rect 119062 706202 119146 706438
rect 119382 706202 154826 706438
rect 155062 706202 155146 706438
rect 155382 706202 190826 706438
rect 191062 706202 191146 706438
rect 191382 706202 226826 706438
rect 227062 706202 227146 706438
rect 227382 706202 262826 706438
rect 263062 706202 263146 706438
rect 263382 706202 298826 706438
rect 299062 706202 299146 706438
rect 299382 706202 334826 706438
rect 335062 706202 335146 706438
rect 335382 706202 370826 706438
rect 371062 706202 371146 706438
rect 371382 706202 406826 706438
rect 407062 706202 407146 706438
rect 407382 706202 442826 706438
rect 443062 706202 443146 706438
rect 443382 706202 478826 706438
rect 479062 706202 479146 706438
rect 479382 706202 514826 706438
rect 515062 706202 515146 706438
rect 515382 706202 550826 706438
rect 551062 706202 551146 706438
rect 551382 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect -3926 706170 587850 706202
rect -2966 705798 586890 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 6326 705798
rect 6562 705562 6646 705798
rect 6882 705562 42326 705798
rect 42562 705562 42646 705798
rect 42882 705562 78326 705798
rect 78562 705562 78646 705798
rect 78882 705562 114326 705798
rect 114562 705562 114646 705798
rect 114882 705562 150326 705798
rect 150562 705562 150646 705798
rect 150882 705562 186326 705798
rect 186562 705562 186646 705798
rect 186882 705562 222326 705798
rect 222562 705562 222646 705798
rect 222882 705562 258326 705798
rect 258562 705562 258646 705798
rect 258882 705562 294326 705798
rect 294562 705562 294646 705798
rect 294882 705562 330326 705798
rect 330562 705562 330646 705798
rect 330882 705562 366326 705798
rect 366562 705562 366646 705798
rect 366882 705562 402326 705798
rect 402562 705562 402646 705798
rect 402882 705562 438326 705798
rect 438562 705562 438646 705798
rect 438882 705562 474326 705798
rect 474562 705562 474646 705798
rect 474882 705562 510326 705798
rect 510562 705562 510646 705798
rect 510882 705562 546326 705798
rect 546562 705562 546646 705798
rect 546882 705562 582326 705798
rect 582562 705562 582646 705798
rect 582882 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect -2966 705478 586890 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 6326 705478
rect 6562 705242 6646 705478
rect 6882 705242 42326 705478
rect 42562 705242 42646 705478
rect 42882 705242 78326 705478
rect 78562 705242 78646 705478
rect 78882 705242 114326 705478
rect 114562 705242 114646 705478
rect 114882 705242 150326 705478
rect 150562 705242 150646 705478
rect 150882 705242 186326 705478
rect 186562 705242 186646 705478
rect 186882 705242 222326 705478
rect 222562 705242 222646 705478
rect 222882 705242 258326 705478
rect 258562 705242 258646 705478
rect 258882 705242 294326 705478
rect 294562 705242 294646 705478
rect 294882 705242 330326 705478
rect 330562 705242 330646 705478
rect 330882 705242 366326 705478
rect 366562 705242 366646 705478
rect 366882 705242 402326 705478
rect 402562 705242 402646 705478
rect 402882 705242 438326 705478
rect 438562 705242 438646 705478
rect 438882 705242 474326 705478
rect 474562 705242 474646 705478
rect 474882 705242 510326 705478
rect 510562 705242 510646 705478
rect 510882 705242 546326 705478
rect 546562 705242 546646 705478
rect 546882 705242 582326 705478
rect 582562 705242 582646 705478
rect 582882 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect -2966 705210 586890 705242
rect -2006 704838 585930 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect -2006 704518 585930 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect -2006 704250 585930 704282
rect -8726 700954 592650 700986
rect -8726 700718 -4854 700954
rect -4618 700718 -4534 700954
rect -4298 700718 15326 700954
rect 15562 700718 15646 700954
rect 15882 700718 51326 700954
rect 51562 700718 51646 700954
rect 51882 700718 87326 700954
rect 87562 700718 87646 700954
rect 87882 700718 123326 700954
rect 123562 700718 123646 700954
rect 123882 700718 159326 700954
rect 159562 700718 159646 700954
rect 159882 700718 195326 700954
rect 195562 700718 195646 700954
rect 195882 700718 231326 700954
rect 231562 700718 231646 700954
rect 231882 700718 267326 700954
rect 267562 700718 267646 700954
rect 267882 700718 303326 700954
rect 303562 700718 303646 700954
rect 303882 700718 339326 700954
rect 339562 700718 339646 700954
rect 339882 700718 375326 700954
rect 375562 700718 375646 700954
rect 375882 700718 411326 700954
rect 411562 700718 411646 700954
rect 411882 700718 447326 700954
rect 447562 700718 447646 700954
rect 447882 700718 483326 700954
rect 483562 700718 483646 700954
rect 483882 700718 519326 700954
rect 519562 700718 519646 700954
rect 519882 700718 555326 700954
rect 555562 700718 555646 700954
rect 555882 700718 588222 700954
rect 588458 700718 588542 700954
rect 588778 700718 592650 700954
rect -8726 700634 592650 700718
rect -8726 700398 -4854 700634
rect -4618 700398 -4534 700634
rect -4298 700398 15326 700634
rect 15562 700398 15646 700634
rect 15882 700398 51326 700634
rect 51562 700398 51646 700634
rect 51882 700398 87326 700634
rect 87562 700398 87646 700634
rect 87882 700398 123326 700634
rect 123562 700398 123646 700634
rect 123882 700398 159326 700634
rect 159562 700398 159646 700634
rect 159882 700398 195326 700634
rect 195562 700398 195646 700634
rect 195882 700398 231326 700634
rect 231562 700398 231646 700634
rect 231882 700398 267326 700634
rect 267562 700398 267646 700634
rect 267882 700398 303326 700634
rect 303562 700398 303646 700634
rect 303882 700398 339326 700634
rect 339562 700398 339646 700634
rect 339882 700398 375326 700634
rect 375562 700398 375646 700634
rect 375882 700398 411326 700634
rect 411562 700398 411646 700634
rect 411882 700398 447326 700634
rect 447562 700398 447646 700634
rect 447882 700398 483326 700634
rect 483562 700398 483646 700634
rect 483882 700398 519326 700634
rect 519562 700398 519646 700634
rect 519882 700398 555326 700634
rect 555562 700398 555646 700634
rect 555882 700398 588222 700634
rect 588458 700398 588542 700634
rect 588778 700398 592650 700634
rect -8726 700366 592650 700398
rect -8726 696454 592650 696486
rect -8726 696218 -3894 696454
rect -3658 696218 -3574 696454
rect -3338 696218 10826 696454
rect 11062 696218 11146 696454
rect 11382 696218 46826 696454
rect 47062 696218 47146 696454
rect 47382 696218 82826 696454
rect 83062 696218 83146 696454
rect 83382 696218 118826 696454
rect 119062 696218 119146 696454
rect 119382 696218 154826 696454
rect 155062 696218 155146 696454
rect 155382 696218 190826 696454
rect 191062 696218 191146 696454
rect 191382 696218 226826 696454
rect 227062 696218 227146 696454
rect 227382 696218 262826 696454
rect 263062 696218 263146 696454
rect 263382 696218 298826 696454
rect 299062 696218 299146 696454
rect 299382 696218 334826 696454
rect 335062 696218 335146 696454
rect 335382 696218 370826 696454
rect 371062 696218 371146 696454
rect 371382 696218 406826 696454
rect 407062 696218 407146 696454
rect 407382 696218 442826 696454
rect 443062 696218 443146 696454
rect 443382 696218 478826 696454
rect 479062 696218 479146 696454
rect 479382 696218 514826 696454
rect 515062 696218 515146 696454
rect 515382 696218 550826 696454
rect 551062 696218 551146 696454
rect 551382 696218 587262 696454
rect 587498 696218 587582 696454
rect 587818 696218 592650 696454
rect -8726 696134 592650 696218
rect -8726 695898 -3894 696134
rect -3658 695898 -3574 696134
rect -3338 695898 10826 696134
rect 11062 695898 11146 696134
rect 11382 695898 46826 696134
rect 47062 695898 47146 696134
rect 47382 695898 82826 696134
rect 83062 695898 83146 696134
rect 83382 695898 118826 696134
rect 119062 695898 119146 696134
rect 119382 695898 154826 696134
rect 155062 695898 155146 696134
rect 155382 695898 190826 696134
rect 191062 695898 191146 696134
rect 191382 695898 226826 696134
rect 227062 695898 227146 696134
rect 227382 695898 262826 696134
rect 263062 695898 263146 696134
rect 263382 695898 298826 696134
rect 299062 695898 299146 696134
rect 299382 695898 334826 696134
rect 335062 695898 335146 696134
rect 335382 695898 370826 696134
rect 371062 695898 371146 696134
rect 371382 695898 406826 696134
rect 407062 695898 407146 696134
rect 407382 695898 442826 696134
rect 443062 695898 443146 696134
rect 443382 695898 478826 696134
rect 479062 695898 479146 696134
rect 479382 695898 514826 696134
rect 515062 695898 515146 696134
rect 515382 695898 550826 696134
rect 551062 695898 551146 696134
rect 551382 695898 587262 696134
rect 587498 695898 587582 696134
rect 587818 695898 592650 696134
rect -8726 695866 592650 695898
rect -8726 691954 592650 691986
rect -8726 691718 -2934 691954
rect -2698 691718 -2614 691954
rect -2378 691718 6326 691954
rect 6562 691718 6646 691954
rect 6882 691718 42326 691954
rect 42562 691718 42646 691954
rect 42882 691718 78326 691954
rect 78562 691718 78646 691954
rect 78882 691718 114326 691954
rect 114562 691718 114646 691954
rect 114882 691718 150326 691954
rect 150562 691718 150646 691954
rect 150882 691718 186326 691954
rect 186562 691718 186646 691954
rect 186882 691718 222326 691954
rect 222562 691718 222646 691954
rect 222882 691718 258326 691954
rect 258562 691718 258646 691954
rect 258882 691718 294326 691954
rect 294562 691718 294646 691954
rect 294882 691718 330326 691954
rect 330562 691718 330646 691954
rect 330882 691718 366326 691954
rect 366562 691718 366646 691954
rect 366882 691718 402326 691954
rect 402562 691718 402646 691954
rect 402882 691718 438326 691954
rect 438562 691718 438646 691954
rect 438882 691718 474326 691954
rect 474562 691718 474646 691954
rect 474882 691718 510326 691954
rect 510562 691718 510646 691954
rect 510882 691718 546326 691954
rect 546562 691718 546646 691954
rect 546882 691718 582326 691954
rect 582562 691718 582646 691954
rect 582882 691718 586302 691954
rect 586538 691718 586622 691954
rect 586858 691718 592650 691954
rect -8726 691634 592650 691718
rect -8726 691398 -2934 691634
rect -2698 691398 -2614 691634
rect -2378 691398 6326 691634
rect 6562 691398 6646 691634
rect 6882 691398 42326 691634
rect 42562 691398 42646 691634
rect 42882 691398 78326 691634
rect 78562 691398 78646 691634
rect 78882 691398 114326 691634
rect 114562 691398 114646 691634
rect 114882 691398 150326 691634
rect 150562 691398 150646 691634
rect 150882 691398 186326 691634
rect 186562 691398 186646 691634
rect 186882 691398 222326 691634
rect 222562 691398 222646 691634
rect 222882 691398 258326 691634
rect 258562 691398 258646 691634
rect 258882 691398 294326 691634
rect 294562 691398 294646 691634
rect 294882 691398 330326 691634
rect 330562 691398 330646 691634
rect 330882 691398 366326 691634
rect 366562 691398 366646 691634
rect 366882 691398 402326 691634
rect 402562 691398 402646 691634
rect 402882 691398 438326 691634
rect 438562 691398 438646 691634
rect 438882 691398 474326 691634
rect 474562 691398 474646 691634
rect 474882 691398 510326 691634
rect 510562 691398 510646 691634
rect 510882 691398 546326 691634
rect 546562 691398 546646 691634
rect 546882 691398 582326 691634
rect 582562 691398 582646 691634
rect 582882 691398 586302 691634
rect 586538 691398 586622 691634
rect 586858 691398 592650 691634
rect -8726 691366 592650 691398
rect -8726 687454 592650 687486
rect -8726 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 592650 687454
rect -8726 687134 592650 687218
rect -8726 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 592650 687134
rect -8726 686866 592650 686898
rect -8726 682954 592650 682986
rect -8726 682718 -8694 682954
rect -8458 682718 -8374 682954
rect -8138 682718 33326 682954
rect 33562 682718 33646 682954
rect 33882 682718 69326 682954
rect 69562 682718 69646 682954
rect 69882 682718 105326 682954
rect 105562 682718 105646 682954
rect 105882 682718 141326 682954
rect 141562 682718 141646 682954
rect 141882 682718 177326 682954
rect 177562 682718 177646 682954
rect 177882 682718 213326 682954
rect 213562 682718 213646 682954
rect 213882 682718 249326 682954
rect 249562 682718 249646 682954
rect 249882 682718 285326 682954
rect 285562 682718 285646 682954
rect 285882 682718 321326 682954
rect 321562 682718 321646 682954
rect 321882 682718 357326 682954
rect 357562 682718 357646 682954
rect 357882 682718 393326 682954
rect 393562 682718 393646 682954
rect 393882 682718 429326 682954
rect 429562 682718 429646 682954
rect 429882 682718 465326 682954
rect 465562 682718 465646 682954
rect 465882 682718 501326 682954
rect 501562 682718 501646 682954
rect 501882 682718 537326 682954
rect 537562 682718 537646 682954
rect 537882 682718 573326 682954
rect 573562 682718 573646 682954
rect 573882 682718 592062 682954
rect 592298 682718 592382 682954
rect 592618 682718 592650 682954
rect -8726 682634 592650 682718
rect -8726 682398 -8694 682634
rect -8458 682398 -8374 682634
rect -8138 682398 33326 682634
rect 33562 682398 33646 682634
rect 33882 682398 69326 682634
rect 69562 682398 69646 682634
rect 69882 682398 105326 682634
rect 105562 682398 105646 682634
rect 105882 682398 141326 682634
rect 141562 682398 141646 682634
rect 141882 682398 177326 682634
rect 177562 682398 177646 682634
rect 177882 682398 213326 682634
rect 213562 682398 213646 682634
rect 213882 682398 249326 682634
rect 249562 682398 249646 682634
rect 249882 682398 285326 682634
rect 285562 682398 285646 682634
rect 285882 682398 321326 682634
rect 321562 682398 321646 682634
rect 321882 682398 357326 682634
rect 357562 682398 357646 682634
rect 357882 682398 393326 682634
rect 393562 682398 393646 682634
rect 393882 682398 429326 682634
rect 429562 682398 429646 682634
rect 429882 682398 465326 682634
rect 465562 682398 465646 682634
rect 465882 682398 501326 682634
rect 501562 682398 501646 682634
rect 501882 682398 537326 682634
rect 537562 682398 537646 682634
rect 537882 682398 573326 682634
rect 573562 682398 573646 682634
rect 573882 682398 592062 682634
rect 592298 682398 592382 682634
rect 592618 682398 592650 682634
rect -8726 682366 592650 682398
rect -8726 678454 592650 678486
rect -8726 678218 -7734 678454
rect -7498 678218 -7414 678454
rect -7178 678218 28826 678454
rect 29062 678218 29146 678454
rect 29382 678218 64826 678454
rect 65062 678218 65146 678454
rect 65382 678218 100826 678454
rect 101062 678218 101146 678454
rect 101382 678218 136826 678454
rect 137062 678218 137146 678454
rect 137382 678218 172826 678454
rect 173062 678218 173146 678454
rect 173382 678218 208826 678454
rect 209062 678218 209146 678454
rect 209382 678218 244826 678454
rect 245062 678218 245146 678454
rect 245382 678218 280826 678454
rect 281062 678218 281146 678454
rect 281382 678218 316826 678454
rect 317062 678218 317146 678454
rect 317382 678218 352826 678454
rect 353062 678218 353146 678454
rect 353382 678218 388826 678454
rect 389062 678218 389146 678454
rect 389382 678218 424826 678454
rect 425062 678218 425146 678454
rect 425382 678218 460826 678454
rect 461062 678218 461146 678454
rect 461382 678218 496826 678454
rect 497062 678218 497146 678454
rect 497382 678218 532826 678454
rect 533062 678218 533146 678454
rect 533382 678218 568826 678454
rect 569062 678218 569146 678454
rect 569382 678218 591102 678454
rect 591338 678218 591422 678454
rect 591658 678218 592650 678454
rect -8726 678134 592650 678218
rect -8726 677898 -7734 678134
rect -7498 677898 -7414 678134
rect -7178 677898 28826 678134
rect 29062 677898 29146 678134
rect 29382 677898 64826 678134
rect 65062 677898 65146 678134
rect 65382 677898 100826 678134
rect 101062 677898 101146 678134
rect 101382 677898 136826 678134
rect 137062 677898 137146 678134
rect 137382 677898 172826 678134
rect 173062 677898 173146 678134
rect 173382 677898 208826 678134
rect 209062 677898 209146 678134
rect 209382 677898 244826 678134
rect 245062 677898 245146 678134
rect 245382 677898 280826 678134
rect 281062 677898 281146 678134
rect 281382 677898 316826 678134
rect 317062 677898 317146 678134
rect 317382 677898 352826 678134
rect 353062 677898 353146 678134
rect 353382 677898 388826 678134
rect 389062 677898 389146 678134
rect 389382 677898 424826 678134
rect 425062 677898 425146 678134
rect 425382 677898 460826 678134
rect 461062 677898 461146 678134
rect 461382 677898 496826 678134
rect 497062 677898 497146 678134
rect 497382 677898 532826 678134
rect 533062 677898 533146 678134
rect 533382 677898 568826 678134
rect 569062 677898 569146 678134
rect 569382 677898 591102 678134
rect 591338 677898 591422 678134
rect 591658 677898 592650 678134
rect -8726 677866 592650 677898
rect -8726 673954 592650 673986
rect -8726 673718 -6774 673954
rect -6538 673718 -6454 673954
rect -6218 673718 24326 673954
rect 24562 673718 24646 673954
rect 24882 673718 60326 673954
rect 60562 673718 60646 673954
rect 60882 673718 96326 673954
rect 96562 673718 96646 673954
rect 96882 673718 132326 673954
rect 132562 673718 132646 673954
rect 132882 673718 168326 673954
rect 168562 673718 168646 673954
rect 168882 673718 204326 673954
rect 204562 673718 204646 673954
rect 204882 673718 240326 673954
rect 240562 673718 240646 673954
rect 240882 673718 276326 673954
rect 276562 673718 276646 673954
rect 276882 673718 312326 673954
rect 312562 673718 312646 673954
rect 312882 673718 348326 673954
rect 348562 673718 348646 673954
rect 348882 673718 384326 673954
rect 384562 673718 384646 673954
rect 384882 673718 420326 673954
rect 420562 673718 420646 673954
rect 420882 673718 456326 673954
rect 456562 673718 456646 673954
rect 456882 673718 492326 673954
rect 492562 673718 492646 673954
rect 492882 673718 528326 673954
rect 528562 673718 528646 673954
rect 528882 673718 564326 673954
rect 564562 673718 564646 673954
rect 564882 673718 590142 673954
rect 590378 673718 590462 673954
rect 590698 673718 592650 673954
rect -8726 673634 592650 673718
rect -8726 673398 -6774 673634
rect -6538 673398 -6454 673634
rect -6218 673398 24326 673634
rect 24562 673398 24646 673634
rect 24882 673398 60326 673634
rect 60562 673398 60646 673634
rect 60882 673398 96326 673634
rect 96562 673398 96646 673634
rect 96882 673398 132326 673634
rect 132562 673398 132646 673634
rect 132882 673398 168326 673634
rect 168562 673398 168646 673634
rect 168882 673398 204326 673634
rect 204562 673398 204646 673634
rect 204882 673398 240326 673634
rect 240562 673398 240646 673634
rect 240882 673398 276326 673634
rect 276562 673398 276646 673634
rect 276882 673398 312326 673634
rect 312562 673398 312646 673634
rect 312882 673398 348326 673634
rect 348562 673398 348646 673634
rect 348882 673398 384326 673634
rect 384562 673398 384646 673634
rect 384882 673398 420326 673634
rect 420562 673398 420646 673634
rect 420882 673398 456326 673634
rect 456562 673398 456646 673634
rect 456882 673398 492326 673634
rect 492562 673398 492646 673634
rect 492882 673398 528326 673634
rect 528562 673398 528646 673634
rect 528882 673398 564326 673634
rect 564562 673398 564646 673634
rect 564882 673398 590142 673634
rect 590378 673398 590462 673634
rect 590698 673398 592650 673634
rect -8726 673366 592650 673398
rect -8726 669454 592650 669486
rect -8726 669218 -5814 669454
rect -5578 669218 -5494 669454
rect -5258 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 55826 669454
rect 56062 669218 56146 669454
rect 56382 669218 91826 669454
rect 92062 669218 92146 669454
rect 92382 669218 127826 669454
rect 128062 669218 128146 669454
rect 128382 669218 163826 669454
rect 164062 669218 164146 669454
rect 164382 669218 199826 669454
rect 200062 669218 200146 669454
rect 200382 669218 235826 669454
rect 236062 669218 236146 669454
rect 236382 669218 271826 669454
rect 272062 669218 272146 669454
rect 272382 669218 307826 669454
rect 308062 669218 308146 669454
rect 308382 669218 343826 669454
rect 344062 669218 344146 669454
rect 344382 669218 379826 669454
rect 380062 669218 380146 669454
rect 380382 669218 415826 669454
rect 416062 669218 416146 669454
rect 416382 669218 451826 669454
rect 452062 669218 452146 669454
rect 452382 669218 487826 669454
rect 488062 669218 488146 669454
rect 488382 669218 523826 669454
rect 524062 669218 524146 669454
rect 524382 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 589182 669454
rect 589418 669218 589502 669454
rect 589738 669218 592650 669454
rect -8726 669134 592650 669218
rect -8726 668898 -5814 669134
rect -5578 668898 -5494 669134
rect -5258 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 55826 669134
rect 56062 668898 56146 669134
rect 56382 668898 91826 669134
rect 92062 668898 92146 669134
rect 92382 668898 127826 669134
rect 128062 668898 128146 669134
rect 128382 668898 163826 669134
rect 164062 668898 164146 669134
rect 164382 668898 199826 669134
rect 200062 668898 200146 669134
rect 200382 668898 235826 669134
rect 236062 668898 236146 669134
rect 236382 668898 271826 669134
rect 272062 668898 272146 669134
rect 272382 668898 307826 669134
rect 308062 668898 308146 669134
rect 308382 668898 343826 669134
rect 344062 668898 344146 669134
rect 344382 668898 379826 669134
rect 380062 668898 380146 669134
rect 380382 668898 415826 669134
rect 416062 668898 416146 669134
rect 416382 668898 451826 669134
rect 452062 668898 452146 669134
rect 452382 668898 487826 669134
rect 488062 668898 488146 669134
rect 488382 668898 523826 669134
rect 524062 668898 524146 669134
rect 524382 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 589182 669134
rect 589418 668898 589502 669134
rect 589738 668898 592650 669134
rect -8726 668866 592650 668898
rect -8726 664954 592650 664986
rect -8726 664718 -4854 664954
rect -4618 664718 -4534 664954
rect -4298 664718 15326 664954
rect 15562 664718 15646 664954
rect 15882 664718 51326 664954
rect 51562 664718 51646 664954
rect 51882 664718 87326 664954
rect 87562 664718 87646 664954
rect 87882 664718 123326 664954
rect 123562 664718 123646 664954
rect 123882 664718 159326 664954
rect 159562 664718 159646 664954
rect 159882 664718 195326 664954
rect 195562 664718 195646 664954
rect 195882 664718 231326 664954
rect 231562 664718 231646 664954
rect 231882 664718 267326 664954
rect 267562 664718 267646 664954
rect 267882 664718 303326 664954
rect 303562 664718 303646 664954
rect 303882 664718 339326 664954
rect 339562 664718 339646 664954
rect 339882 664718 375326 664954
rect 375562 664718 375646 664954
rect 375882 664718 411326 664954
rect 411562 664718 411646 664954
rect 411882 664718 447326 664954
rect 447562 664718 447646 664954
rect 447882 664718 483326 664954
rect 483562 664718 483646 664954
rect 483882 664718 519326 664954
rect 519562 664718 519646 664954
rect 519882 664718 555326 664954
rect 555562 664718 555646 664954
rect 555882 664718 588222 664954
rect 588458 664718 588542 664954
rect 588778 664718 592650 664954
rect -8726 664634 592650 664718
rect -8726 664398 -4854 664634
rect -4618 664398 -4534 664634
rect -4298 664398 15326 664634
rect 15562 664398 15646 664634
rect 15882 664398 51326 664634
rect 51562 664398 51646 664634
rect 51882 664398 87326 664634
rect 87562 664398 87646 664634
rect 87882 664398 123326 664634
rect 123562 664398 123646 664634
rect 123882 664398 159326 664634
rect 159562 664398 159646 664634
rect 159882 664398 195326 664634
rect 195562 664398 195646 664634
rect 195882 664398 231326 664634
rect 231562 664398 231646 664634
rect 231882 664398 267326 664634
rect 267562 664398 267646 664634
rect 267882 664398 303326 664634
rect 303562 664398 303646 664634
rect 303882 664398 339326 664634
rect 339562 664398 339646 664634
rect 339882 664398 375326 664634
rect 375562 664398 375646 664634
rect 375882 664398 411326 664634
rect 411562 664398 411646 664634
rect 411882 664398 447326 664634
rect 447562 664398 447646 664634
rect 447882 664398 483326 664634
rect 483562 664398 483646 664634
rect 483882 664398 519326 664634
rect 519562 664398 519646 664634
rect 519882 664398 555326 664634
rect 555562 664398 555646 664634
rect 555882 664398 588222 664634
rect 588458 664398 588542 664634
rect 588778 664398 592650 664634
rect -8726 664366 592650 664398
rect -8726 660454 592650 660486
rect -8726 660218 -3894 660454
rect -3658 660218 -3574 660454
rect -3338 660218 10826 660454
rect 11062 660218 11146 660454
rect 11382 660218 46826 660454
rect 47062 660218 47146 660454
rect 47382 660218 82826 660454
rect 83062 660218 83146 660454
rect 83382 660218 118826 660454
rect 119062 660218 119146 660454
rect 119382 660218 154826 660454
rect 155062 660218 155146 660454
rect 155382 660218 190826 660454
rect 191062 660218 191146 660454
rect 191382 660218 226826 660454
rect 227062 660218 227146 660454
rect 227382 660218 262826 660454
rect 263062 660218 263146 660454
rect 263382 660218 298826 660454
rect 299062 660218 299146 660454
rect 299382 660218 334826 660454
rect 335062 660218 335146 660454
rect 335382 660218 370826 660454
rect 371062 660218 371146 660454
rect 371382 660218 406826 660454
rect 407062 660218 407146 660454
rect 407382 660218 442826 660454
rect 443062 660218 443146 660454
rect 443382 660218 478826 660454
rect 479062 660218 479146 660454
rect 479382 660218 514826 660454
rect 515062 660218 515146 660454
rect 515382 660218 550826 660454
rect 551062 660218 551146 660454
rect 551382 660218 587262 660454
rect 587498 660218 587582 660454
rect 587818 660218 592650 660454
rect -8726 660134 592650 660218
rect -8726 659898 -3894 660134
rect -3658 659898 -3574 660134
rect -3338 659898 10826 660134
rect 11062 659898 11146 660134
rect 11382 659898 46826 660134
rect 47062 659898 47146 660134
rect 47382 659898 82826 660134
rect 83062 659898 83146 660134
rect 83382 659898 118826 660134
rect 119062 659898 119146 660134
rect 119382 659898 154826 660134
rect 155062 659898 155146 660134
rect 155382 659898 190826 660134
rect 191062 659898 191146 660134
rect 191382 659898 226826 660134
rect 227062 659898 227146 660134
rect 227382 659898 262826 660134
rect 263062 659898 263146 660134
rect 263382 659898 298826 660134
rect 299062 659898 299146 660134
rect 299382 659898 334826 660134
rect 335062 659898 335146 660134
rect 335382 659898 370826 660134
rect 371062 659898 371146 660134
rect 371382 659898 406826 660134
rect 407062 659898 407146 660134
rect 407382 659898 442826 660134
rect 443062 659898 443146 660134
rect 443382 659898 478826 660134
rect 479062 659898 479146 660134
rect 479382 659898 514826 660134
rect 515062 659898 515146 660134
rect 515382 659898 550826 660134
rect 551062 659898 551146 660134
rect 551382 659898 587262 660134
rect 587498 659898 587582 660134
rect 587818 659898 592650 660134
rect -8726 659866 592650 659898
rect -8726 655954 592650 655986
rect -8726 655718 -2934 655954
rect -2698 655718 -2614 655954
rect -2378 655718 6326 655954
rect 6562 655718 6646 655954
rect 6882 655718 42326 655954
rect 42562 655718 42646 655954
rect 42882 655718 78326 655954
rect 78562 655718 78646 655954
rect 78882 655718 114326 655954
rect 114562 655718 114646 655954
rect 114882 655718 150326 655954
rect 150562 655718 150646 655954
rect 150882 655718 186326 655954
rect 186562 655718 186646 655954
rect 186882 655718 222326 655954
rect 222562 655718 222646 655954
rect 222882 655718 258326 655954
rect 258562 655718 258646 655954
rect 258882 655718 294326 655954
rect 294562 655718 294646 655954
rect 294882 655718 330326 655954
rect 330562 655718 330646 655954
rect 330882 655718 366326 655954
rect 366562 655718 366646 655954
rect 366882 655718 402326 655954
rect 402562 655718 402646 655954
rect 402882 655718 438326 655954
rect 438562 655718 438646 655954
rect 438882 655718 474326 655954
rect 474562 655718 474646 655954
rect 474882 655718 510326 655954
rect 510562 655718 510646 655954
rect 510882 655718 546326 655954
rect 546562 655718 546646 655954
rect 546882 655718 582326 655954
rect 582562 655718 582646 655954
rect 582882 655718 586302 655954
rect 586538 655718 586622 655954
rect 586858 655718 592650 655954
rect -8726 655634 592650 655718
rect -8726 655398 -2934 655634
rect -2698 655398 -2614 655634
rect -2378 655398 6326 655634
rect 6562 655398 6646 655634
rect 6882 655398 42326 655634
rect 42562 655398 42646 655634
rect 42882 655398 78326 655634
rect 78562 655398 78646 655634
rect 78882 655398 114326 655634
rect 114562 655398 114646 655634
rect 114882 655398 150326 655634
rect 150562 655398 150646 655634
rect 150882 655398 186326 655634
rect 186562 655398 186646 655634
rect 186882 655398 222326 655634
rect 222562 655398 222646 655634
rect 222882 655398 258326 655634
rect 258562 655398 258646 655634
rect 258882 655398 294326 655634
rect 294562 655398 294646 655634
rect 294882 655398 330326 655634
rect 330562 655398 330646 655634
rect 330882 655398 366326 655634
rect 366562 655398 366646 655634
rect 366882 655398 402326 655634
rect 402562 655398 402646 655634
rect 402882 655398 438326 655634
rect 438562 655398 438646 655634
rect 438882 655398 474326 655634
rect 474562 655398 474646 655634
rect 474882 655398 510326 655634
rect 510562 655398 510646 655634
rect 510882 655398 546326 655634
rect 546562 655398 546646 655634
rect 546882 655398 582326 655634
rect 582562 655398 582646 655634
rect 582882 655398 586302 655634
rect 586538 655398 586622 655634
rect 586858 655398 592650 655634
rect -8726 655366 592650 655398
rect -8726 651454 592650 651486
rect -8726 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 109826 651454
rect 110062 651218 110146 651454
rect 110382 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 592650 651454
rect -8726 651134 592650 651218
rect -8726 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 109826 651134
rect 110062 650898 110146 651134
rect 110382 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 592650 651134
rect -8726 650866 592650 650898
rect -8726 646954 592650 646986
rect -8726 646718 -8694 646954
rect -8458 646718 -8374 646954
rect -8138 646718 33326 646954
rect 33562 646718 33646 646954
rect 33882 646718 69326 646954
rect 69562 646718 69646 646954
rect 69882 646718 105326 646954
rect 105562 646718 105646 646954
rect 105882 646718 141326 646954
rect 141562 646718 141646 646954
rect 141882 646718 177326 646954
rect 177562 646718 177646 646954
rect 177882 646718 213326 646954
rect 213562 646718 213646 646954
rect 213882 646718 249326 646954
rect 249562 646718 249646 646954
rect 249882 646718 285326 646954
rect 285562 646718 285646 646954
rect 285882 646718 321326 646954
rect 321562 646718 321646 646954
rect 321882 646718 357326 646954
rect 357562 646718 357646 646954
rect 357882 646718 393326 646954
rect 393562 646718 393646 646954
rect 393882 646718 429326 646954
rect 429562 646718 429646 646954
rect 429882 646718 465326 646954
rect 465562 646718 465646 646954
rect 465882 646718 501326 646954
rect 501562 646718 501646 646954
rect 501882 646718 537326 646954
rect 537562 646718 537646 646954
rect 537882 646718 573326 646954
rect 573562 646718 573646 646954
rect 573882 646718 592062 646954
rect 592298 646718 592382 646954
rect 592618 646718 592650 646954
rect -8726 646634 592650 646718
rect -8726 646398 -8694 646634
rect -8458 646398 -8374 646634
rect -8138 646398 33326 646634
rect 33562 646398 33646 646634
rect 33882 646398 69326 646634
rect 69562 646398 69646 646634
rect 69882 646398 105326 646634
rect 105562 646398 105646 646634
rect 105882 646398 141326 646634
rect 141562 646398 141646 646634
rect 141882 646398 177326 646634
rect 177562 646398 177646 646634
rect 177882 646398 213326 646634
rect 213562 646398 213646 646634
rect 213882 646398 249326 646634
rect 249562 646398 249646 646634
rect 249882 646398 285326 646634
rect 285562 646398 285646 646634
rect 285882 646398 321326 646634
rect 321562 646398 321646 646634
rect 321882 646398 357326 646634
rect 357562 646398 357646 646634
rect 357882 646398 393326 646634
rect 393562 646398 393646 646634
rect 393882 646398 429326 646634
rect 429562 646398 429646 646634
rect 429882 646398 465326 646634
rect 465562 646398 465646 646634
rect 465882 646398 501326 646634
rect 501562 646398 501646 646634
rect 501882 646398 537326 646634
rect 537562 646398 537646 646634
rect 537882 646398 573326 646634
rect 573562 646398 573646 646634
rect 573882 646398 592062 646634
rect 592298 646398 592382 646634
rect 592618 646398 592650 646634
rect -8726 646366 592650 646398
rect -8726 642454 592650 642486
rect -8726 642218 -7734 642454
rect -7498 642218 -7414 642454
rect -7178 642218 28826 642454
rect 29062 642218 29146 642454
rect 29382 642218 64826 642454
rect 65062 642218 65146 642454
rect 65382 642218 100826 642454
rect 101062 642218 101146 642454
rect 101382 642218 136826 642454
rect 137062 642218 137146 642454
rect 137382 642218 172826 642454
rect 173062 642218 173146 642454
rect 173382 642218 208826 642454
rect 209062 642218 209146 642454
rect 209382 642218 244826 642454
rect 245062 642218 245146 642454
rect 245382 642218 280826 642454
rect 281062 642218 281146 642454
rect 281382 642218 316826 642454
rect 317062 642218 317146 642454
rect 317382 642218 352826 642454
rect 353062 642218 353146 642454
rect 353382 642218 388826 642454
rect 389062 642218 389146 642454
rect 389382 642218 424826 642454
rect 425062 642218 425146 642454
rect 425382 642218 460826 642454
rect 461062 642218 461146 642454
rect 461382 642218 496826 642454
rect 497062 642218 497146 642454
rect 497382 642218 532826 642454
rect 533062 642218 533146 642454
rect 533382 642218 568826 642454
rect 569062 642218 569146 642454
rect 569382 642218 591102 642454
rect 591338 642218 591422 642454
rect 591658 642218 592650 642454
rect -8726 642134 592650 642218
rect -8726 641898 -7734 642134
rect -7498 641898 -7414 642134
rect -7178 641898 28826 642134
rect 29062 641898 29146 642134
rect 29382 641898 64826 642134
rect 65062 641898 65146 642134
rect 65382 641898 100826 642134
rect 101062 641898 101146 642134
rect 101382 641898 136826 642134
rect 137062 641898 137146 642134
rect 137382 641898 172826 642134
rect 173062 641898 173146 642134
rect 173382 641898 208826 642134
rect 209062 641898 209146 642134
rect 209382 641898 244826 642134
rect 245062 641898 245146 642134
rect 245382 641898 280826 642134
rect 281062 641898 281146 642134
rect 281382 641898 316826 642134
rect 317062 641898 317146 642134
rect 317382 641898 352826 642134
rect 353062 641898 353146 642134
rect 353382 641898 388826 642134
rect 389062 641898 389146 642134
rect 389382 641898 424826 642134
rect 425062 641898 425146 642134
rect 425382 641898 460826 642134
rect 461062 641898 461146 642134
rect 461382 641898 496826 642134
rect 497062 641898 497146 642134
rect 497382 641898 532826 642134
rect 533062 641898 533146 642134
rect 533382 641898 568826 642134
rect 569062 641898 569146 642134
rect 569382 641898 591102 642134
rect 591338 641898 591422 642134
rect 591658 641898 592650 642134
rect -8726 641866 592650 641898
rect -8726 637954 592650 637986
rect -8726 637718 -6774 637954
rect -6538 637718 -6454 637954
rect -6218 637718 24326 637954
rect 24562 637718 24646 637954
rect 24882 637718 60326 637954
rect 60562 637718 60646 637954
rect 60882 637718 96326 637954
rect 96562 637718 96646 637954
rect 96882 637718 132326 637954
rect 132562 637718 132646 637954
rect 132882 637718 168326 637954
rect 168562 637718 168646 637954
rect 168882 637718 204326 637954
rect 204562 637718 204646 637954
rect 204882 637718 240326 637954
rect 240562 637718 240646 637954
rect 240882 637718 276326 637954
rect 276562 637718 276646 637954
rect 276882 637718 312326 637954
rect 312562 637718 312646 637954
rect 312882 637718 348326 637954
rect 348562 637718 348646 637954
rect 348882 637718 384326 637954
rect 384562 637718 384646 637954
rect 384882 637718 420326 637954
rect 420562 637718 420646 637954
rect 420882 637718 456326 637954
rect 456562 637718 456646 637954
rect 456882 637718 492326 637954
rect 492562 637718 492646 637954
rect 492882 637718 528326 637954
rect 528562 637718 528646 637954
rect 528882 637718 564326 637954
rect 564562 637718 564646 637954
rect 564882 637718 590142 637954
rect 590378 637718 590462 637954
rect 590698 637718 592650 637954
rect -8726 637634 592650 637718
rect -8726 637398 -6774 637634
rect -6538 637398 -6454 637634
rect -6218 637398 24326 637634
rect 24562 637398 24646 637634
rect 24882 637398 60326 637634
rect 60562 637398 60646 637634
rect 60882 637398 96326 637634
rect 96562 637398 96646 637634
rect 96882 637398 132326 637634
rect 132562 637398 132646 637634
rect 132882 637398 168326 637634
rect 168562 637398 168646 637634
rect 168882 637398 204326 637634
rect 204562 637398 204646 637634
rect 204882 637398 240326 637634
rect 240562 637398 240646 637634
rect 240882 637398 276326 637634
rect 276562 637398 276646 637634
rect 276882 637398 312326 637634
rect 312562 637398 312646 637634
rect 312882 637398 348326 637634
rect 348562 637398 348646 637634
rect 348882 637398 384326 637634
rect 384562 637398 384646 637634
rect 384882 637398 420326 637634
rect 420562 637398 420646 637634
rect 420882 637398 456326 637634
rect 456562 637398 456646 637634
rect 456882 637398 492326 637634
rect 492562 637398 492646 637634
rect 492882 637398 528326 637634
rect 528562 637398 528646 637634
rect 528882 637398 564326 637634
rect 564562 637398 564646 637634
rect 564882 637398 590142 637634
rect 590378 637398 590462 637634
rect 590698 637398 592650 637634
rect -8726 637366 592650 637398
rect -8726 633454 592650 633486
rect -8726 633218 -5814 633454
rect -5578 633218 -5494 633454
rect -5258 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 55826 633454
rect 56062 633218 56146 633454
rect 56382 633218 91826 633454
rect 92062 633218 92146 633454
rect 92382 633218 127826 633454
rect 128062 633218 128146 633454
rect 128382 633218 163826 633454
rect 164062 633218 164146 633454
rect 164382 633218 199826 633454
rect 200062 633218 200146 633454
rect 200382 633218 235826 633454
rect 236062 633218 236146 633454
rect 236382 633218 271826 633454
rect 272062 633218 272146 633454
rect 272382 633218 307826 633454
rect 308062 633218 308146 633454
rect 308382 633218 343826 633454
rect 344062 633218 344146 633454
rect 344382 633218 379826 633454
rect 380062 633218 380146 633454
rect 380382 633218 415826 633454
rect 416062 633218 416146 633454
rect 416382 633218 451826 633454
rect 452062 633218 452146 633454
rect 452382 633218 487826 633454
rect 488062 633218 488146 633454
rect 488382 633218 523826 633454
rect 524062 633218 524146 633454
rect 524382 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 589182 633454
rect 589418 633218 589502 633454
rect 589738 633218 592650 633454
rect -8726 633134 592650 633218
rect -8726 632898 -5814 633134
rect -5578 632898 -5494 633134
rect -5258 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 55826 633134
rect 56062 632898 56146 633134
rect 56382 632898 91826 633134
rect 92062 632898 92146 633134
rect 92382 632898 127826 633134
rect 128062 632898 128146 633134
rect 128382 632898 163826 633134
rect 164062 632898 164146 633134
rect 164382 632898 199826 633134
rect 200062 632898 200146 633134
rect 200382 632898 235826 633134
rect 236062 632898 236146 633134
rect 236382 632898 271826 633134
rect 272062 632898 272146 633134
rect 272382 632898 307826 633134
rect 308062 632898 308146 633134
rect 308382 632898 343826 633134
rect 344062 632898 344146 633134
rect 344382 632898 379826 633134
rect 380062 632898 380146 633134
rect 380382 632898 415826 633134
rect 416062 632898 416146 633134
rect 416382 632898 451826 633134
rect 452062 632898 452146 633134
rect 452382 632898 487826 633134
rect 488062 632898 488146 633134
rect 488382 632898 523826 633134
rect 524062 632898 524146 633134
rect 524382 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 589182 633134
rect 589418 632898 589502 633134
rect 589738 632898 592650 633134
rect -8726 632866 592650 632898
rect -8726 628954 592650 628986
rect -8726 628718 -4854 628954
rect -4618 628718 -4534 628954
rect -4298 628718 15326 628954
rect 15562 628718 15646 628954
rect 15882 628718 51326 628954
rect 51562 628718 51646 628954
rect 51882 628718 87326 628954
rect 87562 628718 87646 628954
rect 87882 628718 123326 628954
rect 123562 628718 123646 628954
rect 123882 628718 159326 628954
rect 159562 628718 159646 628954
rect 159882 628718 195326 628954
rect 195562 628718 195646 628954
rect 195882 628718 231326 628954
rect 231562 628718 231646 628954
rect 231882 628718 267326 628954
rect 267562 628718 267646 628954
rect 267882 628718 303326 628954
rect 303562 628718 303646 628954
rect 303882 628718 339326 628954
rect 339562 628718 339646 628954
rect 339882 628718 375326 628954
rect 375562 628718 375646 628954
rect 375882 628718 411326 628954
rect 411562 628718 411646 628954
rect 411882 628718 447326 628954
rect 447562 628718 447646 628954
rect 447882 628718 483326 628954
rect 483562 628718 483646 628954
rect 483882 628718 519326 628954
rect 519562 628718 519646 628954
rect 519882 628718 555326 628954
rect 555562 628718 555646 628954
rect 555882 628718 588222 628954
rect 588458 628718 588542 628954
rect 588778 628718 592650 628954
rect -8726 628634 592650 628718
rect -8726 628398 -4854 628634
rect -4618 628398 -4534 628634
rect -4298 628398 15326 628634
rect 15562 628398 15646 628634
rect 15882 628398 51326 628634
rect 51562 628398 51646 628634
rect 51882 628398 87326 628634
rect 87562 628398 87646 628634
rect 87882 628398 123326 628634
rect 123562 628398 123646 628634
rect 123882 628398 159326 628634
rect 159562 628398 159646 628634
rect 159882 628398 195326 628634
rect 195562 628398 195646 628634
rect 195882 628398 231326 628634
rect 231562 628398 231646 628634
rect 231882 628398 267326 628634
rect 267562 628398 267646 628634
rect 267882 628398 303326 628634
rect 303562 628398 303646 628634
rect 303882 628398 339326 628634
rect 339562 628398 339646 628634
rect 339882 628398 375326 628634
rect 375562 628398 375646 628634
rect 375882 628398 411326 628634
rect 411562 628398 411646 628634
rect 411882 628398 447326 628634
rect 447562 628398 447646 628634
rect 447882 628398 483326 628634
rect 483562 628398 483646 628634
rect 483882 628398 519326 628634
rect 519562 628398 519646 628634
rect 519882 628398 555326 628634
rect 555562 628398 555646 628634
rect 555882 628398 588222 628634
rect 588458 628398 588542 628634
rect 588778 628398 592650 628634
rect -8726 628366 592650 628398
rect -8726 624454 592650 624486
rect -8726 624218 -3894 624454
rect -3658 624218 -3574 624454
rect -3338 624218 10826 624454
rect 11062 624218 11146 624454
rect 11382 624218 46826 624454
rect 47062 624218 47146 624454
rect 47382 624218 82826 624454
rect 83062 624218 83146 624454
rect 83382 624218 118826 624454
rect 119062 624218 119146 624454
rect 119382 624218 154826 624454
rect 155062 624218 155146 624454
rect 155382 624218 190826 624454
rect 191062 624218 191146 624454
rect 191382 624218 226826 624454
rect 227062 624218 227146 624454
rect 227382 624218 262826 624454
rect 263062 624218 263146 624454
rect 263382 624218 298826 624454
rect 299062 624218 299146 624454
rect 299382 624218 334826 624454
rect 335062 624218 335146 624454
rect 335382 624218 370826 624454
rect 371062 624218 371146 624454
rect 371382 624218 406826 624454
rect 407062 624218 407146 624454
rect 407382 624218 442826 624454
rect 443062 624218 443146 624454
rect 443382 624218 478826 624454
rect 479062 624218 479146 624454
rect 479382 624218 514826 624454
rect 515062 624218 515146 624454
rect 515382 624218 550826 624454
rect 551062 624218 551146 624454
rect 551382 624218 587262 624454
rect 587498 624218 587582 624454
rect 587818 624218 592650 624454
rect -8726 624134 592650 624218
rect -8726 623898 -3894 624134
rect -3658 623898 -3574 624134
rect -3338 623898 10826 624134
rect 11062 623898 11146 624134
rect 11382 623898 46826 624134
rect 47062 623898 47146 624134
rect 47382 623898 82826 624134
rect 83062 623898 83146 624134
rect 83382 623898 118826 624134
rect 119062 623898 119146 624134
rect 119382 623898 154826 624134
rect 155062 623898 155146 624134
rect 155382 623898 190826 624134
rect 191062 623898 191146 624134
rect 191382 623898 226826 624134
rect 227062 623898 227146 624134
rect 227382 623898 262826 624134
rect 263062 623898 263146 624134
rect 263382 623898 298826 624134
rect 299062 623898 299146 624134
rect 299382 623898 334826 624134
rect 335062 623898 335146 624134
rect 335382 623898 370826 624134
rect 371062 623898 371146 624134
rect 371382 623898 406826 624134
rect 407062 623898 407146 624134
rect 407382 623898 442826 624134
rect 443062 623898 443146 624134
rect 443382 623898 478826 624134
rect 479062 623898 479146 624134
rect 479382 623898 514826 624134
rect 515062 623898 515146 624134
rect 515382 623898 550826 624134
rect 551062 623898 551146 624134
rect 551382 623898 587262 624134
rect 587498 623898 587582 624134
rect 587818 623898 592650 624134
rect -8726 623866 592650 623898
rect -8726 619954 592650 619986
rect -8726 619718 -2934 619954
rect -2698 619718 -2614 619954
rect -2378 619718 6326 619954
rect 6562 619718 6646 619954
rect 6882 619718 42326 619954
rect 42562 619718 42646 619954
rect 42882 619718 78326 619954
rect 78562 619718 78646 619954
rect 78882 619718 114326 619954
rect 114562 619718 114646 619954
rect 114882 619718 150326 619954
rect 150562 619718 150646 619954
rect 150882 619718 186326 619954
rect 186562 619718 186646 619954
rect 186882 619718 222326 619954
rect 222562 619718 222646 619954
rect 222882 619718 258326 619954
rect 258562 619718 258646 619954
rect 258882 619718 294326 619954
rect 294562 619718 294646 619954
rect 294882 619718 330326 619954
rect 330562 619718 330646 619954
rect 330882 619718 366326 619954
rect 366562 619718 366646 619954
rect 366882 619718 402326 619954
rect 402562 619718 402646 619954
rect 402882 619718 438326 619954
rect 438562 619718 438646 619954
rect 438882 619718 474326 619954
rect 474562 619718 474646 619954
rect 474882 619718 510326 619954
rect 510562 619718 510646 619954
rect 510882 619718 546326 619954
rect 546562 619718 546646 619954
rect 546882 619718 582326 619954
rect 582562 619718 582646 619954
rect 582882 619718 586302 619954
rect 586538 619718 586622 619954
rect 586858 619718 592650 619954
rect -8726 619634 592650 619718
rect -8726 619398 -2934 619634
rect -2698 619398 -2614 619634
rect -2378 619398 6326 619634
rect 6562 619398 6646 619634
rect 6882 619398 42326 619634
rect 42562 619398 42646 619634
rect 42882 619398 78326 619634
rect 78562 619398 78646 619634
rect 78882 619398 114326 619634
rect 114562 619398 114646 619634
rect 114882 619398 150326 619634
rect 150562 619398 150646 619634
rect 150882 619398 186326 619634
rect 186562 619398 186646 619634
rect 186882 619398 222326 619634
rect 222562 619398 222646 619634
rect 222882 619398 258326 619634
rect 258562 619398 258646 619634
rect 258882 619398 294326 619634
rect 294562 619398 294646 619634
rect 294882 619398 330326 619634
rect 330562 619398 330646 619634
rect 330882 619398 366326 619634
rect 366562 619398 366646 619634
rect 366882 619398 402326 619634
rect 402562 619398 402646 619634
rect 402882 619398 438326 619634
rect 438562 619398 438646 619634
rect 438882 619398 474326 619634
rect 474562 619398 474646 619634
rect 474882 619398 510326 619634
rect 510562 619398 510646 619634
rect 510882 619398 546326 619634
rect 546562 619398 546646 619634
rect 546882 619398 582326 619634
rect 582562 619398 582646 619634
rect 582882 619398 586302 619634
rect 586538 619398 586622 619634
rect 586858 619398 592650 619634
rect -8726 619366 592650 619398
rect -8726 615454 592650 615486
rect -8726 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 73826 615454
rect 74062 615218 74146 615454
rect 74382 615218 109826 615454
rect 110062 615218 110146 615454
rect 110382 615218 145826 615454
rect 146062 615218 146146 615454
rect 146382 615218 181826 615454
rect 182062 615218 182146 615454
rect 182382 615218 217826 615454
rect 218062 615218 218146 615454
rect 218382 615218 253826 615454
rect 254062 615218 254146 615454
rect 254382 615218 289826 615454
rect 290062 615218 290146 615454
rect 290382 615218 325826 615454
rect 326062 615218 326146 615454
rect 326382 615218 361826 615454
rect 362062 615218 362146 615454
rect 362382 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 469826 615454
rect 470062 615218 470146 615454
rect 470382 615218 505826 615454
rect 506062 615218 506146 615454
rect 506382 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 592650 615454
rect -8726 615134 592650 615218
rect -8726 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 73826 615134
rect 74062 614898 74146 615134
rect 74382 614898 109826 615134
rect 110062 614898 110146 615134
rect 110382 614898 145826 615134
rect 146062 614898 146146 615134
rect 146382 614898 181826 615134
rect 182062 614898 182146 615134
rect 182382 614898 217826 615134
rect 218062 614898 218146 615134
rect 218382 614898 253826 615134
rect 254062 614898 254146 615134
rect 254382 614898 289826 615134
rect 290062 614898 290146 615134
rect 290382 614898 325826 615134
rect 326062 614898 326146 615134
rect 326382 614898 361826 615134
rect 362062 614898 362146 615134
rect 362382 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 469826 615134
rect 470062 614898 470146 615134
rect 470382 614898 505826 615134
rect 506062 614898 506146 615134
rect 506382 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 592650 615134
rect -8726 614866 592650 614898
rect -8726 610954 592650 610986
rect -8726 610718 -8694 610954
rect -8458 610718 -8374 610954
rect -8138 610718 33326 610954
rect 33562 610718 33646 610954
rect 33882 610718 69326 610954
rect 69562 610718 69646 610954
rect 69882 610718 105326 610954
rect 105562 610718 105646 610954
rect 105882 610718 141326 610954
rect 141562 610718 141646 610954
rect 141882 610718 177326 610954
rect 177562 610718 177646 610954
rect 177882 610718 213326 610954
rect 213562 610718 213646 610954
rect 213882 610718 249326 610954
rect 249562 610718 249646 610954
rect 249882 610718 285326 610954
rect 285562 610718 285646 610954
rect 285882 610718 321326 610954
rect 321562 610718 321646 610954
rect 321882 610718 357326 610954
rect 357562 610718 357646 610954
rect 357882 610718 393326 610954
rect 393562 610718 393646 610954
rect 393882 610718 429326 610954
rect 429562 610718 429646 610954
rect 429882 610718 465326 610954
rect 465562 610718 465646 610954
rect 465882 610718 501326 610954
rect 501562 610718 501646 610954
rect 501882 610718 537326 610954
rect 537562 610718 537646 610954
rect 537882 610718 573326 610954
rect 573562 610718 573646 610954
rect 573882 610718 592062 610954
rect 592298 610718 592382 610954
rect 592618 610718 592650 610954
rect -8726 610634 592650 610718
rect -8726 610398 -8694 610634
rect -8458 610398 -8374 610634
rect -8138 610398 33326 610634
rect 33562 610398 33646 610634
rect 33882 610398 69326 610634
rect 69562 610398 69646 610634
rect 69882 610398 105326 610634
rect 105562 610398 105646 610634
rect 105882 610398 141326 610634
rect 141562 610398 141646 610634
rect 141882 610398 177326 610634
rect 177562 610398 177646 610634
rect 177882 610398 213326 610634
rect 213562 610398 213646 610634
rect 213882 610398 249326 610634
rect 249562 610398 249646 610634
rect 249882 610398 285326 610634
rect 285562 610398 285646 610634
rect 285882 610398 321326 610634
rect 321562 610398 321646 610634
rect 321882 610398 357326 610634
rect 357562 610398 357646 610634
rect 357882 610398 393326 610634
rect 393562 610398 393646 610634
rect 393882 610398 429326 610634
rect 429562 610398 429646 610634
rect 429882 610398 465326 610634
rect 465562 610398 465646 610634
rect 465882 610398 501326 610634
rect 501562 610398 501646 610634
rect 501882 610398 537326 610634
rect 537562 610398 537646 610634
rect 537882 610398 573326 610634
rect 573562 610398 573646 610634
rect 573882 610398 592062 610634
rect 592298 610398 592382 610634
rect 592618 610398 592650 610634
rect -8726 610366 592650 610398
rect -8726 606454 592650 606486
rect -8726 606218 -7734 606454
rect -7498 606218 -7414 606454
rect -7178 606218 28826 606454
rect 29062 606218 29146 606454
rect 29382 606218 64826 606454
rect 65062 606218 65146 606454
rect 65382 606218 100826 606454
rect 101062 606218 101146 606454
rect 101382 606218 136826 606454
rect 137062 606218 137146 606454
rect 137382 606218 172826 606454
rect 173062 606218 173146 606454
rect 173382 606218 208826 606454
rect 209062 606218 209146 606454
rect 209382 606218 244826 606454
rect 245062 606218 245146 606454
rect 245382 606218 280826 606454
rect 281062 606218 281146 606454
rect 281382 606218 316826 606454
rect 317062 606218 317146 606454
rect 317382 606218 352826 606454
rect 353062 606218 353146 606454
rect 353382 606218 388826 606454
rect 389062 606218 389146 606454
rect 389382 606218 424826 606454
rect 425062 606218 425146 606454
rect 425382 606218 460826 606454
rect 461062 606218 461146 606454
rect 461382 606218 496826 606454
rect 497062 606218 497146 606454
rect 497382 606218 532826 606454
rect 533062 606218 533146 606454
rect 533382 606218 568826 606454
rect 569062 606218 569146 606454
rect 569382 606218 591102 606454
rect 591338 606218 591422 606454
rect 591658 606218 592650 606454
rect -8726 606134 592650 606218
rect -8726 605898 -7734 606134
rect -7498 605898 -7414 606134
rect -7178 605898 28826 606134
rect 29062 605898 29146 606134
rect 29382 605898 64826 606134
rect 65062 605898 65146 606134
rect 65382 605898 100826 606134
rect 101062 605898 101146 606134
rect 101382 605898 136826 606134
rect 137062 605898 137146 606134
rect 137382 605898 172826 606134
rect 173062 605898 173146 606134
rect 173382 605898 208826 606134
rect 209062 605898 209146 606134
rect 209382 605898 244826 606134
rect 245062 605898 245146 606134
rect 245382 605898 280826 606134
rect 281062 605898 281146 606134
rect 281382 605898 316826 606134
rect 317062 605898 317146 606134
rect 317382 605898 352826 606134
rect 353062 605898 353146 606134
rect 353382 605898 388826 606134
rect 389062 605898 389146 606134
rect 389382 605898 424826 606134
rect 425062 605898 425146 606134
rect 425382 605898 460826 606134
rect 461062 605898 461146 606134
rect 461382 605898 496826 606134
rect 497062 605898 497146 606134
rect 497382 605898 532826 606134
rect 533062 605898 533146 606134
rect 533382 605898 568826 606134
rect 569062 605898 569146 606134
rect 569382 605898 591102 606134
rect 591338 605898 591422 606134
rect 591658 605898 592650 606134
rect -8726 605866 592650 605898
rect -8726 601954 592650 601986
rect -8726 601718 -6774 601954
rect -6538 601718 -6454 601954
rect -6218 601718 24326 601954
rect 24562 601718 24646 601954
rect 24882 601718 60326 601954
rect 60562 601718 60646 601954
rect 60882 601718 96326 601954
rect 96562 601718 96646 601954
rect 96882 601718 132326 601954
rect 132562 601718 132646 601954
rect 132882 601718 168326 601954
rect 168562 601718 168646 601954
rect 168882 601718 204326 601954
rect 204562 601718 204646 601954
rect 204882 601718 240326 601954
rect 240562 601718 240646 601954
rect 240882 601718 276326 601954
rect 276562 601718 276646 601954
rect 276882 601718 312326 601954
rect 312562 601718 312646 601954
rect 312882 601718 348326 601954
rect 348562 601718 348646 601954
rect 348882 601718 384326 601954
rect 384562 601718 384646 601954
rect 384882 601718 420326 601954
rect 420562 601718 420646 601954
rect 420882 601718 456326 601954
rect 456562 601718 456646 601954
rect 456882 601718 492326 601954
rect 492562 601718 492646 601954
rect 492882 601718 528326 601954
rect 528562 601718 528646 601954
rect 528882 601718 564326 601954
rect 564562 601718 564646 601954
rect 564882 601718 590142 601954
rect 590378 601718 590462 601954
rect 590698 601718 592650 601954
rect -8726 601634 592650 601718
rect -8726 601398 -6774 601634
rect -6538 601398 -6454 601634
rect -6218 601398 24326 601634
rect 24562 601398 24646 601634
rect 24882 601398 60326 601634
rect 60562 601398 60646 601634
rect 60882 601398 96326 601634
rect 96562 601398 96646 601634
rect 96882 601398 132326 601634
rect 132562 601398 132646 601634
rect 132882 601398 168326 601634
rect 168562 601398 168646 601634
rect 168882 601398 204326 601634
rect 204562 601398 204646 601634
rect 204882 601398 240326 601634
rect 240562 601398 240646 601634
rect 240882 601398 276326 601634
rect 276562 601398 276646 601634
rect 276882 601398 312326 601634
rect 312562 601398 312646 601634
rect 312882 601398 348326 601634
rect 348562 601398 348646 601634
rect 348882 601398 384326 601634
rect 384562 601398 384646 601634
rect 384882 601398 420326 601634
rect 420562 601398 420646 601634
rect 420882 601398 456326 601634
rect 456562 601398 456646 601634
rect 456882 601398 492326 601634
rect 492562 601398 492646 601634
rect 492882 601398 528326 601634
rect 528562 601398 528646 601634
rect 528882 601398 564326 601634
rect 564562 601398 564646 601634
rect 564882 601398 590142 601634
rect 590378 601398 590462 601634
rect 590698 601398 592650 601634
rect -8726 601366 592650 601398
rect -8726 597454 592650 597486
rect -8726 597218 -5814 597454
rect -5578 597218 -5494 597454
rect -5258 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 55826 597454
rect 56062 597218 56146 597454
rect 56382 597218 91826 597454
rect 92062 597218 92146 597454
rect 92382 597218 127826 597454
rect 128062 597218 128146 597454
rect 128382 597218 163826 597454
rect 164062 597218 164146 597454
rect 164382 597218 199826 597454
rect 200062 597218 200146 597454
rect 200382 597218 235826 597454
rect 236062 597218 236146 597454
rect 236382 597218 271826 597454
rect 272062 597218 272146 597454
rect 272382 597218 307826 597454
rect 308062 597218 308146 597454
rect 308382 597218 343826 597454
rect 344062 597218 344146 597454
rect 344382 597218 379826 597454
rect 380062 597218 380146 597454
rect 380382 597218 415826 597454
rect 416062 597218 416146 597454
rect 416382 597218 451826 597454
rect 452062 597218 452146 597454
rect 452382 597218 487826 597454
rect 488062 597218 488146 597454
rect 488382 597218 523826 597454
rect 524062 597218 524146 597454
rect 524382 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 589182 597454
rect 589418 597218 589502 597454
rect 589738 597218 592650 597454
rect -8726 597134 592650 597218
rect -8726 596898 -5814 597134
rect -5578 596898 -5494 597134
rect -5258 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 55826 597134
rect 56062 596898 56146 597134
rect 56382 596898 91826 597134
rect 92062 596898 92146 597134
rect 92382 596898 127826 597134
rect 128062 596898 128146 597134
rect 128382 596898 163826 597134
rect 164062 596898 164146 597134
rect 164382 596898 199826 597134
rect 200062 596898 200146 597134
rect 200382 596898 235826 597134
rect 236062 596898 236146 597134
rect 236382 596898 271826 597134
rect 272062 596898 272146 597134
rect 272382 596898 307826 597134
rect 308062 596898 308146 597134
rect 308382 596898 343826 597134
rect 344062 596898 344146 597134
rect 344382 596898 379826 597134
rect 380062 596898 380146 597134
rect 380382 596898 415826 597134
rect 416062 596898 416146 597134
rect 416382 596898 451826 597134
rect 452062 596898 452146 597134
rect 452382 596898 487826 597134
rect 488062 596898 488146 597134
rect 488382 596898 523826 597134
rect 524062 596898 524146 597134
rect 524382 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 589182 597134
rect 589418 596898 589502 597134
rect 589738 596898 592650 597134
rect -8726 596866 592650 596898
rect -8726 592954 592650 592986
rect -8726 592718 -4854 592954
rect -4618 592718 -4534 592954
rect -4298 592718 15326 592954
rect 15562 592718 15646 592954
rect 15882 592718 51326 592954
rect 51562 592718 51646 592954
rect 51882 592718 87326 592954
rect 87562 592718 87646 592954
rect 87882 592718 123326 592954
rect 123562 592718 123646 592954
rect 123882 592718 159326 592954
rect 159562 592718 159646 592954
rect 159882 592718 195326 592954
rect 195562 592718 195646 592954
rect 195882 592718 231326 592954
rect 231562 592718 231646 592954
rect 231882 592718 267326 592954
rect 267562 592718 267646 592954
rect 267882 592718 303326 592954
rect 303562 592718 303646 592954
rect 303882 592718 339326 592954
rect 339562 592718 339646 592954
rect 339882 592718 375326 592954
rect 375562 592718 375646 592954
rect 375882 592718 411326 592954
rect 411562 592718 411646 592954
rect 411882 592718 447326 592954
rect 447562 592718 447646 592954
rect 447882 592718 483326 592954
rect 483562 592718 483646 592954
rect 483882 592718 519326 592954
rect 519562 592718 519646 592954
rect 519882 592718 555326 592954
rect 555562 592718 555646 592954
rect 555882 592718 588222 592954
rect 588458 592718 588542 592954
rect 588778 592718 592650 592954
rect -8726 592634 592650 592718
rect -8726 592398 -4854 592634
rect -4618 592398 -4534 592634
rect -4298 592398 15326 592634
rect 15562 592398 15646 592634
rect 15882 592398 51326 592634
rect 51562 592398 51646 592634
rect 51882 592398 87326 592634
rect 87562 592398 87646 592634
rect 87882 592398 123326 592634
rect 123562 592398 123646 592634
rect 123882 592398 159326 592634
rect 159562 592398 159646 592634
rect 159882 592398 195326 592634
rect 195562 592398 195646 592634
rect 195882 592398 231326 592634
rect 231562 592398 231646 592634
rect 231882 592398 267326 592634
rect 267562 592398 267646 592634
rect 267882 592398 303326 592634
rect 303562 592398 303646 592634
rect 303882 592398 339326 592634
rect 339562 592398 339646 592634
rect 339882 592398 375326 592634
rect 375562 592398 375646 592634
rect 375882 592398 411326 592634
rect 411562 592398 411646 592634
rect 411882 592398 447326 592634
rect 447562 592398 447646 592634
rect 447882 592398 483326 592634
rect 483562 592398 483646 592634
rect 483882 592398 519326 592634
rect 519562 592398 519646 592634
rect 519882 592398 555326 592634
rect 555562 592398 555646 592634
rect 555882 592398 588222 592634
rect 588458 592398 588542 592634
rect 588778 592398 592650 592634
rect -8726 592366 592650 592398
rect -8726 588454 592650 588486
rect -8726 588218 -3894 588454
rect -3658 588218 -3574 588454
rect -3338 588218 10826 588454
rect 11062 588218 11146 588454
rect 11382 588218 46826 588454
rect 47062 588218 47146 588454
rect 47382 588218 82826 588454
rect 83062 588218 83146 588454
rect 83382 588218 118826 588454
rect 119062 588218 119146 588454
rect 119382 588218 154826 588454
rect 155062 588218 155146 588454
rect 155382 588218 190826 588454
rect 191062 588218 191146 588454
rect 191382 588218 226826 588454
rect 227062 588218 227146 588454
rect 227382 588218 262826 588454
rect 263062 588218 263146 588454
rect 263382 588218 298826 588454
rect 299062 588218 299146 588454
rect 299382 588218 334826 588454
rect 335062 588218 335146 588454
rect 335382 588218 370826 588454
rect 371062 588218 371146 588454
rect 371382 588218 406826 588454
rect 407062 588218 407146 588454
rect 407382 588218 442826 588454
rect 443062 588218 443146 588454
rect 443382 588218 478826 588454
rect 479062 588218 479146 588454
rect 479382 588218 514826 588454
rect 515062 588218 515146 588454
rect 515382 588218 550826 588454
rect 551062 588218 551146 588454
rect 551382 588218 587262 588454
rect 587498 588218 587582 588454
rect 587818 588218 592650 588454
rect -8726 588134 592650 588218
rect -8726 587898 -3894 588134
rect -3658 587898 -3574 588134
rect -3338 587898 10826 588134
rect 11062 587898 11146 588134
rect 11382 587898 46826 588134
rect 47062 587898 47146 588134
rect 47382 587898 82826 588134
rect 83062 587898 83146 588134
rect 83382 587898 118826 588134
rect 119062 587898 119146 588134
rect 119382 587898 154826 588134
rect 155062 587898 155146 588134
rect 155382 587898 190826 588134
rect 191062 587898 191146 588134
rect 191382 587898 226826 588134
rect 227062 587898 227146 588134
rect 227382 587898 262826 588134
rect 263062 587898 263146 588134
rect 263382 587898 298826 588134
rect 299062 587898 299146 588134
rect 299382 587898 334826 588134
rect 335062 587898 335146 588134
rect 335382 587898 370826 588134
rect 371062 587898 371146 588134
rect 371382 587898 406826 588134
rect 407062 587898 407146 588134
rect 407382 587898 442826 588134
rect 443062 587898 443146 588134
rect 443382 587898 478826 588134
rect 479062 587898 479146 588134
rect 479382 587898 514826 588134
rect 515062 587898 515146 588134
rect 515382 587898 550826 588134
rect 551062 587898 551146 588134
rect 551382 587898 587262 588134
rect 587498 587898 587582 588134
rect 587818 587898 592650 588134
rect -8726 587866 592650 587898
rect -8726 583954 592650 583986
rect -8726 583718 -2934 583954
rect -2698 583718 -2614 583954
rect -2378 583718 6326 583954
rect 6562 583718 6646 583954
rect 6882 583718 42326 583954
rect 42562 583718 42646 583954
rect 42882 583718 78326 583954
rect 78562 583718 78646 583954
rect 78882 583718 114326 583954
rect 114562 583718 114646 583954
rect 114882 583718 150326 583954
rect 150562 583718 150646 583954
rect 150882 583718 186326 583954
rect 186562 583718 186646 583954
rect 186882 583718 222326 583954
rect 222562 583718 222646 583954
rect 222882 583718 258326 583954
rect 258562 583718 258646 583954
rect 258882 583718 294326 583954
rect 294562 583718 294646 583954
rect 294882 583718 330326 583954
rect 330562 583718 330646 583954
rect 330882 583718 366326 583954
rect 366562 583718 366646 583954
rect 366882 583718 402326 583954
rect 402562 583718 402646 583954
rect 402882 583718 438326 583954
rect 438562 583718 438646 583954
rect 438882 583718 474326 583954
rect 474562 583718 474646 583954
rect 474882 583718 510326 583954
rect 510562 583718 510646 583954
rect 510882 583718 546326 583954
rect 546562 583718 546646 583954
rect 546882 583718 582326 583954
rect 582562 583718 582646 583954
rect 582882 583718 586302 583954
rect 586538 583718 586622 583954
rect 586858 583718 592650 583954
rect -8726 583634 592650 583718
rect -8726 583398 -2934 583634
rect -2698 583398 -2614 583634
rect -2378 583398 6326 583634
rect 6562 583398 6646 583634
rect 6882 583398 42326 583634
rect 42562 583398 42646 583634
rect 42882 583398 78326 583634
rect 78562 583398 78646 583634
rect 78882 583398 114326 583634
rect 114562 583398 114646 583634
rect 114882 583398 150326 583634
rect 150562 583398 150646 583634
rect 150882 583398 186326 583634
rect 186562 583398 186646 583634
rect 186882 583398 222326 583634
rect 222562 583398 222646 583634
rect 222882 583398 258326 583634
rect 258562 583398 258646 583634
rect 258882 583398 294326 583634
rect 294562 583398 294646 583634
rect 294882 583398 330326 583634
rect 330562 583398 330646 583634
rect 330882 583398 366326 583634
rect 366562 583398 366646 583634
rect 366882 583398 402326 583634
rect 402562 583398 402646 583634
rect 402882 583398 438326 583634
rect 438562 583398 438646 583634
rect 438882 583398 474326 583634
rect 474562 583398 474646 583634
rect 474882 583398 510326 583634
rect 510562 583398 510646 583634
rect 510882 583398 546326 583634
rect 546562 583398 546646 583634
rect 546882 583398 582326 583634
rect 582562 583398 582646 583634
rect 582882 583398 586302 583634
rect 586538 583398 586622 583634
rect 586858 583398 592650 583634
rect -8726 583366 592650 583398
rect -8726 579454 592650 579486
rect -8726 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 73826 579454
rect 74062 579218 74146 579454
rect 74382 579218 109826 579454
rect 110062 579218 110146 579454
rect 110382 579218 145826 579454
rect 146062 579218 146146 579454
rect 146382 579218 181826 579454
rect 182062 579218 182146 579454
rect 182382 579218 217826 579454
rect 218062 579218 218146 579454
rect 218382 579218 253826 579454
rect 254062 579218 254146 579454
rect 254382 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 325826 579454
rect 326062 579218 326146 579454
rect 326382 579218 361826 579454
rect 362062 579218 362146 579454
rect 362382 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 592650 579454
rect -8726 579134 592650 579218
rect -8726 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 73826 579134
rect 74062 578898 74146 579134
rect 74382 578898 109826 579134
rect 110062 578898 110146 579134
rect 110382 578898 145826 579134
rect 146062 578898 146146 579134
rect 146382 578898 181826 579134
rect 182062 578898 182146 579134
rect 182382 578898 217826 579134
rect 218062 578898 218146 579134
rect 218382 578898 253826 579134
rect 254062 578898 254146 579134
rect 254382 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 325826 579134
rect 326062 578898 326146 579134
rect 326382 578898 361826 579134
rect 362062 578898 362146 579134
rect 362382 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 592650 579134
rect -8726 578866 592650 578898
rect -8726 574954 592650 574986
rect -8726 574718 -8694 574954
rect -8458 574718 -8374 574954
rect -8138 574718 33326 574954
rect 33562 574718 33646 574954
rect 33882 574718 69326 574954
rect 69562 574718 69646 574954
rect 69882 574718 105326 574954
rect 105562 574718 105646 574954
rect 105882 574718 141326 574954
rect 141562 574718 141646 574954
rect 141882 574718 177326 574954
rect 177562 574718 177646 574954
rect 177882 574718 213326 574954
rect 213562 574718 213646 574954
rect 213882 574718 249326 574954
rect 249562 574718 249646 574954
rect 249882 574718 285326 574954
rect 285562 574718 285646 574954
rect 285882 574718 321326 574954
rect 321562 574718 321646 574954
rect 321882 574718 357326 574954
rect 357562 574718 357646 574954
rect 357882 574718 393326 574954
rect 393562 574718 393646 574954
rect 393882 574718 429326 574954
rect 429562 574718 429646 574954
rect 429882 574718 465326 574954
rect 465562 574718 465646 574954
rect 465882 574718 501326 574954
rect 501562 574718 501646 574954
rect 501882 574718 537326 574954
rect 537562 574718 537646 574954
rect 537882 574718 573326 574954
rect 573562 574718 573646 574954
rect 573882 574718 592062 574954
rect 592298 574718 592382 574954
rect 592618 574718 592650 574954
rect -8726 574634 592650 574718
rect -8726 574398 -8694 574634
rect -8458 574398 -8374 574634
rect -8138 574398 33326 574634
rect 33562 574398 33646 574634
rect 33882 574398 69326 574634
rect 69562 574398 69646 574634
rect 69882 574398 105326 574634
rect 105562 574398 105646 574634
rect 105882 574398 141326 574634
rect 141562 574398 141646 574634
rect 141882 574398 177326 574634
rect 177562 574398 177646 574634
rect 177882 574398 213326 574634
rect 213562 574398 213646 574634
rect 213882 574398 249326 574634
rect 249562 574398 249646 574634
rect 249882 574398 285326 574634
rect 285562 574398 285646 574634
rect 285882 574398 321326 574634
rect 321562 574398 321646 574634
rect 321882 574398 357326 574634
rect 357562 574398 357646 574634
rect 357882 574398 393326 574634
rect 393562 574398 393646 574634
rect 393882 574398 429326 574634
rect 429562 574398 429646 574634
rect 429882 574398 465326 574634
rect 465562 574398 465646 574634
rect 465882 574398 501326 574634
rect 501562 574398 501646 574634
rect 501882 574398 537326 574634
rect 537562 574398 537646 574634
rect 537882 574398 573326 574634
rect 573562 574398 573646 574634
rect 573882 574398 592062 574634
rect 592298 574398 592382 574634
rect 592618 574398 592650 574634
rect -8726 574366 592650 574398
rect -8726 570454 592650 570486
rect -8726 570218 -7734 570454
rect -7498 570218 -7414 570454
rect -7178 570218 28826 570454
rect 29062 570218 29146 570454
rect 29382 570218 64826 570454
rect 65062 570218 65146 570454
rect 65382 570218 100826 570454
rect 101062 570218 101146 570454
rect 101382 570218 136826 570454
rect 137062 570218 137146 570454
rect 137382 570218 172826 570454
rect 173062 570218 173146 570454
rect 173382 570218 208826 570454
rect 209062 570218 209146 570454
rect 209382 570218 244826 570454
rect 245062 570218 245146 570454
rect 245382 570218 280826 570454
rect 281062 570218 281146 570454
rect 281382 570218 316826 570454
rect 317062 570218 317146 570454
rect 317382 570218 352826 570454
rect 353062 570218 353146 570454
rect 353382 570218 388826 570454
rect 389062 570218 389146 570454
rect 389382 570218 424826 570454
rect 425062 570218 425146 570454
rect 425382 570218 460826 570454
rect 461062 570218 461146 570454
rect 461382 570218 496826 570454
rect 497062 570218 497146 570454
rect 497382 570218 532826 570454
rect 533062 570218 533146 570454
rect 533382 570218 568826 570454
rect 569062 570218 569146 570454
rect 569382 570218 591102 570454
rect 591338 570218 591422 570454
rect 591658 570218 592650 570454
rect -8726 570134 592650 570218
rect -8726 569898 -7734 570134
rect -7498 569898 -7414 570134
rect -7178 569898 28826 570134
rect 29062 569898 29146 570134
rect 29382 569898 64826 570134
rect 65062 569898 65146 570134
rect 65382 569898 100826 570134
rect 101062 569898 101146 570134
rect 101382 569898 136826 570134
rect 137062 569898 137146 570134
rect 137382 569898 172826 570134
rect 173062 569898 173146 570134
rect 173382 569898 208826 570134
rect 209062 569898 209146 570134
rect 209382 569898 244826 570134
rect 245062 569898 245146 570134
rect 245382 569898 280826 570134
rect 281062 569898 281146 570134
rect 281382 569898 316826 570134
rect 317062 569898 317146 570134
rect 317382 569898 352826 570134
rect 353062 569898 353146 570134
rect 353382 569898 388826 570134
rect 389062 569898 389146 570134
rect 389382 569898 424826 570134
rect 425062 569898 425146 570134
rect 425382 569898 460826 570134
rect 461062 569898 461146 570134
rect 461382 569898 496826 570134
rect 497062 569898 497146 570134
rect 497382 569898 532826 570134
rect 533062 569898 533146 570134
rect 533382 569898 568826 570134
rect 569062 569898 569146 570134
rect 569382 569898 591102 570134
rect 591338 569898 591422 570134
rect 591658 569898 592650 570134
rect -8726 569866 592650 569898
rect -8726 565954 592650 565986
rect -8726 565718 -6774 565954
rect -6538 565718 -6454 565954
rect -6218 565718 24326 565954
rect 24562 565718 24646 565954
rect 24882 565718 60326 565954
rect 60562 565718 60646 565954
rect 60882 565718 96326 565954
rect 96562 565718 96646 565954
rect 96882 565718 132326 565954
rect 132562 565718 132646 565954
rect 132882 565718 168326 565954
rect 168562 565718 168646 565954
rect 168882 565718 204326 565954
rect 204562 565718 204646 565954
rect 204882 565718 240326 565954
rect 240562 565718 240646 565954
rect 240882 565718 276326 565954
rect 276562 565718 276646 565954
rect 276882 565718 312326 565954
rect 312562 565718 312646 565954
rect 312882 565718 348326 565954
rect 348562 565718 348646 565954
rect 348882 565718 384326 565954
rect 384562 565718 384646 565954
rect 384882 565718 420326 565954
rect 420562 565718 420646 565954
rect 420882 565718 456326 565954
rect 456562 565718 456646 565954
rect 456882 565718 492326 565954
rect 492562 565718 492646 565954
rect 492882 565718 528326 565954
rect 528562 565718 528646 565954
rect 528882 565718 564326 565954
rect 564562 565718 564646 565954
rect 564882 565718 590142 565954
rect 590378 565718 590462 565954
rect 590698 565718 592650 565954
rect -8726 565634 592650 565718
rect -8726 565398 -6774 565634
rect -6538 565398 -6454 565634
rect -6218 565398 24326 565634
rect 24562 565398 24646 565634
rect 24882 565398 60326 565634
rect 60562 565398 60646 565634
rect 60882 565398 96326 565634
rect 96562 565398 96646 565634
rect 96882 565398 132326 565634
rect 132562 565398 132646 565634
rect 132882 565398 168326 565634
rect 168562 565398 168646 565634
rect 168882 565398 204326 565634
rect 204562 565398 204646 565634
rect 204882 565398 240326 565634
rect 240562 565398 240646 565634
rect 240882 565398 276326 565634
rect 276562 565398 276646 565634
rect 276882 565398 312326 565634
rect 312562 565398 312646 565634
rect 312882 565398 348326 565634
rect 348562 565398 348646 565634
rect 348882 565398 384326 565634
rect 384562 565398 384646 565634
rect 384882 565398 420326 565634
rect 420562 565398 420646 565634
rect 420882 565398 456326 565634
rect 456562 565398 456646 565634
rect 456882 565398 492326 565634
rect 492562 565398 492646 565634
rect 492882 565398 528326 565634
rect 528562 565398 528646 565634
rect 528882 565398 564326 565634
rect 564562 565398 564646 565634
rect 564882 565398 590142 565634
rect 590378 565398 590462 565634
rect 590698 565398 592650 565634
rect -8726 565366 592650 565398
rect -8726 561454 592650 561486
rect -8726 561218 -5814 561454
rect -5578 561218 -5494 561454
rect -5258 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 55826 561454
rect 56062 561218 56146 561454
rect 56382 561218 91826 561454
rect 92062 561218 92146 561454
rect 92382 561218 127826 561454
rect 128062 561218 128146 561454
rect 128382 561218 163826 561454
rect 164062 561218 164146 561454
rect 164382 561218 199826 561454
rect 200062 561218 200146 561454
rect 200382 561218 235826 561454
rect 236062 561218 236146 561454
rect 236382 561218 271826 561454
rect 272062 561218 272146 561454
rect 272382 561218 307826 561454
rect 308062 561218 308146 561454
rect 308382 561218 343826 561454
rect 344062 561218 344146 561454
rect 344382 561218 379826 561454
rect 380062 561218 380146 561454
rect 380382 561218 415826 561454
rect 416062 561218 416146 561454
rect 416382 561218 451826 561454
rect 452062 561218 452146 561454
rect 452382 561218 487826 561454
rect 488062 561218 488146 561454
rect 488382 561218 523826 561454
rect 524062 561218 524146 561454
rect 524382 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 589182 561454
rect 589418 561218 589502 561454
rect 589738 561218 592650 561454
rect -8726 561134 592650 561218
rect -8726 560898 -5814 561134
rect -5578 560898 -5494 561134
rect -5258 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 55826 561134
rect 56062 560898 56146 561134
rect 56382 560898 91826 561134
rect 92062 560898 92146 561134
rect 92382 560898 127826 561134
rect 128062 560898 128146 561134
rect 128382 560898 163826 561134
rect 164062 560898 164146 561134
rect 164382 560898 199826 561134
rect 200062 560898 200146 561134
rect 200382 560898 235826 561134
rect 236062 560898 236146 561134
rect 236382 560898 271826 561134
rect 272062 560898 272146 561134
rect 272382 560898 307826 561134
rect 308062 560898 308146 561134
rect 308382 560898 343826 561134
rect 344062 560898 344146 561134
rect 344382 560898 379826 561134
rect 380062 560898 380146 561134
rect 380382 560898 415826 561134
rect 416062 560898 416146 561134
rect 416382 560898 451826 561134
rect 452062 560898 452146 561134
rect 452382 560898 487826 561134
rect 488062 560898 488146 561134
rect 488382 560898 523826 561134
rect 524062 560898 524146 561134
rect 524382 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 589182 561134
rect 589418 560898 589502 561134
rect 589738 560898 592650 561134
rect -8726 560866 592650 560898
rect -8726 556954 592650 556986
rect -8726 556718 -4854 556954
rect -4618 556718 -4534 556954
rect -4298 556718 15326 556954
rect 15562 556718 15646 556954
rect 15882 556718 51326 556954
rect 51562 556718 51646 556954
rect 51882 556718 87326 556954
rect 87562 556718 87646 556954
rect 87882 556718 123326 556954
rect 123562 556718 123646 556954
rect 123882 556718 159326 556954
rect 159562 556718 159646 556954
rect 159882 556718 195326 556954
rect 195562 556718 195646 556954
rect 195882 556718 231326 556954
rect 231562 556718 231646 556954
rect 231882 556718 267326 556954
rect 267562 556718 267646 556954
rect 267882 556718 303326 556954
rect 303562 556718 303646 556954
rect 303882 556718 339326 556954
rect 339562 556718 339646 556954
rect 339882 556718 375326 556954
rect 375562 556718 375646 556954
rect 375882 556718 411326 556954
rect 411562 556718 411646 556954
rect 411882 556718 447326 556954
rect 447562 556718 447646 556954
rect 447882 556718 483326 556954
rect 483562 556718 483646 556954
rect 483882 556718 519326 556954
rect 519562 556718 519646 556954
rect 519882 556718 555326 556954
rect 555562 556718 555646 556954
rect 555882 556718 588222 556954
rect 588458 556718 588542 556954
rect 588778 556718 592650 556954
rect -8726 556634 592650 556718
rect -8726 556398 -4854 556634
rect -4618 556398 -4534 556634
rect -4298 556398 15326 556634
rect 15562 556398 15646 556634
rect 15882 556398 51326 556634
rect 51562 556398 51646 556634
rect 51882 556398 87326 556634
rect 87562 556398 87646 556634
rect 87882 556398 123326 556634
rect 123562 556398 123646 556634
rect 123882 556398 159326 556634
rect 159562 556398 159646 556634
rect 159882 556398 195326 556634
rect 195562 556398 195646 556634
rect 195882 556398 231326 556634
rect 231562 556398 231646 556634
rect 231882 556398 267326 556634
rect 267562 556398 267646 556634
rect 267882 556398 303326 556634
rect 303562 556398 303646 556634
rect 303882 556398 339326 556634
rect 339562 556398 339646 556634
rect 339882 556398 375326 556634
rect 375562 556398 375646 556634
rect 375882 556398 411326 556634
rect 411562 556398 411646 556634
rect 411882 556398 447326 556634
rect 447562 556398 447646 556634
rect 447882 556398 483326 556634
rect 483562 556398 483646 556634
rect 483882 556398 519326 556634
rect 519562 556398 519646 556634
rect 519882 556398 555326 556634
rect 555562 556398 555646 556634
rect 555882 556398 588222 556634
rect 588458 556398 588542 556634
rect 588778 556398 592650 556634
rect -8726 556366 592650 556398
rect -8726 552454 592650 552486
rect -8726 552218 -3894 552454
rect -3658 552218 -3574 552454
rect -3338 552218 10826 552454
rect 11062 552218 11146 552454
rect 11382 552218 46826 552454
rect 47062 552218 47146 552454
rect 47382 552218 82826 552454
rect 83062 552218 83146 552454
rect 83382 552218 118826 552454
rect 119062 552218 119146 552454
rect 119382 552218 154826 552454
rect 155062 552218 155146 552454
rect 155382 552218 190826 552454
rect 191062 552218 191146 552454
rect 191382 552218 226826 552454
rect 227062 552218 227146 552454
rect 227382 552218 262826 552454
rect 263062 552218 263146 552454
rect 263382 552218 298826 552454
rect 299062 552218 299146 552454
rect 299382 552218 334826 552454
rect 335062 552218 335146 552454
rect 335382 552218 370826 552454
rect 371062 552218 371146 552454
rect 371382 552218 406826 552454
rect 407062 552218 407146 552454
rect 407382 552218 442826 552454
rect 443062 552218 443146 552454
rect 443382 552218 478826 552454
rect 479062 552218 479146 552454
rect 479382 552218 514826 552454
rect 515062 552218 515146 552454
rect 515382 552218 550826 552454
rect 551062 552218 551146 552454
rect 551382 552218 587262 552454
rect 587498 552218 587582 552454
rect 587818 552218 592650 552454
rect -8726 552134 592650 552218
rect -8726 551898 -3894 552134
rect -3658 551898 -3574 552134
rect -3338 551898 10826 552134
rect 11062 551898 11146 552134
rect 11382 551898 46826 552134
rect 47062 551898 47146 552134
rect 47382 551898 82826 552134
rect 83062 551898 83146 552134
rect 83382 551898 118826 552134
rect 119062 551898 119146 552134
rect 119382 551898 154826 552134
rect 155062 551898 155146 552134
rect 155382 551898 190826 552134
rect 191062 551898 191146 552134
rect 191382 551898 226826 552134
rect 227062 551898 227146 552134
rect 227382 551898 262826 552134
rect 263062 551898 263146 552134
rect 263382 551898 298826 552134
rect 299062 551898 299146 552134
rect 299382 551898 334826 552134
rect 335062 551898 335146 552134
rect 335382 551898 370826 552134
rect 371062 551898 371146 552134
rect 371382 551898 406826 552134
rect 407062 551898 407146 552134
rect 407382 551898 442826 552134
rect 443062 551898 443146 552134
rect 443382 551898 478826 552134
rect 479062 551898 479146 552134
rect 479382 551898 514826 552134
rect 515062 551898 515146 552134
rect 515382 551898 550826 552134
rect 551062 551898 551146 552134
rect 551382 551898 587262 552134
rect 587498 551898 587582 552134
rect 587818 551898 592650 552134
rect -8726 551866 592650 551898
rect -8726 547954 592650 547986
rect -8726 547718 -2934 547954
rect -2698 547718 -2614 547954
rect -2378 547718 6326 547954
rect 6562 547718 6646 547954
rect 6882 547718 42326 547954
rect 42562 547718 42646 547954
rect 42882 547718 78326 547954
rect 78562 547718 78646 547954
rect 78882 547718 114326 547954
rect 114562 547718 114646 547954
rect 114882 547718 150326 547954
rect 150562 547718 150646 547954
rect 150882 547718 186326 547954
rect 186562 547718 186646 547954
rect 186882 547718 222326 547954
rect 222562 547718 222646 547954
rect 222882 547718 258326 547954
rect 258562 547718 258646 547954
rect 258882 547718 294326 547954
rect 294562 547718 294646 547954
rect 294882 547718 330326 547954
rect 330562 547718 330646 547954
rect 330882 547718 366326 547954
rect 366562 547718 366646 547954
rect 366882 547718 402326 547954
rect 402562 547718 402646 547954
rect 402882 547718 438326 547954
rect 438562 547718 438646 547954
rect 438882 547718 474326 547954
rect 474562 547718 474646 547954
rect 474882 547718 510326 547954
rect 510562 547718 510646 547954
rect 510882 547718 546326 547954
rect 546562 547718 546646 547954
rect 546882 547718 582326 547954
rect 582562 547718 582646 547954
rect 582882 547718 586302 547954
rect 586538 547718 586622 547954
rect 586858 547718 592650 547954
rect -8726 547634 592650 547718
rect -8726 547398 -2934 547634
rect -2698 547398 -2614 547634
rect -2378 547398 6326 547634
rect 6562 547398 6646 547634
rect 6882 547398 42326 547634
rect 42562 547398 42646 547634
rect 42882 547398 78326 547634
rect 78562 547398 78646 547634
rect 78882 547398 114326 547634
rect 114562 547398 114646 547634
rect 114882 547398 150326 547634
rect 150562 547398 150646 547634
rect 150882 547398 186326 547634
rect 186562 547398 186646 547634
rect 186882 547398 222326 547634
rect 222562 547398 222646 547634
rect 222882 547398 258326 547634
rect 258562 547398 258646 547634
rect 258882 547398 294326 547634
rect 294562 547398 294646 547634
rect 294882 547398 330326 547634
rect 330562 547398 330646 547634
rect 330882 547398 366326 547634
rect 366562 547398 366646 547634
rect 366882 547398 402326 547634
rect 402562 547398 402646 547634
rect 402882 547398 438326 547634
rect 438562 547398 438646 547634
rect 438882 547398 474326 547634
rect 474562 547398 474646 547634
rect 474882 547398 510326 547634
rect 510562 547398 510646 547634
rect 510882 547398 546326 547634
rect 546562 547398 546646 547634
rect 546882 547398 582326 547634
rect 582562 547398 582646 547634
rect 582882 547398 586302 547634
rect 586538 547398 586622 547634
rect 586858 547398 592650 547634
rect -8726 547366 592650 547398
rect -8726 543454 592650 543486
rect -8726 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 73826 543454
rect 74062 543218 74146 543454
rect 74382 543218 109826 543454
rect 110062 543218 110146 543454
rect 110382 543218 145826 543454
rect 146062 543218 146146 543454
rect 146382 543218 181826 543454
rect 182062 543218 182146 543454
rect 182382 543218 217826 543454
rect 218062 543218 218146 543454
rect 218382 543218 253826 543454
rect 254062 543218 254146 543454
rect 254382 543218 289826 543454
rect 290062 543218 290146 543454
rect 290382 543218 325826 543454
rect 326062 543218 326146 543454
rect 326382 543218 361826 543454
rect 362062 543218 362146 543454
rect 362382 543218 397826 543454
rect 398062 543218 398146 543454
rect 398382 543218 433826 543454
rect 434062 543218 434146 543454
rect 434382 543218 469826 543454
rect 470062 543218 470146 543454
rect 470382 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 592650 543454
rect -8726 543134 592650 543218
rect -8726 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 73826 543134
rect 74062 542898 74146 543134
rect 74382 542898 109826 543134
rect 110062 542898 110146 543134
rect 110382 542898 145826 543134
rect 146062 542898 146146 543134
rect 146382 542898 181826 543134
rect 182062 542898 182146 543134
rect 182382 542898 217826 543134
rect 218062 542898 218146 543134
rect 218382 542898 253826 543134
rect 254062 542898 254146 543134
rect 254382 542898 289826 543134
rect 290062 542898 290146 543134
rect 290382 542898 325826 543134
rect 326062 542898 326146 543134
rect 326382 542898 361826 543134
rect 362062 542898 362146 543134
rect 362382 542898 397826 543134
rect 398062 542898 398146 543134
rect 398382 542898 433826 543134
rect 434062 542898 434146 543134
rect 434382 542898 469826 543134
rect 470062 542898 470146 543134
rect 470382 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 592650 543134
rect -8726 542866 592650 542898
rect -8726 538954 592650 538986
rect -8726 538718 -8694 538954
rect -8458 538718 -8374 538954
rect -8138 538718 33326 538954
rect 33562 538718 33646 538954
rect 33882 538718 69326 538954
rect 69562 538718 69646 538954
rect 69882 538718 105326 538954
rect 105562 538718 105646 538954
rect 105882 538718 141326 538954
rect 141562 538718 141646 538954
rect 141882 538718 177326 538954
rect 177562 538718 177646 538954
rect 177882 538718 213326 538954
rect 213562 538718 213646 538954
rect 213882 538718 249326 538954
rect 249562 538718 249646 538954
rect 249882 538718 285326 538954
rect 285562 538718 285646 538954
rect 285882 538718 321326 538954
rect 321562 538718 321646 538954
rect 321882 538718 357326 538954
rect 357562 538718 357646 538954
rect 357882 538718 393326 538954
rect 393562 538718 393646 538954
rect 393882 538718 429326 538954
rect 429562 538718 429646 538954
rect 429882 538718 465326 538954
rect 465562 538718 465646 538954
rect 465882 538718 501326 538954
rect 501562 538718 501646 538954
rect 501882 538718 537326 538954
rect 537562 538718 537646 538954
rect 537882 538718 573326 538954
rect 573562 538718 573646 538954
rect 573882 538718 592062 538954
rect 592298 538718 592382 538954
rect 592618 538718 592650 538954
rect -8726 538634 592650 538718
rect -8726 538398 -8694 538634
rect -8458 538398 -8374 538634
rect -8138 538398 33326 538634
rect 33562 538398 33646 538634
rect 33882 538398 69326 538634
rect 69562 538398 69646 538634
rect 69882 538398 105326 538634
rect 105562 538398 105646 538634
rect 105882 538398 141326 538634
rect 141562 538398 141646 538634
rect 141882 538398 177326 538634
rect 177562 538398 177646 538634
rect 177882 538398 213326 538634
rect 213562 538398 213646 538634
rect 213882 538398 249326 538634
rect 249562 538398 249646 538634
rect 249882 538398 285326 538634
rect 285562 538398 285646 538634
rect 285882 538398 321326 538634
rect 321562 538398 321646 538634
rect 321882 538398 357326 538634
rect 357562 538398 357646 538634
rect 357882 538398 393326 538634
rect 393562 538398 393646 538634
rect 393882 538398 429326 538634
rect 429562 538398 429646 538634
rect 429882 538398 465326 538634
rect 465562 538398 465646 538634
rect 465882 538398 501326 538634
rect 501562 538398 501646 538634
rect 501882 538398 537326 538634
rect 537562 538398 537646 538634
rect 537882 538398 573326 538634
rect 573562 538398 573646 538634
rect 573882 538398 592062 538634
rect 592298 538398 592382 538634
rect 592618 538398 592650 538634
rect -8726 538366 592650 538398
rect -8726 534454 592650 534486
rect -8726 534218 -7734 534454
rect -7498 534218 -7414 534454
rect -7178 534218 28826 534454
rect 29062 534218 29146 534454
rect 29382 534218 64826 534454
rect 65062 534218 65146 534454
rect 65382 534218 100826 534454
rect 101062 534218 101146 534454
rect 101382 534218 136826 534454
rect 137062 534218 137146 534454
rect 137382 534218 172826 534454
rect 173062 534218 173146 534454
rect 173382 534218 208826 534454
rect 209062 534218 209146 534454
rect 209382 534218 244826 534454
rect 245062 534218 245146 534454
rect 245382 534218 280826 534454
rect 281062 534218 281146 534454
rect 281382 534218 316826 534454
rect 317062 534218 317146 534454
rect 317382 534218 352826 534454
rect 353062 534218 353146 534454
rect 353382 534218 388826 534454
rect 389062 534218 389146 534454
rect 389382 534218 424826 534454
rect 425062 534218 425146 534454
rect 425382 534218 460826 534454
rect 461062 534218 461146 534454
rect 461382 534218 496826 534454
rect 497062 534218 497146 534454
rect 497382 534218 532826 534454
rect 533062 534218 533146 534454
rect 533382 534218 568826 534454
rect 569062 534218 569146 534454
rect 569382 534218 591102 534454
rect 591338 534218 591422 534454
rect 591658 534218 592650 534454
rect -8726 534134 592650 534218
rect -8726 533898 -7734 534134
rect -7498 533898 -7414 534134
rect -7178 533898 28826 534134
rect 29062 533898 29146 534134
rect 29382 533898 64826 534134
rect 65062 533898 65146 534134
rect 65382 533898 100826 534134
rect 101062 533898 101146 534134
rect 101382 533898 136826 534134
rect 137062 533898 137146 534134
rect 137382 533898 172826 534134
rect 173062 533898 173146 534134
rect 173382 533898 208826 534134
rect 209062 533898 209146 534134
rect 209382 533898 244826 534134
rect 245062 533898 245146 534134
rect 245382 533898 280826 534134
rect 281062 533898 281146 534134
rect 281382 533898 316826 534134
rect 317062 533898 317146 534134
rect 317382 533898 352826 534134
rect 353062 533898 353146 534134
rect 353382 533898 388826 534134
rect 389062 533898 389146 534134
rect 389382 533898 424826 534134
rect 425062 533898 425146 534134
rect 425382 533898 460826 534134
rect 461062 533898 461146 534134
rect 461382 533898 496826 534134
rect 497062 533898 497146 534134
rect 497382 533898 532826 534134
rect 533062 533898 533146 534134
rect 533382 533898 568826 534134
rect 569062 533898 569146 534134
rect 569382 533898 591102 534134
rect 591338 533898 591422 534134
rect 591658 533898 592650 534134
rect -8726 533866 592650 533898
rect -8726 529954 592650 529986
rect -8726 529718 -6774 529954
rect -6538 529718 -6454 529954
rect -6218 529718 24326 529954
rect 24562 529718 24646 529954
rect 24882 529718 60326 529954
rect 60562 529718 60646 529954
rect 60882 529718 96326 529954
rect 96562 529718 96646 529954
rect 96882 529718 132326 529954
rect 132562 529718 132646 529954
rect 132882 529718 168326 529954
rect 168562 529718 168646 529954
rect 168882 529718 204326 529954
rect 204562 529718 204646 529954
rect 204882 529718 240326 529954
rect 240562 529718 240646 529954
rect 240882 529718 276326 529954
rect 276562 529718 276646 529954
rect 276882 529718 312326 529954
rect 312562 529718 312646 529954
rect 312882 529718 348326 529954
rect 348562 529718 348646 529954
rect 348882 529718 384326 529954
rect 384562 529718 384646 529954
rect 384882 529718 420326 529954
rect 420562 529718 420646 529954
rect 420882 529718 456326 529954
rect 456562 529718 456646 529954
rect 456882 529718 492326 529954
rect 492562 529718 492646 529954
rect 492882 529718 528326 529954
rect 528562 529718 528646 529954
rect 528882 529718 564326 529954
rect 564562 529718 564646 529954
rect 564882 529718 590142 529954
rect 590378 529718 590462 529954
rect 590698 529718 592650 529954
rect -8726 529634 592650 529718
rect -8726 529398 -6774 529634
rect -6538 529398 -6454 529634
rect -6218 529398 24326 529634
rect 24562 529398 24646 529634
rect 24882 529398 60326 529634
rect 60562 529398 60646 529634
rect 60882 529398 96326 529634
rect 96562 529398 96646 529634
rect 96882 529398 132326 529634
rect 132562 529398 132646 529634
rect 132882 529398 168326 529634
rect 168562 529398 168646 529634
rect 168882 529398 204326 529634
rect 204562 529398 204646 529634
rect 204882 529398 240326 529634
rect 240562 529398 240646 529634
rect 240882 529398 276326 529634
rect 276562 529398 276646 529634
rect 276882 529398 312326 529634
rect 312562 529398 312646 529634
rect 312882 529398 348326 529634
rect 348562 529398 348646 529634
rect 348882 529398 384326 529634
rect 384562 529398 384646 529634
rect 384882 529398 420326 529634
rect 420562 529398 420646 529634
rect 420882 529398 456326 529634
rect 456562 529398 456646 529634
rect 456882 529398 492326 529634
rect 492562 529398 492646 529634
rect 492882 529398 528326 529634
rect 528562 529398 528646 529634
rect 528882 529398 564326 529634
rect 564562 529398 564646 529634
rect 564882 529398 590142 529634
rect 590378 529398 590462 529634
rect 590698 529398 592650 529634
rect -8726 529366 592650 529398
rect -8726 525454 592650 525486
rect -8726 525218 -5814 525454
rect -5578 525218 -5494 525454
rect -5258 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 55826 525454
rect 56062 525218 56146 525454
rect 56382 525218 91826 525454
rect 92062 525218 92146 525454
rect 92382 525218 127826 525454
rect 128062 525218 128146 525454
rect 128382 525218 163826 525454
rect 164062 525218 164146 525454
rect 164382 525218 199826 525454
rect 200062 525218 200146 525454
rect 200382 525218 235826 525454
rect 236062 525218 236146 525454
rect 236382 525218 271826 525454
rect 272062 525218 272146 525454
rect 272382 525218 307826 525454
rect 308062 525218 308146 525454
rect 308382 525218 343826 525454
rect 344062 525218 344146 525454
rect 344382 525218 379826 525454
rect 380062 525218 380146 525454
rect 380382 525218 415826 525454
rect 416062 525218 416146 525454
rect 416382 525218 451826 525454
rect 452062 525218 452146 525454
rect 452382 525218 487826 525454
rect 488062 525218 488146 525454
rect 488382 525218 523826 525454
rect 524062 525218 524146 525454
rect 524382 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 589182 525454
rect 589418 525218 589502 525454
rect 589738 525218 592650 525454
rect -8726 525134 592650 525218
rect -8726 524898 -5814 525134
rect -5578 524898 -5494 525134
rect -5258 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 55826 525134
rect 56062 524898 56146 525134
rect 56382 524898 91826 525134
rect 92062 524898 92146 525134
rect 92382 524898 127826 525134
rect 128062 524898 128146 525134
rect 128382 524898 163826 525134
rect 164062 524898 164146 525134
rect 164382 524898 199826 525134
rect 200062 524898 200146 525134
rect 200382 524898 235826 525134
rect 236062 524898 236146 525134
rect 236382 524898 271826 525134
rect 272062 524898 272146 525134
rect 272382 524898 307826 525134
rect 308062 524898 308146 525134
rect 308382 524898 343826 525134
rect 344062 524898 344146 525134
rect 344382 524898 379826 525134
rect 380062 524898 380146 525134
rect 380382 524898 415826 525134
rect 416062 524898 416146 525134
rect 416382 524898 451826 525134
rect 452062 524898 452146 525134
rect 452382 524898 487826 525134
rect 488062 524898 488146 525134
rect 488382 524898 523826 525134
rect 524062 524898 524146 525134
rect 524382 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 589182 525134
rect 589418 524898 589502 525134
rect 589738 524898 592650 525134
rect -8726 524866 592650 524898
rect -8726 520954 592650 520986
rect -8726 520718 -4854 520954
rect -4618 520718 -4534 520954
rect -4298 520718 15326 520954
rect 15562 520718 15646 520954
rect 15882 520718 51326 520954
rect 51562 520718 51646 520954
rect 51882 520718 87326 520954
rect 87562 520718 87646 520954
rect 87882 520718 123326 520954
rect 123562 520718 123646 520954
rect 123882 520718 159326 520954
rect 159562 520718 159646 520954
rect 159882 520718 195326 520954
rect 195562 520718 195646 520954
rect 195882 520718 231326 520954
rect 231562 520718 231646 520954
rect 231882 520718 267326 520954
rect 267562 520718 267646 520954
rect 267882 520718 303326 520954
rect 303562 520718 303646 520954
rect 303882 520718 339326 520954
rect 339562 520718 339646 520954
rect 339882 520718 375326 520954
rect 375562 520718 375646 520954
rect 375882 520718 411326 520954
rect 411562 520718 411646 520954
rect 411882 520718 447326 520954
rect 447562 520718 447646 520954
rect 447882 520718 483326 520954
rect 483562 520718 483646 520954
rect 483882 520718 519326 520954
rect 519562 520718 519646 520954
rect 519882 520718 555326 520954
rect 555562 520718 555646 520954
rect 555882 520718 588222 520954
rect 588458 520718 588542 520954
rect 588778 520718 592650 520954
rect -8726 520634 592650 520718
rect -8726 520398 -4854 520634
rect -4618 520398 -4534 520634
rect -4298 520398 15326 520634
rect 15562 520398 15646 520634
rect 15882 520398 51326 520634
rect 51562 520398 51646 520634
rect 51882 520398 87326 520634
rect 87562 520398 87646 520634
rect 87882 520398 123326 520634
rect 123562 520398 123646 520634
rect 123882 520398 159326 520634
rect 159562 520398 159646 520634
rect 159882 520398 195326 520634
rect 195562 520398 195646 520634
rect 195882 520398 231326 520634
rect 231562 520398 231646 520634
rect 231882 520398 267326 520634
rect 267562 520398 267646 520634
rect 267882 520398 303326 520634
rect 303562 520398 303646 520634
rect 303882 520398 339326 520634
rect 339562 520398 339646 520634
rect 339882 520398 375326 520634
rect 375562 520398 375646 520634
rect 375882 520398 411326 520634
rect 411562 520398 411646 520634
rect 411882 520398 447326 520634
rect 447562 520398 447646 520634
rect 447882 520398 483326 520634
rect 483562 520398 483646 520634
rect 483882 520398 519326 520634
rect 519562 520398 519646 520634
rect 519882 520398 555326 520634
rect 555562 520398 555646 520634
rect 555882 520398 588222 520634
rect 588458 520398 588542 520634
rect 588778 520398 592650 520634
rect -8726 520366 592650 520398
rect -8726 516454 592650 516486
rect -8726 516218 -3894 516454
rect -3658 516218 -3574 516454
rect -3338 516218 10826 516454
rect 11062 516218 11146 516454
rect 11382 516218 46826 516454
rect 47062 516218 47146 516454
rect 47382 516218 82826 516454
rect 83062 516218 83146 516454
rect 83382 516218 118826 516454
rect 119062 516218 119146 516454
rect 119382 516218 154826 516454
rect 155062 516218 155146 516454
rect 155382 516218 190826 516454
rect 191062 516218 191146 516454
rect 191382 516218 226826 516454
rect 227062 516218 227146 516454
rect 227382 516218 262826 516454
rect 263062 516218 263146 516454
rect 263382 516218 298826 516454
rect 299062 516218 299146 516454
rect 299382 516218 334826 516454
rect 335062 516218 335146 516454
rect 335382 516218 370826 516454
rect 371062 516218 371146 516454
rect 371382 516218 406826 516454
rect 407062 516218 407146 516454
rect 407382 516218 442826 516454
rect 443062 516218 443146 516454
rect 443382 516218 478826 516454
rect 479062 516218 479146 516454
rect 479382 516218 514826 516454
rect 515062 516218 515146 516454
rect 515382 516218 550826 516454
rect 551062 516218 551146 516454
rect 551382 516218 587262 516454
rect 587498 516218 587582 516454
rect 587818 516218 592650 516454
rect -8726 516134 592650 516218
rect -8726 515898 -3894 516134
rect -3658 515898 -3574 516134
rect -3338 515898 10826 516134
rect 11062 515898 11146 516134
rect 11382 515898 46826 516134
rect 47062 515898 47146 516134
rect 47382 515898 82826 516134
rect 83062 515898 83146 516134
rect 83382 515898 118826 516134
rect 119062 515898 119146 516134
rect 119382 515898 154826 516134
rect 155062 515898 155146 516134
rect 155382 515898 190826 516134
rect 191062 515898 191146 516134
rect 191382 515898 226826 516134
rect 227062 515898 227146 516134
rect 227382 515898 262826 516134
rect 263062 515898 263146 516134
rect 263382 515898 298826 516134
rect 299062 515898 299146 516134
rect 299382 515898 334826 516134
rect 335062 515898 335146 516134
rect 335382 515898 370826 516134
rect 371062 515898 371146 516134
rect 371382 515898 406826 516134
rect 407062 515898 407146 516134
rect 407382 515898 442826 516134
rect 443062 515898 443146 516134
rect 443382 515898 478826 516134
rect 479062 515898 479146 516134
rect 479382 515898 514826 516134
rect 515062 515898 515146 516134
rect 515382 515898 550826 516134
rect 551062 515898 551146 516134
rect 551382 515898 587262 516134
rect 587498 515898 587582 516134
rect 587818 515898 592650 516134
rect -8726 515866 592650 515898
rect -8726 511954 592650 511986
rect -8726 511718 -2934 511954
rect -2698 511718 -2614 511954
rect -2378 511718 6326 511954
rect 6562 511718 6646 511954
rect 6882 511718 42326 511954
rect 42562 511718 42646 511954
rect 42882 511718 78326 511954
rect 78562 511718 78646 511954
rect 78882 511718 114326 511954
rect 114562 511718 114646 511954
rect 114882 511718 150326 511954
rect 150562 511718 150646 511954
rect 150882 511718 186326 511954
rect 186562 511718 186646 511954
rect 186882 511718 222326 511954
rect 222562 511718 222646 511954
rect 222882 511718 258326 511954
rect 258562 511718 258646 511954
rect 258882 511718 294326 511954
rect 294562 511718 294646 511954
rect 294882 511718 330326 511954
rect 330562 511718 330646 511954
rect 330882 511718 366326 511954
rect 366562 511718 366646 511954
rect 366882 511718 402326 511954
rect 402562 511718 402646 511954
rect 402882 511718 438326 511954
rect 438562 511718 438646 511954
rect 438882 511718 474326 511954
rect 474562 511718 474646 511954
rect 474882 511718 510326 511954
rect 510562 511718 510646 511954
rect 510882 511718 546326 511954
rect 546562 511718 546646 511954
rect 546882 511718 582326 511954
rect 582562 511718 582646 511954
rect 582882 511718 586302 511954
rect 586538 511718 586622 511954
rect 586858 511718 592650 511954
rect -8726 511634 592650 511718
rect -8726 511398 -2934 511634
rect -2698 511398 -2614 511634
rect -2378 511398 6326 511634
rect 6562 511398 6646 511634
rect 6882 511398 42326 511634
rect 42562 511398 42646 511634
rect 42882 511398 78326 511634
rect 78562 511398 78646 511634
rect 78882 511398 114326 511634
rect 114562 511398 114646 511634
rect 114882 511398 150326 511634
rect 150562 511398 150646 511634
rect 150882 511398 186326 511634
rect 186562 511398 186646 511634
rect 186882 511398 222326 511634
rect 222562 511398 222646 511634
rect 222882 511398 258326 511634
rect 258562 511398 258646 511634
rect 258882 511398 294326 511634
rect 294562 511398 294646 511634
rect 294882 511398 330326 511634
rect 330562 511398 330646 511634
rect 330882 511398 366326 511634
rect 366562 511398 366646 511634
rect 366882 511398 402326 511634
rect 402562 511398 402646 511634
rect 402882 511398 438326 511634
rect 438562 511398 438646 511634
rect 438882 511398 474326 511634
rect 474562 511398 474646 511634
rect 474882 511398 510326 511634
rect 510562 511398 510646 511634
rect 510882 511398 546326 511634
rect 546562 511398 546646 511634
rect 546882 511398 582326 511634
rect 582562 511398 582646 511634
rect 582882 511398 586302 511634
rect 586538 511398 586622 511634
rect 586858 511398 592650 511634
rect -8726 511366 592650 511398
rect -8726 507454 592650 507486
rect -8726 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 73826 507454
rect 74062 507218 74146 507454
rect 74382 507218 109826 507454
rect 110062 507218 110146 507454
rect 110382 507218 145826 507454
rect 146062 507218 146146 507454
rect 146382 507218 181826 507454
rect 182062 507218 182146 507454
rect 182382 507218 217826 507454
rect 218062 507218 218146 507454
rect 218382 507218 253826 507454
rect 254062 507218 254146 507454
rect 254382 507218 289826 507454
rect 290062 507218 290146 507454
rect 290382 507218 325826 507454
rect 326062 507218 326146 507454
rect 326382 507218 361826 507454
rect 362062 507218 362146 507454
rect 362382 507218 397826 507454
rect 398062 507218 398146 507454
rect 398382 507218 433826 507454
rect 434062 507218 434146 507454
rect 434382 507218 469826 507454
rect 470062 507218 470146 507454
rect 470382 507218 505826 507454
rect 506062 507218 506146 507454
rect 506382 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 592650 507454
rect -8726 507134 592650 507218
rect -8726 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 73826 507134
rect 74062 506898 74146 507134
rect 74382 506898 109826 507134
rect 110062 506898 110146 507134
rect 110382 506898 145826 507134
rect 146062 506898 146146 507134
rect 146382 506898 181826 507134
rect 182062 506898 182146 507134
rect 182382 506898 217826 507134
rect 218062 506898 218146 507134
rect 218382 506898 253826 507134
rect 254062 506898 254146 507134
rect 254382 506898 289826 507134
rect 290062 506898 290146 507134
rect 290382 506898 325826 507134
rect 326062 506898 326146 507134
rect 326382 506898 361826 507134
rect 362062 506898 362146 507134
rect 362382 506898 397826 507134
rect 398062 506898 398146 507134
rect 398382 506898 433826 507134
rect 434062 506898 434146 507134
rect 434382 506898 469826 507134
rect 470062 506898 470146 507134
rect 470382 506898 505826 507134
rect 506062 506898 506146 507134
rect 506382 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 592650 507134
rect -8726 506866 592650 506898
rect -8726 502954 592650 502986
rect -8726 502718 -8694 502954
rect -8458 502718 -8374 502954
rect -8138 502718 33326 502954
rect 33562 502718 33646 502954
rect 33882 502718 69326 502954
rect 69562 502718 69646 502954
rect 69882 502718 105326 502954
rect 105562 502718 105646 502954
rect 105882 502718 141326 502954
rect 141562 502718 141646 502954
rect 141882 502718 177326 502954
rect 177562 502718 177646 502954
rect 177882 502718 213326 502954
rect 213562 502718 213646 502954
rect 213882 502718 249326 502954
rect 249562 502718 249646 502954
rect 249882 502718 285326 502954
rect 285562 502718 285646 502954
rect 285882 502718 321326 502954
rect 321562 502718 321646 502954
rect 321882 502718 357326 502954
rect 357562 502718 357646 502954
rect 357882 502718 393326 502954
rect 393562 502718 393646 502954
rect 393882 502718 429326 502954
rect 429562 502718 429646 502954
rect 429882 502718 465326 502954
rect 465562 502718 465646 502954
rect 465882 502718 501326 502954
rect 501562 502718 501646 502954
rect 501882 502718 537326 502954
rect 537562 502718 537646 502954
rect 537882 502718 573326 502954
rect 573562 502718 573646 502954
rect 573882 502718 592062 502954
rect 592298 502718 592382 502954
rect 592618 502718 592650 502954
rect -8726 502634 592650 502718
rect -8726 502398 -8694 502634
rect -8458 502398 -8374 502634
rect -8138 502398 33326 502634
rect 33562 502398 33646 502634
rect 33882 502398 69326 502634
rect 69562 502398 69646 502634
rect 69882 502398 105326 502634
rect 105562 502398 105646 502634
rect 105882 502398 141326 502634
rect 141562 502398 141646 502634
rect 141882 502398 177326 502634
rect 177562 502398 177646 502634
rect 177882 502398 213326 502634
rect 213562 502398 213646 502634
rect 213882 502398 249326 502634
rect 249562 502398 249646 502634
rect 249882 502398 285326 502634
rect 285562 502398 285646 502634
rect 285882 502398 321326 502634
rect 321562 502398 321646 502634
rect 321882 502398 357326 502634
rect 357562 502398 357646 502634
rect 357882 502398 393326 502634
rect 393562 502398 393646 502634
rect 393882 502398 429326 502634
rect 429562 502398 429646 502634
rect 429882 502398 465326 502634
rect 465562 502398 465646 502634
rect 465882 502398 501326 502634
rect 501562 502398 501646 502634
rect 501882 502398 537326 502634
rect 537562 502398 537646 502634
rect 537882 502398 573326 502634
rect 573562 502398 573646 502634
rect 573882 502398 592062 502634
rect 592298 502398 592382 502634
rect 592618 502398 592650 502634
rect -8726 502366 592650 502398
rect -8726 498454 592650 498486
rect -8726 498218 -7734 498454
rect -7498 498218 -7414 498454
rect -7178 498218 28826 498454
rect 29062 498218 29146 498454
rect 29382 498218 64826 498454
rect 65062 498218 65146 498454
rect 65382 498218 100826 498454
rect 101062 498218 101146 498454
rect 101382 498218 136826 498454
rect 137062 498218 137146 498454
rect 137382 498218 172826 498454
rect 173062 498218 173146 498454
rect 173382 498218 208826 498454
rect 209062 498218 209146 498454
rect 209382 498218 244826 498454
rect 245062 498218 245146 498454
rect 245382 498218 280826 498454
rect 281062 498218 281146 498454
rect 281382 498218 316826 498454
rect 317062 498218 317146 498454
rect 317382 498218 352826 498454
rect 353062 498218 353146 498454
rect 353382 498218 388826 498454
rect 389062 498218 389146 498454
rect 389382 498218 424826 498454
rect 425062 498218 425146 498454
rect 425382 498218 460826 498454
rect 461062 498218 461146 498454
rect 461382 498218 496826 498454
rect 497062 498218 497146 498454
rect 497382 498218 532826 498454
rect 533062 498218 533146 498454
rect 533382 498218 568826 498454
rect 569062 498218 569146 498454
rect 569382 498218 591102 498454
rect 591338 498218 591422 498454
rect 591658 498218 592650 498454
rect -8726 498134 592650 498218
rect -8726 497898 -7734 498134
rect -7498 497898 -7414 498134
rect -7178 497898 28826 498134
rect 29062 497898 29146 498134
rect 29382 497898 64826 498134
rect 65062 497898 65146 498134
rect 65382 497898 100826 498134
rect 101062 497898 101146 498134
rect 101382 497898 136826 498134
rect 137062 497898 137146 498134
rect 137382 497898 172826 498134
rect 173062 497898 173146 498134
rect 173382 497898 208826 498134
rect 209062 497898 209146 498134
rect 209382 497898 244826 498134
rect 245062 497898 245146 498134
rect 245382 497898 280826 498134
rect 281062 497898 281146 498134
rect 281382 497898 316826 498134
rect 317062 497898 317146 498134
rect 317382 497898 352826 498134
rect 353062 497898 353146 498134
rect 353382 497898 388826 498134
rect 389062 497898 389146 498134
rect 389382 497898 424826 498134
rect 425062 497898 425146 498134
rect 425382 497898 460826 498134
rect 461062 497898 461146 498134
rect 461382 497898 496826 498134
rect 497062 497898 497146 498134
rect 497382 497898 532826 498134
rect 533062 497898 533146 498134
rect 533382 497898 568826 498134
rect 569062 497898 569146 498134
rect 569382 497898 591102 498134
rect 591338 497898 591422 498134
rect 591658 497898 592650 498134
rect -8726 497866 592650 497898
rect -8726 493954 592650 493986
rect -8726 493718 -6774 493954
rect -6538 493718 -6454 493954
rect -6218 493718 24326 493954
rect 24562 493718 24646 493954
rect 24882 493718 60326 493954
rect 60562 493718 60646 493954
rect 60882 493718 96326 493954
rect 96562 493718 96646 493954
rect 96882 493718 132326 493954
rect 132562 493718 132646 493954
rect 132882 493718 168326 493954
rect 168562 493718 168646 493954
rect 168882 493718 204326 493954
rect 204562 493718 204646 493954
rect 204882 493718 240326 493954
rect 240562 493718 240646 493954
rect 240882 493718 276326 493954
rect 276562 493718 276646 493954
rect 276882 493718 312326 493954
rect 312562 493718 312646 493954
rect 312882 493718 348326 493954
rect 348562 493718 348646 493954
rect 348882 493718 384326 493954
rect 384562 493718 384646 493954
rect 384882 493718 420326 493954
rect 420562 493718 420646 493954
rect 420882 493718 456326 493954
rect 456562 493718 456646 493954
rect 456882 493718 492326 493954
rect 492562 493718 492646 493954
rect 492882 493718 528326 493954
rect 528562 493718 528646 493954
rect 528882 493718 564326 493954
rect 564562 493718 564646 493954
rect 564882 493718 590142 493954
rect 590378 493718 590462 493954
rect 590698 493718 592650 493954
rect -8726 493634 592650 493718
rect -8726 493398 -6774 493634
rect -6538 493398 -6454 493634
rect -6218 493398 24326 493634
rect 24562 493398 24646 493634
rect 24882 493398 60326 493634
rect 60562 493398 60646 493634
rect 60882 493398 96326 493634
rect 96562 493398 96646 493634
rect 96882 493398 132326 493634
rect 132562 493398 132646 493634
rect 132882 493398 168326 493634
rect 168562 493398 168646 493634
rect 168882 493398 204326 493634
rect 204562 493398 204646 493634
rect 204882 493398 240326 493634
rect 240562 493398 240646 493634
rect 240882 493398 276326 493634
rect 276562 493398 276646 493634
rect 276882 493398 312326 493634
rect 312562 493398 312646 493634
rect 312882 493398 348326 493634
rect 348562 493398 348646 493634
rect 348882 493398 384326 493634
rect 384562 493398 384646 493634
rect 384882 493398 420326 493634
rect 420562 493398 420646 493634
rect 420882 493398 456326 493634
rect 456562 493398 456646 493634
rect 456882 493398 492326 493634
rect 492562 493398 492646 493634
rect 492882 493398 528326 493634
rect 528562 493398 528646 493634
rect 528882 493398 564326 493634
rect 564562 493398 564646 493634
rect 564882 493398 590142 493634
rect 590378 493398 590462 493634
rect 590698 493398 592650 493634
rect -8726 493366 592650 493398
rect -8726 489454 592650 489486
rect -8726 489218 -5814 489454
rect -5578 489218 -5494 489454
rect -5258 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 55826 489454
rect 56062 489218 56146 489454
rect 56382 489218 91826 489454
rect 92062 489218 92146 489454
rect 92382 489218 127826 489454
rect 128062 489218 128146 489454
rect 128382 489218 163826 489454
rect 164062 489218 164146 489454
rect 164382 489218 199826 489454
rect 200062 489218 200146 489454
rect 200382 489218 235826 489454
rect 236062 489218 236146 489454
rect 236382 489218 271826 489454
rect 272062 489218 272146 489454
rect 272382 489218 307826 489454
rect 308062 489218 308146 489454
rect 308382 489218 343826 489454
rect 344062 489218 344146 489454
rect 344382 489218 379826 489454
rect 380062 489218 380146 489454
rect 380382 489218 415826 489454
rect 416062 489218 416146 489454
rect 416382 489218 451826 489454
rect 452062 489218 452146 489454
rect 452382 489218 487826 489454
rect 488062 489218 488146 489454
rect 488382 489218 523826 489454
rect 524062 489218 524146 489454
rect 524382 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 589182 489454
rect 589418 489218 589502 489454
rect 589738 489218 592650 489454
rect -8726 489134 592650 489218
rect -8726 488898 -5814 489134
rect -5578 488898 -5494 489134
rect -5258 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 55826 489134
rect 56062 488898 56146 489134
rect 56382 488898 91826 489134
rect 92062 488898 92146 489134
rect 92382 488898 127826 489134
rect 128062 488898 128146 489134
rect 128382 488898 163826 489134
rect 164062 488898 164146 489134
rect 164382 488898 199826 489134
rect 200062 488898 200146 489134
rect 200382 488898 235826 489134
rect 236062 488898 236146 489134
rect 236382 488898 271826 489134
rect 272062 488898 272146 489134
rect 272382 488898 307826 489134
rect 308062 488898 308146 489134
rect 308382 488898 343826 489134
rect 344062 488898 344146 489134
rect 344382 488898 379826 489134
rect 380062 488898 380146 489134
rect 380382 488898 415826 489134
rect 416062 488898 416146 489134
rect 416382 488898 451826 489134
rect 452062 488898 452146 489134
rect 452382 488898 487826 489134
rect 488062 488898 488146 489134
rect 488382 488898 523826 489134
rect 524062 488898 524146 489134
rect 524382 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 589182 489134
rect 589418 488898 589502 489134
rect 589738 488898 592650 489134
rect -8726 488866 592650 488898
rect -8726 484954 592650 484986
rect -8726 484718 -4854 484954
rect -4618 484718 -4534 484954
rect -4298 484718 15326 484954
rect 15562 484718 15646 484954
rect 15882 484718 51326 484954
rect 51562 484718 51646 484954
rect 51882 484718 87326 484954
rect 87562 484718 87646 484954
rect 87882 484718 123326 484954
rect 123562 484718 123646 484954
rect 123882 484718 159326 484954
rect 159562 484718 159646 484954
rect 159882 484718 195326 484954
rect 195562 484718 195646 484954
rect 195882 484718 231326 484954
rect 231562 484718 231646 484954
rect 231882 484718 267326 484954
rect 267562 484718 267646 484954
rect 267882 484718 303326 484954
rect 303562 484718 303646 484954
rect 303882 484718 339326 484954
rect 339562 484718 339646 484954
rect 339882 484718 375326 484954
rect 375562 484718 375646 484954
rect 375882 484718 411326 484954
rect 411562 484718 411646 484954
rect 411882 484718 447326 484954
rect 447562 484718 447646 484954
rect 447882 484718 483326 484954
rect 483562 484718 483646 484954
rect 483882 484718 519326 484954
rect 519562 484718 519646 484954
rect 519882 484718 555326 484954
rect 555562 484718 555646 484954
rect 555882 484718 588222 484954
rect 588458 484718 588542 484954
rect 588778 484718 592650 484954
rect -8726 484634 592650 484718
rect -8726 484398 -4854 484634
rect -4618 484398 -4534 484634
rect -4298 484398 15326 484634
rect 15562 484398 15646 484634
rect 15882 484398 51326 484634
rect 51562 484398 51646 484634
rect 51882 484398 87326 484634
rect 87562 484398 87646 484634
rect 87882 484398 123326 484634
rect 123562 484398 123646 484634
rect 123882 484398 159326 484634
rect 159562 484398 159646 484634
rect 159882 484398 195326 484634
rect 195562 484398 195646 484634
rect 195882 484398 231326 484634
rect 231562 484398 231646 484634
rect 231882 484398 267326 484634
rect 267562 484398 267646 484634
rect 267882 484398 303326 484634
rect 303562 484398 303646 484634
rect 303882 484398 339326 484634
rect 339562 484398 339646 484634
rect 339882 484398 375326 484634
rect 375562 484398 375646 484634
rect 375882 484398 411326 484634
rect 411562 484398 411646 484634
rect 411882 484398 447326 484634
rect 447562 484398 447646 484634
rect 447882 484398 483326 484634
rect 483562 484398 483646 484634
rect 483882 484398 519326 484634
rect 519562 484398 519646 484634
rect 519882 484398 555326 484634
rect 555562 484398 555646 484634
rect 555882 484398 588222 484634
rect 588458 484398 588542 484634
rect 588778 484398 592650 484634
rect -8726 484366 592650 484398
rect -8726 480454 592650 480486
rect -8726 480218 -3894 480454
rect -3658 480218 -3574 480454
rect -3338 480218 10826 480454
rect 11062 480218 11146 480454
rect 11382 480218 46826 480454
rect 47062 480218 47146 480454
rect 47382 480218 82826 480454
rect 83062 480218 83146 480454
rect 83382 480218 118826 480454
rect 119062 480218 119146 480454
rect 119382 480218 154826 480454
rect 155062 480218 155146 480454
rect 155382 480218 190826 480454
rect 191062 480218 191146 480454
rect 191382 480218 226826 480454
rect 227062 480218 227146 480454
rect 227382 480218 262826 480454
rect 263062 480218 263146 480454
rect 263382 480218 298826 480454
rect 299062 480218 299146 480454
rect 299382 480218 334826 480454
rect 335062 480218 335146 480454
rect 335382 480218 370826 480454
rect 371062 480218 371146 480454
rect 371382 480218 406826 480454
rect 407062 480218 407146 480454
rect 407382 480218 442826 480454
rect 443062 480218 443146 480454
rect 443382 480218 478826 480454
rect 479062 480218 479146 480454
rect 479382 480218 514826 480454
rect 515062 480218 515146 480454
rect 515382 480218 550826 480454
rect 551062 480218 551146 480454
rect 551382 480218 587262 480454
rect 587498 480218 587582 480454
rect 587818 480218 592650 480454
rect -8726 480134 592650 480218
rect -8726 479898 -3894 480134
rect -3658 479898 -3574 480134
rect -3338 479898 10826 480134
rect 11062 479898 11146 480134
rect 11382 479898 46826 480134
rect 47062 479898 47146 480134
rect 47382 479898 82826 480134
rect 83062 479898 83146 480134
rect 83382 479898 118826 480134
rect 119062 479898 119146 480134
rect 119382 479898 154826 480134
rect 155062 479898 155146 480134
rect 155382 479898 190826 480134
rect 191062 479898 191146 480134
rect 191382 479898 226826 480134
rect 227062 479898 227146 480134
rect 227382 479898 262826 480134
rect 263062 479898 263146 480134
rect 263382 479898 298826 480134
rect 299062 479898 299146 480134
rect 299382 479898 334826 480134
rect 335062 479898 335146 480134
rect 335382 479898 370826 480134
rect 371062 479898 371146 480134
rect 371382 479898 406826 480134
rect 407062 479898 407146 480134
rect 407382 479898 442826 480134
rect 443062 479898 443146 480134
rect 443382 479898 478826 480134
rect 479062 479898 479146 480134
rect 479382 479898 514826 480134
rect 515062 479898 515146 480134
rect 515382 479898 550826 480134
rect 551062 479898 551146 480134
rect 551382 479898 587262 480134
rect 587498 479898 587582 480134
rect 587818 479898 592650 480134
rect -8726 479866 592650 479898
rect -8726 475954 592650 475986
rect -8726 475718 -2934 475954
rect -2698 475718 -2614 475954
rect -2378 475718 6326 475954
rect 6562 475718 6646 475954
rect 6882 475718 42326 475954
rect 42562 475718 42646 475954
rect 42882 475718 78326 475954
rect 78562 475718 78646 475954
rect 78882 475718 114326 475954
rect 114562 475718 114646 475954
rect 114882 475718 150326 475954
rect 150562 475718 150646 475954
rect 150882 475718 186326 475954
rect 186562 475718 186646 475954
rect 186882 475718 222326 475954
rect 222562 475718 222646 475954
rect 222882 475718 258326 475954
rect 258562 475718 258646 475954
rect 258882 475718 294326 475954
rect 294562 475718 294646 475954
rect 294882 475718 330326 475954
rect 330562 475718 330646 475954
rect 330882 475718 366326 475954
rect 366562 475718 366646 475954
rect 366882 475718 402326 475954
rect 402562 475718 402646 475954
rect 402882 475718 438326 475954
rect 438562 475718 438646 475954
rect 438882 475718 474326 475954
rect 474562 475718 474646 475954
rect 474882 475718 510326 475954
rect 510562 475718 510646 475954
rect 510882 475718 546326 475954
rect 546562 475718 546646 475954
rect 546882 475718 582326 475954
rect 582562 475718 582646 475954
rect 582882 475718 586302 475954
rect 586538 475718 586622 475954
rect 586858 475718 592650 475954
rect -8726 475634 592650 475718
rect -8726 475398 -2934 475634
rect -2698 475398 -2614 475634
rect -2378 475398 6326 475634
rect 6562 475398 6646 475634
rect 6882 475398 42326 475634
rect 42562 475398 42646 475634
rect 42882 475398 78326 475634
rect 78562 475398 78646 475634
rect 78882 475398 114326 475634
rect 114562 475398 114646 475634
rect 114882 475398 150326 475634
rect 150562 475398 150646 475634
rect 150882 475398 186326 475634
rect 186562 475398 186646 475634
rect 186882 475398 222326 475634
rect 222562 475398 222646 475634
rect 222882 475398 258326 475634
rect 258562 475398 258646 475634
rect 258882 475398 294326 475634
rect 294562 475398 294646 475634
rect 294882 475398 330326 475634
rect 330562 475398 330646 475634
rect 330882 475398 366326 475634
rect 366562 475398 366646 475634
rect 366882 475398 402326 475634
rect 402562 475398 402646 475634
rect 402882 475398 438326 475634
rect 438562 475398 438646 475634
rect 438882 475398 474326 475634
rect 474562 475398 474646 475634
rect 474882 475398 510326 475634
rect 510562 475398 510646 475634
rect 510882 475398 546326 475634
rect 546562 475398 546646 475634
rect 546882 475398 582326 475634
rect 582562 475398 582646 475634
rect 582882 475398 586302 475634
rect 586538 475398 586622 475634
rect 586858 475398 592650 475634
rect -8726 475366 592650 475398
rect -8726 471454 592650 471486
rect -8726 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 73826 471454
rect 74062 471218 74146 471454
rect 74382 471218 109826 471454
rect 110062 471218 110146 471454
rect 110382 471218 145826 471454
rect 146062 471218 146146 471454
rect 146382 471218 181826 471454
rect 182062 471218 182146 471454
rect 182382 471218 217826 471454
rect 218062 471218 218146 471454
rect 218382 471218 253826 471454
rect 254062 471218 254146 471454
rect 254382 471218 289826 471454
rect 290062 471218 290146 471454
rect 290382 471218 325826 471454
rect 326062 471218 326146 471454
rect 326382 471218 361826 471454
rect 362062 471218 362146 471454
rect 362382 471218 397826 471454
rect 398062 471218 398146 471454
rect 398382 471218 433826 471454
rect 434062 471218 434146 471454
rect 434382 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 592650 471454
rect -8726 471134 592650 471218
rect -8726 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 73826 471134
rect 74062 470898 74146 471134
rect 74382 470898 109826 471134
rect 110062 470898 110146 471134
rect 110382 470898 145826 471134
rect 146062 470898 146146 471134
rect 146382 470898 181826 471134
rect 182062 470898 182146 471134
rect 182382 470898 217826 471134
rect 218062 470898 218146 471134
rect 218382 470898 253826 471134
rect 254062 470898 254146 471134
rect 254382 470898 289826 471134
rect 290062 470898 290146 471134
rect 290382 470898 325826 471134
rect 326062 470898 326146 471134
rect 326382 470898 361826 471134
rect 362062 470898 362146 471134
rect 362382 470898 397826 471134
rect 398062 470898 398146 471134
rect 398382 470898 433826 471134
rect 434062 470898 434146 471134
rect 434382 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 592650 471134
rect -8726 470866 592650 470898
rect -8726 466954 592650 466986
rect -8726 466718 -8694 466954
rect -8458 466718 -8374 466954
rect -8138 466718 33326 466954
rect 33562 466718 33646 466954
rect 33882 466718 69326 466954
rect 69562 466718 69646 466954
rect 69882 466718 105326 466954
rect 105562 466718 105646 466954
rect 105882 466718 141326 466954
rect 141562 466718 141646 466954
rect 141882 466718 177326 466954
rect 177562 466718 177646 466954
rect 177882 466718 213326 466954
rect 213562 466718 213646 466954
rect 213882 466718 249326 466954
rect 249562 466718 249646 466954
rect 249882 466718 285326 466954
rect 285562 466718 285646 466954
rect 285882 466718 321326 466954
rect 321562 466718 321646 466954
rect 321882 466718 357326 466954
rect 357562 466718 357646 466954
rect 357882 466718 393326 466954
rect 393562 466718 393646 466954
rect 393882 466718 429326 466954
rect 429562 466718 429646 466954
rect 429882 466718 465326 466954
rect 465562 466718 465646 466954
rect 465882 466718 501326 466954
rect 501562 466718 501646 466954
rect 501882 466718 537326 466954
rect 537562 466718 537646 466954
rect 537882 466718 573326 466954
rect 573562 466718 573646 466954
rect 573882 466718 592062 466954
rect 592298 466718 592382 466954
rect 592618 466718 592650 466954
rect -8726 466634 592650 466718
rect -8726 466398 -8694 466634
rect -8458 466398 -8374 466634
rect -8138 466398 33326 466634
rect 33562 466398 33646 466634
rect 33882 466398 69326 466634
rect 69562 466398 69646 466634
rect 69882 466398 105326 466634
rect 105562 466398 105646 466634
rect 105882 466398 141326 466634
rect 141562 466398 141646 466634
rect 141882 466398 177326 466634
rect 177562 466398 177646 466634
rect 177882 466398 213326 466634
rect 213562 466398 213646 466634
rect 213882 466398 249326 466634
rect 249562 466398 249646 466634
rect 249882 466398 285326 466634
rect 285562 466398 285646 466634
rect 285882 466398 321326 466634
rect 321562 466398 321646 466634
rect 321882 466398 357326 466634
rect 357562 466398 357646 466634
rect 357882 466398 393326 466634
rect 393562 466398 393646 466634
rect 393882 466398 429326 466634
rect 429562 466398 429646 466634
rect 429882 466398 465326 466634
rect 465562 466398 465646 466634
rect 465882 466398 501326 466634
rect 501562 466398 501646 466634
rect 501882 466398 537326 466634
rect 537562 466398 537646 466634
rect 537882 466398 573326 466634
rect 573562 466398 573646 466634
rect 573882 466398 592062 466634
rect 592298 466398 592382 466634
rect 592618 466398 592650 466634
rect -8726 466366 592650 466398
rect -8726 462454 592650 462486
rect -8726 462218 -7734 462454
rect -7498 462218 -7414 462454
rect -7178 462218 28826 462454
rect 29062 462218 29146 462454
rect 29382 462218 64826 462454
rect 65062 462218 65146 462454
rect 65382 462218 100826 462454
rect 101062 462218 101146 462454
rect 101382 462218 136826 462454
rect 137062 462218 137146 462454
rect 137382 462218 172826 462454
rect 173062 462218 173146 462454
rect 173382 462218 208826 462454
rect 209062 462218 209146 462454
rect 209382 462218 244826 462454
rect 245062 462218 245146 462454
rect 245382 462218 280826 462454
rect 281062 462218 281146 462454
rect 281382 462218 316826 462454
rect 317062 462218 317146 462454
rect 317382 462218 352826 462454
rect 353062 462218 353146 462454
rect 353382 462218 388826 462454
rect 389062 462218 389146 462454
rect 389382 462218 424826 462454
rect 425062 462218 425146 462454
rect 425382 462218 460826 462454
rect 461062 462218 461146 462454
rect 461382 462218 496826 462454
rect 497062 462218 497146 462454
rect 497382 462218 532826 462454
rect 533062 462218 533146 462454
rect 533382 462218 568826 462454
rect 569062 462218 569146 462454
rect 569382 462218 591102 462454
rect 591338 462218 591422 462454
rect 591658 462218 592650 462454
rect -8726 462134 592650 462218
rect -8726 461898 -7734 462134
rect -7498 461898 -7414 462134
rect -7178 461898 28826 462134
rect 29062 461898 29146 462134
rect 29382 461898 64826 462134
rect 65062 461898 65146 462134
rect 65382 461898 100826 462134
rect 101062 461898 101146 462134
rect 101382 461898 136826 462134
rect 137062 461898 137146 462134
rect 137382 461898 172826 462134
rect 173062 461898 173146 462134
rect 173382 461898 208826 462134
rect 209062 461898 209146 462134
rect 209382 461898 244826 462134
rect 245062 461898 245146 462134
rect 245382 461898 280826 462134
rect 281062 461898 281146 462134
rect 281382 461898 316826 462134
rect 317062 461898 317146 462134
rect 317382 461898 352826 462134
rect 353062 461898 353146 462134
rect 353382 461898 388826 462134
rect 389062 461898 389146 462134
rect 389382 461898 424826 462134
rect 425062 461898 425146 462134
rect 425382 461898 460826 462134
rect 461062 461898 461146 462134
rect 461382 461898 496826 462134
rect 497062 461898 497146 462134
rect 497382 461898 532826 462134
rect 533062 461898 533146 462134
rect 533382 461898 568826 462134
rect 569062 461898 569146 462134
rect 569382 461898 591102 462134
rect 591338 461898 591422 462134
rect 591658 461898 592650 462134
rect -8726 461866 592650 461898
rect -8726 457954 592650 457986
rect -8726 457718 -6774 457954
rect -6538 457718 -6454 457954
rect -6218 457718 24326 457954
rect 24562 457718 24646 457954
rect 24882 457718 60326 457954
rect 60562 457718 60646 457954
rect 60882 457718 96326 457954
rect 96562 457718 96646 457954
rect 96882 457718 132326 457954
rect 132562 457718 132646 457954
rect 132882 457718 168326 457954
rect 168562 457718 168646 457954
rect 168882 457718 204326 457954
rect 204562 457718 204646 457954
rect 204882 457718 240326 457954
rect 240562 457718 240646 457954
rect 240882 457718 276326 457954
rect 276562 457718 276646 457954
rect 276882 457718 312326 457954
rect 312562 457718 312646 457954
rect 312882 457718 348326 457954
rect 348562 457718 348646 457954
rect 348882 457718 384326 457954
rect 384562 457718 384646 457954
rect 384882 457718 420326 457954
rect 420562 457718 420646 457954
rect 420882 457718 456326 457954
rect 456562 457718 456646 457954
rect 456882 457718 492326 457954
rect 492562 457718 492646 457954
rect 492882 457718 528326 457954
rect 528562 457718 528646 457954
rect 528882 457718 564326 457954
rect 564562 457718 564646 457954
rect 564882 457718 590142 457954
rect 590378 457718 590462 457954
rect 590698 457718 592650 457954
rect -8726 457634 592650 457718
rect -8726 457398 -6774 457634
rect -6538 457398 -6454 457634
rect -6218 457398 24326 457634
rect 24562 457398 24646 457634
rect 24882 457398 60326 457634
rect 60562 457398 60646 457634
rect 60882 457398 96326 457634
rect 96562 457398 96646 457634
rect 96882 457398 132326 457634
rect 132562 457398 132646 457634
rect 132882 457398 168326 457634
rect 168562 457398 168646 457634
rect 168882 457398 204326 457634
rect 204562 457398 204646 457634
rect 204882 457398 240326 457634
rect 240562 457398 240646 457634
rect 240882 457398 276326 457634
rect 276562 457398 276646 457634
rect 276882 457398 312326 457634
rect 312562 457398 312646 457634
rect 312882 457398 348326 457634
rect 348562 457398 348646 457634
rect 348882 457398 384326 457634
rect 384562 457398 384646 457634
rect 384882 457398 420326 457634
rect 420562 457398 420646 457634
rect 420882 457398 456326 457634
rect 456562 457398 456646 457634
rect 456882 457398 492326 457634
rect 492562 457398 492646 457634
rect 492882 457398 528326 457634
rect 528562 457398 528646 457634
rect 528882 457398 564326 457634
rect 564562 457398 564646 457634
rect 564882 457398 590142 457634
rect 590378 457398 590462 457634
rect 590698 457398 592650 457634
rect -8726 457366 592650 457398
rect -8726 453454 592650 453486
rect -8726 453218 -5814 453454
rect -5578 453218 -5494 453454
rect -5258 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 55826 453454
rect 56062 453218 56146 453454
rect 56382 453218 91826 453454
rect 92062 453218 92146 453454
rect 92382 453218 127826 453454
rect 128062 453218 128146 453454
rect 128382 453218 163826 453454
rect 164062 453218 164146 453454
rect 164382 453218 199826 453454
rect 200062 453218 200146 453454
rect 200382 453218 235826 453454
rect 236062 453218 236146 453454
rect 236382 453218 271826 453454
rect 272062 453218 272146 453454
rect 272382 453218 307826 453454
rect 308062 453218 308146 453454
rect 308382 453218 343826 453454
rect 344062 453218 344146 453454
rect 344382 453218 379826 453454
rect 380062 453218 380146 453454
rect 380382 453218 415826 453454
rect 416062 453218 416146 453454
rect 416382 453218 451826 453454
rect 452062 453218 452146 453454
rect 452382 453218 487826 453454
rect 488062 453218 488146 453454
rect 488382 453218 523826 453454
rect 524062 453218 524146 453454
rect 524382 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 589182 453454
rect 589418 453218 589502 453454
rect 589738 453218 592650 453454
rect -8726 453134 592650 453218
rect -8726 452898 -5814 453134
rect -5578 452898 -5494 453134
rect -5258 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 55826 453134
rect 56062 452898 56146 453134
rect 56382 452898 91826 453134
rect 92062 452898 92146 453134
rect 92382 452898 127826 453134
rect 128062 452898 128146 453134
rect 128382 452898 163826 453134
rect 164062 452898 164146 453134
rect 164382 452898 199826 453134
rect 200062 452898 200146 453134
rect 200382 452898 235826 453134
rect 236062 452898 236146 453134
rect 236382 452898 271826 453134
rect 272062 452898 272146 453134
rect 272382 452898 307826 453134
rect 308062 452898 308146 453134
rect 308382 452898 343826 453134
rect 344062 452898 344146 453134
rect 344382 452898 379826 453134
rect 380062 452898 380146 453134
rect 380382 452898 415826 453134
rect 416062 452898 416146 453134
rect 416382 452898 451826 453134
rect 452062 452898 452146 453134
rect 452382 452898 487826 453134
rect 488062 452898 488146 453134
rect 488382 452898 523826 453134
rect 524062 452898 524146 453134
rect 524382 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 589182 453134
rect 589418 452898 589502 453134
rect 589738 452898 592650 453134
rect -8726 452866 592650 452898
rect -8726 448954 592650 448986
rect -8726 448718 -4854 448954
rect -4618 448718 -4534 448954
rect -4298 448718 15326 448954
rect 15562 448718 15646 448954
rect 15882 448718 51326 448954
rect 51562 448718 51646 448954
rect 51882 448718 87326 448954
rect 87562 448718 87646 448954
rect 87882 448718 123326 448954
rect 123562 448718 123646 448954
rect 123882 448718 159326 448954
rect 159562 448718 159646 448954
rect 159882 448718 195326 448954
rect 195562 448718 195646 448954
rect 195882 448718 231326 448954
rect 231562 448718 231646 448954
rect 231882 448718 267326 448954
rect 267562 448718 267646 448954
rect 267882 448718 303326 448954
rect 303562 448718 303646 448954
rect 303882 448718 339326 448954
rect 339562 448718 339646 448954
rect 339882 448718 375326 448954
rect 375562 448718 375646 448954
rect 375882 448718 411326 448954
rect 411562 448718 411646 448954
rect 411882 448718 447326 448954
rect 447562 448718 447646 448954
rect 447882 448718 483326 448954
rect 483562 448718 483646 448954
rect 483882 448718 519326 448954
rect 519562 448718 519646 448954
rect 519882 448718 555326 448954
rect 555562 448718 555646 448954
rect 555882 448718 588222 448954
rect 588458 448718 588542 448954
rect 588778 448718 592650 448954
rect -8726 448634 592650 448718
rect -8726 448398 -4854 448634
rect -4618 448398 -4534 448634
rect -4298 448398 15326 448634
rect 15562 448398 15646 448634
rect 15882 448398 51326 448634
rect 51562 448398 51646 448634
rect 51882 448398 87326 448634
rect 87562 448398 87646 448634
rect 87882 448398 123326 448634
rect 123562 448398 123646 448634
rect 123882 448398 159326 448634
rect 159562 448398 159646 448634
rect 159882 448398 195326 448634
rect 195562 448398 195646 448634
rect 195882 448398 231326 448634
rect 231562 448398 231646 448634
rect 231882 448398 267326 448634
rect 267562 448398 267646 448634
rect 267882 448398 303326 448634
rect 303562 448398 303646 448634
rect 303882 448398 339326 448634
rect 339562 448398 339646 448634
rect 339882 448398 375326 448634
rect 375562 448398 375646 448634
rect 375882 448398 411326 448634
rect 411562 448398 411646 448634
rect 411882 448398 447326 448634
rect 447562 448398 447646 448634
rect 447882 448398 483326 448634
rect 483562 448398 483646 448634
rect 483882 448398 519326 448634
rect 519562 448398 519646 448634
rect 519882 448398 555326 448634
rect 555562 448398 555646 448634
rect 555882 448398 588222 448634
rect 588458 448398 588542 448634
rect 588778 448398 592650 448634
rect -8726 448366 592650 448398
rect -8726 444454 592650 444486
rect -8726 444218 -3894 444454
rect -3658 444218 -3574 444454
rect -3338 444218 10826 444454
rect 11062 444218 11146 444454
rect 11382 444218 46826 444454
rect 47062 444218 47146 444454
rect 47382 444218 82826 444454
rect 83062 444218 83146 444454
rect 83382 444218 118826 444454
rect 119062 444218 119146 444454
rect 119382 444218 154826 444454
rect 155062 444218 155146 444454
rect 155382 444218 190826 444454
rect 191062 444218 191146 444454
rect 191382 444218 226826 444454
rect 227062 444218 227146 444454
rect 227382 444218 262826 444454
rect 263062 444218 263146 444454
rect 263382 444218 298826 444454
rect 299062 444218 299146 444454
rect 299382 444218 334826 444454
rect 335062 444218 335146 444454
rect 335382 444218 370826 444454
rect 371062 444218 371146 444454
rect 371382 444218 406826 444454
rect 407062 444218 407146 444454
rect 407382 444218 442826 444454
rect 443062 444218 443146 444454
rect 443382 444218 478826 444454
rect 479062 444218 479146 444454
rect 479382 444218 514826 444454
rect 515062 444218 515146 444454
rect 515382 444218 550826 444454
rect 551062 444218 551146 444454
rect 551382 444218 587262 444454
rect 587498 444218 587582 444454
rect 587818 444218 592650 444454
rect -8726 444134 592650 444218
rect -8726 443898 -3894 444134
rect -3658 443898 -3574 444134
rect -3338 443898 10826 444134
rect 11062 443898 11146 444134
rect 11382 443898 46826 444134
rect 47062 443898 47146 444134
rect 47382 443898 82826 444134
rect 83062 443898 83146 444134
rect 83382 443898 118826 444134
rect 119062 443898 119146 444134
rect 119382 443898 154826 444134
rect 155062 443898 155146 444134
rect 155382 443898 190826 444134
rect 191062 443898 191146 444134
rect 191382 443898 226826 444134
rect 227062 443898 227146 444134
rect 227382 443898 262826 444134
rect 263062 443898 263146 444134
rect 263382 443898 298826 444134
rect 299062 443898 299146 444134
rect 299382 443898 334826 444134
rect 335062 443898 335146 444134
rect 335382 443898 370826 444134
rect 371062 443898 371146 444134
rect 371382 443898 406826 444134
rect 407062 443898 407146 444134
rect 407382 443898 442826 444134
rect 443062 443898 443146 444134
rect 443382 443898 478826 444134
rect 479062 443898 479146 444134
rect 479382 443898 514826 444134
rect 515062 443898 515146 444134
rect 515382 443898 550826 444134
rect 551062 443898 551146 444134
rect 551382 443898 587262 444134
rect 587498 443898 587582 444134
rect 587818 443898 592650 444134
rect -8726 443866 592650 443898
rect -8726 439954 592650 439986
rect -8726 439718 -2934 439954
rect -2698 439718 -2614 439954
rect -2378 439718 6326 439954
rect 6562 439718 6646 439954
rect 6882 439718 42326 439954
rect 42562 439718 42646 439954
rect 42882 439718 78326 439954
rect 78562 439718 78646 439954
rect 78882 439718 114326 439954
rect 114562 439718 114646 439954
rect 114882 439718 150326 439954
rect 150562 439718 150646 439954
rect 150882 439718 186326 439954
rect 186562 439718 186646 439954
rect 186882 439718 222326 439954
rect 222562 439718 222646 439954
rect 222882 439718 258326 439954
rect 258562 439718 258646 439954
rect 258882 439718 294326 439954
rect 294562 439718 294646 439954
rect 294882 439718 330326 439954
rect 330562 439718 330646 439954
rect 330882 439718 366326 439954
rect 366562 439718 366646 439954
rect 366882 439718 402326 439954
rect 402562 439718 402646 439954
rect 402882 439718 438326 439954
rect 438562 439718 438646 439954
rect 438882 439718 474326 439954
rect 474562 439718 474646 439954
rect 474882 439718 510326 439954
rect 510562 439718 510646 439954
rect 510882 439718 546326 439954
rect 546562 439718 546646 439954
rect 546882 439718 582326 439954
rect 582562 439718 582646 439954
rect 582882 439718 586302 439954
rect 586538 439718 586622 439954
rect 586858 439718 592650 439954
rect -8726 439634 592650 439718
rect -8726 439398 -2934 439634
rect -2698 439398 -2614 439634
rect -2378 439398 6326 439634
rect 6562 439398 6646 439634
rect 6882 439398 42326 439634
rect 42562 439398 42646 439634
rect 42882 439398 78326 439634
rect 78562 439398 78646 439634
rect 78882 439398 114326 439634
rect 114562 439398 114646 439634
rect 114882 439398 150326 439634
rect 150562 439398 150646 439634
rect 150882 439398 186326 439634
rect 186562 439398 186646 439634
rect 186882 439398 222326 439634
rect 222562 439398 222646 439634
rect 222882 439398 258326 439634
rect 258562 439398 258646 439634
rect 258882 439398 294326 439634
rect 294562 439398 294646 439634
rect 294882 439398 330326 439634
rect 330562 439398 330646 439634
rect 330882 439398 366326 439634
rect 366562 439398 366646 439634
rect 366882 439398 402326 439634
rect 402562 439398 402646 439634
rect 402882 439398 438326 439634
rect 438562 439398 438646 439634
rect 438882 439398 474326 439634
rect 474562 439398 474646 439634
rect 474882 439398 510326 439634
rect 510562 439398 510646 439634
rect 510882 439398 546326 439634
rect 546562 439398 546646 439634
rect 546882 439398 582326 439634
rect 582562 439398 582646 439634
rect 582882 439398 586302 439634
rect 586538 439398 586622 439634
rect 586858 439398 592650 439634
rect -8726 439366 592650 439398
rect -8726 435454 592650 435486
rect -8726 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 73826 435454
rect 74062 435218 74146 435454
rect 74382 435218 109826 435454
rect 110062 435218 110146 435454
rect 110382 435218 145826 435454
rect 146062 435218 146146 435454
rect 146382 435218 181826 435454
rect 182062 435218 182146 435454
rect 182382 435218 217826 435454
rect 218062 435218 218146 435454
rect 218382 435218 253826 435454
rect 254062 435218 254146 435454
rect 254382 435218 289826 435454
rect 290062 435218 290146 435454
rect 290382 435218 325826 435454
rect 326062 435218 326146 435454
rect 326382 435218 361826 435454
rect 362062 435218 362146 435454
rect 362382 435218 397826 435454
rect 398062 435218 398146 435454
rect 398382 435218 433826 435454
rect 434062 435218 434146 435454
rect 434382 435218 469826 435454
rect 470062 435218 470146 435454
rect 470382 435218 505826 435454
rect 506062 435218 506146 435454
rect 506382 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 592650 435454
rect -8726 435134 592650 435218
rect -8726 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 73826 435134
rect 74062 434898 74146 435134
rect 74382 434898 109826 435134
rect 110062 434898 110146 435134
rect 110382 434898 145826 435134
rect 146062 434898 146146 435134
rect 146382 434898 181826 435134
rect 182062 434898 182146 435134
rect 182382 434898 217826 435134
rect 218062 434898 218146 435134
rect 218382 434898 253826 435134
rect 254062 434898 254146 435134
rect 254382 434898 289826 435134
rect 290062 434898 290146 435134
rect 290382 434898 325826 435134
rect 326062 434898 326146 435134
rect 326382 434898 361826 435134
rect 362062 434898 362146 435134
rect 362382 434898 397826 435134
rect 398062 434898 398146 435134
rect 398382 434898 433826 435134
rect 434062 434898 434146 435134
rect 434382 434898 469826 435134
rect 470062 434898 470146 435134
rect 470382 434898 505826 435134
rect 506062 434898 506146 435134
rect 506382 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 592650 435134
rect -8726 434866 592650 434898
rect -8726 430954 592650 430986
rect -8726 430718 -8694 430954
rect -8458 430718 -8374 430954
rect -8138 430718 33326 430954
rect 33562 430718 33646 430954
rect 33882 430718 69326 430954
rect 69562 430718 69646 430954
rect 69882 430718 105326 430954
rect 105562 430718 105646 430954
rect 105882 430718 141326 430954
rect 141562 430718 141646 430954
rect 141882 430718 177326 430954
rect 177562 430718 177646 430954
rect 177882 430718 213326 430954
rect 213562 430718 213646 430954
rect 213882 430718 249326 430954
rect 249562 430718 249646 430954
rect 249882 430718 285326 430954
rect 285562 430718 285646 430954
rect 285882 430718 321326 430954
rect 321562 430718 321646 430954
rect 321882 430718 357326 430954
rect 357562 430718 357646 430954
rect 357882 430718 393326 430954
rect 393562 430718 393646 430954
rect 393882 430718 429326 430954
rect 429562 430718 429646 430954
rect 429882 430718 465326 430954
rect 465562 430718 465646 430954
rect 465882 430718 501326 430954
rect 501562 430718 501646 430954
rect 501882 430718 537326 430954
rect 537562 430718 537646 430954
rect 537882 430718 573326 430954
rect 573562 430718 573646 430954
rect 573882 430718 592062 430954
rect 592298 430718 592382 430954
rect 592618 430718 592650 430954
rect -8726 430634 592650 430718
rect -8726 430398 -8694 430634
rect -8458 430398 -8374 430634
rect -8138 430398 33326 430634
rect 33562 430398 33646 430634
rect 33882 430398 69326 430634
rect 69562 430398 69646 430634
rect 69882 430398 105326 430634
rect 105562 430398 105646 430634
rect 105882 430398 141326 430634
rect 141562 430398 141646 430634
rect 141882 430398 177326 430634
rect 177562 430398 177646 430634
rect 177882 430398 213326 430634
rect 213562 430398 213646 430634
rect 213882 430398 249326 430634
rect 249562 430398 249646 430634
rect 249882 430398 285326 430634
rect 285562 430398 285646 430634
rect 285882 430398 321326 430634
rect 321562 430398 321646 430634
rect 321882 430398 357326 430634
rect 357562 430398 357646 430634
rect 357882 430398 393326 430634
rect 393562 430398 393646 430634
rect 393882 430398 429326 430634
rect 429562 430398 429646 430634
rect 429882 430398 465326 430634
rect 465562 430398 465646 430634
rect 465882 430398 501326 430634
rect 501562 430398 501646 430634
rect 501882 430398 537326 430634
rect 537562 430398 537646 430634
rect 537882 430398 573326 430634
rect 573562 430398 573646 430634
rect 573882 430398 592062 430634
rect 592298 430398 592382 430634
rect 592618 430398 592650 430634
rect -8726 430366 592650 430398
rect -8726 426454 592650 426486
rect -8726 426218 -7734 426454
rect -7498 426218 -7414 426454
rect -7178 426218 28826 426454
rect 29062 426218 29146 426454
rect 29382 426218 64826 426454
rect 65062 426218 65146 426454
rect 65382 426218 100826 426454
rect 101062 426218 101146 426454
rect 101382 426218 136826 426454
rect 137062 426218 137146 426454
rect 137382 426218 172826 426454
rect 173062 426218 173146 426454
rect 173382 426218 208826 426454
rect 209062 426218 209146 426454
rect 209382 426218 244826 426454
rect 245062 426218 245146 426454
rect 245382 426218 280826 426454
rect 281062 426218 281146 426454
rect 281382 426218 316826 426454
rect 317062 426218 317146 426454
rect 317382 426218 352826 426454
rect 353062 426218 353146 426454
rect 353382 426218 388826 426454
rect 389062 426218 389146 426454
rect 389382 426218 424826 426454
rect 425062 426218 425146 426454
rect 425382 426218 460826 426454
rect 461062 426218 461146 426454
rect 461382 426218 496826 426454
rect 497062 426218 497146 426454
rect 497382 426218 532826 426454
rect 533062 426218 533146 426454
rect 533382 426218 568826 426454
rect 569062 426218 569146 426454
rect 569382 426218 591102 426454
rect 591338 426218 591422 426454
rect 591658 426218 592650 426454
rect -8726 426134 592650 426218
rect -8726 425898 -7734 426134
rect -7498 425898 -7414 426134
rect -7178 425898 28826 426134
rect 29062 425898 29146 426134
rect 29382 425898 64826 426134
rect 65062 425898 65146 426134
rect 65382 425898 100826 426134
rect 101062 425898 101146 426134
rect 101382 425898 136826 426134
rect 137062 425898 137146 426134
rect 137382 425898 172826 426134
rect 173062 425898 173146 426134
rect 173382 425898 208826 426134
rect 209062 425898 209146 426134
rect 209382 425898 244826 426134
rect 245062 425898 245146 426134
rect 245382 425898 280826 426134
rect 281062 425898 281146 426134
rect 281382 425898 316826 426134
rect 317062 425898 317146 426134
rect 317382 425898 352826 426134
rect 353062 425898 353146 426134
rect 353382 425898 388826 426134
rect 389062 425898 389146 426134
rect 389382 425898 424826 426134
rect 425062 425898 425146 426134
rect 425382 425898 460826 426134
rect 461062 425898 461146 426134
rect 461382 425898 496826 426134
rect 497062 425898 497146 426134
rect 497382 425898 532826 426134
rect 533062 425898 533146 426134
rect 533382 425898 568826 426134
rect 569062 425898 569146 426134
rect 569382 425898 591102 426134
rect 591338 425898 591422 426134
rect 591658 425898 592650 426134
rect -8726 425866 592650 425898
rect -8726 421954 592650 421986
rect -8726 421718 -6774 421954
rect -6538 421718 -6454 421954
rect -6218 421718 24326 421954
rect 24562 421718 24646 421954
rect 24882 421718 60326 421954
rect 60562 421718 60646 421954
rect 60882 421718 96326 421954
rect 96562 421718 96646 421954
rect 96882 421718 132326 421954
rect 132562 421718 132646 421954
rect 132882 421718 168326 421954
rect 168562 421718 168646 421954
rect 168882 421718 204326 421954
rect 204562 421718 204646 421954
rect 204882 421718 240326 421954
rect 240562 421718 240646 421954
rect 240882 421718 276326 421954
rect 276562 421718 276646 421954
rect 276882 421718 312326 421954
rect 312562 421718 312646 421954
rect 312882 421718 348326 421954
rect 348562 421718 348646 421954
rect 348882 421718 384326 421954
rect 384562 421718 384646 421954
rect 384882 421718 420326 421954
rect 420562 421718 420646 421954
rect 420882 421718 456326 421954
rect 456562 421718 456646 421954
rect 456882 421718 492326 421954
rect 492562 421718 492646 421954
rect 492882 421718 528326 421954
rect 528562 421718 528646 421954
rect 528882 421718 564326 421954
rect 564562 421718 564646 421954
rect 564882 421718 590142 421954
rect 590378 421718 590462 421954
rect 590698 421718 592650 421954
rect -8726 421634 592650 421718
rect -8726 421398 -6774 421634
rect -6538 421398 -6454 421634
rect -6218 421398 24326 421634
rect 24562 421398 24646 421634
rect 24882 421398 60326 421634
rect 60562 421398 60646 421634
rect 60882 421398 96326 421634
rect 96562 421398 96646 421634
rect 96882 421398 132326 421634
rect 132562 421398 132646 421634
rect 132882 421398 168326 421634
rect 168562 421398 168646 421634
rect 168882 421398 204326 421634
rect 204562 421398 204646 421634
rect 204882 421398 240326 421634
rect 240562 421398 240646 421634
rect 240882 421398 276326 421634
rect 276562 421398 276646 421634
rect 276882 421398 312326 421634
rect 312562 421398 312646 421634
rect 312882 421398 348326 421634
rect 348562 421398 348646 421634
rect 348882 421398 384326 421634
rect 384562 421398 384646 421634
rect 384882 421398 420326 421634
rect 420562 421398 420646 421634
rect 420882 421398 456326 421634
rect 456562 421398 456646 421634
rect 456882 421398 492326 421634
rect 492562 421398 492646 421634
rect 492882 421398 528326 421634
rect 528562 421398 528646 421634
rect 528882 421398 564326 421634
rect 564562 421398 564646 421634
rect 564882 421398 590142 421634
rect 590378 421398 590462 421634
rect 590698 421398 592650 421634
rect -8726 421366 592650 421398
rect -8726 417454 592650 417486
rect -8726 417218 -5814 417454
rect -5578 417218 -5494 417454
rect -5258 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 55826 417454
rect 56062 417218 56146 417454
rect 56382 417218 91826 417454
rect 92062 417218 92146 417454
rect 92382 417218 127826 417454
rect 128062 417218 128146 417454
rect 128382 417218 163826 417454
rect 164062 417218 164146 417454
rect 164382 417218 199826 417454
rect 200062 417218 200146 417454
rect 200382 417218 235826 417454
rect 236062 417218 236146 417454
rect 236382 417218 271826 417454
rect 272062 417218 272146 417454
rect 272382 417218 307826 417454
rect 308062 417218 308146 417454
rect 308382 417218 343826 417454
rect 344062 417218 344146 417454
rect 344382 417218 379826 417454
rect 380062 417218 380146 417454
rect 380382 417218 415826 417454
rect 416062 417218 416146 417454
rect 416382 417218 451826 417454
rect 452062 417218 452146 417454
rect 452382 417218 487826 417454
rect 488062 417218 488146 417454
rect 488382 417218 523826 417454
rect 524062 417218 524146 417454
rect 524382 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 589182 417454
rect 589418 417218 589502 417454
rect 589738 417218 592650 417454
rect -8726 417134 592650 417218
rect -8726 416898 -5814 417134
rect -5578 416898 -5494 417134
rect -5258 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 55826 417134
rect 56062 416898 56146 417134
rect 56382 416898 91826 417134
rect 92062 416898 92146 417134
rect 92382 416898 127826 417134
rect 128062 416898 128146 417134
rect 128382 416898 163826 417134
rect 164062 416898 164146 417134
rect 164382 416898 199826 417134
rect 200062 416898 200146 417134
rect 200382 416898 235826 417134
rect 236062 416898 236146 417134
rect 236382 416898 271826 417134
rect 272062 416898 272146 417134
rect 272382 416898 307826 417134
rect 308062 416898 308146 417134
rect 308382 416898 343826 417134
rect 344062 416898 344146 417134
rect 344382 416898 379826 417134
rect 380062 416898 380146 417134
rect 380382 416898 415826 417134
rect 416062 416898 416146 417134
rect 416382 416898 451826 417134
rect 452062 416898 452146 417134
rect 452382 416898 487826 417134
rect 488062 416898 488146 417134
rect 488382 416898 523826 417134
rect 524062 416898 524146 417134
rect 524382 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 589182 417134
rect 589418 416898 589502 417134
rect 589738 416898 592650 417134
rect -8726 416866 592650 416898
rect -8726 412954 592650 412986
rect -8726 412718 -4854 412954
rect -4618 412718 -4534 412954
rect -4298 412718 15326 412954
rect 15562 412718 15646 412954
rect 15882 412718 51326 412954
rect 51562 412718 51646 412954
rect 51882 412718 87326 412954
rect 87562 412718 87646 412954
rect 87882 412718 123326 412954
rect 123562 412718 123646 412954
rect 123882 412718 159326 412954
rect 159562 412718 159646 412954
rect 159882 412718 195326 412954
rect 195562 412718 195646 412954
rect 195882 412718 231326 412954
rect 231562 412718 231646 412954
rect 231882 412718 267326 412954
rect 267562 412718 267646 412954
rect 267882 412718 303326 412954
rect 303562 412718 303646 412954
rect 303882 412718 339326 412954
rect 339562 412718 339646 412954
rect 339882 412718 375326 412954
rect 375562 412718 375646 412954
rect 375882 412718 411326 412954
rect 411562 412718 411646 412954
rect 411882 412718 447326 412954
rect 447562 412718 447646 412954
rect 447882 412718 483326 412954
rect 483562 412718 483646 412954
rect 483882 412718 519326 412954
rect 519562 412718 519646 412954
rect 519882 412718 555326 412954
rect 555562 412718 555646 412954
rect 555882 412718 588222 412954
rect 588458 412718 588542 412954
rect 588778 412718 592650 412954
rect -8726 412634 592650 412718
rect -8726 412398 -4854 412634
rect -4618 412398 -4534 412634
rect -4298 412398 15326 412634
rect 15562 412398 15646 412634
rect 15882 412398 51326 412634
rect 51562 412398 51646 412634
rect 51882 412398 87326 412634
rect 87562 412398 87646 412634
rect 87882 412398 123326 412634
rect 123562 412398 123646 412634
rect 123882 412398 159326 412634
rect 159562 412398 159646 412634
rect 159882 412398 195326 412634
rect 195562 412398 195646 412634
rect 195882 412398 231326 412634
rect 231562 412398 231646 412634
rect 231882 412398 267326 412634
rect 267562 412398 267646 412634
rect 267882 412398 303326 412634
rect 303562 412398 303646 412634
rect 303882 412398 339326 412634
rect 339562 412398 339646 412634
rect 339882 412398 375326 412634
rect 375562 412398 375646 412634
rect 375882 412398 411326 412634
rect 411562 412398 411646 412634
rect 411882 412398 447326 412634
rect 447562 412398 447646 412634
rect 447882 412398 483326 412634
rect 483562 412398 483646 412634
rect 483882 412398 519326 412634
rect 519562 412398 519646 412634
rect 519882 412398 555326 412634
rect 555562 412398 555646 412634
rect 555882 412398 588222 412634
rect 588458 412398 588542 412634
rect 588778 412398 592650 412634
rect -8726 412366 592650 412398
rect -8726 408454 592650 408486
rect -8726 408218 -3894 408454
rect -3658 408218 -3574 408454
rect -3338 408218 10826 408454
rect 11062 408218 11146 408454
rect 11382 408218 46826 408454
rect 47062 408218 47146 408454
rect 47382 408218 82826 408454
rect 83062 408218 83146 408454
rect 83382 408218 118826 408454
rect 119062 408218 119146 408454
rect 119382 408218 154826 408454
rect 155062 408218 155146 408454
rect 155382 408218 190826 408454
rect 191062 408218 191146 408454
rect 191382 408218 226826 408454
rect 227062 408218 227146 408454
rect 227382 408218 262826 408454
rect 263062 408218 263146 408454
rect 263382 408218 298826 408454
rect 299062 408218 299146 408454
rect 299382 408218 334826 408454
rect 335062 408218 335146 408454
rect 335382 408218 370826 408454
rect 371062 408218 371146 408454
rect 371382 408218 406826 408454
rect 407062 408218 407146 408454
rect 407382 408218 442826 408454
rect 443062 408218 443146 408454
rect 443382 408218 478826 408454
rect 479062 408218 479146 408454
rect 479382 408218 514826 408454
rect 515062 408218 515146 408454
rect 515382 408218 550826 408454
rect 551062 408218 551146 408454
rect 551382 408218 587262 408454
rect 587498 408218 587582 408454
rect 587818 408218 592650 408454
rect -8726 408134 592650 408218
rect -8726 407898 -3894 408134
rect -3658 407898 -3574 408134
rect -3338 407898 10826 408134
rect 11062 407898 11146 408134
rect 11382 407898 46826 408134
rect 47062 407898 47146 408134
rect 47382 407898 82826 408134
rect 83062 407898 83146 408134
rect 83382 407898 118826 408134
rect 119062 407898 119146 408134
rect 119382 407898 154826 408134
rect 155062 407898 155146 408134
rect 155382 407898 190826 408134
rect 191062 407898 191146 408134
rect 191382 407898 226826 408134
rect 227062 407898 227146 408134
rect 227382 407898 262826 408134
rect 263062 407898 263146 408134
rect 263382 407898 298826 408134
rect 299062 407898 299146 408134
rect 299382 407898 334826 408134
rect 335062 407898 335146 408134
rect 335382 407898 370826 408134
rect 371062 407898 371146 408134
rect 371382 407898 406826 408134
rect 407062 407898 407146 408134
rect 407382 407898 442826 408134
rect 443062 407898 443146 408134
rect 443382 407898 478826 408134
rect 479062 407898 479146 408134
rect 479382 407898 514826 408134
rect 515062 407898 515146 408134
rect 515382 407898 550826 408134
rect 551062 407898 551146 408134
rect 551382 407898 587262 408134
rect 587498 407898 587582 408134
rect 587818 407898 592650 408134
rect -8726 407866 592650 407898
rect -8726 403954 592650 403986
rect -8726 403718 -2934 403954
rect -2698 403718 -2614 403954
rect -2378 403718 6326 403954
rect 6562 403718 6646 403954
rect 6882 403718 42326 403954
rect 42562 403718 42646 403954
rect 42882 403718 78326 403954
rect 78562 403718 78646 403954
rect 78882 403718 114326 403954
rect 114562 403718 114646 403954
rect 114882 403718 150326 403954
rect 150562 403718 150646 403954
rect 150882 403718 186326 403954
rect 186562 403718 186646 403954
rect 186882 403718 222326 403954
rect 222562 403718 222646 403954
rect 222882 403718 258326 403954
rect 258562 403718 258646 403954
rect 258882 403718 294326 403954
rect 294562 403718 294646 403954
rect 294882 403718 330326 403954
rect 330562 403718 330646 403954
rect 330882 403718 366326 403954
rect 366562 403718 366646 403954
rect 366882 403718 402326 403954
rect 402562 403718 402646 403954
rect 402882 403718 438326 403954
rect 438562 403718 438646 403954
rect 438882 403718 474326 403954
rect 474562 403718 474646 403954
rect 474882 403718 510326 403954
rect 510562 403718 510646 403954
rect 510882 403718 546326 403954
rect 546562 403718 546646 403954
rect 546882 403718 582326 403954
rect 582562 403718 582646 403954
rect 582882 403718 586302 403954
rect 586538 403718 586622 403954
rect 586858 403718 592650 403954
rect -8726 403634 592650 403718
rect -8726 403398 -2934 403634
rect -2698 403398 -2614 403634
rect -2378 403398 6326 403634
rect 6562 403398 6646 403634
rect 6882 403398 42326 403634
rect 42562 403398 42646 403634
rect 42882 403398 78326 403634
rect 78562 403398 78646 403634
rect 78882 403398 114326 403634
rect 114562 403398 114646 403634
rect 114882 403398 150326 403634
rect 150562 403398 150646 403634
rect 150882 403398 186326 403634
rect 186562 403398 186646 403634
rect 186882 403398 222326 403634
rect 222562 403398 222646 403634
rect 222882 403398 258326 403634
rect 258562 403398 258646 403634
rect 258882 403398 294326 403634
rect 294562 403398 294646 403634
rect 294882 403398 330326 403634
rect 330562 403398 330646 403634
rect 330882 403398 366326 403634
rect 366562 403398 366646 403634
rect 366882 403398 402326 403634
rect 402562 403398 402646 403634
rect 402882 403398 438326 403634
rect 438562 403398 438646 403634
rect 438882 403398 474326 403634
rect 474562 403398 474646 403634
rect 474882 403398 510326 403634
rect 510562 403398 510646 403634
rect 510882 403398 546326 403634
rect 546562 403398 546646 403634
rect 546882 403398 582326 403634
rect 582562 403398 582646 403634
rect 582882 403398 586302 403634
rect 586538 403398 586622 403634
rect 586858 403398 592650 403634
rect -8726 403366 592650 403398
rect -8726 399454 592650 399486
rect -8726 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 73826 399454
rect 74062 399218 74146 399454
rect 74382 399218 109826 399454
rect 110062 399218 110146 399454
rect 110382 399218 145826 399454
rect 146062 399218 146146 399454
rect 146382 399218 181826 399454
rect 182062 399218 182146 399454
rect 182382 399218 217826 399454
rect 218062 399218 218146 399454
rect 218382 399218 253826 399454
rect 254062 399218 254146 399454
rect 254382 399218 289826 399454
rect 290062 399218 290146 399454
rect 290382 399218 325826 399454
rect 326062 399218 326146 399454
rect 326382 399218 361826 399454
rect 362062 399218 362146 399454
rect 362382 399218 397826 399454
rect 398062 399218 398146 399454
rect 398382 399218 433826 399454
rect 434062 399218 434146 399454
rect 434382 399218 469826 399454
rect 470062 399218 470146 399454
rect 470382 399218 505826 399454
rect 506062 399218 506146 399454
rect 506382 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 592650 399454
rect -8726 399134 592650 399218
rect -8726 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 73826 399134
rect 74062 398898 74146 399134
rect 74382 398898 109826 399134
rect 110062 398898 110146 399134
rect 110382 398898 145826 399134
rect 146062 398898 146146 399134
rect 146382 398898 181826 399134
rect 182062 398898 182146 399134
rect 182382 398898 217826 399134
rect 218062 398898 218146 399134
rect 218382 398898 253826 399134
rect 254062 398898 254146 399134
rect 254382 398898 289826 399134
rect 290062 398898 290146 399134
rect 290382 398898 325826 399134
rect 326062 398898 326146 399134
rect 326382 398898 361826 399134
rect 362062 398898 362146 399134
rect 362382 398898 397826 399134
rect 398062 398898 398146 399134
rect 398382 398898 433826 399134
rect 434062 398898 434146 399134
rect 434382 398898 469826 399134
rect 470062 398898 470146 399134
rect 470382 398898 505826 399134
rect 506062 398898 506146 399134
rect 506382 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 592650 399134
rect -8726 398866 592650 398898
rect -8726 394954 592650 394986
rect -8726 394718 -8694 394954
rect -8458 394718 -8374 394954
rect -8138 394718 33326 394954
rect 33562 394718 33646 394954
rect 33882 394718 69326 394954
rect 69562 394718 69646 394954
rect 69882 394718 105326 394954
rect 105562 394718 105646 394954
rect 105882 394718 141326 394954
rect 141562 394718 141646 394954
rect 141882 394718 177326 394954
rect 177562 394718 177646 394954
rect 177882 394718 213326 394954
rect 213562 394718 213646 394954
rect 213882 394718 249326 394954
rect 249562 394718 249646 394954
rect 249882 394718 285326 394954
rect 285562 394718 285646 394954
rect 285882 394718 321326 394954
rect 321562 394718 321646 394954
rect 321882 394718 357326 394954
rect 357562 394718 357646 394954
rect 357882 394718 393326 394954
rect 393562 394718 393646 394954
rect 393882 394718 429326 394954
rect 429562 394718 429646 394954
rect 429882 394718 465326 394954
rect 465562 394718 465646 394954
rect 465882 394718 501326 394954
rect 501562 394718 501646 394954
rect 501882 394718 537326 394954
rect 537562 394718 537646 394954
rect 537882 394718 573326 394954
rect 573562 394718 573646 394954
rect 573882 394718 592062 394954
rect 592298 394718 592382 394954
rect 592618 394718 592650 394954
rect -8726 394634 592650 394718
rect -8726 394398 -8694 394634
rect -8458 394398 -8374 394634
rect -8138 394398 33326 394634
rect 33562 394398 33646 394634
rect 33882 394398 69326 394634
rect 69562 394398 69646 394634
rect 69882 394398 105326 394634
rect 105562 394398 105646 394634
rect 105882 394398 141326 394634
rect 141562 394398 141646 394634
rect 141882 394398 177326 394634
rect 177562 394398 177646 394634
rect 177882 394398 213326 394634
rect 213562 394398 213646 394634
rect 213882 394398 249326 394634
rect 249562 394398 249646 394634
rect 249882 394398 285326 394634
rect 285562 394398 285646 394634
rect 285882 394398 321326 394634
rect 321562 394398 321646 394634
rect 321882 394398 357326 394634
rect 357562 394398 357646 394634
rect 357882 394398 393326 394634
rect 393562 394398 393646 394634
rect 393882 394398 429326 394634
rect 429562 394398 429646 394634
rect 429882 394398 465326 394634
rect 465562 394398 465646 394634
rect 465882 394398 501326 394634
rect 501562 394398 501646 394634
rect 501882 394398 537326 394634
rect 537562 394398 537646 394634
rect 537882 394398 573326 394634
rect 573562 394398 573646 394634
rect 573882 394398 592062 394634
rect 592298 394398 592382 394634
rect 592618 394398 592650 394634
rect -8726 394366 592650 394398
rect -8726 390454 592650 390486
rect -8726 390218 -7734 390454
rect -7498 390218 -7414 390454
rect -7178 390218 28826 390454
rect 29062 390218 29146 390454
rect 29382 390218 64826 390454
rect 65062 390218 65146 390454
rect 65382 390218 100826 390454
rect 101062 390218 101146 390454
rect 101382 390218 136826 390454
rect 137062 390218 137146 390454
rect 137382 390218 172826 390454
rect 173062 390218 173146 390454
rect 173382 390218 208826 390454
rect 209062 390218 209146 390454
rect 209382 390218 244826 390454
rect 245062 390218 245146 390454
rect 245382 390218 280826 390454
rect 281062 390218 281146 390454
rect 281382 390218 316826 390454
rect 317062 390218 317146 390454
rect 317382 390218 352826 390454
rect 353062 390218 353146 390454
rect 353382 390218 388826 390454
rect 389062 390218 389146 390454
rect 389382 390218 424826 390454
rect 425062 390218 425146 390454
rect 425382 390218 460826 390454
rect 461062 390218 461146 390454
rect 461382 390218 496826 390454
rect 497062 390218 497146 390454
rect 497382 390218 532826 390454
rect 533062 390218 533146 390454
rect 533382 390218 568826 390454
rect 569062 390218 569146 390454
rect 569382 390218 591102 390454
rect 591338 390218 591422 390454
rect 591658 390218 592650 390454
rect -8726 390134 592650 390218
rect -8726 389898 -7734 390134
rect -7498 389898 -7414 390134
rect -7178 389898 28826 390134
rect 29062 389898 29146 390134
rect 29382 389898 64826 390134
rect 65062 389898 65146 390134
rect 65382 389898 100826 390134
rect 101062 389898 101146 390134
rect 101382 389898 136826 390134
rect 137062 389898 137146 390134
rect 137382 389898 172826 390134
rect 173062 389898 173146 390134
rect 173382 389898 208826 390134
rect 209062 389898 209146 390134
rect 209382 389898 244826 390134
rect 245062 389898 245146 390134
rect 245382 389898 280826 390134
rect 281062 389898 281146 390134
rect 281382 389898 316826 390134
rect 317062 389898 317146 390134
rect 317382 389898 352826 390134
rect 353062 389898 353146 390134
rect 353382 389898 388826 390134
rect 389062 389898 389146 390134
rect 389382 389898 424826 390134
rect 425062 389898 425146 390134
rect 425382 389898 460826 390134
rect 461062 389898 461146 390134
rect 461382 389898 496826 390134
rect 497062 389898 497146 390134
rect 497382 389898 532826 390134
rect 533062 389898 533146 390134
rect 533382 389898 568826 390134
rect 569062 389898 569146 390134
rect 569382 389898 591102 390134
rect 591338 389898 591422 390134
rect 591658 389898 592650 390134
rect -8726 389866 592650 389898
rect -8726 385954 592650 385986
rect -8726 385718 -6774 385954
rect -6538 385718 -6454 385954
rect -6218 385718 24326 385954
rect 24562 385718 24646 385954
rect 24882 385718 60326 385954
rect 60562 385718 60646 385954
rect 60882 385718 96326 385954
rect 96562 385718 96646 385954
rect 96882 385718 132326 385954
rect 132562 385718 132646 385954
rect 132882 385718 168326 385954
rect 168562 385718 168646 385954
rect 168882 385718 204326 385954
rect 204562 385718 204646 385954
rect 204882 385718 240326 385954
rect 240562 385718 240646 385954
rect 240882 385718 276326 385954
rect 276562 385718 276646 385954
rect 276882 385718 312326 385954
rect 312562 385718 312646 385954
rect 312882 385718 348326 385954
rect 348562 385718 348646 385954
rect 348882 385718 384326 385954
rect 384562 385718 384646 385954
rect 384882 385718 420326 385954
rect 420562 385718 420646 385954
rect 420882 385718 456326 385954
rect 456562 385718 456646 385954
rect 456882 385718 492326 385954
rect 492562 385718 492646 385954
rect 492882 385718 528326 385954
rect 528562 385718 528646 385954
rect 528882 385718 564326 385954
rect 564562 385718 564646 385954
rect 564882 385718 590142 385954
rect 590378 385718 590462 385954
rect 590698 385718 592650 385954
rect -8726 385634 592650 385718
rect -8726 385398 -6774 385634
rect -6538 385398 -6454 385634
rect -6218 385398 24326 385634
rect 24562 385398 24646 385634
rect 24882 385398 60326 385634
rect 60562 385398 60646 385634
rect 60882 385398 96326 385634
rect 96562 385398 96646 385634
rect 96882 385398 132326 385634
rect 132562 385398 132646 385634
rect 132882 385398 168326 385634
rect 168562 385398 168646 385634
rect 168882 385398 204326 385634
rect 204562 385398 204646 385634
rect 204882 385398 240326 385634
rect 240562 385398 240646 385634
rect 240882 385398 276326 385634
rect 276562 385398 276646 385634
rect 276882 385398 312326 385634
rect 312562 385398 312646 385634
rect 312882 385398 348326 385634
rect 348562 385398 348646 385634
rect 348882 385398 384326 385634
rect 384562 385398 384646 385634
rect 384882 385398 420326 385634
rect 420562 385398 420646 385634
rect 420882 385398 456326 385634
rect 456562 385398 456646 385634
rect 456882 385398 492326 385634
rect 492562 385398 492646 385634
rect 492882 385398 528326 385634
rect 528562 385398 528646 385634
rect 528882 385398 564326 385634
rect 564562 385398 564646 385634
rect 564882 385398 590142 385634
rect 590378 385398 590462 385634
rect 590698 385398 592650 385634
rect -8726 385366 592650 385398
rect -8726 381454 592650 381486
rect -8726 381218 -5814 381454
rect -5578 381218 -5494 381454
rect -5258 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 55826 381454
rect 56062 381218 56146 381454
rect 56382 381218 91826 381454
rect 92062 381218 92146 381454
rect 92382 381218 127826 381454
rect 128062 381218 128146 381454
rect 128382 381218 163826 381454
rect 164062 381218 164146 381454
rect 164382 381218 199826 381454
rect 200062 381218 200146 381454
rect 200382 381218 235826 381454
rect 236062 381218 236146 381454
rect 236382 381218 271826 381454
rect 272062 381218 272146 381454
rect 272382 381218 307826 381454
rect 308062 381218 308146 381454
rect 308382 381218 343826 381454
rect 344062 381218 344146 381454
rect 344382 381218 379826 381454
rect 380062 381218 380146 381454
rect 380382 381218 415826 381454
rect 416062 381218 416146 381454
rect 416382 381218 451826 381454
rect 452062 381218 452146 381454
rect 452382 381218 487826 381454
rect 488062 381218 488146 381454
rect 488382 381218 523826 381454
rect 524062 381218 524146 381454
rect 524382 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 589182 381454
rect 589418 381218 589502 381454
rect 589738 381218 592650 381454
rect -8726 381134 592650 381218
rect -8726 380898 -5814 381134
rect -5578 380898 -5494 381134
rect -5258 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 55826 381134
rect 56062 380898 56146 381134
rect 56382 380898 91826 381134
rect 92062 380898 92146 381134
rect 92382 380898 127826 381134
rect 128062 380898 128146 381134
rect 128382 380898 163826 381134
rect 164062 380898 164146 381134
rect 164382 380898 199826 381134
rect 200062 380898 200146 381134
rect 200382 380898 235826 381134
rect 236062 380898 236146 381134
rect 236382 380898 271826 381134
rect 272062 380898 272146 381134
rect 272382 380898 307826 381134
rect 308062 380898 308146 381134
rect 308382 380898 343826 381134
rect 344062 380898 344146 381134
rect 344382 380898 379826 381134
rect 380062 380898 380146 381134
rect 380382 380898 415826 381134
rect 416062 380898 416146 381134
rect 416382 380898 451826 381134
rect 452062 380898 452146 381134
rect 452382 380898 487826 381134
rect 488062 380898 488146 381134
rect 488382 380898 523826 381134
rect 524062 380898 524146 381134
rect 524382 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 589182 381134
rect 589418 380898 589502 381134
rect 589738 380898 592650 381134
rect -8726 380866 592650 380898
rect -8726 376954 592650 376986
rect -8726 376718 -4854 376954
rect -4618 376718 -4534 376954
rect -4298 376718 15326 376954
rect 15562 376718 15646 376954
rect 15882 376718 51326 376954
rect 51562 376718 51646 376954
rect 51882 376718 87326 376954
rect 87562 376718 87646 376954
rect 87882 376718 123326 376954
rect 123562 376718 123646 376954
rect 123882 376718 159326 376954
rect 159562 376718 159646 376954
rect 159882 376718 195326 376954
rect 195562 376718 195646 376954
rect 195882 376718 231326 376954
rect 231562 376718 231646 376954
rect 231882 376718 267326 376954
rect 267562 376718 267646 376954
rect 267882 376718 303326 376954
rect 303562 376718 303646 376954
rect 303882 376718 339326 376954
rect 339562 376718 339646 376954
rect 339882 376718 375326 376954
rect 375562 376718 375646 376954
rect 375882 376718 411326 376954
rect 411562 376718 411646 376954
rect 411882 376718 447326 376954
rect 447562 376718 447646 376954
rect 447882 376718 483326 376954
rect 483562 376718 483646 376954
rect 483882 376718 519326 376954
rect 519562 376718 519646 376954
rect 519882 376718 555326 376954
rect 555562 376718 555646 376954
rect 555882 376718 588222 376954
rect 588458 376718 588542 376954
rect 588778 376718 592650 376954
rect -8726 376634 592650 376718
rect -8726 376398 -4854 376634
rect -4618 376398 -4534 376634
rect -4298 376398 15326 376634
rect 15562 376398 15646 376634
rect 15882 376398 51326 376634
rect 51562 376398 51646 376634
rect 51882 376398 87326 376634
rect 87562 376398 87646 376634
rect 87882 376398 123326 376634
rect 123562 376398 123646 376634
rect 123882 376398 159326 376634
rect 159562 376398 159646 376634
rect 159882 376398 195326 376634
rect 195562 376398 195646 376634
rect 195882 376398 231326 376634
rect 231562 376398 231646 376634
rect 231882 376398 267326 376634
rect 267562 376398 267646 376634
rect 267882 376398 303326 376634
rect 303562 376398 303646 376634
rect 303882 376398 339326 376634
rect 339562 376398 339646 376634
rect 339882 376398 375326 376634
rect 375562 376398 375646 376634
rect 375882 376398 411326 376634
rect 411562 376398 411646 376634
rect 411882 376398 447326 376634
rect 447562 376398 447646 376634
rect 447882 376398 483326 376634
rect 483562 376398 483646 376634
rect 483882 376398 519326 376634
rect 519562 376398 519646 376634
rect 519882 376398 555326 376634
rect 555562 376398 555646 376634
rect 555882 376398 588222 376634
rect 588458 376398 588542 376634
rect 588778 376398 592650 376634
rect -8726 376366 592650 376398
rect -8726 372454 592650 372486
rect -8726 372218 -3894 372454
rect -3658 372218 -3574 372454
rect -3338 372218 10826 372454
rect 11062 372218 11146 372454
rect 11382 372218 46826 372454
rect 47062 372218 47146 372454
rect 47382 372218 82826 372454
rect 83062 372218 83146 372454
rect 83382 372218 118826 372454
rect 119062 372218 119146 372454
rect 119382 372218 154826 372454
rect 155062 372218 155146 372454
rect 155382 372218 190826 372454
rect 191062 372218 191146 372454
rect 191382 372218 226826 372454
rect 227062 372218 227146 372454
rect 227382 372218 262826 372454
rect 263062 372218 263146 372454
rect 263382 372218 298826 372454
rect 299062 372218 299146 372454
rect 299382 372218 334826 372454
rect 335062 372218 335146 372454
rect 335382 372218 370826 372454
rect 371062 372218 371146 372454
rect 371382 372218 406826 372454
rect 407062 372218 407146 372454
rect 407382 372218 442826 372454
rect 443062 372218 443146 372454
rect 443382 372218 478826 372454
rect 479062 372218 479146 372454
rect 479382 372218 514826 372454
rect 515062 372218 515146 372454
rect 515382 372218 550826 372454
rect 551062 372218 551146 372454
rect 551382 372218 587262 372454
rect 587498 372218 587582 372454
rect 587818 372218 592650 372454
rect -8726 372134 592650 372218
rect -8726 371898 -3894 372134
rect -3658 371898 -3574 372134
rect -3338 371898 10826 372134
rect 11062 371898 11146 372134
rect 11382 371898 46826 372134
rect 47062 371898 47146 372134
rect 47382 371898 82826 372134
rect 83062 371898 83146 372134
rect 83382 371898 118826 372134
rect 119062 371898 119146 372134
rect 119382 371898 154826 372134
rect 155062 371898 155146 372134
rect 155382 371898 190826 372134
rect 191062 371898 191146 372134
rect 191382 371898 226826 372134
rect 227062 371898 227146 372134
rect 227382 371898 262826 372134
rect 263062 371898 263146 372134
rect 263382 371898 298826 372134
rect 299062 371898 299146 372134
rect 299382 371898 334826 372134
rect 335062 371898 335146 372134
rect 335382 371898 370826 372134
rect 371062 371898 371146 372134
rect 371382 371898 406826 372134
rect 407062 371898 407146 372134
rect 407382 371898 442826 372134
rect 443062 371898 443146 372134
rect 443382 371898 478826 372134
rect 479062 371898 479146 372134
rect 479382 371898 514826 372134
rect 515062 371898 515146 372134
rect 515382 371898 550826 372134
rect 551062 371898 551146 372134
rect 551382 371898 587262 372134
rect 587498 371898 587582 372134
rect 587818 371898 592650 372134
rect -8726 371866 592650 371898
rect -8726 367954 592650 367986
rect -8726 367718 -2934 367954
rect -2698 367718 -2614 367954
rect -2378 367718 6326 367954
rect 6562 367718 6646 367954
rect 6882 367718 42326 367954
rect 42562 367718 42646 367954
rect 42882 367718 78326 367954
rect 78562 367718 78646 367954
rect 78882 367718 114326 367954
rect 114562 367718 114646 367954
rect 114882 367718 150326 367954
rect 150562 367718 150646 367954
rect 150882 367718 186326 367954
rect 186562 367718 186646 367954
rect 186882 367718 222326 367954
rect 222562 367718 222646 367954
rect 222882 367718 258326 367954
rect 258562 367718 258646 367954
rect 258882 367718 294326 367954
rect 294562 367718 294646 367954
rect 294882 367718 330326 367954
rect 330562 367718 330646 367954
rect 330882 367718 366326 367954
rect 366562 367718 366646 367954
rect 366882 367718 402326 367954
rect 402562 367718 402646 367954
rect 402882 367718 438326 367954
rect 438562 367718 438646 367954
rect 438882 367718 474326 367954
rect 474562 367718 474646 367954
rect 474882 367718 510326 367954
rect 510562 367718 510646 367954
rect 510882 367718 546326 367954
rect 546562 367718 546646 367954
rect 546882 367718 582326 367954
rect 582562 367718 582646 367954
rect 582882 367718 586302 367954
rect 586538 367718 586622 367954
rect 586858 367718 592650 367954
rect -8726 367634 592650 367718
rect -8726 367398 -2934 367634
rect -2698 367398 -2614 367634
rect -2378 367398 6326 367634
rect 6562 367398 6646 367634
rect 6882 367398 42326 367634
rect 42562 367398 42646 367634
rect 42882 367398 78326 367634
rect 78562 367398 78646 367634
rect 78882 367398 114326 367634
rect 114562 367398 114646 367634
rect 114882 367398 150326 367634
rect 150562 367398 150646 367634
rect 150882 367398 186326 367634
rect 186562 367398 186646 367634
rect 186882 367398 222326 367634
rect 222562 367398 222646 367634
rect 222882 367398 258326 367634
rect 258562 367398 258646 367634
rect 258882 367398 294326 367634
rect 294562 367398 294646 367634
rect 294882 367398 330326 367634
rect 330562 367398 330646 367634
rect 330882 367398 366326 367634
rect 366562 367398 366646 367634
rect 366882 367398 402326 367634
rect 402562 367398 402646 367634
rect 402882 367398 438326 367634
rect 438562 367398 438646 367634
rect 438882 367398 474326 367634
rect 474562 367398 474646 367634
rect 474882 367398 510326 367634
rect 510562 367398 510646 367634
rect 510882 367398 546326 367634
rect 546562 367398 546646 367634
rect 546882 367398 582326 367634
rect 582562 367398 582646 367634
rect 582882 367398 586302 367634
rect 586538 367398 586622 367634
rect 586858 367398 592650 367634
rect -8726 367366 592650 367398
rect -8726 363454 592650 363486
rect -8726 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 73826 363454
rect 74062 363218 74146 363454
rect 74382 363218 109826 363454
rect 110062 363218 110146 363454
rect 110382 363218 145826 363454
rect 146062 363218 146146 363454
rect 146382 363218 181826 363454
rect 182062 363218 182146 363454
rect 182382 363218 217826 363454
rect 218062 363218 218146 363454
rect 218382 363218 253826 363454
rect 254062 363218 254146 363454
rect 254382 363218 289826 363454
rect 290062 363218 290146 363454
rect 290382 363218 325826 363454
rect 326062 363218 326146 363454
rect 326382 363218 361826 363454
rect 362062 363218 362146 363454
rect 362382 363218 397826 363454
rect 398062 363218 398146 363454
rect 398382 363218 433826 363454
rect 434062 363218 434146 363454
rect 434382 363218 469826 363454
rect 470062 363218 470146 363454
rect 470382 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 592650 363454
rect -8726 363134 592650 363218
rect -8726 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 73826 363134
rect 74062 362898 74146 363134
rect 74382 362898 109826 363134
rect 110062 362898 110146 363134
rect 110382 362898 145826 363134
rect 146062 362898 146146 363134
rect 146382 362898 181826 363134
rect 182062 362898 182146 363134
rect 182382 362898 217826 363134
rect 218062 362898 218146 363134
rect 218382 362898 253826 363134
rect 254062 362898 254146 363134
rect 254382 362898 289826 363134
rect 290062 362898 290146 363134
rect 290382 362898 325826 363134
rect 326062 362898 326146 363134
rect 326382 362898 361826 363134
rect 362062 362898 362146 363134
rect 362382 362898 397826 363134
rect 398062 362898 398146 363134
rect 398382 362898 433826 363134
rect 434062 362898 434146 363134
rect 434382 362898 469826 363134
rect 470062 362898 470146 363134
rect 470382 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 592650 363134
rect -8726 362866 592650 362898
rect -8726 358954 592650 358986
rect -8726 358718 -8694 358954
rect -8458 358718 -8374 358954
rect -8138 358718 33326 358954
rect 33562 358718 33646 358954
rect 33882 358718 69326 358954
rect 69562 358718 69646 358954
rect 69882 358718 105326 358954
rect 105562 358718 105646 358954
rect 105882 358718 141326 358954
rect 141562 358718 141646 358954
rect 141882 358718 177326 358954
rect 177562 358718 177646 358954
rect 177882 358718 213326 358954
rect 213562 358718 213646 358954
rect 213882 358718 249326 358954
rect 249562 358718 249646 358954
rect 249882 358718 285326 358954
rect 285562 358718 285646 358954
rect 285882 358718 321326 358954
rect 321562 358718 321646 358954
rect 321882 358718 357326 358954
rect 357562 358718 357646 358954
rect 357882 358718 393326 358954
rect 393562 358718 393646 358954
rect 393882 358718 429326 358954
rect 429562 358718 429646 358954
rect 429882 358718 465326 358954
rect 465562 358718 465646 358954
rect 465882 358718 501326 358954
rect 501562 358718 501646 358954
rect 501882 358718 537326 358954
rect 537562 358718 537646 358954
rect 537882 358718 573326 358954
rect 573562 358718 573646 358954
rect 573882 358718 592062 358954
rect 592298 358718 592382 358954
rect 592618 358718 592650 358954
rect -8726 358634 592650 358718
rect -8726 358398 -8694 358634
rect -8458 358398 -8374 358634
rect -8138 358398 33326 358634
rect 33562 358398 33646 358634
rect 33882 358398 69326 358634
rect 69562 358398 69646 358634
rect 69882 358398 105326 358634
rect 105562 358398 105646 358634
rect 105882 358398 141326 358634
rect 141562 358398 141646 358634
rect 141882 358398 177326 358634
rect 177562 358398 177646 358634
rect 177882 358398 213326 358634
rect 213562 358398 213646 358634
rect 213882 358398 249326 358634
rect 249562 358398 249646 358634
rect 249882 358398 285326 358634
rect 285562 358398 285646 358634
rect 285882 358398 321326 358634
rect 321562 358398 321646 358634
rect 321882 358398 357326 358634
rect 357562 358398 357646 358634
rect 357882 358398 393326 358634
rect 393562 358398 393646 358634
rect 393882 358398 429326 358634
rect 429562 358398 429646 358634
rect 429882 358398 465326 358634
rect 465562 358398 465646 358634
rect 465882 358398 501326 358634
rect 501562 358398 501646 358634
rect 501882 358398 537326 358634
rect 537562 358398 537646 358634
rect 537882 358398 573326 358634
rect 573562 358398 573646 358634
rect 573882 358398 592062 358634
rect 592298 358398 592382 358634
rect 592618 358398 592650 358634
rect -8726 358366 592650 358398
rect -8726 354454 592650 354486
rect -8726 354218 -7734 354454
rect -7498 354218 -7414 354454
rect -7178 354218 28826 354454
rect 29062 354218 29146 354454
rect 29382 354218 64826 354454
rect 65062 354218 65146 354454
rect 65382 354218 100826 354454
rect 101062 354218 101146 354454
rect 101382 354218 136826 354454
rect 137062 354218 137146 354454
rect 137382 354218 172826 354454
rect 173062 354218 173146 354454
rect 173382 354218 208826 354454
rect 209062 354218 209146 354454
rect 209382 354218 244826 354454
rect 245062 354218 245146 354454
rect 245382 354218 280826 354454
rect 281062 354218 281146 354454
rect 281382 354218 316826 354454
rect 317062 354218 317146 354454
rect 317382 354218 352826 354454
rect 353062 354218 353146 354454
rect 353382 354218 388826 354454
rect 389062 354218 389146 354454
rect 389382 354218 424826 354454
rect 425062 354218 425146 354454
rect 425382 354218 460826 354454
rect 461062 354218 461146 354454
rect 461382 354218 496826 354454
rect 497062 354218 497146 354454
rect 497382 354218 532826 354454
rect 533062 354218 533146 354454
rect 533382 354218 568826 354454
rect 569062 354218 569146 354454
rect 569382 354218 591102 354454
rect 591338 354218 591422 354454
rect 591658 354218 592650 354454
rect -8726 354134 592650 354218
rect -8726 353898 -7734 354134
rect -7498 353898 -7414 354134
rect -7178 353898 28826 354134
rect 29062 353898 29146 354134
rect 29382 353898 64826 354134
rect 65062 353898 65146 354134
rect 65382 353898 100826 354134
rect 101062 353898 101146 354134
rect 101382 353898 136826 354134
rect 137062 353898 137146 354134
rect 137382 353898 172826 354134
rect 173062 353898 173146 354134
rect 173382 353898 208826 354134
rect 209062 353898 209146 354134
rect 209382 353898 244826 354134
rect 245062 353898 245146 354134
rect 245382 353898 280826 354134
rect 281062 353898 281146 354134
rect 281382 353898 316826 354134
rect 317062 353898 317146 354134
rect 317382 353898 352826 354134
rect 353062 353898 353146 354134
rect 353382 353898 388826 354134
rect 389062 353898 389146 354134
rect 389382 353898 424826 354134
rect 425062 353898 425146 354134
rect 425382 353898 460826 354134
rect 461062 353898 461146 354134
rect 461382 353898 496826 354134
rect 497062 353898 497146 354134
rect 497382 353898 532826 354134
rect 533062 353898 533146 354134
rect 533382 353898 568826 354134
rect 569062 353898 569146 354134
rect 569382 353898 591102 354134
rect 591338 353898 591422 354134
rect 591658 353898 592650 354134
rect -8726 353866 592650 353898
rect -8726 349954 592650 349986
rect -8726 349718 -6774 349954
rect -6538 349718 -6454 349954
rect -6218 349718 24326 349954
rect 24562 349718 24646 349954
rect 24882 349718 60326 349954
rect 60562 349718 60646 349954
rect 60882 349718 96326 349954
rect 96562 349718 96646 349954
rect 96882 349718 132326 349954
rect 132562 349718 132646 349954
rect 132882 349718 168326 349954
rect 168562 349718 168646 349954
rect 168882 349718 204326 349954
rect 204562 349718 204646 349954
rect 204882 349718 240326 349954
rect 240562 349718 240646 349954
rect 240882 349718 276326 349954
rect 276562 349718 276646 349954
rect 276882 349718 312326 349954
rect 312562 349718 312646 349954
rect 312882 349718 348326 349954
rect 348562 349718 348646 349954
rect 348882 349718 384326 349954
rect 384562 349718 384646 349954
rect 384882 349718 420326 349954
rect 420562 349718 420646 349954
rect 420882 349718 456326 349954
rect 456562 349718 456646 349954
rect 456882 349718 492326 349954
rect 492562 349718 492646 349954
rect 492882 349718 528326 349954
rect 528562 349718 528646 349954
rect 528882 349718 564326 349954
rect 564562 349718 564646 349954
rect 564882 349718 590142 349954
rect 590378 349718 590462 349954
rect 590698 349718 592650 349954
rect -8726 349634 592650 349718
rect -8726 349398 -6774 349634
rect -6538 349398 -6454 349634
rect -6218 349398 24326 349634
rect 24562 349398 24646 349634
rect 24882 349398 60326 349634
rect 60562 349398 60646 349634
rect 60882 349398 96326 349634
rect 96562 349398 96646 349634
rect 96882 349398 132326 349634
rect 132562 349398 132646 349634
rect 132882 349398 168326 349634
rect 168562 349398 168646 349634
rect 168882 349398 204326 349634
rect 204562 349398 204646 349634
rect 204882 349398 240326 349634
rect 240562 349398 240646 349634
rect 240882 349398 276326 349634
rect 276562 349398 276646 349634
rect 276882 349398 312326 349634
rect 312562 349398 312646 349634
rect 312882 349398 348326 349634
rect 348562 349398 348646 349634
rect 348882 349398 384326 349634
rect 384562 349398 384646 349634
rect 384882 349398 420326 349634
rect 420562 349398 420646 349634
rect 420882 349398 456326 349634
rect 456562 349398 456646 349634
rect 456882 349398 492326 349634
rect 492562 349398 492646 349634
rect 492882 349398 528326 349634
rect 528562 349398 528646 349634
rect 528882 349398 564326 349634
rect 564562 349398 564646 349634
rect 564882 349398 590142 349634
rect 590378 349398 590462 349634
rect 590698 349398 592650 349634
rect -8726 349366 592650 349398
rect -8726 345454 592650 345486
rect -8726 345218 -5814 345454
rect -5578 345218 -5494 345454
rect -5258 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 55826 345454
rect 56062 345218 56146 345454
rect 56382 345218 91826 345454
rect 92062 345218 92146 345454
rect 92382 345218 127826 345454
rect 128062 345218 128146 345454
rect 128382 345218 163826 345454
rect 164062 345218 164146 345454
rect 164382 345218 199826 345454
rect 200062 345218 200146 345454
rect 200382 345218 235826 345454
rect 236062 345218 236146 345454
rect 236382 345218 271826 345454
rect 272062 345218 272146 345454
rect 272382 345218 307826 345454
rect 308062 345218 308146 345454
rect 308382 345218 343826 345454
rect 344062 345218 344146 345454
rect 344382 345218 379826 345454
rect 380062 345218 380146 345454
rect 380382 345218 415826 345454
rect 416062 345218 416146 345454
rect 416382 345218 451826 345454
rect 452062 345218 452146 345454
rect 452382 345218 487826 345454
rect 488062 345218 488146 345454
rect 488382 345218 523826 345454
rect 524062 345218 524146 345454
rect 524382 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 589182 345454
rect 589418 345218 589502 345454
rect 589738 345218 592650 345454
rect -8726 345134 592650 345218
rect -8726 344898 -5814 345134
rect -5578 344898 -5494 345134
rect -5258 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 55826 345134
rect 56062 344898 56146 345134
rect 56382 344898 91826 345134
rect 92062 344898 92146 345134
rect 92382 344898 127826 345134
rect 128062 344898 128146 345134
rect 128382 344898 163826 345134
rect 164062 344898 164146 345134
rect 164382 344898 199826 345134
rect 200062 344898 200146 345134
rect 200382 344898 235826 345134
rect 236062 344898 236146 345134
rect 236382 344898 271826 345134
rect 272062 344898 272146 345134
rect 272382 344898 307826 345134
rect 308062 344898 308146 345134
rect 308382 344898 343826 345134
rect 344062 344898 344146 345134
rect 344382 344898 379826 345134
rect 380062 344898 380146 345134
rect 380382 344898 415826 345134
rect 416062 344898 416146 345134
rect 416382 344898 451826 345134
rect 452062 344898 452146 345134
rect 452382 344898 487826 345134
rect 488062 344898 488146 345134
rect 488382 344898 523826 345134
rect 524062 344898 524146 345134
rect 524382 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 589182 345134
rect 589418 344898 589502 345134
rect 589738 344898 592650 345134
rect -8726 344866 592650 344898
rect -8726 340954 592650 340986
rect -8726 340718 -4854 340954
rect -4618 340718 -4534 340954
rect -4298 340718 15326 340954
rect 15562 340718 15646 340954
rect 15882 340718 51326 340954
rect 51562 340718 51646 340954
rect 51882 340718 87326 340954
rect 87562 340718 87646 340954
rect 87882 340718 123326 340954
rect 123562 340718 123646 340954
rect 123882 340718 159326 340954
rect 159562 340718 159646 340954
rect 159882 340718 195326 340954
rect 195562 340718 195646 340954
rect 195882 340718 231326 340954
rect 231562 340718 231646 340954
rect 231882 340718 267326 340954
rect 267562 340718 267646 340954
rect 267882 340718 303326 340954
rect 303562 340718 303646 340954
rect 303882 340718 339326 340954
rect 339562 340718 339646 340954
rect 339882 340718 375326 340954
rect 375562 340718 375646 340954
rect 375882 340718 411326 340954
rect 411562 340718 411646 340954
rect 411882 340718 447326 340954
rect 447562 340718 447646 340954
rect 447882 340718 483326 340954
rect 483562 340718 483646 340954
rect 483882 340718 519326 340954
rect 519562 340718 519646 340954
rect 519882 340718 555326 340954
rect 555562 340718 555646 340954
rect 555882 340718 588222 340954
rect 588458 340718 588542 340954
rect 588778 340718 592650 340954
rect -8726 340634 592650 340718
rect -8726 340398 -4854 340634
rect -4618 340398 -4534 340634
rect -4298 340398 15326 340634
rect 15562 340398 15646 340634
rect 15882 340398 51326 340634
rect 51562 340398 51646 340634
rect 51882 340398 87326 340634
rect 87562 340398 87646 340634
rect 87882 340398 123326 340634
rect 123562 340398 123646 340634
rect 123882 340398 159326 340634
rect 159562 340398 159646 340634
rect 159882 340398 195326 340634
rect 195562 340398 195646 340634
rect 195882 340398 231326 340634
rect 231562 340398 231646 340634
rect 231882 340398 267326 340634
rect 267562 340398 267646 340634
rect 267882 340398 303326 340634
rect 303562 340398 303646 340634
rect 303882 340398 339326 340634
rect 339562 340398 339646 340634
rect 339882 340398 375326 340634
rect 375562 340398 375646 340634
rect 375882 340398 411326 340634
rect 411562 340398 411646 340634
rect 411882 340398 447326 340634
rect 447562 340398 447646 340634
rect 447882 340398 483326 340634
rect 483562 340398 483646 340634
rect 483882 340398 519326 340634
rect 519562 340398 519646 340634
rect 519882 340398 555326 340634
rect 555562 340398 555646 340634
rect 555882 340398 588222 340634
rect 588458 340398 588542 340634
rect 588778 340398 592650 340634
rect -8726 340366 592650 340398
rect -8726 336454 592650 336486
rect -8726 336218 -3894 336454
rect -3658 336218 -3574 336454
rect -3338 336218 10826 336454
rect 11062 336218 11146 336454
rect 11382 336218 46826 336454
rect 47062 336218 47146 336454
rect 47382 336218 82826 336454
rect 83062 336218 83146 336454
rect 83382 336218 118826 336454
rect 119062 336218 119146 336454
rect 119382 336218 154826 336454
rect 155062 336218 155146 336454
rect 155382 336218 190826 336454
rect 191062 336218 191146 336454
rect 191382 336218 226826 336454
rect 227062 336218 227146 336454
rect 227382 336218 262826 336454
rect 263062 336218 263146 336454
rect 263382 336218 298826 336454
rect 299062 336218 299146 336454
rect 299382 336218 334826 336454
rect 335062 336218 335146 336454
rect 335382 336218 370826 336454
rect 371062 336218 371146 336454
rect 371382 336218 406826 336454
rect 407062 336218 407146 336454
rect 407382 336218 442826 336454
rect 443062 336218 443146 336454
rect 443382 336218 478826 336454
rect 479062 336218 479146 336454
rect 479382 336218 514826 336454
rect 515062 336218 515146 336454
rect 515382 336218 550826 336454
rect 551062 336218 551146 336454
rect 551382 336218 587262 336454
rect 587498 336218 587582 336454
rect 587818 336218 592650 336454
rect -8726 336134 592650 336218
rect -8726 335898 -3894 336134
rect -3658 335898 -3574 336134
rect -3338 335898 10826 336134
rect 11062 335898 11146 336134
rect 11382 335898 46826 336134
rect 47062 335898 47146 336134
rect 47382 335898 82826 336134
rect 83062 335898 83146 336134
rect 83382 335898 118826 336134
rect 119062 335898 119146 336134
rect 119382 335898 154826 336134
rect 155062 335898 155146 336134
rect 155382 335898 190826 336134
rect 191062 335898 191146 336134
rect 191382 335898 226826 336134
rect 227062 335898 227146 336134
rect 227382 335898 262826 336134
rect 263062 335898 263146 336134
rect 263382 335898 298826 336134
rect 299062 335898 299146 336134
rect 299382 335898 334826 336134
rect 335062 335898 335146 336134
rect 335382 335898 370826 336134
rect 371062 335898 371146 336134
rect 371382 335898 406826 336134
rect 407062 335898 407146 336134
rect 407382 335898 442826 336134
rect 443062 335898 443146 336134
rect 443382 335898 478826 336134
rect 479062 335898 479146 336134
rect 479382 335898 514826 336134
rect 515062 335898 515146 336134
rect 515382 335898 550826 336134
rect 551062 335898 551146 336134
rect 551382 335898 587262 336134
rect 587498 335898 587582 336134
rect 587818 335898 592650 336134
rect -8726 335866 592650 335898
rect -8726 331954 592650 331986
rect -8726 331718 -2934 331954
rect -2698 331718 -2614 331954
rect -2378 331718 6326 331954
rect 6562 331718 6646 331954
rect 6882 331718 42326 331954
rect 42562 331718 42646 331954
rect 42882 331718 78326 331954
rect 78562 331718 78646 331954
rect 78882 331718 114326 331954
rect 114562 331718 114646 331954
rect 114882 331718 150326 331954
rect 150562 331718 150646 331954
rect 150882 331718 186326 331954
rect 186562 331718 186646 331954
rect 186882 331718 222326 331954
rect 222562 331718 222646 331954
rect 222882 331718 258326 331954
rect 258562 331718 258646 331954
rect 258882 331718 294326 331954
rect 294562 331718 294646 331954
rect 294882 331718 330326 331954
rect 330562 331718 330646 331954
rect 330882 331718 366326 331954
rect 366562 331718 366646 331954
rect 366882 331718 402326 331954
rect 402562 331718 402646 331954
rect 402882 331718 438326 331954
rect 438562 331718 438646 331954
rect 438882 331718 474326 331954
rect 474562 331718 474646 331954
rect 474882 331718 510326 331954
rect 510562 331718 510646 331954
rect 510882 331718 546326 331954
rect 546562 331718 546646 331954
rect 546882 331718 582326 331954
rect 582562 331718 582646 331954
rect 582882 331718 586302 331954
rect 586538 331718 586622 331954
rect 586858 331718 592650 331954
rect -8726 331634 592650 331718
rect -8726 331398 -2934 331634
rect -2698 331398 -2614 331634
rect -2378 331398 6326 331634
rect 6562 331398 6646 331634
rect 6882 331398 42326 331634
rect 42562 331398 42646 331634
rect 42882 331398 78326 331634
rect 78562 331398 78646 331634
rect 78882 331398 114326 331634
rect 114562 331398 114646 331634
rect 114882 331398 150326 331634
rect 150562 331398 150646 331634
rect 150882 331398 186326 331634
rect 186562 331398 186646 331634
rect 186882 331398 222326 331634
rect 222562 331398 222646 331634
rect 222882 331398 258326 331634
rect 258562 331398 258646 331634
rect 258882 331398 294326 331634
rect 294562 331398 294646 331634
rect 294882 331398 330326 331634
rect 330562 331398 330646 331634
rect 330882 331398 366326 331634
rect 366562 331398 366646 331634
rect 366882 331398 402326 331634
rect 402562 331398 402646 331634
rect 402882 331398 438326 331634
rect 438562 331398 438646 331634
rect 438882 331398 474326 331634
rect 474562 331398 474646 331634
rect 474882 331398 510326 331634
rect 510562 331398 510646 331634
rect 510882 331398 546326 331634
rect 546562 331398 546646 331634
rect 546882 331398 582326 331634
rect 582562 331398 582646 331634
rect 582882 331398 586302 331634
rect 586538 331398 586622 331634
rect 586858 331398 592650 331634
rect -8726 331366 592650 331398
rect -8726 327454 592650 327486
rect -8726 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 73826 327454
rect 74062 327218 74146 327454
rect 74382 327218 109826 327454
rect 110062 327218 110146 327454
rect 110382 327218 145826 327454
rect 146062 327218 146146 327454
rect 146382 327218 181826 327454
rect 182062 327218 182146 327454
rect 182382 327218 217826 327454
rect 218062 327218 218146 327454
rect 218382 327218 253826 327454
rect 254062 327218 254146 327454
rect 254382 327218 289826 327454
rect 290062 327218 290146 327454
rect 290382 327218 325826 327454
rect 326062 327218 326146 327454
rect 326382 327218 361826 327454
rect 362062 327218 362146 327454
rect 362382 327218 397826 327454
rect 398062 327218 398146 327454
rect 398382 327218 433826 327454
rect 434062 327218 434146 327454
rect 434382 327218 469826 327454
rect 470062 327218 470146 327454
rect 470382 327218 505826 327454
rect 506062 327218 506146 327454
rect 506382 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 592650 327454
rect -8726 327134 592650 327218
rect -8726 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 73826 327134
rect 74062 326898 74146 327134
rect 74382 326898 109826 327134
rect 110062 326898 110146 327134
rect 110382 326898 145826 327134
rect 146062 326898 146146 327134
rect 146382 326898 181826 327134
rect 182062 326898 182146 327134
rect 182382 326898 217826 327134
rect 218062 326898 218146 327134
rect 218382 326898 253826 327134
rect 254062 326898 254146 327134
rect 254382 326898 289826 327134
rect 290062 326898 290146 327134
rect 290382 326898 325826 327134
rect 326062 326898 326146 327134
rect 326382 326898 361826 327134
rect 362062 326898 362146 327134
rect 362382 326898 397826 327134
rect 398062 326898 398146 327134
rect 398382 326898 433826 327134
rect 434062 326898 434146 327134
rect 434382 326898 469826 327134
rect 470062 326898 470146 327134
rect 470382 326898 505826 327134
rect 506062 326898 506146 327134
rect 506382 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 592650 327134
rect -8726 326866 592650 326898
rect -8726 322954 592650 322986
rect -8726 322718 -8694 322954
rect -8458 322718 -8374 322954
rect -8138 322718 33326 322954
rect 33562 322718 33646 322954
rect 33882 322718 69326 322954
rect 69562 322718 69646 322954
rect 69882 322718 105326 322954
rect 105562 322718 105646 322954
rect 105882 322718 141326 322954
rect 141562 322718 141646 322954
rect 141882 322718 177326 322954
rect 177562 322718 177646 322954
rect 177882 322718 213326 322954
rect 213562 322718 213646 322954
rect 213882 322718 249326 322954
rect 249562 322718 249646 322954
rect 249882 322718 285326 322954
rect 285562 322718 285646 322954
rect 285882 322718 321326 322954
rect 321562 322718 321646 322954
rect 321882 322718 357326 322954
rect 357562 322718 357646 322954
rect 357882 322718 393326 322954
rect 393562 322718 393646 322954
rect 393882 322718 429326 322954
rect 429562 322718 429646 322954
rect 429882 322718 465326 322954
rect 465562 322718 465646 322954
rect 465882 322718 501326 322954
rect 501562 322718 501646 322954
rect 501882 322718 537326 322954
rect 537562 322718 537646 322954
rect 537882 322718 573326 322954
rect 573562 322718 573646 322954
rect 573882 322718 592062 322954
rect 592298 322718 592382 322954
rect 592618 322718 592650 322954
rect -8726 322634 592650 322718
rect -8726 322398 -8694 322634
rect -8458 322398 -8374 322634
rect -8138 322398 33326 322634
rect 33562 322398 33646 322634
rect 33882 322398 69326 322634
rect 69562 322398 69646 322634
rect 69882 322398 105326 322634
rect 105562 322398 105646 322634
rect 105882 322398 141326 322634
rect 141562 322398 141646 322634
rect 141882 322398 177326 322634
rect 177562 322398 177646 322634
rect 177882 322398 213326 322634
rect 213562 322398 213646 322634
rect 213882 322398 249326 322634
rect 249562 322398 249646 322634
rect 249882 322398 285326 322634
rect 285562 322398 285646 322634
rect 285882 322398 321326 322634
rect 321562 322398 321646 322634
rect 321882 322398 357326 322634
rect 357562 322398 357646 322634
rect 357882 322398 393326 322634
rect 393562 322398 393646 322634
rect 393882 322398 429326 322634
rect 429562 322398 429646 322634
rect 429882 322398 465326 322634
rect 465562 322398 465646 322634
rect 465882 322398 501326 322634
rect 501562 322398 501646 322634
rect 501882 322398 537326 322634
rect 537562 322398 537646 322634
rect 537882 322398 573326 322634
rect 573562 322398 573646 322634
rect 573882 322398 592062 322634
rect 592298 322398 592382 322634
rect 592618 322398 592650 322634
rect -8726 322366 592650 322398
rect -8726 318454 592650 318486
rect -8726 318218 -7734 318454
rect -7498 318218 -7414 318454
rect -7178 318218 28826 318454
rect 29062 318218 29146 318454
rect 29382 318218 64826 318454
rect 65062 318218 65146 318454
rect 65382 318218 100826 318454
rect 101062 318218 101146 318454
rect 101382 318218 136826 318454
rect 137062 318218 137146 318454
rect 137382 318218 172826 318454
rect 173062 318218 173146 318454
rect 173382 318218 208826 318454
rect 209062 318218 209146 318454
rect 209382 318218 244826 318454
rect 245062 318218 245146 318454
rect 245382 318218 280826 318454
rect 281062 318218 281146 318454
rect 281382 318218 316826 318454
rect 317062 318218 317146 318454
rect 317382 318218 352826 318454
rect 353062 318218 353146 318454
rect 353382 318218 388826 318454
rect 389062 318218 389146 318454
rect 389382 318218 424826 318454
rect 425062 318218 425146 318454
rect 425382 318218 460826 318454
rect 461062 318218 461146 318454
rect 461382 318218 496826 318454
rect 497062 318218 497146 318454
rect 497382 318218 532826 318454
rect 533062 318218 533146 318454
rect 533382 318218 568826 318454
rect 569062 318218 569146 318454
rect 569382 318218 591102 318454
rect 591338 318218 591422 318454
rect 591658 318218 592650 318454
rect -8726 318134 592650 318218
rect -8726 317898 -7734 318134
rect -7498 317898 -7414 318134
rect -7178 317898 28826 318134
rect 29062 317898 29146 318134
rect 29382 317898 64826 318134
rect 65062 317898 65146 318134
rect 65382 317898 100826 318134
rect 101062 317898 101146 318134
rect 101382 317898 136826 318134
rect 137062 317898 137146 318134
rect 137382 317898 172826 318134
rect 173062 317898 173146 318134
rect 173382 317898 208826 318134
rect 209062 317898 209146 318134
rect 209382 317898 244826 318134
rect 245062 317898 245146 318134
rect 245382 317898 280826 318134
rect 281062 317898 281146 318134
rect 281382 317898 316826 318134
rect 317062 317898 317146 318134
rect 317382 317898 352826 318134
rect 353062 317898 353146 318134
rect 353382 317898 388826 318134
rect 389062 317898 389146 318134
rect 389382 317898 424826 318134
rect 425062 317898 425146 318134
rect 425382 317898 460826 318134
rect 461062 317898 461146 318134
rect 461382 317898 496826 318134
rect 497062 317898 497146 318134
rect 497382 317898 532826 318134
rect 533062 317898 533146 318134
rect 533382 317898 568826 318134
rect 569062 317898 569146 318134
rect 569382 317898 591102 318134
rect 591338 317898 591422 318134
rect 591658 317898 592650 318134
rect -8726 317866 592650 317898
rect -8726 313954 592650 313986
rect -8726 313718 -6774 313954
rect -6538 313718 -6454 313954
rect -6218 313718 24326 313954
rect 24562 313718 24646 313954
rect 24882 313718 60326 313954
rect 60562 313718 60646 313954
rect 60882 313718 96326 313954
rect 96562 313718 96646 313954
rect 96882 313718 132326 313954
rect 132562 313718 132646 313954
rect 132882 313718 168326 313954
rect 168562 313718 168646 313954
rect 168882 313718 204326 313954
rect 204562 313718 204646 313954
rect 204882 313718 240326 313954
rect 240562 313718 240646 313954
rect 240882 313718 276326 313954
rect 276562 313718 276646 313954
rect 276882 313718 312326 313954
rect 312562 313718 312646 313954
rect 312882 313718 348326 313954
rect 348562 313718 348646 313954
rect 348882 313718 384326 313954
rect 384562 313718 384646 313954
rect 384882 313718 420326 313954
rect 420562 313718 420646 313954
rect 420882 313718 456326 313954
rect 456562 313718 456646 313954
rect 456882 313718 492326 313954
rect 492562 313718 492646 313954
rect 492882 313718 528326 313954
rect 528562 313718 528646 313954
rect 528882 313718 564326 313954
rect 564562 313718 564646 313954
rect 564882 313718 590142 313954
rect 590378 313718 590462 313954
rect 590698 313718 592650 313954
rect -8726 313634 592650 313718
rect -8726 313398 -6774 313634
rect -6538 313398 -6454 313634
rect -6218 313398 24326 313634
rect 24562 313398 24646 313634
rect 24882 313398 60326 313634
rect 60562 313398 60646 313634
rect 60882 313398 96326 313634
rect 96562 313398 96646 313634
rect 96882 313398 132326 313634
rect 132562 313398 132646 313634
rect 132882 313398 168326 313634
rect 168562 313398 168646 313634
rect 168882 313398 204326 313634
rect 204562 313398 204646 313634
rect 204882 313398 240326 313634
rect 240562 313398 240646 313634
rect 240882 313398 276326 313634
rect 276562 313398 276646 313634
rect 276882 313398 312326 313634
rect 312562 313398 312646 313634
rect 312882 313398 348326 313634
rect 348562 313398 348646 313634
rect 348882 313398 384326 313634
rect 384562 313398 384646 313634
rect 384882 313398 420326 313634
rect 420562 313398 420646 313634
rect 420882 313398 456326 313634
rect 456562 313398 456646 313634
rect 456882 313398 492326 313634
rect 492562 313398 492646 313634
rect 492882 313398 528326 313634
rect 528562 313398 528646 313634
rect 528882 313398 564326 313634
rect 564562 313398 564646 313634
rect 564882 313398 590142 313634
rect 590378 313398 590462 313634
rect 590698 313398 592650 313634
rect -8726 313366 592650 313398
rect -8726 309454 592650 309486
rect -8726 309218 -5814 309454
rect -5578 309218 -5494 309454
rect -5258 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 55826 309454
rect 56062 309218 56146 309454
rect 56382 309218 91826 309454
rect 92062 309218 92146 309454
rect 92382 309218 127826 309454
rect 128062 309218 128146 309454
rect 128382 309218 163826 309454
rect 164062 309218 164146 309454
rect 164382 309218 199826 309454
rect 200062 309218 200146 309454
rect 200382 309218 235826 309454
rect 236062 309218 236146 309454
rect 236382 309218 271826 309454
rect 272062 309218 272146 309454
rect 272382 309218 307826 309454
rect 308062 309218 308146 309454
rect 308382 309218 343826 309454
rect 344062 309218 344146 309454
rect 344382 309218 379826 309454
rect 380062 309218 380146 309454
rect 380382 309218 415826 309454
rect 416062 309218 416146 309454
rect 416382 309218 451826 309454
rect 452062 309218 452146 309454
rect 452382 309218 487826 309454
rect 488062 309218 488146 309454
rect 488382 309218 523826 309454
rect 524062 309218 524146 309454
rect 524382 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 589182 309454
rect 589418 309218 589502 309454
rect 589738 309218 592650 309454
rect -8726 309134 592650 309218
rect -8726 308898 -5814 309134
rect -5578 308898 -5494 309134
rect -5258 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 55826 309134
rect 56062 308898 56146 309134
rect 56382 308898 91826 309134
rect 92062 308898 92146 309134
rect 92382 308898 127826 309134
rect 128062 308898 128146 309134
rect 128382 308898 163826 309134
rect 164062 308898 164146 309134
rect 164382 308898 199826 309134
rect 200062 308898 200146 309134
rect 200382 308898 235826 309134
rect 236062 308898 236146 309134
rect 236382 308898 271826 309134
rect 272062 308898 272146 309134
rect 272382 308898 307826 309134
rect 308062 308898 308146 309134
rect 308382 308898 343826 309134
rect 344062 308898 344146 309134
rect 344382 308898 379826 309134
rect 380062 308898 380146 309134
rect 380382 308898 415826 309134
rect 416062 308898 416146 309134
rect 416382 308898 451826 309134
rect 452062 308898 452146 309134
rect 452382 308898 487826 309134
rect 488062 308898 488146 309134
rect 488382 308898 523826 309134
rect 524062 308898 524146 309134
rect 524382 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 589182 309134
rect 589418 308898 589502 309134
rect 589738 308898 592650 309134
rect -8726 308866 592650 308898
rect -8726 304954 592650 304986
rect -8726 304718 -4854 304954
rect -4618 304718 -4534 304954
rect -4298 304718 15326 304954
rect 15562 304718 15646 304954
rect 15882 304718 51326 304954
rect 51562 304718 51646 304954
rect 51882 304718 87326 304954
rect 87562 304718 87646 304954
rect 87882 304718 123326 304954
rect 123562 304718 123646 304954
rect 123882 304718 159326 304954
rect 159562 304718 159646 304954
rect 159882 304718 195326 304954
rect 195562 304718 195646 304954
rect 195882 304718 231326 304954
rect 231562 304718 231646 304954
rect 231882 304718 267326 304954
rect 267562 304718 267646 304954
rect 267882 304718 303326 304954
rect 303562 304718 303646 304954
rect 303882 304718 339326 304954
rect 339562 304718 339646 304954
rect 339882 304718 375326 304954
rect 375562 304718 375646 304954
rect 375882 304718 411326 304954
rect 411562 304718 411646 304954
rect 411882 304718 447326 304954
rect 447562 304718 447646 304954
rect 447882 304718 483326 304954
rect 483562 304718 483646 304954
rect 483882 304718 519326 304954
rect 519562 304718 519646 304954
rect 519882 304718 555326 304954
rect 555562 304718 555646 304954
rect 555882 304718 588222 304954
rect 588458 304718 588542 304954
rect 588778 304718 592650 304954
rect -8726 304634 592650 304718
rect -8726 304398 -4854 304634
rect -4618 304398 -4534 304634
rect -4298 304398 15326 304634
rect 15562 304398 15646 304634
rect 15882 304398 51326 304634
rect 51562 304398 51646 304634
rect 51882 304398 87326 304634
rect 87562 304398 87646 304634
rect 87882 304398 123326 304634
rect 123562 304398 123646 304634
rect 123882 304398 159326 304634
rect 159562 304398 159646 304634
rect 159882 304398 195326 304634
rect 195562 304398 195646 304634
rect 195882 304398 231326 304634
rect 231562 304398 231646 304634
rect 231882 304398 267326 304634
rect 267562 304398 267646 304634
rect 267882 304398 303326 304634
rect 303562 304398 303646 304634
rect 303882 304398 339326 304634
rect 339562 304398 339646 304634
rect 339882 304398 375326 304634
rect 375562 304398 375646 304634
rect 375882 304398 411326 304634
rect 411562 304398 411646 304634
rect 411882 304398 447326 304634
rect 447562 304398 447646 304634
rect 447882 304398 483326 304634
rect 483562 304398 483646 304634
rect 483882 304398 519326 304634
rect 519562 304398 519646 304634
rect 519882 304398 555326 304634
rect 555562 304398 555646 304634
rect 555882 304398 588222 304634
rect 588458 304398 588542 304634
rect 588778 304398 592650 304634
rect -8726 304366 592650 304398
rect -8726 300454 592650 300486
rect -8726 300218 -3894 300454
rect -3658 300218 -3574 300454
rect -3338 300218 10826 300454
rect 11062 300218 11146 300454
rect 11382 300218 46826 300454
rect 47062 300218 47146 300454
rect 47382 300218 82826 300454
rect 83062 300218 83146 300454
rect 83382 300218 118826 300454
rect 119062 300218 119146 300454
rect 119382 300218 154826 300454
rect 155062 300218 155146 300454
rect 155382 300218 190826 300454
rect 191062 300218 191146 300454
rect 191382 300218 226826 300454
rect 227062 300218 227146 300454
rect 227382 300218 262826 300454
rect 263062 300218 263146 300454
rect 263382 300218 298826 300454
rect 299062 300218 299146 300454
rect 299382 300218 334826 300454
rect 335062 300218 335146 300454
rect 335382 300218 370826 300454
rect 371062 300218 371146 300454
rect 371382 300218 406826 300454
rect 407062 300218 407146 300454
rect 407382 300218 442826 300454
rect 443062 300218 443146 300454
rect 443382 300218 478826 300454
rect 479062 300218 479146 300454
rect 479382 300218 514826 300454
rect 515062 300218 515146 300454
rect 515382 300218 550826 300454
rect 551062 300218 551146 300454
rect 551382 300218 587262 300454
rect 587498 300218 587582 300454
rect 587818 300218 592650 300454
rect -8726 300134 592650 300218
rect -8726 299898 -3894 300134
rect -3658 299898 -3574 300134
rect -3338 299898 10826 300134
rect 11062 299898 11146 300134
rect 11382 299898 46826 300134
rect 47062 299898 47146 300134
rect 47382 299898 82826 300134
rect 83062 299898 83146 300134
rect 83382 299898 118826 300134
rect 119062 299898 119146 300134
rect 119382 299898 154826 300134
rect 155062 299898 155146 300134
rect 155382 299898 190826 300134
rect 191062 299898 191146 300134
rect 191382 299898 226826 300134
rect 227062 299898 227146 300134
rect 227382 299898 262826 300134
rect 263062 299898 263146 300134
rect 263382 299898 298826 300134
rect 299062 299898 299146 300134
rect 299382 299898 334826 300134
rect 335062 299898 335146 300134
rect 335382 299898 370826 300134
rect 371062 299898 371146 300134
rect 371382 299898 406826 300134
rect 407062 299898 407146 300134
rect 407382 299898 442826 300134
rect 443062 299898 443146 300134
rect 443382 299898 478826 300134
rect 479062 299898 479146 300134
rect 479382 299898 514826 300134
rect 515062 299898 515146 300134
rect 515382 299898 550826 300134
rect 551062 299898 551146 300134
rect 551382 299898 587262 300134
rect 587498 299898 587582 300134
rect 587818 299898 592650 300134
rect -8726 299866 592650 299898
rect -8726 295954 592650 295986
rect -8726 295718 -2934 295954
rect -2698 295718 -2614 295954
rect -2378 295718 6326 295954
rect 6562 295718 6646 295954
rect 6882 295718 42326 295954
rect 42562 295718 42646 295954
rect 42882 295718 78326 295954
rect 78562 295718 78646 295954
rect 78882 295718 114326 295954
rect 114562 295718 114646 295954
rect 114882 295718 150326 295954
rect 150562 295718 150646 295954
rect 150882 295718 186326 295954
rect 186562 295718 186646 295954
rect 186882 295718 222326 295954
rect 222562 295718 222646 295954
rect 222882 295718 258326 295954
rect 258562 295718 258646 295954
rect 258882 295718 294326 295954
rect 294562 295718 294646 295954
rect 294882 295718 330326 295954
rect 330562 295718 330646 295954
rect 330882 295718 366326 295954
rect 366562 295718 366646 295954
rect 366882 295718 402326 295954
rect 402562 295718 402646 295954
rect 402882 295718 438326 295954
rect 438562 295718 438646 295954
rect 438882 295718 474326 295954
rect 474562 295718 474646 295954
rect 474882 295718 510326 295954
rect 510562 295718 510646 295954
rect 510882 295718 546326 295954
rect 546562 295718 546646 295954
rect 546882 295718 582326 295954
rect 582562 295718 582646 295954
rect 582882 295718 586302 295954
rect 586538 295718 586622 295954
rect 586858 295718 592650 295954
rect -8726 295634 592650 295718
rect -8726 295398 -2934 295634
rect -2698 295398 -2614 295634
rect -2378 295398 6326 295634
rect 6562 295398 6646 295634
rect 6882 295398 42326 295634
rect 42562 295398 42646 295634
rect 42882 295398 78326 295634
rect 78562 295398 78646 295634
rect 78882 295398 114326 295634
rect 114562 295398 114646 295634
rect 114882 295398 150326 295634
rect 150562 295398 150646 295634
rect 150882 295398 186326 295634
rect 186562 295398 186646 295634
rect 186882 295398 222326 295634
rect 222562 295398 222646 295634
rect 222882 295398 258326 295634
rect 258562 295398 258646 295634
rect 258882 295398 294326 295634
rect 294562 295398 294646 295634
rect 294882 295398 330326 295634
rect 330562 295398 330646 295634
rect 330882 295398 366326 295634
rect 366562 295398 366646 295634
rect 366882 295398 402326 295634
rect 402562 295398 402646 295634
rect 402882 295398 438326 295634
rect 438562 295398 438646 295634
rect 438882 295398 474326 295634
rect 474562 295398 474646 295634
rect 474882 295398 510326 295634
rect 510562 295398 510646 295634
rect 510882 295398 546326 295634
rect 546562 295398 546646 295634
rect 546882 295398 582326 295634
rect 582562 295398 582646 295634
rect 582882 295398 586302 295634
rect 586538 295398 586622 295634
rect 586858 295398 592650 295634
rect -8726 295366 592650 295398
rect -8726 291454 592650 291486
rect -8726 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 73826 291454
rect 74062 291218 74146 291454
rect 74382 291218 109826 291454
rect 110062 291218 110146 291454
rect 110382 291218 145826 291454
rect 146062 291218 146146 291454
rect 146382 291218 181826 291454
rect 182062 291218 182146 291454
rect 182382 291218 217826 291454
rect 218062 291218 218146 291454
rect 218382 291218 253826 291454
rect 254062 291218 254146 291454
rect 254382 291218 289826 291454
rect 290062 291218 290146 291454
rect 290382 291218 325826 291454
rect 326062 291218 326146 291454
rect 326382 291218 361826 291454
rect 362062 291218 362146 291454
rect 362382 291218 397826 291454
rect 398062 291218 398146 291454
rect 398382 291218 433826 291454
rect 434062 291218 434146 291454
rect 434382 291218 469826 291454
rect 470062 291218 470146 291454
rect 470382 291218 505826 291454
rect 506062 291218 506146 291454
rect 506382 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 592650 291454
rect -8726 291134 592650 291218
rect -8726 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 73826 291134
rect 74062 290898 74146 291134
rect 74382 290898 109826 291134
rect 110062 290898 110146 291134
rect 110382 290898 145826 291134
rect 146062 290898 146146 291134
rect 146382 290898 181826 291134
rect 182062 290898 182146 291134
rect 182382 290898 217826 291134
rect 218062 290898 218146 291134
rect 218382 290898 253826 291134
rect 254062 290898 254146 291134
rect 254382 290898 289826 291134
rect 290062 290898 290146 291134
rect 290382 290898 325826 291134
rect 326062 290898 326146 291134
rect 326382 290898 361826 291134
rect 362062 290898 362146 291134
rect 362382 290898 397826 291134
rect 398062 290898 398146 291134
rect 398382 290898 433826 291134
rect 434062 290898 434146 291134
rect 434382 290898 469826 291134
rect 470062 290898 470146 291134
rect 470382 290898 505826 291134
rect 506062 290898 506146 291134
rect 506382 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 592650 291134
rect -8726 290866 592650 290898
rect -8726 286954 592650 286986
rect -8726 286718 -8694 286954
rect -8458 286718 -8374 286954
rect -8138 286718 33326 286954
rect 33562 286718 33646 286954
rect 33882 286718 69326 286954
rect 69562 286718 69646 286954
rect 69882 286718 105326 286954
rect 105562 286718 105646 286954
rect 105882 286718 141326 286954
rect 141562 286718 141646 286954
rect 141882 286718 177326 286954
rect 177562 286718 177646 286954
rect 177882 286718 213326 286954
rect 213562 286718 213646 286954
rect 213882 286718 249326 286954
rect 249562 286718 249646 286954
rect 249882 286718 285326 286954
rect 285562 286718 285646 286954
rect 285882 286718 321326 286954
rect 321562 286718 321646 286954
rect 321882 286718 357326 286954
rect 357562 286718 357646 286954
rect 357882 286718 393326 286954
rect 393562 286718 393646 286954
rect 393882 286718 429326 286954
rect 429562 286718 429646 286954
rect 429882 286718 465326 286954
rect 465562 286718 465646 286954
rect 465882 286718 501326 286954
rect 501562 286718 501646 286954
rect 501882 286718 537326 286954
rect 537562 286718 537646 286954
rect 537882 286718 573326 286954
rect 573562 286718 573646 286954
rect 573882 286718 592062 286954
rect 592298 286718 592382 286954
rect 592618 286718 592650 286954
rect -8726 286634 592650 286718
rect -8726 286398 -8694 286634
rect -8458 286398 -8374 286634
rect -8138 286398 33326 286634
rect 33562 286398 33646 286634
rect 33882 286398 69326 286634
rect 69562 286398 69646 286634
rect 69882 286398 105326 286634
rect 105562 286398 105646 286634
rect 105882 286398 141326 286634
rect 141562 286398 141646 286634
rect 141882 286398 177326 286634
rect 177562 286398 177646 286634
rect 177882 286398 213326 286634
rect 213562 286398 213646 286634
rect 213882 286398 249326 286634
rect 249562 286398 249646 286634
rect 249882 286398 285326 286634
rect 285562 286398 285646 286634
rect 285882 286398 321326 286634
rect 321562 286398 321646 286634
rect 321882 286398 357326 286634
rect 357562 286398 357646 286634
rect 357882 286398 393326 286634
rect 393562 286398 393646 286634
rect 393882 286398 429326 286634
rect 429562 286398 429646 286634
rect 429882 286398 465326 286634
rect 465562 286398 465646 286634
rect 465882 286398 501326 286634
rect 501562 286398 501646 286634
rect 501882 286398 537326 286634
rect 537562 286398 537646 286634
rect 537882 286398 573326 286634
rect 573562 286398 573646 286634
rect 573882 286398 592062 286634
rect 592298 286398 592382 286634
rect 592618 286398 592650 286634
rect -8726 286366 592650 286398
rect -8726 282454 592650 282486
rect -8726 282218 -7734 282454
rect -7498 282218 -7414 282454
rect -7178 282218 28826 282454
rect 29062 282218 29146 282454
rect 29382 282218 64826 282454
rect 65062 282218 65146 282454
rect 65382 282218 100826 282454
rect 101062 282218 101146 282454
rect 101382 282218 136826 282454
rect 137062 282218 137146 282454
rect 137382 282218 172826 282454
rect 173062 282218 173146 282454
rect 173382 282218 208826 282454
rect 209062 282218 209146 282454
rect 209382 282218 244826 282454
rect 245062 282218 245146 282454
rect 245382 282218 280826 282454
rect 281062 282218 281146 282454
rect 281382 282218 316826 282454
rect 317062 282218 317146 282454
rect 317382 282218 352826 282454
rect 353062 282218 353146 282454
rect 353382 282218 388826 282454
rect 389062 282218 389146 282454
rect 389382 282218 424826 282454
rect 425062 282218 425146 282454
rect 425382 282218 460826 282454
rect 461062 282218 461146 282454
rect 461382 282218 496826 282454
rect 497062 282218 497146 282454
rect 497382 282218 532826 282454
rect 533062 282218 533146 282454
rect 533382 282218 568826 282454
rect 569062 282218 569146 282454
rect 569382 282218 591102 282454
rect 591338 282218 591422 282454
rect 591658 282218 592650 282454
rect -8726 282134 592650 282218
rect -8726 281898 -7734 282134
rect -7498 281898 -7414 282134
rect -7178 281898 28826 282134
rect 29062 281898 29146 282134
rect 29382 281898 64826 282134
rect 65062 281898 65146 282134
rect 65382 281898 100826 282134
rect 101062 281898 101146 282134
rect 101382 281898 136826 282134
rect 137062 281898 137146 282134
rect 137382 281898 172826 282134
rect 173062 281898 173146 282134
rect 173382 281898 208826 282134
rect 209062 281898 209146 282134
rect 209382 281898 244826 282134
rect 245062 281898 245146 282134
rect 245382 281898 280826 282134
rect 281062 281898 281146 282134
rect 281382 281898 316826 282134
rect 317062 281898 317146 282134
rect 317382 281898 352826 282134
rect 353062 281898 353146 282134
rect 353382 281898 388826 282134
rect 389062 281898 389146 282134
rect 389382 281898 424826 282134
rect 425062 281898 425146 282134
rect 425382 281898 460826 282134
rect 461062 281898 461146 282134
rect 461382 281898 496826 282134
rect 497062 281898 497146 282134
rect 497382 281898 532826 282134
rect 533062 281898 533146 282134
rect 533382 281898 568826 282134
rect 569062 281898 569146 282134
rect 569382 281898 591102 282134
rect 591338 281898 591422 282134
rect 591658 281898 592650 282134
rect -8726 281866 592650 281898
rect -8726 277954 592650 277986
rect -8726 277718 -6774 277954
rect -6538 277718 -6454 277954
rect -6218 277718 24326 277954
rect 24562 277718 24646 277954
rect 24882 277718 60326 277954
rect 60562 277718 60646 277954
rect 60882 277718 96326 277954
rect 96562 277718 96646 277954
rect 96882 277718 132326 277954
rect 132562 277718 132646 277954
rect 132882 277718 168326 277954
rect 168562 277718 168646 277954
rect 168882 277718 204326 277954
rect 204562 277718 204646 277954
rect 204882 277718 240326 277954
rect 240562 277718 240646 277954
rect 240882 277718 276326 277954
rect 276562 277718 276646 277954
rect 276882 277718 312326 277954
rect 312562 277718 312646 277954
rect 312882 277718 348326 277954
rect 348562 277718 348646 277954
rect 348882 277718 384326 277954
rect 384562 277718 384646 277954
rect 384882 277718 420326 277954
rect 420562 277718 420646 277954
rect 420882 277718 456326 277954
rect 456562 277718 456646 277954
rect 456882 277718 492326 277954
rect 492562 277718 492646 277954
rect 492882 277718 528326 277954
rect 528562 277718 528646 277954
rect 528882 277718 564326 277954
rect 564562 277718 564646 277954
rect 564882 277718 590142 277954
rect 590378 277718 590462 277954
rect 590698 277718 592650 277954
rect -8726 277634 592650 277718
rect -8726 277398 -6774 277634
rect -6538 277398 -6454 277634
rect -6218 277398 24326 277634
rect 24562 277398 24646 277634
rect 24882 277398 60326 277634
rect 60562 277398 60646 277634
rect 60882 277398 96326 277634
rect 96562 277398 96646 277634
rect 96882 277398 132326 277634
rect 132562 277398 132646 277634
rect 132882 277398 168326 277634
rect 168562 277398 168646 277634
rect 168882 277398 204326 277634
rect 204562 277398 204646 277634
rect 204882 277398 240326 277634
rect 240562 277398 240646 277634
rect 240882 277398 276326 277634
rect 276562 277398 276646 277634
rect 276882 277398 312326 277634
rect 312562 277398 312646 277634
rect 312882 277398 348326 277634
rect 348562 277398 348646 277634
rect 348882 277398 384326 277634
rect 384562 277398 384646 277634
rect 384882 277398 420326 277634
rect 420562 277398 420646 277634
rect 420882 277398 456326 277634
rect 456562 277398 456646 277634
rect 456882 277398 492326 277634
rect 492562 277398 492646 277634
rect 492882 277398 528326 277634
rect 528562 277398 528646 277634
rect 528882 277398 564326 277634
rect 564562 277398 564646 277634
rect 564882 277398 590142 277634
rect 590378 277398 590462 277634
rect 590698 277398 592650 277634
rect -8726 277366 592650 277398
rect -8726 273454 592650 273486
rect -8726 273218 -5814 273454
rect -5578 273218 -5494 273454
rect -5258 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 55826 273454
rect 56062 273218 56146 273454
rect 56382 273218 91826 273454
rect 92062 273218 92146 273454
rect 92382 273218 127826 273454
rect 128062 273218 128146 273454
rect 128382 273218 163826 273454
rect 164062 273218 164146 273454
rect 164382 273218 199826 273454
rect 200062 273218 200146 273454
rect 200382 273218 235826 273454
rect 236062 273218 236146 273454
rect 236382 273218 271826 273454
rect 272062 273218 272146 273454
rect 272382 273218 307826 273454
rect 308062 273218 308146 273454
rect 308382 273218 343826 273454
rect 344062 273218 344146 273454
rect 344382 273218 379826 273454
rect 380062 273218 380146 273454
rect 380382 273218 415826 273454
rect 416062 273218 416146 273454
rect 416382 273218 451826 273454
rect 452062 273218 452146 273454
rect 452382 273218 487826 273454
rect 488062 273218 488146 273454
rect 488382 273218 523826 273454
rect 524062 273218 524146 273454
rect 524382 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 589182 273454
rect 589418 273218 589502 273454
rect 589738 273218 592650 273454
rect -8726 273134 592650 273218
rect -8726 272898 -5814 273134
rect -5578 272898 -5494 273134
rect -5258 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 55826 273134
rect 56062 272898 56146 273134
rect 56382 272898 91826 273134
rect 92062 272898 92146 273134
rect 92382 272898 127826 273134
rect 128062 272898 128146 273134
rect 128382 272898 163826 273134
rect 164062 272898 164146 273134
rect 164382 272898 199826 273134
rect 200062 272898 200146 273134
rect 200382 272898 235826 273134
rect 236062 272898 236146 273134
rect 236382 272898 271826 273134
rect 272062 272898 272146 273134
rect 272382 272898 307826 273134
rect 308062 272898 308146 273134
rect 308382 272898 343826 273134
rect 344062 272898 344146 273134
rect 344382 272898 379826 273134
rect 380062 272898 380146 273134
rect 380382 272898 415826 273134
rect 416062 272898 416146 273134
rect 416382 272898 451826 273134
rect 452062 272898 452146 273134
rect 452382 272898 487826 273134
rect 488062 272898 488146 273134
rect 488382 272898 523826 273134
rect 524062 272898 524146 273134
rect 524382 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 589182 273134
rect 589418 272898 589502 273134
rect 589738 272898 592650 273134
rect -8726 272866 592650 272898
rect -8726 268954 592650 268986
rect -8726 268718 -4854 268954
rect -4618 268718 -4534 268954
rect -4298 268718 15326 268954
rect 15562 268718 15646 268954
rect 15882 268718 51326 268954
rect 51562 268718 51646 268954
rect 51882 268718 87326 268954
rect 87562 268718 87646 268954
rect 87882 268718 123326 268954
rect 123562 268718 123646 268954
rect 123882 268718 159326 268954
rect 159562 268718 159646 268954
rect 159882 268718 195326 268954
rect 195562 268718 195646 268954
rect 195882 268718 231326 268954
rect 231562 268718 231646 268954
rect 231882 268718 267326 268954
rect 267562 268718 267646 268954
rect 267882 268718 303326 268954
rect 303562 268718 303646 268954
rect 303882 268718 339326 268954
rect 339562 268718 339646 268954
rect 339882 268718 375326 268954
rect 375562 268718 375646 268954
rect 375882 268718 411326 268954
rect 411562 268718 411646 268954
rect 411882 268718 447326 268954
rect 447562 268718 447646 268954
rect 447882 268718 483326 268954
rect 483562 268718 483646 268954
rect 483882 268718 519326 268954
rect 519562 268718 519646 268954
rect 519882 268718 555326 268954
rect 555562 268718 555646 268954
rect 555882 268718 588222 268954
rect 588458 268718 588542 268954
rect 588778 268718 592650 268954
rect -8726 268634 592650 268718
rect -8726 268398 -4854 268634
rect -4618 268398 -4534 268634
rect -4298 268398 15326 268634
rect 15562 268398 15646 268634
rect 15882 268398 51326 268634
rect 51562 268398 51646 268634
rect 51882 268398 87326 268634
rect 87562 268398 87646 268634
rect 87882 268398 123326 268634
rect 123562 268398 123646 268634
rect 123882 268398 159326 268634
rect 159562 268398 159646 268634
rect 159882 268398 195326 268634
rect 195562 268398 195646 268634
rect 195882 268398 231326 268634
rect 231562 268398 231646 268634
rect 231882 268398 267326 268634
rect 267562 268398 267646 268634
rect 267882 268398 303326 268634
rect 303562 268398 303646 268634
rect 303882 268398 339326 268634
rect 339562 268398 339646 268634
rect 339882 268398 375326 268634
rect 375562 268398 375646 268634
rect 375882 268398 411326 268634
rect 411562 268398 411646 268634
rect 411882 268398 447326 268634
rect 447562 268398 447646 268634
rect 447882 268398 483326 268634
rect 483562 268398 483646 268634
rect 483882 268398 519326 268634
rect 519562 268398 519646 268634
rect 519882 268398 555326 268634
rect 555562 268398 555646 268634
rect 555882 268398 588222 268634
rect 588458 268398 588542 268634
rect 588778 268398 592650 268634
rect -8726 268366 592650 268398
rect -8726 264454 592650 264486
rect -8726 264218 -3894 264454
rect -3658 264218 -3574 264454
rect -3338 264218 10826 264454
rect 11062 264218 11146 264454
rect 11382 264218 46826 264454
rect 47062 264218 47146 264454
rect 47382 264218 82826 264454
rect 83062 264218 83146 264454
rect 83382 264218 118826 264454
rect 119062 264218 119146 264454
rect 119382 264218 154826 264454
rect 155062 264218 155146 264454
rect 155382 264218 190826 264454
rect 191062 264218 191146 264454
rect 191382 264218 226826 264454
rect 227062 264218 227146 264454
rect 227382 264218 262826 264454
rect 263062 264218 263146 264454
rect 263382 264218 298826 264454
rect 299062 264218 299146 264454
rect 299382 264218 334826 264454
rect 335062 264218 335146 264454
rect 335382 264218 370826 264454
rect 371062 264218 371146 264454
rect 371382 264218 406826 264454
rect 407062 264218 407146 264454
rect 407382 264218 442826 264454
rect 443062 264218 443146 264454
rect 443382 264218 478826 264454
rect 479062 264218 479146 264454
rect 479382 264218 514826 264454
rect 515062 264218 515146 264454
rect 515382 264218 550826 264454
rect 551062 264218 551146 264454
rect 551382 264218 587262 264454
rect 587498 264218 587582 264454
rect 587818 264218 592650 264454
rect -8726 264134 592650 264218
rect -8726 263898 -3894 264134
rect -3658 263898 -3574 264134
rect -3338 263898 10826 264134
rect 11062 263898 11146 264134
rect 11382 263898 46826 264134
rect 47062 263898 47146 264134
rect 47382 263898 82826 264134
rect 83062 263898 83146 264134
rect 83382 263898 118826 264134
rect 119062 263898 119146 264134
rect 119382 263898 154826 264134
rect 155062 263898 155146 264134
rect 155382 263898 190826 264134
rect 191062 263898 191146 264134
rect 191382 263898 226826 264134
rect 227062 263898 227146 264134
rect 227382 263898 262826 264134
rect 263062 263898 263146 264134
rect 263382 263898 298826 264134
rect 299062 263898 299146 264134
rect 299382 263898 334826 264134
rect 335062 263898 335146 264134
rect 335382 263898 370826 264134
rect 371062 263898 371146 264134
rect 371382 263898 406826 264134
rect 407062 263898 407146 264134
rect 407382 263898 442826 264134
rect 443062 263898 443146 264134
rect 443382 263898 478826 264134
rect 479062 263898 479146 264134
rect 479382 263898 514826 264134
rect 515062 263898 515146 264134
rect 515382 263898 550826 264134
rect 551062 263898 551146 264134
rect 551382 263898 587262 264134
rect 587498 263898 587582 264134
rect 587818 263898 592650 264134
rect -8726 263866 592650 263898
rect -8726 259954 592650 259986
rect -8726 259718 -2934 259954
rect -2698 259718 -2614 259954
rect -2378 259718 6326 259954
rect 6562 259718 6646 259954
rect 6882 259718 42326 259954
rect 42562 259718 42646 259954
rect 42882 259718 78326 259954
rect 78562 259718 78646 259954
rect 78882 259718 114326 259954
rect 114562 259718 114646 259954
rect 114882 259718 222326 259954
rect 222562 259718 222646 259954
rect 222882 259718 258326 259954
rect 258562 259718 258646 259954
rect 258882 259718 294326 259954
rect 294562 259718 294646 259954
rect 294882 259718 330326 259954
rect 330562 259718 330646 259954
rect 330882 259718 366326 259954
rect 366562 259718 366646 259954
rect 366882 259718 402326 259954
rect 402562 259718 402646 259954
rect 402882 259718 438326 259954
rect 438562 259718 438646 259954
rect 438882 259718 474326 259954
rect 474562 259718 474646 259954
rect 474882 259718 510326 259954
rect 510562 259718 510646 259954
rect 510882 259718 546326 259954
rect 546562 259718 546646 259954
rect 546882 259718 582326 259954
rect 582562 259718 582646 259954
rect 582882 259718 586302 259954
rect 586538 259718 586622 259954
rect 586858 259718 592650 259954
rect -8726 259634 592650 259718
rect -8726 259398 -2934 259634
rect -2698 259398 -2614 259634
rect -2378 259398 6326 259634
rect 6562 259398 6646 259634
rect 6882 259398 42326 259634
rect 42562 259398 42646 259634
rect 42882 259398 78326 259634
rect 78562 259398 78646 259634
rect 78882 259398 114326 259634
rect 114562 259398 114646 259634
rect 114882 259398 222326 259634
rect 222562 259398 222646 259634
rect 222882 259398 258326 259634
rect 258562 259398 258646 259634
rect 258882 259398 294326 259634
rect 294562 259398 294646 259634
rect 294882 259398 330326 259634
rect 330562 259398 330646 259634
rect 330882 259398 366326 259634
rect 366562 259398 366646 259634
rect 366882 259398 402326 259634
rect 402562 259398 402646 259634
rect 402882 259398 438326 259634
rect 438562 259398 438646 259634
rect 438882 259398 474326 259634
rect 474562 259398 474646 259634
rect 474882 259398 510326 259634
rect 510562 259398 510646 259634
rect 510882 259398 546326 259634
rect 546562 259398 546646 259634
rect 546882 259398 582326 259634
rect 582562 259398 582646 259634
rect 582882 259398 586302 259634
rect 586538 259398 586622 259634
rect 586858 259398 592650 259634
rect -8726 259366 592650 259398
rect -8726 255454 592650 255486
rect -8726 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 73826 255454
rect 74062 255218 74146 255454
rect 74382 255218 109826 255454
rect 110062 255218 110146 255454
rect 110382 255218 124250 255454
rect 124486 255218 154970 255454
rect 155206 255218 185690 255454
rect 185926 255218 217826 255454
rect 218062 255218 218146 255454
rect 218382 255218 253826 255454
rect 254062 255218 254146 255454
rect 254382 255218 289826 255454
rect 290062 255218 290146 255454
rect 290382 255218 325826 255454
rect 326062 255218 326146 255454
rect 326382 255218 361826 255454
rect 362062 255218 362146 255454
rect 362382 255218 397826 255454
rect 398062 255218 398146 255454
rect 398382 255218 433826 255454
rect 434062 255218 434146 255454
rect 434382 255218 469826 255454
rect 470062 255218 470146 255454
rect 470382 255218 505826 255454
rect 506062 255218 506146 255454
rect 506382 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 592650 255454
rect -8726 255134 592650 255218
rect -8726 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 73826 255134
rect 74062 254898 74146 255134
rect 74382 254898 109826 255134
rect 110062 254898 110146 255134
rect 110382 254898 124250 255134
rect 124486 254898 154970 255134
rect 155206 254898 185690 255134
rect 185926 254898 217826 255134
rect 218062 254898 218146 255134
rect 218382 254898 253826 255134
rect 254062 254898 254146 255134
rect 254382 254898 289826 255134
rect 290062 254898 290146 255134
rect 290382 254898 325826 255134
rect 326062 254898 326146 255134
rect 326382 254898 361826 255134
rect 362062 254898 362146 255134
rect 362382 254898 397826 255134
rect 398062 254898 398146 255134
rect 398382 254898 433826 255134
rect 434062 254898 434146 255134
rect 434382 254898 469826 255134
rect 470062 254898 470146 255134
rect 470382 254898 505826 255134
rect 506062 254898 506146 255134
rect 506382 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 592650 255134
rect -8726 254866 592650 254898
rect -8726 250954 592650 250986
rect -8726 250718 -8694 250954
rect -8458 250718 -8374 250954
rect -8138 250718 33326 250954
rect 33562 250718 33646 250954
rect 33882 250718 69326 250954
rect 69562 250718 69646 250954
rect 69882 250718 105326 250954
rect 105562 250718 105646 250954
rect 105882 250718 213326 250954
rect 213562 250718 213646 250954
rect 213882 250718 249326 250954
rect 249562 250718 249646 250954
rect 249882 250718 285326 250954
rect 285562 250718 285646 250954
rect 285882 250718 321326 250954
rect 321562 250718 321646 250954
rect 321882 250718 357326 250954
rect 357562 250718 357646 250954
rect 357882 250718 393326 250954
rect 393562 250718 393646 250954
rect 393882 250718 429326 250954
rect 429562 250718 429646 250954
rect 429882 250718 465326 250954
rect 465562 250718 465646 250954
rect 465882 250718 501326 250954
rect 501562 250718 501646 250954
rect 501882 250718 537326 250954
rect 537562 250718 537646 250954
rect 537882 250718 573326 250954
rect 573562 250718 573646 250954
rect 573882 250718 592062 250954
rect 592298 250718 592382 250954
rect 592618 250718 592650 250954
rect -8726 250634 592650 250718
rect -8726 250398 -8694 250634
rect -8458 250398 -8374 250634
rect -8138 250398 33326 250634
rect 33562 250398 33646 250634
rect 33882 250398 69326 250634
rect 69562 250398 69646 250634
rect 69882 250398 105326 250634
rect 105562 250398 105646 250634
rect 105882 250398 213326 250634
rect 213562 250398 213646 250634
rect 213882 250398 249326 250634
rect 249562 250398 249646 250634
rect 249882 250398 285326 250634
rect 285562 250398 285646 250634
rect 285882 250398 321326 250634
rect 321562 250398 321646 250634
rect 321882 250398 357326 250634
rect 357562 250398 357646 250634
rect 357882 250398 393326 250634
rect 393562 250398 393646 250634
rect 393882 250398 429326 250634
rect 429562 250398 429646 250634
rect 429882 250398 465326 250634
rect 465562 250398 465646 250634
rect 465882 250398 501326 250634
rect 501562 250398 501646 250634
rect 501882 250398 537326 250634
rect 537562 250398 537646 250634
rect 537882 250398 573326 250634
rect 573562 250398 573646 250634
rect 573882 250398 592062 250634
rect 592298 250398 592382 250634
rect 592618 250398 592650 250634
rect -8726 250366 592650 250398
rect -8726 246454 592650 246486
rect -8726 246218 -7734 246454
rect -7498 246218 -7414 246454
rect -7178 246218 28826 246454
rect 29062 246218 29146 246454
rect 29382 246218 64826 246454
rect 65062 246218 65146 246454
rect 65382 246218 100826 246454
rect 101062 246218 101146 246454
rect 101382 246218 208826 246454
rect 209062 246218 209146 246454
rect 209382 246218 244826 246454
rect 245062 246218 245146 246454
rect 245382 246218 280826 246454
rect 281062 246218 281146 246454
rect 281382 246218 316826 246454
rect 317062 246218 317146 246454
rect 317382 246218 352826 246454
rect 353062 246218 353146 246454
rect 353382 246218 388826 246454
rect 389062 246218 389146 246454
rect 389382 246218 424826 246454
rect 425062 246218 425146 246454
rect 425382 246218 460826 246454
rect 461062 246218 461146 246454
rect 461382 246218 496826 246454
rect 497062 246218 497146 246454
rect 497382 246218 532826 246454
rect 533062 246218 533146 246454
rect 533382 246218 568826 246454
rect 569062 246218 569146 246454
rect 569382 246218 591102 246454
rect 591338 246218 591422 246454
rect 591658 246218 592650 246454
rect -8726 246134 592650 246218
rect -8726 245898 -7734 246134
rect -7498 245898 -7414 246134
rect -7178 245898 28826 246134
rect 29062 245898 29146 246134
rect 29382 245898 64826 246134
rect 65062 245898 65146 246134
rect 65382 245898 100826 246134
rect 101062 245898 101146 246134
rect 101382 245898 208826 246134
rect 209062 245898 209146 246134
rect 209382 245898 244826 246134
rect 245062 245898 245146 246134
rect 245382 245898 280826 246134
rect 281062 245898 281146 246134
rect 281382 245898 316826 246134
rect 317062 245898 317146 246134
rect 317382 245898 352826 246134
rect 353062 245898 353146 246134
rect 353382 245898 388826 246134
rect 389062 245898 389146 246134
rect 389382 245898 424826 246134
rect 425062 245898 425146 246134
rect 425382 245898 460826 246134
rect 461062 245898 461146 246134
rect 461382 245898 496826 246134
rect 497062 245898 497146 246134
rect 497382 245898 532826 246134
rect 533062 245898 533146 246134
rect 533382 245898 568826 246134
rect 569062 245898 569146 246134
rect 569382 245898 591102 246134
rect 591338 245898 591422 246134
rect 591658 245898 592650 246134
rect -8726 245866 592650 245898
rect -8726 241954 592650 241986
rect -8726 241718 -6774 241954
rect -6538 241718 -6454 241954
rect -6218 241718 24326 241954
rect 24562 241718 24646 241954
rect 24882 241718 60326 241954
rect 60562 241718 60646 241954
rect 60882 241718 96326 241954
rect 96562 241718 96646 241954
rect 96882 241718 204326 241954
rect 204562 241718 204646 241954
rect 204882 241718 240326 241954
rect 240562 241718 240646 241954
rect 240882 241718 276326 241954
rect 276562 241718 276646 241954
rect 276882 241718 312326 241954
rect 312562 241718 312646 241954
rect 312882 241718 348326 241954
rect 348562 241718 348646 241954
rect 348882 241718 384326 241954
rect 384562 241718 384646 241954
rect 384882 241718 420326 241954
rect 420562 241718 420646 241954
rect 420882 241718 456326 241954
rect 456562 241718 456646 241954
rect 456882 241718 492326 241954
rect 492562 241718 492646 241954
rect 492882 241718 528326 241954
rect 528562 241718 528646 241954
rect 528882 241718 564326 241954
rect 564562 241718 564646 241954
rect 564882 241718 590142 241954
rect 590378 241718 590462 241954
rect 590698 241718 592650 241954
rect -8726 241634 592650 241718
rect -8726 241398 -6774 241634
rect -6538 241398 -6454 241634
rect -6218 241398 24326 241634
rect 24562 241398 24646 241634
rect 24882 241398 60326 241634
rect 60562 241398 60646 241634
rect 60882 241398 96326 241634
rect 96562 241398 96646 241634
rect 96882 241398 204326 241634
rect 204562 241398 204646 241634
rect 204882 241398 240326 241634
rect 240562 241398 240646 241634
rect 240882 241398 276326 241634
rect 276562 241398 276646 241634
rect 276882 241398 312326 241634
rect 312562 241398 312646 241634
rect 312882 241398 348326 241634
rect 348562 241398 348646 241634
rect 348882 241398 384326 241634
rect 384562 241398 384646 241634
rect 384882 241398 420326 241634
rect 420562 241398 420646 241634
rect 420882 241398 456326 241634
rect 456562 241398 456646 241634
rect 456882 241398 492326 241634
rect 492562 241398 492646 241634
rect 492882 241398 528326 241634
rect 528562 241398 528646 241634
rect 528882 241398 564326 241634
rect 564562 241398 564646 241634
rect 564882 241398 590142 241634
rect 590378 241398 590462 241634
rect 590698 241398 592650 241634
rect -8726 241366 592650 241398
rect -8726 237454 592650 237486
rect -8726 237218 -5814 237454
rect -5578 237218 -5494 237454
rect -5258 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 55826 237454
rect 56062 237218 56146 237454
rect 56382 237218 91826 237454
rect 92062 237218 92146 237454
rect 92382 237218 199826 237454
rect 200062 237218 200146 237454
rect 200382 237218 235826 237454
rect 236062 237218 236146 237454
rect 236382 237218 271826 237454
rect 272062 237218 272146 237454
rect 272382 237218 307826 237454
rect 308062 237218 308146 237454
rect 308382 237218 343826 237454
rect 344062 237218 344146 237454
rect 344382 237218 379826 237454
rect 380062 237218 380146 237454
rect 380382 237218 415826 237454
rect 416062 237218 416146 237454
rect 416382 237218 451826 237454
rect 452062 237218 452146 237454
rect 452382 237218 487826 237454
rect 488062 237218 488146 237454
rect 488382 237218 523826 237454
rect 524062 237218 524146 237454
rect 524382 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 589182 237454
rect 589418 237218 589502 237454
rect 589738 237218 592650 237454
rect -8726 237134 592650 237218
rect -8726 236898 -5814 237134
rect -5578 236898 -5494 237134
rect -5258 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 55826 237134
rect 56062 236898 56146 237134
rect 56382 236898 91826 237134
rect 92062 236898 92146 237134
rect 92382 236898 199826 237134
rect 200062 236898 200146 237134
rect 200382 236898 235826 237134
rect 236062 236898 236146 237134
rect 236382 236898 271826 237134
rect 272062 236898 272146 237134
rect 272382 236898 307826 237134
rect 308062 236898 308146 237134
rect 308382 236898 343826 237134
rect 344062 236898 344146 237134
rect 344382 236898 379826 237134
rect 380062 236898 380146 237134
rect 380382 236898 415826 237134
rect 416062 236898 416146 237134
rect 416382 236898 451826 237134
rect 452062 236898 452146 237134
rect 452382 236898 487826 237134
rect 488062 236898 488146 237134
rect 488382 236898 523826 237134
rect 524062 236898 524146 237134
rect 524382 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 589182 237134
rect 589418 236898 589502 237134
rect 589738 236898 592650 237134
rect -8726 236866 592650 236898
rect -8726 232954 592650 232986
rect -8726 232718 -4854 232954
rect -4618 232718 -4534 232954
rect -4298 232718 15326 232954
rect 15562 232718 15646 232954
rect 15882 232718 51326 232954
rect 51562 232718 51646 232954
rect 51882 232718 87326 232954
rect 87562 232718 87646 232954
rect 87882 232718 195326 232954
rect 195562 232718 195646 232954
rect 195882 232718 231326 232954
rect 231562 232718 231646 232954
rect 231882 232718 267326 232954
rect 267562 232718 267646 232954
rect 267882 232718 303326 232954
rect 303562 232718 303646 232954
rect 303882 232718 339326 232954
rect 339562 232718 339646 232954
rect 339882 232718 375326 232954
rect 375562 232718 375646 232954
rect 375882 232718 411326 232954
rect 411562 232718 411646 232954
rect 411882 232718 447326 232954
rect 447562 232718 447646 232954
rect 447882 232718 483326 232954
rect 483562 232718 483646 232954
rect 483882 232718 519326 232954
rect 519562 232718 519646 232954
rect 519882 232718 555326 232954
rect 555562 232718 555646 232954
rect 555882 232718 588222 232954
rect 588458 232718 588542 232954
rect 588778 232718 592650 232954
rect -8726 232634 592650 232718
rect -8726 232398 -4854 232634
rect -4618 232398 -4534 232634
rect -4298 232398 15326 232634
rect 15562 232398 15646 232634
rect 15882 232398 51326 232634
rect 51562 232398 51646 232634
rect 51882 232398 87326 232634
rect 87562 232398 87646 232634
rect 87882 232398 195326 232634
rect 195562 232398 195646 232634
rect 195882 232398 231326 232634
rect 231562 232398 231646 232634
rect 231882 232398 267326 232634
rect 267562 232398 267646 232634
rect 267882 232398 303326 232634
rect 303562 232398 303646 232634
rect 303882 232398 339326 232634
rect 339562 232398 339646 232634
rect 339882 232398 375326 232634
rect 375562 232398 375646 232634
rect 375882 232398 411326 232634
rect 411562 232398 411646 232634
rect 411882 232398 447326 232634
rect 447562 232398 447646 232634
rect 447882 232398 483326 232634
rect 483562 232398 483646 232634
rect 483882 232398 519326 232634
rect 519562 232398 519646 232634
rect 519882 232398 555326 232634
rect 555562 232398 555646 232634
rect 555882 232398 588222 232634
rect 588458 232398 588542 232634
rect 588778 232398 592650 232634
rect -8726 232366 592650 232398
rect -8726 228454 592650 228486
rect -8726 228218 -3894 228454
rect -3658 228218 -3574 228454
rect -3338 228218 10826 228454
rect 11062 228218 11146 228454
rect 11382 228218 46826 228454
rect 47062 228218 47146 228454
rect 47382 228218 82826 228454
rect 83062 228218 83146 228454
rect 83382 228218 226826 228454
rect 227062 228218 227146 228454
rect 227382 228218 262826 228454
rect 263062 228218 263146 228454
rect 263382 228218 298826 228454
rect 299062 228218 299146 228454
rect 299382 228218 334826 228454
rect 335062 228218 335146 228454
rect 335382 228218 370826 228454
rect 371062 228218 371146 228454
rect 371382 228218 406826 228454
rect 407062 228218 407146 228454
rect 407382 228218 442826 228454
rect 443062 228218 443146 228454
rect 443382 228218 478826 228454
rect 479062 228218 479146 228454
rect 479382 228218 514826 228454
rect 515062 228218 515146 228454
rect 515382 228218 550826 228454
rect 551062 228218 551146 228454
rect 551382 228218 587262 228454
rect 587498 228218 587582 228454
rect 587818 228218 592650 228454
rect -8726 228134 592650 228218
rect -8726 227898 -3894 228134
rect -3658 227898 -3574 228134
rect -3338 227898 10826 228134
rect 11062 227898 11146 228134
rect 11382 227898 46826 228134
rect 47062 227898 47146 228134
rect 47382 227898 82826 228134
rect 83062 227898 83146 228134
rect 83382 227898 226826 228134
rect 227062 227898 227146 228134
rect 227382 227898 262826 228134
rect 263062 227898 263146 228134
rect 263382 227898 298826 228134
rect 299062 227898 299146 228134
rect 299382 227898 334826 228134
rect 335062 227898 335146 228134
rect 335382 227898 370826 228134
rect 371062 227898 371146 228134
rect 371382 227898 406826 228134
rect 407062 227898 407146 228134
rect 407382 227898 442826 228134
rect 443062 227898 443146 228134
rect 443382 227898 478826 228134
rect 479062 227898 479146 228134
rect 479382 227898 514826 228134
rect 515062 227898 515146 228134
rect 515382 227898 550826 228134
rect 551062 227898 551146 228134
rect 551382 227898 587262 228134
rect 587498 227898 587582 228134
rect 587818 227898 592650 228134
rect -8726 227866 592650 227898
rect -8726 223954 592650 223986
rect -8726 223718 -2934 223954
rect -2698 223718 -2614 223954
rect -2378 223718 6326 223954
rect 6562 223718 6646 223954
rect 6882 223718 42326 223954
rect 42562 223718 42646 223954
rect 42882 223718 78326 223954
rect 78562 223718 78646 223954
rect 78882 223718 114326 223954
rect 114562 223718 114646 223954
rect 114882 223718 139610 223954
rect 139846 223718 170330 223954
rect 170566 223718 222326 223954
rect 222562 223718 222646 223954
rect 222882 223718 258326 223954
rect 258562 223718 258646 223954
rect 258882 223718 294326 223954
rect 294562 223718 294646 223954
rect 294882 223718 330326 223954
rect 330562 223718 330646 223954
rect 330882 223718 366326 223954
rect 366562 223718 366646 223954
rect 366882 223718 402326 223954
rect 402562 223718 402646 223954
rect 402882 223718 438326 223954
rect 438562 223718 438646 223954
rect 438882 223718 474326 223954
rect 474562 223718 474646 223954
rect 474882 223718 510326 223954
rect 510562 223718 510646 223954
rect 510882 223718 546326 223954
rect 546562 223718 546646 223954
rect 546882 223718 582326 223954
rect 582562 223718 582646 223954
rect 582882 223718 586302 223954
rect 586538 223718 586622 223954
rect 586858 223718 592650 223954
rect -8726 223634 592650 223718
rect -8726 223398 -2934 223634
rect -2698 223398 -2614 223634
rect -2378 223398 6326 223634
rect 6562 223398 6646 223634
rect 6882 223398 42326 223634
rect 42562 223398 42646 223634
rect 42882 223398 78326 223634
rect 78562 223398 78646 223634
rect 78882 223398 114326 223634
rect 114562 223398 114646 223634
rect 114882 223398 139610 223634
rect 139846 223398 170330 223634
rect 170566 223398 222326 223634
rect 222562 223398 222646 223634
rect 222882 223398 258326 223634
rect 258562 223398 258646 223634
rect 258882 223398 294326 223634
rect 294562 223398 294646 223634
rect 294882 223398 330326 223634
rect 330562 223398 330646 223634
rect 330882 223398 366326 223634
rect 366562 223398 366646 223634
rect 366882 223398 402326 223634
rect 402562 223398 402646 223634
rect 402882 223398 438326 223634
rect 438562 223398 438646 223634
rect 438882 223398 474326 223634
rect 474562 223398 474646 223634
rect 474882 223398 510326 223634
rect 510562 223398 510646 223634
rect 510882 223398 546326 223634
rect 546562 223398 546646 223634
rect 546882 223398 582326 223634
rect 582562 223398 582646 223634
rect 582882 223398 586302 223634
rect 586538 223398 586622 223634
rect 586858 223398 592650 223634
rect -8726 223366 592650 223398
rect -8726 219454 592650 219486
rect -8726 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 73826 219454
rect 74062 219218 74146 219454
rect 74382 219218 109826 219454
rect 110062 219218 110146 219454
rect 110382 219218 124250 219454
rect 124486 219218 154970 219454
rect 155206 219218 185690 219454
rect 185926 219218 217826 219454
rect 218062 219218 218146 219454
rect 218382 219218 253826 219454
rect 254062 219218 254146 219454
rect 254382 219218 289826 219454
rect 290062 219218 290146 219454
rect 290382 219218 325826 219454
rect 326062 219218 326146 219454
rect 326382 219218 361826 219454
rect 362062 219218 362146 219454
rect 362382 219218 397826 219454
rect 398062 219218 398146 219454
rect 398382 219218 433826 219454
rect 434062 219218 434146 219454
rect 434382 219218 469826 219454
rect 470062 219218 470146 219454
rect 470382 219218 505826 219454
rect 506062 219218 506146 219454
rect 506382 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 592650 219454
rect -8726 219134 592650 219218
rect -8726 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 73826 219134
rect 74062 218898 74146 219134
rect 74382 218898 109826 219134
rect 110062 218898 110146 219134
rect 110382 218898 124250 219134
rect 124486 218898 154970 219134
rect 155206 218898 185690 219134
rect 185926 218898 217826 219134
rect 218062 218898 218146 219134
rect 218382 218898 253826 219134
rect 254062 218898 254146 219134
rect 254382 218898 289826 219134
rect 290062 218898 290146 219134
rect 290382 218898 325826 219134
rect 326062 218898 326146 219134
rect 326382 218898 361826 219134
rect 362062 218898 362146 219134
rect 362382 218898 397826 219134
rect 398062 218898 398146 219134
rect 398382 218898 433826 219134
rect 434062 218898 434146 219134
rect 434382 218898 469826 219134
rect 470062 218898 470146 219134
rect 470382 218898 505826 219134
rect 506062 218898 506146 219134
rect 506382 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 592650 219134
rect -8726 218866 592650 218898
rect -8726 214954 592650 214986
rect -8726 214718 -8694 214954
rect -8458 214718 -8374 214954
rect -8138 214718 33326 214954
rect 33562 214718 33646 214954
rect 33882 214718 69326 214954
rect 69562 214718 69646 214954
rect 69882 214718 105326 214954
rect 105562 214718 105646 214954
rect 105882 214718 213326 214954
rect 213562 214718 213646 214954
rect 213882 214718 249326 214954
rect 249562 214718 249646 214954
rect 249882 214718 285326 214954
rect 285562 214718 285646 214954
rect 285882 214718 321326 214954
rect 321562 214718 321646 214954
rect 321882 214718 357326 214954
rect 357562 214718 357646 214954
rect 357882 214718 393326 214954
rect 393562 214718 393646 214954
rect 393882 214718 429326 214954
rect 429562 214718 429646 214954
rect 429882 214718 465326 214954
rect 465562 214718 465646 214954
rect 465882 214718 501326 214954
rect 501562 214718 501646 214954
rect 501882 214718 537326 214954
rect 537562 214718 537646 214954
rect 537882 214718 573326 214954
rect 573562 214718 573646 214954
rect 573882 214718 592062 214954
rect 592298 214718 592382 214954
rect 592618 214718 592650 214954
rect -8726 214634 592650 214718
rect -8726 214398 -8694 214634
rect -8458 214398 -8374 214634
rect -8138 214398 33326 214634
rect 33562 214398 33646 214634
rect 33882 214398 69326 214634
rect 69562 214398 69646 214634
rect 69882 214398 105326 214634
rect 105562 214398 105646 214634
rect 105882 214398 213326 214634
rect 213562 214398 213646 214634
rect 213882 214398 249326 214634
rect 249562 214398 249646 214634
rect 249882 214398 285326 214634
rect 285562 214398 285646 214634
rect 285882 214398 321326 214634
rect 321562 214398 321646 214634
rect 321882 214398 357326 214634
rect 357562 214398 357646 214634
rect 357882 214398 393326 214634
rect 393562 214398 393646 214634
rect 393882 214398 429326 214634
rect 429562 214398 429646 214634
rect 429882 214398 465326 214634
rect 465562 214398 465646 214634
rect 465882 214398 501326 214634
rect 501562 214398 501646 214634
rect 501882 214398 537326 214634
rect 537562 214398 537646 214634
rect 537882 214398 573326 214634
rect 573562 214398 573646 214634
rect 573882 214398 592062 214634
rect 592298 214398 592382 214634
rect 592618 214398 592650 214634
rect -8726 214366 592650 214398
rect -8726 210454 592650 210486
rect -8726 210218 -7734 210454
rect -7498 210218 -7414 210454
rect -7178 210218 28826 210454
rect 29062 210218 29146 210454
rect 29382 210218 64826 210454
rect 65062 210218 65146 210454
rect 65382 210218 100826 210454
rect 101062 210218 101146 210454
rect 101382 210218 208826 210454
rect 209062 210218 209146 210454
rect 209382 210218 244826 210454
rect 245062 210218 245146 210454
rect 245382 210218 280826 210454
rect 281062 210218 281146 210454
rect 281382 210218 316826 210454
rect 317062 210218 317146 210454
rect 317382 210218 352826 210454
rect 353062 210218 353146 210454
rect 353382 210218 388826 210454
rect 389062 210218 389146 210454
rect 389382 210218 424826 210454
rect 425062 210218 425146 210454
rect 425382 210218 460826 210454
rect 461062 210218 461146 210454
rect 461382 210218 496826 210454
rect 497062 210218 497146 210454
rect 497382 210218 532826 210454
rect 533062 210218 533146 210454
rect 533382 210218 568826 210454
rect 569062 210218 569146 210454
rect 569382 210218 591102 210454
rect 591338 210218 591422 210454
rect 591658 210218 592650 210454
rect -8726 210134 592650 210218
rect -8726 209898 -7734 210134
rect -7498 209898 -7414 210134
rect -7178 209898 28826 210134
rect 29062 209898 29146 210134
rect 29382 209898 64826 210134
rect 65062 209898 65146 210134
rect 65382 209898 100826 210134
rect 101062 209898 101146 210134
rect 101382 209898 208826 210134
rect 209062 209898 209146 210134
rect 209382 209898 244826 210134
rect 245062 209898 245146 210134
rect 245382 209898 280826 210134
rect 281062 209898 281146 210134
rect 281382 209898 316826 210134
rect 317062 209898 317146 210134
rect 317382 209898 352826 210134
rect 353062 209898 353146 210134
rect 353382 209898 388826 210134
rect 389062 209898 389146 210134
rect 389382 209898 424826 210134
rect 425062 209898 425146 210134
rect 425382 209898 460826 210134
rect 461062 209898 461146 210134
rect 461382 209898 496826 210134
rect 497062 209898 497146 210134
rect 497382 209898 532826 210134
rect 533062 209898 533146 210134
rect 533382 209898 568826 210134
rect 569062 209898 569146 210134
rect 569382 209898 591102 210134
rect 591338 209898 591422 210134
rect 591658 209898 592650 210134
rect -8726 209866 592650 209898
rect -8726 205954 592650 205986
rect -8726 205718 -6774 205954
rect -6538 205718 -6454 205954
rect -6218 205718 24326 205954
rect 24562 205718 24646 205954
rect 24882 205718 60326 205954
rect 60562 205718 60646 205954
rect 60882 205718 96326 205954
rect 96562 205718 96646 205954
rect 96882 205718 204326 205954
rect 204562 205718 204646 205954
rect 204882 205718 240326 205954
rect 240562 205718 240646 205954
rect 240882 205718 276326 205954
rect 276562 205718 276646 205954
rect 276882 205718 312326 205954
rect 312562 205718 312646 205954
rect 312882 205718 348326 205954
rect 348562 205718 348646 205954
rect 348882 205718 384326 205954
rect 384562 205718 384646 205954
rect 384882 205718 420326 205954
rect 420562 205718 420646 205954
rect 420882 205718 456326 205954
rect 456562 205718 456646 205954
rect 456882 205718 492326 205954
rect 492562 205718 492646 205954
rect 492882 205718 528326 205954
rect 528562 205718 528646 205954
rect 528882 205718 564326 205954
rect 564562 205718 564646 205954
rect 564882 205718 590142 205954
rect 590378 205718 590462 205954
rect 590698 205718 592650 205954
rect -8726 205634 592650 205718
rect -8726 205398 -6774 205634
rect -6538 205398 -6454 205634
rect -6218 205398 24326 205634
rect 24562 205398 24646 205634
rect 24882 205398 60326 205634
rect 60562 205398 60646 205634
rect 60882 205398 96326 205634
rect 96562 205398 96646 205634
rect 96882 205398 204326 205634
rect 204562 205398 204646 205634
rect 204882 205398 240326 205634
rect 240562 205398 240646 205634
rect 240882 205398 276326 205634
rect 276562 205398 276646 205634
rect 276882 205398 312326 205634
rect 312562 205398 312646 205634
rect 312882 205398 348326 205634
rect 348562 205398 348646 205634
rect 348882 205398 384326 205634
rect 384562 205398 384646 205634
rect 384882 205398 420326 205634
rect 420562 205398 420646 205634
rect 420882 205398 456326 205634
rect 456562 205398 456646 205634
rect 456882 205398 492326 205634
rect 492562 205398 492646 205634
rect 492882 205398 528326 205634
rect 528562 205398 528646 205634
rect 528882 205398 564326 205634
rect 564562 205398 564646 205634
rect 564882 205398 590142 205634
rect 590378 205398 590462 205634
rect 590698 205398 592650 205634
rect -8726 205366 592650 205398
rect -8726 201454 592650 201486
rect -8726 201218 -5814 201454
rect -5578 201218 -5494 201454
rect -5258 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 55826 201454
rect 56062 201218 56146 201454
rect 56382 201218 91826 201454
rect 92062 201218 92146 201454
rect 92382 201218 199826 201454
rect 200062 201218 200146 201454
rect 200382 201218 235826 201454
rect 236062 201218 236146 201454
rect 236382 201218 271826 201454
rect 272062 201218 272146 201454
rect 272382 201218 307826 201454
rect 308062 201218 308146 201454
rect 308382 201218 343826 201454
rect 344062 201218 344146 201454
rect 344382 201218 379826 201454
rect 380062 201218 380146 201454
rect 380382 201218 415826 201454
rect 416062 201218 416146 201454
rect 416382 201218 451826 201454
rect 452062 201218 452146 201454
rect 452382 201218 487826 201454
rect 488062 201218 488146 201454
rect 488382 201218 523826 201454
rect 524062 201218 524146 201454
rect 524382 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 589182 201454
rect 589418 201218 589502 201454
rect 589738 201218 592650 201454
rect -8726 201134 592650 201218
rect -8726 200898 -5814 201134
rect -5578 200898 -5494 201134
rect -5258 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 55826 201134
rect 56062 200898 56146 201134
rect 56382 200898 91826 201134
rect 92062 200898 92146 201134
rect 92382 200898 199826 201134
rect 200062 200898 200146 201134
rect 200382 200898 235826 201134
rect 236062 200898 236146 201134
rect 236382 200898 271826 201134
rect 272062 200898 272146 201134
rect 272382 200898 307826 201134
rect 308062 200898 308146 201134
rect 308382 200898 343826 201134
rect 344062 200898 344146 201134
rect 344382 200898 379826 201134
rect 380062 200898 380146 201134
rect 380382 200898 415826 201134
rect 416062 200898 416146 201134
rect 416382 200898 451826 201134
rect 452062 200898 452146 201134
rect 452382 200898 487826 201134
rect 488062 200898 488146 201134
rect 488382 200898 523826 201134
rect 524062 200898 524146 201134
rect 524382 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 589182 201134
rect 589418 200898 589502 201134
rect 589738 200898 592650 201134
rect -8726 200866 592650 200898
rect -8726 196954 592650 196986
rect -8726 196718 -4854 196954
rect -4618 196718 -4534 196954
rect -4298 196718 15326 196954
rect 15562 196718 15646 196954
rect 15882 196718 51326 196954
rect 51562 196718 51646 196954
rect 51882 196718 87326 196954
rect 87562 196718 87646 196954
rect 87882 196718 123326 196954
rect 123562 196718 123646 196954
rect 123882 196718 159326 196954
rect 159562 196718 159646 196954
rect 159882 196718 195326 196954
rect 195562 196718 195646 196954
rect 195882 196718 231326 196954
rect 231562 196718 231646 196954
rect 231882 196718 267326 196954
rect 267562 196718 267646 196954
rect 267882 196718 303326 196954
rect 303562 196718 303646 196954
rect 303882 196718 339326 196954
rect 339562 196718 339646 196954
rect 339882 196718 375326 196954
rect 375562 196718 375646 196954
rect 375882 196718 411326 196954
rect 411562 196718 411646 196954
rect 411882 196718 447326 196954
rect 447562 196718 447646 196954
rect 447882 196718 483326 196954
rect 483562 196718 483646 196954
rect 483882 196718 519326 196954
rect 519562 196718 519646 196954
rect 519882 196718 555326 196954
rect 555562 196718 555646 196954
rect 555882 196718 588222 196954
rect 588458 196718 588542 196954
rect 588778 196718 592650 196954
rect -8726 196634 592650 196718
rect -8726 196398 -4854 196634
rect -4618 196398 -4534 196634
rect -4298 196398 15326 196634
rect 15562 196398 15646 196634
rect 15882 196398 51326 196634
rect 51562 196398 51646 196634
rect 51882 196398 87326 196634
rect 87562 196398 87646 196634
rect 87882 196398 123326 196634
rect 123562 196398 123646 196634
rect 123882 196398 159326 196634
rect 159562 196398 159646 196634
rect 159882 196398 195326 196634
rect 195562 196398 195646 196634
rect 195882 196398 231326 196634
rect 231562 196398 231646 196634
rect 231882 196398 267326 196634
rect 267562 196398 267646 196634
rect 267882 196398 303326 196634
rect 303562 196398 303646 196634
rect 303882 196398 339326 196634
rect 339562 196398 339646 196634
rect 339882 196398 375326 196634
rect 375562 196398 375646 196634
rect 375882 196398 411326 196634
rect 411562 196398 411646 196634
rect 411882 196398 447326 196634
rect 447562 196398 447646 196634
rect 447882 196398 483326 196634
rect 483562 196398 483646 196634
rect 483882 196398 519326 196634
rect 519562 196398 519646 196634
rect 519882 196398 555326 196634
rect 555562 196398 555646 196634
rect 555882 196398 588222 196634
rect 588458 196398 588542 196634
rect 588778 196398 592650 196634
rect -8726 196366 592650 196398
rect -8726 192454 592650 192486
rect -8726 192218 -3894 192454
rect -3658 192218 -3574 192454
rect -3338 192218 10826 192454
rect 11062 192218 11146 192454
rect 11382 192218 46826 192454
rect 47062 192218 47146 192454
rect 47382 192218 82826 192454
rect 83062 192218 83146 192454
rect 83382 192218 118826 192454
rect 119062 192218 119146 192454
rect 119382 192218 154826 192454
rect 155062 192218 155146 192454
rect 155382 192218 190826 192454
rect 191062 192218 191146 192454
rect 191382 192218 226826 192454
rect 227062 192218 227146 192454
rect 227382 192218 262826 192454
rect 263062 192218 263146 192454
rect 263382 192218 298826 192454
rect 299062 192218 299146 192454
rect 299382 192218 334826 192454
rect 335062 192218 335146 192454
rect 335382 192218 370826 192454
rect 371062 192218 371146 192454
rect 371382 192218 406826 192454
rect 407062 192218 407146 192454
rect 407382 192218 442826 192454
rect 443062 192218 443146 192454
rect 443382 192218 478826 192454
rect 479062 192218 479146 192454
rect 479382 192218 514826 192454
rect 515062 192218 515146 192454
rect 515382 192218 550826 192454
rect 551062 192218 551146 192454
rect 551382 192218 587262 192454
rect 587498 192218 587582 192454
rect 587818 192218 592650 192454
rect -8726 192134 592650 192218
rect -8726 191898 -3894 192134
rect -3658 191898 -3574 192134
rect -3338 191898 10826 192134
rect 11062 191898 11146 192134
rect 11382 191898 46826 192134
rect 47062 191898 47146 192134
rect 47382 191898 82826 192134
rect 83062 191898 83146 192134
rect 83382 191898 118826 192134
rect 119062 191898 119146 192134
rect 119382 191898 154826 192134
rect 155062 191898 155146 192134
rect 155382 191898 190826 192134
rect 191062 191898 191146 192134
rect 191382 191898 226826 192134
rect 227062 191898 227146 192134
rect 227382 191898 262826 192134
rect 263062 191898 263146 192134
rect 263382 191898 298826 192134
rect 299062 191898 299146 192134
rect 299382 191898 334826 192134
rect 335062 191898 335146 192134
rect 335382 191898 370826 192134
rect 371062 191898 371146 192134
rect 371382 191898 406826 192134
rect 407062 191898 407146 192134
rect 407382 191898 442826 192134
rect 443062 191898 443146 192134
rect 443382 191898 478826 192134
rect 479062 191898 479146 192134
rect 479382 191898 514826 192134
rect 515062 191898 515146 192134
rect 515382 191898 550826 192134
rect 551062 191898 551146 192134
rect 551382 191898 587262 192134
rect 587498 191898 587582 192134
rect 587818 191898 592650 192134
rect -8726 191866 592650 191898
rect -8726 187954 592650 187986
rect -8726 187718 -2934 187954
rect -2698 187718 -2614 187954
rect -2378 187718 6326 187954
rect 6562 187718 6646 187954
rect 6882 187718 42326 187954
rect 42562 187718 42646 187954
rect 42882 187718 78326 187954
rect 78562 187718 78646 187954
rect 78882 187718 114326 187954
rect 114562 187718 114646 187954
rect 114882 187718 150326 187954
rect 150562 187718 150646 187954
rect 150882 187718 186326 187954
rect 186562 187718 186646 187954
rect 186882 187718 222326 187954
rect 222562 187718 222646 187954
rect 222882 187718 258326 187954
rect 258562 187718 258646 187954
rect 258882 187718 294326 187954
rect 294562 187718 294646 187954
rect 294882 187718 330326 187954
rect 330562 187718 330646 187954
rect 330882 187718 366326 187954
rect 366562 187718 366646 187954
rect 366882 187718 402326 187954
rect 402562 187718 402646 187954
rect 402882 187718 438326 187954
rect 438562 187718 438646 187954
rect 438882 187718 474326 187954
rect 474562 187718 474646 187954
rect 474882 187718 510326 187954
rect 510562 187718 510646 187954
rect 510882 187718 546326 187954
rect 546562 187718 546646 187954
rect 546882 187718 582326 187954
rect 582562 187718 582646 187954
rect 582882 187718 586302 187954
rect 586538 187718 586622 187954
rect 586858 187718 592650 187954
rect -8726 187634 592650 187718
rect -8726 187398 -2934 187634
rect -2698 187398 -2614 187634
rect -2378 187398 6326 187634
rect 6562 187398 6646 187634
rect 6882 187398 42326 187634
rect 42562 187398 42646 187634
rect 42882 187398 78326 187634
rect 78562 187398 78646 187634
rect 78882 187398 114326 187634
rect 114562 187398 114646 187634
rect 114882 187398 150326 187634
rect 150562 187398 150646 187634
rect 150882 187398 186326 187634
rect 186562 187398 186646 187634
rect 186882 187398 222326 187634
rect 222562 187398 222646 187634
rect 222882 187398 258326 187634
rect 258562 187398 258646 187634
rect 258882 187398 294326 187634
rect 294562 187398 294646 187634
rect 294882 187398 330326 187634
rect 330562 187398 330646 187634
rect 330882 187398 366326 187634
rect 366562 187398 366646 187634
rect 366882 187398 402326 187634
rect 402562 187398 402646 187634
rect 402882 187398 438326 187634
rect 438562 187398 438646 187634
rect 438882 187398 474326 187634
rect 474562 187398 474646 187634
rect 474882 187398 510326 187634
rect 510562 187398 510646 187634
rect 510882 187398 546326 187634
rect 546562 187398 546646 187634
rect 546882 187398 582326 187634
rect 582562 187398 582646 187634
rect 582882 187398 586302 187634
rect 586538 187398 586622 187634
rect 586858 187398 592650 187634
rect -8726 187366 592650 187398
rect -8726 183454 592650 183486
rect -8726 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 73826 183454
rect 74062 183218 74146 183454
rect 74382 183218 109826 183454
rect 110062 183218 110146 183454
rect 110382 183218 145826 183454
rect 146062 183218 146146 183454
rect 146382 183218 181826 183454
rect 182062 183218 182146 183454
rect 182382 183218 217826 183454
rect 218062 183218 218146 183454
rect 218382 183218 253826 183454
rect 254062 183218 254146 183454
rect 254382 183218 289826 183454
rect 290062 183218 290146 183454
rect 290382 183218 325826 183454
rect 326062 183218 326146 183454
rect 326382 183218 361826 183454
rect 362062 183218 362146 183454
rect 362382 183218 397826 183454
rect 398062 183218 398146 183454
rect 398382 183218 433826 183454
rect 434062 183218 434146 183454
rect 434382 183218 469826 183454
rect 470062 183218 470146 183454
rect 470382 183218 505826 183454
rect 506062 183218 506146 183454
rect 506382 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 592650 183454
rect -8726 183134 592650 183218
rect -8726 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 73826 183134
rect 74062 182898 74146 183134
rect 74382 182898 109826 183134
rect 110062 182898 110146 183134
rect 110382 182898 145826 183134
rect 146062 182898 146146 183134
rect 146382 182898 181826 183134
rect 182062 182898 182146 183134
rect 182382 182898 217826 183134
rect 218062 182898 218146 183134
rect 218382 182898 253826 183134
rect 254062 182898 254146 183134
rect 254382 182898 289826 183134
rect 290062 182898 290146 183134
rect 290382 182898 325826 183134
rect 326062 182898 326146 183134
rect 326382 182898 361826 183134
rect 362062 182898 362146 183134
rect 362382 182898 397826 183134
rect 398062 182898 398146 183134
rect 398382 182898 433826 183134
rect 434062 182898 434146 183134
rect 434382 182898 469826 183134
rect 470062 182898 470146 183134
rect 470382 182898 505826 183134
rect 506062 182898 506146 183134
rect 506382 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 592650 183134
rect -8726 182866 592650 182898
rect -8726 178954 592650 178986
rect -8726 178718 -8694 178954
rect -8458 178718 -8374 178954
rect -8138 178718 33326 178954
rect 33562 178718 33646 178954
rect 33882 178718 69326 178954
rect 69562 178718 69646 178954
rect 69882 178718 105326 178954
rect 105562 178718 105646 178954
rect 105882 178718 141326 178954
rect 141562 178718 141646 178954
rect 141882 178718 177326 178954
rect 177562 178718 177646 178954
rect 177882 178718 213326 178954
rect 213562 178718 213646 178954
rect 213882 178718 249326 178954
rect 249562 178718 249646 178954
rect 249882 178718 285326 178954
rect 285562 178718 285646 178954
rect 285882 178718 321326 178954
rect 321562 178718 321646 178954
rect 321882 178718 357326 178954
rect 357562 178718 357646 178954
rect 357882 178718 393326 178954
rect 393562 178718 393646 178954
rect 393882 178718 429326 178954
rect 429562 178718 429646 178954
rect 429882 178718 465326 178954
rect 465562 178718 465646 178954
rect 465882 178718 501326 178954
rect 501562 178718 501646 178954
rect 501882 178718 537326 178954
rect 537562 178718 537646 178954
rect 537882 178718 573326 178954
rect 573562 178718 573646 178954
rect 573882 178718 592062 178954
rect 592298 178718 592382 178954
rect 592618 178718 592650 178954
rect -8726 178634 592650 178718
rect -8726 178398 -8694 178634
rect -8458 178398 -8374 178634
rect -8138 178398 33326 178634
rect 33562 178398 33646 178634
rect 33882 178398 69326 178634
rect 69562 178398 69646 178634
rect 69882 178398 105326 178634
rect 105562 178398 105646 178634
rect 105882 178398 141326 178634
rect 141562 178398 141646 178634
rect 141882 178398 177326 178634
rect 177562 178398 177646 178634
rect 177882 178398 213326 178634
rect 213562 178398 213646 178634
rect 213882 178398 249326 178634
rect 249562 178398 249646 178634
rect 249882 178398 285326 178634
rect 285562 178398 285646 178634
rect 285882 178398 321326 178634
rect 321562 178398 321646 178634
rect 321882 178398 357326 178634
rect 357562 178398 357646 178634
rect 357882 178398 393326 178634
rect 393562 178398 393646 178634
rect 393882 178398 429326 178634
rect 429562 178398 429646 178634
rect 429882 178398 465326 178634
rect 465562 178398 465646 178634
rect 465882 178398 501326 178634
rect 501562 178398 501646 178634
rect 501882 178398 537326 178634
rect 537562 178398 537646 178634
rect 537882 178398 573326 178634
rect 573562 178398 573646 178634
rect 573882 178398 592062 178634
rect 592298 178398 592382 178634
rect 592618 178398 592650 178634
rect -8726 178366 592650 178398
rect -8726 174454 592650 174486
rect -8726 174218 -7734 174454
rect -7498 174218 -7414 174454
rect -7178 174218 28826 174454
rect 29062 174218 29146 174454
rect 29382 174218 64826 174454
rect 65062 174218 65146 174454
rect 65382 174218 100826 174454
rect 101062 174218 101146 174454
rect 101382 174218 208826 174454
rect 209062 174218 209146 174454
rect 209382 174218 244826 174454
rect 245062 174218 245146 174454
rect 245382 174218 280826 174454
rect 281062 174218 281146 174454
rect 281382 174218 316826 174454
rect 317062 174218 317146 174454
rect 317382 174218 352826 174454
rect 353062 174218 353146 174454
rect 353382 174218 388826 174454
rect 389062 174218 389146 174454
rect 389382 174218 424826 174454
rect 425062 174218 425146 174454
rect 425382 174218 460826 174454
rect 461062 174218 461146 174454
rect 461382 174218 496826 174454
rect 497062 174218 497146 174454
rect 497382 174218 532826 174454
rect 533062 174218 533146 174454
rect 533382 174218 568826 174454
rect 569062 174218 569146 174454
rect 569382 174218 591102 174454
rect 591338 174218 591422 174454
rect 591658 174218 592650 174454
rect -8726 174134 592650 174218
rect -8726 173898 -7734 174134
rect -7498 173898 -7414 174134
rect -7178 173898 28826 174134
rect 29062 173898 29146 174134
rect 29382 173898 64826 174134
rect 65062 173898 65146 174134
rect 65382 173898 100826 174134
rect 101062 173898 101146 174134
rect 101382 173898 208826 174134
rect 209062 173898 209146 174134
rect 209382 173898 244826 174134
rect 245062 173898 245146 174134
rect 245382 173898 280826 174134
rect 281062 173898 281146 174134
rect 281382 173898 316826 174134
rect 317062 173898 317146 174134
rect 317382 173898 352826 174134
rect 353062 173898 353146 174134
rect 353382 173898 388826 174134
rect 389062 173898 389146 174134
rect 389382 173898 424826 174134
rect 425062 173898 425146 174134
rect 425382 173898 460826 174134
rect 461062 173898 461146 174134
rect 461382 173898 496826 174134
rect 497062 173898 497146 174134
rect 497382 173898 532826 174134
rect 533062 173898 533146 174134
rect 533382 173898 568826 174134
rect 569062 173898 569146 174134
rect 569382 173898 591102 174134
rect 591338 173898 591422 174134
rect 591658 173898 592650 174134
rect -8726 173866 592650 173898
rect -8726 169954 592650 169986
rect -8726 169718 -6774 169954
rect -6538 169718 -6454 169954
rect -6218 169718 24326 169954
rect 24562 169718 24646 169954
rect 24882 169718 60326 169954
rect 60562 169718 60646 169954
rect 60882 169718 96326 169954
rect 96562 169718 96646 169954
rect 96882 169718 204326 169954
rect 204562 169718 204646 169954
rect 204882 169718 240326 169954
rect 240562 169718 240646 169954
rect 240882 169718 276326 169954
rect 276562 169718 276646 169954
rect 276882 169718 312326 169954
rect 312562 169718 312646 169954
rect 312882 169718 348326 169954
rect 348562 169718 348646 169954
rect 348882 169718 384326 169954
rect 384562 169718 384646 169954
rect 384882 169718 420326 169954
rect 420562 169718 420646 169954
rect 420882 169718 456326 169954
rect 456562 169718 456646 169954
rect 456882 169718 492326 169954
rect 492562 169718 492646 169954
rect 492882 169718 528326 169954
rect 528562 169718 528646 169954
rect 528882 169718 564326 169954
rect 564562 169718 564646 169954
rect 564882 169718 590142 169954
rect 590378 169718 590462 169954
rect 590698 169718 592650 169954
rect -8726 169634 592650 169718
rect -8726 169398 -6774 169634
rect -6538 169398 -6454 169634
rect -6218 169398 24326 169634
rect 24562 169398 24646 169634
rect 24882 169398 60326 169634
rect 60562 169398 60646 169634
rect 60882 169398 96326 169634
rect 96562 169398 96646 169634
rect 96882 169398 204326 169634
rect 204562 169398 204646 169634
rect 204882 169398 240326 169634
rect 240562 169398 240646 169634
rect 240882 169398 276326 169634
rect 276562 169398 276646 169634
rect 276882 169398 312326 169634
rect 312562 169398 312646 169634
rect 312882 169398 348326 169634
rect 348562 169398 348646 169634
rect 348882 169398 384326 169634
rect 384562 169398 384646 169634
rect 384882 169398 420326 169634
rect 420562 169398 420646 169634
rect 420882 169398 456326 169634
rect 456562 169398 456646 169634
rect 456882 169398 492326 169634
rect 492562 169398 492646 169634
rect 492882 169398 528326 169634
rect 528562 169398 528646 169634
rect 528882 169398 564326 169634
rect 564562 169398 564646 169634
rect 564882 169398 590142 169634
rect 590378 169398 590462 169634
rect 590698 169398 592650 169634
rect -8726 169366 592650 169398
rect -8726 165454 592650 165486
rect -8726 165218 -5814 165454
rect -5578 165218 -5494 165454
rect -5258 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 55826 165454
rect 56062 165218 56146 165454
rect 56382 165218 91826 165454
rect 92062 165218 92146 165454
rect 92382 165218 199826 165454
rect 200062 165218 200146 165454
rect 200382 165218 235826 165454
rect 236062 165218 236146 165454
rect 236382 165218 271826 165454
rect 272062 165218 272146 165454
rect 272382 165218 307826 165454
rect 308062 165218 308146 165454
rect 308382 165218 343826 165454
rect 344062 165218 344146 165454
rect 344382 165218 379826 165454
rect 380062 165218 380146 165454
rect 380382 165218 415826 165454
rect 416062 165218 416146 165454
rect 416382 165218 451826 165454
rect 452062 165218 452146 165454
rect 452382 165218 487826 165454
rect 488062 165218 488146 165454
rect 488382 165218 523826 165454
rect 524062 165218 524146 165454
rect 524382 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 589182 165454
rect 589418 165218 589502 165454
rect 589738 165218 592650 165454
rect -8726 165134 592650 165218
rect -8726 164898 -5814 165134
rect -5578 164898 -5494 165134
rect -5258 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 55826 165134
rect 56062 164898 56146 165134
rect 56382 164898 91826 165134
rect 92062 164898 92146 165134
rect 92382 164898 199826 165134
rect 200062 164898 200146 165134
rect 200382 164898 235826 165134
rect 236062 164898 236146 165134
rect 236382 164898 271826 165134
rect 272062 164898 272146 165134
rect 272382 164898 307826 165134
rect 308062 164898 308146 165134
rect 308382 164898 343826 165134
rect 344062 164898 344146 165134
rect 344382 164898 379826 165134
rect 380062 164898 380146 165134
rect 380382 164898 415826 165134
rect 416062 164898 416146 165134
rect 416382 164898 451826 165134
rect 452062 164898 452146 165134
rect 452382 164898 487826 165134
rect 488062 164898 488146 165134
rect 488382 164898 523826 165134
rect 524062 164898 524146 165134
rect 524382 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 589182 165134
rect 589418 164898 589502 165134
rect 589738 164898 592650 165134
rect -8726 164866 592650 164898
rect -8726 160954 592650 160986
rect -8726 160718 -4854 160954
rect -4618 160718 -4534 160954
rect -4298 160718 15326 160954
rect 15562 160718 15646 160954
rect 15882 160718 51326 160954
rect 51562 160718 51646 160954
rect 51882 160718 87326 160954
rect 87562 160718 87646 160954
rect 87882 160718 123326 160954
rect 123562 160718 123646 160954
rect 123882 160718 159326 160954
rect 159562 160718 159646 160954
rect 159882 160718 195326 160954
rect 195562 160718 195646 160954
rect 195882 160718 231326 160954
rect 231562 160718 231646 160954
rect 231882 160718 267326 160954
rect 267562 160718 267646 160954
rect 267882 160718 303326 160954
rect 303562 160718 303646 160954
rect 303882 160718 339326 160954
rect 339562 160718 339646 160954
rect 339882 160718 375326 160954
rect 375562 160718 375646 160954
rect 375882 160718 411326 160954
rect 411562 160718 411646 160954
rect 411882 160718 447326 160954
rect 447562 160718 447646 160954
rect 447882 160718 483326 160954
rect 483562 160718 483646 160954
rect 483882 160718 519326 160954
rect 519562 160718 519646 160954
rect 519882 160718 555326 160954
rect 555562 160718 555646 160954
rect 555882 160718 588222 160954
rect 588458 160718 588542 160954
rect 588778 160718 592650 160954
rect -8726 160634 592650 160718
rect -8726 160398 -4854 160634
rect -4618 160398 -4534 160634
rect -4298 160398 15326 160634
rect 15562 160398 15646 160634
rect 15882 160398 51326 160634
rect 51562 160398 51646 160634
rect 51882 160398 87326 160634
rect 87562 160398 87646 160634
rect 87882 160398 123326 160634
rect 123562 160398 123646 160634
rect 123882 160398 159326 160634
rect 159562 160398 159646 160634
rect 159882 160398 195326 160634
rect 195562 160398 195646 160634
rect 195882 160398 231326 160634
rect 231562 160398 231646 160634
rect 231882 160398 267326 160634
rect 267562 160398 267646 160634
rect 267882 160398 303326 160634
rect 303562 160398 303646 160634
rect 303882 160398 339326 160634
rect 339562 160398 339646 160634
rect 339882 160398 375326 160634
rect 375562 160398 375646 160634
rect 375882 160398 411326 160634
rect 411562 160398 411646 160634
rect 411882 160398 447326 160634
rect 447562 160398 447646 160634
rect 447882 160398 483326 160634
rect 483562 160398 483646 160634
rect 483882 160398 519326 160634
rect 519562 160398 519646 160634
rect 519882 160398 555326 160634
rect 555562 160398 555646 160634
rect 555882 160398 588222 160634
rect 588458 160398 588542 160634
rect 588778 160398 592650 160634
rect -8726 160366 592650 160398
rect -8726 156454 592650 156486
rect -8726 156218 -3894 156454
rect -3658 156218 -3574 156454
rect -3338 156218 10826 156454
rect 11062 156218 11146 156454
rect 11382 156218 46826 156454
rect 47062 156218 47146 156454
rect 47382 156218 82826 156454
rect 83062 156218 83146 156454
rect 83382 156218 118826 156454
rect 119062 156218 119146 156454
rect 119382 156218 154826 156454
rect 155062 156218 155146 156454
rect 155382 156218 190826 156454
rect 191062 156218 191146 156454
rect 191382 156218 226826 156454
rect 227062 156218 227146 156454
rect 227382 156218 262826 156454
rect 263062 156218 263146 156454
rect 263382 156218 298826 156454
rect 299062 156218 299146 156454
rect 299382 156218 334826 156454
rect 335062 156218 335146 156454
rect 335382 156218 370826 156454
rect 371062 156218 371146 156454
rect 371382 156218 406826 156454
rect 407062 156218 407146 156454
rect 407382 156218 442826 156454
rect 443062 156218 443146 156454
rect 443382 156218 478826 156454
rect 479062 156218 479146 156454
rect 479382 156218 514826 156454
rect 515062 156218 515146 156454
rect 515382 156218 550826 156454
rect 551062 156218 551146 156454
rect 551382 156218 587262 156454
rect 587498 156218 587582 156454
rect 587818 156218 592650 156454
rect -8726 156134 592650 156218
rect -8726 155898 -3894 156134
rect -3658 155898 -3574 156134
rect -3338 155898 10826 156134
rect 11062 155898 11146 156134
rect 11382 155898 46826 156134
rect 47062 155898 47146 156134
rect 47382 155898 82826 156134
rect 83062 155898 83146 156134
rect 83382 155898 118826 156134
rect 119062 155898 119146 156134
rect 119382 155898 154826 156134
rect 155062 155898 155146 156134
rect 155382 155898 190826 156134
rect 191062 155898 191146 156134
rect 191382 155898 226826 156134
rect 227062 155898 227146 156134
rect 227382 155898 262826 156134
rect 263062 155898 263146 156134
rect 263382 155898 298826 156134
rect 299062 155898 299146 156134
rect 299382 155898 334826 156134
rect 335062 155898 335146 156134
rect 335382 155898 370826 156134
rect 371062 155898 371146 156134
rect 371382 155898 406826 156134
rect 407062 155898 407146 156134
rect 407382 155898 442826 156134
rect 443062 155898 443146 156134
rect 443382 155898 478826 156134
rect 479062 155898 479146 156134
rect 479382 155898 514826 156134
rect 515062 155898 515146 156134
rect 515382 155898 550826 156134
rect 551062 155898 551146 156134
rect 551382 155898 587262 156134
rect 587498 155898 587582 156134
rect 587818 155898 592650 156134
rect -8726 155866 592650 155898
rect -8726 151954 592650 151986
rect -8726 151718 -2934 151954
rect -2698 151718 -2614 151954
rect -2378 151718 6326 151954
rect 6562 151718 6646 151954
rect 6882 151718 42326 151954
rect 42562 151718 42646 151954
rect 42882 151718 78326 151954
rect 78562 151718 78646 151954
rect 78882 151718 114326 151954
rect 114562 151718 114646 151954
rect 114882 151718 150326 151954
rect 150562 151718 150646 151954
rect 150882 151718 186326 151954
rect 186562 151718 186646 151954
rect 186882 151718 222326 151954
rect 222562 151718 222646 151954
rect 222882 151718 258326 151954
rect 258562 151718 258646 151954
rect 258882 151718 294326 151954
rect 294562 151718 294646 151954
rect 294882 151718 330326 151954
rect 330562 151718 330646 151954
rect 330882 151718 366326 151954
rect 366562 151718 366646 151954
rect 366882 151718 402326 151954
rect 402562 151718 402646 151954
rect 402882 151718 438326 151954
rect 438562 151718 438646 151954
rect 438882 151718 474326 151954
rect 474562 151718 474646 151954
rect 474882 151718 510326 151954
rect 510562 151718 510646 151954
rect 510882 151718 546326 151954
rect 546562 151718 546646 151954
rect 546882 151718 582326 151954
rect 582562 151718 582646 151954
rect 582882 151718 586302 151954
rect 586538 151718 586622 151954
rect 586858 151718 592650 151954
rect -8726 151634 592650 151718
rect -8726 151398 -2934 151634
rect -2698 151398 -2614 151634
rect -2378 151398 6326 151634
rect 6562 151398 6646 151634
rect 6882 151398 42326 151634
rect 42562 151398 42646 151634
rect 42882 151398 78326 151634
rect 78562 151398 78646 151634
rect 78882 151398 114326 151634
rect 114562 151398 114646 151634
rect 114882 151398 150326 151634
rect 150562 151398 150646 151634
rect 150882 151398 186326 151634
rect 186562 151398 186646 151634
rect 186882 151398 222326 151634
rect 222562 151398 222646 151634
rect 222882 151398 258326 151634
rect 258562 151398 258646 151634
rect 258882 151398 294326 151634
rect 294562 151398 294646 151634
rect 294882 151398 330326 151634
rect 330562 151398 330646 151634
rect 330882 151398 366326 151634
rect 366562 151398 366646 151634
rect 366882 151398 402326 151634
rect 402562 151398 402646 151634
rect 402882 151398 438326 151634
rect 438562 151398 438646 151634
rect 438882 151398 474326 151634
rect 474562 151398 474646 151634
rect 474882 151398 510326 151634
rect 510562 151398 510646 151634
rect 510882 151398 546326 151634
rect 546562 151398 546646 151634
rect 546882 151398 582326 151634
rect 582562 151398 582646 151634
rect 582882 151398 586302 151634
rect 586538 151398 586622 151634
rect 586858 151398 592650 151634
rect -8726 151366 592650 151398
rect -8726 147454 592650 147486
rect -8726 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 73826 147454
rect 74062 147218 74146 147454
rect 74382 147218 109826 147454
rect 110062 147218 110146 147454
rect 110382 147218 145826 147454
rect 146062 147218 146146 147454
rect 146382 147218 181826 147454
rect 182062 147218 182146 147454
rect 182382 147218 217826 147454
rect 218062 147218 218146 147454
rect 218382 147218 253826 147454
rect 254062 147218 254146 147454
rect 254382 147218 289826 147454
rect 290062 147218 290146 147454
rect 290382 147218 325826 147454
rect 326062 147218 326146 147454
rect 326382 147218 361826 147454
rect 362062 147218 362146 147454
rect 362382 147218 397826 147454
rect 398062 147218 398146 147454
rect 398382 147218 433826 147454
rect 434062 147218 434146 147454
rect 434382 147218 469826 147454
rect 470062 147218 470146 147454
rect 470382 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 592650 147454
rect -8726 147134 592650 147218
rect -8726 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 73826 147134
rect 74062 146898 74146 147134
rect 74382 146898 109826 147134
rect 110062 146898 110146 147134
rect 110382 146898 145826 147134
rect 146062 146898 146146 147134
rect 146382 146898 181826 147134
rect 182062 146898 182146 147134
rect 182382 146898 217826 147134
rect 218062 146898 218146 147134
rect 218382 146898 253826 147134
rect 254062 146898 254146 147134
rect 254382 146898 289826 147134
rect 290062 146898 290146 147134
rect 290382 146898 325826 147134
rect 326062 146898 326146 147134
rect 326382 146898 361826 147134
rect 362062 146898 362146 147134
rect 362382 146898 397826 147134
rect 398062 146898 398146 147134
rect 398382 146898 433826 147134
rect 434062 146898 434146 147134
rect 434382 146898 469826 147134
rect 470062 146898 470146 147134
rect 470382 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 592650 147134
rect -8726 146866 592650 146898
rect -8726 142954 592650 142986
rect -8726 142718 -8694 142954
rect -8458 142718 -8374 142954
rect -8138 142718 33326 142954
rect 33562 142718 33646 142954
rect 33882 142718 69326 142954
rect 69562 142718 69646 142954
rect 69882 142718 105326 142954
rect 105562 142718 105646 142954
rect 105882 142718 141326 142954
rect 141562 142718 141646 142954
rect 141882 142718 177326 142954
rect 177562 142718 177646 142954
rect 177882 142718 213326 142954
rect 213562 142718 213646 142954
rect 213882 142718 249326 142954
rect 249562 142718 249646 142954
rect 249882 142718 285326 142954
rect 285562 142718 285646 142954
rect 285882 142718 321326 142954
rect 321562 142718 321646 142954
rect 321882 142718 357326 142954
rect 357562 142718 357646 142954
rect 357882 142718 393326 142954
rect 393562 142718 393646 142954
rect 393882 142718 429326 142954
rect 429562 142718 429646 142954
rect 429882 142718 465326 142954
rect 465562 142718 465646 142954
rect 465882 142718 501326 142954
rect 501562 142718 501646 142954
rect 501882 142718 537326 142954
rect 537562 142718 537646 142954
rect 537882 142718 573326 142954
rect 573562 142718 573646 142954
rect 573882 142718 592062 142954
rect 592298 142718 592382 142954
rect 592618 142718 592650 142954
rect -8726 142634 592650 142718
rect -8726 142398 -8694 142634
rect -8458 142398 -8374 142634
rect -8138 142398 33326 142634
rect 33562 142398 33646 142634
rect 33882 142398 69326 142634
rect 69562 142398 69646 142634
rect 69882 142398 105326 142634
rect 105562 142398 105646 142634
rect 105882 142398 141326 142634
rect 141562 142398 141646 142634
rect 141882 142398 177326 142634
rect 177562 142398 177646 142634
rect 177882 142398 213326 142634
rect 213562 142398 213646 142634
rect 213882 142398 249326 142634
rect 249562 142398 249646 142634
rect 249882 142398 285326 142634
rect 285562 142398 285646 142634
rect 285882 142398 321326 142634
rect 321562 142398 321646 142634
rect 321882 142398 357326 142634
rect 357562 142398 357646 142634
rect 357882 142398 393326 142634
rect 393562 142398 393646 142634
rect 393882 142398 429326 142634
rect 429562 142398 429646 142634
rect 429882 142398 465326 142634
rect 465562 142398 465646 142634
rect 465882 142398 501326 142634
rect 501562 142398 501646 142634
rect 501882 142398 537326 142634
rect 537562 142398 537646 142634
rect 537882 142398 573326 142634
rect 573562 142398 573646 142634
rect 573882 142398 592062 142634
rect 592298 142398 592382 142634
rect 592618 142398 592650 142634
rect -8726 142366 592650 142398
rect -8726 138454 592650 138486
rect -8726 138218 -7734 138454
rect -7498 138218 -7414 138454
rect -7178 138218 28826 138454
rect 29062 138218 29146 138454
rect 29382 138218 64826 138454
rect 65062 138218 65146 138454
rect 65382 138218 100826 138454
rect 101062 138218 101146 138454
rect 101382 138218 208826 138454
rect 209062 138218 209146 138454
rect 209382 138218 244826 138454
rect 245062 138218 245146 138454
rect 245382 138218 280826 138454
rect 281062 138218 281146 138454
rect 281382 138218 316826 138454
rect 317062 138218 317146 138454
rect 317382 138218 352826 138454
rect 353062 138218 353146 138454
rect 353382 138218 388826 138454
rect 389062 138218 389146 138454
rect 389382 138218 424826 138454
rect 425062 138218 425146 138454
rect 425382 138218 460826 138454
rect 461062 138218 461146 138454
rect 461382 138218 496826 138454
rect 497062 138218 497146 138454
rect 497382 138218 532826 138454
rect 533062 138218 533146 138454
rect 533382 138218 568826 138454
rect 569062 138218 569146 138454
rect 569382 138218 591102 138454
rect 591338 138218 591422 138454
rect 591658 138218 592650 138454
rect -8726 138134 592650 138218
rect -8726 137898 -7734 138134
rect -7498 137898 -7414 138134
rect -7178 137898 28826 138134
rect 29062 137898 29146 138134
rect 29382 137898 64826 138134
rect 65062 137898 65146 138134
rect 65382 137898 100826 138134
rect 101062 137898 101146 138134
rect 101382 137898 208826 138134
rect 209062 137898 209146 138134
rect 209382 137898 244826 138134
rect 245062 137898 245146 138134
rect 245382 137898 280826 138134
rect 281062 137898 281146 138134
rect 281382 137898 316826 138134
rect 317062 137898 317146 138134
rect 317382 137898 352826 138134
rect 353062 137898 353146 138134
rect 353382 137898 388826 138134
rect 389062 137898 389146 138134
rect 389382 137898 424826 138134
rect 425062 137898 425146 138134
rect 425382 137898 460826 138134
rect 461062 137898 461146 138134
rect 461382 137898 496826 138134
rect 497062 137898 497146 138134
rect 497382 137898 532826 138134
rect 533062 137898 533146 138134
rect 533382 137898 568826 138134
rect 569062 137898 569146 138134
rect 569382 137898 591102 138134
rect 591338 137898 591422 138134
rect 591658 137898 592650 138134
rect -8726 137866 592650 137898
rect -8726 133954 592650 133986
rect -8726 133718 -6774 133954
rect -6538 133718 -6454 133954
rect -6218 133718 24326 133954
rect 24562 133718 24646 133954
rect 24882 133718 60326 133954
rect 60562 133718 60646 133954
rect 60882 133718 96326 133954
rect 96562 133718 96646 133954
rect 96882 133718 204326 133954
rect 204562 133718 204646 133954
rect 204882 133718 240326 133954
rect 240562 133718 240646 133954
rect 240882 133718 276326 133954
rect 276562 133718 276646 133954
rect 276882 133718 312326 133954
rect 312562 133718 312646 133954
rect 312882 133718 348326 133954
rect 348562 133718 348646 133954
rect 348882 133718 384326 133954
rect 384562 133718 384646 133954
rect 384882 133718 420326 133954
rect 420562 133718 420646 133954
rect 420882 133718 456326 133954
rect 456562 133718 456646 133954
rect 456882 133718 492326 133954
rect 492562 133718 492646 133954
rect 492882 133718 528326 133954
rect 528562 133718 528646 133954
rect 528882 133718 564326 133954
rect 564562 133718 564646 133954
rect 564882 133718 590142 133954
rect 590378 133718 590462 133954
rect 590698 133718 592650 133954
rect -8726 133634 592650 133718
rect -8726 133398 -6774 133634
rect -6538 133398 -6454 133634
rect -6218 133398 24326 133634
rect 24562 133398 24646 133634
rect 24882 133398 60326 133634
rect 60562 133398 60646 133634
rect 60882 133398 96326 133634
rect 96562 133398 96646 133634
rect 96882 133398 204326 133634
rect 204562 133398 204646 133634
rect 204882 133398 240326 133634
rect 240562 133398 240646 133634
rect 240882 133398 276326 133634
rect 276562 133398 276646 133634
rect 276882 133398 312326 133634
rect 312562 133398 312646 133634
rect 312882 133398 348326 133634
rect 348562 133398 348646 133634
rect 348882 133398 384326 133634
rect 384562 133398 384646 133634
rect 384882 133398 420326 133634
rect 420562 133398 420646 133634
rect 420882 133398 456326 133634
rect 456562 133398 456646 133634
rect 456882 133398 492326 133634
rect 492562 133398 492646 133634
rect 492882 133398 528326 133634
rect 528562 133398 528646 133634
rect 528882 133398 564326 133634
rect 564562 133398 564646 133634
rect 564882 133398 590142 133634
rect 590378 133398 590462 133634
rect 590698 133398 592650 133634
rect -8726 133366 592650 133398
rect -8726 129454 592650 129486
rect -8726 129218 -5814 129454
rect -5578 129218 -5494 129454
rect -5258 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 55826 129454
rect 56062 129218 56146 129454
rect 56382 129218 91826 129454
rect 92062 129218 92146 129454
rect 92382 129218 199826 129454
rect 200062 129218 200146 129454
rect 200382 129218 235826 129454
rect 236062 129218 236146 129454
rect 236382 129218 271826 129454
rect 272062 129218 272146 129454
rect 272382 129218 307826 129454
rect 308062 129218 308146 129454
rect 308382 129218 343826 129454
rect 344062 129218 344146 129454
rect 344382 129218 379826 129454
rect 380062 129218 380146 129454
rect 380382 129218 415826 129454
rect 416062 129218 416146 129454
rect 416382 129218 451826 129454
rect 452062 129218 452146 129454
rect 452382 129218 487826 129454
rect 488062 129218 488146 129454
rect 488382 129218 523826 129454
rect 524062 129218 524146 129454
rect 524382 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 589182 129454
rect 589418 129218 589502 129454
rect 589738 129218 592650 129454
rect -8726 129134 592650 129218
rect -8726 128898 -5814 129134
rect -5578 128898 -5494 129134
rect -5258 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 55826 129134
rect 56062 128898 56146 129134
rect 56382 128898 91826 129134
rect 92062 128898 92146 129134
rect 92382 128898 199826 129134
rect 200062 128898 200146 129134
rect 200382 128898 235826 129134
rect 236062 128898 236146 129134
rect 236382 128898 271826 129134
rect 272062 128898 272146 129134
rect 272382 128898 307826 129134
rect 308062 128898 308146 129134
rect 308382 128898 343826 129134
rect 344062 128898 344146 129134
rect 344382 128898 379826 129134
rect 380062 128898 380146 129134
rect 380382 128898 415826 129134
rect 416062 128898 416146 129134
rect 416382 128898 451826 129134
rect 452062 128898 452146 129134
rect 452382 128898 487826 129134
rect 488062 128898 488146 129134
rect 488382 128898 523826 129134
rect 524062 128898 524146 129134
rect 524382 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 589182 129134
rect 589418 128898 589502 129134
rect 589738 128898 592650 129134
rect -8726 128866 592650 128898
rect -8726 124954 592650 124986
rect -8726 124718 -4854 124954
rect -4618 124718 -4534 124954
rect -4298 124718 15326 124954
rect 15562 124718 15646 124954
rect 15882 124718 51326 124954
rect 51562 124718 51646 124954
rect 51882 124718 87326 124954
rect 87562 124718 87646 124954
rect 87882 124718 195326 124954
rect 195562 124718 195646 124954
rect 195882 124718 231326 124954
rect 231562 124718 231646 124954
rect 231882 124718 267326 124954
rect 267562 124718 267646 124954
rect 267882 124718 303326 124954
rect 303562 124718 303646 124954
rect 303882 124718 339326 124954
rect 339562 124718 339646 124954
rect 339882 124718 375326 124954
rect 375562 124718 375646 124954
rect 375882 124718 411326 124954
rect 411562 124718 411646 124954
rect 411882 124718 447326 124954
rect 447562 124718 447646 124954
rect 447882 124718 483326 124954
rect 483562 124718 483646 124954
rect 483882 124718 519326 124954
rect 519562 124718 519646 124954
rect 519882 124718 555326 124954
rect 555562 124718 555646 124954
rect 555882 124718 588222 124954
rect 588458 124718 588542 124954
rect 588778 124718 592650 124954
rect -8726 124634 592650 124718
rect -8726 124398 -4854 124634
rect -4618 124398 -4534 124634
rect -4298 124398 15326 124634
rect 15562 124398 15646 124634
rect 15882 124398 51326 124634
rect 51562 124398 51646 124634
rect 51882 124398 87326 124634
rect 87562 124398 87646 124634
rect 87882 124398 195326 124634
rect 195562 124398 195646 124634
rect 195882 124398 231326 124634
rect 231562 124398 231646 124634
rect 231882 124398 267326 124634
rect 267562 124398 267646 124634
rect 267882 124398 303326 124634
rect 303562 124398 303646 124634
rect 303882 124398 339326 124634
rect 339562 124398 339646 124634
rect 339882 124398 375326 124634
rect 375562 124398 375646 124634
rect 375882 124398 411326 124634
rect 411562 124398 411646 124634
rect 411882 124398 447326 124634
rect 447562 124398 447646 124634
rect 447882 124398 483326 124634
rect 483562 124398 483646 124634
rect 483882 124398 519326 124634
rect 519562 124398 519646 124634
rect 519882 124398 555326 124634
rect 555562 124398 555646 124634
rect 555882 124398 588222 124634
rect 588458 124398 588542 124634
rect 588778 124398 592650 124634
rect -8726 124366 592650 124398
rect -8726 120454 592650 120486
rect -8726 120218 -3894 120454
rect -3658 120218 -3574 120454
rect -3338 120218 10826 120454
rect 11062 120218 11146 120454
rect 11382 120218 46826 120454
rect 47062 120218 47146 120454
rect 47382 120218 82826 120454
rect 83062 120218 83146 120454
rect 83382 120218 226826 120454
rect 227062 120218 227146 120454
rect 227382 120218 262826 120454
rect 263062 120218 263146 120454
rect 263382 120218 298826 120454
rect 299062 120218 299146 120454
rect 299382 120218 334826 120454
rect 335062 120218 335146 120454
rect 335382 120218 370826 120454
rect 371062 120218 371146 120454
rect 371382 120218 406826 120454
rect 407062 120218 407146 120454
rect 407382 120218 442826 120454
rect 443062 120218 443146 120454
rect 443382 120218 478826 120454
rect 479062 120218 479146 120454
rect 479382 120218 514826 120454
rect 515062 120218 515146 120454
rect 515382 120218 550826 120454
rect 551062 120218 551146 120454
rect 551382 120218 587262 120454
rect 587498 120218 587582 120454
rect 587818 120218 592650 120454
rect -8726 120134 592650 120218
rect -8726 119898 -3894 120134
rect -3658 119898 -3574 120134
rect -3338 119898 10826 120134
rect 11062 119898 11146 120134
rect 11382 119898 46826 120134
rect 47062 119898 47146 120134
rect 47382 119898 82826 120134
rect 83062 119898 83146 120134
rect 83382 119898 226826 120134
rect 227062 119898 227146 120134
rect 227382 119898 262826 120134
rect 263062 119898 263146 120134
rect 263382 119898 298826 120134
rect 299062 119898 299146 120134
rect 299382 119898 334826 120134
rect 335062 119898 335146 120134
rect 335382 119898 370826 120134
rect 371062 119898 371146 120134
rect 371382 119898 406826 120134
rect 407062 119898 407146 120134
rect 407382 119898 442826 120134
rect 443062 119898 443146 120134
rect 443382 119898 478826 120134
rect 479062 119898 479146 120134
rect 479382 119898 514826 120134
rect 515062 119898 515146 120134
rect 515382 119898 550826 120134
rect 551062 119898 551146 120134
rect 551382 119898 587262 120134
rect 587498 119898 587582 120134
rect 587818 119898 592650 120134
rect -8726 119866 592650 119898
rect -8726 115954 592650 115986
rect -8726 115718 -2934 115954
rect -2698 115718 -2614 115954
rect -2378 115718 6326 115954
rect 6562 115718 6646 115954
rect 6882 115718 42326 115954
rect 42562 115718 42646 115954
rect 42882 115718 78326 115954
rect 78562 115718 78646 115954
rect 78882 115718 114326 115954
rect 114562 115718 114646 115954
rect 114882 115718 139610 115954
rect 139846 115718 170330 115954
rect 170566 115718 222326 115954
rect 222562 115718 222646 115954
rect 222882 115718 258326 115954
rect 258562 115718 258646 115954
rect 258882 115718 294326 115954
rect 294562 115718 294646 115954
rect 294882 115718 330326 115954
rect 330562 115718 330646 115954
rect 330882 115718 366326 115954
rect 366562 115718 366646 115954
rect 366882 115718 402326 115954
rect 402562 115718 402646 115954
rect 402882 115718 438326 115954
rect 438562 115718 438646 115954
rect 438882 115718 474326 115954
rect 474562 115718 474646 115954
rect 474882 115718 510326 115954
rect 510562 115718 510646 115954
rect 510882 115718 546326 115954
rect 546562 115718 546646 115954
rect 546882 115718 582326 115954
rect 582562 115718 582646 115954
rect 582882 115718 586302 115954
rect 586538 115718 586622 115954
rect 586858 115718 592650 115954
rect -8726 115634 592650 115718
rect -8726 115398 -2934 115634
rect -2698 115398 -2614 115634
rect -2378 115398 6326 115634
rect 6562 115398 6646 115634
rect 6882 115398 42326 115634
rect 42562 115398 42646 115634
rect 42882 115398 78326 115634
rect 78562 115398 78646 115634
rect 78882 115398 114326 115634
rect 114562 115398 114646 115634
rect 114882 115398 139610 115634
rect 139846 115398 170330 115634
rect 170566 115398 222326 115634
rect 222562 115398 222646 115634
rect 222882 115398 258326 115634
rect 258562 115398 258646 115634
rect 258882 115398 294326 115634
rect 294562 115398 294646 115634
rect 294882 115398 330326 115634
rect 330562 115398 330646 115634
rect 330882 115398 366326 115634
rect 366562 115398 366646 115634
rect 366882 115398 402326 115634
rect 402562 115398 402646 115634
rect 402882 115398 438326 115634
rect 438562 115398 438646 115634
rect 438882 115398 474326 115634
rect 474562 115398 474646 115634
rect 474882 115398 510326 115634
rect 510562 115398 510646 115634
rect 510882 115398 546326 115634
rect 546562 115398 546646 115634
rect 546882 115398 582326 115634
rect 582562 115398 582646 115634
rect 582882 115398 586302 115634
rect 586538 115398 586622 115634
rect 586858 115398 592650 115634
rect -8726 115366 592650 115398
rect -8726 111454 592650 111486
rect -8726 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 73826 111454
rect 74062 111218 74146 111454
rect 74382 111218 109826 111454
rect 110062 111218 110146 111454
rect 110382 111218 124250 111454
rect 124486 111218 154970 111454
rect 155206 111218 185690 111454
rect 185926 111218 217826 111454
rect 218062 111218 218146 111454
rect 218382 111218 253826 111454
rect 254062 111218 254146 111454
rect 254382 111218 289826 111454
rect 290062 111218 290146 111454
rect 290382 111218 325826 111454
rect 326062 111218 326146 111454
rect 326382 111218 361826 111454
rect 362062 111218 362146 111454
rect 362382 111218 397826 111454
rect 398062 111218 398146 111454
rect 398382 111218 433826 111454
rect 434062 111218 434146 111454
rect 434382 111218 469826 111454
rect 470062 111218 470146 111454
rect 470382 111218 505826 111454
rect 506062 111218 506146 111454
rect 506382 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 592650 111454
rect -8726 111134 592650 111218
rect -8726 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 73826 111134
rect 74062 110898 74146 111134
rect 74382 110898 109826 111134
rect 110062 110898 110146 111134
rect 110382 110898 124250 111134
rect 124486 110898 154970 111134
rect 155206 110898 185690 111134
rect 185926 110898 217826 111134
rect 218062 110898 218146 111134
rect 218382 110898 253826 111134
rect 254062 110898 254146 111134
rect 254382 110898 289826 111134
rect 290062 110898 290146 111134
rect 290382 110898 325826 111134
rect 326062 110898 326146 111134
rect 326382 110898 361826 111134
rect 362062 110898 362146 111134
rect 362382 110898 397826 111134
rect 398062 110898 398146 111134
rect 398382 110898 433826 111134
rect 434062 110898 434146 111134
rect 434382 110898 469826 111134
rect 470062 110898 470146 111134
rect 470382 110898 505826 111134
rect 506062 110898 506146 111134
rect 506382 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 592650 111134
rect -8726 110866 592650 110898
rect -8726 106954 592650 106986
rect -8726 106718 -8694 106954
rect -8458 106718 -8374 106954
rect -8138 106718 33326 106954
rect 33562 106718 33646 106954
rect 33882 106718 69326 106954
rect 69562 106718 69646 106954
rect 69882 106718 105326 106954
rect 105562 106718 105646 106954
rect 105882 106718 213326 106954
rect 213562 106718 213646 106954
rect 213882 106718 249326 106954
rect 249562 106718 249646 106954
rect 249882 106718 285326 106954
rect 285562 106718 285646 106954
rect 285882 106718 321326 106954
rect 321562 106718 321646 106954
rect 321882 106718 357326 106954
rect 357562 106718 357646 106954
rect 357882 106718 393326 106954
rect 393562 106718 393646 106954
rect 393882 106718 429326 106954
rect 429562 106718 429646 106954
rect 429882 106718 465326 106954
rect 465562 106718 465646 106954
rect 465882 106718 501326 106954
rect 501562 106718 501646 106954
rect 501882 106718 537326 106954
rect 537562 106718 537646 106954
rect 537882 106718 573326 106954
rect 573562 106718 573646 106954
rect 573882 106718 592062 106954
rect 592298 106718 592382 106954
rect 592618 106718 592650 106954
rect -8726 106634 592650 106718
rect -8726 106398 -8694 106634
rect -8458 106398 -8374 106634
rect -8138 106398 33326 106634
rect 33562 106398 33646 106634
rect 33882 106398 69326 106634
rect 69562 106398 69646 106634
rect 69882 106398 105326 106634
rect 105562 106398 105646 106634
rect 105882 106398 213326 106634
rect 213562 106398 213646 106634
rect 213882 106398 249326 106634
rect 249562 106398 249646 106634
rect 249882 106398 285326 106634
rect 285562 106398 285646 106634
rect 285882 106398 321326 106634
rect 321562 106398 321646 106634
rect 321882 106398 357326 106634
rect 357562 106398 357646 106634
rect 357882 106398 393326 106634
rect 393562 106398 393646 106634
rect 393882 106398 429326 106634
rect 429562 106398 429646 106634
rect 429882 106398 465326 106634
rect 465562 106398 465646 106634
rect 465882 106398 501326 106634
rect 501562 106398 501646 106634
rect 501882 106398 537326 106634
rect 537562 106398 537646 106634
rect 537882 106398 573326 106634
rect 573562 106398 573646 106634
rect 573882 106398 592062 106634
rect 592298 106398 592382 106634
rect 592618 106398 592650 106634
rect -8726 106366 592650 106398
rect -8726 102454 592650 102486
rect -8726 102218 -7734 102454
rect -7498 102218 -7414 102454
rect -7178 102218 28826 102454
rect 29062 102218 29146 102454
rect 29382 102218 64826 102454
rect 65062 102218 65146 102454
rect 65382 102218 100826 102454
rect 101062 102218 101146 102454
rect 101382 102218 208826 102454
rect 209062 102218 209146 102454
rect 209382 102218 244826 102454
rect 245062 102218 245146 102454
rect 245382 102218 280826 102454
rect 281062 102218 281146 102454
rect 281382 102218 316826 102454
rect 317062 102218 317146 102454
rect 317382 102218 352826 102454
rect 353062 102218 353146 102454
rect 353382 102218 388826 102454
rect 389062 102218 389146 102454
rect 389382 102218 424826 102454
rect 425062 102218 425146 102454
rect 425382 102218 460826 102454
rect 461062 102218 461146 102454
rect 461382 102218 496826 102454
rect 497062 102218 497146 102454
rect 497382 102218 532826 102454
rect 533062 102218 533146 102454
rect 533382 102218 568826 102454
rect 569062 102218 569146 102454
rect 569382 102218 591102 102454
rect 591338 102218 591422 102454
rect 591658 102218 592650 102454
rect -8726 102134 592650 102218
rect -8726 101898 -7734 102134
rect -7498 101898 -7414 102134
rect -7178 101898 28826 102134
rect 29062 101898 29146 102134
rect 29382 101898 64826 102134
rect 65062 101898 65146 102134
rect 65382 101898 100826 102134
rect 101062 101898 101146 102134
rect 101382 101898 208826 102134
rect 209062 101898 209146 102134
rect 209382 101898 244826 102134
rect 245062 101898 245146 102134
rect 245382 101898 280826 102134
rect 281062 101898 281146 102134
rect 281382 101898 316826 102134
rect 317062 101898 317146 102134
rect 317382 101898 352826 102134
rect 353062 101898 353146 102134
rect 353382 101898 388826 102134
rect 389062 101898 389146 102134
rect 389382 101898 424826 102134
rect 425062 101898 425146 102134
rect 425382 101898 460826 102134
rect 461062 101898 461146 102134
rect 461382 101898 496826 102134
rect 497062 101898 497146 102134
rect 497382 101898 532826 102134
rect 533062 101898 533146 102134
rect 533382 101898 568826 102134
rect 569062 101898 569146 102134
rect 569382 101898 591102 102134
rect 591338 101898 591422 102134
rect 591658 101898 592650 102134
rect -8726 101866 592650 101898
rect -8726 97954 592650 97986
rect -8726 97718 -6774 97954
rect -6538 97718 -6454 97954
rect -6218 97718 24326 97954
rect 24562 97718 24646 97954
rect 24882 97718 60326 97954
rect 60562 97718 60646 97954
rect 60882 97718 96326 97954
rect 96562 97718 96646 97954
rect 96882 97718 204326 97954
rect 204562 97718 204646 97954
rect 204882 97718 240326 97954
rect 240562 97718 240646 97954
rect 240882 97718 276326 97954
rect 276562 97718 276646 97954
rect 276882 97718 312326 97954
rect 312562 97718 312646 97954
rect 312882 97718 348326 97954
rect 348562 97718 348646 97954
rect 348882 97718 384326 97954
rect 384562 97718 384646 97954
rect 384882 97718 420326 97954
rect 420562 97718 420646 97954
rect 420882 97718 456326 97954
rect 456562 97718 456646 97954
rect 456882 97718 492326 97954
rect 492562 97718 492646 97954
rect 492882 97718 528326 97954
rect 528562 97718 528646 97954
rect 528882 97718 564326 97954
rect 564562 97718 564646 97954
rect 564882 97718 590142 97954
rect 590378 97718 590462 97954
rect 590698 97718 592650 97954
rect -8726 97634 592650 97718
rect -8726 97398 -6774 97634
rect -6538 97398 -6454 97634
rect -6218 97398 24326 97634
rect 24562 97398 24646 97634
rect 24882 97398 60326 97634
rect 60562 97398 60646 97634
rect 60882 97398 96326 97634
rect 96562 97398 96646 97634
rect 96882 97398 204326 97634
rect 204562 97398 204646 97634
rect 204882 97398 240326 97634
rect 240562 97398 240646 97634
rect 240882 97398 276326 97634
rect 276562 97398 276646 97634
rect 276882 97398 312326 97634
rect 312562 97398 312646 97634
rect 312882 97398 348326 97634
rect 348562 97398 348646 97634
rect 348882 97398 384326 97634
rect 384562 97398 384646 97634
rect 384882 97398 420326 97634
rect 420562 97398 420646 97634
rect 420882 97398 456326 97634
rect 456562 97398 456646 97634
rect 456882 97398 492326 97634
rect 492562 97398 492646 97634
rect 492882 97398 528326 97634
rect 528562 97398 528646 97634
rect 528882 97398 564326 97634
rect 564562 97398 564646 97634
rect 564882 97398 590142 97634
rect 590378 97398 590462 97634
rect 590698 97398 592650 97634
rect -8726 97366 592650 97398
rect -8726 93454 592650 93486
rect -8726 93218 -5814 93454
rect -5578 93218 -5494 93454
rect -5258 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 55826 93454
rect 56062 93218 56146 93454
rect 56382 93218 91826 93454
rect 92062 93218 92146 93454
rect 92382 93218 199826 93454
rect 200062 93218 200146 93454
rect 200382 93218 235826 93454
rect 236062 93218 236146 93454
rect 236382 93218 271826 93454
rect 272062 93218 272146 93454
rect 272382 93218 307826 93454
rect 308062 93218 308146 93454
rect 308382 93218 343826 93454
rect 344062 93218 344146 93454
rect 344382 93218 379826 93454
rect 380062 93218 380146 93454
rect 380382 93218 415826 93454
rect 416062 93218 416146 93454
rect 416382 93218 451826 93454
rect 452062 93218 452146 93454
rect 452382 93218 487826 93454
rect 488062 93218 488146 93454
rect 488382 93218 523826 93454
rect 524062 93218 524146 93454
rect 524382 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 589182 93454
rect 589418 93218 589502 93454
rect 589738 93218 592650 93454
rect -8726 93134 592650 93218
rect -8726 92898 -5814 93134
rect -5578 92898 -5494 93134
rect -5258 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 55826 93134
rect 56062 92898 56146 93134
rect 56382 92898 91826 93134
rect 92062 92898 92146 93134
rect 92382 92898 199826 93134
rect 200062 92898 200146 93134
rect 200382 92898 235826 93134
rect 236062 92898 236146 93134
rect 236382 92898 271826 93134
rect 272062 92898 272146 93134
rect 272382 92898 307826 93134
rect 308062 92898 308146 93134
rect 308382 92898 343826 93134
rect 344062 92898 344146 93134
rect 344382 92898 379826 93134
rect 380062 92898 380146 93134
rect 380382 92898 415826 93134
rect 416062 92898 416146 93134
rect 416382 92898 451826 93134
rect 452062 92898 452146 93134
rect 452382 92898 487826 93134
rect 488062 92898 488146 93134
rect 488382 92898 523826 93134
rect 524062 92898 524146 93134
rect 524382 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 589182 93134
rect 589418 92898 589502 93134
rect 589738 92898 592650 93134
rect -8726 92866 592650 92898
rect -8726 88954 592650 88986
rect -8726 88718 -4854 88954
rect -4618 88718 -4534 88954
rect -4298 88718 15326 88954
rect 15562 88718 15646 88954
rect 15882 88718 51326 88954
rect 51562 88718 51646 88954
rect 51882 88718 87326 88954
rect 87562 88718 87646 88954
rect 87882 88718 195326 88954
rect 195562 88718 195646 88954
rect 195882 88718 231326 88954
rect 231562 88718 231646 88954
rect 231882 88718 267326 88954
rect 267562 88718 267646 88954
rect 267882 88718 303326 88954
rect 303562 88718 303646 88954
rect 303882 88718 339326 88954
rect 339562 88718 339646 88954
rect 339882 88718 375326 88954
rect 375562 88718 375646 88954
rect 375882 88718 411326 88954
rect 411562 88718 411646 88954
rect 411882 88718 447326 88954
rect 447562 88718 447646 88954
rect 447882 88718 483326 88954
rect 483562 88718 483646 88954
rect 483882 88718 519326 88954
rect 519562 88718 519646 88954
rect 519882 88718 555326 88954
rect 555562 88718 555646 88954
rect 555882 88718 588222 88954
rect 588458 88718 588542 88954
rect 588778 88718 592650 88954
rect -8726 88634 592650 88718
rect -8726 88398 -4854 88634
rect -4618 88398 -4534 88634
rect -4298 88398 15326 88634
rect 15562 88398 15646 88634
rect 15882 88398 51326 88634
rect 51562 88398 51646 88634
rect 51882 88398 87326 88634
rect 87562 88398 87646 88634
rect 87882 88398 195326 88634
rect 195562 88398 195646 88634
rect 195882 88398 231326 88634
rect 231562 88398 231646 88634
rect 231882 88398 267326 88634
rect 267562 88398 267646 88634
rect 267882 88398 303326 88634
rect 303562 88398 303646 88634
rect 303882 88398 339326 88634
rect 339562 88398 339646 88634
rect 339882 88398 375326 88634
rect 375562 88398 375646 88634
rect 375882 88398 411326 88634
rect 411562 88398 411646 88634
rect 411882 88398 447326 88634
rect 447562 88398 447646 88634
rect 447882 88398 483326 88634
rect 483562 88398 483646 88634
rect 483882 88398 519326 88634
rect 519562 88398 519646 88634
rect 519882 88398 555326 88634
rect 555562 88398 555646 88634
rect 555882 88398 588222 88634
rect 588458 88398 588542 88634
rect 588778 88398 592650 88634
rect -8726 88366 592650 88398
rect -8726 84454 592650 84486
rect -8726 84218 -3894 84454
rect -3658 84218 -3574 84454
rect -3338 84218 10826 84454
rect 11062 84218 11146 84454
rect 11382 84218 46826 84454
rect 47062 84218 47146 84454
rect 47382 84218 82826 84454
rect 83062 84218 83146 84454
rect 83382 84218 226826 84454
rect 227062 84218 227146 84454
rect 227382 84218 262826 84454
rect 263062 84218 263146 84454
rect 263382 84218 298826 84454
rect 299062 84218 299146 84454
rect 299382 84218 334826 84454
rect 335062 84218 335146 84454
rect 335382 84218 370826 84454
rect 371062 84218 371146 84454
rect 371382 84218 406826 84454
rect 407062 84218 407146 84454
rect 407382 84218 442826 84454
rect 443062 84218 443146 84454
rect 443382 84218 478826 84454
rect 479062 84218 479146 84454
rect 479382 84218 514826 84454
rect 515062 84218 515146 84454
rect 515382 84218 550826 84454
rect 551062 84218 551146 84454
rect 551382 84218 587262 84454
rect 587498 84218 587582 84454
rect 587818 84218 592650 84454
rect -8726 84134 592650 84218
rect -8726 83898 -3894 84134
rect -3658 83898 -3574 84134
rect -3338 83898 10826 84134
rect 11062 83898 11146 84134
rect 11382 83898 46826 84134
rect 47062 83898 47146 84134
rect 47382 83898 82826 84134
rect 83062 83898 83146 84134
rect 83382 83898 226826 84134
rect 227062 83898 227146 84134
rect 227382 83898 262826 84134
rect 263062 83898 263146 84134
rect 263382 83898 298826 84134
rect 299062 83898 299146 84134
rect 299382 83898 334826 84134
rect 335062 83898 335146 84134
rect 335382 83898 370826 84134
rect 371062 83898 371146 84134
rect 371382 83898 406826 84134
rect 407062 83898 407146 84134
rect 407382 83898 442826 84134
rect 443062 83898 443146 84134
rect 443382 83898 478826 84134
rect 479062 83898 479146 84134
rect 479382 83898 514826 84134
rect 515062 83898 515146 84134
rect 515382 83898 550826 84134
rect 551062 83898 551146 84134
rect 551382 83898 587262 84134
rect 587498 83898 587582 84134
rect 587818 83898 592650 84134
rect -8726 83866 592650 83898
rect -8726 79954 592650 79986
rect -8726 79718 -2934 79954
rect -2698 79718 -2614 79954
rect -2378 79718 6326 79954
rect 6562 79718 6646 79954
rect 6882 79718 42326 79954
rect 42562 79718 42646 79954
rect 42882 79718 78326 79954
rect 78562 79718 78646 79954
rect 78882 79718 114326 79954
rect 114562 79718 114646 79954
rect 114882 79718 222326 79954
rect 222562 79718 222646 79954
rect 222882 79718 258326 79954
rect 258562 79718 258646 79954
rect 258882 79718 294326 79954
rect 294562 79718 294646 79954
rect 294882 79718 330326 79954
rect 330562 79718 330646 79954
rect 330882 79718 366326 79954
rect 366562 79718 366646 79954
rect 366882 79718 402326 79954
rect 402562 79718 402646 79954
rect 402882 79718 438326 79954
rect 438562 79718 438646 79954
rect 438882 79718 474326 79954
rect 474562 79718 474646 79954
rect 474882 79718 510326 79954
rect 510562 79718 510646 79954
rect 510882 79718 546326 79954
rect 546562 79718 546646 79954
rect 546882 79718 582326 79954
rect 582562 79718 582646 79954
rect 582882 79718 586302 79954
rect 586538 79718 586622 79954
rect 586858 79718 592650 79954
rect -8726 79634 592650 79718
rect -8726 79398 -2934 79634
rect -2698 79398 -2614 79634
rect -2378 79398 6326 79634
rect 6562 79398 6646 79634
rect 6882 79398 42326 79634
rect 42562 79398 42646 79634
rect 42882 79398 78326 79634
rect 78562 79398 78646 79634
rect 78882 79398 114326 79634
rect 114562 79398 114646 79634
rect 114882 79398 222326 79634
rect 222562 79398 222646 79634
rect 222882 79398 258326 79634
rect 258562 79398 258646 79634
rect 258882 79398 294326 79634
rect 294562 79398 294646 79634
rect 294882 79398 330326 79634
rect 330562 79398 330646 79634
rect 330882 79398 366326 79634
rect 366562 79398 366646 79634
rect 366882 79398 402326 79634
rect 402562 79398 402646 79634
rect 402882 79398 438326 79634
rect 438562 79398 438646 79634
rect 438882 79398 474326 79634
rect 474562 79398 474646 79634
rect 474882 79398 510326 79634
rect 510562 79398 510646 79634
rect 510882 79398 546326 79634
rect 546562 79398 546646 79634
rect 546882 79398 582326 79634
rect 582562 79398 582646 79634
rect 582882 79398 586302 79634
rect 586538 79398 586622 79634
rect 586858 79398 592650 79634
rect -8726 79366 592650 79398
rect -8726 75454 592650 75486
rect -8726 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 73826 75454
rect 74062 75218 74146 75454
rect 74382 75218 109826 75454
rect 110062 75218 110146 75454
rect 110382 75218 145826 75454
rect 146062 75218 146146 75454
rect 146382 75218 181826 75454
rect 182062 75218 182146 75454
rect 182382 75218 217826 75454
rect 218062 75218 218146 75454
rect 218382 75218 253826 75454
rect 254062 75218 254146 75454
rect 254382 75218 289826 75454
rect 290062 75218 290146 75454
rect 290382 75218 325826 75454
rect 326062 75218 326146 75454
rect 326382 75218 361826 75454
rect 362062 75218 362146 75454
rect 362382 75218 397826 75454
rect 398062 75218 398146 75454
rect 398382 75218 433826 75454
rect 434062 75218 434146 75454
rect 434382 75218 469826 75454
rect 470062 75218 470146 75454
rect 470382 75218 505826 75454
rect 506062 75218 506146 75454
rect 506382 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 592650 75454
rect -8726 75134 592650 75218
rect -8726 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 73826 75134
rect 74062 74898 74146 75134
rect 74382 74898 109826 75134
rect 110062 74898 110146 75134
rect 110382 74898 145826 75134
rect 146062 74898 146146 75134
rect 146382 74898 181826 75134
rect 182062 74898 182146 75134
rect 182382 74898 217826 75134
rect 218062 74898 218146 75134
rect 218382 74898 253826 75134
rect 254062 74898 254146 75134
rect 254382 74898 289826 75134
rect 290062 74898 290146 75134
rect 290382 74898 325826 75134
rect 326062 74898 326146 75134
rect 326382 74898 361826 75134
rect 362062 74898 362146 75134
rect 362382 74898 397826 75134
rect 398062 74898 398146 75134
rect 398382 74898 433826 75134
rect 434062 74898 434146 75134
rect 434382 74898 469826 75134
rect 470062 74898 470146 75134
rect 470382 74898 505826 75134
rect 506062 74898 506146 75134
rect 506382 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 592650 75134
rect -8726 74866 592650 74898
rect -8726 70954 592650 70986
rect -8726 70718 -8694 70954
rect -8458 70718 -8374 70954
rect -8138 70718 33326 70954
rect 33562 70718 33646 70954
rect 33882 70718 69326 70954
rect 69562 70718 69646 70954
rect 69882 70718 105326 70954
rect 105562 70718 105646 70954
rect 105882 70718 141326 70954
rect 141562 70718 141646 70954
rect 141882 70718 177326 70954
rect 177562 70718 177646 70954
rect 177882 70718 213326 70954
rect 213562 70718 213646 70954
rect 213882 70718 249326 70954
rect 249562 70718 249646 70954
rect 249882 70718 285326 70954
rect 285562 70718 285646 70954
rect 285882 70718 321326 70954
rect 321562 70718 321646 70954
rect 321882 70718 357326 70954
rect 357562 70718 357646 70954
rect 357882 70718 393326 70954
rect 393562 70718 393646 70954
rect 393882 70718 429326 70954
rect 429562 70718 429646 70954
rect 429882 70718 465326 70954
rect 465562 70718 465646 70954
rect 465882 70718 501326 70954
rect 501562 70718 501646 70954
rect 501882 70718 537326 70954
rect 537562 70718 537646 70954
rect 537882 70718 573326 70954
rect 573562 70718 573646 70954
rect 573882 70718 592062 70954
rect 592298 70718 592382 70954
rect 592618 70718 592650 70954
rect -8726 70634 592650 70718
rect -8726 70398 -8694 70634
rect -8458 70398 -8374 70634
rect -8138 70398 33326 70634
rect 33562 70398 33646 70634
rect 33882 70398 69326 70634
rect 69562 70398 69646 70634
rect 69882 70398 105326 70634
rect 105562 70398 105646 70634
rect 105882 70398 141326 70634
rect 141562 70398 141646 70634
rect 141882 70398 177326 70634
rect 177562 70398 177646 70634
rect 177882 70398 213326 70634
rect 213562 70398 213646 70634
rect 213882 70398 249326 70634
rect 249562 70398 249646 70634
rect 249882 70398 285326 70634
rect 285562 70398 285646 70634
rect 285882 70398 321326 70634
rect 321562 70398 321646 70634
rect 321882 70398 357326 70634
rect 357562 70398 357646 70634
rect 357882 70398 393326 70634
rect 393562 70398 393646 70634
rect 393882 70398 429326 70634
rect 429562 70398 429646 70634
rect 429882 70398 465326 70634
rect 465562 70398 465646 70634
rect 465882 70398 501326 70634
rect 501562 70398 501646 70634
rect 501882 70398 537326 70634
rect 537562 70398 537646 70634
rect 537882 70398 573326 70634
rect 573562 70398 573646 70634
rect 573882 70398 592062 70634
rect 592298 70398 592382 70634
rect 592618 70398 592650 70634
rect -8726 70366 592650 70398
rect -8726 66454 592650 66486
rect -8726 66218 -7734 66454
rect -7498 66218 -7414 66454
rect -7178 66218 28826 66454
rect 29062 66218 29146 66454
rect 29382 66218 64826 66454
rect 65062 66218 65146 66454
rect 65382 66218 100826 66454
rect 101062 66218 101146 66454
rect 101382 66218 136826 66454
rect 137062 66218 137146 66454
rect 137382 66218 172826 66454
rect 173062 66218 173146 66454
rect 173382 66218 208826 66454
rect 209062 66218 209146 66454
rect 209382 66218 244826 66454
rect 245062 66218 245146 66454
rect 245382 66218 280826 66454
rect 281062 66218 281146 66454
rect 281382 66218 316826 66454
rect 317062 66218 317146 66454
rect 317382 66218 352826 66454
rect 353062 66218 353146 66454
rect 353382 66218 388826 66454
rect 389062 66218 389146 66454
rect 389382 66218 424826 66454
rect 425062 66218 425146 66454
rect 425382 66218 460826 66454
rect 461062 66218 461146 66454
rect 461382 66218 496826 66454
rect 497062 66218 497146 66454
rect 497382 66218 532826 66454
rect 533062 66218 533146 66454
rect 533382 66218 568826 66454
rect 569062 66218 569146 66454
rect 569382 66218 591102 66454
rect 591338 66218 591422 66454
rect 591658 66218 592650 66454
rect -8726 66134 592650 66218
rect -8726 65898 -7734 66134
rect -7498 65898 -7414 66134
rect -7178 65898 28826 66134
rect 29062 65898 29146 66134
rect 29382 65898 64826 66134
rect 65062 65898 65146 66134
rect 65382 65898 100826 66134
rect 101062 65898 101146 66134
rect 101382 65898 136826 66134
rect 137062 65898 137146 66134
rect 137382 65898 172826 66134
rect 173062 65898 173146 66134
rect 173382 65898 208826 66134
rect 209062 65898 209146 66134
rect 209382 65898 244826 66134
rect 245062 65898 245146 66134
rect 245382 65898 280826 66134
rect 281062 65898 281146 66134
rect 281382 65898 316826 66134
rect 317062 65898 317146 66134
rect 317382 65898 352826 66134
rect 353062 65898 353146 66134
rect 353382 65898 388826 66134
rect 389062 65898 389146 66134
rect 389382 65898 424826 66134
rect 425062 65898 425146 66134
rect 425382 65898 460826 66134
rect 461062 65898 461146 66134
rect 461382 65898 496826 66134
rect 497062 65898 497146 66134
rect 497382 65898 532826 66134
rect 533062 65898 533146 66134
rect 533382 65898 568826 66134
rect 569062 65898 569146 66134
rect 569382 65898 591102 66134
rect 591338 65898 591422 66134
rect 591658 65898 592650 66134
rect -8726 65866 592650 65898
rect -8726 61954 592650 61986
rect -8726 61718 -6774 61954
rect -6538 61718 -6454 61954
rect -6218 61718 24326 61954
rect 24562 61718 24646 61954
rect 24882 61718 60326 61954
rect 60562 61718 60646 61954
rect 60882 61718 96326 61954
rect 96562 61718 96646 61954
rect 96882 61718 132326 61954
rect 132562 61718 132646 61954
rect 132882 61718 168326 61954
rect 168562 61718 168646 61954
rect 168882 61718 204326 61954
rect 204562 61718 204646 61954
rect 204882 61718 240326 61954
rect 240562 61718 240646 61954
rect 240882 61718 276326 61954
rect 276562 61718 276646 61954
rect 276882 61718 312326 61954
rect 312562 61718 312646 61954
rect 312882 61718 348326 61954
rect 348562 61718 348646 61954
rect 348882 61718 384326 61954
rect 384562 61718 384646 61954
rect 384882 61718 420326 61954
rect 420562 61718 420646 61954
rect 420882 61718 456326 61954
rect 456562 61718 456646 61954
rect 456882 61718 492326 61954
rect 492562 61718 492646 61954
rect 492882 61718 528326 61954
rect 528562 61718 528646 61954
rect 528882 61718 564326 61954
rect 564562 61718 564646 61954
rect 564882 61718 590142 61954
rect 590378 61718 590462 61954
rect 590698 61718 592650 61954
rect -8726 61634 592650 61718
rect -8726 61398 -6774 61634
rect -6538 61398 -6454 61634
rect -6218 61398 24326 61634
rect 24562 61398 24646 61634
rect 24882 61398 60326 61634
rect 60562 61398 60646 61634
rect 60882 61398 96326 61634
rect 96562 61398 96646 61634
rect 96882 61398 132326 61634
rect 132562 61398 132646 61634
rect 132882 61398 168326 61634
rect 168562 61398 168646 61634
rect 168882 61398 204326 61634
rect 204562 61398 204646 61634
rect 204882 61398 240326 61634
rect 240562 61398 240646 61634
rect 240882 61398 276326 61634
rect 276562 61398 276646 61634
rect 276882 61398 312326 61634
rect 312562 61398 312646 61634
rect 312882 61398 348326 61634
rect 348562 61398 348646 61634
rect 348882 61398 384326 61634
rect 384562 61398 384646 61634
rect 384882 61398 420326 61634
rect 420562 61398 420646 61634
rect 420882 61398 456326 61634
rect 456562 61398 456646 61634
rect 456882 61398 492326 61634
rect 492562 61398 492646 61634
rect 492882 61398 528326 61634
rect 528562 61398 528646 61634
rect 528882 61398 564326 61634
rect 564562 61398 564646 61634
rect 564882 61398 590142 61634
rect 590378 61398 590462 61634
rect 590698 61398 592650 61634
rect -8726 61366 592650 61398
rect -8726 57454 592650 57486
rect -8726 57218 -5814 57454
rect -5578 57218 -5494 57454
rect -5258 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 55826 57454
rect 56062 57218 56146 57454
rect 56382 57218 91826 57454
rect 92062 57218 92146 57454
rect 92382 57218 127826 57454
rect 128062 57218 128146 57454
rect 128382 57218 163826 57454
rect 164062 57218 164146 57454
rect 164382 57218 199826 57454
rect 200062 57218 200146 57454
rect 200382 57218 235826 57454
rect 236062 57218 236146 57454
rect 236382 57218 271826 57454
rect 272062 57218 272146 57454
rect 272382 57218 307826 57454
rect 308062 57218 308146 57454
rect 308382 57218 343826 57454
rect 344062 57218 344146 57454
rect 344382 57218 379826 57454
rect 380062 57218 380146 57454
rect 380382 57218 415826 57454
rect 416062 57218 416146 57454
rect 416382 57218 451826 57454
rect 452062 57218 452146 57454
rect 452382 57218 487826 57454
rect 488062 57218 488146 57454
rect 488382 57218 523826 57454
rect 524062 57218 524146 57454
rect 524382 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 589182 57454
rect 589418 57218 589502 57454
rect 589738 57218 592650 57454
rect -8726 57134 592650 57218
rect -8726 56898 -5814 57134
rect -5578 56898 -5494 57134
rect -5258 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 55826 57134
rect 56062 56898 56146 57134
rect 56382 56898 91826 57134
rect 92062 56898 92146 57134
rect 92382 56898 127826 57134
rect 128062 56898 128146 57134
rect 128382 56898 163826 57134
rect 164062 56898 164146 57134
rect 164382 56898 199826 57134
rect 200062 56898 200146 57134
rect 200382 56898 235826 57134
rect 236062 56898 236146 57134
rect 236382 56898 271826 57134
rect 272062 56898 272146 57134
rect 272382 56898 307826 57134
rect 308062 56898 308146 57134
rect 308382 56898 343826 57134
rect 344062 56898 344146 57134
rect 344382 56898 379826 57134
rect 380062 56898 380146 57134
rect 380382 56898 415826 57134
rect 416062 56898 416146 57134
rect 416382 56898 451826 57134
rect 452062 56898 452146 57134
rect 452382 56898 487826 57134
rect 488062 56898 488146 57134
rect 488382 56898 523826 57134
rect 524062 56898 524146 57134
rect 524382 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 589182 57134
rect 589418 56898 589502 57134
rect 589738 56898 592650 57134
rect -8726 56866 592650 56898
rect -8726 52954 592650 52986
rect -8726 52718 -4854 52954
rect -4618 52718 -4534 52954
rect -4298 52718 15326 52954
rect 15562 52718 15646 52954
rect 15882 52718 51326 52954
rect 51562 52718 51646 52954
rect 51882 52718 87326 52954
rect 87562 52718 87646 52954
rect 87882 52718 123326 52954
rect 123562 52718 123646 52954
rect 123882 52718 159326 52954
rect 159562 52718 159646 52954
rect 159882 52718 195326 52954
rect 195562 52718 195646 52954
rect 195882 52718 231326 52954
rect 231562 52718 231646 52954
rect 231882 52718 267326 52954
rect 267562 52718 267646 52954
rect 267882 52718 303326 52954
rect 303562 52718 303646 52954
rect 303882 52718 339326 52954
rect 339562 52718 339646 52954
rect 339882 52718 375326 52954
rect 375562 52718 375646 52954
rect 375882 52718 411326 52954
rect 411562 52718 411646 52954
rect 411882 52718 447326 52954
rect 447562 52718 447646 52954
rect 447882 52718 483326 52954
rect 483562 52718 483646 52954
rect 483882 52718 519326 52954
rect 519562 52718 519646 52954
rect 519882 52718 555326 52954
rect 555562 52718 555646 52954
rect 555882 52718 588222 52954
rect 588458 52718 588542 52954
rect 588778 52718 592650 52954
rect -8726 52634 592650 52718
rect -8726 52398 -4854 52634
rect -4618 52398 -4534 52634
rect -4298 52398 15326 52634
rect 15562 52398 15646 52634
rect 15882 52398 51326 52634
rect 51562 52398 51646 52634
rect 51882 52398 87326 52634
rect 87562 52398 87646 52634
rect 87882 52398 123326 52634
rect 123562 52398 123646 52634
rect 123882 52398 159326 52634
rect 159562 52398 159646 52634
rect 159882 52398 195326 52634
rect 195562 52398 195646 52634
rect 195882 52398 231326 52634
rect 231562 52398 231646 52634
rect 231882 52398 267326 52634
rect 267562 52398 267646 52634
rect 267882 52398 303326 52634
rect 303562 52398 303646 52634
rect 303882 52398 339326 52634
rect 339562 52398 339646 52634
rect 339882 52398 375326 52634
rect 375562 52398 375646 52634
rect 375882 52398 411326 52634
rect 411562 52398 411646 52634
rect 411882 52398 447326 52634
rect 447562 52398 447646 52634
rect 447882 52398 483326 52634
rect 483562 52398 483646 52634
rect 483882 52398 519326 52634
rect 519562 52398 519646 52634
rect 519882 52398 555326 52634
rect 555562 52398 555646 52634
rect 555882 52398 588222 52634
rect 588458 52398 588542 52634
rect 588778 52398 592650 52634
rect -8726 52366 592650 52398
rect -8726 48454 592650 48486
rect -8726 48218 -3894 48454
rect -3658 48218 -3574 48454
rect -3338 48218 10826 48454
rect 11062 48218 11146 48454
rect 11382 48218 46826 48454
rect 47062 48218 47146 48454
rect 47382 48218 82826 48454
rect 83062 48218 83146 48454
rect 83382 48218 118826 48454
rect 119062 48218 119146 48454
rect 119382 48218 154826 48454
rect 155062 48218 155146 48454
rect 155382 48218 190826 48454
rect 191062 48218 191146 48454
rect 191382 48218 226826 48454
rect 227062 48218 227146 48454
rect 227382 48218 262826 48454
rect 263062 48218 263146 48454
rect 263382 48218 298826 48454
rect 299062 48218 299146 48454
rect 299382 48218 334826 48454
rect 335062 48218 335146 48454
rect 335382 48218 370826 48454
rect 371062 48218 371146 48454
rect 371382 48218 406826 48454
rect 407062 48218 407146 48454
rect 407382 48218 442826 48454
rect 443062 48218 443146 48454
rect 443382 48218 478826 48454
rect 479062 48218 479146 48454
rect 479382 48218 514826 48454
rect 515062 48218 515146 48454
rect 515382 48218 550826 48454
rect 551062 48218 551146 48454
rect 551382 48218 587262 48454
rect 587498 48218 587582 48454
rect 587818 48218 592650 48454
rect -8726 48134 592650 48218
rect -8726 47898 -3894 48134
rect -3658 47898 -3574 48134
rect -3338 47898 10826 48134
rect 11062 47898 11146 48134
rect 11382 47898 46826 48134
rect 47062 47898 47146 48134
rect 47382 47898 82826 48134
rect 83062 47898 83146 48134
rect 83382 47898 118826 48134
rect 119062 47898 119146 48134
rect 119382 47898 154826 48134
rect 155062 47898 155146 48134
rect 155382 47898 190826 48134
rect 191062 47898 191146 48134
rect 191382 47898 226826 48134
rect 227062 47898 227146 48134
rect 227382 47898 262826 48134
rect 263062 47898 263146 48134
rect 263382 47898 298826 48134
rect 299062 47898 299146 48134
rect 299382 47898 334826 48134
rect 335062 47898 335146 48134
rect 335382 47898 370826 48134
rect 371062 47898 371146 48134
rect 371382 47898 406826 48134
rect 407062 47898 407146 48134
rect 407382 47898 442826 48134
rect 443062 47898 443146 48134
rect 443382 47898 478826 48134
rect 479062 47898 479146 48134
rect 479382 47898 514826 48134
rect 515062 47898 515146 48134
rect 515382 47898 550826 48134
rect 551062 47898 551146 48134
rect 551382 47898 587262 48134
rect 587498 47898 587582 48134
rect 587818 47898 592650 48134
rect -8726 47866 592650 47898
rect -8726 43954 592650 43986
rect -8726 43718 -2934 43954
rect -2698 43718 -2614 43954
rect -2378 43718 6326 43954
rect 6562 43718 6646 43954
rect 6882 43718 42326 43954
rect 42562 43718 42646 43954
rect 42882 43718 78326 43954
rect 78562 43718 78646 43954
rect 78882 43718 114326 43954
rect 114562 43718 114646 43954
rect 114882 43718 150326 43954
rect 150562 43718 150646 43954
rect 150882 43718 186326 43954
rect 186562 43718 186646 43954
rect 186882 43718 222326 43954
rect 222562 43718 222646 43954
rect 222882 43718 258326 43954
rect 258562 43718 258646 43954
rect 258882 43718 294326 43954
rect 294562 43718 294646 43954
rect 294882 43718 330326 43954
rect 330562 43718 330646 43954
rect 330882 43718 366326 43954
rect 366562 43718 366646 43954
rect 366882 43718 402326 43954
rect 402562 43718 402646 43954
rect 402882 43718 438326 43954
rect 438562 43718 438646 43954
rect 438882 43718 474326 43954
rect 474562 43718 474646 43954
rect 474882 43718 510326 43954
rect 510562 43718 510646 43954
rect 510882 43718 546326 43954
rect 546562 43718 546646 43954
rect 546882 43718 582326 43954
rect 582562 43718 582646 43954
rect 582882 43718 586302 43954
rect 586538 43718 586622 43954
rect 586858 43718 592650 43954
rect -8726 43634 592650 43718
rect -8726 43398 -2934 43634
rect -2698 43398 -2614 43634
rect -2378 43398 6326 43634
rect 6562 43398 6646 43634
rect 6882 43398 42326 43634
rect 42562 43398 42646 43634
rect 42882 43398 78326 43634
rect 78562 43398 78646 43634
rect 78882 43398 114326 43634
rect 114562 43398 114646 43634
rect 114882 43398 150326 43634
rect 150562 43398 150646 43634
rect 150882 43398 186326 43634
rect 186562 43398 186646 43634
rect 186882 43398 222326 43634
rect 222562 43398 222646 43634
rect 222882 43398 258326 43634
rect 258562 43398 258646 43634
rect 258882 43398 294326 43634
rect 294562 43398 294646 43634
rect 294882 43398 330326 43634
rect 330562 43398 330646 43634
rect 330882 43398 366326 43634
rect 366562 43398 366646 43634
rect 366882 43398 402326 43634
rect 402562 43398 402646 43634
rect 402882 43398 438326 43634
rect 438562 43398 438646 43634
rect 438882 43398 474326 43634
rect 474562 43398 474646 43634
rect 474882 43398 510326 43634
rect 510562 43398 510646 43634
rect 510882 43398 546326 43634
rect 546562 43398 546646 43634
rect 546882 43398 582326 43634
rect 582562 43398 582646 43634
rect 582882 43398 586302 43634
rect 586538 43398 586622 43634
rect 586858 43398 592650 43634
rect -8726 43366 592650 43398
rect -8726 39454 592650 39486
rect -8726 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 592650 39454
rect -8726 39134 592650 39218
rect -8726 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 592650 39134
rect -8726 38866 592650 38898
rect -8726 34954 592650 34986
rect -8726 34718 -8694 34954
rect -8458 34718 -8374 34954
rect -8138 34718 33326 34954
rect 33562 34718 33646 34954
rect 33882 34718 69326 34954
rect 69562 34718 69646 34954
rect 69882 34718 105326 34954
rect 105562 34718 105646 34954
rect 105882 34718 141326 34954
rect 141562 34718 141646 34954
rect 141882 34718 177326 34954
rect 177562 34718 177646 34954
rect 177882 34718 213326 34954
rect 213562 34718 213646 34954
rect 213882 34718 249326 34954
rect 249562 34718 249646 34954
rect 249882 34718 285326 34954
rect 285562 34718 285646 34954
rect 285882 34718 321326 34954
rect 321562 34718 321646 34954
rect 321882 34718 357326 34954
rect 357562 34718 357646 34954
rect 357882 34718 393326 34954
rect 393562 34718 393646 34954
rect 393882 34718 429326 34954
rect 429562 34718 429646 34954
rect 429882 34718 465326 34954
rect 465562 34718 465646 34954
rect 465882 34718 501326 34954
rect 501562 34718 501646 34954
rect 501882 34718 537326 34954
rect 537562 34718 537646 34954
rect 537882 34718 573326 34954
rect 573562 34718 573646 34954
rect 573882 34718 592062 34954
rect 592298 34718 592382 34954
rect 592618 34718 592650 34954
rect -8726 34634 592650 34718
rect -8726 34398 -8694 34634
rect -8458 34398 -8374 34634
rect -8138 34398 33326 34634
rect 33562 34398 33646 34634
rect 33882 34398 69326 34634
rect 69562 34398 69646 34634
rect 69882 34398 105326 34634
rect 105562 34398 105646 34634
rect 105882 34398 141326 34634
rect 141562 34398 141646 34634
rect 141882 34398 177326 34634
rect 177562 34398 177646 34634
rect 177882 34398 213326 34634
rect 213562 34398 213646 34634
rect 213882 34398 249326 34634
rect 249562 34398 249646 34634
rect 249882 34398 285326 34634
rect 285562 34398 285646 34634
rect 285882 34398 321326 34634
rect 321562 34398 321646 34634
rect 321882 34398 357326 34634
rect 357562 34398 357646 34634
rect 357882 34398 393326 34634
rect 393562 34398 393646 34634
rect 393882 34398 429326 34634
rect 429562 34398 429646 34634
rect 429882 34398 465326 34634
rect 465562 34398 465646 34634
rect 465882 34398 501326 34634
rect 501562 34398 501646 34634
rect 501882 34398 537326 34634
rect 537562 34398 537646 34634
rect 537882 34398 573326 34634
rect 573562 34398 573646 34634
rect 573882 34398 592062 34634
rect 592298 34398 592382 34634
rect 592618 34398 592650 34634
rect -8726 34366 592650 34398
rect -8726 30454 592650 30486
rect -8726 30218 -7734 30454
rect -7498 30218 -7414 30454
rect -7178 30218 28826 30454
rect 29062 30218 29146 30454
rect 29382 30218 64826 30454
rect 65062 30218 65146 30454
rect 65382 30218 100826 30454
rect 101062 30218 101146 30454
rect 101382 30218 136826 30454
rect 137062 30218 137146 30454
rect 137382 30218 172826 30454
rect 173062 30218 173146 30454
rect 173382 30218 208826 30454
rect 209062 30218 209146 30454
rect 209382 30218 244826 30454
rect 245062 30218 245146 30454
rect 245382 30218 280826 30454
rect 281062 30218 281146 30454
rect 281382 30218 316826 30454
rect 317062 30218 317146 30454
rect 317382 30218 352826 30454
rect 353062 30218 353146 30454
rect 353382 30218 388826 30454
rect 389062 30218 389146 30454
rect 389382 30218 424826 30454
rect 425062 30218 425146 30454
rect 425382 30218 460826 30454
rect 461062 30218 461146 30454
rect 461382 30218 496826 30454
rect 497062 30218 497146 30454
rect 497382 30218 532826 30454
rect 533062 30218 533146 30454
rect 533382 30218 568826 30454
rect 569062 30218 569146 30454
rect 569382 30218 591102 30454
rect 591338 30218 591422 30454
rect 591658 30218 592650 30454
rect -8726 30134 592650 30218
rect -8726 29898 -7734 30134
rect -7498 29898 -7414 30134
rect -7178 29898 28826 30134
rect 29062 29898 29146 30134
rect 29382 29898 64826 30134
rect 65062 29898 65146 30134
rect 65382 29898 100826 30134
rect 101062 29898 101146 30134
rect 101382 29898 136826 30134
rect 137062 29898 137146 30134
rect 137382 29898 172826 30134
rect 173062 29898 173146 30134
rect 173382 29898 208826 30134
rect 209062 29898 209146 30134
rect 209382 29898 244826 30134
rect 245062 29898 245146 30134
rect 245382 29898 280826 30134
rect 281062 29898 281146 30134
rect 281382 29898 316826 30134
rect 317062 29898 317146 30134
rect 317382 29898 352826 30134
rect 353062 29898 353146 30134
rect 353382 29898 388826 30134
rect 389062 29898 389146 30134
rect 389382 29898 424826 30134
rect 425062 29898 425146 30134
rect 425382 29898 460826 30134
rect 461062 29898 461146 30134
rect 461382 29898 496826 30134
rect 497062 29898 497146 30134
rect 497382 29898 532826 30134
rect 533062 29898 533146 30134
rect 533382 29898 568826 30134
rect 569062 29898 569146 30134
rect 569382 29898 591102 30134
rect 591338 29898 591422 30134
rect 591658 29898 592650 30134
rect -8726 29866 592650 29898
rect -8726 25954 592650 25986
rect -8726 25718 -6774 25954
rect -6538 25718 -6454 25954
rect -6218 25718 24326 25954
rect 24562 25718 24646 25954
rect 24882 25718 60326 25954
rect 60562 25718 60646 25954
rect 60882 25718 96326 25954
rect 96562 25718 96646 25954
rect 96882 25718 132326 25954
rect 132562 25718 132646 25954
rect 132882 25718 168326 25954
rect 168562 25718 168646 25954
rect 168882 25718 204326 25954
rect 204562 25718 204646 25954
rect 204882 25718 240326 25954
rect 240562 25718 240646 25954
rect 240882 25718 276326 25954
rect 276562 25718 276646 25954
rect 276882 25718 312326 25954
rect 312562 25718 312646 25954
rect 312882 25718 348326 25954
rect 348562 25718 348646 25954
rect 348882 25718 384326 25954
rect 384562 25718 384646 25954
rect 384882 25718 420326 25954
rect 420562 25718 420646 25954
rect 420882 25718 456326 25954
rect 456562 25718 456646 25954
rect 456882 25718 492326 25954
rect 492562 25718 492646 25954
rect 492882 25718 528326 25954
rect 528562 25718 528646 25954
rect 528882 25718 564326 25954
rect 564562 25718 564646 25954
rect 564882 25718 590142 25954
rect 590378 25718 590462 25954
rect 590698 25718 592650 25954
rect -8726 25634 592650 25718
rect -8726 25398 -6774 25634
rect -6538 25398 -6454 25634
rect -6218 25398 24326 25634
rect 24562 25398 24646 25634
rect 24882 25398 60326 25634
rect 60562 25398 60646 25634
rect 60882 25398 96326 25634
rect 96562 25398 96646 25634
rect 96882 25398 132326 25634
rect 132562 25398 132646 25634
rect 132882 25398 168326 25634
rect 168562 25398 168646 25634
rect 168882 25398 204326 25634
rect 204562 25398 204646 25634
rect 204882 25398 240326 25634
rect 240562 25398 240646 25634
rect 240882 25398 276326 25634
rect 276562 25398 276646 25634
rect 276882 25398 312326 25634
rect 312562 25398 312646 25634
rect 312882 25398 348326 25634
rect 348562 25398 348646 25634
rect 348882 25398 384326 25634
rect 384562 25398 384646 25634
rect 384882 25398 420326 25634
rect 420562 25398 420646 25634
rect 420882 25398 456326 25634
rect 456562 25398 456646 25634
rect 456882 25398 492326 25634
rect 492562 25398 492646 25634
rect 492882 25398 528326 25634
rect 528562 25398 528646 25634
rect 528882 25398 564326 25634
rect 564562 25398 564646 25634
rect 564882 25398 590142 25634
rect 590378 25398 590462 25634
rect 590698 25398 592650 25634
rect -8726 25366 592650 25398
rect -8726 21454 592650 21486
rect -8726 21218 -5814 21454
rect -5578 21218 -5494 21454
rect -5258 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 589182 21454
rect 589418 21218 589502 21454
rect 589738 21218 592650 21454
rect -8726 21134 592650 21218
rect -8726 20898 -5814 21134
rect -5578 20898 -5494 21134
rect -5258 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 589182 21134
rect 589418 20898 589502 21134
rect 589738 20898 592650 21134
rect -8726 20866 592650 20898
rect -8726 16954 592650 16986
rect -8726 16718 -4854 16954
rect -4618 16718 -4534 16954
rect -4298 16718 15326 16954
rect 15562 16718 15646 16954
rect 15882 16718 51326 16954
rect 51562 16718 51646 16954
rect 51882 16718 87326 16954
rect 87562 16718 87646 16954
rect 87882 16718 123326 16954
rect 123562 16718 123646 16954
rect 123882 16718 159326 16954
rect 159562 16718 159646 16954
rect 159882 16718 195326 16954
rect 195562 16718 195646 16954
rect 195882 16718 231326 16954
rect 231562 16718 231646 16954
rect 231882 16718 267326 16954
rect 267562 16718 267646 16954
rect 267882 16718 303326 16954
rect 303562 16718 303646 16954
rect 303882 16718 339326 16954
rect 339562 16718 339646 16954
rect 339882 16718 375326 16954
rect 375562 16718 375646 16954
rect 375882 16718 411326 16954
rect 411562 16718 411646 16954
rect 411882 16718 447326 16954
rect 447562 16718 447646 16954
rect 447882 16718 483326 16954
rect 483562 16718 483646 16954
rect 483882 16718 519326 16954
rect 519562 16718 519646 16954
rect 519882 16718 555326 16954
rect 555562 16718 555646 16954
rect 555882 16718 588222 16954
rect 588458 16718 588542 16954
rect 588778 16718 592650 16954
rect -8726 16634 592650 16718
rect -8726 16398 -4854 16634
rect -4618 16398 -4534 16634
rect -4298 16398 15326 16634
rect 15562 16398 15646 16634
rect 15882 16398 51326 16634
rect 51562 16398 51646 16634
rect 51882 16398 87326 16634
rect 87562 16398 87646 16634
rect 87882 16398 123326 16634
rect 123562 16398 123646 16634
rect 123882 16398 159326 16634
rect 159562 16398 159646 16634
rect 159882 16398 195326 16634
rect 195562 16398 195646 16634
rect 195882 16398 231326 16634
rect 231562 16398 231646 16634
rect 231882 16398 267326 16634
rect 267562 16398 267646 16634
rect 267882 16398 303326 16634
rect 303562 16398 303646 16634
rect 303882 16398 339326 16634
rect 339562 16398 339646 16634
rect 339882 16398 375326 16634
rect 375562 16398 375646 16634
rect 375882 16398 411326 16634
rect 411562 16398 411646 16634
rect 411882 16398 447326 16634
rect 447562 16398 447646 16634
rect 447882 16398 483326 16634
rect 483562 16398 483646 16634
rect 483882 16398 519326 16634
rect 519562 16398 519646 16634
rect 519882 16398 555326 16634
rect 555562 16398 555646 16634
rect 555882 16398 588222 16634
rect 588458 16398 588542 16634
rect 588778 16398 592650 16634
rect -8726 16366 592650 16398
rect -8726 12454 592650 12486
rect -8726 12218 -3894 12454
rect -3658 12218 -3574 12454
rect -3338 12218 10826 12454
rect 11062 12218 11146 12454
rect 11382 12218 46826 12454
rect 47062 12218 47146 12454
rect 47382 12218 82826 12454
rect 83062 12218 83146 12454
rect 83382 12218 118826 12454
rect 119062 12218 119146 12454
rect 119382 12218 154826 12454
rect 155062 12218 155146 12454
rect 155382 12218 190826 12454
rect 191062 12218 191146 12454
rect 191382 12218 226826 12454
rect 227062 12218 227146 12454
rect 227382 12218 262826 12454
rect 263062 12218 263146 12454
rect 263382 12218 298826 12454
rect 299062 12218 299146 12454
rect 299382 12218 334826 12454
rect 335062 12218 335146 12454
rect 335382 12218 370826 12454
rect 371062 12218 371146 12454
rect 371382 12218 406826 12454
rect 407062 12218 407146 12454
rect 407382 12218 442826 12454
rect 443062 12218 443146 12454
rect 443382 12218 478826 12454
rect 479062 12218 479146 12454
rect 479382 12218 514826 12454
rect 515062 12218 515146 12454
rect 515382 12218 550826 12454
rect 551062 12218 551146 12454
rect 551382 12218 587262 12454
rect 587498 12218 587582 12454
rect 587818 12218 592650 12454
rect -8726 12134 592650 12218
rect -8726 11898 -3894 12134
rect -3658 11898 -3574 12134
rect -3338 11898 10826 12134
rect 11062 11898 11146 12134
rect 11382 11898 46826 12134
rect 47062 11898 47146 12134
rect 47382 11898 82826 12134
rect 83062 11898 83146 12134
rect 83382 11898 118826 12134
rect 119062 11898 119146 12134
rect 119382 11898 154826 12134
rect 155062 11898 155146 12134
rect 155382 11898 190826 12134
rect 191062 11898 191146 12134
rect 191382 11898 226826 12134
rect 227062 11898 227146 12134
rect 227382 11898 262826 12134
rect 263062 11898 263146 12134
rect 263382 11898 298826 12134
rect 299062 11898 299146 12134
rect 299382 11898 334826 12134
rect 335062 11898 335146 12134
rect 335382 11898 370826 12134
rect 371062 11898 371146 12134
rect 371382 11898 406826 12134
rect 407062 11898 407146 12134
rect 407382 11898 442826 12134
rect 443062 11898 443146 12134
rect 443382 11898 478826 12134
rect 479062 11898 479146 12134
rect 479382 11898 514826 12134
rect 515062 11898 515146 12134
rect 515382 11898 550826 12134
rect 551062 11898 551146 12134
rect 551382 11898 587262 12134
rect 587498 11898 587582 12134
rect 587818 11898 592650 12134
rect -8726 11866 592650 11898
rect -8726 7954 592650 7986
rect -8726 7718 -2934 7954
rect -2698 7718 -2614 7954
rect -2378 7718 6326 7954
rect 6562 7718 6646 7954
rect 6882 7718 42326 7954
rect 42562 7718 42646 7954
rect 42882 7718 78326 7954
rect 78562 7718 78646 7954
rect 78882 7718 114326 7954
rect 114562 7718 114646 7954
rect 114882 7718 150326 7954
rect 150562 7718 150646 7954
rect 150882 7718 186326 7954
rect 186562 7718 186646 7954
rect 186882 7718 222326 7954
rect 222562 7718 222646 7954
rect 222882 7718 258326 7954
rect 258562 7718 258646 7954
rect 258882 7718 294326 7954
rect 294562 7718 294646 7954
rect 294882 7718 330326 7954
rect 330562 7718 330646 7954
rect 330882 7718 366326 7954
rect 366562 7718 366646 7954
rect 366882 7718 402326 7954
rect 402562 7718 402646 7954
rect 402882 7718 438326 7954
rect 438562 7718 438646 7954
rect 438882 7718 474326 7954
rect 474562 7718 474646 7954
rect 474882 7718 510326 7954
rect 510562 7718 510646 7954
rect 510882 7718 546326 7954
rect 546562 7718 546646 7954
rect 546882 7718 582326 7954
rect 582562 7718 582646 7954
rect 582882 7718 586302 7954
rect 586538 7718 586622 7954
rect 586858 7718 592650 7954
rect -8726 7634 592650 7718
rect -8726 7398 -2934 7634
rect -2698 7398 -2614 7634
rect -2378 7398 6326 7634
rect 6562 7398 6646 7634
rect 6882 7398 42326 7634
rect 42562 7398 42646 7634
rect 42882 7398 78326 7634
rect 78562 7398 78646 7634
rect 78882 7398 114326 7634
rect 114562 7398 114646 7634
rect 114882 7398 150326 7634
rect 150562 7398 150646 7634
rect 150882 7398 186326 7634
rect 186562 7398 186646 7634
rect 186882 7398 222326 7634
rect 222562 7398 222646 7634
rect 222882 7398 258326 7634
rect 258562 7398 258646 7634
rect 258882 7398 294326 7634
rect 294562 7398 294646 7634
rect 294882 7398 330326 7634
rect 330562 7398 330646 7634
rect 330882 7398 366326 7634
rect 366562 7398 366646 7634
rect 366882 7398 402326 7634
rect 402562 7398 402646 7634
rect 402882 7398 438326 7634
rect 438562 7398 438646 7634
rect 438882 7398 474326 7634
rect 474562 7398 474646 7634
rect 474882 7398 510326 7634
rect 510562 7398 510646 7634
rect 510882 7398 546326 7634
rect 546562 7398 546646 7634
rect 546882 7398 582326 7634
rect 582562 7398 582646 7634
rect 582882 7398 586302 7634
rect 586538 7398 586622 7634
rect 586858 7398 592650 7634
rect -8726 7366 592650 7398
rect -8726 3454 592650 3486
rect -8726 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 592650 3454
rect -8726 3134 592650 3218
rect -8726 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 592650 3134
rect -8726 2866 592650 2898
rect -2006 -346 585930 -314
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect -2006 -666 585930 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect -2006 -934 585930 -902
rect -2966 -1306 586890 -1274
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 6326 -1306
rect 6562 -1542 6646 -1306
rect 6882 -1542 42326 -1306
rect 42562 -1542 42646 -1306
rect 42882 -1542 78326 -1306
rect 78562 -1542 78646 -1306
rect 78882 -1542 114326 -1306
rect 114562 -1542 114646 -1306
rect 114882 -1542 150326 -1306
rect 150562 -1542 150646 -1306
rect 150882 -1542 186326 -1306
rect 186562 -1542 186646 -1306
rect 186882 -1542 222326 -1306
rect 222562 -1542 222646 -1306
rect 222882 -1542 258326 -1306
rect 258562 -1542 258646 -1306
rect 258882 -1542 294326 -1306
rect 294562 -1542 294646 -1306
rect 294882 -1542 330326 -1306
rect 330562 -1542 330646 -1306
rect 330882 -1542 366326 -1306
rect 366562 -1542 366646 -1306
rect 366882 -1542 402326 -1306
rect 402562 -1542 402646 -1306
rect 402882 -1542 438326 -1306
rect 438562 -1542 438646 -1306
rect 438882 -1542 474326 -1306
rect 474562 -1542 474646 -1306
rect 474882 -1542 510326 -1306
rect 510562 -1542 510646 -1306
rect 510882 -1542 546326 -1306
rect 546562 -1542 546646 -1306
rect 546882 -1542 582326 -1306
rect 582562 -1542 582646 -1306
rect 582882 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect -2966 -1626 586890 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 6326 -1626
rect 6562 -1862 6646 -1626
rect 6882 -1862 42326 -1626
rect 42562 -1862 42646 -1626
rect 42882 -1862 78326 -1626
rect 78562 -1862 78646 -1626
rect 78882 -1862 114326 -1626
rect 114562 -1862 114646 -1626
rect 114882 -1862 150326 -1626
rect 150562 -1862 150646 -1626
rect 150882 -1862 186326 -1626
rect 186562 -1862 186646 -1626
rect 186882 -1862 222326 -1626
rect 222562 -1862 222646 -1626
rect 222882 -1862 258326 -1626
rect 258562 -1862 258646 -1626
rect 258882 -1862 294326 -1626
rect 294562 -1862 294646 -1626
rect 294882 -1862 330326 -1626
rect 330562 -1862 330646 -1626
rect 330882 -1862 366326 -1626
rect 366562 -1862 366646 -1626
rect 366882 -1862 402326 -1626
rect 402562 -1862 402646 -1626
rect 402882 -1862 438326 -1626
rect 438562 -1862 438646 -1626
rect 438882 -1862 474326 -1626
rect 474562 -1862 474646 -1626
rect 474882 -1862 510326 -1626
rect 510562 -1862 510646 -1626
rect 510882 -1862 546326 -1626
rect 546562 -1862 546646 -1626
rect 546882 -1862 582326 -1626
rect 582562 -1862 582646 -1626
rect 582882 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect -2966 -1894 586890 -1862
rect -3926 -2266 587850 -2234
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 10826 -2266
rect 11062 -2502 11146 -2266
rect 11382 -2502 46826 -2266
rect 47062 -2502 47146 -2266
rect 47382 -2502 82826 -2266
rect 83062 -2502 83146 -2266
rect 83382 -2502 118826 -2266
rect 119062 -2502 119146 -2266
rect 119382 -2502 154826 -2266
rect 155062 -2502 155146 -2266
rect 155382 -2502 190826 -2266
rect 191062 -2502 191146 -2266
rect 191382 -2502 226826 -2266
rect 227062 -2502 227146 -2266
rect 227382 -2502 262826 -2266
rect 263062 -2502 263146 -2266
rect 263382 -2502 298826 -2266
rect 299062 -2502 299146 -2266
rect 299382 -2502 334826 -2266
rect 335062 -2502 335146 -2266
rect 335382 -2502 370826 -2266
rect 371062 -2502 371146 -2266
rect 371382 -2502 406826 -2266
rect 407062 -2502 407146 -2266
rect 407382 -2502 442826 -2266
rect 443062 -2502 443146 -2266
rect 443382 -2502 478826 -2266
rect 479062 -2502 479146 -2266
rect 479382 -2502 514826 -2266
rect 515062 -2502 515146 -2266
rect 515382 -2502 550826 -2266
rect 551062 -2502 551146 -2266
rect 551382 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect -3926 -2586 587850 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 10826 -2586
rect 11062 -2822 11146 -2586
rect 11382 -2822 46826 -2586
rect 47062 -2822 47146 -2586
rect 47382 -2822 82826 -2586
rect 83062 -2822 83146 -2586
rect 83382 -2822 118826 -2586
rect 119062 -2822 119146 -2586
rect 119382 -2822 154826 -2586
rect 155062 -2822 155146 -2586
rect 155382 -2822 190826 -2586
rect 191062 -2822 191146 -2586
rect 191382 -2822 226826 -2586
rect 227062 -2822 227146 -2586
rect 227382 -2822 262826 -2586
rect 263062 -2822 263146 -2586
rect 263382 -2822 298826 -2586
rect 299062 -2822 299146 -2586
rect 299382 -2822 334826 -2586
rect 335062 -2822 335146 -2586
rect 335382 -2822 370826 -2586
rect 371062 -2822 371146 -2586
rect 371382 -2822 406826 -2586
rect 407062 -2822 407146 -2586
rect 407382 -2822 442826 -2586
rect 443062 -2822 443146 -2586
rect 443382 -2822 478826 -2586
rect 479062 -2822 479146 -2586
rect 479382 -2822 514826 -2586
rect 515062 -2822 515146 -2586
rect 515382 -2822 550826 -2586
rect 551062 -2822 551146 -2586
rect 551382 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect -3926 -2854 587850 -2822
rect -4886 -3226 588810 -3194
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 15326 -3226
rect 15562 -3462 15646 -3226
rect 15882 -3462 51326 -3226
rect 51562 -3462 51646 -3226
rect 51882 -3462 87326 -3226
rect 87562 -3462 87646 -3226
rect 87882 -3462 123326 -3226
rect 123562 -3462 123646 -3226
rect 123882 -3462 159326 -3226
rect 159562 -3462 159646 -3226
rect 159882 -3462 195326 -3226
rect 195562 -3462 195646 -3226
rect 195882 -3462 231326 -3226
rect 231562 -3462 231646 -3226
rect 231882 -3462 267326 -3226
rect 267562 -3462 267646 -3226
rect 267882 -3462 303326 -3226
rect 303562 -3462 303646 -3226
rect 303882 -3462 339326 -3226
rect 339562 -3462 339646 -3226
rect 339882 -3462 375326 -3226
rect 375562 -3462 375646 -3226
rect 375882 -3462 411326 -3226
rect 411562 -3462 411646 -3226
rect 411882 -3462 447326 -3226
rect 447562 -3462 447646 -3226
rect 447882 -3462 483326 -3226
rect 483562 -3462 483646 -3226
rect 483882 -3462 519326 -3226
rect 519562 -3462 519646 -3226
rect 519882 -3462 555326 -3226
rect 555562 -3462 555646 -3226
rect 555882 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect -4886 -3546 588810 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 15326 -3546
rect 15562 -3782 15646 -3546
rect 15882 -3782 51326 -3546
rect 51562 -3782 51646 -3546
rect 51882 -3782 87326 -3546
rect 87562 -3782 87646 -3546
rect 87882 -3782 123326 -3546
rect 123562 -3782 123646 -3546
rect 123882 -3782 159326 -3546
rect 159562 -3782 159646 -3546
rect 159882 -3782 195326 -3546
rect 195562 -3782 195646 -3546
rect 195882 -3782 231326 -3546
rect 231562 -3782 231646 -3546
rect 231882 -3782 267326 -3546
rect 267562 -3782 267646 -3546
rect 267882 -3782 303326 -3546
rect 303562 -3782 303646 -3546
rect 303882 -3782 339326 -3546
rect 339562 -3782 339646 -3546
rect 339882 -3782 375326 -3546
rect 375562 -3782 375646 -3546
rect 375882 -3782 411326 -3546
rect 411562 -3782 411646 -3546
rect 411882 -3782 447326 -3546
rect 447562 -3782 447646 -3546
rect 447882 -3782 483326 -3546
rect 483562 -3782 483646 -3546
rect 483882 -3782 519326 -3546
rect 519562 -3782 519646 -3546
rect 519882 -3782 555326 -3546
rect 555562 -3782 555646 -3546
rect 555882 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect -4886 -3814 588810 -3782
rect -5846 -4186 589770 -4154
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 19826 -4186
rect 20062 -4422 20146 -4186
rect 20382 -4422 55826 -4186
rect 56062 -4422 56146 -4186
rect 56382 -4422 91826 -4186
rect 92062 -4422 92146 -4186
rect 92382 -4422 127826 -4186
rect 128062 -4422 128146 -4186
rect 128382 -4422 163826 -4186
rect 164062 -4422 164146 -4186
rect 164382 -4422 199826 -4186
rect 200062 -4422 200146 -4186
rect 200382 -4422 235826 -4186
rect 236062 -4422 236146 -4186
rect 236382 -4422 271826 -4186
rect 272062 -4422 272146 -4186
rect 272382 -4422 307826 -4186
rect 308062 -4422 308146 -4186
rect 308382 -4422 343826 -4186
rect 344062 -4422 344146 -4186
rect 344382 -4422 379826 -4186
rect 380062 -4422 380146 -4186
rect 380382 -4422 415826 -4186
rect 416062 -4422 416146 -4186
rect 416382 -4422 451826 -4186
rect 452062 -4422 452146 -4186
rect 452382 -4422 487826 -4186
rect 488062 -4422 488146 -4186
rect 488382 -4422 523826 -4186
rect 524062 -4422 524146 -4186
rect 524382 -4422 559826 -4186
rect 560062 -4422 560146 -4186
rect 560382 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect -5846 -4506 589770 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 19826 -4506
rect 20062 -4742 20146 -4506
rect 20382 -4742 55826 -4506
rect 56062 -4742 56146 -4506
rect 56382 -4742 91826 -4506
rect 92062 -4742 92146 -4506
rect 92382 -4742 127826 -4506
rect 128062 -4742 128146 -4506
rect 128382 -4742 163826 -4506
rect 164062 -4742 164146 -4506
rect 164382 -4742 199826 -4506
rect 200062 -4742 200146 -4506
rect 200382 -4742 235826 -4506
rect 236062 -4742 236146 -4506
rect 236382 -4742 271826 -4506
rect 272062 -4742 272146 -4506
rect 272382 -4742 307826 -4506
rect 308062 -4742 308146 -4506
rect 308382 -4742 343826 -4506
rect 344062 -4742 344146 -4506
rect 344382 -4742 379826 -4506
rect 380062 -4742 380146 -4506
rect 380382 -4742 415826 -4506
rect 416062 -4742 416146 -4506
rect 416382 -4742 451826 -4506
rect 452062 -4742 452146 -4506
rect 452382 -4742 487826 -4506
rect 488062 -4742 488146 -4506
rect 488382 -4742 523826 -4506
rect 524062 -4742 524146 -4506
rect 524382 -4742 559826 -4506
rect 560062 -4742 560146 -4506
rect 560382 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect -5846 -4774 589770 -4742
rect -6806 -5146 590730 -5114
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 24326 -5146
rect 24562 -5382 24646 -5146
rect 24882 -5382 60326 -5146
rect 60562 -5382 60646 -5146
rect 60882 -5382 96326 -5146
rect 96562 -5382 96646 -5146
rect 96882 -5382 132326 -5146
rect 132562 -5382 132646 -5146
rect 132882 -5382 168326 -5146
rect 168562 -5382 168646 -5146
rect 168882 -5382 204326 -5146
rect 204562 -5382 204646 -5146
rect 204882 -5382 240326 -5146
rect 240562 -5382 240646 -5146
rect 240882 -5382 276326 -5146
rect 276562 -5382 276646 -5146
rect 276882 -5382 312326 -5146
rect 312562 -5382 312646 -5146
rect 312882 -5382 348326 -5146
rect 348562 -5382 348646 -5146
rect 348882 -5382 384326 -5146
rect 384562 -5382 384646 -5146
rect 384882 -5382 420326 -5146
rect 420562 -5382 420646 -5146
rect 420882 -5382 456326 -5146
rect 456562 -5382 456646 -5146
rect 456882 -5382 492326 -5146
rect 492562 -5382 492646 -5146
rect 492882 -5382 528326 -5146
rect 528562 -5382 528646 -5146
rect 528882 -5382 564326 -5146
rect 564562 -5382 564646 -5146
rect 564882 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect -6806 -5466 590730 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 24326 -5466
rect 24562 -5702 24646 -5466
rect 24882 -5702 60326 -5466
rect 60562 -5702 60646 -5466
rect 60882 -5702 96326 -5466
rect 96562 -5702 96646 -5466
rect 96882 -5702 132326 -5466
rect 132562 -5702 132646 -5466
rect 132882 -5702 168326 -5466
rect 168562 -5702 168646 -5466
rect 168882 -5702 204326 -5466
rect 204562 -5702 204646 -5466
rect 204882 -5702 240326 -5466
rect 240562 -5702 240646 -5466
rect 240882 -5702 276326 -5466
rect 276562 -5702 276646 -5466
rect 276882 -5702 312326 -5466
rect 312562 -5702 312646 -5466
rect 312882 -5702 348326 -5466
rect 348562 -5702 348646 -5466
rect 348882 -5702 384326 -5466
rect 384562 -5702 384646 -5466
rect 384882 -5702 420326 -5466
rect 420562 -5702 420646 -5466
rect 420882 -5702 456326 -5466
rect 456562 -5702 456646 -5466
rect 456882 -5702 492326 -5466
rect 492562 -5702 492646 -5466
rect 492882 -5702 528326 -5466
rect 528562 -5702 528646 -5466
rect 528882 -5702 564326 -5466
rect 564562 -5702 564646 -5466
rect 564882 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect -6806 -5734 590730 -5702
rect -7766 -6106 591690 -6074
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 28826 -6106
rect 29062 -6342 29146 -6106
rect 29382 -6342 64826 -6106
rect 65062 -6342 65146 -6106
rect 65382 -6342 100826 -6106
rect 101062 -6342 101146 -6106
rect 101382 -6342 136826 -6106
rect 137062 -6342 137146 -6106
rect 137382 -6342 172826 -6106
rect 173062 -6342 173146 -6106
rect 173382 -6342 208826 -6106
rect 209062 -6342 209146 -6106
rect 209382 -6342 244826 -6106
rect 245062 -6342 245146 -6106
rect 245382 -6342 280826 -6106
rect 281062 -6342 281146 -6106
rect 281382 -6342 316826 -6106
rect 317062 -6342 317146 -6106
rect 317382 -6342 352826 -6106
rect 353062 -6342 353146 -6106
rect 353382 -6342 388826 -6106
rect 389062 -6342 389146 -6106
rect 389382 -6342 424826 -6106
rect 425062 -6342 425146 -6106
rect 425382 -6342 460826 -6106
rect 461062 -6342 461146 -6106
rect 461382 -6342 496826 -6106
rect 497062 -6342 497146 -6106
rect 497382 -6342 532826 -6106
rect 533062 -6342 533146 -6106
rect 533382 -6342 568826 -6106
rect 569062 -6342 569146 -6106
rect 569382 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect -7766 -6426 591690 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 28826 -6426
rect 29062 -6662 29146 -6426
rect 29382 -6662 64826 -6426
rect 65062 -6662 65146 -6426
rect 65382 -6662 100826 -6426
rect 101062 -6662 101146 -6426
rect 101382 -6662 136826 -6426
rect 137062 -6662 137146 -6426
rect 137382 -6662 172826 -6426
rect 173062 -6662 173146 -6426
rect 173382 -6662 208826 -6426
rect 209062 -6662 209146 -6426
rect 209382 -6662 244826 -6426
rect 245062 -6662 245146 -6426
rect 245382 -6662 280826 -6426
rect 281062 -6662 281146 -6426
rect 281382 -6662 316826 -6426
rect 317062 -6662 317146 -6426
rect 317382 -6662 352826 -6426
rect 353062 -6662 353146 -6426
rect 353382 -6662 388826 -6426
rect 389062 -6662 389146 -6426
rect 389382 -6662 424826 -6426
rect 425062 -6662 425146 -6426
rect 425382 -6662 460826 -6426
rect 461062 -6662 461146 -6426
rect 461382 -6662 496826 -6426
rect 497062 -6662 497146 -6426
rect 497382 -6662 532826 -6426
rect 533062 -6662 533146 -6426
rect 533382 -6662 568826 -6426
rect 569062 -6662 569146 -6426
rect 569382 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect -7766 -6694 591690 -6662
rect -8726 -7066 592650 -7034
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 33326 -7066
rect 33562 -7302 33646 -7066
rect 33882 -7302 69326 -7066
rect 69562 -7302 69646 -7066
rect 69882 -7302 105326 -7066
rect 105562 -7302 105646 -7066
rect 105882 -7302 141326 -7066
rect 141562 -7302 141646 -7066
rect 141882 -7302 177326 -7066
rect 177562 -7302 177646 -7066
rect 177882 -7302 213326 -7066
rect 213562 -7302 213646 -7066
rect 213882 -7302 249326 -7066
rect 249562 -7302 249646 -7066
rect 249882 -7302 285326 -7066
rect 285562 -7302 285646 -7066
rect 285882 -7302 321326 -7066
rect 321562 -7302 321646 -7066
rect 321882 -7302 357326 -7066
rect 357562 -7302 357646 -7066
rect 357882 -7302 393326 -7066
rect 393562 -7302 393646 -7066
rect 393882 -7302 429326 -7066
rect 429562 -7302 429646 -7066
rect 429882 -7302 465326 -7066
rect 465562 -7302 465646 -7066
rect 465882 -7302 501326 -7066
rect 501562 -7302 501646 -7066
rect 501882 -7302 537326 -7066
rect 537562 -7302 537646 -7066
rect 537882 -7302 573326 -7066
rect 573562 -7302 573646 -7066
rect 573882 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect -8726 -7386 592650 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 33326 -7386
rect 33562 -7622 33646 -7386
rect 33882 -7622 69326 -7386
rect 69562 -7622 69646 -7386
rect 69882 -7622 105326 -7386
rect 105562 -7622 105646 -7386
rect 105882 -7622 141326 -7386
rect 141562 -7622 141646 -7386
rect 141882 -7622 177326 -7386
rect 177562 -7622 177646 -7386
rect 177882 -7622 213326 -7386
rect 213562 -7622 213646 -7386
rect 213882 -7622 249326 -7386
rect 249562 -7622 249646 -7386
rect 249882 -7622 285326 -7386
rect 285562 -7622 285646 -7386
rect 285882 -7622 321326 -7386
rect 321562 -7622 321646 -7386
rect 321882 -7622 357326 -7386
rect 357562 -7622 357646 -7386
rect 357882 -7622 393326 -7386
rect 393562 -7622 393646 -7386
rect 393882 -7622 429326 -7386
rect 429562 -7622 429646 -7386
rect 429882 -7622 465326 -7386
rect 465562 -7622 465646 -7386
rect 465882 -7622 501326 -7386
rect 501562 -7622 501646 -7386
rect 501882 -7622 537326 -7386
rect 537562 -7622 537646 -7386
rect 537882 -7622 573326 -7386
rect 573562 -7622 573646 -7386
rect 573882 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect -8726 -7654 592650 -7622
use pixel_macro  pixel_macro0
timestamp 0
transform 1 0 120000 0 1 200000
box 1066 0 68854 60000
use rlbp_macro  rlbp_macro0
timestamp 0
transform 1 0 120000 0 1 80000
box 1066 0 68854 60000
<< labels >>
flabel metal3 s 583520 285276 584960 285516 0 FreeSans 960 0 0 0 analog_io[0]
port 0 nsew signal bidirectional
flabel metal2 s 446098 703520 446210 704960 0 FreeSans 448 90 0 0 analog_io[10]
port 1 nsew signal bidirectional
flabel metal2 s 381146 703520 381258 704960 0 FreeSans 448 90 0 0 analog_io[11]
port 2 nsew signal bidirectional
flabel metal2 s 316286 703520 316398 704960 0 FreeSans 448 90 0 0 analog_io[12]
port 3 nsew signal bidirectional
flabel metal2 s 251426 703520 251538 704960 0 FreeSans 448 90 0 0 analog_io[13]
port 4 nsew signal bidirectional
flabel metal2 s 186474 703520 186586 704960 0 FreeSans 448 90 0 0 analog_io[14]
port 5 nsew signal bidirectional
flabel metal2 s 121614 703520 121726 704960 0 FreeSans 448 90 0 0 analog_io[15]
port 6 nsew signal bidirectional
flabel metal2 s 56754 703520 56866 704960 0 FreeSans 448 90 0 0 analog_io[16]
port 7 nsew signal bidirectional
flabel metal3 s -960 697220 480 697460 0 FreeSans 960 0 0 0 analog_io[17]
port 8 nsew signal bidirectional
flabel metal3 s -960 644996 480 645236 0 FreeSans 960 0 0 0 analog_io[18]
port 9 nsew signal bidirectional
flabel metal3 s -960 592908 480 593148 0 FreeSans 960 0 0 0 analog_io[19]
port 10 nsew signal bidirectional
flabel metal3 s 583520 338452 584960 338692 0 FreeSans 960 0 0 0 analog_io[1]
port 11 nsew signal bidirectional
flabel metal3 s -960 540684 480 540924 0 FreeSans 960 0 0 0 analog_io[20]
port 12 nsew signal bidirectional
flabel metal3 s -960 488596 480 488836 0 FreeSans 960 0 0 0 analog_io[21]
port 13 nsew signal bidirectional
flabel metal3 s -960 436508 480 436748 0 FreeSans 960 0 0 0 analog_io[22]
port 14 nsew signal bidirectional
flabel metal3 s -960 384284 480 384524 0 FreeSans 960 0 0 0 analog_io[23]
port 15 nsew signal bidirectional
flabel metal3 s -960 332196 480 332436 0 FreeSans 960 0 0 0 analog_io[24]
port 16 nsew signal bidirectional
flabel metal3 s -960 279972 480 280212 0 FreeSans 960 0 0 0 analog_io[25]
port 17 nsew signal bidirectional
flabel metal3 s -960 227884 480 228124 0 FreeSans 960 0 0 0 analog_io[26]
port 18 nsew signal bidirectional
flabel metal3 s -960 175796 480 176036 0 FreeSans 960 0 0 0 analog_io[27]
port 19 nsew signal bidirectional
flabel metal3 s -960 123572 480 123812 0 FreeSans 960 0 0 0 analog_io[28]
port 20 nsew signal bidirectional
flabel metal3 s 583520 391628 584960 391868 0 FreeSans 960 0 0 0 analog_io[2]
port 21 nsew signal bidirectional
flabel metal3 s 583520 444668 584960 444908 0 FreeSans 960 0 0 0 analog_io[3]
port 22 nsew signal bidirectional
flabel metal3 s 583520 497844 584960 498084 0 FreeSans 960 0 0 0 analog_io[4]
port 23 nsew signal bidirectional
flabel metal3 s 583520 551020 584960 551260 0 FreeSans 960 0 0 0 analog_io[5]
port 24 nsew signal bidirectional
flabel metal3 s 583520 604060 584960 604300 0 FreeSans 960 0 0 0 analog_io[6]
port 25 nsew signal bidirectional
flabel metal3 s 583520 657236 584960 657476 0 FreeSans 960 0 0 0 analog_io[7]
port 26 nsew signal bidirectional
flabel metal2 s 575818 703520 575930 704960 0 FreeSans 448 90 0 0 analog_io[8]
port 27 nsew signal bidirectional
flabel metal2 s 510958 703520 511070 704960 0 FreeSans 448 90 0 0 analog_io[9]
port 28 nsew signal bidirectional
flabel metal3 s 583520 6476 584960 6716 0 FreeSans 960 0 0 0 io_in[0]
port 29 nsew signal input
flabel metal3 s 583520 457996 584960 458236 0 FreeSans 960 0 0 0 io_in[10]
port 30 nsew signal input
flabel metal3 s 583520 511172 584960 511412 0 FreeSans 960 0 0 0 io_in[11]
port 31 nsew signal input
flabel metal3 s 583520 564212 584960 564452 0 FreeSans 960 0 0 0 io_in[12]
port 32 nsew signal input
flabel metal3 s 583520 617388 584960 617628 0 FreeSans 960 0 0 0 io_in[13]
port 33 nsew signal input
flabel metal3 s 583520 670564 584960 670804 0 FreeSans 960 0 0 0 io_in[14]
port 34 nsew signal input
flabel metal2 s 559626 703520 559738 704960 0 FreeSans 448 90 0 0 io_in[15]
port 35 nsew signal input
flabel metal2 s 494766 703520 494878 704960 0 FreeSans 448 90 0 0 io_in[16]
port 36 nsew signal input
flabel metal2 s 429814 703520 429926 704960 0 FreeSans 448 90 0 0 io_in[17]
port 37 nsew signal input
flabel metal2 s 364954 703520 365066 704960 0 FreeSans 448 90 0 0 io_in[18]
port 38 nsew signal input
flabel metal2 s 300094 703520 300206 704960 0 FreeSans 448 90 0 0 io_in[19]
port 39 nsew signal input
flabel metal3 s 583520 46188 584960 46428 0 FreeSans 960 0 0 0 io_in[1]
port 40 nsew signal input
flabel metal2 s 235142 703520 235254 704960 0 FreeSans 448 90 0 0 io_in[20]
port 41 nsew signal input
flabel metal2 s 170282 703520 170394 704960 0 FreeSans 448 90 0 0 io_in[21]
port 42 nsew signal input
flabel metal2 s 105422 703520 105534 704960 0 FreeSans 448 90 0 0 io_in[22]
port 43 nsew signal input
flabel metal2 s 40470 703520 40582 704960 0 FreeSans 448 90 0 0 io_in[23]
port 44 nsew signal input
flabel metal3 s -960 684164 480 684404 0 FreeSans 960 0 0 0 io_in[24]
port 45 nsew signal input
flabel metal3 s -960 631940 480 632180 0 FreeSans 960 0 0 0 io_in[25]
port 46 nsew signal input
flabel metal3 s -960 579852 480 580092 0 FreeSans 960 0 0 0 io_in[26]
port 47 nsew signal input
flabel metal3 s -960 527764 480 528004 0 FreeSans 960 0 0 0 io_in[27]
port 48 nsew signal input
flabel metal3 s -960 475540 480 475780 0 FreeSans 960 0 0 0 io_in[28]
port 49 nsew signal input
flabel metal3 s -960 423452 480 423692 0 FreeSans 960 0 0 0 io_in[29]
port 50 nsew signal input
flabel metal3 s 583520 86036 584960 86276 0 FreeSans 960 0 0 0 io_in[2]
port 51 nsew signal input
flabel metal3 s -960 371228 480 371468 0 FreeSans 960 0 0 0 io_in[30]
port 52 nsew signal input
flabel metal3 s -960 319140 480 319380 0 FreeSans 960 0 0 0 io_in[31]
port 53 nsew signal input
flabel metal3 s -960 267052 480 267292 0 FreeSans 960 0 0 0 io_in[32]
port 54 nsew signal input
flabel metal3 s -960 214828 480 215068 0 FreeSans 960 0 0 0 io_in[33]
port 55 nsew signal input
flabel metal3 s -960 162740 480 162980 0 FreeSans 960 0 0 0 io_in[34]
port 56 nsew signal input
flabel metal3 s -960 110516 480 110756 0 FreeSans 960 0 0 0 io_in[35]
port 57 nsew signal input
flabel metal3 s -960 71484 480 71724 0 FreeSans 960 0 0 0 io_in[36]
port 58 nsew signal input
flabel metal3 s -960 32316 480 32556 0 FreeSans 960 0 0 0 io_in[37]
port 59 nsew signal input
flabel metal3 s 583520 125884 584960 126124 0 FreeSans 960 0 0 0 io_in[3]
port 60 nsew signal input
flabel metal3 s 583520 165732 584960 165972 0 FreeSans 960 0 0 0 io_in[4]
port 61 nsew signal input
flabel metal3 s 583520 205580 584960 205820 0 FreeSans 960 0 0 0 io_in[5]
port 62 nsew signal input
flabel metal3 s 583520 245428 584960 245668 0 FreeSans 960 0 0 0 io_in[6]
port 63 nsew signal input
flabel metal3 s 583520 298604 584960 298844 0 FreeSans 960 0 0 0 io_in[7]
port 64 nsew signal input
flabel metal3 s 583520 351780 584960 352020 0 FreeSans 960 0 0 0 io_in[8]
port 65 nsew signal input
flabel metal3 s 583520 404820 584960 405060 0 FreeSans 960 0 0 0 io_in[9]
port 66 nsew signal input
flabel metal3 s 583520 32996 584960 33236 0 FreeSans 960 0 0 0 io_oeb[0]
port 67 nsew signal tristate
flabel metal3 s 583520 484516 584960 484756 0 FreeSans 960 0 0 0 io_oeb[10]
port 68 nsew signal tristate
flabel metal3 s 583520 537692 584960 537932 0 FreeSans 960 0 0 0 io_oeb[11]
port 69 nsew signal tristate
flabel metal3 s 583520 590868 584960 591108 0 FreeSans 960 0 0 0 io_oeb[12]
port 70 nsew signal tristate
flabel metal3 s 583520 643908 584960 644148 0 FreeSans 960 0 0 0 io_oeb[13]
port 71 nsew signal tristate
flabel metal3 s 583520 697084 584960 697324 0 FreeSans 960 0 0 0 io_oeb[14]
port 72 nsew signal tristate
flabel metal2 s 527150 703520 527262 704960 0 FreeSans 448 90 0 0 io_oeb[15]
port 73 nsew signal tristate
flabel metal2 s 462290 703520 462402 704960 0 FreeSans 448 90 0 0 io_oeb[16]
port 74 nsew signal tristate
flabel metal2 s 397430 703520 397542 704960 0 FreeSans 448 90 0 0 io_oeb[17]
port 75 nsew signal tristate
flabel metal2 s 332478 703520 332590 704960 0 FreeSans 448 90 0 0 io_oeb[18]
port 76 nsew signal tristate
flabel metal2 s 267618 703520 267730 704960 0 FreeSans 448 90 0 0 io_oeb[19]
port 77 nsew signal tristate
flabel metal3 s 583520 72844 584960 73084 0 FreeSans 960 0 0 0 io_oeb[1]
port 78 nsew signal tristate
flabel metal2 s 202758 703520 202870 704960 0 FreeSans 448 90 0 0 io_oeb[20]
port 79 nsew signal tristate
flabel metal2 s 137806 703520 137918 704960 0 FreeSans 448 90 0 0 io_oeb[21]
port 80 nsew signal tristate
flabel metal2 s 72946 703520 73058 704960 0 FreeSans 448 90 0 0 io_oeb[22]
port 81 nsew signal tristate
flabel metal2 s 8086 703520 8198 704960 0 FreeSans 448 90 0 0 io_oeb[23]
port 82 nsew signal tristate
flabel metal3 s -960 658052 480 658292 0 FreeSans 960 0 0 0 io_oeb[24]
port 83 nsew signal tristate
flabel metal3 s -960 605964 480 606204 0 FreeSans 960 0 0 0 io_oeb[25]
port 84 nsew signal tristate
flabel metal3 s -960 553740 480 553980 0 FreeSans 960 0 0 0 io_oeb[26]
port 85 nsew signal tristate
flabel metal3 s -960 501652 480 501892 0 FreeSans 960 0 0 0 io_oeb[27]
port 86 nsew signal tristate
flabel metal3 s -960 449428 480 449668 0 FreeSans 960 0 0 0 io_oeb[28]
port 87 nsew signal tristate
flabel metal3 s -960 397340 480 397580 0 FreeSans 960 0 0 0 io_oeb[29]
port 88 nsew signal tristate
flabel metal3 s 583520 112692 584960 112932 0 FreeSans 960 0 0 0 io_oeb[2]
port 89 nsew signal tristate
flabel metal3 s -960 345252 480 345492 0 FreeSans 960 0 0 0 io_oeb[30]
port 90 nsew signal tristate
flabel metal3 s -960 293028 480 293268 0 FreeSans 960 0 0 0 io_oeb[31]
port 91 nsew signal tristate
flabel metal3 s -960 240940 480 241180 0 FreeSans 960 0 0 0 io_oeb[32]
port 92 nsew signal tristate
flabel metal3 s -960 188716 480 188956 0 FreeSans 960 0 0 0 io_oeb[33]
port 93 nsew signal tristate
flabel metal3 s -960 136628 480 136868 0 FreeSans 960 0 0 0 io_oeb[34]
port 94 nsew signal tristate
flabel metal3 s -960 84540 480 84780 0 FreeSans 960 0 0 0 io_oeb[35]
port 95 nsew signal tristate
flabel metal3 s -960 45372 480 45612 0 FreeSans 960 0 0 0 io_oeb[36]
port 96 nsew signal tristate
flabel metal3 s -960 6340 480 6580 0 FreeSans 960 0 0 0 io_oeb[37]
port 97 nsew signal tristate
flabel metal3 s 583520 152540 584960 152780 0 FreeSans 960 0 0 0 io_oeb[3]
port 98 nsew signal tristate
flabel metal3 s 583520 192388 584960 192628 0 FreeSans 960 0 0 0 io_oeb[4]
port 99 nsew signal tristate
flabel metal3 s 583520 232236 584960 232476 0 FreeSans 960 0 0 0 io_oeb[5]
port 100 nsew signal tristate
flabel metal3 s 583520 272084 584960 272324 0 FreeSans 960 0 0 0 io_oeb[6]
port 101 nsew signal tristate
flabel metal3 s 583520 325124 584960 325364 0 FreeSans 960 0 0 0 io_oeb[7]
port 102 nsew signal tristate
flabel metal3 s 583520 378300 584960 378540 0 FreeSans 960 0 0 0 io_oeb[8]
port 103 nsew signal tristate
flabel metal3 s 583520 431476 584960 431716 0 FreeSans 960 0 0 0 io_oeb[9]
port 104 nsew signal tristate
flabel metal3 s 583520 19668 584960 19908 0 FreeSans 960 0 0 0 io_out[0]
port 105 nsew signal tristate
flabel metal3 s 583520 471324 584960 471564 0 FreeSans 960 0 0 0 io_out[10]
port 106 nsew signal tristate
flabel metal3 s 583520 524364 584960 524604 0 FreeSans 960 0 0 0 io_out[11]
port 107 nsew signal tristate
flabel metal3 s 583520 577540 584960 577780 0 FreeSans 960 0 0 0 io_out[12]
port 108 nsew signal tristate
flabel metal3 s 583520 630716 584960 630956 0 FreeSans 960 0 0 0 io_out[13]
port 109 nsew signal tristate
flabel metal3 s 583520 683756 584960 683996 0 FreeSans 960 0 0 0 io_out[14]
port 110 nsew signal tristate
flabel metal2 s 543434 703520 543546 704960 0 FreeSans 448 90 0 0 io_out[15]
port 111 nsew signal tristate
flabel metal2 s 478482 703520 478594 704960 0 FreeSans 448 90 0 0 io_out[16]
port 112 nsew signal tristate
flabel metal2 s 413622 703520 413734 704960 0 FreeSans 448 90 0 0 io_out[17]
port 113 nsew signal tristate
flabel metal2 s 348762 703520 348874 704960 0 FreeSans 448 90 0 0 io_out[18]
port 114 nsew signal tristate
flabel metal2 s 283810 703520 283922 704960 0 FreeSans 448 90 0 0 io_out[19]
port 115 nsew signal tristate
flabel metal3 s 583520 59516 584960 59756 0 FreeSans 960 0 0 0 io_out[1]
port 116 nsew signal tristate
flabel metal2 s 218950 703520 219062 704960 0 FreeSans 448 90 0 0 io_out[20]
port 117 nsew signal tristate
flabel metal2 s 154090 703520 154202 704960 0 FreeSans 448 90 0 0 io_out[21]
port 118 nsew signal tristate
flabel metal2 s 89138 703520 89250 704960 0 FreeSans 448 90 0 0 io_out[22]
port 119 nsew signal tristate
flabel metal2 s 24278 703520 24390 704960 0 FreeSans 448 90 0 0 io_out[23]
port 120 nsew signal tristate
flabel metal3 s -960 671108 480 671348 0 FreeSans 960 0 0 0 io_out[24]
port 121 nsew signal tristate
flabel metal3 s -960 619020 480 619260 0 FreeSans 960 0 0 0 io_out[25]
port 122 nsew signal tristate
flabel metal3 s -960 566796 480 567036 0 FreeSans 960 0 0 0 io_out[26]
port 123 nsew signal tristate
flabel metal3 s -960 514708 480 514948 0 FreeSans 960 0 0 0 io_out[27]
port 124 nsew signal tristate
flabel metal3 s -960 462484 480 462724 0 FreeSans 960 0 0 0 io_out[28]
port 125 nsew signal tristate
flabel metal3 s -960 410396 480 410636 0 FreeSans 960 0 0 0 io_out[29]
port 126 nsew signal tristate
flabel metal3 s 583520 99364 584960 99604 0 FreeSans 960 0 0 0 io_out[2]
port 127 nsew signal tristate
flabel metal3 s -960 358308 480 358548 0 FreeSans 960 0 0 0 io_out[30]
port 128 nsew signal tristate
flabel metal3 s -960 306084 480 306324 0 FreeSans 960 0 0 0 io_out[31]
port 129 nsew signal tristate
flabel metal3 s -960 253996 480 254236 0 FreeSans 960 0 0 0 io_out[32]
port 130 nsew signal tristate
flabel metal3 s -960 201772 480 202012 0 FreeSans 960 0 0 0 io_out[33]
port 131 nsew signal tristate
flabel metal3 s -960 149684 480 149924 0 FreeSans 960 0 0 0 io_out[34]
port 132 nsew signal tristate
flabel metal3 s -960 97460 480 97700 0 FreeSans 960 0 0 0 io_out[35]
port 133 nsew signal tristate
flabel metal3 s -960 58428 480 58668 0 FreeSans 960 0 0 0 io_out[36]
port 134 nsew signal tristate
flabel metal3 s -960 19260 480 19500 0 FreeSans 960 0 0 0 io_out[37]
port 135 nsew signal tristate
flabel metal3 s 583520 139212 584960 139452 0 FreeSans 960 0 0 0 io_out[3]
port 136 nsew signal tristate
flabel metal3 s 583520 179060 584960 179300 0 FreeSans 960 0 0 0 io_out[4]
port 137 nsew signal tristate
flabel metal3 s 583520 218908 584960 219148 0 FreeSans 960 0 0 0 io_out[5]
port 138 nsew signal tristate
flabel metal3 s 583520 258756 584960 258996 0 FreeSans 960 0 0 0 io_out[6]
port 139 nsew signal tristate
flabel metal3 s 583520 311932 584960 312172 0 FreeSans 960 0 0 0 io_out[7]
port 140 nsew signal tristate
flabel metal3 s 583520 364972 584960 365212 0 FreeSans 960 0 0 0 io_out[8]
port 141 nsew signal tristate
flabel metal3 s 583520 418148 584960 418388 0 FreeSans 960 0 0 0 io_out[9]
port 142 nsew signal tristate
flabel metal2 s 125846 -960 125958 480 0 FreeSans 448 90 0 0 la_data_in[0]
port 143 nsew signal input
flabel metal2 s 480506 -960 480618 480 0 FreeSans 448 90 0 0 la_data_in[100]
port 144 nsew signal input
flabel metal2 s 484002 -960 484114 480 0 FreeSans 448 90 0 0 la_data_in[101]
port 145 nsew signal input
flabel metal2 s 487590 -960 487702 480 0 FreeSans 448 90 0 0 la_data_in[102]
port 146 nsew signal input
flabel metal2 s 491086 -960 491198 480 0 FreeSans 448 90 0 0 la_data_in[103]
port 147 nsew signal input
flabel metal2 s 494674 -960 494786 480 0 FreeSans 448 90 0 0 la_data_in[104]
port 148 nsew signal input
flabel metal2 s 498170 -960 498282 480 0 FreeSans 448 90 0 0 la_data_in[105]
port 149 nsew signal input
flabel metal2 s 501758 -960 501870 480 0 FreeSans 448 90 0 0 la_data_in[106]
port 150 nsew signal input
flabel metal2 s 505346 -960 505458 480 0 FreeSans 448 90 0 0 la_data_in[107]
port 151 nsew signal input
flabel metal2 s 508842 -960 508954 480 0 FreeSans 448 90 0 0 la_data_in[108]
port 152 nsew signal input
flabel metal2 s 512430 -960 512542 480 0 FreeSans 448 90 0 0 la_data_in[109]
port 153 nsew signal input
flabel metal2 s 161266 -960 161378 480 0 FreeSans 448 90 0 0 la_data_in[10]
port 154 nsew signal input
flabel metal2 s 515926 -960 516038 480 0 FreeSans 448 90 0 0 la_data_in[110]
port 155 nsew signal input
flabel metal2 s 519514 -960 519626 480 0 FreeSans 448 90 0 0 la_data_in[111]
port 156 nsew signal input
flabel metal2 s 523010 -960 523122 480 0 FreeSans 448 90 0 0 la_data_in[112]
port 157 nsew signal input
flabel metal2 s 526598 -960 526710 480 0 FreeSans 448 90 0 0 la_data_in[113]
port 158 nsew signal input
flabel metal2 s 530094 -960 530206 480 0 FreeSans 448 90 0 0 la_data_in[114]
port 159 nsew signal input
flabel metal2 s 533682 -960 533794 480 0 FreeSans 448 90 0 0 la_data_in[115]
port 160 nsew signal input
flabel metal2 s 537178 -960 537290 480 0 FreeSans 448 90 0 0 la_data_in[116]
port 161 nsew signal input
flabel metal2 s 540766 -960 540878 480 0 FreeSans 448 90 0 0 la_data_in[117]
port 162 nsew signal input
flabel metal2 s 544354 -960 544466 480 0 FreeSans 448 90 0 0 la_data_in[118]
port 163 nsew signal input
flabel metal2 s 547850 -960 547962 480 0 FreeSans 448 90 0 0 la_data_in[119]
port 164 nsew signal input
flabel metal2 s 164854 -960 164966 480 0 FreeSans 448 90 0 0 la_data_in[11]
port 165 nsew signal input
flabel metal2 s 551438 -960 551550 480 0 FreeSans 448 90 0 0 la_data_in[120]
port 166 nsew signal input
flabel metal2 s 554934 -960 555046 480 0 FreeSans 448 90 0 0 la_data_in[121]
port 167 nsew signal input
flabel metal2 s 558522 -960 558634 480 0 FreeSans 448 90 0 0 la_data_in[122]
port 168 nsew signal input
flabel metal2 s 562018 -960 562130 480 0 FreeSans 448 90 0 0 la_data_in[123]
port 169 nsew signal input
flabel metal2 s 565606 -960 565718 480 0 FreeSans 448 90 0 0 la_data_in[124]
port 170 nsew signal input
flabel metal2 s 569102 -960 569214 480 0 FreeSans 448 90 0 0 la_data_in[125]
port 171 nsew signal input
flabel metal2 s 572690 -960 572802 480 0 FreeSans 448 90 0 0 la_data_in[126]
port 172 nsew signal input
flabel metal2 s 576278 -960 576390 480 0 FreeSans 448 90 0 0 la_data_in[127]
port 173 nsew signal input
flabel metal2 s 168350 -960 168462 480 0 FreeSans 448 90 0 0 la_data_in[12]
port 174 nsew signal input
flabel metal2 s 171938 -960 172050 480 0 FreeSans 448 90 0 0 la_data_in[13]
port 175 nsew signal input
flabel metal2 s 175434 -960 175546 480 0 FreeSans 448 90 0 0 la_data_in[14]
port 176 nsew signal input
flabel metal2 s 179022 -960 179134 480 0 FreeSans 448 90 0 0 la_data_in[15]
port 177 nsew signal input
flabel metal2 s 182518 -960 182630 480 0 FreeSans 448 90 0 0 la_data_in[16]
port 178 nsew signal input
flabel metal2 s 186106 -960 186218 480 0 FreeSans 448 90 0 0 la_data_in[17]
port 179 nsew signal input
flabel metal2 s 189694 -960 189806 480 0 FreeSans 448 90 0 0 la_data_in[18]
port 180 nsew signal input
flabel metal2 s 193190 -960 193302 480 0 FreeSans 448 90 0 0 la_data_in[19]
port 181 nsew signal input
flabel metal2 s 129342 -960 129454 480 0 FreeSans 448 90 0 0 la_data_in[1]
port 182 nsew signal input
flabel metal2 s 196778 -960 196890 480 0 FreeSans 448 90 0 0 la_data_in[20]
port 183 nsew signal input
flabel metal2 s 200274 -960 200386 480 0 FreeSans 448 90 0 0 la_data_in[21]
port 184 nsew signal input
flabel metal2 s 203862 -960 203974 480 0 FreeSans 448 90 0 0 la_data_in[22]
port 185 nsew signal input
flabel metal2 s 207358 -960 207470 480 0 FreeSans 448 90 0 0 la_data_in[23]
port 186 nsew signal input
flabel metal2 s 210946 -960 211058 480 0 FreeSans 448 90 0 0 la_data_in[24]
port 187 nsew signal input
flabel metal2 s 214442 -960 214554 480 0 FreeSans 448 90 0 0 la_data_in[25]
port 188 nsew signal input
flabel metal2 s 218030 -960 218142 480 0 FreeSans 448 90 0 0 la_data_in[26]
port 189 nsew signal input
flabel metal2 s 221526 -960 221638 480 0 FreeSans 448 90 0 0 la_data_in[27]
port 190 nsew signal input
flabel metal2 s 225114 -960 225226 480 0 FreeSans 448 90 0 0 la_data_in[28]
port 191 nsew signal input
flabel metal2 s 228702 -960 228814 480 0 FreeSans 448 90 0 0 la_data_in[29]
port 192 nsew signal input
flabel metal2 s 132930 -960 133042 480 0 FreeSans 448 90 0 0 la_data_in[2]
port 193 nsew signal input
flabel metal2 s 232198 -960 232310 480 0 FreeSans 448 90 0 0 la_data_in[30]
port 194 nsew signal input
flabel metal2 s 235786 -960 235898 480 0 FreeSans 448 90 0 0 la_data_in[31]
port 195 nsew signal input
flabel metal2 s 239282 -960 239394 480 0 FreeSans 448 90 0 0 la_data_in[32]
port 196 nsew signal input
flabel metal2 s 242870 -960 242982 480 0 FreeSans 448 90 0 0 la_data_in[33]
port 197 nsew signal input
flabel metal2 s 246366 -960 246478 480 0 FreeSans 448 90 0 0 la_data_in[34]
port 198 nsew signal input
flabel metal2 s 249954 -960 250066 480 0 FreeSans 448 90 0 0 la_data_in[35]
port 199 nsew signal input
flabel metal2 s 253450 -960 253562 480 0 FreeSans 448 90 0 0 la_data_in[36]
port 200 nsew signal input
flabel metal2 s 257038 -960 257150 480 0 FreeSans 448 90 0 0 la_data_in[37]
port 201 nsew signal input
flabel metal2 s 260626 -960 260738 480 0 FreeSans 448 90 0 0 la_data_in[38]
port 202 nsew signal input
flabel metal2 s 264122 -960 264234 480 0 FreeSans 448 90 0 0 la_data_in[39]
port 203 nsew signal input
flabel metal2 s 136426 -960 136538 480 0 FreeSans 448 90 0 0 la_data_in[3]
port 204 nsew signal input
flabel metal2 s 267710 -960 267822 480 0 FreeSans 448 90 0 0 la_data_in[40]
port 205 nsew signal input
flabel metal2 s 271206 -960 271318 480 0 FreeSans 448 90 0 0 la_data_in[41]
port 206 nsew signal input
flabel metal2 s 274794 -960 274906 480 0 FreeSans 448 90 0 0 la_data_in[42]
port 207 nsew signal input
flabel metal2 s 278290 -960 278402 480 0 FreeSans 448 90 0 0 la_data_in[43]
port 208 nsew signal input
flabel metal2 s 281878 -960 281990 480 0 FreeSans 448 90 0 0 la_data_in[44]
port 209 nsew signal input
flabel metal2 s 285374 -960 285486 480 0 FreeSans 448 90 0 0 la_data_in[45]
port 210 nsew signal input
flabel metal2 s 288962 -960 289074 480 0 FreeSans 448 90 0 0 la_data_in[46]
port 211 nsew signal input
flabel metal2 s 292550 -960 292662 480 0 FreeSans 448 90 0 0 la_data_in[47]
port 212 nsew signal input
flabel metal2 s 296046 -960 296158 480 0 FreeSans 448 90 0 0 la_data_in[48]
port 213 nsew signal input
flabel metal2 s 299634 -960 299746 480 0 FreeSans 448 90 0 0 la_data_in[49]
port 214 nsew signal input
flabel metal2 s 140014 -960 140126 480 0 FreeSans 448 90 0 0 la_data_in[4]
port 215 nsew signal input
flabel metal2 s 303130 -960 303242 480 0 FreeSans 448 90 0 0 la_data_in[50]
port 216 nsew signal input
flabel metal2 s 306718 -960 306830 480 0 FreeSans 448 90 0 0 la_data_in[51]
port 217 nsew signal input
flabel metal2 s 310214 -960 310326 480 0 FreeSans 448 90 0 0 la_data_in[52]
port 218 nsew signal input
flabel metal2 s 313802 -960 313914 480 0 FreeSans 448 90 0 0 la_data_in[53]
port 219 nsew signal input
flabel metal2 s 317298 -960 317410 480 0 FreeSans 448 90 0 0 la_data_in[54]
port 220 nsew signal input
flabel metal2 s 320886 -960 320998 480 0 FreeSans 448 90 0 0 la_data_in[55]
port 221 nsew signal input
flabel metal2 s 324382 -960 324494 480 0 FreeSans 448 90 0 0 la_data_in[56]
port 222 nsew signal input
flabel metal2 s 327970 -960 328082 480 0 FreeSans 448 90 0 0 la_data_in[57]
port 223 nsew signal input
flabel metal2 s 331558 -960 331670 480 0 FreeSans 448 90 0 0 la_data_in[58]
port 224 nsew signal input
flabel metal2 s 335054 -960 335166 480 0 FreeSans 448 90 0 0 la_data_in[59]
port 225 nsew signal input
flabel metal2 s 143510 -960 143622 480 0 FreeSans 448 90 0 0 la_data_in[5]
port 226 nsew signal input
flabel metal2 s 338642 -960 338754 480 0 FreeSans 448 90 0 0 la_data_in[60]
port 227 nsew signal input
flabel metal2 s 342138 -960 342250 480 0 FreeSans 448 90 0 0 la_data_in[61]
port 228 nsew signal input
flabel metal2 s 345726 -960 345838 480 0 FreeSans 448 90 0 0 la_data_in[62]
port 229 nsew signal input
flabel metal2 s 349222 -960 349334 480 0 FreeSans 448 90 0 0 la_data_in[63]
port 230 nsew signal input
flabel metal2 s 352810 -960 352922 480 0 FreeSans 448 90 0 0 la_data_in[64]
port 231 nsew signal input
flabel metal2 s 356306 -960 356418 480 0 FreeSans 448 90 0 0 la_data_in[65]
port 232 nsew signal input
flabel metal2 s 359894 -960 360006 480 0 FreeSans 448 90 0 0 la_data_in[66]
port 233 nsew signal input
flabel metal2 s 363482 -960 363594 480 0 FreeSans 448 90 0 0 la_data_in[67]
port 234 nsew signal input
flabel metal2 s 366978 -960 367090 480 0 FreeSans 448 90 0 0 la_data_in[68]
port 235 nsew signal input
flabel metal2 s 370566 -960 370678 480 0 FreeSans 448 90 0 0 la_data_in[69]
port 236 nsew signal input
flabel metal2 s 147098 -960 147210 480 0 FreeSans 448 90 0 0 la_data_in[6]
port 237 nsew signal input
flabel metal2 s 374062 -960 374174 480 0 FreeSans 448 90 0 0 la_data_in[70]
port 238 nsew signal input
flabel metal2 s 377650 -960 377762 480 0 FreeSans 448 90 0 0 la_data_in[71]
port 239 nsew signal input
flabel metal2 s 381146 -960 381258 480 0 FreeSans 448 90 0 0 la_data_in[72]
port 240 nsew signal input
flabel metal2 s 384734 -960 384846 480 0 FreeSans 448 90 0 0 la_data_in[73]
port 241 nsew signal input
flabel metal2 s 388230 -960 388342 480 0 FreeSans 448 90 0 0 la_data_in[74]
port 242 nsew signal input
flabel metal2 s 391818 -960 391930 480 0 FreeSans 448 90 0 0 la_data_in[75]
port 243 nsew signal input
flabel metal2 s 395314 -960 395426 480 0 FreeSans 448 90 0 0 la_data_in[76]
port 244 nsew signal input
flabel metal2 s 398902 -960 399014 480 0 FreeSans 448 90 0 0 la_data_in[77]
port 245 nsew signal input
flabel metal2 s 402490 -960 402602 480 0 FreeSans 448 90 0 0 la_data_in[78]
port 246 nsew signal input
flabel metal2 s 405986 -960 406098 480 0 FreeSans 448 90 0 0 la_data_in[79]
port 247 nsew signal input
flabel metal2 s 150594 -960 150706 480 0 FreeSans 448 90 0 0 la_data_in[7]
port 248 nsew signal input
flabel metal2 s 409574 -960 409686 480 0 FreeSans 448 90 0 0 la_data_in[80]
port 249 nsew signal input
flabel metal2 s 413070 -960 413182 480 0 FreeSans 448 90 0 0 la_data_in[81]
port 250 nsew signal input
flabel metal2 s 416658 -960 416770 480 0 FreeSans 448 90 0 0 la_data_in[82]
port 251 nsew signal input
flabel metal2 s 420154 -960 420266 480 0 FreeSans 448 90 0 0 la_data_in[83]
port 252 nsew signal input
flabel metal2 s 423742 -960 423854 480 0 FreeSans 448 90 0 0 la_data_in[84]
port 253 nsew signal input
flabel metal2 s 427238 -960 427350 480 0 FreeSans 448 90 0 0 la_data_in[85]
port 254 nsew signal input
flabel metal2 s 430826 -960 430938 480 0 FreeSans 448 90 0 0 la_data_in[86]
port 255 nsew signal input
flabel metal2 s 434414 -960 434526 480 0 FreeSans 448 90 0 0 la_data_in[87]
port 256 nsew signal input
flabel metal2 s 437910 -960 438022 480 0 FreeSans 448 90 0 0 la_data_in[88]
port 257 nsew signal input
flabel metal2 s 441498 -960 441610 480 0 FreeSans 448 90 0 0 la_data_in[89]
port 258 nsew signal input
flabel metal2 s 154182 -960 154294 480 0 FreeSans 448 90 0 0 la_data_in[8]
port 259 nsew signal input
flabel metal2 s 444994 -960 445106 480 0 FreeSans 448 90 0 0 la_data_in[90]
port 260 nsew signal input
flabel metal2 s 448582 -960 448694 480 0 FreeSans 448 90 0 0 la_data_in[91]
port 261 nsew signal input
flabel metal2 s 452078 -960 452190 480 0 FreeSans 448 90 0 0 la_data_in[92]
port 262 nsew signal input
flabel metal2 s 455666 -960 455778 480 0 FreeSans 448 90 0 0 la_data_in[93]
port 263 nsew signal input
flabel metal2 s 459162 -960 459274 480 0 FreeSans 448 90 0 0 la_data_in[94]
port 264 nsew signal input
flabel metal2 s 462750 -960 462862 480 0 FreeSans 448 90 0 0 la_data_in[95]
port 265 nsew signal input
flabel metal2 s 466246 -960 466358 480 0 FreeSans 448 90 0 0 la_data_in[96]
port 266 nsew signal input
flabel metal2 s 469834 -960 469946 480 0 FreeSans 448 90 0 0 la_data_in[97]
port 267 nsew signal input
flabel metal2 s 473422 -960 473534 480 0 FreeSans 448 90 0 0 la_data_in[98]
port 268 nsew signal input
flabel metal2 s 476918 -960 477030 480 0 FreeSans 448 90 0 0 la_data_in[99]
port 269 nsew signal input
flabel metal2 s 157770 -960 157882 480 0 FreeSans 448 90 0 0 la_data_in[9]
port 270 nsew signal input
flabel metal2 s 126950 -960 127062 480 0 FreeSans 448 90 0 0 la_data_out[0]
port 271 nsew signal tristate
flabel metal2 s 481702 -960 481814 480 0 FreeSans 448 90 0 0 la_data_out[100]
port 272 nsew signal tristate
flabel metal2 s 485198 -960 485310 480 0 FreeSans 448 90 0 0 la_data_out[101]
port 273 nsew signal tristate
flabel metal2 s 488786 -960 488898 480 0 FreeSans 448 90 0 0 la_data_out[102]
port 274 nsew signal tristate
flabel metal2 s 492282 -960 492394 480 0 FreeSans 448 90 0 0 la_data_out[103]
port 275 nsew signal tristate
flabel metal2 s 495870 -960 495982 480 0 FreeSans 448 90 0 0 la_data_out[104]
port 276 nsew signal tristate
flabel metal2 s 499366 -960 499478 480 0 FreeSans 448 90 0 0 la_data_out[105]
port 277 nsew signal tristate
flabel metal2 s 502954 -960 503066 480 0 FreeSans 448 90 0 0 la_data_out[106]
port 278 nsew signal tristate
flabel metal2 s 506450 -960 506562 480 0 FreeSans 448 90 0 0 la_data_out[107]
port 279 nsew signal tristate
flabel metal2 s 510038 -960 510150 480 0 FreeSans 448 90 0 0 la_data_out[108]
port 280 nsew signal tristate
flabel metal2 s 513534 -960 513646 480 0 FreeSans 448 90 0 0 la_data_out[109]
port 281 nsew signal tristate
flabel metal2 s 162462 -960 162574 480 0 FreeSans 448 90 0 0 la_data_out[10]
port 282 nsew signal tristate
flabel metal2 s 517122 -960 517234 480 0 FreeSans 448 90 0 0 la_data_out[110]
port 283 nsew signal tristate
flabel metal2 s 520710 -960 520822 480 0 FreeSans 448 90 0 0 la_data_out[111]
port 284 nsew signal tristate
flabel metal2 s 524206 -960 524318 480 0 FreeSans 448 90 0 0 la_data_out[112]
port 285 nsew signal tristate
flabel metal2 s 527794 -960 527906 480 0 FreeSans 448 90 0 0 la_data_out[113]
port 286 nsew signal tristate
flabel metal2 s 531290 -960 531402 480 0 FreeSans 448 90 0 0 la_data_out[114]
port 287 nsew signal tristate
flabel metal2 s 534878 -960 534990 480 0 FreeSans 448 90 0 0 la_data_out[115]
port 288 nsew signal tristate
flabel metal2 s 538374 -960 538486 480 0 FreeSans 448 90 0 0 la_data_out[116]
port 289 nsew signal tristate
flabel metal2 s 541962 -960 542074 480 0 FreeSans 448 90 0 0 la_data_out[117]
port 290 nsew signal tristate
flabel metal2 s 545458 -960 545570 480 0 FreeSans 448 90 0 0 la_data_out[118]
port 291 nsew signal tristate
flabel metal2 s 549046 -960 549158 480 0 FreeSans 448 90 0 0 la_data_out[119]
port 292 nsew signal tristate
flabel metal2 s 166050 -960 166162 480 0 FreeSans 448 90 0 0 la_data_out[11]
port 293 nsew signal tristate
flabel metal2 s 552634 -960 552746 480 0 FreeSans 448 90 0 0 la_data_out[120]
port 294 nsew signal tristate
flabel metal2 s 556130 -960 556242 480 0 FreeSans 448 90 0 0 la_data_out[121]
port 295 nsew signal tristate
flabel metal2 s 559718 -960 559830 480 0 FreeSans 448 90 0 0 la_data_out[122]
port 296 nsew signal tristate
flabel metal2 s 563214 -960 563326 480 0 FreeSans 448 90 0 0 la_data_out[123]
port 297 nsew signal tristate
flabel metal2 s 566802 -960 566914 480 0 FreeSans 448 90 0 0 la_data_out[124]
port 298 nsew signal tristate
flabel metal2 s 570298 -960 570410 480 0 FreeSans 448 90 0 0 la_data_out[125]
port 299 nsew signal tristate
flabel metal2 s 573886 -960 573998 480 0 FreeSans 448 90 0 0 la_data_out[126]
port 300 nsew signal tristate
flabel metal2 s 577382 -960 577494 480 0 FreeSans 448 90 0 0 la_data_out[127]
port 301 nsew signal tristate
flabel metal2 s 169546 -960 169658 480 0 FreeSans 448 90 0 0 la_data_out[12]
port 302 nsew signal tristate
flabel metal2 s 173134 -960 173246 480 0 FreeSans 448 90 0 0 la_data_out[13]
port 303 nsew signal tristate
flabel metal2 s 176630 -960 176742 480 0 FreeSans 448 90 0 0 la_data_out[14]
port 304 nsew signal tristate
flabel metal2 s 180218 -960 180330 480 0 FreeSans 448 90 0 0 la_data_out[15]
port 305 nsew signal tristate
flabel metal2 s 183714 -960 183826 480 0 FreeSans 448 90 0 0 la_data_out[16]
port 306 nsew signal tristate
flabel metal2 s 187302 -960 187414 480 0 FreeSans 448 90 0 0 la_data_out[17]
port 307 nsew signal tristate
flabel metal2 s 190798 -960 190910 480 0 FreeSans 448 90 0 0 la_data_out[18]
port 308 nsew signal tristate
flabel metal2 s 194386 -960 194498 480 0 FreeSans 448 90 0 0 la_data_out[19]
port 309 nsew signal tristate
flabel metal2 s 130538 -960 130650 480 0 FreeSans 448 90 0 0 la_data_out[1]
port 310 nsew signal tristate
flabel metal2 s 197882 -960 197994 480 0 FreeSans 448 90 0 0 la_data_out[20]
port 311 nsew signal tristate
flabel metal2 s 201470 -960 201582 480 0 FreeSans 448 90 0 0 la_data_out[21]
port 312 nsew signal tristate
flabel metal2 s 205058 -960 205170 480 0 FreeSans 448 90 0 0 la_data_out[22]
port 313 nsew signal tristate
flabel metal2 s 208554 -960 208666 480 0 FreeSans 448 90 0 0 la_data_out[23]
port 314 nsew signal tristate
flabel metal2 s 212142 -960 212254 480 0 FreeSans 448 90 0 0 la_data_out[24]
port 315 nsew signal tristate
flabel metal2 s 215638 -960 215750 480 0 FreeSans 448 90 0 0 la_data_out[25]
port 316 nsew signal tristate
flabel metal2 s 219226 -960 219338 480 0 FreeSans 448 90 0 0 la_data_out[26]
port 317 nsew signal tristate
flabel metal2 s 222722 -960 222834 480 0 FreeSans 448 90 0 0 la_data_out[27]
port 318 nsew signal tristate
flabel metal2 s 226310 -960 226422 480 0 FreeSans 448 90 0 0 la_data_out[28]
port 319 nsew signal tristate
flabel metal2 s 229806 -960 229918 480 0 FreeSans 448 90 0 0 la_data_out[29]
port 320 nsew signal tristate
flabel metal2 s 134126 -960 134238 480 0 FreeSans 448 90 0 0 la_data_out[2]
port 321 nsew signal tristate
flabel metal2 s 233394 -960 233506 480 0 FreeSans 448 90 0 0 la_data_out[30]
port 322 nsew signal tristate
flabel metal2 s 236982 -960 237094 480 0 FreeSans 448 90 0 0 la_data_out[31]
port 323 nsew signal tristate
flabel metal2 s 240478 -960 240590 480 0 FreeSans 448 90 0 0 la_data_out[32]
port 324 nsew signal tristate
flabel metal2 s 244066 -960 244178 480 0 FreeSans 448 90 0 0 la_data_out[33]
port 325 nsew signal tristate
flabel metal2 s 247562 -960 247674 480 0 FreeSans 448 90 0 0 la_data_out[34]
port 326 nsew signal tristate
flabel metal2 s 251150 -960 251262 480 0 FreeSans 448 90 0 0 la_data_out[35]
port 327 nsew signal tristate
flabel metal2 s 254646 -960 254758 480 0 FreeSans 448 90 0 0 la_data_out[36]
port 328 nsew signal tristate
flabel metal2 s 258234 -960 258346 480 0 FreeSans 448 90 0 0 la_data_out[37]
port 329 nsew signal tristate
flabel metal2 s 261730 -960 261842 480 0 FreeSans 448 90 0 0 la_data_out[38]
port 330 nsew signal tristate
flabel metal2 s 265318 -960 265430 480 0 FreeSans 448 90 0 0 la_data_out[39]
port 331 nsew signal tristate
flabel metal2 s 137622 -960 137734 480 0 FreeSans 448 90 0 0 la_data_out[3]
port 332 nsew signal tristate
flabel metal2 s 268814 -960 268926 480 0 FreeSans 448 90 0 0 la_data_out[40]
port 333 nsew signal tristate
flabel metal2 s 272402 -960 272514 480 0 FreeSans 448 90 0 0 la_data_out[41]
port 334 nsew signal tristate
flabel metal2 s 275990 -960 276102 480 0 FreeSans 448 90 0 0 la_data_out[42]
port 335 nsew signal tristate
flabel metal2 s 279486 -960 279598 480 0 FreeSans 448 90 0 0 la_data_out[43]
port 336 nsew signal tristate
flabel metal2 s 283074 -960 283186 480 0 FreeSans 448 90 0 0 la_data_out[44]
port 337 nsew signal tristate
flabel metal2 s 286570 -960 286682 480 0 FreeSans 448 90 0 0 la_data_out[45]
port 338 nsew signal tristate
flabel metal2 s 290158 -960 290270 480 0 FreeSans 448 90 0 0 la_data_out[46]
port 339 nsew signal tristate
flabel metal2 s 293654 -960 293766 480 0 FreeSans 448 90 0 0 la_data_out[47]
port 340 nsew signal tristate
flabel metal2 s 297242 -960 297354 480 0 FreeSans 448 90 0 0 la_data_out[48]
port 341 nsew signal tristate
flabel metal2 s 300738 -960 300850 480 0 FreeSans 448 90 0 0 la_data_out[49]
port 342 nsew signal tristate
flabel metal2 s 141210 -960 141322 480 0 FreeSans 448 90 0 0 la_data_out[4]
port 343 nsew signal tristate
flabel metal2 s 304326 -960 304438 480 0 FreeSans 448 90 0 0 la_data_out[50]
port 344 nsew signal tristate
flabel metal2 s 307914 -960 308026 480 0 FreeSans 448 90 0 0 la_data_out[51]
port 345 nsew signal tristate
flabel metal2 s 311410 -960 311522 480 0 FreeSans 448 90 0 0 la_data_out[52]
port 346 nsew signal tristate
flabel metal2 s 314998 -960 315110 480 0 FreeSans 448 90 0 0 la_data_out[53]
port 347 nsew signal tristate
flabel metal2 s 318494 -960 318606 480 0 FreeSans 448 90 0 0 la_data_out[54]
port 348 nsew signal tristate
flabel metal2 s 322082 -960 322194 480 0 FreeSans 448 90 0 0 la_data_out[55]
port 349 nsew signal tristate
flabel metal2 s 325578 -960 325690 480 0 FreeSans 448 90 0 0 la_data_out[56]
port 350 nsew signal tristate
flabel metal2 s 329166 -960 329278 480 0 FreeSans 448 90 0 0 la_data_out[57]
port 351 nsew signal tristate
flabel metal2 s 332662 -960 332774 480 0 FreeSans 448 90 0 0 la_data_out[58]
port 352 nsew signal tristate
flabel metal2 s 336250 -960 336362 480 0 FreeSans 448 90 0 0 la_data_out[59]
port 353 nsew signal tristate
flabel metal2 s 144706 -960 144818 480 0 FreeSans 448 90 0 0 la_data_out[5]
port 354 nsew signal tristate
flabel metal2 s 339838 -960 339950 480 0 FreeSans 448 90 0 0 la_data_out[60]
port 355 nsew signal tristate
flabel metal2 s 343334 -960 343446 480 0 FreeSans 448 90 0 0 la_data_out[61]
port 356 nsew signal tristate
flabel metal2 s 346922 -960 347034 480 0 FreeSans 448 90 0 0 la_data_out[62]
port 357 nsew signal tristate
flabel metal2 s 350418 -960 350530 480 0 FreeSans 448 90 0 0 la_data_out[63]
port 358 nsew signal tristate
flabel metal2 s 354006 -960 354118 480 0 FreeSans 448 90 0 0 la_data_out[64]
port 359 nsew signal tristate
flabel metal2 s 357502 -960 357614 480 0 FreeSans 448 90 0 0 la_data_out[65]
port 360 nsew signal tristate
flabel metal2 s 361090 -960 361202 480 0 FreeSans 448 90 0 0 la_data_out[66]
port 361 nsew signal tristate
flabel metal2 s 364586 -960 364698 480 0 FreeSans 448 90 0 0 la_data_out[67]
port 362 nsew signal tristate
flabel metal2 s 368174 -960 368286 480 0 FreeSans 448 90 0 0 la_data_out[68]
port 363 nsew signal tristate
flabel metal2 s 371670 -960 371782 480 0 FreeSans 448 90 0 0 la_data_out[69]
port 364 nsew signal tristate
flabel metal2 s 148294 -960 148406 480 0 FreeSans 448 90 0 0 la_data_out[6]
port 365 nsew signal tristate
flabel metal2 s 375258 -960 375370 480 0 FreeSans 448 90 0 0 la_data_out[70]
port 366 nsew signal tristate
flabel metal2 s 378846 -960 378958 480 0 FreeSans 448 90 0 0 la_data_out[71]
port 367 nsew signal tristate
flabel metal2 s 382342 -960 382454 480 0 FreeSans 448 90 0 0 la_data_out[72]
port 368 nsew signal tristate
flabel metal2 s 385930 -960 386042 480 0 FreeSans 448 90 0 0 la_data_out[73]
port 369 nsew signal tristate
flabel metal2 s 389426 -960 389538 480 0 FreeSans 448 90 0 0 la_data_out[74]
port 370 nsew signal tristate
flabel metal2 s 393014 -960 393126 480 0 FreeSans 448 90 0 0 la_data_out[75]
port 371 nsew signal tristate
flabel metal2 s 396510 -960 396622 480 0 FreeSans 448 90 0 0 la_data_out[76]
port 372 nsew signal tristate
flabel metal2 s 400098 -960 400210 480 0 FreeSans 448 90 0 0 la_data_out[77]
port 373 nsew signal tristate
flabel metal2 s 403594 -960 403706 480 0 FreeSans 448 90 0 0 la_data_out[78]
port 374 nsew signal tristate
flabel metal2 s 407182 -960 407294 480 0 FreeSans 448 90 0 0 la_data_out[79]
port 375 nsew signal tristate
flabel metal2 s 151790 -960 151902 480 0 FreeSans 448 90 0 0 la_data_out[7]
port 376 nsew signal tristate
flabel metal2 s 410770 -960 410882 480 0 FreeSans 448 90 0 0 la_data_out[80]
port 377 nsew signal tristate
flabel metal2 s 414266 -960 414378 480 0 FreeSans 448 90 0 0 la_data_out[81]
port 378 nsew signal tristate
flabel metal2 s 417854 -960 417966 480 0 FreeSans 448 90 0 0 la_data_out[82]
port 379 nsew signal tristate
flabel metal2 s 421350 -960 421462 480 0 FreeSans 448 90 0 0 la_data_out[83]
port 380 nsew signal tristate
flabel metal2 s 424938 -960 425050 480 0 FreeSans 448 90 0 0 la_data_out[84]
port 381 nsew signal tristate
flabel metal2 s 428434 -960 428546 480 0 FreeSans 448 90 0 0 la_data_out[85]
port 382 nsew signal tristate
flabel metal2 s 432022 -960 432134 480 0 FreeSans 448 90 0 0 la_data_out[86]
port 383 nsew signal tristate
flabel metal2 s 435518 -960 435630 480 0 FreeSans 448 90 0 0 la_data_out[87]
port 384 nsew signal tristate
flabel metal2 s 439106 -960 439218 480 0 FreeSans 448 90 0 0 la_data_out[88]
port 385 nsew signal tristate
flabel metal2 s 442602 -960 442714 480 0 FreeSans 448 90 0 0 la_data_out[89]
port 386 nsew signal tristate
flabel metal2 s 155378 -960 155490 480 0 FreeSans 448 90 0 0 la_data_out[8]
port 387 nsew signal tristate
flabel metal2 s 446190 -960 446302 480 0 FreeSans 448 90 0 0 la_data_out[90]
port 388 nsew signal tristate
flabel metal2 s 449778 -960 449890 480 0 FreeSans 448 90 0 0 la_data_out[91]
port 389 nsew signal tristate
flabel metal2 s 453274 -960 453386 480 0 FreeSans 448 90 0 0 la_data_out[92]
port 390 nsew signal tristate
flabel metal2 s 456862 -960 456974 480 0 FreeSans 448 90 0 0 la_data_out[93]
port 391 nsew signal tristate
flabel metal2 s 460358 -960 460470 480 0 FreeSans 448 90 0 0 la_data_out[94]
port 392 nsew signal tristate
flabel metal2 s 463946 -960 464058 480 0 FreeSans 448 90 0 0 la_data_out[95]
port 393 nsew signal tristate
flabel metal2 s 467442 -960 467554 480 0 FreeSans 448 90 0 0 la_data_out[96]
port 394 nsew signal tristate
flabel metal2 s 471030 -960 471142 480 0 FreeSans 448 90 0 0 la_data_out[97]
port 395 nsew signal tristate
flabel metal2 s 474526 -960 474638 480 0 FreeSans 448 90 0 0 la_data_out[98]
port 396 nsew signal tristate
flabel metal2 s 478114 -960 478226 480 0 FreeSans 448 90 0 0 la_data_out[99]
port 397 nsew signal tristate
flabel metal2 s 158874 -960 158986 480 0 FreeSans 448 90 0 0 la_data_out[9]
port 398 nsew signal tristate
flabel metal2 s 128146 -960 128258 480 0 FreeSans 448 90 0 0 la_oenb[0]
port 399 nsew signal input
flabel metal2 s 482806 -960 482918 480 0 FreeSans 448 90 0 0 la_oenb[100]
port 400 nsew signal input
flabel metal2 s 486394 -960 486506 480 0 FreeSans 448 90 0 0 la_oenb[101]
port 401 nsew signal input
flabel metal2 s 489890 -960 490002 480 0 FreeSans 448 90 0 0 la_oenb[102]
port 402 nsew signal input
flabel metal2 s 493478 -960 493590 480 0 FreeSans 448 90 0 0 la_oenb[103]
port 403 nsew signal input
flabel metal2 s 497066 -960 497178 480 0 FreeSans 448 90 0 0 la_oenb[104]
port 404 nsew signal input
flabel metal2 s 500562 -960 500674 480 0 FreeSans 448 90 0 0 la_oenb[105]
port 405 nsew signal input
flabel metal2 s 504150 -960 504262 480 0 FreeSans 448 90 0 0 la_oenb[106]
port 406 nsew signal input
flabel metal2 s 507646 -960 507758 480 0 FreeSans 448 90 0 0 la_oenb[107]
port 407 nsew signal input
flabel metal2 s 511234 -960 511346 480 0 FreeSans 448 90 0 0 la_oenb[108]
port 408 nsew signal input
flabel metal2 s 514730 -960 514842 480 0 FreeSans 448 90 0 0 la_oenb[109]
port 409 nsew signal input
flabel metal2 s 163658 -960 163770 480 0 FreeSans 448 90 0 0 la_oenb[10]
port 410 nsew signal input
flabel metal2 s 518318 -960 518430 480 0 FreeSans 448 90 0 0 la_oenb[110]
port 411 nsew signal input
flabel metal2 s 521814 -960 521926 480 0 FreeSans 448 90 0 0 la_oenb[111]
port 412 nsew signal input
flabel metal2 s 525402 -960 525514 480 0 FreeSans 448 90 0 0 la_oenb[112]
port 413 nsew signal input
flabel metal2 s 528990 -960 529102 480 0 FreeSans 448 90 0 0 la_oenb[113]
port 414 nsew signal input
flabel metal2 s 532486 -960 532598 480 0 FreeSans 448 90 0 0 la_oenb[114]
port 415 nsew signal input
flabel metal2 s 536074 -960 536186 480 0 FreeSans 448 90 0 0 la_oenb[115]
port 416 nsew signal input
flabel metal2 s 539570 -960 539682 480 0 FreeSans 448 90 0 0 la_oenb[116]
port 417 nsew signal input
flabel metal2 s 543158 -960 543270 480 0 FreeSans 448 90 0 0 la_oenb[117]
port 418 nsew signal input
flabel metal2 s 546654 -960 546766 480 0 FreeSans 448 90 0 0 la_oenb[118]
port 419 nsew signal input
flabel metal2 s 550242 -960 550354 480 0 FreeSans 448 90 0 0 la_oenb[119]
port 420 nsew signal input
flabel metal2 s 167154 -960 167266 480 0 FreeSans 448 90 0 0 la_oenb[11]
port 421 nsew signal input
flabel metal2 s 553738 -960 553850 480 0 FreeSans 448 90 0 0 la_oenb[120]
port 422 nsew signal input
flabel metal2 s 557326 -960 557438 480 0 FreeSans 448 90 0 0 la_oenb[121]
port 423 nsew signal input
flabel metal2 s 560822 -960 560934 480 0 FreeSans 448 90 0 0 la_oenb[122]
port 424 nsew signal input
flabel metal2 s 564410 -960 564522 480 0 FreeSans 448 90 0 0 la_oenb[123]
port 425 nsew signal input
flabel metal2 s 567998 -960 568110 480 0 FreeSans 448 90 0 0 la_oenb[124]
port 426 nsew signal input
flabel metal2 s 571494 -960 571606 480 0 FreeSans 448 90 0 0 la_oenb[125]
port 427 nsew signal input
flabel metal2 s 575082 -960 575194 480 0 FreeSans 448 90 0 0 la_oenb[126]
port 428 nsew signal input
flabel metal2 s 578578 -960 578690 480 0 FreeSans 448 90 0 0 la_oenb[127]
port 429 nsew signal input
flabel metal2 s 170742 -960 170854 480 0 FreeSans 448 90 0 0 la_oenb[12]
port 430 nsew signal input
flabel metal2 s 174238 -960 174350 480 0 FreeSans 448 90 0 0 la_oenb[13]
port 431 nsew signal input
flabel metal2 s 177826 -960 177938 480 0 FreeSans 448 90 0 0 la_oenb[14]
port 432 nsew signal input
flabel metal2 s 181414 -960 181526 480 0 FreeSans 448 90 0 0 la_oenb[15]
port 433 nsew signal input
flabel metal2 s 184910 -960 185022 480 0 FreeSans 448 90 0 0 la_oenb[16]
port 434 nsew signal input
flabel metal2 s 188498 -960 188610 480 0 FreeSans 448 90 0 0 la_oenb[17]
port 435 nsew signal input
flabel metal2 s 191994 -960 192106 480 0 FreeSans 448 90 0 0 la_oenb[18]
port 436 nsew signal input
flabel metal2 s 195582 -960 195694 480 0 FreeSans 448 90 0 0 la_oenb[19]
port 437 nsew signal input
flabel metal2 s 131734 -960 131846 480 0 FreeSans 448 90 0 0 la_oenb[1]
port 438 nsew signal input
flabel metal2 s 199078 -960 199190 480 0 FreeSans 448 90 0 0 la_oenb[20]
port 439 nsew signal input
flabel metal2 s 202666 -960 202778 480 0 FreeSans 448 90 0 0 la_oenb[21]
port 440 nsew signal input
flabel metal2 s 206162 -960 206274 480 0 FreeSans 448 90 0 0 la_oenb[22]
port 441 nsew signal input
flabel metal2 s 209750 -960 209862 480 0 FreeSans 448 90 0 0 la_oenb[23]
port 442 nsew signal input
flabel metal2 s 213338 -960 213450 480 0 FreeSans 448 90 0 0 la_oenb[24]
port 443 nsew signal input
flabel metal2 s 216834 -960 216946 480 0 FreeSans 448 90 0 0 la_oenb[25]
port 444 nsew signal input
flabel metal2 s 220422 -960 220534 480 0 FreeSans 448 90 0 0 la_oenb[26]
port 445 nsew signal input
flabel metal2 s 223918 -960 224030 480 0 FreeSans 448 90 0 0 la_oenb[27]
port 446 nsew signal input
flabel metal2 s 227506 -960 227618 480 0 FreeSans 448 90 0 0 la_oenb[28]
port 447 nsew signal input
flabel metal2 s 231002 -960 231114 480 0 FreeSans 448 90 0 0 la_oenb[29]
port 448 nsew signal input
flabel metal2 s 135230 -960 135342 480 0 FreeSans 448 90 0 0 la_oenb[2]
port 449 nsew signal input
flabel metal2 s 234590 -960 234702 480 0 FreeSans 448 90 0 0 la_oenb[30]
port 450 nsew signal input
flabel metal2 s 238086 -960 238198 480 0 FreeSans 448 90 0 0 la_oenb[31]
port 451 nsew signal input
flabel metal2 s 241674 -960 241786 480 0 FreeSans 448 90 0 0 la_oenb[32]
port 452 nsew signal input
flabel metal2 s 245170 -960 245282 480 0 FreeSans 448 90 0 0 la_oenb[33]
port 453 nsew signal input
flabel metal2 s 248758 -960 248870 480 0 FreeSans 448 90 0 0 la_oenb[34]
port 454 nsew signal input
flabel metal2 s 252346 -960 252458 480 0 FreeSans 448 90 0 0 la_oenb[35]
port 455 nsew signal input
flabel metal2 s 255842 -960 255954 480 0 FreeSans 448 90 0 0 la_oenb[36]
port 456 nsew signal input
flabel metal2 s 259430 -960 259542 480 0 FreeSans 448 90 0 0 la_oenb[37]
port 457 nsew signal input
flabel metal2 s 262926 -960 263038 480 0 FreeSans 448 90 0 0 la_oenb[38]
port 458 nsew signal input
flabel metal2 s 266514 -960 266626 480 0 FreeSans 448 90 0 0 la_oenb[39]
port 459 nsew signal input
flabel metal2 s 138818 -960 138930 480 0 FreeSans 448 90 0 0 la_oenb[3]
port 460 nsew signal input
flabel metal2 s 270010 -960 270122 480 0 FreeSans 448 90 0 0 la_oenb[40]
port 461 nsew signal input
flabel metal2 s 273598 -960 273710 480 0 FreeSans 448 90 0 0 la_oenb[41]
port 462 nsew signal input
flabel metal2 s 277094 -960 277206 480 0 FreeSans 448 90 0 0 la_oenb[42]
port 463 nsew signal input
flabel metal2 s 280682 -960 280794 480 0 FreeSans 448 90 0 0 la_oenb[43]
port 464 nsew signal input
flabel metal2 s 284270 -960 284382 480 0 FreeSans 448 90 0 0 la_oenb[44]
port 465 nsew signal input
flabel metal2 s 287766 -960 287878 480 0 FreeSans 448 90 0 0 la_oenb[45]
port 466 nsew signal input
flabel metal2 s 291354 -960 291466 480 0 FreeSans 448 90 0 0 la_oenb[46]
port 467 nsew signal input
flabel metal2 s 294850 -960 294962 480 0 FreeSans 448 90 0 0 la_oenb[47]
port 468 nsew signal input
flabel metal2 s 298438 -960 298550 480 0 FreeSans 448 90 0 0 la_oenb[48]
port 469 nsew signal input
flabel metal2 s 301934 -960 302046 480 0 FreeSans 448 90 0 0 la_oenb[49]
port 470 nsew signal input
flabel metal2 s 142406 -960 142518 480 0 FreeSans 448 90 0 0 la_oenb[4]
port 471 nsew signal input
flabel metal2 s 305522 -960 305634 480 0 FreeSans 448 90 0 0 la_oenb[50]
port 472 nsew signal input
flabel metal2 s 309018 -960 309130 480 0 FreeSans 448 90 0 0 la_oenb[51]
port 473 nsew signal input
flabel metal2 s 312606 -960 312718 480 0 FreeSans 448 90 0 0 la_oenb[52]
port 474 nsew signal input
flabel metal2 s 316194 -960 316306 480 0 FreeSans 448 90 0 0 la_oenb[53]
port 475 nsew signal input
flabel metal2 s 319690 -960 319802 480 0 FreeSans 448 90 0 0 la_oenb[54]
port 476 nsew signal input
flabel metal2 s 323278 -960 323390 480 0 FreeSans 448 90 0 0 la_oenb[55]
port 477 nsew signal input
flabel metal2 s 326774 -960 326886 480 0 FreeSans 448 90 0 0 la_oenb[56]
port 478 nsew signal input
flabel metal2 s 330362 -960 330474 480 0 FreeSans 448 90 0 0 la_oenb[57]
port 479 nsew signal input
flabel metal2 s 333858 -960 333970 480 0 FreeSans 448 90 0 0 la_oenb[58]
port 480 nsew signal input
flabel metal2 s 337446 -960 337558 480 0 FreeSans 448 90 0 0 la_oenb[59]
port 481 nsew signal input
flabel metal2 s 145902 -960 146014 480 0 FreeSans 448 90 0 0 la_oenb[5]
port 482 nsew signal input
flabel metal2 s 340942 -960 341054 480 0 FreeSans 448 90 0 0 la_oenb[60]
port 483 nsew signal input
flabel metal2 s 344530 -960 344642 480 0 FreeSans 448 90 0 0 la_oenb[61]
port 484 nsew signal input
flabel metal2 s 348026 -960 348138 480 0 FreeSans 448 90 0 0 la_oenb[62]
port 485 nsew signal input
flabel metal2 s 351614 -960 351726 480 0 FreeSans 448 90 0 0 la_oenb[63]
port 486 nsew signal input
flabel metal2 s 355202 -960 355314 480 0 FreeSans 448 90 0 0 la_oenb[64]
port 487 nsew signal input
flabel metal2 s 358698 -960 358810 480 0 FreeSans 448 90 0 0 la_oenb[65]
port 488 nsew signal input
flabel metal2 s 362286 -960 362398 480 0 FreeSans 448 90 0 0 la_oenb[66]
port 489 nsew signal input
flabel metal2 s 365782 -960 365894 480 0 FreeSans 448 90 0 0 la_oenb[67]
port 490 nsew signal input
flabel metal2 s 369370 -960 369482 480 0 FreeSans 448 90 0 0 la_oenb[68]
port 491 nsew signal input
flabel metal2 s 372866 -960 372978 480 0 FreeSans 448 90 0 0 la_oenb[69]
port 492 nsew signal input
flabel metal2 s 149490 -960 149602 480 0 FreeSans 448 90 0 0 la_oenb[6]
port 493 nsew signal input
flabel metal2 s 376454 -960 376566 480 0 FreeSans 448 90 0 0 la_oenb[70]
port 494 nsew signal input
flabel metal2 s 379950 -960 380062 480 0 FreeSans 448 90 0 0 la_oenb[71]
port 495 nsew signal input
flabel metal2 s 383538 -960 383650 480 0 FreeSans 448 90 0 0 la_oenb[72]
port 496 nsew signal input
flabel metal2 s 387126 -960 387238 480 0 FreeSans 448 90 0 0 la_oenb[73]
port 497 nsew signal input
flabel metal2 s 390622 -960 390734 480 0 FreeSans 448 90 0 0 la_oenb[74]
port 498 nsew signal input
flabel metal2 s 394210 -960 394322 480 0 FreeSans 448 90 0 0 la_oenb[75]
port 499 nsew signal input
flabel metal2 s 397706 -960 397818 480 0 FreeSans 448 90 0 0 la_oenb[76]
port 500 nsew signal input
flabel metal2 s 401294 -960 401406 480 0 FreeSans 448 90 0 0 la_oenb[77]
port 501 nsew signal input
flabel metal2 s 404790 -960 404902 480 0 FreeSans 448 90 0 0 la_oenb[78]
port 502 nsew signal input
flabel metal2 s 408378 -960 408490 480 0 FreeSans 448 90 0 0 la_oenb[79]
port 503 nsew signal input
flabel metal2 s 152986 -960 153098 480 0 FreeSans 448 90 0 0 la_oenb[7]
port 504 nsew signal input
flabel metal2 s 411874 -960 411986 480 0 FreeSans 448 90 0 0 la_oenb[80]
port 505 nsew signal input
flabel metal2 s 415462 -960 415574 480 0 FreeSans 448 90 0 0 la_oenb[81]
port 506 nsew signal input
flabel metal2 s 418958 -960 419070 480 0 FreeSans 448 90 0 0 la_oenb[82]
port 507 nsew signal input
flabel metal2 s 422546 -960 422658 480 0 FreeSans 448 90 0 0 la_oenb[83]
port 508 nsew signal input
flabel metal2 s 426134 -960 426246 480 0 FreeSans 448 90 0 0 la_oenb[84]
port 509 nsew signal input
flabel metal2 s 429630 -960 429742 480 0 FreeSans 448 90 0 0 la_oenb[85]
port 510 nsew signal input
flabel metal2 s 433218 -960 433330 480 0 FreeSans 448 90 0 0 la_oenb[86]
port 511 nsew signal input
flabel metal2 s 436714 -960 436826 480 0 FreeSans 448 90 0 0 la_oenb[87]
port 512 nsew signal input
flabel metal2 s 440302 -960 440414 480 0 FreeSans 448 90 0 0 la_oenb[88]
port 513 nsew signal input
flabel metal2 s 443798 -960 443910 480 0 FreeSans 448 90 0 0 la_oenb[89]
port 514 nsew signal input
flabel metal2 s 156574 -960 156686 480 0 FreeSans 448 90 0 0 la_oenb[8]
port 515 nsew signal input
flabel metal2 s 447386 -960 447498 480 0 FreeSans 448 90 0 0 la_oenb[90]
port 516 nsew signal input
flabel metal2 s 450882 -960 450994 480 0 FreeSans 448 90 0 0 la_oenb[91]
port 517 nsew signal input
flabel metal2 s 454470 -960 454582 480 0 FreeSans 448 90 0 0 la_oenb[92]
port 518 nsew signal input
flabel metal2 s 458058 -960 458170 480 0 FreeSans 448 90 0 0 la_oenb[93]
port 519 nsew signal input
flabel metal2 s 461554 -960 461666 480 0 FreeSans 448 90 0 0 la_oenb[94]
port 520 nsew signal input
flabel metal2 s 465142 -960 465254 480 0 FreeSans 448 90 0 0 la_oenb[95]
port 521 nsew signal input
flabel metal2 s 468638 -960 468750 480 0 FreeSans 448 90 0 0 la_oenb[96]
port 522 nsew signal input
flabel metal2 s 472226 -960 472338 480 0 FreeSans 448 90 0 0 la_oenb[97]
port 523 nsew signal input
flabel metal2 s 475722 -960 475834 480 0 FreeSans 448 90 0 0 la_oenb[98]
port 524 nsew signal input
flabel metal2 s 479310 -960 479422 480 0 FreeSans 448 90 0 0 la_oenb[99]
port 525 nsew signal input
flabel metal2 s 160070 -960 160182 480 0 FreeSans 448 90 0 0 la_oenb[9]
port 526 nsew signal input
flabel metal2 s 579774 -960 579886 480 0 FreeSans 448 90 0 0 user_clock2
port 527 nsew signal input
flabel metal2 s 580970 -960 581082 480 0 FreeSans 448 90 0 0 user_irq[0]
port 528 nsew signal tristate
flabel metal2 s 582166 -960 582278 480 0 FreeSans 448 90 0 0 user_irq[1]
port 529 nsew signal tristate
flabel metal2 s 583362 -960 583474 480 0 FreeSans 448 90 0 0 user_irq[2]
port 530 nsew signal tristate
flabel metal4 s -2006 -934 -1386 704870 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -2006 -934 585930 -314 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -2006 704250 585930 704870 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 585310 -934 585930 704870 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 1794 -7654 2414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 37794 -7654 38414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 73794 -7654 74414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 109794 -7654 110414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 145794 -7654 146414 78000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 145794 142000 146414 198000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 145794 262000 146414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 181794 -7654 182414 78000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 181794 142000 182414 198000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 181794 262000 182414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 217794 -7654 218414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 253794 -7654 254414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 289794 -7654 290414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 325794 -7654 326414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 361794 -7654 362414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 397794 -7654 398414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 433794 -7654 434414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 469794 -7654 470414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 505794 -7654 506414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 541794 -7654 542414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 577794 -7654 578414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 2866 592650 3486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 38866 592650 39486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 74866 592650 75486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 110866 592650 111486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 146866 592650 147486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 182866 592650 183486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 218866 592650 219486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 254866 592650 255486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 290866 592650 291486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 326866 592650 327486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 362866 592650 363486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 398866 592650 399486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 434866 592650 435486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 470866 592650 471486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 506866 592650 507486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 542866 592650 543486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 578866 592650 579486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 614866 592650 615486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 650866 592650 651486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 686866 592650 687486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s -3926 -2854 -3306 706790 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -3926 -2854 587850 -2234 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -3926 706170 587850 706790 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 587230 -2854 587850 706790 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 10794 -7654 11414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 46794 -7654 47414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 82794 -7654 83414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 118794 -7654 119414 78000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 118794 142000 119414 198000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 118794 262000 119414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 154794 -7654 155414 78000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 154794 142000 155414 198000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 154794 262000 155414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 190794 -7654 191414 78000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 190794 142000 191414 198000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 190794 262000 191414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 226794 -7654 227414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 262794 -7654 263414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 298794 -7654 299414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 334794 -7654 335414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 370794 -7654 371414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 406794 -7654 407414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 442794 -7654 443414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 478794 -7654 479414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 514794 -7654 515414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 550794 -7654 551414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 11866 592650 12486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 47866 592650 48486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 83866 592650 84486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 119866 592650 120486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 155866 592650 156486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 191866 592650 192486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 227866 592650 228486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 263866 592650 264486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 299866 592650 300486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 335866 592650 336486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 371866 592650 372486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 407866 592650 408486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 443866 592650 444486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 479866 592650 480486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 515866 592650 516486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 551866 592650 552486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 587866 592650 588486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 623866 592650 624486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 659866 592650 660486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 695866 592650 696486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s -5846 -4774 -5226 708710 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -5846 -4774 589770 -4154 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -5846 708090 589770 708710 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 589150 -4774 589770 708710 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 19794 -7654 20414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 55794 -7654 56414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 91794 -7654 92414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 127794 -7654 128414 78000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 127794 262000 128414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 163794 -7654 164414 78000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 163794 262000 164414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 199794 -7654 200414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 235794 -7654 236414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 271794 -7654 272414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 307794 -7654 308414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 343794 -7654 344414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 379794 -7654 380414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 415794 -7654 416414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 451794 -7654 452414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 487794 -7654 488414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 523794 -7654 524414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 559794 -7654 560414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 20866 592650 21486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 56866 592650 57486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 92866 592650 93486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 128866 592650 129486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 164866 592650 165486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 200866 592650 201486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 236866 592650 237486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 272866 592650 273486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 308866 592650 309486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 344866 592650 345486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 380866 592650 381486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 416866 592650 417486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 452866 592650 453486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 488866 592650 489486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 524866 592650 525486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 560866 592650 561486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 596866 592650 597486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 632866 592650 633486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 668866 592650 669486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s -7766 -6694 -7146 710630 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -7766 -6694 591690 -6074 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -7766 710010 591690 710630 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 591070 -6694 591690 710630 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 28794 -7654 29414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 64794 -7654 65414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 100794 -7654 101414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 136794 -7654 137414 78000 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 136794 262000 137414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 172794 -7654 173414 78000 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 172794 262000 173414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 208794 -7654 209414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 244794 -7654 245414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 280794 -7654 281414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 316794 -7654 317414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 352794 -7654 353414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 388794 -7654 389414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 424794 -7654 425414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 460794 -7654 461414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 496794 -7654 497414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 532794 -7654 533414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 568794 -7654 569414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 29866 592650 30486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 65866 592650 66486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 101866 592650 102486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 137866 592650 138486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 173866 592650 174486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 209866 592650 210486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 245866 592650 246486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 281866 592650 282486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 317866 592650 318486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 353866 592650 354486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 389866 592650 390486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 425866 592650 426486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 461866 592650 462486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 497866 592650 498486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 533866 592650 534486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 569866 592650 570486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 605866 592650 606486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 641866 592650 642486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 677866 592650 678486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s -6806 -5734 -6186 709670 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -6806 -5734 590730 -5114 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -6806 709050 590730 709670 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 590110 -5734 590730 709670 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 24294 -7654 24914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 60294 -7654 60914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 96294 -7654 96914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 132294 -7654 132914 78000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 132294 262000 132914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 168294 -7654 168914 78000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 168294 262000 168914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 204294 -7654 204914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 240294 -7654 240914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 276294 -7654 276914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 312294 -7654 312914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 348294 -7654 348914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 384294 -7654 384914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 420294 -7654 420914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 456294 -7654 456914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 492294 -7654 492914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 528294 -7654 528914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 564294 -7654 564914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 25366 592650 25986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 61366 592650 61986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 97366 592650 97986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 133366 592650 133986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 169366 592650 169986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 205366 592650 205986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 241366 592650 241986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 277366 592650 277986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 313366 592650 313986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 349366 592650 349986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 385366 592650 385986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 421366 592650 421986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 457366 592650 457986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 493366 592650 493986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 529366 592650 529986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 565366 592650 565986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 601366 592650 601986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 637366 592650 637986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 673366 592650 673986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s -8726 -7654 -8106 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 -7654 592650 -7034 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 710970 592650 711590 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 592030 -7654 592650 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 33294 -7654 33914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 69294 -7654 69914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 105294 -7654 105914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 141294 -7654 141914 78000 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 141294 142000 141914 198000 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 141294 262000 141914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 177294 -7654 177914 78000 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 177294 142000 177914 198000 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 177294 262000 177914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 213294 -7654 213914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 249294 -7654 249914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 285294 -7654 285914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 321294 -7654 321914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 357294 -7654 357914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 393294 -7654 393914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 429294 -7654 429914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 465294 -7654 465914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 501294 -7654 501914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 537294 -7654 537914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 573294 -7654 573914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 34366 592650 34986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 70366 592650 70986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 106366 592650 106986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 142366 592650 142986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 178366 592650 178986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 214366 592650 214986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 250366 592650 250986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 286366 592650 286986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 322366 592650 322986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 358366 592650 358986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 394366 592650 394986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 430366 592650 430986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 466366 592650 466986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 502366 592650 502986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 538366 592650 538986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 574366 592650 574986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 610366 592650 610986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 646366 592650 646986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 682366 592650 682986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s -2966 -1894 -2346 705830 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -2966 -1894 586890 -1274 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -2966 705210 586890 705830 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 586270 -1894 586890 705830 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 6294 -7654 6914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 42294 -7654 42914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 78294 -7654 78914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 114294 -7654 114914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 150294 -7654 150914 78000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 150294 142000 150914 198000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 150294 262000 150914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 186294 -7654 186914 78000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 186294 142000 186914 198000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 186294 262000 186914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 222294 -7654 222914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 258294 -7654 258914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 294294 -7654 294914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 330294 -7654 330914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 366294 -7654 366914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 402294 -7654 402914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 438294 -7654 438914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 474294 -7654 474914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 510294 -7654 510914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 546294 -7654 546914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 582294 -7654 582914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 7366 592650 7986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 43366 592650 43986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 79366 592650 79986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 115366 592650 115986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 151366 592650 151986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 187366 592650 187986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 223366 592650 223986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 259366 592650 259986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 295366 592650 295986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 331366 592650 331986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 367366 592650 367986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 403366 592650 403986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 439366 592650 439986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 475366 592650 475986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 511366 592650 511986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 547366 592650 547986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 583366 592650 583986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 619366 592650 619986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 655366 592650 655986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 691366 592650 691986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s -4886 -3814 -4266 707750 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -4886 -3814 588810 -3194 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -4886 707130 588810 707750 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 588190 -3814 588810 707750 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 15294 -7654 15914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 51294 -7654 51914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 87294 -7654 87914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 123294 -7654 123914 78000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 123294 142000 123914 198000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 123294 262000 123914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 159294 -7654 159914 78000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 159294 142000 159914 198000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 159294 262000 159914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 195294 -7654 195914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 231294 -7654 231914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 267294 -7654 267914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 303294 -7654 303914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 339294 -7654 339914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 375294 -7654 375914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 411294 -7654 411914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 447294 -7654 447914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 483294 -7654 483914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 519294 -7654 519914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 555294 -7654 555914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 16366 592650 16986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 52366 592650 52986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 88366 592650 88986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 124366 592650 124986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 160366 592650 160986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 196366 592650 196986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 232366 592650 232986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 268366 592650 268986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 304366 592650 304986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 340366 592650 340986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 376366 592650 376986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 412366 592650 412986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 448366 592650 448986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 484366 592650 484986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 520366 592650 520986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 556366 592650 556986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 592366 592650 592986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 628366 592650 628986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 664366 592650 664986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 700366 592650 700986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal2 s 542 -960 654 480 0 FreeSans 448 90 0 0 wb_clk_i
port 539 nsew signal input
flabel metal2 s 1646 -960 1758 480 0 FreeSans 448 90 0 0 wb_rst_i
port 540 nsew signal input
flabel metal2 s 2842 -960 2954 480 0 FreeSans 448 90 0 0 wbs_ack_o
port 541 nsew signal tristate
flabel metal2 s 7626 -960 7738 480 0 FreeSans 448 90 0 0 wbs_adr_i[0]
port 542 nsew signal input
flabel metal2 s 47830 -960 47942 480 0 FreeSans 448 90 0 0 wbs_adr_i[10]
port 543 nsew signal input
flabel metal2 s 51326 -960 51438 480 0 FreeSans 448 90 0 0 wbs_adr_i[11]
port 544 nsew signal input
flabel metal2 s 54914 -960 55026 480 0 FreeSans 448 90 0 0 wbs_adr_i[12]
port 545 nsew signal input
flabel metal2 s 58410 -960 58522 480 0 FreeSans 448 90 0 0 wbs_adr_i[13]
port 546 nsew signal input
flabel metal2 s 61998 -960 62110 480 0 FreeSans 448 90 0 0 wbs_adr_i[14]
port 547 nsew signal input
flabel metal2 s 65494 -960 65606 480 0 FreeSans 448 90 0 0 wbs_adr_i[15]
port 548 nsew signal input
flabel metal2 s 69082 -960 69194 480 0 FreeSans 448 90 0 0 wbs_adr_i[16]
port 549 nsew signal input
flabel metal2 s 72578 -960 72690 480 0 FreeSans 448 90 0 0 wbs_adr_i[17]
port 550 nsew signal input
flabel metal2 s 76166 -960 76278 480 0 FreeSans 448 90 0 0 wbs_adr_i[18]
port 551 nsew signal input
flabel metal2 s 79662 -960 79774 480 0 FreeSans 448 90 0 0 wbs_adr_i[19]
port 552 nsew signal input
flabel metal2 s 12318 -960 12430 480 0 FreeSans 448 90 0 0 wbs_adr_i[1]
port 553 nsew signal input
flabel metal2 s 83250 -960 83362 480 0 FreeSans 448 90 0 0 wbs_adr_i[20]
port 554 nsew signal input
flabel metal2 s 86838 -960 86950 480 0 FreeSans 448 90 0 0 wbs_adr_i[21]
port 555 nsew signal input
flabel metal2 s 90334 -960 90446 480 0 FreeSans 448 90 0 0 wbs_adr_i[22]
port 556 nsew signal input
flabel metal2 s 93922 -960 94034 480 0 FreeSans 448 90 0 0 wbs_adr_i[23]
port 557 nsew signal input
flabel metal2 s 97418 -960 97530 480 0 FreeSans 448 90 0 0 wbs_adr_i[24]
port 558 nsew signal input
flabel metal2 s 101006 -960 101118 480 0 FreeSans 448 90 0 0 wbs_adr_i[25]
port 559 nsew signal input
flabel metal2 s 104502 -960 104614 480 0 FreeSans 448 90 0 0 wbs_adr_i[26]
port 560 nsew signal input
flabel metal2 s 108090 -960 108202 480 0 FreeSans 448 90 0 0 wbs_adr_i[27]
port 561 nsew signal input
flabel metal2 s 111586 -960 111698 480 0 FreeSans 448 90 0 0 wbs_adr_i[28]
port 562 nsew signal input
flabel metal2 s 115174 -960 115286 480 0 FreeSans 448 90 0 0 wbs_adr_i[29]
port 563 nsew signal input
flabel metal2 s 17010 -960 17122 480 0 FreeSans 448 90 0 0 wbs_adr_i[2]
port 564 nsew signal input
flabel metal2 s 118762 -960 118874 480 0 FreeSans 448 90 0 0 wbs_adr_i[30]
port 565 nsew signal input
flabel metal2 s 122258 -960 122370 480 0 FreeSans 448 90 0 0 wbs_adr_i[31]
port 566 nsew signal input
flabel metal2 s 21794 -960 21906 480 0 FreeSans 448 90 0 0 wbs_adr_i[3]
port 567 nsew signal input
flabel metal2 s 26486 -960 26598 480 0 FreeSans 448 90 0 0 wbs_adr_i[4]
port 568 nsew signal input
flabel metal2 s 30074 -960 30186 480 0 FreeSans 448 90 0 0 wbs_adr_i[5]
port 569 nsew signal input
flabel metal2 s 33570 -960 33682 480 0 FreeSans 448 90 0 0 wbs_adr_i[6]
port 570 nsew signal input
flabel metal2 s 37158 -960 37270 480 0 FreeSans 448 90 0 0 wbs_adr_i[7]
port 571 nsew signal input
flabel metal2 s 40654 -960 40766 480 0 FreeSans 448 90 0 0 wbs_adr_i[8]
port 572 nsew signal input
flabel metal2 s 44242 -960 44354 480 0 FreeSans 448 90 0 0 wbs_adr_i[9]
port 573 nsew signal input
flabel metal2 s 4038 -960 4150 480 0 FreeSans 448 90 0 0 wbs_cyc_i
port 574 nsew signal input
flabel metal2 s 8730 -960 8842 480 0 FreeSans 448 90 0 0 wbs_dat_i[0]
port 575 nsew signal input
flabel metal2 s 48934 -960 49046 480 0 FreeSans 448 90 0 0 wbs_dat_i[10]
port 576 nsew signal input
flabel metal2 s 52522 -960 52634 480 0 FreeSans 448 90 0 0 wbs_dat_i[11]
port 577 nsew signal input
flabel metal2 s 56018 -960 56130 480 0 FreeSans 448 90 0 0 wbs_dat_i[12]
port 578 nsew signal input
flabel metal2 s 59606 -960 59718 480 0 FreeSans 448 90 0 0 wbs_dat_i[13]
port 579 nsew signal input
flabel metal2 s 63194 -960 63306 480 0 FreeSans 448 90 0 0 wbs_dat_i[14]
port 580 nsew signal input
flabel metal2 s 66690 -960 66802 480 0 FreeSans 448 90 0 0 wbs_dat_i[15]
port 581 nsew signal input
flabel metal2 s 70278 -960 70390 480 0 FreeSans 448 90 0 0 wbs_dat_i[16]
port 582 nsew signal input
flabel metal2 s 73774 -960 73886 480 0 FreeSans 448 90 0 0 wbs_dat_i[17]
port 583 nsew signal input
flabel metal2 s 77362 -960 77474 480 0 FreeSans 448 90 0 0 wbs_dat_i[18]
port 584 nsew signal input
flabel metal2 s 80858 -960 80970 480 0 FreeSans 448 90 0 0 wbs_dat_i[19]
port 585 nsew signal input
flabel metal2 s 13514 -960 13626 480 0 FreeSans 448 90 0 0 wbs_dat_i[1]
port 586 nsew signal input
flabel metal2 s 84446 -960 84558 480 0 FreeSans 448 90 0 0 wbs_dat_i[20]
port 587 nsew signal input
flabel metal2 s 87942 -960 88054 480 0 FreeSans 448 90 0 0 wbs_dat_i[21]
port 588 nsew signal input
flabel metal2 s 91530 -960 91642 480 0 FreeSans 448 90 0 0 wbs_dat_i[22]
port 589 nsew signal input
flabel metal2 s 95118 -960 95230 480 0 FreeSans 448 90 0 0 wbs_dat_i[23]
port 590 nsew signal input
flabel metal2 s 98614 -960 98726 480 0 FreeSans 448 90 0 0 wbs_dat_i[24]
port 591 nsew signal input
flabel metal2 s 102202 -960 102314 480 0 FreeSans 448 90 0 0 wbs_dat_i[25]
port 592 nsew signal input
flabel metal2 s 105698 -960 105810 480 0 FreeSans 448 90 0 0 wbs_dat_i[26]
port 593 nsew signal input
flabel metal2 s 109286 -960 109398 480 0 FreeSans 448 90 0 0 wbs_dat_i[27]
port 594 nsew signal input
flabel metal2 s 112782 -960 112894 480 0 FreeSans 448 90 0 0 wbs_dat_i[28]
port 595 nsew signal input
flabel metal2 s 116370 -960 116482 480 0 FreeSans 448 90 0 0 wbs_dat_i[29]
port 596 nsew signal input
flabel metal2 s 18206 -960 18318 480 0 FreeSans 448 90 0 0 wbs_dat_i[2]
port 597 nsew signal input
flabel metal2 s 119866 -960 119978 480 0 FreeSans 448 90 0 0 wbs_dat_i[30]
port 598 nsew signal input
flabel metal2 s 123454 -960 123566 480 0 FreeSans 448 90 0 0 wbs_dat_i[31]
port 599 nsew signal input
flabel metal2 s 22990 -960 23102 480 0 FreeSans 448 90 0 0 wbs_dat_i[3]
port 600 nsew signal input
flabel metal2 s 27682 -960 27794 480 0 FreeSans 448 90 0 0 wbs_dat_i[4]
port 601 nsew signal input
flabel metal2 s 31270 -960 31382 480 0 FreeSans 448 90 0 0 wbs_dat_i[5]
port 602 nsew signal input
flabel metal2 s 34766 -960 34878 480 0 FreeSans 448 90 0 0 wbs_dat_i[6]
port 603 nsew signal input
flabel metal2 s 38354 -960 38466 480 0 FreeSans 448 90 0 0 wbs_dat_i[7]
port 604 nsew signal input
flabel metal2 s 41850 -960 41962 480 0 FreeSans 448 90 0 0 wbs_dat_i[8]
port 605 nsew signal input
flabel metal2 s 45438 -960 45550 480 0 FreeSans 448 90 0 0 wbs_dat_i[9]
port 606 nsew signal input
flabel metal2 s 9926 -960 10038 480 0 FreeSans 448 90 0 0 wbs_dat_o[0]
port 607 nsew signal tristate
flabel metal2 s 50130 -960 50242 480 0 FreeSans 448 90 0 0 wbs_dat_o[10]
port 608 nsew signal tristate
flabel metal2 s 53718 -960 53830 480 0 FreeSans 448 90 0 0 wbs_dat_o[11]
port 609 nsew signal tristate
flabel metal2 s 57214 -960 57326 480 0 FreeSans 448 90 0 0 wbs_dat_o[12]
port 610 nsew signal tristate
flabel metal2 s 60802 -960 60914 480 0 FreeSans 448 90 0 0 wbs_dat_o[13]
port 611 nsew signal tristate
flabel metal2 s 64298 -960 64410 480 0 FreeSans 448 90 0 0 wbs_dat_o[14]
port 612 nsew signal tristate
flabel metal2 s 67886 -960 67998 480 0 FreeSans 448 90 0 0 wbs_dat_o[15]
port 613 nsew signal tristate
flabel metal2 s 71474 -960 71586 480 0 FreeSans 448 90 0 0 wbs_dat_o[16]
port 614 nsew signal tristate
flabel metal2 s 74970 -960 75082 480 0 FreeSans 448 90 0 0 wbs_dat_o[17]
port 615 nsew signal tristate
flabel metal2 s 78558 -960 78670 480 0 FreeSans 448 90 0 0 wbs_dat_o[18]
port 616 nsew signal tristate
flabel metal2 s 82054 -960 82166 480 0 FreeSans 448 90 0 0 wbs_dat_o[19]
port 617 nsew signal tristate
flabel metal2 s 14710 -960 14822 480 0 FreeSans 448 90 0 0 wbs_dat_o[1]
port 618 nsew signal tristate
flabel metal2 s 85642 -960 85754 480 0 FreeSans 448 90 0 0 wbs_dat_o[20]
port 619 nsew signal tristate
flabel metal2 s 89138 -960 89250 480 0 FreeSans 448 90 0 0 wbs_dat_o[21]
port 620 nsew signal tristate
flabel metal2 s 92726 -960 92838 480 0 FreeSans 448 90 0 0 wbs_dat_o[22]
port 621 nsew signal tristate
flabel metal2 s 96222 -960 96334 480 0 FreeSans 448 90 0 0 wbs_dat_o[23]
port 622 nsew signal tristate
flabel metal2 s 99810 -960 99922 480 0 FreeSans 448 90 0 0 wbs_dat_o[24]
port 623 nsew signal tristate
flabel metal2 s 103306 -960 103418 480 0 FreeSans 448 90 0 0 wbs_dat_o[25]
port 624 nsew signal tristate
flabel metal2 s 106894 -960 107006 480 0 FreeSans 448 90 0 0 wbs_dat_o[26]
port 625 nsew signal tristate
flabel metal2 s 110482 -960 110594 480 0 FreeSans 448 90 0 0 wbs_dat_o[27]
port 626 nsew signal tristate
flabel metal2 s 113978 -960 114090 480 0 FreeSans 448 90 0 0 wbs_dat_o[28]
port 627 nsew signal tristate
flabel metal2 s 117566 -960 117678 480 0 FreeSans 448 90 0 0 wbs_dat_o[29]
port 628 nsew signal tristate
flabel metal2 s 19402 -960 19514 480 0 FreeSans 448 90 0 0 wbs_dat_o[2]
port 629 nsew signal tristate
flabel metal2 s 121062 -960 121174 480 0 FreeSans 448 90 0 0 wbs_dat_o[30]
port 630 nsew signal tristate
flabel metal2 s 124650 -960 124762 480 0 FreeSans 448 90 0 0 wbs_dat_o[31]
port 631 nsew signal tristate
flabel metal2 s 24186 -960 24298 480 0 FreeSans 448 90 0 0 wbs_dat_o[3]
port 632 nsew signal tristate
flabel metal2 s 28878 -960 28990 480 0 FreeSans 448 90 0 0 wbs_dat_o[4]
port 633 nsew signal tristate
flabel metal2 s 32374 -960 32486 480 0 FreeSans 448 90 0 0 wbs_dat_o[5]
port 634 nsew signal tristate
flabel metal2 s 35962 -960 36074 480 0 FreeSans 448 90 0 0 wbs_dat_o[6]
port 635 nsew signal tristate
flabel metal2 s 39550 -960 39662 480 0 FreeSans 448 90 0 0 wbs_dat_o[7]
port 636 nsew signal tristate
flabel metal2 s 43046 -960 43158 480 0 FreeSans 448 90 0 0 wbs_dat_o[8]
port 637 nsew signal tristate
flabel metal2 s 46634 -960 46746 480 0 FreeSans 448 90 0 0 wbs_dat_o[9]
port 638 nsew signal tristate
flabel metal2 s 11122 -960 11234 480 0 FreeSans 448 90 0 0 wbs_sel_i[0]
port 639 nsew signal input
flabel metal2 s 15906 -960 16018 480 0 FreeSans 448 90 0 0 wbs_sel_i[1]
port 640 nsew signal input
flabel metal2 s 20598 -960 20710 480 0 FreeSans 448 90 0 0 wbs_sel_i[2]
port 641 nsew signal input
flabel metal2 s 25290 -960 25402 480 0 FreeSans 448 90 0 0 wbs_sel_i[3]
port 642 nsew signal input
flabel metal2 s 5234 -960 5346 480 0 FreeSans 448 90 0 0 wbs_stb_i
port 643 nsew signal input
flabel metal2 s 6430 -960 6542 480 0 FreeSans 448 90 0 0 wbs_we_i
port 644 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
