magic
tech sky130B
magscale 1 2
timestamp 1662148784
<< viali >>
rect 3893 17289 3927 17323
rect 11713 17289 11747 17323
rect 18153 17289 18187 17323
rect 25329 17289 25363 17323
rect 32597 17289 32631 17323
rect 34069 17289 34103 17323
rect 1409 17153 1443 17187
rect 4077 17153 4111 17187
rect 11529 17153 11563 17187
rect 18337 17153 18371 17187
rect 25513 17153 25547 17187
rect 32413 17153 32447 17187
rect 33885 17153 33919 17187
rect 1685 17085 1719 17119
rect 33333 16949 33367 16983
rect 1409 16745 1443 16779
rect 6561 16541 6595 16575
rect 33885 16541 33919 16575
rect 6745 16405 6779 16439
rect 34069 16405 34103 16439
rect 8493 16201 8527 16235
rect 21833 16201 21867 16235
rect 28181 16201 28215 16235
rect 7021 16133 7055 16167
rect 22293 16133 22327 16167
rect 28273 16133 28307 16167
rect 15209 16065 15243 16099
rect 21005 16065 21039 16099
rect 22201 16065 22235 16099
rect 29285 16065 29319 16099
rect 6745 15997 6779 16031
rect 8953 15997 8987 16031
rect 22385 15997 22419 16031
rect 27997 15997 28031 16031
rect 28641 15929 28675 15963
rect 15025 15861 15059 15895
rect 20821 15861 20855 15895
rect 29101 15861 29135 15895
rect 6469 15657 6503 15691
rect 7941 15657 7975 15691
rect 13461 15657 13495 15691
rect 15853 15657 15887 15691
rect 22109 15657 22143 15691
rect 7021 15521 7055 15555
rect 14105 15521 14139 15555
rect 14381 15521 14415 15555
rect 20637 15521 20671 15555
rect 8033 15453 8067 15487
rect 20361 15453 20395 15487
rect 6929 15385 6963 15419
rect 6837 15317 6871 15351
rect 14381 15113 14415 15147
rect 20545 15113 20579 15147
rect 21005 15113 21039 15147
rect 29929 15113 29963 15147
rect 14289 14977 14323 15011
rect 15117 14977 15151 15011
rect 20913 14977 20947 15011
rect 21189 14909 21223 14943
rect 28181 14909 28215 14943
rect 28457 14909 28491 14943
rect 15209 14841 15243 14875
rect 7297 14773 7331 14807
rect 21925 14773 21959 14807
rect 6653 14433 6687 14467
rect 6469 14365 6503 14399
rect 6377 14297 6411 14331
rect 6009 14229 6043 14263
rect 7297 14229 7331 14263
rect 29837 14025 29871 14059
rect 5181 13889 5215 13923
rect 28089 13889 28123 13923
rect 33885 13889 33919 13923
rect 6837 13821 6871 13855
rect 28365 13821 28399 13855
rect 4997 13685 5031 13719
rect 34069 13685 34103 13719
rect 5917 13481 5951 13515
rect 6469 13481 6503 13515
rect 20177 13481 20211 13515
rect 21741 13481 21775 13515
rect 29745 13481 29779 13515
rect 4169 13345 4203 13379
rect 31493 13345 31527 13379
rect 31585 13345 31619 13379
rect 14289 13277 14323 13311
rect 21649 13277 21683 13311
rect 22293 13277 22327 13311
rect 29929 13277 29963 13311
rect 31401 13277 31435 13311
rect 4445 13209 4479 13243
rect 14197 13141 14231 13175
rect 20729 13141 20763 13175
rect 30481 13141 30515 13175
rect 31033 13141 31067 13175
rect 6469 12937 6503 12971
rect 12909 12937 12943 12971
rect 20913 12937 20947 12971
rect 28549 12937 28583 12971
rect 6561 12801 6595 12835
rect 15209 12801 15243 12835
rect 19809 12801 19843 12835
rect 28457 12801 28491 12835
rect 29101 12801 29135 12835
rect 1409 12733 1443 12767
rect 1685 12733 1719 12767
rect 14933 12733 14967 12767
rect 20729 12733 20763 12767
rect 21097 12733 21131 12767
rect 19625 12665 19659 12699
rect 13461 12597 13495 12631
rect 21097 12597 21131 12631
rect 21925 12597 21959 12631
rect 1409 12393 1443 12427
rect 6653 12393 6687 12427
rect 20729 12393 20763 12427
rect 21281 12257 21315 12291
rect 6837 12189 6871 12223
rect 21097 12121 21131 12155
rect 6009 12053 6043 12087
rect 20269 12053 20303 12087
rect 21189 12053 21223 12087
rect 6377 11713 6411 11747
rect 33885 11713 33919 11747
rect 6837 11577 6871 11611
rect 20545 11577 20579 11611
rect 5733 11509 5767 11543
rect 6469 11509 6503 11543
rect 34069 11509 34103 11543
rect 6101 11305 6135 11339
rect 11253 11305 11287 11339
rect 27905 11305 27939 11339
rect 20453 11237 20487 11271
rect 31033 11237 31067 11271
rect 11805 11169 11839 11203
rect 13553 11169 13587 11203
rect 19441 11169 19475 11203
rect 31585 11169 31619 11203
rect 19717 11101 19751 11135
rect 28457 11101 28491 11135
rect 29929 11101 29963 11135
rect 13277 11033 13311 11067
rect 28549 11033 28583 11067
rect 30481 11033 30515 11067
rect 31401 11033 31435 11067
rect 31493 11033 31527 11067
rect 29745 10965 29779 10999
rect 12725 10761 12759 10795
rect 29745 10761 29779 10795
rect 4445 10625 4479 10659
rect 12817 10625 12851 10659
rect 13277 10625 13311 10659
rect 18245 10625 18279 10659
rect 19993 10625 20027 10659
rect 27997 10625 28031 10659
rect 28273 10557 28307 10591
rect 3893 10421 3927 10455
rect 4629 10421 4663 10455
rect 10885 10217 10919 10251
rect 13093 10217 13127 10251
rect 20269 10217 20303 10251
rect 17693 10081 17727 10115
rect 21281 10081 21315 10115
rect 4905 10013 4939 10047
rect 5549 10013 5583 10047
rect 12173 10013 12207 10047
rect 13277 10013 13311 10047
rect 13553 10013 13587 10047
rect 21005 10013 21039 10047
rect 15945 9945 15979 9979
rect 4997 9877 5031 9911
rect 13461 9877 13495 9911
rect 15393 9877 15427 9911
rect 13737 9673 13771 9707
rect 6469 9605 6503 9639
rect 13645 9537 13679 9571
rect 13829 9537 13863 9571
rect 3985 9469 4019 9503
rect 4261 9469 4295 9503
rect 5733 9333 5767 9367
rect 28089 9129 28123 9163
rect 12725 8993 12759 9027
rect 21741 8993 21775 9027
rect 12357 8925 12391 8959
rect 12633 8925 12667 8959
rect 22017 8925 22051 8959
rect 22845 8925 22879 8959
rect 28641 8925 28675 8959
rect 33885 8925 33919 8959
rect 28733 8789 28767 8823
rect 34069 8789 34103 8823
rect 14289 8585 14323 8619
rect 11805 8449 11839 8483
rect 14197 8449 14231 8483
rect 14381 8449 14415 8483
rect 27813 8449 27847 8483
rect 12081 8381 12115 8415
rect 28089 8381 28123 8415
rect 29561 8313 29595 8347
rect 1593 8041 1627 8075
rect 10885 8041 10919 8075
rect 11805 8041 11839 8075
rect 27445 8041 27479 8075
rect 32413 8041 32447 8075
rect 19993 7905 20027 7939
rect 21281 7905 21315 7939
rect 1409 7837 1443 7871
rect 10793 7837 10827 7871
rect 10977 7837 11011 7871
rect 11437 7837 11471 7871
rect 11713 7837 11747 7871
rect 19717 7837 19751 7871
rect 19809 7837 19843 7871
rect 21189 7837 21223 7871
rect 22109 7837 22143 7871
rect 27261 7837 27295 7871
rect 31401 7837 31435 7871
rect 31677 7837 31711 7871
rect 19993 7769 20027 7803
rect 21925 7769 21959 7803
rect 11989 7701 12023 7735
rect 22293 7701 22327 7735
rect 1409 7497 1443 7531
rect 12173 7497 12207 7531
rect 26433 7497 26467 7531
rect 27353 7497 27387 7531
rect 27721 7497 27755 7531
rect 3617 7361 3651 7395
rect 12357 7361 12391 7395
rect 12449 7361 12483 7395
rect 12725 7361 12759 7395
rect 14565 7361 14599 7395
rect 14749 7361 14783 7395
rect 3893 7293 3927 7327
rect 27077 7293 27111 7327
rect 27261 7293 27295 7327
rect 12633 7225 12667 7259
rect 5365 7157 5399 7191
rect 14657 7157 14691 7191
rect 11989 6953 12023 6987
rect 20821 6953 20855 6987
rect 11897 6885 11931 6919
rect 21005 6885 21039 6919
rect 4721 6817 4755 6851
rect 12127 6817 12161 6851
rect 20085 6817 20119 6851
rect 4629 6749 4663 6783
rect 11805 6749 11839 6783
rect 12265 6749 12299 6783
rect 19993 6749 20027 6783
rect 20177 6749 20211 6783
rect 21465 6749 21499 6783
rect 21649 6749 21683 6783
rect 30389 6749 30423 6783
rect 33885 6749 33919 6783
rect 20637 6681 20671 6715
rect 5549 6613 5583 6647
rect 20837 6613 20871 6647
rect 21649 6613 21683 6647
rect 30573 6613 30607 6647
rect 34069 6613 34103 6647
rect 4905 6409 4939 6443
rect 12265 6409 12299 6443
rect 33149 6409 33183 6443
rect 12449 6273 12483 6307
rect 28089 6273 28123 6307
rect 32413 6273 32447 6307
rect 12633 6205 12667 6239
rect 32137 6205 32171 6239
rect 28273 6069 28307 6103
rect 11713 5729 11747 5763
rect 4721 5661 4755 5695
rect 5181 5661 5215 5695
rect 6193 5661 6227 5695
rect 11437 5661 11471 5695
rect 6009 5593 6043 5627
rect 4629 5525 4663 5559
rect 6377 5525 6411 5559
rect 12357 5321 12391 5355
rect 19809 5253 19843 5287
rect 20361 5253 20395 5287
rect 12265 5185 12299 5219
rect 12449 5185 12483 5219
rect 19625 5185 19659 5219
rect 20545 5185 20579 5219
rect 22937 5185 22971 5219
rect 23213 5185 23247 5219
rect 23949 4981 23983 5015
rect 19625 4777 19659 4811
rect 12725 4641 12759 4675
rect 29561 4641 29595 4675
rect 12357 4573 12391 4607
rect 12541 4573 12575 4607
rect 18337 4573 18371 4607
rect 18521 4573 18555 4607
rect 19257 4573 19291 4607
rect 19441 4573 19475 4607
rect 29837 4573 29871 4607
rect 6377 4505 6411 4539
rect 6469 4437 6503 4471
rect 18521 4437 18555 4471
rect 30573 4437 30607 4471
rect 11529 4097 11563 4131
rect 11713 4097 11747 4131
rect 12173 4097 12207 4131
rect 12449 4097 12483 4131
rect 12725 4097 12759 4131
rect 12817 4097 12851 4131
rect 13185 4097 13219 4131
rect 13645 4097 13679 4131
rect 33885 4097 33919 4131
rect 3525 4029 3559 4063
rect 3801 4029 3835 4063
rect 5273 4029 5307 4063
rect 12265 4029 12299 4063
rect 13737 4029 13771 4063
rect 15393 4029 15427 4063
rect 15853 4029 15887 4063
rect 5733 3961 5767 3995
rect 15669 3961 15703 3995
rect 11713 3893 11747 3927
rect 34069 3893 34103 3927
rect 12909 3689 12943 3723
rect 21741 3689 21775 3723
rect 22569 3689 22603 3723
rect 24593 3689 24627 3723
rect 29653 3689 29687 3723
rect 31585 3689 31619 3723
rect 23673 3621 23707 3655
rect 24777 3621 24811 3655
rect 5089 3553 5123 3587
rect 5549 3553 5583 3587
rect 22937 3553 22971 3587
rect 5181 3485 5215 3519
rect 12357 3485 12391 3519
rect 12725 3485 12759 3519
rect 21925 3485 21959 3519
rect 23857 3485 23891 3519
rect 28549 3485 28583 3519
rect 30389 3485 30423 3519
rect 30665 3485 30699 3519
rect 31677 3485 31711 3519
rect 12541 3417 12575 3451
rect 12633 3417 12667 3451
rect 22569 3417 22603 3451
rect 24409 3417 24443 3451
rect 22385 3349 22419 3383
rect 24609 3349 24643 3383
rect 28733 3349 28767 3383
rect 31217 3349 31251 3383
rect 12541 3145 12575 3179
rect 23765 3145 23799 3179
rect 30757 3145 30791 3179
rect 23581 3077 23615 3111
rect 12173 3009 12207 3043
rect 12357 3009 12391 3043
rect 23213 3009 23247 3043
rect 30941 3009 30975 3043
rect 1777 2805 1811 2839
rect 12357 2805 12391 2839
rect 23581 2805 23615 2839
rect 2053 2533 2087 2567
rect 4537 2533 4571 2567
rect 6837 2533 6871 2567
rect 33425 2465 33459 2499
rect 1869 2397 1903 2431
rect 4353 2397 4387 2431
rect 4997 2397 5031 2431
rect 7021 2397 7055 2431
rect 7481 2397 7515 2431
rect 9321 2397 9355 2431
rect 9965 2397 9999 2431
rect 14565 2397 14599 2431
rect 21833 2397 21867 2431
rect 29837 2397 29871 2431
rect 30297 2397 30331 2431
rect 33885 2397 33919 2431
rect 9505 2261 9539 2295
rect 14381 2261 14415 2295
rect 22017 2261 22051 2295
rect 29653 2261 29687 2295
rect 34069 2261 34103 2295
<< metal1 >>
rect 1104 17434 34868 17456
rect 1104 17382 9398 17434
rect 9450 17382 9462 17434
rect 9514 17382 9526 17434
rect 9578 17382 9590 17434
rect 9642 17382 9654 17434
rect 9706 17382 17846 17434
rect 17898 17382 17910 17434
rect 17962 17382 17974 17434
rect 18026 17382 18038 17434
rect 18090 17382 18102 17434
rect 18154 17382 26294 17434
rect 26346 17382 26358 17434
rect 26410 17382 26422 17434
rect 26474 17382 26486 17434
rect 26538 17382 26550 17434
rect 26602 17382 34868 17434
rect 1104 17360 34868 17382
rect 3602 17280 3608 17332
rect 3660 17320 3666 17332
rect 3881 17323 3939 17329
rect 3881 17320 3893 17323
rect 3660 17292 3893 17320
rect 3660 17280 3666 17292
rect 3881 17289 3893 17292
rect 3927 17289 3939 17323
rect 3881 17283 3939 17289
rect 10778 17280 10784 17332
rect 10836 17320 10842 17332
rect 11701 17323 11759 17329
rect 11701 17320 11713 17323
rect 10836 17292 11713 17320
rect 10836 17280 10842 17292
rect 11701 17289 11713 17292
rect 11747 17289 11759 17323
rect 11701 17283 11759 17289
rect 18141 17323 18199 17329
rect 18141 17289 18153 17323
rect 18187 17320 18199 17323
rect 18230 17320 18236 17332
rect 18187 17292 18236 17320
rect 18187 17289 18199 17292
rect 18141 17283 18199 17289
rect 18230 17280 18236 17292
rect 18288 17280 18294 17332
rect 25130 17280 25136 17332
rect 25188 17320 25194 17332
rect 25317 17323 25375 17329
rect 25317 17320 25329 17323
rect 25188 17292 25329 17320
rect 25188 17280 25194 17292
rect 25317 17289 25329 17292
rect 25363 17289 25375 17323
rect 25317 17283 25375 17289
rect 32306 17280 32312 17332
rect 32364 17320 32370 17332
rect 32585 17323 32643 17329
rect 32585 17320 32597 17323
rect 32364 17292 32597 17320
rect 32364 17280 32370 17292
rect 32585 17289 32597 17292
rect 32631 17289 32643 17323
rect 34054 17320 34060 17332
rect 34015 17292 34060 17320
rect 32585 17283 32643 17289
rect 34054 17280 34060 17292
rect 34112 17280 34118 17332
rect 1394 17184 1400 17196
rect 1355 17156 1400 17184
rect 1394 17144 1400 17156
rect 1452 17144 1458 17196
rect 4065 17187 4123 17193
rect 4065 17153 4077 17187
rect 4111 17184 4123 17187
rect 6822 17184 6828 17196
rect 4111 17156 6828 17184
rect 4111 17153 4123 17156
rect 4065 17147 4123 17153
rect 6822 17144 6828 17156
rect 6880 17144 6886 17196
rect 11514 17184 11520 17196
rect 11475 17156 11520 17184
rect 11514 17144 11520 17156
rect 11572 17144 11578 17196
rect 18322 17184 18328 17196
rect 18283 17156 18328 17184
rect 18322 17144 18328 17156
rect 18380 17144 18386 17196
rect 25498 17184 25504 17196
rect 25459 17156 25504 17184
rect 25498 17144 25504 17156
rect 25556 17144 25562 17196
rect 29914 17144 29920 17196
rect 29972 17184 29978 17196
rect 32401 17187 32459 17193
rect 32401 17184 32413 17187
rect 29972 17156 32413 17184
rect 29972 17144 29978 17156
rect 32401 17153 32413 17156
rect 32447 17153 32459 17187
rect 32401 17147 32459 17153
rect 33318 17144 33324 17196
rect 33376 17184 33382 17196
rect 33873 17187 33931 17193
rect 33873 17184 33885 17187
rect 33376 17156 33885 17184
rect 33376 17144 33382 17156
rect 33873 17153 33885 17156
rect 33919 17153 33931 17187
rect 33873 17147 33931 17153
rect 1673 17119 1731 17125
rect 1673 17085 1685 17119
rect 1719 17116 1731 17119
rect 1719 17088 6914 17116
rect 1719 17085 1731 17088
rect 1673 17079 1731 17085
rect 6886 17048 6914 17088
rect 20070 17048 20076 17060
rect 6886 17020 20076 17048
rect 20070 17008 20076 17020
rect 20128 17008 20134 17060
rect 33318 16980 33324 16992
rect 33279 16952 33324 16980
rect 33318 16940 33324 16952
rect 33376 16940 33382 16992
rect 1104 16890 34868 16912
rect 1104 16838 5174 16890
rect 5226 16838 5238 16890
rect 5290 16838 5302 16890
rect 5354 16838 5366 16890
rect 5418 16838 5430 16890
rect 5482 16838 13622 16890
rect 13674 16838 13686 16890
rect 13738 16838 13750 16890
rect 13802 16838 13814 16890
rect 13866 16838 13878 16890
rect 13930 16838 22070 16890
rect 22122 16838 22134 16890
rect 22186 16838 22198 16890
rect 22250 16838 22262 16890
rect 22314 16838 22326 16890
rect 22378 16838 30518 16890
rect 30570 16838 30582 16890
rect 30634 16838 30646 16890
rect 30698 16838 30710 16890
rect 30762 16838 30774 16890
rect 30826 16838 34868 16890
rect 1104 16816 34868 16838
rect 1394 16776 1400 16788
rect 1355 16748 1400 16776
rect 1394 16736 1400 16748
rect 1452 16736 1458 16788
rect 6546 16572 6552 16584
rect 6507 16544 6552 16572
rect 6546 16532 6552 16544
rect 6604 16532 6610 16584
rect 31386 16532 31392 16584
rect 31444 16572 31450 16584
rect 33873 16575 33931 16581
rect 33873 16572 33885 16575
rect 31444 16544 33885 16572
rect 31444 16532 31450 16544
rect 33873 16541 33885 16544
rect 33919 16541 33931 16575
rect 33873 16535 33931 16541
rect 6733 16439 6791 16445
rect 6733 16405 6745 16439
rect 6779 16436 6791 16439
rect 7006 16436 7012 16448
rect 6779 16408 7012 16436
rect 6779 16405 6791 16408
rect 6733 16399 6791 16405
rect 7006 16396 7012 16408
rect 7064 16396 7070 16448
rect 34054 16436 34060 16448
rect 34015 16408 34060 16436
rect 34054 16396 34060 16408
rect 34112 16396 34118 16448
rect 1104 16346 34868 16368
rect 1104 16294 9398 16346
rect 9450 16294 9462 16346
rect 9514 16294 9526 16346
rect 9578 16294 9590 16346
rect 9642 16294 9654 16346
rect 9706 16294 17846 16346
rect 17898 16294 17910 16346
rect 17962 16294 17974 16346
rect 18026 16294 18038 16346
rect 18090 16294 18102 16346
rect 18154 16294 26294 16346
rect 26346 16294 26358 16346
rect 26410 16294 26422 16346
rect 26474 16294 26486 16346
rect 26538 16294 26550 16346
rect 26602 16294 34868 16346
rect 1104 16272 34868 16294
rect 6914 16192 6920 16244
rect 6972 16232 6978 16244
rect 8481 16235 8539 16241
rect 8481 16232 8493 16235
rect 6972 16204 8493 16232
rect 6972 16192 6978 16204
rect 8481 16201 8493 16204
rect 8527 16232 8539 16235
rect 11514 16232 11520 16244
rect 8527 16204 11520 16232
rect 8527 16201 8539 16204
rect 8481 16195 8539 16201
rect 11514 16192 11520 16204
rect 11572 16192 11578 16244
rect 21821 16235 21879 16241
rect 21821 16201 21833 16235
rect 21867 16201 21879 16235
rect 21821 16195 21879 16201
rect 28169 16235 28227 16241
rect 28169 16201 28181 16235
rect 28215 16232 28227 16235
rect 29914 16232 29920 16244
rect 28215 16204 29920 16232
rect 28215 16201 28227 16204
rect 28169 16195 28227 16201
rect 7006 16164 7012 16176
rect 6967 16136 7012 16164
rect 7006 16124 7012 16136
rect 7064 16124 7070 16176
rect 8018 16124 8024 16176
rect 8076 16124 8082 16176
rect 15197 16099 15255 16105
rect 15197 16065 15209 16099
rect 15243 16096 15255 16099
rect 17770 16096 17776 16108
rect 15243 16068 17776 16096
rect 15243 16065 15255 16068
rect 15197 16059 15255 16065
rect 17770 16056 17776 16068
rect 17828 16056 17834 16108
rect 20993 16099 21051 16105
rect 20993 16065 21005 16099
rect 21039 16096 21051 16099
rect 21836 16096 21864 16195
rect 29914 16192 29920 16204
rect 29972 16192 29978 16244
rect 22281 16167 22339 16173
rect 22281 16133 22293 16167
rect 22327 16164 22339 16167
rect 22462 16164 22468 16176
rect 22327 16136 22468 16164
rect 22327 16133 22339 16136
rect 22281 16127 22339 16133
rect 22462 16124 22468 16136
rect 22520 16164 22526 16176
rect 25498 16164 25504 16176
rect 22520 16136 25504 16164
rect 22520 16124 22526 16136
rect 25498 16124 25504 16136
rect 25556 16164 25562 16176
rect 28261 16167 28319 16173
rect 28261 16164 28273 16167
rect 25556 16136 28273 16164
rect 25556 16124 25562 16136
rect 28261 16133 28273 16136
rect 28307 16133 28319 16167
rect 28261 16127 28319 16133
rect 21039 16068 21864 16096
rect 21039 16065 21051 16068
rect 20993 16059 21051 16065
rect 21910 16056 21916 16108
rect 21968 16096 21974 16108
rect 22189 16099 22247 16105
rect 22189 16096 22201 16099
rect 21968 16068 22201 16096
rect 21968 16056 21974 16068
rect 22189 16065 22201 16068
rect 22235 16065 22247 16099
rect 29273 16099 29331 16105
rect 29273 16096 29285 16099
rect 22189 16059 22247 16065
rect 28644 16068 29285 16096
rect 6454 15988 6460 16040
rect 6512 16028 6518 16040
rect 6733 16031 6791 16037
rect 6733 16028 6745 16031
rect 6512 16000 6745 16028
rect 6512 15988 6518 16000
rect 6733 15997 6745 16000
rect 6779 16028 6791 16031
rect 8941 16031 8999 16037
rect 8941 16028 8953 16031
rect 6779 16000 8953 16028
rect 6779 15997 6791 16000
rect 6733 15991 6791 15997
rect 8941 15997 8953 16000
rect 8987 16028 8999 16031
rect 13446 16028 13452 16040
rect 8987 16000 13452 16028
rect 8987 15997 8999 16000
rect 8941 15991 8999 15997
rect 13446 15988 13452 16000
rect 13504 15988 13510 16040
rect 18322 15988 18328 16040
rect 18380 16028 18386 16040
rect 21928 16028 21956 16056
rect 18380 16000 21956 16028
rect 22373 16031 22431 16037
rect 18380 15988 18386 16000
rect 22373 15997 22385 16031
rect 22419 16028 22431 16031
rect 27985 16031 28043 16037
rect 27985 16028 27997 16031
rect 22419 16000 27997 16028
rect 22419 15997 22431 16000
rect 22373 15991 22431 15997
rect 27985 15997 27997 16000
rect 28031 15997 28043 16031
rect 27985 15991 28043 15997
rect 14366 15852 14372 15904
rect 14424 15892 14430 15904
rect 15013 15895 15071 15901
rect 15013 15892 15025 15895
rect 14424 15864 15025 15892
rect 14424 15852 14430 15864
rect 15013 15861 15025 15864
rect 15059 15861 15071 15895
rect 15013 15855 15071 15861
rect 20622 15852 20628 15904
rect 20680 15892 20686 15904
rect 20809 15895 20867 15901
rect 20809 15892 20821 15895
rect 20680 15864 20821 15892
rect 20680 15852 20686 15864
rect 20809 15861 20821 15864
rect 20855 15861 20867 15895
rect 20809 15855 20867 15861
rect 21174 15852 21180 15904
rect 21232 15892 21238 15904
rect 22388 15892 22416 15991
rect 28644 15969 28672 16068
rect 29273 16065 29285 16068
rect 29319 16065 29331 16099
rect 29273 16059 29331 16065
rect 28629 15963 28687 15969
rect 28629 15929 28641 15963
rect 28675 15929 28687 15963
rect 28629 15923 28687 15929
rect 29086 15892 29092 15904
rect 21232 15864 22416 15892
rect 29047 15864 29092 15892
rect 21232 15852 21238 15864
rect 29086 15852 29092 15864
rect 29144 15852 29150 15904
rect 1104 15802 34868 15824
rect 1104 15750 5174 15802
rect 5226 15750 5238 15802
rect 5290 15750 5302 15802
rect 5354 15750 5366 15802
rect 5418 15750 5430 15802
rect 5482 15750 13622 15802
rect 13674 15750 13686 15802
rect 13738 15750 13750 15802
rect 13802 15750 13814 15802
rect 13866 15750 13878 15802
rect 13930 15750 22070 15802
rect 22122 15750 22134 15802
rect 22186 15750 22198 15802
rect 22250 15750 22262 15802
rect 22314 15750 22326 15802
rect 22378 15750 30518 15802
rect 30570 15750 30582 15802
rect 30634 15750 30646 15802
rect 30698 15750 30710 15802
rect 30762 15750 30774 15802
rect 30826 15750 34868 15802
rect 1104 15728 34868 15750
rect 6457 15691 6515 15697
rect 6457 15657 6469 15691
rect 6503 15688 6515 15691
rect 6546 15688 6552 15700
rect 6503 15660 6552 15688
rect 6503 15657 6515 15660
rect 6457 15651 6515 15657
rect 6546 15648 6552 15660
rect 6604 15648 6610 15700
rect 7929 15691 7987 15697
rect 7929 15657 7941 15691
rect 7975 15688 7987 15691
rect 8018 15688 8024 15700
rect 7975 15660 8024 15688
rect 7975 15657 7987 15660
rect 7929 15651 7987 15657
rect 8018 15648 8024 15660
rect 8076 15648 8082 15700
rect 13446 15688 13452 15700
rect 13407 15660 13452 15688
rect 13446 15648 13452 15660
rect 13504 15648 13510 15700
rect 15841 15691 15899 15697
rect 15841 15657 15853 15691
rect 15887 15688 15899 15691
rect 18322 15688 18328 15700
rect 15887 15660 18328 15688
rect 15887 15657 15899 15660
rect 15841 15651 15899 15657
rect 18322 15648 18328 15660
rect 18380 15648 18386 15700
rect 22097 15691 22155 15697
rect 22097 15657 22109 15691
rect 22143 15688 22155 15691
rect 22462 15688 22468 15700
rect 22143 15660 22468 15688
rect 22143 15657 22155 15660
rect 22097 15651 22155 15657
rect 22462 15648 22468 15660
rect 22520 15648 22526 15700
rect 6638 15512 6644 15564
rect 6696 15552 6702 15564
rect 7009 15555 7067 15561
rect 7009 15552 7021 15555
rect 6696 15524 7021 15552
rect 6696 15512 6702 15524
rect 7009 15521 7021 15524
rect 7055 15521 7067 15555
rect 13464 15552 13492 15648
rect 14093 15555 14151 15561
rect 14093 15552 14105 15555
rect 13464 15524 14105 15552
rect 7009 15515 7067 15521
rect 14093 15521 14105 15524
rect 14139 15521 14151 15555
rect 14366 15552 14372 15564
rect 14327 15524 14372 15552
rect 14093 15515 14151 15521
rect 14366 15512 14372 15524
rect 14424 15512 14430 15564
rect 20622 15552 20628 15564
rect 20583 15524 20628 15552
rect 20622 15512 20628 15524
rect 20680 15512 20686 15564
rect 6822 15444 6828 15496
rect 6880 15484 6886 15496
rect 8021 15487 8079 15493
rect 8021 15484 8033 15487
rect 6880 15456 8033 15484
rect 6880 15444 6886 15456
rect 8021 15453 8033 15456
rect 8067 15453 8079 15487
rect 20346 15484 20352 15496
rect 20307 15456 20352 15484
rect 8021 15447 8079 15453
rect 20346 15444 20352 15456
rect 20404 15444 20410 15496
rect 6914 15376 6920 15428
rect 6972 15416 6978 15428
rect 6972 15388 7017 15416
rect 6972 15376 6978 15388
rect 15378 15376 15384 15428
rect 15436 15376 15442 15428
rect 19334 15376 19340 15428
rect 19392 15416 19398 15428
rect 19392 15388 21114 15416
rect 19392 15376 19398 15388
rect 6730 15308 6736 15360
rect 6788 15348 6794 15360
rect 6825 15351 6883 15357
rect 6825 15348 6837 15351
rect 6788 15320 6837 15348
rect 6788 15308 6794 15320
rect 6825 15317 6837 15320
rect 6871 15317 6883 15351
rect 6825 15311 6883 15317
rect 1104 15258 34868 15280
rect 1104 15206 9398 15258
rect 9450 15206 9462 15258
rect 9514 15206 9526 15258
rect 9578 15206 9590 15258
rect 9642 15206 9654 15258
rect 9706 15206 17846 15258
rect 17898 15206 17910 15258
rect 17962 15206 17974 15258
rect 18026 15206 18038 15258
rect 18090 15206 18102 15258
rect 18154 15206 26294 15258
rect 26346 15206 26358 15258
rect 26410 15206 26422 15258
rect 26474 15206 26486 15258
rect 26538 15206 26550 15258
rect 26602 15206 34868 15258
rect 1104 15184 34868 15206
rect 14369 15147 14427 15153
rect 14369 15113 14381 15147
rect 14415 15144 14427 15147
rect 15378 15144 15384 15156
rect 14415 15116 15384 15144
rect 14415 15113 14427 15116
rect 14369 15107 14427 15113
rect 15378 15104 15384 15116
rect 15436 15104 15442 15156
rect 17770 15104 17776 15156
rect 17828 15144 17834 15156
rect 20533 15147 20591 15153
rect 20533 15144 20545 15147
rect 17828 15116 20545 15144
rect 17828 15104 17834 15116
rect 20533 15113 20545 15116
rect 20579 15113 20591 15147
rect 20533 15107 20591 15113
rect 20993 15147 21051 15153
rect 20993 15113 21005 15147
rect 21039 15144 21051 15147
rect 21910 15144 21916 15156
rect 21039 15116 21916 15144
rect 21039 15113 21051 15116
rect 20993 15107 21051 15113
rect 21910 15104 21916 15116
rect 21968 15104 21974 15156
rect 29914 15144 29920 15156
rect 29875 15116 29920 15144
rect 29914 15104 29920 15116
rect 29972 15104 29978 15156
rect 24854 15036 24860 15088
rect 24912 15076 24918 15088
rect 24912 15048 28934 15076
rect 24912 15036 24918 15048
rect 14274 15008 14280 15020
rect 14235 14980 14280 15008
rect 14274 14968 14280 14980
rect 14332 15008 14338 15020
rect 15105 15011 15163 15017
rect 15105 15008 15117 15011
rect 14332 14980 15117 15008
rect 14332 14968 14338 14980
rect 15105 14977 15117 14980
rect 15151 14977 15163 15011
rect 15105 14971 15163 14977
rect 20901 15011 20959 15017
rect 20901 14977 20913 15011
rect 20947 15008 20959 15011
rect 20947 14980 21956 15008
rect 20947 14977 20959 14980
rect 20901 14971 20959 14977
rect 21174 14940 21180 14952
rect 21135 14912 21180 14940
rect 21174 14900 21180 14912
rect 21232 14900 21238 14952
rect 15197 14875 15255 14881
rect 15197 14841 15209 14875
rect 15243 14872 15255 14875
rect 19334 14872 19340 14884
rect 15243 14844 19340 14872
rect 15243 14841 15255 14844
rect 15197 14835 15255 14841
rect 19334 14832 19340 14844
rect 19392 14832 19398 14884
rect 6638 14764 6644 14816
rect 6696 14804 6702 14816
rect 21928 14813 21956 14980
rect 28074 14900 28080 14952
rect 28132 14940 28138 14952
rect 28169 14943 28227 14949
rect 28169 14940 28181 14943
rect 28132 14912 28181 14940
rect 28132 14900 28138 14912
rect 28169 14909 28181 14912
rect 28215 14909 28227 14943
rect 28169 14903 28227 14909
rect 28445 14943 28503 14949
rect 28445 14909 28457 14943
rect 28491 14940 28503 14943
rect 29086 14940 29092 14952
rect 28491 14912 29092 14940
rect 28491 14909 28503 14912
rect 28445 14903 28503 14909
rect 29086 14900 29092 14912
rect 29144 14900 29150 14952
rect 7285 14807 7343 14813
rect 7285 14804 7297 14807
rect 6696 14776 7297 14804
rect 6696 14764 6702 14776
rect 7285 14773 7297 14776
rect 7331 14773 7343 14807
rect 7285 14767 7343 14773
rect 21913 14807 21971 14813
rect 21913 14773 21925 14807
rect 21959 14804 21971 14807
rect 29638 14804 29644 14816
rect 21959 14776 29644 14804
rect 21959 14773 21971 14776
rect 21913 14767 21971 14773
rect 29638 14764 29644 14776
rect 29696 14764 29702 14816
rect 1104 14714 34868 14736
rect 1104 14662 5174 14714
rect 5226 14662 5238 14714
rect 5290 14662 5302 14714
rect 5354 14662 5366 14714
rect 5418 14662 5430 14714
rect 5482 14662 13622 14714
rect 13674 14662 13686 14714
rect 13738 14662 13750 14714
rect 13802 14662 13814 14714
rect 13866 14662 13878 14714
rect 13930 14662 22070 14714
rect 22122 14662 22134 14714
rect 22186 14662 22198 14714
rect 22250 14662 22262 14714
rect 22314 14662 22326 14714
rect 22378 14662 30518 14714
rect 30570 14662 30582 14714
rect 30634 14662 30646 14714
rect 30698 14662 30710 14714
rect 30762 14662 30774 14714
rect 30826 14662 34868 14714
rect 1104 14640 34868 14662
rect 6638 14464 6644 14476
rect 6599 14436 6644 14464
rect 6638 14424 6644 14436
rect 6696 14424 6702 14476
rect 5902 14356 5908 14408
rect 5960 14396 5966 14408
rect 6457 14399 6515 14405
rect 6457 14396 6469 14399
rect 5960 14368 6469 14396
rect 5960 14356 5966 14368
rect 6457 14365 6469 14368
rect 6503 14396 6515 14399
rect 6730 14396 6736 14408
rect 6503 14368 6736 14396
rect 6503 14365 6515 14368
rect 6457 14359 6515 14365
rect 6730 14356 6736 14368
rect 6788 14356 6794 14408
rect 6365 14331 6423 14337
rect 6365 14297 6377 14331
rect 6411 14328 6423 14331
rect 6411 14300 6914 14328
rect 6411 14297 6423 14300
rect 6365 14291 6423 14297
rect 5166 14220 5172 14272
rect 5224 14260 5230 14272
rect 5997 14263 6055 14269
rect 5997 14260 6009 14263
rect 5224 14232 6009 14260
rect 5224 14220 5230 14232
rect 5997 14229 6009 14232
rect 6043 14229 6055 14263
rect 6886 14260 6914 14300
rect 7285 14263 7343 14269
rect 7285 14260 7297 14263
rect 6886 14232 7297 14260
rect 5997 14223 6055 14229
rect 7285 14229 7297 14232
rect 7331 14260 7343 14263
rect 12434 14260 12440 14272
rect 7331 14232 12440 14260
rect 7331 14229 7343 14232
rect 7285 14223 7343 14229
rect 12434 14220 12440 14232
rect 12492 14220 12498 14272
rect 1104 14170 34868 14192
rect 1104 14118 9398 14170
rect 9450 14118 9462 14170
rect 9514 14118 9526 14170
rect 9578 14118 9590 14170
rect 9642 14118 9654 14170
rect 9706 14118 17846 14170
rect 17898 14118 17910 14170
rect 17962 14118 17974 14170
rect 18026 14118 18038 14170
rect 18090 14118 18102 14170
rect 18154 14118 26294 14170
rect 26346 14118 26358 14170
rect 26410 14118 26422 14170
rect 26474 14118 26486 14170
rect 26538 14118 26550 14170
rect 26602 14118 34868 14170
rect 1104 14096 34868 14118
rect 29825 14059 29883 14065
rect 29825 14025 29837 14059
rect 29871 14056 29883 14059
rect 31386 14056 31392 14068
rect 29871 14028 31392 14056
rect 29871 14025 29883 14028
rect 29825 14019 29883 14025
rect 31386 14016 31392 14028
rect 31444 14016 31450 14068
rect 28994 13948 29000 14000
rect 29052 13948 29058 14000
rect 5166 13920 5172 13932
rect 5127 13892 5172 13920
rect 5166 13880 5172 13892
rect 5224 13880 5230 13932
rect 28074 13920 28080 13932
rect 28035 13892 28080 13920
rect 28074 13880 28080 13892
rect 28132 13880 28138 13932
rect 31478 13880 31484 13932
rect 31536 13920 31542 13932
rect 33873 13923 33931 13929
rect 33873 13920 33885 13923
rect 31536 13892 33885 13920
rect 31536 13880 31542 13892
rect 33873 13889 33885 13892
rect 33919 13889 33931 13923
rect 33873 13883 33931 13889
rect 6730 13812 6736 13864
rect 6788 13852 6794 13864
rect 6825 13855 6883 13861
rect 6825 13852 6837 13855
rect 6788 13824 6837 13852
rect 6788 13812 6794 13824
rect 6825 13821 6837 13824
rect 6871 13821 6883 13855
rect 28350 13852 28356 13864
rect 28311 13824 28356 13852
rect 6825 13815 6883 13821
rect 28350 13812 28356 13824
rect 28408 13812 28414 13864
rect 4430 13676 4436 13728
rect 4488 13716 4494 13728
rect 4985 13719 5043 13725
rect 4985 13716 4997 13719
rect 4488 13688 4997 13716
rect 4488 13676 4494 13688
rect 4985 13685 4997 13688
rect 5031 13685 5043 13719
rect 34054 13716 34060 13728
rect 34015 13688 34060 13716
rect 4985 13679 5043 13685
rect 34054 13676 34060 13688
rect 34112 13676 34118 13728
rect 1104 13626 34868 13648
rect 1104 13574 5174 13626
rect 5226 13574 5238 13626
rect 5290 13574 5302 13626
rect 5354 13574 5366 13626
rect 5418 13574 5430 13626
rect 5482 13574 13622 13626
rect 13674 13574 13686 13626
rect 13738 13574 13750 13626
rect 13802 13574 13814 13626
rect 13866 13574 13878 13626
rect 13930 13574 22070 13626
rect 22122 13574 22134 13626
rect 22186 13574 22198 13626
rect 22250 13574 22262 13626
rect 22314 13574 22326 13626
rect 22378 13574 30518 13626
rect 30570 13574 30582 13626
rect 30634 13574 30646 13626
rect 30698 13574 30710 13626
rect 30762 13574 30774 13626
rect 30826 13574 34868 13626
rect 1104 13552 34868 13574
rect 5902 13512 5908 13524
rect 5863 13484 5908 13512
rect 5902 13472 5908 13484
rect 5960 13472 5966 13524
rect 6454 13512 6460 13524
rect 6415 13484 6460 13512
rect 6454 13472 6460 13484
rect 6512 13472 6518 13524
rect 20070 13472 20076 13524
rect 20128 13512 20134 13524
rect 20165 13515 20223 13521
rect 20165 13512 20177 13515
rect 20128 13484 20177 13512
rect 20128 13472 20134 13484
rect 20165 13481 20177 13484
rect 20211 13481 20223 13515
rect 20165 13475 20223 13481
rect 21729 13515 21787 13521
rect 21729 13481 21741 13515
rect 21775 13512 21787 13515
rect 24854 13512 24860 13524
rect 21775 13484 24860 13512
rect 21775 13481 21787 13484
rect 21729 13475 21787 13481
rect 24854 13472 24860 13484
rect 24912 13472 24918 13524
rect 28350 13472 28356 13524
rect 28408 13512 28414 13524
rect 29733 13515 29791 13521
rect 29733 13512 29745 13515
rect 28408 13484 29745 13512
rect 28408 13472 28414 13484
rect 29733 13481 29745 13484
rect 29779 13481 29791 13515
rect 29733 13475 29791 13481
rect 4157 13379 4215 13385
rect 4157 13345 4169 13379
rect 4203 13376 4215 13379
rect 6472 13376 6500 13472
rect 30374 13404 30380 13456
rect 30432 13444 30438 13456
rect 30432 13416 31616 13444
rect 30432 13404 30438 13416
rect 31478 13376 31484 13388
rect 4203 13348 6500 13376
rect 31439 13348 31484 13376
rect 4203 13345 4215 13348
rect 4157 13339 4215 13345
rect 31478 13336 31484 13348
rect 31536 13336 31542 13388
rect 31588 13385 31616 13416
rect 31573 13379 31631 13385
rect 31573 13345 31585 13379
rect 31619 13345 31631 13379
rect 31573 13339 31631 13345
rect 14274 13308 14280 13320
rect 14235 13280 14280 13308
rect 14274 13268 14280 13280
rect 14332 13268 14338 13320
rect 19242 13268 19248 13320
rect 19300 13308 19306 13320
rect 21637 13311 21695 13317
rect 21637 13308 21649 13311
rect 19300 13280 21649 13308
rect 19300 13268 19306 13280
rect 21637 13277 21649 13280
rect 21683 13308 21695 13311
rect 22281 13311 22339 13317
rect 22281 13308 22293 13311
rect 21683 13280 22293 13308
rect 21683 13277 21695 13280
rect 21637 13271 21695 13277
rect 22281 13277 22293 13280
rect 22327 13277 22339 13311
rect 22281 13271 22339 13277
rect 29917 13311 29975 13317
rect 29917 13277 29929 13311
rect 29963 13308 29975 13311
rect 31386 13308 31392 13320
rect 29963 13280 31064 13308
rect 31347 13280 31392 13308
rect 29963 13277 29975 13280
rect 29917 13271 29975 13277
rect 4430 13240 4436 13252
rect 4391 13212 4436 13240
rect 4430 13200 4436 13212
rect 4488 13200 4494 13252
rect 6362 13240 6368 13252
rect 5658 13212 6368 13240
rect 6362 13200 6368 13212
rect 6420 13200 6426 13252
rect 14182 13172 14188 13184
rect 14143 13144 14188 13172
rect 14182 13132 14188 13144
rect 14240 13132 14246 13184
rect 20714 13172 20720 13184
rect 20675 13144 20720 13172
rect 20714 13132 20720 13144
rect 20772 13132 20778 13184
rect 30374 13132 30380 13184
rect 30432 13172 30438 13184
rect 31036 13181 31064 13280
rect 31386 13268 31392 13280
rect 31444 13268 31450 13320
rect 30469 13175 30527 13181
rect 30469 13172 30481 13175
rect 30432 13144 30481 13172
rect 30432 13132 30438 13144
rect 30469 13141 30481 13144
rect 30515 13141 30527 13175
rect 30469 13135 30527 13141
rect 31021 13175 31079 13181
rect 31021 13141 31033 13175
rect 31067 13141 31079 13175
rect 31021 13135 31079 13141
rect 1104 13082 34868 13104
rect 1104 13030 9398 13082
rect 9450 13030 9462 13082
rect 9514 13030 9526 13082
rect 9578 13030 9590 13082
rect 9642 13030 9654 13082
rect 9706 13030 17846 13082
rect 17898 13030 17910 13082
rect 17962 13030 17974 13082
rect 18026 13030 18038 13082
rect 18090 13030 18102 13082
rect 18154 13030 26294 13082
rect 26346 13030 26358 13082
rect 26410 13030 26422 13082
rect 26474 13030 26486 13082
rect 26538 13030 26550 13082
rect 26602 13030 34868 13082
rect 1104 13008 34868 13030
rect 6362 12928 6368 12980
rect 6420 12968 6426 12980
rect 6457 12971 6515 12977
rect 6457 12968 6469 12971
rect 6420 12940 6469 12968
rect 6420 12928 6426 12940
rect 6457 12937 6469 12940
rect 6503 12937 6515 12971
rect 12894 12968 12900 12980
rect 12807 12940 12900 12968
rect 6457 12931 6515 12937
rect 12894 12928 12900 12940
rect 12952 12968 12958 12980
rect 13446 12968 13452 12980
rect 12952 12940 13452 12968
rect 12952 12928 12958 12940
rect 13446 12928 13452 12940
rect 13504 12968 13510 12980
rect 13504 12940 15240 12968
rect 13504 12928 13510 12940
rect 14182 12860 14188 12912
rect 14240 12860 14246 12912
rect 6549 12835 6607 12841
rect 6549 12801 6561 12835
rect 6595 12832 6607 12835
rect 6822 12832 6828 12844
rect 6595 12804 6828 12832
rect 6595 12801 6607 12804
rect 6549 12795 6607 12801
rect 6822 12792 6828 12804
rect 6880 12832 6886 12844
rect 15212 12841 15240 12940
rect 15286 12928 15292 12980
rect 15344 12968 15350 12980
rect 20254 12968 20260 12980
rect 15344 12940 20260 12968
rect 15344 12928 15350 12940
rect 20254 12928 20260 12940
rect 20312 12928 20318 12980
rect 20901 12971 20959 12977
rect 20901 12937 20913 12971
rect 20947 12968 20959 12971
rect 21174 12968 21180 12980
rect 20947 12940 21180 12968
rect 20947 12937 20959 12940
rect 20901 12931 20959 12937
rect 21174 12928 21180 12940
rect 21232 12928 21238 12980
rect 28537 12971 28595 12977
rect 28537 12937 28549 12971
rect 28583 12968 28595 12971
rect 28994 12968 29000 12980
rect 28583 12940 29000 12968
rect 28583 12937 28595 12940
rect 28537 12931 28595 12937
rect 28994 12928 29000 12940
rect 29052 12928 29058 12980
rect 15197 12835 15255 12841
rect 6880 12792 6914 12832
rect 15197 12801 15209 12835
rect 15243 12801 15255 12835
rect 15197 12795 15255 12801
rect 19797 12835 19855 12841
rect 19797 12801 19809 12835
rect 19843 12832 19855 12835
rect 20806 12832 20812 12844
rect 19843 12804 20812 12832
rect 19843 12801 19855 12804
rect 19797 12795 19855 12801
rect 20806 12792 20812 12804
rect 20864 12792 20870 12844
rect 27890 12792 27896 12844
rect 27948 12832 27954 12844
rect 28445 12835 28503 12841
rect 28445 12832 28457 12835
rect 27948 12804 28457 12832
rect 27948 12792 27954 12804
rect 28445 12801 28457 12804
rect 28491 12832 28503 12835
rect 29089 12835 29147 12841
rect 29089 12832 29101 12835
rect 28491 12804 29101 12832
rect 28491 12801 28503 12804
rect 28445 12795 28503 12801
rect 29089 12801 29101 12804
rect 29135 12801 29147 12835
rect 29089 12795 29147 12801
rect 1394 12764 1400 12776
rect 1355 12736 1400 12764
rect 1394 12724 1400 12736
rect 1452 12724 1458 12776
rect 1673 12767 1731 12773
rect 1673 12733 1685 12767
rect 1719 12764 1731 12767
rect 6362 12764 6368 12776
rect 1719 12736 6368 12764
rect 1719 12733 1731 12736
rect 1673 12727 1731 12733
rect 6362 12724 6368 12736
rect 6420 12724 6426 12776
rect 6886 12764 6914 12792
rect 14274 12764 14280 12776
rect 6886 12736 14280 12764
rect 14274 12724 14280 12736
rect 14332 12724 14338 12776
rect 14921 12767 14979 12773
rect 14921 12733 14933 12767
rect 14967 12764 14979 12767
rect 14967 12736 16574 12764
rect 14967 12733 14979 12736
rect 14921 12727 14979 12733
rect 16546 12696 16574 12736
rect 20070 12724 20076 12776
rect 20128 12764 20134 12776
rect 20717 12767 20775 12773
rect 20717 12764 20729 12767
rect 20128 12736 20729 12764
rect 20128 12724 20134 12736
rect 20717 12733 20729 12736
rect 20763 12733 20775 12767
rect 21082 12764 21088 12776
rect 20995 12736 21088 12764
rect 20717 12727 20775 12733
rect 21082 12724 21088 12736
rect 21140 12764 21146 12776
rect 21140 12736 21956 12764
rect 21140 12724 21146 12736
rect 19613 12699 19671 12705
rect 19613 12696 19625 12699
rect 16546 12668 19625 12696
rect 19613 12665 19625 12668
rect 19659 12665 19671 12699
rect 19613 12659 19671 12665
rect 12434 12588 12440 12640
rect 12492 12628 12498 12640
rect 13449 12631 13507 12637
rect 13449 12628 13461 12631
rect 12492 12600 13461 12628
rect 12492 12588 12498 12600
rect 13449 12597 13461 12600
rect 13495 12628 13507 12631
rect 15286 12628 15292 12640
rect 13495 12600 15292 12628
rect 13495 12597 13507 12600
rect 13449 12591 13507 12597
rect 15286 12588 15292 12600
rect 15344 12588 15350 12640
rect 20714 12588 20720 12640
rect 20772 12628 20778 12640
rect 21928 12637 21956 12736
rect 21085 12631 21143 12637
rect 21085 12628 21097 12631
rect 20772 12600 21097 12628
rect 20772 12588 20778 12600
rect 21085 12597 21097 12600
rect 21131 12597 21143 12631
rect 21085 12591 21143 12597
rect 21913 12631 21971 12637
rect 21913 12597 21925 12631
rect 21959 12628 21971 12631
rect 22830 12628 22836 12640
rect 21959 12600 22836 12628
rect 21959 12597 21971 12600
rect 21913 12591 21971 12597
rect 22830 12588 22836 12600
rect 22888 12588 22894 12640
rect 1104 12538 34868 12560
rect 1104 12486 5174 12538
rect 5226 12486 5238 12538
rect 5290 12486 5302 12538
rect 5354 12486 5366 12538
rect 5418 12486 5430 12538
rect 5482 12486 13622 12538
rect 13674 12486 13686 12538
rect 13738 12486 13750 12538
rect 13802 12486 13814 12538
rect 13866 12486 13878 12538
rect 13930 12486 22070 12538
rect 22122 12486 22134 12538
rect 22186 12486 22198 12538
rect 22250 12486 22262 12538
rect 22314 12486 22326 12538
rect 22378 12486 30518 12538
rect 30570 12486 30582 12538
rect 30634 12486 30646 12538
rect 30698 12486 30710 12538
rect 30762 12486 30774 12538
rect 30826 12486 34868 12538
rect 1104 12464 34868 12486
rect 1394 12424 1400 12436
rect 1355 12396 1400 12424
rect 1394 12384 1400 12396
rect 1452 12384 1458 12436
rect 6641 12427 6699 12433
rect 6641 12393 6653 12427
rect 6687 12424 6699 12427
rect 6822 12424 6828 12436
rect 6687 12396 6828 12424
rect 6687 12393 6699 12396
rect 6641 12387 6699 12393
rect 6822 12384 6828 12396
rect 6880 12384 6886 12436
rect 20717 12427 20775 12433
rect 20717 12393 20729 12427
rect 20763 12424 20775 12427
rect 20806 12424 20812 12436
rect 20763 12396 20812 12424
rect 20763 12393 20775 12396
rect 20717 12387 20775 12393
rect 20806 12384 20812 12396
rect 20864 12384 20870 12436
rect 21266 12288 21272 12300
rect 21227 12260 21272 12288
rect 21266 12248 21272 12260
rect 21324 12248 21330 12300
rect 6825 12223 6883 12229
rect 6825 12220 6837 12223
rect 6012 12192 6837 12220
rect 6012 12096 6040 12192
rect 6825 12189 6837 12192
rect 6871 12220 6883 12223
rect 27890 12220 27896 12232
rect 6871 12192 27896 12220
rect 6871 12189 6883 12192
rect 6825 12183 6883 12189
rect 27890 12180 27896 12192
rect 27948 12180 27954 12232
rect 21085 12155 21143 12161
rect 21085 12121 21097 12155
rect 21131 12152 21143 12155
rect 21634 12152 21640 12164
rect 21131 12124 21640 12152
rect 21131 12121 21143 12124
rect 21085 12115 21143 12121
rect 21634 12112 21640 12124
rect 21692 12112 21698 12164
rect 5994 12084 6000 12096
rect 5955 12056 6000 12084
rect 5994 12044 6000 12056
rect 6052 12044 6058 12096
rect 20254 12084 20260 12096
rect 20167 12056 20260 12084
rect 20254 12044 20260 12056
rect 20312 12084 20318 12096
rect 21177 12087 21235 12093
rect 21177 12084 21189 12087
rect 20312 12056 21189 12084
rect 20312 12044 20318 12056
rect 21177 12053 21189 12056
rect 21223 12084 21235 12087
rect 33318 12084 33324 12096
rect 21223 12056 33324 12084
rect 21223 12053 21235 12056
rect 21177 12047 21235 12053
rect 33318 12044 33324 12056
rect 33376 12044 33382 12096
rect 1104 11994 34868 12016
rect 1104 11942 9398 11994
rect 9450 11942 9462 11994
rect 9514 11942 9526 11994
rect 9578 11942 9590 11994
rect 9642 11942 9654 11994
rect 9706 11942 17846 11994
rect 17898 11942 17910 11994
rect 17962 11942 17974 11994
rect 18026 11942 18038 11994
rect 18090 11942 18102 11994
rect 18154 11942 26294 11994
rect 26346 11942 26358 11994
rect 26410 11942 26422 11994
rect 26474 11942 26486 11994
rect 26538 11942 26550 11994
rect 26602 11942 34868 11994
rect 1104 11920 34868 11942
rect 6362 11744 6368 11756
rect 6323 11716 6368 11744
rect 6362 11704 6368 11716
rect 6420 11744 6426 11756
rect 20714 11744 20720 11756
rect 6420 11716 20720 11744
rect 6420 11704 6426 11716
rect 20714 11704 20720 11716
rect 20772 11704 20778 11756
rect 31478 11704 31484 11756
rect 31536 11744 31542 11756
rect 33873 11747 33931 11753
rect 33873 11744 33885 11747
rect 31536 11716 33885 11744
rect 31536 11704 31542 11716
rect 33873 11713 33885 11716
rect 33919 11713 33931 11747
rect 33873 11707 33931 11713
rect 6730 11568 6736 11620
rect 6788 11608 6794 11620
rect 6825 11611 6883 11617
rect 6825 11608 6837 11611
rect 6788 11580 6837 11608
rect 6788 11568 6794 11580
rect 6825 11577 6837 11580
rect 6871 11608 6883 11611
rect 20533 11611 20591 11617
rect 20533 11608 20545 11611
rect 6871 11580 20545 11608
rect 6871 11577 6883 11580
rect 6825 11571 6883 11577
rect 20533 11577 20545 11580
rect 20579 11608 20591 11611
rect 21266 11608 21272 11620
rect 20579 11580 21272 11608
rect 20579 11577 20591 11580
rect 20533 11571 20591 11577
rect 21266 11568 21272 11580
rect 21324 11568 21330 11620
rect 5718 11540 5724 11552
rect 5679 11512 5724 11540
rect 5718 11500 5724 11512
rect 5776 11540 5782 11552
rect 6457 11543 6515 11549
rect 6457 11540 6469 11543
rect 5776 11512 6469 11540
rect 5776 11500 5782 11512
rect 6457 11509 6469 11512
rect 6503 11540 6515 11543
rect 21082 11540 21088 11552
rect 6503 11512 21088 11540
rect 6503 11509 6515 11512
rect 6457 11503 6515 11509
rect 21082 11500 21088 11512
rect 21140 11500 21146 11552
rect 34054 11540 34060 11552
rect 34015 11512 34060 11540
rect 34054 11500 34060 11512
rect 34112 11500 34118 11552
rect 1104 11450 34868 11472
rect 1104 11398 5174 11450
rect 5226 11398 5238 11450
rect 5290 11398 5302 11450
rect 5354 11398 5366 11450
rect 5418 11398 5430 11450
rect 5482 11398 13622 11450
rect 13674 11398 13686 11450
rect 13738 11398 13750 11450
rect 13802 11398 13814 11450
rect 13866 11398 13878 11450
rect 13930 11398 22070 11450
rect 22122 11398 22134 11450
rect 22186 11398 22198 11450
rect 22250 11398 22262 11450
rect 22314 11398 22326 11450
rect 22378 11398 30518 11450
rect 30570 11398 30582 11450
rect 30634 11398 30646 11450
rect 30698 11398 30710 11450
rect 30762 11398 30774 11450
rect 30826 11398 34868 11450
rect 1104 11376 34868 11398
rect 6089 11339 6147 11345
rect 6089 11305 6101 11339
rect 6135 11336 6147 11339
rect 6362 11336 6368 11348
rect 6135 11308 6368 11336
rect 6135 11305 6147 11308
rect 6089 11299 6147 11305
rect 6362 11296 6368 11308
rect 6420 11296 6426 11348
rect 11238 11336 11244 11348
rect 11151 11308 11244 11336
rect 11238 11296 11244 11308
rect 11296 11336 11302 11348
rect 12894 11336 12900 11348
rect 11296 11308 12900 11336
rect 11296 11296 11302 11308
rect 12894 11296 12900 11308
rect 12952 11336 12958 11348
rect 21266 11336 21272 11348
rect 12952 11308 13584 11336
rect 12952 11296 12958 11308
rect 11793 11203 11851 11209
rect 11793 11169 11805 11203
rect 11839 11200 11851 11203
rect 12618 11200 12624 11212
rect 11839 11172 12624 11200
rect 11839 11169 11851 11172
rect 11793 11163 11851 11169
rect 12618 11160 12624 11172
rect 12676 11160 12682 11212
rect 13556 11209 13584 11308
rect 19444 11308 21272 11336
rect 19444 11209 19472 11308
rect 21266 11296 21272 11308
rect 21324 11296 21330 11348
rect 27890 11336 27896 11348
rect 27851 11308 27896 11336
rect 27890 11296 27896 11308
rect 27948 11296 27954 11348
rect 20441 11271 20499 11277
rect 20441 11237 20453 11271
rect 20487 11268 20499 11271
rect 20714 11268 20720 11280
rect 20487 11240 20720 11268
rect 20487 11237 20499 11240
rect 20441 11231 20499 11237
rect 20714 11228 20720 11240
rect 20772 11228 20778 11280
rect 31021 11271 31079 11277
rect 31021 11237 31033 11271
rect 31067 11237 31079 11271
rect 31021 11231 31079 11237
rect 13541 11203 13599 11209
rect 13541 11169 13553 11203
rect 13587 11169 13599 11203
rect 13541 11163 13599 11169
rect 19429 11203 19487 11209
rect 19429 11169 19441 11203
rect 19475 11169 19487 11203
rect 19429 11163 19487 11169
rect 19705 11135 19763 11141
rect 19705 11101 19717 11135
rect 19751 11101 19763 11135
rect 19705 11095 19763 11101
rect 12710 11024 12716 11076
rect 12768 11024 12774 11076
rect 13262 11064 13268 11076
rect 13223 11036 13268 11064
rect 13262 11024 13268 11036
rect 13320 11024 13326 11076
rect 14366 11024 14372 11076
rect 14424 11064 14430 11076
rect 19720 11064 19748 11095
rect 27890 11092 27896 11144
rect 27948 11132 27954 11144
rect 28445 11135 28503 11141
rect 28445 11132 28457 11135
rect 27948 11104 28457 11132
rect 27948 11092 27954 11104
rect 28445 11101 28457 11104
rect 28491 11101 28503 11135
rect 28445 11095 28503 11101
rect 29917 11135 29975 11141
rect 29917 11101 29929 11135
rect 29963 11132 29975 11135
rect 31036 11132 31064 11231
rect 31573 11203 31631 11209
rect 31573 11200 31585 11203
rect 29963 11104 31064 11132
rect 31128 11172 31585 11200
rect 29963 11101 29975 11104
rect 29917 11095 29975 11101
rect 14424 11036 19748 11064
rect 28537 11067 28595 11073
rect 14424 11024 14430 11036
rect 28537 11033 28549 11067
rect 28583 11064 28595 11067
rect 28994 11064 29000 11076
rect 28583 11036 29000 11064
rect 28583 11033 28595 11036
rect 28537 11027 28595 11033
rect 28994 11024 29000 11036
rect 29052 11024 29058 11076
rect 30374 11024 30380 11076
rect 30432 11064 30438 11076
rect 30469 11067 30527 11073
rect 30469 11064 30481 11067
rect 30432 11036 30481 11064
rect 30432 11024 30438 11036
rect 30469 11033 30481 11036
rect 30515 11064 30527 11067
rect 31128 11064 31156 11172
rect 31573 11169 31585 11172
rect 31619 11169 31631 11203
rect 31573 11163 31631 11169
rect 31386 11064 31392 11076
rect 30515 11036 31156 11064
rect 31347 11036 31392 11064
rect 30515 11033 30527 11036
rect 30469 11027 30527 11033
rect 31386 11024 31392 11036
rect 31444 11024 31450 11076
rect 31478 11024 31484 11076
rect 31536 11064 31542 11076
rect 31536 11036 31581 11064
rect 31536 11024 31542 11036
rect 29730 10996 29736 11008
rect 29691 10968 29736 10996
rect 29730 10956 29736 10968
rect 29788 10956 29794 11008
rect 1104 10906 34868 10928
rect 1104 10854 9398 10906
rect 9450 10854 9462 10906
rect 9514 10854 9526 10906
rect 9578 10854 9590 10906
rect 9642 10854 9654 10906
rect 9706 10854 17846 10906
rect 17898 10854 17910 10906
rect 17962 10854 17974 10906
rect 18026 10854 18038 10906
rect 18090 10854 18102 10906
rect 18154 10854 26294 10906
rect 26346 10854 26358 10906
rect 26410 10854 26422 10906
rect 26474 10854 26486 10906
rect 26538 10854 26550 10906
rect 26602 10854 34868 10906
rect 1104 10832 34868 10854
rect 12710 10792 12716 10804
rect 12671 10764 12716 10792
rect 12710 10752 12716 10764
rect 12768 10752 12774 10804
rect 19242 10792 19248 10804
rect 16546 10764 19248 10792
rect 3878 10616 3884 10668
rect 3936 10656 3942 10668
rect 4433 10659 4491 10665
rect 4433 10656 4445 10659
rect 3936 10628 4445 10656
rect 3936 10616 3942 10628
rect 4433 10625 4445 10628
rect 4479 10656 4491 10659
rect 5994 10656 6000 10668
rect 4479 10628 6000 10656
rect 4479 10625 4491 10628
rect 4433 10619 4491 10625
rect 5994 10616 6000 10628
rect 6052 10616 6058 10668
rect 12802 10656 12808 10668
rect 12763 10628 12808 10656
rect 12802 10616 12808 10628
rect 12860 10656 12866 10668
rect 13265 10659 13323 10665
rect 13265 10656 13277 10659
rect 12860 10628 13277 10656
rect 12860 10616 12866 10628
rect 13265 10625 13277 10628
rect 13311 10656 13323 10659
rect 16546 10656 16574 10764
rect 19242 10752 19248 10764
rect 19300 10752 19306 10804
rect 29733 10795 29791 10801
rect 29733 10761 29745 10795
rect 29779 10792 29791 10795
rect 31386 10792 31392 10804
rect 29779 10764 31392 10792
rect 29779 10761 29791 10764
rect 29733 10755 29791 10761
rect 31386 10752 31392 10764
rect 31444 10752 31450 10804
rect 28994 10684 29000 10736
rect 29052 10684 29058 10736
rect 13311 10628 16574 10656
rect 13311 10625 13323 10628
rect 13265 10619 13323 10625
rect 17678 10616 17684 10668
rect 17736 10656 17742 10668
rect 18233 10659 18291 10665
rect 18233 10656 18245 10659
rect 17736 10628 18245 10656
rect 17736 10616 17742 10628
rect 18233 10625 18245 10628
rect 18279 10625 18291 10659
rect 18233 10619 18291 10625
rect 19981 10659 20039 10665
rect 19981 10625 19993 10659
rect 20027 10656 20039 10659
rect 20346 10656 20352 10668
rect 20027 10628 20352 10656
rect 20027 10625 20039 10628
rect 19981 10619 20039 10625
rect 20346 10616 20352 10628
rect 20404 10656 20410 10668
rect 27798 10656 27804 10668
rect 20404 10628 27804 10656
rect 20404 10616 20410 10628
rect 27798 10616 27804 10628
rect 27856 10656 27862 10668
rect 27982 10656 27988 10668
rect 27856 10628 27988 10656
rect 27856 10616 27862 10628
rect 27982 10616 27988 10628
rect 28040 10616 28046 10668
rect 28261 10591 28319 10597
rect 28261 10557 28273 10591
rect 28307 10588 28319 10591
rect 29730 10588 29736 10600
rect 28307 10560 29736 10588
rect 28307 10557 28319 10560
rect 28261 10551 28319 10557
rect 29730 10548 29736 10560
rect 29788 10548 29794 10600
rect 3878 10452 3884 10464
rect 3839 10424 3884 10452
rect 3878 10412 3884 10424
rect 3936 10412 3942 10464
rect 4617 10455 4675 10461
rect 4617 10421 4629 10455
rect 4663 10452 4675 10455
rect 4798 10452 4804 10464
rect 4663 10424 4804 10452
rect 4663 10421 4675 10424
rect 4617 10415 4675 10421
rect 4798 10412 4804 10424
rect 4856 10412 4862 10464
rect 1104 10362 34868 10384
rect 1104 10310 5174 10362
rect 5226 10310 5238 10362
rect 5290 10310 5302 10362
rect 5354 10310 5366 10362
rect 5418 10310 5430 10362
rect 5482 10310 13622 10362
rect 13674 10310 13686 10362
rect 13738 10310 13750 10362
rect 13802 10310 13814 10362
rect 13866 10310 13878 10362
rect 13930 10310 22070 10362
rect 22122 10310 22134 10362
rect 22186 10310 22198 10362
rect 22250 10310 22262 10362
rect 22314 10310 22326 10362
rect 22378 10310 30518 10362
rect 30570 10310 30582 10362
rect 30634 10310 30646 10362
rect 30698 10310 30710 10362
rect 30762 10310 30774 10362
rect 30826 10310 34868 10362
rect 1104 10288 34868 10310
rect 10873 10251 10931 10257
rect 10873 10217 10885 10251
rect 10919 10248 10931 10251
rect 11238 10248 11244 10260
rect 10919 10220 11244 10248
rect 10919 10217 10931 10220
rect 10873 10211 10931 10217
rect 11238 10208 11244 10220
rect 11296 10208 11302 10260
rect 13081 10251 13139 10257
rect 13081 10217 13093 10251
rect 13127 10248 13139 10251
rect 13262 10248 13268 10260
rect 13127 10220 13268 10248
rect 13127 10217 13139 10220
rect 13081 10211 13139 10217
rect 13262 10208 13268 10220
rect 13320 10208 13326 10260
rect 20070 10208 20076 10260
rect 20128 10248 20134 10260
rect 20257 10251 20315 10257
rect 20257 10248 20269 10251
rect 20128 10220 20269 10248
rect 20128 10208 20134 10220
rect 20257 10217 20269 10220
rect 20303 10217 20315 10251
rect 20257 10211 20315 10217
rect 17678 10112 17684 10124
rect 12176 10084 17684 10112
rect 4798 10004 4804 10056
rect 4856 10044 4862 10056
rect 12176 10053 12204 10084
rect 17678 10072 17684 10084
rect 17736 10072 17742 10124
rect 21266 10072 21272 10124
rect 21324 10112 21330 10124
rect 21324 10084 21369 10112
rect 21324 10072 21330 10084
rect 4893 10047 4951 10053
rect 4893 10044 4905 10047
rect 4856 10016 4905 10044
rect 4856 10004 4862 10016
rect 4893 10013 4905 10016
rect 4939 10044 4951 10047
rect 5537 10047 5595 10053
rect 5537 10044 5549 10047
rect 4939 10016 5549 10044
rect 4939 10013 4951 10016
rect 4893 10007 4951 10013
rect 5537 10013 5549 10016
rect 5583 10013 5595 10047
rect 5537 10007 5595 10013
rect 12161 10047 12219 10053
rect 12161 10013 12173 10047
rect 12207 10013 12219 10047
rect 12161 10007 12219 10013
rect 13265 10047 13323 10053
rect 13265 10013 13277 10047
rect 13311 10013 13323 10047
rect 13265 10007 13323 10013
rect 13541 10047 13599 10053
rect 13541 10013 13553 10047
rect 13587 10044 13599 10047
rect 14274 10044 14280 10056
rect 13587 10016 14280 10044
rect 13587 10013 13599 10016
rect 13541 10007 13599 10013
rect 13280 9976 13308 10007
rect 14274 10004 14280 10016
rect 14332 10004 14338 10056
rect 20990 10044 20996 10056
rect 20951 10016 20996 10044
rect 20990 10004 20996 10016
rect 21048 10004 21054 10056
rect 14366 9976 14372 9988
rect 13280 9948 14372 9976
rect 14366 9936 14372 9948
rect 14424 9936 14430 9988
rect 15933 9979 15991 9985
rect 15933 9945 15945 9979
rect 15979 9945 15991 9979
rect 15933 9939 15991 9945
rect 4982 9908 4988 9920
rect 4943 9880 4988 9908
rect 4982 9868 4988 9880
rect 5040 9868 5046 9920
rect 13449 9911 13507 9917
rect 13449 9877 13461 9911
rect 13495 9908 13507 9911
rect 13630 9908 13636 9920
rect 13495 9880 13636 9908
rect 13495 9877 13507 9880
rect 13449 9871 13507 9877
rect 13630 9868 13636 9880
rect 13688 9868 13694 9920
rect 15378 9908 15384 9920
rect 15339 9880 15384 9908
rect 15378 9868 15384 9880
rect 15436 9908 15442 9920
rect 15948 9908 15976 9939
rect 15436 9880 15976 9908
rect 15436 9868 15442 9880
rect 1104 9818 34868 9840
rect 1104 9766 9398 9818
rect 9450 9766 9462 9818
rect 9514 9766 9526 9818
rect 9578 9766 9590 9818
rect 9642 9766 9654 9818
rect 9706 9766 17846 9818
rect 17898 9766 17910 9818
rect 17962 9766 17974 9818
rect 18026 9766 18038 9818
rect 18090 9766 18102 9818
rect 18154 9766 26294 9818
rect 26346 9766 26358 9818
rect 26410 9766 26422 9818
rect 26474 9766 26486 9818
rect 26538 9766 26550 9818
rect 26602 9766 34868 9818
rect 1104 9744 34868 9766
rect 4890 9664 4896 9716
rect 4948 9704 4954 9716
rect 12802 9704 12808 9716
rect 4948 9676 12808 9704
rect 4948 9664 4954 9676
rect 12802 9664 12808 9676
rect 12860 9664 12866 9716
rect 13725 9707 13783 9713
rect 13725 9673 13737 9707
rect 13771 9704 13783 9707
rect 14366 9704 14372 9716
rect 13771 9676 14372 9704
rect 13771 9673 13783 9676
rect 13725 9667 13783 9673
rect 14366 9664 14372 9676
rect 14424 9664 14430 9716
rect 4982 9596 4988 9648
rect 5040 9596 5046 9648
rect 6454 9636 6460 9648
rect 6415 9608 6460 9636
rect 6454 9596 6460 9608
rect 6512 9596 6518 9648
rect 12250 9528 12256 9580
rect 12308 9568 12314 9580
rect 13630 9568 13636 9580
rect 12308 9540 13636 9568
rect 12308 9528 12314 9540
rect 13630 9528 13636 9540
rect 13688 9528 13694 9580
rect 13817 9571 13875 9577
rect 13817 9537 13829 9571
rect 13863 9537 13875 9571
rect 13817 9531 13875 9537
rect 3973 9503 4031 9509
rect 3973 9469 3985 9503
rect 4019 9469 4031 9503
rect 4246 9500 4252 9512
rect 4207 9472 4252 9500
rect 3973 9463 4031 9469
rect 3602 9324 3608 9376
rect 3660 9364 3666 9376
rect 3988 9364 4016 9463
rect 4246 9460 4252 9472
rect 4304 9460 4310 9512
rect 12710 9460 12716 9512
rect 12768 9500 12774 9512
rect 13832 9500 13860 9531
rect 12768 9472 13860 9500
rect 12768 9460 12774 9472
rect 5534 9432 5540 9444
rect 5276 9404 5540 9432
rect 5276 9364 5304 9404
rect 5534 9392 5540 9404
rect 5592 9432 5598 9444
rect 6454 9432 6460 9444
rect 5592 9404 6460 9432
rect 5592 9392 5598 9404
rect 6454 9392 6460 9404
rect 6512 9392 6518 9444
rect 3660 9336 5304 9364
rect 5721 9367 5779 9373
rect 3660 9324 3666 9336
rect 5721 9333 5733 9367
rect 5767 9364 5779 9367
rect 11790 9364 11796 9376
rect 5767 9336 11796 9364
rect 5767 9333 5779 9336
rect 5721 9327 5779 9333
rect 11790 9324 11796 9336
rect 11848 9324 11854 9376
rect 1104 9274 34868 9296
rect 1104 9222 5174 9274
rect 5226 9222 5238 9274
rect 5290 9222 5302 9274
rect 5354 9222 5366 9274
rect 5418 9222 5430 9274
rect 5482 9222 13622 9274
rect 13674 9222 13686 9274
rect 13738 9222 13750 9274
rect 13802 9222 13814 9274
rect 13866 9222 13878 9274
rect 13930 9222 22070 9274
rect 22122 9222 22134 9274
rect 22186 9222 22198 9274
rect 22250 9222 22262 9274
rect 22314 9222 22326 9274
rect 22378 9222 30518 9274
rect 30570 9222 30582 9274
rect 30634 9222 30646 9274
rect 30698 9222 30710 9274
rect 30762 9222 30774 9274
rect 30826 9222 34868 9274
rect 1104 9200 34868 9222
rect 4246 9120 4252 9172
rect 4304 9160 4310 9172
rect 10870 9160 10876 9172
rect 4304 9132 10876 9160
rect 4304 9120 4310 9132
rect 10870 9120 10876 9132
rect 10928 9120 10934 9172
rect 27890 9120 27896 9172
rect 27948 9160 27954 9172
rect 28077 9163 28135 9169
rect 28077 9160 28089 9163
rect 27948 9132 28089 9160
rect 27948 9120 27954 9132
rect 28077 9129 28089 9132
rect 28123 9129 28135 9163
rect 28077 9123 28135 9129
rect 12710 9024 12716 9036
rect 12671 8996 12716 9024
rect 12710 8984 12716 8996
rect 12768 8984 12774 9036
rect 21266 8984 21272 9036
rect 21324 9024 21330 9036
rect 21726 9024 21732 9036
rect 21324 8996 21732 9024
rect 21324 8984 21330 8996
rect 21726 8984 21732 8996
rect 21784 8984 21790 9036
rect 11790 8916 11796 8968
rect 11848 8956 11854 8968
rect 12345 8959 12403 8965
rect 12345 8956 12357 8959
rect 11848 8928 12357 8956
rect 11848 8916 11854 8928
rect 12345 8925 12357 8928
rect 12391 8925 12403 8959
rect 12618 8956 12624 8968
rect 12579 8928 12624 8956
rect 12345 8919 12403 8925
rect 12618 8916 12624 8928
rect 12676 8916 12682 8968
rect 21910 8916 21916 8968
rect 21968 8956 21974 8968
rect 22005 8959 22063 8965
rect 22005 8956 22017 8959
rect 21968 8928 22017 8956
rect 21968 8916 21974 8928
rect 22005 8925 22017 8928
rect 22051 8925 22063 8959
rect 22830 8956 22836 8968
rect 22791 8928 22836 8956
rect 22005 8919 22063 8925
rect 22830 8916 22836 8928
rect 22888 8956 22894 8968
rect 26694 8956 26700 8968
rect 22888 8928 26700 8956
rect 22888 8916 22894 8928
rect 26694 8916 26700 8928
rect 26752 8916 26758 8968
rect 28092 8956 28120 9123
rect 28629 8959 28687 8965
rect 28629 8956 28641 8959
rect 28092 8928 28641 8956
rect 28629 8925 28641 8928
rect 28675 8925 28687 8959
rect 33870 8956 33876 8968
rect 33831 8928 33876 8956
rect 28629 8919 28687 8925
rect 33870 8916 33876 8928
rect 33928 8916 33934 8968
rect 28718 8820 28724 8832
rect 28679 8792 28724 8820
rect 28718 8780 28724 8792
rect 28776 8780 28782 8832
rect 34054 8820 34060 8832
rect 34015 8792 34060 8820
rect 34054 8780 34060 8792
rect 34112 8780 34118 8832
rect 1104 8730 34868 8752
rect 1104 8678 9398 8730
rect 9450 8678 9462 8730
rect 9514 8678 9526 8730
rect 9578 8678 9590 8730
rect 9642 8678 9654 8730
rect 9706 8678 17846 8730
rect 17898 8678 17910 8730
rect 17962 8678 17974 8730
rect 18026 8678 18038 8730
rect 18090 8678 18102 8730
rect 18154 8678 26294 8730
rect 26346 8678 26358 8730
rect 26410 8678 26422 8730
rect 26474 8678 26486 8730
rect 26538 8678 26550 8730
rect 26602 8678 34868 8730
rect 1104 8656 34868 8678
rect 14274 8616 14280 8628
rect 14235 8588 14280 8616
rect 14274 8576 14280 8588
rect 14332 8576 14338 8628
rect 28718 8508 28724 8560
rect 28776 8508 28782 8560
rect 11790 8480 11796 8492
rect 11751 8452 11796 8480
rect 11790 8440 11796 8452
rect 11848 8440 11854 8492
rect 12618 8440 12624 8492
rect 12676 8480 12682 8492
rect 13538 8480 13544 8492
rect 12676 8452 13544 8480
rect 12676 8440 12682 8452
rect 13538 8440 13544 8452
rect 13596 8480 13602 8492
rect 14185 8483 14243 8489
rect 14185 8480 14197 8483
rect 13596 8452 14197 8480
rect 13596 8440 13602 8452
rect 14185 8449 14197 8452
rect 14231 8449 14243 8483
rect 14185 8443 14243 8449
rect 14369 8483 14427 8489
rect 14369 8449 14381 8483
rect 14415 8449 14427 8483
rect 27798 8480 27804 8492
rect 27759 8452 27804 8480
rect 14369 8443 14427 8449
rect 11974 8372 11980 8424
rect 12032 8412 12038 8424
rect 12069 8415 12127 8421
rect 12069 8412 12081 8415
rect 12032 8384 12081 8412
rect 12032 8372 12038 8384
rect 12069 8381 12081 8384
rect 12115 8412 12127 8415
rect 14384 8412 14412 8443
rect 27798 8440 27804 8452
rect 27856 8440 27862 8492
rect 28074 8412 28080 8424
rect 12115 8384 14412 8412
rect 28035 8384 28080 8412
rect 12115 8381 12127 8384
rect 12069 8375 12127 8381
rect 28074 8372 28080 8384
rect 28132 8372 28138 8424
rect 29549 8347 29607 8353
rect 29549 8313 29561 8347
rect 29595 8344 29607 8347
rect 31478 8344 31484 8356
rect 29595 8316 31484 8344
rect 29595 8313 29607 8316
rect 29549 8307 29607 8313
rect 27338 8236 27344 8288
rect 27396 8276 27402 8288
rect 29564 8276 29592 8307
rect 31478 8304 31484 8316
rect 31536 8304 31542 8356
rect 27396 8248 29592 8276
rect 27396 8236 27402 8248
rect 1104 8186 34868 8208
rect 1104 8134 5174 8186
rect 5226 8134 5238 8186
rect 5290 8134 5302 8186
rect 5354 8134 5366 8186
rect 5418 8134 5430 8186
rect 5482 8134 13622 8186
rect 13674 8134 13686 8186
rect 13738 8134 13750 8186
rect 13802 8134 13814 8186
rect 13866 8134 13878 8186
rect 13930 8134 22070 8186
rect 22122 8134 22134 8186
rect 22186 8134 22198 8186
rect 22250 8134 22262 8186
rect 22314 8134 22326 8186
rect 22378 8134 30518 8186
rect 30570 8134 30582 8186
rect 30634 8134 30646 8186
rect 30698 8134 30710 8186
rect 30762 8134 30774 8186
rect 30826 8134 34868 8186
rect 1104 8112 34868 8134
rect 1581 8075 1639 8081
rect 1581 8041 1593 8075
rect 1627 8072 1639 8075
rect 5718 8072 5724 8084
rect 1627 8044 5724 8072
rect 1627 8041 1639 8044
rect 1581 8035 1639 8041
rect 5718 8032 5724 8044
rect 5776 8032 5782 8084
rect 10870 8072 10876 8084
rect 10831 8044 10876 8072
rect 10870 8032 10876 8044
rect 10928 8032 10934 8084
rect 11793 8075 11851 8081
rect 11793 8041 11805 8075
rect 11839 8072 11851 8075
rect 12618 8072 12624 8084
rect 11839 8044 12624 8072
rect 11839 8041 11851 8044
rect 11793 8035 11851 8041
rect 12618 8032 12624 8044
rect 12676 8032 12682 8084
rect 27433 8075 27491 8081
rect 27433 8041 27445 8075
rect 27479 8072 27491 8075
rect 28074 8072 28080 8084
rect 27479 8044 28080 8072
rect 27479 8041 27491 8044
rect 27433 8035 27491 8041
rect 28074 8032 28080 8044
rect 28132 8032 28138 8084
rect 32401 8075 32459 8081
rect 32401 8041 32413 8075
rect 32447 8072 32459 8075
rect 33870 8072 33876 8084
rect 32447 8044 33876 8072
rect 32447 8041 32459 8044
rect 32401 8035 32459 8041
rect 33870 8032 33876 8044
rect 33928 8032 33934 8084
rect 26694 7964 26700 8016
rect 26752 8004 26758 8016
rect 30374 8004 30380 8016
rect 26752 7976 30380 8004
rect 26752 7964 26758 7976
rect 30374 7964 30380 7976
rect 30432 7964 30438 8016
rect 11790 7936 11796 7948
rect 11440 7908 11796 7936
rect 1394 7868 1400 7880
rect 1355 7840 1400 7868
rect 1394 7828 1400 7840
rect 1452 7828 1458 7880
rect 10781 7871 10839 7877
rect 10781 7837 10793 7871
rect 10827 7837 10839 7871
rect 10962 7868 10968 7880
rect 10923 7840 10968 7868
rect 10781 7831 10839 7837
rect 10796 7800 10824 7831
rect 10962 7828 10968 7840
rect 11020 7828 11026 7880
rect 11440 7877 11468 7908
rect 11790 7896 11796 7908
rect 11848 7896 11854 7948
rect 19981 7939 20039 7945
rect 19981 7905 19993 7939
rect 20027 7936 20039 7939
rect 20254 7936 20260 7948
rect 20027 7908 20260 7936
rect 20027 7905 20039 7908
rect 19981 7899 20039 7905
rect 20254 7896 20260 7908
rect 20312 7896 20318 7948
rect 21269 7939 21327 7945
rect 21269 7905 21281 7939
rect 21315 7936 21327 7939
rect 21910 7936 21916 7948
rect 21315 7908 21916 7936
rect 21315 7905 21327 7908
rect 21269 7899 21327 7905
rect 21910 7896 21916 7908
rect 21968 7936 21974 7948
rect 21968 7908 22140 7936
rect 21968 7896 21974 7908
rect 11425 7871 11483 7877
rect 11425 7837 11437 7871
rect 11471 7837 11483 7871
rect 11698 7868 11704 7880
rect 11659 7840 11704 7868
rect 11425 7831 11483 7837
rect 11698 7828 11704 7840
rect 11756 7828 11762 7880
rect 19334 7828 19340 7880
rect 19392 7868 19398 7880
rect 19705 7871 19763 7877
rect 19705 7868 19717 7871
rect 19392 7840 19717 7868
rect 19392 7828 19398 7840
rect 19705 7837 19717 7840
rect 19751 7837 19763 7871
rect 19705 7831 19763 7837
rect 19794 7828 19800 7880
rect 19852 7868 19858 7880
rect 19852 7840 19897 7868
rect 19852 7828 19858 7840
rect 20806 7828 20812 7880
rect 20864 7868 20870 7880
rect 22112 7877 22140 7908
rect 21177 7871 21235 7877
rect 21177 7868 21189 7871
rect 20864 7840 21189 7868
rect 20864 7828 20870 7840
rect 21177 7837 21189 7840
rect 21223 7837 21235 7871
rect 21177 7831 21235 7837
rect 22097 7871 22155 7877
rect 22097 7837 22109 7871
rect 22143 7837 22155 7871
rect 22097 7831 22155 7837
rect 27249 7871 27307 7877
rect 27249 7837 27261 7871
rect 27295 7868 27307 7871
rect 27706 7868 27712 7880
rect 27295 7840 27712 7868
rect 27295 7837 27307 7840
rect 27249 7831 27307 7837
rect 27706 7828 27712 7840
rect 27764 7828 27770 7880
rect 31389 7871 31447 7877
rect 31389 7837 31401 7871
rect 31435 7837 31447 7871
rect 31662 7868 31668 7880
rect 31623 7840 31668 7868
rect 31389 7831 31447 7837
rect 11790 7800 11796 7812
rect 10796 7772 11796 7800
rect 11790 7760 11796 7772
rect 11848 7760 11854 7812
rect 19981 7803 20039 7809
rect 19981 7769 19993 7803
rect 20027 7800 20039 7803
rect 20990 7800 20996 7812
rect 20027 7772 20996 7800
rect 20027 7769 20039 7772
rect 19981 7763 20039 7769
rect 20990 7760 20996 7772
rect 21048 7800 21054 7812
rect 21913 7803 21971 7809
rect 21913 7800 21925 7803
rect 21048 7772 21925 7800
rect 21048 7760 21054 7772
rect 21913 7769 21925 7772
rect 21959 7769 21971 7803
rect 31404 7800 31432 7831
rect 31662 7828 31668 7840
rect 31720 7828 31726 7880
rect 32122 7800 32128 7812
rect 31404 7772 32128 7800
rect 21913 7763 21971 7769
rect 32122 7760 32128 7772
rect 32180 7760 32186 7812
rect 11977 7735 12035 7741
rect 11977 7701 11989 7735
rect 12023 7732 12035 7735
rect 12342 7732 12348 7744
rect 12023 7704 12348 7732
rect 12023 7701 12035 7704
rect 11977 7695 12035 7701
rect 12342 7692 12348 7704
rect 12400 7692 12406 7744
rect 22281 7735 22339 7741
rect 22281 7701 22293 7735
rect 22327 7732 22339 7735
rect 24762 7732 24768 7744
rect 22327 7704 24768 7732
rect 22327 7701 22339 7704
rect 22281 7695 22339 7701
rect 24762 7692 24768 7704
rect 24820 7692 24826 7744
rect 1104 7642 34868 7664
rect 1104 7590 9398 7642
rect 9450 7590 9462 7642
rect 9514 7590 9526 7642
rect 9578 7590 9590 7642
rect 9642 7590 9654 7642
rect 9706 7590 17846 7642
rect 17898 7590 17910 7642
rect 17962 7590 17974 7642
rect 18026 7590 18038 7642
rect 18090 7590 18102 7642
rect 18154 7590 26294 7642
rect 26346 7590 26358 7642
rect 26410 7590 26422 7642
rect 26474 7590 26486 7642
rect 26538 7590 26550 7642
rect 26602 7590 34868 7642
rect 1104 7568 34868 7590
rect 1394 7528 1400 7540
rect 1355 7500 1400 7528
rect 1394 7488 1400 7500
rect 1452 7488 1458 7540
rect 10962 7488 10968 7540
rect 11020 7528 11026 7540
rect 12161 7531 12219 7537
rect 12161 7528 12173 7531
rect 11020 7500 12173 7528
rect 11020 7488 11026 7500
rect 12161 7497 12173 7500
rect 12207 7497 12219 7531
rect 12161 7491 12219 7497
rect 26421 7531 26479 7537
rect 26421 7497 26433 7531
rect 26467 7528 26479 7531
rect 26694 7528 26700 7540
rect 26467 7500 26700 7528
rect 26467 7497 26479 7500
rect 26421 7491 26479 7497
rect 26694 7488 26700 7500
rect 26752 7488 26758 7540
rect 27338 7528 27344 7540
rect 27299 7500 27344 7528
rect 27338 7488 27344 7500
rect 27396 7488 27402 7540
rect 27706 7528 27712 7540
rect 27667 7500 27712 7528
rect 27706 7488 27712 7500
rect 27764 7488 27770 7540
rect 4890 7420 4896 7472
rect 4948 7420 4954 7472
rect 3602 7392 3608 7404
rect 3563 7364 3608 7392
rect 3602 7352 3608 7364
rect 3660 7352 3666 7404
rect 12342 7392 12348 7404
rect 12303 7364 12348 7392
rect 12342 7352 12348 7364
rect 12400 7352 12406 7404
rect 12437 7395 12495 7401
rect 12437 7361 12449 7395
rect 12483 7392 12495 7395
rect 12526 7392 12532 7404
rect 12483 7364 12532 7392
rect 12483 7361 12495 7364
rect 12437 7355 12495 7361
rect 12526 7352 12532 7364
rect 12584 7352 12590 7404
rect 12618 7352 12624 7404
rect 12676 7392 12682 7404
rect 12713 7395 12771 7401
rect 12713 7392 12725 7395
rect 12676 7364 12725 7392
rect 12676 7352 12682 7364
rect 12713 7361 12725 7364
rect 12759 7361 12771 7395
rect 12713 7355 12771 7361
rect 14274 7352 14280 7404
rect 14332 7392 14338 7404
rect 14553 7395 14611 7401
rect 14553 7392 14565 7395
rect 14332 7364 14565 7392
rect 14332 7352 14338 7364
rect 14553 7361 14565 7364
rect 14599 7361 14611 7395
rect 14734 7392 14740 7404
rect 14695 7364 14740 7392
rect 14553 7355 14611 7361
rect 14734 7352 14740 7364
rect 14792 7352 14798 7404
rect 3881 7327 3939 7333
rect 3881 7293 3893 7327
rect 3927 7324 3939 7327
rect 5626 7324 5632 7336
rect 3927 7296 5632 7324
rect 3927 7293 3939 7296
rect 3881 7287 3939 7293
rect 5626 7284 5632 7296
rect 5684 7284 5690 7336
rect 26694 7284 26700 7336
rect 26752 7324 26758 7336
rect 27065 7327 27123 7333
rect 27065 7324 27077 7327
rect 26752 7296 27077 7324
rect 26752 7284 26758 7296
rect 27065 7293 27077 7296
rect 27111 7293 27123 7327
rect 27246 7324 27252 7336
rect 27207 7296 27252 7324
rect 27065 7287 27123 7293
rect 27246 7284 27252 7296
rect 27304 7284 27310 7336
rect 12621 7259 12679 7265
rect 12621 7225 12633 7259
rect 12667 7256 12679 7259
rect 12710 7256 12716 7268
rect 12667 7228 12716 7256
rect 12667 7225 12679 7228
rect 12621 7219 12679 7225
rect 12710 7216 12716 7228
rect 12768 7256 12774 7268
rect 19794 7256 19800 7268
rect 12768 7228 19800 7256
rect 12768 7216 12774 7228
rect 19794 7216 19800 7228
rect 19852 7256 19858 7268
rect 20346 7256 20352 7268
rect 19852 7228 20352 7256
rect 19852 7216 19858 7228
rect 20346 7216 20352 7228
rect 20404 7216 20410 7268
rect 5353 7191 5411 7197
rect 5353 7157 5365 7191
rect 5399 7188 5411 7191
rect 6178 7188 6184 7200
rect 5399 7160 6184 7188
rect 5399 7157 5411 7160
rect 5353 7151 5411 7157
rect 6178 7148 6184 7160
rect 6236 7148 6242 7200
rect 14645 7191 14703 7197
rect 14645 7157 14657 7191
rect 14691 7188 14703 7191
rect 20806 7188 20812 7200
rect 14691 7160 20812 7188
rect 14691 7157 14703 7160
rect 14645 7151 14703 7157
rect 20806 7148 20812 7160
rect 20864 7148 20870 7200
rect 1104 7098 34868 7120
rect 1104 7046 5174 7098
rect 5226 7046 5238 7098
rect 5290 7046 5302 7098
rect 5354 7046 5366 7098
rect 5418 7046 5430 7098
rect 5482 7046 13622 7098
rect 13674 7046 13686 7098
rect 13738 7046 13750 7098
rect 13802 7046 13814 7098
rect 13866 7046 13878 7098
rect 13930 7046 22070 7098
rect 22122 7046 22134 7098
rect 22186 7046 22198 7098
rect 22250 7046 22262 7098
rect 22314 7046 22326 7098
rect 22378 7046 30518 7098
rect 30570 7046 30582 7098
rect 30634 7046 30646 7098
rect 30698 7046 30710 7098
rect 30762 7046 30774 7098
rect 30826 7046 34868 7098
rect 1104 7024 34868 7046
rect 5534 6944 5540 6996
rect 5592 6944 5598 6996
rect 11977 6987 12035 6993
rect 11977 6953 11989 6987
rect 12023 6984 12035 6987
rect 12250 6984 12256 6996
rect 12023 6956 12256 6984
rect 12023 6953 12035 6956
rect 11977 6947 12035 6953
rect 12250 6944 12256 6956
rect 12308 6944 12314 6996
rect 12342 6944 12348 6996
rect 12400 6984 12406 6996
rect 20254 6984 20260 6996
rect 12400 6956 20260 6984
rect 12400 6944 12406 6956
rect 20254 6944 20260 6956
rect 20312 6944 20318 6996
rect 20806 6984 20812 6996
rect 20767 6956 20812 6984
rect 20806 6944 20812 6956
rect 20864 6944 20870 6996
rect 5552 6860 5580 6944
rect 5626 6876 5632 6928
rect 5684 6916 5690 6928
rect 11885 6919 11943 6925
rect 11885 6916 11897 6919
rect 5684 6888 11897 6916
rect 5684 6876 5690 6888
rect 11885 6885 11897 6888
rect 11931 6885 11943 6919
rect 11885 6879 11943 6885
rect 20993 6919 21051 6925
rect 20993 6885 21005 6919
rect 21039 6916 21051 6919
rect 21039 6888 21956 6916
rect 21039 6885 21051 6888
rect 20993 6879 21051 6885
rect 4709 6851 4767 6857
rect 4709 6817 4721 6851
rect 4755 6848 4767 6851
rect 4890 6848 4896 6860
rect 4755 6820 4896 6848
rect 4755 6817 4767 6820
rect 4709 6811 4767 6817
rect 4890 6808 4896 6820
rect 4948 6808 4954 6860
rect 5534 6808 5540 6860
rect 5592 6808 5598 6860
rect 12115 6851 12173 6857
rect 12115 6817 12127 6851
rect 12161 6848 12173 6851
rect 12342 6848 12348 6860
rect 12161 6820 12348 6848
rect 12161 6817 12173 6820
rect 12115 6811 12173 6817
rect 12342 6808 12348 6820
rect 12400 6848 12406 6860
rect 20073 6851 20131 6857
rect 12400 6820 16574 6848
rect 12400 6808 12406 6820
rect 4617 6783 4675 6789
rect 4617 6749 4629 6783
rect 4663 6780 4675 6783
rect 4798 6780 4804 6792
rect 4663 6752 4804 6780
rect 4663 6749 4675 6752
rect 4617 6743 4675 6749
rect 4798 6740 4804 6752
rect 4856 6740 4862 6792
rect 11790 6780 11796 6792
rect 11751 6752 11796 6780
rect 11790 6740 11796 6752
rect 11848 6740 11854 6792
rect 11974 6740 11980 6792
rect 12032 6780 12038 6792
rect 12253 6783 12311 6789
rect 12253 6780 12265 6783
rect 12032 6752 12265 6780
rect 12032 6740 12038 6752
rect 12253 6749 12265 6752
rect 12299 6749 12311 6783
rect 16546 6780 16574 6820
rect 20073 6817 20085 6851
rect 20119 6848 20131 6851
rect 21928 6848 21956 6888
rect 20119 6820 21772 6848
rect 21928 6820 22094 6848
rect 20119 6817 20131 6820
rect 20073 6811 20131 6817
rect 19981 6783 20039 6789
rect 19981 6780 19993 6783
rect 16546 6752 19993 6780
rect 12253 6743 12311 6749
rect 19981 6749 19993 6752
rect 20027 6749 20039 6783
rect 20162 6780 20168 6792
rect 20123 6752 20168 6780
rect 19981 6743 20039 6749
rect 20162 6740 20168 6752
rect 20220 6740 20226 6792
rect 20254 6740 20260 6792
rect 20312 6780 20318 6792
rect 21453 6783 21511 6789
rect 21453 6780 21465 6783
rect 20312 6752 21465 6780
rect 20312 6740 20318 6752
rect 21453 6749 21465 6752
rect 21499 6749 21511 6783
rect 21637 6783 21695 6789
rect 21637 6780 21649 6783
rect 21453 6743 21511 6749
rect 21560 6752 21649 6780
rect 20180 6712 20208 6740
rect 20625 6715 20683 6721
rect 20625 6712 20637 6715
rect 20180 6684 20637 6712
rect 20625 6681 20637 6684
rect 20671 6681 20683 6715
rect 20625 6675 20683 6681
rect 5534 6644 5540 6656
rect 5495 6616 5540 6644
rect 5534 6604 5540 6616
rect 5592 6604 5598 6656
rect 20346 6604 20352 6656
rect 20404 6644 20410 6656
rect 20825 6647 20883 6653
rect 20825 6644 20837 6647
rect 20404 6616 20837 6644
rect 20404 6604 20410 6616
rect 20825 6613 20837 6616
rect 20871 6644 20883 6647
rect 21560 6644 21588 6752
rect 21637 6749 21649 6752
rect 21683 6749 21695 6783
rect 21637 6743 21695 6749
rect 21744 6712 21772 6820
rect 22066 6780 22094 6820
rect 30377 6783 30435 6789
rect 30377 6780 30389 6783
rect 22066 6752 30389 6780
rect 30377 6749 30389 6752
rect 30423 6749 30435 6783
rect 30377 6743 30435 6749
rect 33134 6740 33140 6792
rect 33192 6780 33198 6792
rect 33873 6783 33931 6789
rect 33873 6780 33885 6783
rect 33192 6752 33885 6780
rect 33192 6740 33198 6752
rect 33873 6749 33885 6752
rect 33919 6749 33931 6783
rect 33873 6743 33931 6749
rect 31662 6712 31668 6724
rect 21744 6684 31668 6712
rect 31662 6672 31668 6684
rect 31720 6672 31726 6724
rect 20871 6616 21588 6644
rect 21637 6647 21695 6653
rect 20871 6613 20883 6616
rect 20825 6607 20883 6613
rect 21637 6613 21649 6647
rect 21683 6644 21695 6647
rect 23198 6644 23204 6656
rect 21683 6616 23204 6644
rect 21683 6613 21695 6616
rect 21637 6607 21695 6613
rect 23198 6604 23204 6616
rect 23256 6604 23262 6656
rect 30558 6644 30564 6656
rect 30519 6616 30564 6644
rect 30558 6604 30564 6616
rect 30616 6604 30622 6656
rect 34054 6644 34060 6656
rect 34015 6616 34060 6644
rect 34054 6604 34060 6616
rect 34112 6604 34118 6656
rect 1104 6554 34868 6576
rect 1104 6502 9398 6554
rect 9450 6502 9462 6554
rect 9514 6502 9526 6554
rect 9578 6502 9590 6554
rect 9642 6502 9654 6554
rect 9706 6502 17846 6554
rect 17898 6502 17910 6554
rect 17962 6502 17974 6554
rect 18026 6502 18038 6554
rect 18090 6502 18102 6554
rect 18154 6502 26294 6554
rect 26346 6502 26358 6554
rect 26410 6502 26422 6554
rect 26474 6502 26486 6554
rect 26538 6502 26550 6554
rect 26602 6502 34868 6554
rect 1104 6480 34868 6502
rect 4798 6400 4804 6452
rect 4856 6440 4862 6452
rect 4893 6443 4951 6449
rect 4893 6440 4905 6443
rect 4856 6412 4905 6440
rect 4856 6400 4862 6412
rect 4893 6409 4905 6412
rect 4939 6409 4951 6443
rect 12250 6440 12256 6452
rect 12211 6412 12256 6440
rect 4893 6403 4951 6409
rect 12250 6400 12256 6412
rect 12308 6400 12314 6452
rect 33134 6440 33140 6452
rect 33095 6412 33140 6440
rect 33134 6400 33140 6412
rect 33192 6400 33198 6452
rect 12437 6307 12495 6313
rect 12437 6273 12449 6307
rect 12483 6304 12495 6307
rect 12526 6304 12532 6316
rect 12483 6276 12532 6304
rect 12483 6273 12495 6276
rect 12437 6267 12495 6273
rect 12526 6264 12532 6276
rect 12584 6264 12590 6316
rect 24762 6264 24768 6316
rect 24820 6304 24826 6316
rect 28077 6307 28135 6313
rect 28077 6304 28089 6307
rect 24820 6276 28089 6304
rect 24820 6264 24826 6276
rect 28077 6273 28089 6276
rect 28123 6273 28135 6307
rect 28077 6267 28135 6273
rect 30558 6264 30564 6316
rect 30616 6304 30622 6316
rect 32401 6307 32459 6313
rect 32401 6304 32413 6307
rect 30616 6276 32413 6304
rect 30616 6264 30622 6276
rect 32401 6273 32413 6276
rect 32447 6273 32459 6307
rect 32401 6267 32459 6273
rect 12621 6239 12679 6245
rect 12621 6236 12633 6239
rect 12452 6208 12633 6236
rect 12452 6180 12480 6208
rect 12621 6205 12633 6208
rect 12667 6205 12679 6239
rect 32122 6236 32128 6248
rect 32083 6208 32128 6236
rect 12621 6199 12679 6205
rect 32122 6196 32128 6208
rect 32180 6196 32186 6248
rect 12434 6128 12440 6180
rect 12492 6128 12498 6180
rect 28261 6103 28319 6109
rect 28261 6069 28273 6103
rect 28307 6100 28319 6103
rect 29822 6100 29828 6112
rect 28307 6072 29828 6100
rect 28307 6069 28319 6072
rect 28261 6063 28319 6069
rect 29822 6060 29828 6072
rect 29880 6060 29886 6112
rect 1104 6010 34868 6032
rect 1104 5958 5174 6010
rect 5226 5958 5238 6010
rect 5290 5958 5302 6010
rect 5354 5958 5366 6010
rect 5418 5958 5430 6010
rect 5482 5958 13622 6010
rect 13674 5958 13686 6010
rect 13738 5958 13750 6010
rect 13802 5958 13814 6010
rect 13866 5958 13878 6010
rect 13930 5958 22070 6010
rect 22122 5958 22134 6010
rect 22186 5958 22198 6010
rect 22250 5958 22262 6010
rect 22314 5958 22326 6010
rect 22378 5958 30518 6010
rect 30570 5958 30582 6010
rect 30634 5958 30646 6010
rect 30698 5958 30710 6010
rect 30762 5958 30774 6010
rect 30826 5958 34868 6010
rect 1104 5936 34868 5958
rect 11698 5760 11704 5772
rect 6886 5732 11704 5760
rect 4709 5695 4767 5701
rect 4709 5661 4721 5695
rect 4755 5692 4767 5695
rect 4798 5692 4804 5704
rect 4755 5664 4804 5692
rect 4755 5661 4767 5664
rect 4709 5655 4767 5661
rect 4798 5652 4804 5664
rect 4856 5692 4862 5704
rect 5169 5695 5227 5701
rect 5169 5692 5181 5695
rect 4856 5664 5181 5692
rect 4856 5652 4862 5664
rect 5169 5661 5181 5664
rect 5215 5661 5227 5695
rect 6178 5692 6184 5704
rect 6139 5664 6184 5692
rect 5169 5655 5227 5661
rect 6178 5652 6184 5664
rect 6236 5692 6242 5704
rect 6886 5692 6914 5732
rect 11698 5720 11704 5732
rect 11756 5720 11762 5772
rect 6236 5664 6914 5692
rect 11425 5695 11483 5701
rect 6236 5652 6242 5664
rect 11425 5661 11437 5695
rect 11471 5692 11483 5695
rect 12434 5692 12440 5704
rect 11471 5664 12440 5692
rect 11471 5661 11483 5664
rect 11425 5655 11483 5661
rect 12434 5652 12440 5664
rect 12492 5652 12498 5704
rect 5997 5627 6055 5633
rect 5997 5593 6009 5627
rect 6043 5624 6055 5627
rect 6270 5624 6276 5636
rect 6043 5596 6276 5624
rect 6043 5593 6055 5596
rect 5997 5587 6055 5593
rect 6270 5584 6276 5596
rect 6328 5584 6334 5636
rect 4522 5516 4528 5568
rect 4580 5556 4586 5568
rect 4617 5559 4675 5565
rect 4617 5556 4629 5559
rect 4580 5528 4629 5556
rect 4580 5516 4586 5528
rect 4617 5525 4629 5528
rect 4663 5525 4675 5559
rect 4617 5519 4675 5525
rect 6365 5559 6423 5565
rect 6365 5525 6377 5559
rect 6411 5556 6423 5559
rect 12158 5556 12164 5568
rect 6411 5528 12164 5556
rect 6411 5525 6423 5528
rect 6365 5519 6423 5525
rect 12158 5516 12164 5528
rect 12216 5516 12222 5568
rect 1104 5466 34868 5488
rect 1104 5414 9398 5466
rect 9450 5414 9462 5466
rect 9514 5414 9526 5466
rect 9578 5414 9590 5466
rect 9642 5414 9654 5466
rect 9706 5414 17846 5466
rect 17898 5414 17910 5466
rect 17962 5414 17974 5466
rect 18026 5414 18038 5466
rect 18090 5414 18102 5466
rect 18154 5414 26294 5466
rect 26346 5414 26358 5466
rect 26410 5414 26422 5466
rect 26474 5414 26486 5466
rect 26538 5414 26550 5466
rect 26602 5414 34868 5466
rect 1104 5392 34868 5414
rect 12342 5352 12348 5364
rect 12303 5324 12348 5352
rect 12342 5312 12348 5324
rect 12400 5312 12406 5364
rect 19797 5287 19855 5293
rect 19797 5253 19809 5287
rect 19843 5284 19855 5287
rect 20349 5287 20407 5293
rect 20349 5284 20361 5287
rect 19843 5256 20361 5284
rect 19843 5253 19855 5256
rect 19797 5247 19855 5253
rect 20349 5253 20361 5256
rect 20395 5284 20407 5287
rect 21726 5284 21732 5296
rect 20395 5256 21732 5284
rect 20395 5253 20407 5256
rect 20349 5247 20407 5253
rect 21726 5244 21732 5256
rect 21784 5244 21790 5296
rect 29546 5284 29552 5296
rect 22940 5256 29552 5284
rect 12253 5219 12311 5225
rect 12253 5185 12265 5219
rect 12299 5185 12311 5219
rect 12434 5216 12440 5228
rect 12395 5188 12440 5216
rect 12253 5179 12311 5185
rect 12268 5148 12296 5179
rect 12434 5176 12440 5188
rect 12492 5216 12498 5228
rect 12802 5216 12808 5228
rect 12492 5188 12808 5216
rect 12492 5176 12498 5188
rect 12802 5176 12808 5188
rect 12860 5176 12866 5228
rect 19610 5216 19616 5228
rect 19571 5188 19616 5216
rect 19610 5176 19616 5188
rect 19668 5176 19674 5228
rect 22940 5225 22968 5256
rect 29546 5244 29552 5256
rect 29604 5284 29610 5296
rect 32122 5284 32128 5296
rect 29604 5256 32128 5284
rect 29604 5244 29610 5256
rect 32122 5244 32128 5256
rect 32180 5244 32186 5296
rect 20533 5219 20591 5225
rect 20533 5185 20545 5219
rect 20579 5216 20591 5219
rect 22925 5219 22983 5225
rect 22925 5216 22937 5219
rect 20579 5188 22937 5216
rect 20579 5185 20591 5188
rect 20533 5179 20591 5185
rect 22925 5185 22937 5188
rect 22971 5185 22983 5219
rect 23198 5216 23204 5228
rect 23159 5188 23204 5216
rect 22925 5179 22983 5185
rect 23198 5176 23204 5188
rect 23256 5176 23262 5228
rect 12526 5148 12532 5160
rect 12268 5120 12532 5148
rect 12526 5108 12532 5120
rect 12584 5108 12590 5160
rect 23937 5015 23995 5021
rect 23937 4981 23949 5015
rect 23983 5012 23995 5015
rect 24578 5012 24584 5024
rect 23983 4984 24584 5012
rect 23983 4981 23995 4984
rect 23937 4975 23995 4981
rect 24578 4972 24584 4984
rect 24636 4972 24642 5024
rect 1104 4922 34868 4944
rect 1104 4870 5174 4922
rect 5226 4870 5238 4922
rect 5290 4870 5302 4922
rect 5354 4870 5366 4922
rect 5418 4870 5430 4922
rect 5482 4870 13622 4922
rect 13674 4870 13686 4922
rect 13738 4870 13750 4922
rect 13802 4870 13814 4922
rect 13866 4870 13878 4922
rect 13930 4870 22070 4922
rect 22122 4870 22134 4922
rect 22186 4870 22198 4922
rect 22250 4870 22262 4922
rect 22314 4870 22326 4922
rect 22378 4870 30518 4922
rect 30570 4870 30582 4922
rect 30634 4870 30646 4922
rect 30698 4870 30710 4922
rect 30762 4870 30774 4922
rect 30826 4870 34868 4922
rect 1104 4848 34868 4870
rect 19610 4808 19616 4820
rect 19571 4780 19616 4808
rect 19610 4768 19616 4780
rect 19668 4768 19674 4820
rect 12526 4740 12532 4752
rect 12360 4712 12532 4740
rect 12360 4613 12388 4712
rect 12526 4700 12532 4712
rect 12584 4700 12590 4752
rect 12434 4632 12440 4684
rect 12492 4672 12498 4684
rect 12618 4672 12624 4684
rect 12492 4644 12624 4672
rect 12492 4632 12498 4644
rect 12618 4632 12624 4644
rect 12676 4672 12682 4684
rect 12713 4675 12771 4681
rect 12713 4672 12725 4675
rect 12676 4644 12725 4672
rect 12676 4632 12682 4644
rect 12713 4641 12725 4644
rect 12759 4672 12771 4675
rect 19334 4672 19340 4684
rect 12759 4644 19340 4672
rect 12759 4641 12771 4644
rect 12713 4635 12771 4641
rect 12345 4607 12403 4613
rect 12345 4604 12357 4607
rect 11532 4576 12357 4604
rect 6362 4536 6368 4548
rect 6323 4508 6368 4536
rect 6362 4496 6368 4508
rect 6420 4496 6426 4548
rect 11532 4480 11560 4576
rect 12345 4573 12357 4576
rect 12391 4573 12403 4607
rect 12345 4567 12403 4573
rect 12529 4607 12587 4613
rect 12529 4573 12541 4607
rect 12575 4604 12587 4607
rect 12802 4604 12808 4616
rect 12575 4576 12808 4604
rect 12575 4573 12587 4576
rect 12529 4567 12587 4573
rect 12802 4564 12808 4576
rect 12860 4564 12866 4616
rect 17126 4564 17132 4616
rect 17184 4604 17190 4616
rect 18524 4613 18552 4644
rect 19334 4632 19340 4644
rect 19392 4632 19398 4684
rect 29546 4672 29552 4684
rect 29507 4644 29552 4672
rect 29546 4632 29552 4644
rect 29604 4632 29610 4684
rect 18325 4607 18383 4613
rect 18325 4604 18337 4607
rect 17184 4576 18337 4604
rect 17184 4564 17190 4576
rect 18325 4573 18337 4576
rect 18371 4573 18383 4607
rect 18325 4567 18383 4573
rect 18509 4607 18567 4613
rect 18509 4573 18521 4607
rect 18555 4573 18567 4607
rect 18509 4567 18567 4573
rect 19245 4607 19303 4613
rect 19245 4573 19257 4607
rect 19291 4573 19303 4607
rect 19245 4567 19303 4573
rect 19429 4607 19487 4613
rect 19429 4573 19441 4607
rect 19475 4604 19487 4607
rect 20162 4604 20168 4616
rect 19475 4576 20168 4604
rect 19475 4573 19487 4576
rect 19429 4567 19487 4573
rect 15654 4496 15660 4548
rect 15712 4536 15718 4548
rect 19260 4536 19288 4567
rect 15712 4508 19288 4536
rect 15712 4496 15718 4508
rect 6457 4471 6515 4477
rect 6457 4437 6469 4471
rect 6503 4468 6515 4471
rect 11514 4468 11520 4480
rect 6503 4440 11520 4468
rect 6503 4437 6515 4440
rect 6457 4431 6515 4437
rect 11514 4428 11520 4440
rect 11572 4428 11578 4480
rect 18509 4471 18567 4477
rect 18509 4437 18521 4471
rect 18555 4468 18567 4471
rect 19444 4468 19472 4567
rect 20162 4564 20168 4576
rect 20220 4564 20226 4616
rect 29822 4604 29828 4616
rect 29783 4576 29828 4604
rect 29822 4564 29828 4576
rect 29880 4564 29886 4616
rect 18555 4440 19472 4468
rect 30561 4471 30619 4477
rect 18555 4437 18567 4440
rect 18509 4431 18567 4437
rect 30561 4437 30573 4471
rect 30607 4468 30619 4471
rect 31570 4468 31576 4480
rect 30607 4440 31576 4468
rect 30607 4437 30619 4440
rect 30561 4431 30619 4437
rect 31570 4428 31576 4440
rect 31628 4428 31634 4480
rect 1104 4378 34868 4400
rect 1104 4326 9398 4378
rect 9450 4326 9462 4378
rect 9514 4326 9526 4378
rect 9578 4326 9590 4378
rect 9642 4326 9654 4378
rect 9706 4326 17846 4378
rect 17898 4326 17910 4378
rect 17962 4326 17974 4378
rect 18026 4326 18038 4378
rect 18090 4326 18102 4378
rect 18154 4326 26294 4378
rect 26346 4326 26358 4378
rect 26410 4326 26422 4378
rect 26474 4326 26486 4378
rect 26538 4326 26550 4378
rect 26602 4326 34868 4378
rect 1104 4304 34868 4326
rect 12802 4224 12808 4276
rect 12860 4224 12866 4276
rect 4522 4156 4528 4208
rect 4580 4156 4586 4208
rect 12618 4156 12624 4208
rect 12676 4196 12682 4208
rect 12820 4196 12848 4224
rect 12676 4168 13676 4196
rect 12676 4156 12682 4168
rect 11514 4128 11520 4140
rect 11475 4100 11520 4128
rect 11514 4088 11520 4100
rect 11572 4088 11578 4140
rect 11701 4131 11759 4137
rect 11701 4097 11713 4131
rect 11747 4128 11759 4131
rect 11974 4128 11980 4140
rect 11747 4100 11980 4128
rect 11747 4097 11759 4100
rect 11701 4091 11759 4097
rect 11974 4088 11980 4100
rect 12032 4088 12038 4140
rect 12158 4128 12164 4140
rect 12119 4100 12164 4128
rect 12158 4088 12164 4100
rect 12216 4088 12222 4140
rect 12434 4128 12440 4140
rect 12395 4100 12440 4128
rect 12434 4088 12440 4100
rect 12492 4088 12498 4140
rect 12713 4131 12771 4137
rect 12713 4097 12725 4131
rect 12759 4097 12771 4131
rect 12713 4091 12771 4097
rect 3513 4063 3571 4069
rect 3513 4029 3525 4063
rect 3559 4029 3571 4063
rect 3786 4060 3792 4072
rect 3747 4032 3792 4060
rect 3513 4023 3571 4029
rect 3528 3924 3556 4023
rect 3786 4020 3792 4032
rect 3844 4020 3850 4072
rect 5261 4063 5319 4069
rect 5261 4029 5273 4063
rect 5307 4060 5319 4063
rect 6362 4060 6368 4072
rect 5307 4032 6368 4060
rect 5307 4029 5319 4032
rect 5261 4023 5319 4029
rect 6362 4020 6368 4032
rect 6420 4020 6426 4072
rect 11790 4020 11796 4072
rect 11848 4060 11854 4072
rect 12253 4063 12311 4069
rect 12253 4060 12265 4063
rect 11848 4032 12265 4060
rect 11848 4020 11854 4032
rect 12253 4029 12265 4032
rect 12299 4029 12311 4063
rect 12728 4060 12756 4091
rect 12802 4088 12808 4140
rect 12860 4128 12866 4140
rect 13648 4137 13676 4168
rect 13173 4131 13231 4137
rect 12860 4100 12905 4128
rect 12860 4088 12866 4100
rect 13173 4097 13185 4131
rect 13219 4097 13231 4131
rect 13173 4091 13231 4097
rect 13633 4131 13691 4137
rect 13633 4097 13645 4131
rect 13679 4097 13691 4131
rect 33870 4128 33876 4140
rect 33831 4100 33876 4128
rect 13633 4091 13691 4097
rect 13188 4060 13216 4091
rect 33870 4088 33876 4100
rect 33928 4088 33934 4140
rect 13725 4063 13783 4069
rect 13725 4060 13737 4063
rect 12728 4032 12848 4060
rect 13188 4032 13737 4060
rect 12253 4023 12311 4029
rect 5534 3992 5540 4004
rect 5092 3964 5540 3992
rect 5092 3924 5120 3964
rect 5534 3952 5540 3964
rect 5592 3992 5598 4004
rect 5721 3995 5779 4001
rect 5721 3992 5733 3995
rect 5592 3964 5733 3992
rect 5592 3952 5598 3964
rect 5721 3961 5733 3964
rect 5767 3961 5779 3995
rect 5721 3955 5779 3961
rect 12710 3952 12716 4004
rect 12768 3992 12774 4004
rect 12820 3992 12848 4032
rect 13725 4029 13737 4032
rect 13771 4029 13783 4063
rect 13725 4023 13783 4029
rect 13814 4020 13820 4072
rect 13872 4060 13878 4072
rect 15381 4063 15439 4069
rect 15381 4060 15393 4063
rect 13872 4032 15393 4060
rect 13872 4020 13878 4032
rect 15381 4029 15393 4032
rect 15427 4029 15439 4063
rect 15841 4063 15899 4069
rect 15841 4060 15853 4063
rect 15381 4023 15439 4029
rect 15488 4032 15853 4060
rect 15488 3992 15516 4032
rect 15841 4029 15853 4032
rect 15887 4060 15899 4063
rect 17126 4060 17132 4072
rect 15887 4032 17132 4060
rect 15887 4029 15899 4032
rect 15841 4023 15899 4029
rect 17126 4020 17132 4032
rect 17184 4020 17190 4072
rect 15654 3992 15660 4004
rect 12768 3964 15516 3992
rect 15615 3964 15660 3992
rect 12768 3952 12774 3964
rect 15654 3952 15660 3964
rect 15712 3952 15718 4004
rect 11698 3924 11704 3936
rect 3528 3896 5120 3924
rect 11659 3896 11704 3924
rect 11698 3884 11704 3896
rect 11756 3884 11762 3936
rect 12158 3884 12164 3936
rect 12216 3924 12222 3936
rect 14734 3924 14740 3936
rect 12216 3896 14740 3924
rect 12216 3884 12222 3896
rect 14734 3884 14740 3896
rect 14792 3884 14798 3936
rect 24578 3884 24584 3936
rect 24636 3924 24642 3936
rect 31662 3924 31668 3936
rect 24636 3896 31668 3924
rect 24636 3884 24642 3896
rect 31662 3884 31668 3896
rect 31720 3884 31726 3936
rect 34054 3924 34060 3936
rect 34015 3896 34060 3924
rect 34054 3884 34060 3896
rect 34112 3884 34118 3936
rect 1104 3834 34868 3856
rect 1104 3782 5174 3834
rect 5226 3782 5238 3834
rect 5290 3782 5302 3834
rect 5354 3782 5366 3834
rect 5418 3782 5430 3834
rect 5482 3782 13622 3834
rect 13674 3782 13686 3834
rect 13738 3782 13750 3834
rect 13802 3782 13814 3834
rect 13866 3782 13878 3834
rect 13930 3782 22070 3834
rect 22122 3782 22134 3834
rect 22186 3782 22198 3834
rect 22250 3782 22262 3834
rect 22314 3782 22326 3834
rect 22378 3782 30518 3834
rect 30570 3782 30582 3834
rect 30634 3782 30646 3834
rect 30698 3782 30710 3834
rect 30762 3782 30774 3834
rect 30826 3782 34868 3834
rect 1104 3760 34868 3782
rect 3786 3680 3792 3732
rect 3844 3720 3850 3732
rect 12897 3723 12955 3729
rect 12897 3720 12909 3723
rect 3844 3692 12909 3720
rect 3844 3680 3850 3692
rect 12897 3689 12909 3692
rect 12943 3689 12955 3723
rect 12897 3683 12955 3689
rect 21634 3680 21640 3732
rect 21692 3720 21698 3732
rect 21729 3723 21787 3729
rect 21729 3720 21741 3723
rect 21692 3692 21741 3720
rect 21692 3680 21698 3692
rect 21729 3689 21741 3692
rect 21775 3689 21787 3723
rect 21729 3683 21787 3689
rect 22557 3723 22615 3729
rect 22557 3689 22569 3723
rect 22603 3720 22615 3723
rect 24578 3720 24584 3732
rect 22603 3692 24584 3720
rect 22603 3689 22615 3692
rect 22557 3683 22615 3689
rect 24578 3680 24584 3692
rect 24636 3680 24642 3732
rect 27246 3720 27252 3732
rect 24688 3692 27252 3720
rect 11974 3612 11980 3664
rect 12032 3652 12038 3664
rect 15654 3652 15660 3664
rect 12032 3624 15660 3652
rect 12032 3612 12038 3624
rect 15654 3612 15660 3624
rect 15712 3612 15718 3664
rect 23658 3652 23664 3664
rect 23571 3624 23664 3652
rect 23658 3612 23664 3624
rect 23716 3652 23722 3664
rect 24688 3652 24716 3692
rect 27246 3680 27252 3692
rect 27304 3680 27310 3732
rect 29638 3720 29644 3732
rect 29599 3692 29644 3720
rect 29638 3680 29644 3692
rect 29696 3680 29702 3732
rect 31570 3720 31576 3732
rect 29748 3692 31576 3720
rect 23716 3624 24716 3652
rect 24765 3655 24823 3661
rect 23716 3612 23722 3624
rect 24765 3621 24777 3655
rect 24811 3621 24823 3655
rect 24765 3615 24823 3621
rect 5074 3584 5080 3596
rect 5035 3556 5080 3584
rect 5074 3544 5080 3556
rect 5132 3544 5138 3596
rect 5537 3587 5595 3593
rect 5537 3553 5549 3587
rect 5583 3584 5595 3587
rect 12158 3584 12164 3596
rect 5583 3556 12164 3584
rect 5583 3553 5595 3556
rect 5537 3547 5595 3553
rect 12158 3544 12164 3556
rect 12216 3584 12222 3596
rect 12802 3584 12808 3596
rect 12216 3556 12808 3584
rect 12216 3544 12222 3556
rect 12802 3544 12808 3556
rect 12860 3544 12866 3596
rect 22925 3587 22983 3593
rect 22925 3553 22937 3587
rect 22971 3584 22983 3587
rect 22971 3556 24440 3584
rect 22971 3553 22983 3556
rect 22925 3547 22983 3553
rect 5169 3519 5227 3525
rect 5169 3485 5181 3519
rect 5215 3516 5227 3519
rect 6822 3516 6828 3528
rect 5215 3488 6828 3516
rect 5215 3485 5227 3488
rect 5169 3479 5227 3485
rect 6822 3476 6828 3488
rect 6880 3476 6886 3528
rect 11698 3476 11704 3528
rect 11756 3516 11762 3528
rect 12345 3519 12403 3525
rect 12345 3516 12357 3519
rect 11756 3488 12357 3516
rect 11756 3476 11762 3488
rect 12345 3485 12357 3488
rect 12391 3485 12403 3519
rect 12710 3516 12716 3528
rect 12671 3488 12716 3516
rect 12345 3479 12403 3485
rect 12710 3476 12716 3488
rect 12768 3476 12774 3528
rect 21913 3519 21971 3525
rect 21913 3485 21925 3519
rect 21959 3516 21971 3519
rect 21959 3488 22094 3516
rect 21959 3485 21971 3488
rect 21913 3479 21971 3485
rect 12526 3448 12532 3460
rect 12487 3420 12532 3448
rect 12526 3408 12532 3420
rect 12584 3408 12590 3460
rect 12621 3451 12679 3457
rect 12621 3417 12633 3451
rect 12667 3417 12679 3451
rect 12621 3411 12679 3417
rect 12342 3340 12348 3392
rect 12400 3380 12406 3392
rect 12636 3380 12664 3411
rect 12400 3352 12664 3380
rect 22066 3380 22094 3488
rect 23750 3476 23756 3528
rect 23808 3516 23814 3528
rect 23845 3519 23903 3525
rect 23845 3516 23857 3519
rect 23808 3488 23857 3516
rect 23808 3476 23814 3488
rect 23845 3485 23857 3488
rect 23891 3485 23903 3519
rect 23845 3479 23903 3485
rect 24412 3460 24440 3556
rect 24780 3516 24808 3615
rect 29748 3584 29776 3692
rect 31570 3680 31576 3692
rect 31628 3680 31634 3732
rect 28644 3556 29776 3584
rect 28537 3519 28595 3525
rect 28537 3516 28549 3519
rect 24780 3488 28549 3516
rect 28537 3485 28549 3488
rect 28583 3485 28595 3519
rect 28537 3479 28595 3485
rect 22554 3448 22560 3460
rect 22467 3420 22560 3448
rect 22554 3408 22560 3420
rect 22612 3448 22618 3460
rect 23382 3448 23388 3460
rect 22612 3420 23388 3448
rect 22612 3408 22618 3420
rect 23382 3408 23388 3420
rect 23440 3448 23446 3460
rect 24394 3448 24400 3460
rect 23440 3420 23796 3448
rect 24307 3420 24400 3448
rect 23440 3408 23446 3420
rect 22373 3383 22431 3389
rect 22373 3380 22385 3383
rect 22066 3352 22385 3380
rect 12400 3340 12406 3352
rect 22373 3349 22385 3352
rect 22419 3349 22431 3383
rect 23768 3380 23796 3420
rect 24394 3408 24400 3420
rect 24452 3448 24458 3460
rect 28644 3448 28672 3556
rect 30377 3519 30435 3525
rect 30377 3516 30389 3519
rect 24452 3420 28672 3448
rect 28736 3488 30389 3516
rect 24452 3408 24458 3420
rect 28736 3389 28764 3488
rect 30377 3485 30389 3488
rect 30423 3485 30435 3519
rect 30377 3479 30435 3485
rect 30653 3519 30711 3525
rect 30653 3485 30665 3519
rect 30699 3516 30711 3519
rect 30742 3516 30748 3528
rect 30699 3488 30748 3516
rect 30699 3485 30711 3488
rect 30653 3479 30711 3485
rect 30742 3476 30748 3488
rect 30800 3476 30806 3528
rect 31662 3516 31668 3528
rect 31575 3488 31668 3516
rect 31662 3476 31668 3488
rect 31720 3516 31726 3528
rect 33870 3516 33876 3528
rect 31720 3488 33876 3516
rect 31720 3476 31726 3488
rect 33870 3476 33876 3488
rect 33928 3476 33934 3528
rect 24597 3383 24655 3389
rect 24597 3380 24609 3383
rect 23768 3352 24609 3380
rect 22373 3343 22431 3349
rect 24597 3349 24609 3352
rect 24643 3349 24655 3383
rect 24597 3343 24655 3349
rect 28721 3383 28779 3389
rect 28721 3349 28733 3383
rect 28767 3349 28779 3383
rect 28721 3343 28779 3349
rect 30926 3340 30932 3392
rect 30984 3380 30990 3392
rect 31205 3383 31263 3389
rect 31205 3380 31217 3383
rect 30984 3352 31217 3380
rect 30984 3340 30990 3352
rect 31205 3349 31217 3352
rect 31251 3349 31263 3383
rect 31205 3343 31263 3349
rect 1104 3290 34868 3312
rect 1104 3238 9398 3290
rect 9450 3238 9462 3290
rect 9514 3238 9526 3290
rect 9578 3238 9590 3290
rect 9642 3238 9654 3290
rect 9706 3238 17846 3290
rect 17898 3238 17910 3290
rect 17962 3238 17974 3290
rect 18026 3238 18038 3290
rect 18090 3238 18102 3290
rect 18154 3238 26294 3290
rect 26346 3238 26358 3290
rect 26410 3238 26422 3290
rect 26474 3238 26486 3290
rect 26538 3238 26550 3290
rect 26602 3238 34868 3290
rect 1104 3216 34868 3238
rect 12526 3176 12532 3188
rect 12487 3148 12532 3176
rect 12526 3136 12532 3148
rect 12584 3136 12590 3188
rect 23750 3176 23756 3188
rect 23711 3148 23756 3176
rect 23750 3136 23756 3148
rect 23808 3136 23814 3188
rect 30742 3176 30748 3188
rect 30703 3148 30748 3176
rect 30742 3136 30748 3148
rect 30800 3136 30806 3188
rect 23569 3111 23627 3117
rect 23569 3077 23581 3111
rect 23615 3108 23627 3111
rect 24394 3108 24400 3120
rect 23615 3080 24400 3108
rect 23615 3077 23627 3080
rect 23569 3071 23627 3077
rect 24394 3068 24400 3080
rect 24452 3068 24458 3120
rect 12158 3040 12164 3052
rect 12119 3012 12164 3040
rect 12158 3000 12164 3012
rect 12216 3000 12222 3052
rect 12345 3043 12403 3049
rect 12345 3009 12357 3043
rect 12391 3040 12403 3043
rect 12618 3040 12624 3052
rect 12391 3012 12624 3040
rect 12391 3009 12403 3012
rect 12345 3003 12403 3009
rect 12618 3000 12624 3012
rect 12676 3000 12682 3052
rect 23201 3043 23259 3049
rect 23201 3009 23213 3043
rect 23247 3040 23259 3043
rect 24578 3040 24584 3052
rect 23247 3012 24584 3040
rect 23247 3009 23259 3012
rect 23201 3003 23259 3009
rect 24578 3000 24584 3012
rect 24636 3000 24642 3052
rect 30926 3040 30932 3052
rect 30887 3012 30932 3040
rect 30926 3000 30932 3012
rect 30984 3000 30990 3052
rect 1762 2836 1768 2848
rect 1723 2808 1768 2836
rect 1762 2796 1768 2808
rect 1820 2796 1826 2848
rect 12345 2839 12403 2845
rect 12345 2805 12357 2839
rect 12391 2836 12403 2839
rect 13538 2836 13544 2848
rect 12391 2808 13544 2836
rect 12391 2805 12403 2808
rect 12345 2799 12403 2805
rect 13538 2796 13544 2808
rect 13596 2796 13602 2848
rect 23382 2796 23388 2848
rect 23440 2836 23446 2848
rect 23569 2839 23627 2845
rect 23569 2836 23581 2839
rect 23440 2808 23581 2836
rect 23440 2796 23446 2808
rect 23569 2805 23581 2808
rect 23615 2805 23627 2839
rect 23569 2799 23627 2805
rect 1104 2746 34868 2768
rect 1104 2694 5174 2746
rect 5226 2694 5238 2746
rect 5290 2694 5302 2746
rect 5354 2694 5366 2746
rect 5418 2694 5430 2746
rect 5482 2694 13622 2746
rect 13674 2694 13686 2746
rect 13738 2694 13750 2746
rect 13802 2694 13814 2746
rect 13866 2694 13878 2746
rect 13930 2694 22070 2746
rect 22122 2694 22134 2746
rect 22186 2694 22198 2746
rect 22250 2694 22262 2746
rect 22314 2694 22326 2746
rect 22378 2694 30518 2746
rect 30570 2694 30582 2746
rect 30634 2694 30646 2746
rect 30698 2694 30710 2746
rect 30762 2694 30774 2746
rect 30826 2694 34868 2746
rect 1104 2672 34868 2694
rect 3142 2592 3148 2644
rect 3200 2632 3206 2644
rect 15378 2632 15384 2644
rect 3200 2604 15384 2632
rect 3200 2592 3206 2604
rect 15378 2592 15384 2604
rect 15436 2592 15442 2644
rect 2041 2567 2099 2573
rect 2041 2533 2053 2567
rect 2087 2564 2099 2567
rect 3878 2564 3884 2576
rect 2087 2536 3884 2564
rect 2087 2533 2099 2536
rect 2041 2527 2099 2533
rect 3878 2524 3884 2536
rect 3936 2524 3942 2576
rect 4525 2567 4583 2573
rect 4525 2533 4537 2567
rect 4571 2564 4583 2567
rect 5074 2564 5080 2576
rect 4571 2536 5080 2564
rect 4571 2533 4583 2536
rect 4525 2527 4583 2533
rect 5074 2524 5080 2536
rect 5132 2524 5138 2576
rect 6822 2564 6828 2576
rect 6783 2536 6828 2564
rect 6822 2524 6828 2536
rect 6880 2524 6886 2576
rect 23658 2496 23664 2508
rect 16546 2468 23664 2496
rect 1762 2388 1768 2440
rect 1820 2428 1826 2440
rect 1857 2431 1915 2437
rect 1857 2428 1869 2431
rect 1820 2400 1869 2428
rect 1820 2388 1826 2400
rect 1857 2397 1869 2400
rect 1903 2397 1915 2431
rect 1857 2391 1915 2397
rect 4246 2388 4252 2440
rect 4304 2428 4310 2440
rect 4341 2431 4399 2437
rect 4341 2428 4353 2431
rect 4304 2400 4353 2428
rect 4304 2388 4310 2400
rect 4341 2397 4353 2400
rect 4387 2428 4399 2431
rect 4985 2431 5043 2437
rect 4985 2428 4997 2431
rect 4387 2400 4997 2428
rect 4387 2397 4399 2400
rect 4341 2391 4399 2397
rect 4985 2397 4997 2400
rect 5031 2397 5043 2431
rect 4985 2391 5043 2397
rect 6914 2388 6920 2440
rect 6972 2428 6978 2440
rect 7009 2431 7067 2437
rect 7009 2428 7021 2431
rect 6972 2400 7021 2428
rect 6972 2388 6978 2400
rect 7009 2397 7021 2400
rect 7055 2428 7067 2431
rect 7469 2431 7527 2437
rect 7469 2428 7481 2431
rect 7055 2400 7481 2428
rect 7055 2397 7067 2400
rect 7009 2391 7067 2397
rect 7469 2397 7481 2400
rect 7515 2397 7527 2431
rect 7469 2391 7527 2397
rect 9214 2388 9220 2440
rect 9272 2428 9278 2440
rect 9309 2431 9367 2437
rect 9309 2428 9321 2431
rect 9272 2400 9321 2428
rect 9272 2388 9278 2400
rect 9309 2397 9321 2400
rect 9355 2428 9367 2431
rect 9953 2431 10011 2437
rect 9953 2428 9965 2431
rect 9355 2400 9965 2428
rect 9355 2397 9367 2400
rect 9309 2391 9367 2397
rect 9953 2397 9965 2400
rect 9999 2397 10011 2431
rect 9953 2391 10011 2397
rect 14553 2431 14611 2437
rect 14553 2397 14565 2431
rect 14599 2428 14611 2431
rect 16546 2428 16574 2468
rect 23658 2456 23664 2468
rect 23716 2456 23722 2508
rect 33413 2499 33471 2505
rect 33413 2465 33425 2499
rect 33459 2496 33471 2499
rect 33962 2496 33968 2508
rect 33459 2468 33968 2496
rect 33459 2465 33471 2468
rect 33413 2459 33471 2465
rect 33962 2456 33968 2468
rect 34020 2456 34026 2508
rect 14599 2400 16574 2428
rect 14599 2397 14611 2400
rect 14553 2391 14611 2397
rect 21634 2388 21640 2440
rect 21692 2428 21698 2440
rect 21821 2431 21879 2437
rect 21821 2428 21833 2431
rect 21692 2400 21833 2428
rect 21692 2388 21698 2400
rect 21821 2397 21833 2400
rect 21867 2397 21879 2431
rect 21821 2391 21879 2397
rect 29638 2388 29644 2440
rect 29696 2428 29702 2440
rect 29825 2431 29883 2437
rect 29825 2428 29837 2431
rect 29696 2400 29837 2428
rect 29696 2388 29702 2400
rect 29825 2397 29837 2400
rect 29871 2428 29883 2431
rect 30285 2431 30343 2437
rect 30285 2428 30297 2431
rect 29871 2400 30297 2428
rect 29871 2397 29883 2400
rect 29825 2391 29883 2397
rect 30285 2397 30297 2400
rect 30331 2397 30343 2431
rect 30285 2391 30343 2397
rect 31570 2388 31576 2440
rect 31628 2428 31634 2440
rect 33873 2431 33931 2437
rect 33873 2428 33885 2431
rect 31628 2400 33885 2428
rect 31628 2388 31634 2400
rect 33873 2397 33885 2400
rect 33919 2397 33931 2431
rect 33873 2391 33931 2397
rect 22554 2360 22560 2372
rect 9508 2332 22560 2360
rect 9508 2301 9536 2332
rect 22554 2320 22560 2332
rect 22612 2320 22618 2372
rect 9493 2295 9551 2301
rect 9493 2261 9505 2295
rect 9539 2261 9551 2295
rect 9493 2255 9551 2261
rect 14182 2252 14188 2304
rect 14240 2292 14246 2304
rect 14369 2295 14427 2301
rect 14369 2292 14381 2295
rect 14240 2264 14381 2292
rect 14240 2252 14246 2264
rect 14369 2261 14381 2264
rect 14415 2261 14427 2295
rect 14369 2255 14427 2261
rect 21634 2252 21640 2304
rect 21692 2292 21698 2304
rect 22005 2295 22063 2301
rect 22005 2292 22017 2295
rect 21692 2264 22017 2292
rect 21692 2252 21698 2264
rect 22005 2261 22017 2264
rect 22051 2261 22063 2295
rect 22005 2255 22063 2261
rect 29086 2252 29092 2304
rect 29144 2292 29150 2304
rect 29641 2295 29699 2301
rect 29641 2292 29653 2295
rect 29144 2264 29653 2292
rect 29144 2252 29150 2264
rect 29641 2261 29653 2264
rect 29687 2261 29699 2295
rect 34054 2292 34060 2304
rect 34015 2264 34060 2292
rect 29641 2255 29699 2261
rect 34054 2252 34060 2264
rect 34112 2252 34118 2304
rect 1104 2202 34868 2224
rect 1104 2150 9398 2202
rect 9450 2150 9462 2202
rect 9514 2150 9526 2202
rect 9578 2150 9590 2202
rect 9642 2150 9654 2202
rect 9706 2150 17846 2202
rect 17898 2150 17910 2202
rect 17962 2150 17974 2202
rect 18026 2150 18038 2202
rect 18090 2150 18102 2202
rect 18154 2150 26294 2202
rect 26346 2150 26358 2202
rect 26410 2150 26422 2202
rect 26474 2150 26486 2202
rect 26538 2150 26550 2202
rect 26602 2150 34868 2202
rect 1104 2128 34868 2150
<< via1 >>
rect 9398 17382 9450 17434
rect 9462 17382 9514 17434
rect 9526 17382 9578 17434
rect 9590 17382 9642 17434
rect 9654 17382 9706 17434
rect 17846 17382 17898 17434
rect 17910 17382 17962 17434
rect 17974 17382 18026 17434
rect 18038 17382 18090 17434
rect 18102 17382 18154 17434
rect 26294 17382 26346 17434
rect 26358 17382 26410 17434
rect 26422 17382 26474 17434
rect 26486 17382 26538 17434
rect 26550 17382 26602 17434
rect 3608 17280 3660 17332
rect 10784 17280 10836 17332
rect 18236 17280 18288 17332
rect 25136 17280 25188 17332
rect 32312 17280 32364 17332
rect 34060 17323 34112 17332
rect 34060 17289 34069 17323
rect 34069 17289 34103 17323
rect 34103 17289 34112 17323
rect 34060 17280 34112 17289
rect 1400 17187 1452 17196
rect 1400 17153 1409 17187
rect 1409 17153 1443 17187
rect 1443 17153 1452 17187
rect 1400 17144 1452 17153
rect 6828 17144 6880 17196
rect 11520 17187 11572 17196
rect 11520 17153 11529 17187
rect 11529 17153 11563 17187
rect 11563 17153 11572 17187
rect 11520 17144 11572 17153
rect 18328 17187 18380 17196
rect 18328 17153 18337 17187
rect 18337 17153 18371 17187
rect 18371 17153 18380 17187
rect 18328 17144 18380 17153
rect 25504 17187 25556 17196
rect 25504 17153 25513 17187
rect 25513 17153 25547 17187
rect 25547 17153 25556 17187
rect 25504 17144 25556 17153
rect 29920 17144 29972 17196
rect 33324 17144 33376 17196
rect 20076 17008 20128 17060
rect 33324 16983 33376 16992
rect 33324 16949 33333 16983
rect 33333 16949 33367 16983
rect 33367 16949 33376 16983
rect 33324 16940 33376 16949
rect 5174 16838 5226 16890
rect 5238 16838 5290 16890
rect 5302 16838 5354 16890
rect 5366 16838 5418 16890
rect 5430 16838 5482 16890
rect 13622 16838 13674 16890
rect 13686 16838 13738 16890
rect 13750 16838 13802 16890
rect 13814 16838 13866 16890
rect 13878 16838 13930 16890
rect 22070 16838 22122 16890
rect 22134 16838 22186 16890
rect 22198 16838 22250 16890
rect 22262 16838 22314 16890
rect 22326 16838 22378 16890
rect 30518 16838 30570 16890
rect 30582 16838 30634 16890
rect 30646 16838 30698 16890
rect 30710 16838 30762 16890
rect 30774 16838 30826 16890
rect 1400 16779 1452 16788
rect 1400 16745 1409 16779
rect 1409 16745 1443 16779
rect 1443 16745 1452 16779
rect 1400 16736 1452 16745
rect 6552 16575 6604 16584
rect 6552 16541 6561 16575
rect 6561 16541 6595 16575
rect 6595 16541 6604 16575
rect 6552 16532 6604 16541
rect 31392 16532 31444 16584
rect 7012 16396 7064 16448
rect 34060 16439 34112 16448
rect 34060 16405 34069 16439
rect 34069 16405 34103 16439
rect 34103 16405 34112 16439
rect 34060 16396 34112 16405
rect 9398 16294 9450 16346
rect 9462 16294 9514 16346
rect 9526 16294 9578 16346
rect 9590 16294 9642 16346
rect 9654 16294 9706 16346
rect 17846 16294 17898 16346
rect 17910 16294 17962 16346
rect 17974 16294 18026 16346
rect 18038 16294 18090 16346
rect 18102 16294 18154 16346
rect 26294 16294 26346 16346
rect 26358 16294 26410 16346
rect 26422 16294 26474 16346
rect 26486 16294 26538 16346
rect 26550 16294 26602 16346
rect 6920 16192 6972 16244
rect 11520 16192 11572 16244
rect 7012 16167 7064 16176
rect 7012 16133 7021 16167
rect 7021 16133 7055 16167
rect 7055 16133 7064 16167
rect 7012 16124 7064 16133
rect 8024 16124 8076 16176
rect 17776 16056 17828 16108
rect 29920 16192 29972 16244
rect 22468 16124 22520 16176
rect 25504 16124 25556 16176
rect 21916 16056 21968 16108
rect 6460 15988 6512 16040
rect 13452 15988 13504 16040
rect 18328 15988 18380 16040
rect 14372 15852 14424 15904
rect 20628 15852 20680 15904
rect 21180 15852 21232 15904
rect 29092 15895 29144 15904
rect 29092 15861 29101 15895
rect 29101 15861 29135 15895
rect 29135 15861 29144 15895
rect 29092 15852 29144 15861
rect 5174 15750 5226 15802
rect 5238 15750 5290 15802
rect 5302 15750 5354 15802
rect 5366 15750 5418 15802
rect 5430 15750 5482 15802
rect 13622 15750 13674 15802
rect 13686 15750 13738 15802
rect 13750 15750 13802 15802
rect 13814 15750 13866 15802
rect 13878 15750 13930 15802
rect 22070 15750 22122 15802
rect 22134 15750 22186 15802
rect 22198 15750 22250 15802
rect 22262 15750 22314 15802
rect 22326 15750 22378 15802
rect 30518 15750 30570 15802
rect 30582 15750 30634 15802
rect 30646 15750 30698 15802
rect 30710 15750 30762 15802
rect 30774 15750 30826 15802
rect 6552 15648 6604 15700
rect 8024 15648 8076 15700
rect 13452 15691 13504 15700
rect 13452 15657 13461 15691
rect 13461 15657 13495 15691
rect 13495 15657 13504 15691
rect 13452 15648 13504 15657
rect 18328 15648 18380 15700
rect 22468 15648 22520 15700
rect 6644 15512 6696 15564
rect 14372 15555 14424 15564
rect 14372 15521 14381 15555
rect 14381 15521 14415 15555
rect 14415 15521 14424 15555
rect 14372 15512 14424 15521
rect 20628 15555 20680 15564
rect 20628 15521 20637 15555
rect 20637 15521 20671 15555
rect 20671 15521 20680 15555
rect 20628 15512 20680 15521
rect 6828 15444 6880 15496
rect 20352 15487 20404 15496
rect 20352 15453 20361 15487
rect 20361 15453 20395 15487
rect 20395 15453 20404 15487
rect 20352 15444 20404 15453
rect 6920 15419 6972 15428
rect 6920 15385 6929 15419
rect 6929 15385 6963 15419
rect 6963 15385 6972 15419
rect 6920 15376 6972 15385
rect 15384 15376 15436 15428
rect 19340 15376 19392 15428
rect 6736 15308 6788 15360
rect 9398 15206 9450 15258
rect 9462 15206 9514 15258
rect 9526 15206 9578 15258
rect 9590 15206 9642 15258
rect 9654 15206 9706 15258
rect 17846 15206 17898 15258
rect 17910 15206 17962 15258
rect 17974 15206 18026 15258
rect 18038 15206 18090 15258
rect 18102 15206 18154 15258
rect 26294 15206 26346 15258
rect 26358 15206 26410 15258
rect 26422 15206 26474 15258
rect 26486 15206 26538 15258
rect 26550 15206 26602 15258
rect 15384 15104 15436 15156
rect 17776 15104 17828 15156
rect 21916 15104 21968 15156
rect 29920 15147 29972 15156
rect 29920 15113 29929 15147
rect 29929 15113 29963 15147
rect 29963 15113 29972 15147
rect 29920 15104 29972 15113
rect 24860 15036 24912 15088
rect 14280 15011 14332 15020
rect 14280 14977 14289 15011
rect 14289 14977 14323 15011
rect 14323 14977 14332 15011
rect 14280 14968 14332 14977
rect 21180 14943 21232 14952
rect 21180 14909 21189 14943
rect 21189 14909 21223 14943
rect 21223 14909 21232 14943
rect 21180 14900 21232 14909
rect 19340 14832 19392 14884
rect 6644 14764 6696 14816
rect 28080 14900 28132 14952
rect 29092 14900 29144 14952
rect 29644 14764 29696 14816
rect 5174 14662 5226 14714
rect 5238 14662 5290 14714
rect 5302 14662 5354 14714
rect 5366 14662 5418 14714
rect 5430 14662 5482 14714
rect 13622 14662 13674 14714
rect 13686 14662 13738 14714
rect 13750 14662 13802 14714
rect 13814 14662 13866 14714
rect 13878 14662 13930 14714
rect 22070 14662 22122 14714
rect 22134 14662 22186 14714
rect 22198 14662 22250 14714
rect 22262 14662 22314 14714
rect 22326 14662 22378 14714
rect 30518 14662 30570 14714
rect 30582 14662 30634 14714
rect 30646 14662 30698 14714
rect 30710 14662 30762 14714
rect 30774 14662 30826 14714
rect 6644 14467 6696 14476
rect 6644 14433 6653 14467
rect 6653 14433 6687 14467
rect 6687 14433 6696 14467
rect 6644 14424 6696 14433
rect 5908 14356 5960 14408
rect 6736 14356 6788 14408
rect 5172 14220 5224 14272
rect 12440 14220 12492 14272
rect 9398 14118 9450 14170
rect 9462 14118 9514 14170
rect 9526 14118 9578 14170
rect 9590 14118 9642 14170
rect 9654 14118 9706 14170
rect 17846 14118 17898 14170
rect 17910 14118 17962 14170
rect 17974 14118 18026 14170
rect 18038 14118 18090 14170
rect 18102 14118 18154 14170
rect 26294 14118 26346 14170
rect 26358 14118 26410 14170
rect 26422 14118 26474 14170
rect 26486 14118 26538 14170
rect 26550 14118 26602 14170
rect 31392 14016 31444 14068
rect 29000 13948 29052 14000
rect 5172 13923 5224 13932
rect 5172 13889 5181 13923
rect 5181 13889 5215 13923
rect 5215 13889 5224 13923
rect 5172 13880 5224 13889
rect 28080 13923 28132 13932
rect 28080 13889 28089 13923
rect 28089 13889 28123 13923
rect 28123 13889 28132 13923
rect 28080 13880 28132 13889
rect 31484 13880 31536 13932
rect 6736 13812 6788 13864
rect 28356 13855 28408 13864
rect 28356 13821 28365 13855
rect 28365 13821 28399 13855
rect 28399 13821 28408 13855
rect 28356 13812 28408 13821
rect 4436 13676 4488 13728
rect 34060 13719 34112 13728
rect 34060 13685 34069 13719
rect 34069 13685 34103 13719
rect 34103 13685 34112 13719
rect 34060 13676 34112 13685
rect 5174 13574 5226 13626
rect 5238 13574 5290 13626
rect 5302 13574 5354 13626
rect 5366 13574 5418 13626
rect 5430 13574 5482 13626
rect 13622 13574 13674 13626
rect 13686 13574 13738 13626
rect 13750 13574 13802 13626
rect 13814 13574 13866 13626
rect 13878 13574 13930 13626
rect 22070 13574 22122 13626
rect 22134 13574 22186 13626
rect 22198 13574 22250 13626
rect 22262 13574 22314 13626
rect 22326 13574 22378 13626
rect 30518 13574 30570 13626
rect 30582 13574 30634 13626
rect 30646 13574 30698 13626
rect 30710 13574 30762 13626
rect 30774 13574 30826 13626
rect 5908 13515 5960 13524
rect 5908 13481 5917 13515
rect 5917 13481 5951 13515
rect 5951 13481 5960 13515
rect 5908 13472 5960 13481
rect 6460 13515 6512 13524
rect 6460 13481 6469 13515
rect 6469 13481 6503 13515
rect 6503 13481 6512 13515
rect 6460 13472 6512 13481
rect 20076 13472 20128 13524
rect 24860 13472 24912 13524
rect 28356 13472 28408 13524
rect 30380 13404 30432 13456
rect 31484 13379 31536 13388
rect 31484 13345 31493 13379
rect 31493 13345 31527 13379
rect 31527 13345 31536 13379
rect 31484 13336 31536 13345
rect 14280 13311 14332 13320
rect 14280 13277 14289 13311
rect 14289 13277 14323 13311
rect 14323 13277 14332 13311
rect 14280 13268 14332 13277
rect 19248 13268 19300 13320
rect 31392 13311 31444 13320
rect 4436 13243 4488 13252
rect 4436 13209 4445 13243
rect 4445 13209 4479 13243
rect 4479 13209 4488 13243
rect 4436 13200 4488 13209
rect 6368 13200 6420 13252
rect 14188 13175 14240 13184
rect 14188 13141 14197 13175
rect 14197 13141 14231 13175
rect 14231 13141 14240 13175
rect 14188 13132 14240 13141
rect 20720 13175 20772 13184
rect 20720 13141 20729 13175
rect 20729 13141 20763 13175
rect 20763 13141 20772 13175
rect 20720 13132 20772 13141
rect 30380 13132 30432 13184
rect 31392 13277 31401 13311
rect 31401 13277 31435 13311
rect 31435 13277 31444 13311
rect 31392 13268 31444 13277
rect 9398 13030 9450 13082
rect 9462 13030 9514 13082
rect 9526 13030 9578 13082
rect 9590 13030 9642 13082
rect 9654 13030 9706 13082
rect 17846 13030 17898 13082
rect 17910 13030 17962 13082
rect 17974 13030 18026 13082
rect 18038 13030 18090 13082
rect 18102 13030 18154 13082
rect 26294 13030 26346 13082
rect 26358 13030 26410 13082
rect 26422 13030 26474 13082
rect 26486 13030 26538 13082
rect 26550 13030 26602 13082
rect 6368 12928 6420 12980
rect 12900 12971 12952 12980
rect 12900 12937 12909 12971
rect 12909 12937 12943 12971
rect 12943 12937 12952 12971
rect 12900 12928 12952 12937
rect 13452 12928 13504 12980
rect 14188 12860 14240 12912
rect 6828 12792 6880 12844
rect 15292 12928 15344 12980
rect 20260 12928 20312 12980
rect 21180 12928 21232 12980
rect 29000 12928 29052 12980
rect 20812 12792 20864 12844
rect 27896 12792 27948 12844
rect 1400 12767 1452 12776
rect 1400 12733 1409 12767
rect 1409 12733 1443 12767
rect 1443 12733 1452 12767
rect 1400 12724 1452 12733
rect 6368 12724 6420 12776
rect 14280 12724 14332 12776
rect 20076 12724 20128 12776
rect 21088 12767 21140 12776
rect 21088 12733 21097 12767
rect 21097 12733 21131 12767
rect 21131 12733 21140 12767
rect 21088 12724 21140 12733
rect 12440 12588 12492 12640
rect 15292 12588 15344 12640
rect 20720 12588 20772 12640
rect 22836 12588 22888 12640
rect 5174 12486 5226 12538
rect 5238 12486 5290 12538
rect 5302 12486 5354 12538
rect 5366 12486 5418 12538
rect 5430 12486 5482 12538
rect 13622 12486 13674 12538
rect 13686 12486 13738 12538
rect 13750 12486 13802 12538
rect 13814 12486 13866 12538
rect 13878 12486 13930 12538
rect 22070 12486 22122 12538
rect 22134 12486 22186 12538
rect 22198 12486 22250 12538
rect 22262 12486 22314 12538
rect 22326 12486 22378 12538
rect 30518 12486 30570 12538
rect 30582 12486 30634 12538
rect 30646 12486 30698 12538
rect 30710 12486 30762 12538
rect 30774 12486 30826 12538
rect 1400 12427 1452 12436
rect 1400 12393 1409 12427
rect 1409 12393 1443 12427
rect 1443 12393 1452 12427
rect 1400 12384 1452 12393
rect 6828 12384 6880 12436
rect 20812 12384 20864 12436
rect 21272 12291 21324 12300
rect 21272 12257 21281 12291
rect 21281 12257 21315 12291
rect 21315 12257 21324 12291
rect 21272 12248 21324 12257
rect 27896 12180 27948 12232
rect 21640 12112 21692 12164
rect 6000 12087 6052 12096
rect 6000 12053 6009 12087
rect 6009 12053 6043 12087
rect 6043 12053 6052 12087
rect 6000 12044 6052 12053
rect 20260 12087 20312 12096
rect 20260 12053 20269 12087
rect 20269 12053 20303 12087
rect 20303 12053 20312 12087
rect 20260 12044 20312 12053
rect 33324 12044 33376 12096
rect 9398 11942 9450 11994
rect 9462 11942 9514 11994
rect 9526 11942 9578 11994
rect 9590 11942 9642 11994
rect 9654 11942 9706 11994
rect 17846 11942 17898 11994
rect 17910 11942 17962 11994
rect 17974 11942 18026 11994
rect 18038 11942 18090 11994
rect 18102 11942 18154 11994
rect 26294 11942 26346 11994
rect 26358 11942 26410 11994
rect 26422 11942 26474 11994
rect 26486 11942 26538 11994
rect 26550 11942 26602 11994
rect 6368 11747 6420 11756
rect 6368 11713 6377 11747
rect 6377 11713 6411 11747
rect 6411 11713 6420 11747
rect 6368 11704 6420 11713
rect 20720 11704 20772 11756
rect 31484 11704 31536 11756
rect 6736 11568 6788 11620
rect 21272 11568 21324 11620
rect 5724 11543 5776 11552
rect 5724 11509 5733 11543
rect 5733 11509 5767 11543
rect 5767 11509 5776 11543
rect 5724 11500 5776 11509
rect 21088 11500 21140 11552
rect 34060 11543 34112 11552
rect 34060 11509 34069 11543
rect 34069 11509 34103 11543
rect 34103 11509 34112 11543
rect 34060 11500 34112 11509
rect 5174 11398 5226 11450
rect 5238 11398 5290 11450
rect 5302 11398 5354 11450
rect 5366 11398 5418 11450
rect 5430 11398 5482 11450
rect 13622 11398 13674 11450
rect 13686 11398 13738 11450
rect 13750 11398 13802 11450
rect 13814 11398 13866 11450
rect 13878 11398 13930 11450
rect 22070 11398 22122 11450
rect 22134 11398 22186 11450
rect 22198 11398 22250 11450
rect 22262 11398 22314 11450
rect 22326 11398 22378 11450
rect 30518 11398 30570 11450
rect 30582 11398 30634 11450
rect 30646 11398 30698 11450
rect 30710 11398 30762 11450
rect 30774 11398 30826 11450
rect 6368 11296 6420 11348
rect 11244 11339 11296 11348
rect 11244 11305 11253 11339
rect 11253 11305 11287 11339
rect 11287 11305 11296 11339
rect 11244 11296 11296 11305
rect 12900 11296 12952 11348
rect 12624 11160 12676 11212
rect 21272 11296 21324 11348
rect 27896 11339 27948 11348
rect 27896 11305 27905 11339
rect 27905 11305 27939 11339
rect 27939 11305 27948 11339
rect 27896 11296 27948 11305
rect 20720 11228 20772 11280
rect 12716 11024 12768 11076
rect 13268 11067 13320 11076
rect 13268 11033 13277 11067
rect 13277 11033 13311 11067
rect 13311 11033 13320 11067
rect 13268 11024 13320 11033
rect 14372 11024 14424 11076
rect 27896 11092 27948 11144
rect 29000 11024 29052 11076
rect 30380 11024 30432 11076
rect 31392 11067 31444 11076
rect 31392 11033 31401 11067
rect 31401 11033 31435 11067
rect 31435 11033 31444 11067
rect 31392 11024 31444 11033
rect 31484 11067 31536 11076
rect 31484 11033 31493 11067
rect 31493 11033 31527 11067
rect 31527 11033 31536 11067
rect 31484 11024 31536 11033
rect 29736 10999 29788 11008
rect 29736 10965 29745 10999
rect 29745 10965 29779 10999
rect 29779 10965 29788 10999
rect 29736 10956 29788 10965
rect 9398 10854 9450 10906
rect 9462 10854 9514 10906
rect 9526 10854 9578 10906
rect 9590 10854 9642 10906
rect 9654 10854 9706 10906
rect 17846 10854 17898 10906
rect 17910 10854 17962 10906
rect 17974 10854 18026 10906
rect 18038 10854 18090 10906
rect 18102 10854 18154 10906
rect 26294 10854 26346 10906
rect 26358 10854 26410 10906
rect 26422 10854 26474 10906
rect 26486 10854 26538 10906
rect 26550 10854 26602 10906
rect 12716 10795 12768 10804
rect 12716 10761 12725 10795
rect 12725 10761 12759 10795
rect 12759 10761 12768 10795
rect 12716 10752 12768 10761
rect 3884 10616 3936 10668
rect 6000 10616 6052 10668
rect 12808 10659 12860 10668
rect 12808 10625 12817 10659
rect 12817 10625 12851 10659
rect 12851 10625 12860 10659
rect 12808 10616 12860 10625
rect 19248 10752 19300 10804
rect 31392 10752 31444 10804
rect 29000 10684 29052 10736
rect 17684 10616 17736 10668
rect 20352 10616 20404 10668
rect 27804 10616 27856 10668
rect 27988 10659 28040 10668
rect 27988 10625 27997 10659
rect 27997 10625 28031 10659
rect 28031 10625 28040 10659
rect 27988 10616 28040 10625
rect 29736 10548 29788 10600
rect 3884 10455 3936 10464
rect 3884 10421 3893 10455
rect 3893 10421 3927 10455
rect 3927 10421 3936 10455
rect 3884 10412 3936 10421
rect 4804 10412 4856 10464
rect 5174 10310 5226 10362
rect 5238 10310 5290 10362
rect 5302 10310 5354 10362
rect 5366 10310 5418 10362
rect 5430 10310 5482 10362
rect 13622 10310 13674 10362
rect 13686 10310 13738 10362
rect 13750 10310 13802 10362
rect 13814 10310 13866 10362
rect 13878 10310 13930 10362
rect 22070 10310 22122 10362
rect 22134 10310 22186 10362
rect 22198 10310 22250 10362
rect 22262 10310 22314 10362
rect 22326 10310 22378 10362
rect 30518 10310 30570 10362
rect 30582 10310 30634 10362
rect 30646 10310 30698 10362
rect 30710 10310 30762 10362
rect 30774 10310 30826 10362
rect 11244 10208 11296 10260
rect 13268 10208 13320 10260
rect 20076 10208 20128 10260
rect 17684 10115 17736 10124
rect 4804 10004 4856 10056
rect 17684 10081 17693 10115
rect 17693 10081 17727 10115
rect 17727 10081 17736 10115
rect 17684 10072 17736 10081
rect 21272 10115 21324 10124
rect 21272 10081 21281 10115
rect 21281 10081 21315 10115
rect 21315 10081 21324 10115
rect 21272 10072 21324 10081
rect 14280 10004 14332 10056
rect 20996 10047 21048 10056
rect 20996 10013 21005 10047
rect 21005 10013 21039 10047
rect 21039 10013 21048 10047
rect 20996 10004 21048 10013
rect 14372 9936 14424 9988
rect 4988 9911 5040 9920
rect 4988 9877 4997 9911
rect 4997 9877 5031 9911
rect 5031 9877 5040 9911
rect 4988 9868 5040 9877
rect 13636 9868 13688 9920
rect 15384 9911 15436 9920
rect 15384 9877 15393 9911
rect 15393 9877 15427 9911
rect 15427 9877 15436 9911
rect 15384 9868 15436 9877
rect 9398 9766 9450 9818
rect 9462 9766 9514 9818
rect 9526 9766 9578 9818
rect 9590 9766 9642 9818
rect 9654 9766 9706 9818
rect 17846 9766 17898 9818
rect 17910 9766 17962 9818
rect 17974 9766 18026 9818
rect 18038 9766 18090 9818
rect 18102 9766 18154 9818
rect 26294 9766 26346 9818
rect 26358 9766 26410 9818
rect 26422 9766 26474 9818
rect 26486 9766 26538 9818
rect 26550 9766 26602 9818
rect 4896 9664 4948 9716
rect 12808 9664 12860 9716
rect 14372 9664 14424 9716
rect 4988 9596 5040 9648
rect 6460 9639 6512 9648
rect 6460 9605 6469 9639
rect 6469 9605 6503 9639
rect 6503 9605 6512 9639
rect 6460 9596 6512 9605
rect 12256 9528 12308 9580
rect 13636 9571 13688 9580
rect 13636 9537 13645 9571
rect 13645 9537 13679 9571
rect 13679 9537 13688 9571
rect 13636 9528 13688 9537
rect 4252 9503 4304 9512
rect 3608 9324 3660 9376
rect 4252 9469 4261 9503
rect 4261 9469 4295 9503
rect 4295 9469 4304 9503
rect 4252 9460 4304 9469
rect 12716 9460 12768 9512
rect 5540 9392 5592 9444
rect 6460 9392 6512 9444
rect 11796 9324 11848 9376
rect 5174 9222 5226 9274
rect 5238 9222 5290 9274
rect 5302 9222 5354 9274
rect 5366 9222 5418 9274
rect 5430 9222 5482 9274
rect 13622 9222 13674 9274
rect 13686 9222 13738 9274
rect 13750 9222 13802 9274
rect 13814 9222 13866 9274
rect 13878 9222 13930 9274
rect 22070 9222 22122 9274
rect 22134 9222 22186 9274
rect 22198 9222 22250 9274
rect 22262 9222 22314 9274
rect 22326 9222 22378 9274
rect 30518 9222 30570 9274
rect 30582 9222 30634 9274
rect 30646 9222 30698 9274
rect 30710 9222 30762 9274
rect 30774 9222 30826 9274
rect 4252 9120 4304 9172
rect 10876 9120 10928 9172
rect 27896 9120 27948 9172
rect 12716 9027 12768 9036
rect 12716 8993 12725 9027
rect 12725 8993 12759 9027
rect 12759 8993 12768 9027
rect 12716 8984 12768 8993
rect 21272 8984 21324 9036
rect 21732 9027 21784 9036
rect 21732 8993 21741 9027
rect 21741 8993 21775 9027
rect 21775 8993 21784 9027
rect 21732 8984 21784 8993
rect 11796 8916 11848 8968
rect 12624 8959 12676 8968
rect 12624 8925 12633 8959
rect 12633 8925 12667 8959
rect 12667 8925 12676 8959
rect 12624 8916 12676 8925
rect 21916 8916 21968 8968
rect 22836 8959 22888 8968
rect 22836 8925 22845 8959
rect 22845 8925 22879 8959
rect 22879 8925 22888 8959
rect 22836 8916 22888 8925
rect 26700 8916 26752 8968
rect 33876 8959 33928 8968
rect 33876 8925 33885 8959
rect 33885 8925 33919 8959
rect 33919 8925 33928 8959
rect 33876 8916 33928 8925
rect 28724 8823 28776 8832
rect 28724 8789 28733 8823
rect 28733 8789 28767 8823
rect 28767 8789 28776 8823
rect 28724 8780 28776 8789
rect 34060 8823 34112 8832
rect 34060 8789 34069 8823
rect 34069 8789 34103 8823
rect 34103 8789 34112 8823
rect 34060 8780 34112 8789
rect 9398 8678 9450 8730
rect 9462 8678 9514 8730
rect 9526 8678 9578 8730
rect 9590 8678 9642 8730
rect 9654 8678 9706 8730
rect 17846 8678 17898 8730
rect 17910 8678 17962 8730
rect 17974 8678 18026 8730
rect 18038 8678 18090 8730
rect 18102 8678 18154 8730
rect 26294 8678 26346 8730
rect 26358 8678 26410 8730
rect 26422 8678 26474 8730
rect 26486 8678 26538 8730
rect 26550 8678 26602 8730
rect 14280 8619 14332 8628
rect 14280 8585 14289 8619
rect 14289 8585 14323 8619
rect 14323 8585 14332 8619
rect 14280 8576 14332 8585
rect 28724 8508 28776 8560
rect 11796 8483 11848 8492
rect 11796 8449 11805 8483
rect 11805 8449 11839 8483
rect 11839 8449 11848 8483
rect 11796 8440 11848 8449
rect 12624 8440 12676 8492
rect 13544 8440 13596 8492
rect 27804 8483 27856 8492
rect 11980 8372 12032 8424
rect 27804 8449 27813 8483
rect 27813 8449 27847 8483
rect 27847 8449 27856 8483
rect 27804 8440 27856 8449
rect 28080 8415 28132 8424
rect 28080 8381 28089 8415
rect 28089 8381 28123 8415
rect 28123 8381 28132 8415
rect 28080 8372 28132 8381
rect 27344 8236 27396 8288
rect 31484 8304 31536 8356
rect 5174 8134 5226 8186
rect 5238 8134 5290 8186
rect 5302 8134 5354 8186
rect 5366 8134 5418 8186
rect 5430 8134 5482 8186
rect 13622 8134 13674 8186
rect 13686 8134 13738 8186
rect 13750 8134 13802 8186
rect 13814 8134 13866 8186
rect 13878 8134 13930 8186
rect 22070 8134 22122 8186
rect 22134 8134 22186 8186
rect 22198 8134 22250 8186
rect 22262 8134 22314 8186
rect 22326 8134 22378 8186
rect 30518 8134 30570 8186
rect 30582 8134 30634 8186
rect 30646 8134 30698 8186
rect 30710 8134 30762 8186
rect 30774 8134 30826 8186
rect 5724 8032 5776 8084
rect 10876 8075 10928 8084
rect 10876 8041 10885 8075
rect 10885 8041 10919 8075
rect 10919 8041 10928 8075
rect 10876 8032 10928 8041
rect 12624 8032 12676 8084
rect 28080 8032 28132 8084
rect 33876 8032 33928 8084
rect 26700 7964 26752 8016
rect 30380 7964 30432 8016
rect 1400 7871 1452 7880
rect 1400 7837 1409 7871
rect 1409 7837 1443 7871
rect 1443 7837 1452 7871
rect 1400 7828 1452 7837
rect 10968 7871 11020 7880
rect 10968 7837 10977 7871
rect 10977 7837 11011 7871
rect 11011 7837 11020 7871
rect 10968 7828 11020 7837
rect 11796 7896 11848 7948
rect 20260 7896 20312 7948
rect 21916 7896 21968 7948
rect 11704 7871 11756 7880
rect 11704 7837 11713 7871
rect 11713 7837 11747 7871
rect 11747 7837 11756 7871
rect 11704 7828 11756 7837
rect 19340 7828 19392 7880
rect 19800 7871 19852 7880
rect 19800 7837 19809 7871
rect 19809 7837 19843 7871
rect 19843 7837 19852 7871
rect 19800 7828 19852 7837
rect 20812 7828 20864 7880
rect 27712 7828 27764 7880
rect 31668 7871 31720 7880
rect 11796 7760 11848 7812
rect 20996 7760 21048 7812
rect 31668 7837 31677 7871
rect 31677 7837 31711 7871
rect 31711 7837 31720 7871
rect 31668 7828 31720 7837
rect 32128 7760 32180 7812
rect 12348 7692 12400 7744
rect 24768 7692 24820 7744
rect 9398 7590 9450 7642
rect 9462 7590 9514 7642
rect 9526 7590 9578 7642
rect 9590 7590 9642 7642
rect 9654 7590 9706 7642
rect 17846 7590 17898 7642
rect 17910 7590 17962 7642
rect 17974 7590 18026 7642
rect 18038 7590 18090 7642
rect 18102 7590 18154 7642
rect 26294 7590 26346 7642
rect 26358 7590 26410 7642
rect 26422 7590 26474 7642
rect 26486 7590 26538 7642
rect 26550 7590 26602 7642
rect 1400 7531 1452 7540
rect 1400 7497 1409 7531
rect 1409 7497 1443 7531
rect 1443 7497 1452 7531
rect 1400 7488 1452 7497
rect 10968 7488 11020 7540
rect 26700 7488 26752 7540
rect 27344 7531 27396 7540
rect 27344 7497 27353 7531
rect 27353 7497 27387 7531
rect 27387 7497 27396 7531
rect 27344 7488 27396 7497
rect 27712 7531 27764 7540
rect 27712 7497 27721 7531
rect 27721 7497 27755 7531
rect 27755 7497 27764 7531
rect 27712 7488 27764 7497
rect 4896 7420 4948 7472
rect 3608 7395 3660 7404
rect 3608 7361 3617 7395
rect 3617 7361 3651 7395
rect 3651 7361 3660 7395
rect 3608 7352 3660 7361
rect 12348 7395 12400 7404
rect 12348 7361 12357 7395
rect 12357 7361 12391 7395
rect 12391 7361 12400 7395
rect 12348 7352 12400 7361
rect 12532 7352 12584 7404
rect 12624 7352 12676 7404
rect 14280 7352 14332 7404
rect 14740 7395 14792 7404
rect 14740 7361 14749 7395
rect 14749 7361 14783 7395
rect 14783 7361 14792 7395
rect 14740 7352 14792 7361
rect 5632 7284 5684 7336
rect 26700 7284 26752 7336
rect 27252 7327 27304 7336
rect 27252 7293 27261 7327
rect 27261 7293 27295 7327
rect 27295 7293 27304 7327
rect 27252 7284 27304 7293
rect 12716 7216 12768 7268
rect 19800 7216 19852 7268
rect 20352 7216 20404 7268
rect 6184 7148 6236 7200
rect 20812 7148 20864 7200
rect 5174 7046 5226 7098
rect 5238 7046 5290 7098
rect 5302 7046 5354 7098
rect 5366 7046 5418 7098
rect 5430 7046 5482 7098
rect 13622 7046 13674 7098
rect 13686 7046 13738 7098
rect 13750 7046 13802 7098
rect 13814 7046 13866 7098
rect 13878 7046 13930 7098
rect 22070 7046 22122 7098
rect 22134 7046 22186 7098
rect 22198 7046 22250 7098
rect 22262 7046 22314 7098
rect 22326 7046 22378 7098
rect 30518 7046 30570 7098
rect 30582 7046 30634 7098
rect 30646 7046 30698 7098
rect 30710 7046 30762 7098
rect 30774 7046 30826 7098
rect 5540 6944 5592 6996
rect 12256 6944 12308 6996
rect 12348 6944 12400 6996
rect 20260 6944 20312 6996
rect 20812 6987 20864 6996
rect 20812 6953 20821 6987
rect 20821 6953 20855 6987
rect 20855 6953 20864 6987
rect 20812 6944 20864 6953
rect 5632 6876 5684 6928
rect 4896 6808 4948 6860
rect 5540 6808 5592 6860
rect 12348 6808 12400 6860
rect 4804 6740 4856 6792
rect 11796 6783 11848 6792
rect 11796 6749 11805 6783
rect 11805 6749 11839 6783
rect 11839 6749 11848 6783
rect 11796 6740 11848 6749
rect 11980 6740 12032 6792
rect 20168 6783 20220 6792
rect 20168 6749 20177 6783
rect 20177 6749 20211 6783
rect 20211 6749 20220 6783
rect 20168 6740 20220 6749
rect 20260 6740 20312 6792
rect 5540 6647 5592 6656
rect 5540 6613 5549 6647
rect 5549 6613 5583 6647
rect 5583 6613 5592 6647
rect 5540 6604 5592 6613
rect 20352 6604 20404 6656
rect 33140 6740 33192 6792
rect 31668 6672 31720 6724
rect 23204 6604 23256 6656
rect 30564 6647 30616 6656
rect 30564 6613 30573 6647
rect 30573 6613 30607 6647
rect 30607 6613 30616 6647
rect 30564 6604 30616 6613
rect 34060 6647 34112 6656
rect 34060 6613 34069 6647
rect 34069 6613 34103 6647
rect 34103 6613 34112 6647
rect 34060 6604 34112 6613
rect 9398 6502 9450 6554
rect 9462 6502 9514 6554
rect 9526 6502 9578 6554
rect 9590 6502 9642 6554
rect 9654 6502 9706 6554
rect 17846 6502 17898 6554
rect 17910 6502 17962 6554
rect 17974 6502 18026 6554
rect 18038 6502 18090 6554
rect 18102 6502 18154 6554
rect 26294 6502 26346 6554
rect 26358 6502 26410 6554
rect 26422 6502 26474 6554
rect 26486 6502 26538 6554
rect 26550 6502 26602 6554
rect 4804 6400 4856 6452
rect 12256 6443 12308 6452
rect 12256 6409 12265 6443
rect 12265 6409 12299 6443
rect 12299 6409 12308 6443
rect 12256 6400 12308 6409
rect 33140 6443 33192 6452
rect 33140 6409 33149 6443
rect 33149 6409 33183 6443
rect 33183 6409 33192 6443
rect 33140 6400 33192 6409
rect 12532 6264 12584 6316
rect 24768 6264 24820 6316
rect 30564 6264 30616 6316
rect 32128 6239 32180 6248
rect 32128 6205 32137 6239
rect 32137 6205 32171 6239
rect 32171 6205 32180 6239
rect 32128 6196 32180 6205
rect 12440 6128 12492 6180
rect 29828 6060 29880 6112
rect 5174 5958 5226 6010
rect 5238 5958 5290 6010
rect 5302 5958 5354 6010
rect 5366 5958 5418 6010
rect 5430 5958 5482 6010
rect 13622 5958 13674 6010
rect 13686 5958 13738 6010
rect 13750 5958 13802 6010
rect 13814 5958 13866 6010
rect 13878 5958 13930 6010
rect 22070 5958 22122 6010
rect 22134 5958 22186 6010
rect 22198 5958 22250 6010
rect 22262 5958 22314 6010
rect 22326 5958 22378 6010
rect 30518 5958 30570 6010
rect 30582 5958 30634 6010
rect 30646 5958 30698 6010
rect 30710 5958 30762 6010
rect 30774 5958 30826 6010
rect 11704 5763 11756 5772
rect 4804 5652 4856 5704
rect 6184 5695 6236 5704
rect 6184 5661 6193 5695
rect 6193 5661 6227 5695
rect 6227 5661 6236 5695
rect 11704 5729 11713 5763
rect 11713 5729 11747 5763
rect 11747 5729 11756 5763
rect 11704 5720 11756 5729
rect 6184 5652 6236 5661
rect 12440 5652 12492 5704
rect 6276 5584 6328 5636
rect 4528 5516 4580 5568
rect 12164 5516 12216 5568
rect 9398 5414 9450 5466
rect 9462 5414 9514 5466
rect 9526 5414 9578 5466
rect 9590 5414 9642 5466
rect 9654 5414 9706 5466
rect 17846 5414 17898 5466
rect 17910 5414 17962 5466
rect 17974 5414 18026 5466
rect 18038 5414 18090 5466
rect 18102 5414 18154 5466
rect 26294 5414 26346 5466
rect 26358 5414 26410 5466
rect 26422 5414 26474 5466
rect 26486 5414 26538 5466
rect 26550 5414 26602 5466
rect 12348 5355 12400 5364
rect 12348 5321 12357 5355
rect 12357 5321 12391 5355
rect 12391 5321 12400 5355
rect 12348 5312 12400 5321
rect 21732 5244 21784 5296
rect 12440 5219 12492 5228
rect 12440 5185 12449 5219
rect 12449 5185 12483 5219
rect 12483 5185 12492 5219
rect 12440 5176 12492 5185
rect 12808 5176 12860 5228
rect 19616 5219 19668 5228
rect 19616 5185 19625 5219
rect 19625 5185 19659 5219
rect 19659 5185 19668 5219
rect 19616 5176 19668 5185
rect 29552 5244 29604 5296
rect 32128 5244 32180 5296
rect 23204 5219 23256 5228
rect 23204 5185 23213 5219
rect 23213 5185 23247 5219
rect 23247 5185 23256 5219
rect 23204 5176 23256 5185
rect 12532 5108 12584 5160
rect 24584 4972 24636 5024
rect 5174 4870 5226 4922
rect 5238 4870 5290 4922
rect 5302 4870 5354 4922
rect 5366 4870 5418 4922
rect 5430 4870 5482 4922
rect 13622 4870 13674 4922
rect 13686 4870 13738 4922
rect 13750 4870 13802 4922
rect 13814 4870 13866 4922
rect 13878 4870 13930 4922
rect 22070 4870 22122 4922
rect 22134 4870 22186 4922
rect 22198 4870 22250 4922
rect 22262 4870 22314 4922
rect 22326 4870 22378 4922
rect 30518 4870 30570 4922
rect 30582 4870 30634 4922
rect 30646 4870 30698 4922
rect 30710 4870 30762 4922
rect 30774 4870 30826 4922
rect 19616 4811 19668 4820
rect 19616 4777 19625 4811
rect 19625 4777 19659 4811
rect 19659 4777 19668 4811
rect 19616 4768 19668 4777
rect 12532 4700 12584 4752
rect 12440 4632 12492 4684
rect 12624 4632 12676 4684
rect 6368 4539 6420 4548
rect 6368 4505 6377 4539
rect 6377 4505 6411 4539
rect 6411 4505 6420 4539
rect 6368 4496 6420 4505
rect 12808 4564 12860 4616
rect 17132 4564 17184 4616
rect 19340 4632 19392 4684
rect 29552 4675 29604 4684
rect 29552 4641 29561 4675
rect 29561 4641 29595 4675
rect 29595 4641 29604 4675
rect 29552 4632 29604 4641
rect 15660 4496 15712 4548
rect 11520 4428 11572 4480
rect 20168 4564 20220 4616
rect 29828 4607 29880 4616
rect 29828 4573 29837 4607
rect 29837 4573 29871 4607
rect 29871 4573 29880 4607
rect 29828 4564 29880 4573
rect 31576 4428 31628 4480
rect 9398 4326 9450 4378
rect 9462 4326 9514 4378
rect 9526 4326 9578 4378
rect 9590 4326 9642 4378
rect 9654 4326 9706 4378
rect 17846 4326 17898 4378
rect 17910 4326 17962 4378
rect 17974 4326 18026 4378
rect 18038 4326 18090 4378
rect 18102 4326 18154 4378
rect 26294 4326 26346 4378
rect 26358 4326 26410 4378
rect 26422 4326 26474 4378
rect 26486 4326 26538 4378
rect 26550 4326 26602 4378
rect 12808 4224 12860 4276
rect 4528 4156 4580 4208
rect 12624 4156 12676 4208
rect 11520 4131 11572 4140
rect 11520 4097 11529 4131
rect 11529 4097 11563 4131
rect 11563 4097 11572 4131
rect 11520 4088 11572 4097
rect 11980 4088 12032 4140
rect 12164 4131 12216 4140
rect 12164 4097 12173 4131
rect 12173 4097 12207 4131
rect 12207 4097 12216 4131
rect 12164 4088 12216 4097
rect 12440 4131 12492 4140
rect 12440 4097 12449 4131
rect 12449 4097 12483 4131
rect 12483 4097 12492 4131
rect 12440 4088 12492 4097
rect 3792 4063 3844 4072
rect 3792 4029 3801 4063
rect 3801 4029 3835 4063
rect 3835 4029 3844 4063
rect 3792 4020 3844 4029
rect 6368 4020 6420 4072
rect 11796 4020 11848 4072
rect 12808 4131 12860 4140
rect 12808 4097 12817 4131
rect 12817 4097 12851 4131
rect 12851 4097 12860 4131
rect 12808 4088 12860 4097
rect 33876 4131 33928 4140
rect 33876 4097 33885 4131
rect 33885 4097 33919 4131
rect 33919 4097 33928 4131
rect 33876 4088 33928 4097
rect 5540 3952 5592 4004
rect 12716 3952 12768 4004
rect 13820 4020 13872 4072
rect 17132 4020 17184 4072
rect 15660 3995 15712 4004
rect 15660 3961 15669 3995
rect 15669 3961 15703 3995
rect 15703 3961 15712 3995
rect 15660 3952 15712 3961
rect 11704 3927 11756 3936
rect 11704 3893 11713 3927
rect 11713 3893 11747 3927
rect 11747 3893 11756 3927
rect 11704 3884 11756 3893
rect 12164 3884 12216 3936
rect 14740 3884 14792 3936
rect 24584 3884 24636 3936
rect 31668 3884 31720 3936
rect 34060 3927 34112 3936
rect 34060 3893 34069 3927
rect 34069 3893 34103 3927
rect 34103 3893 34112 3927
rect 34060 3884 34112 3893
rect 5174 3782 5226 3834
rect 5238 3782 5290 3834
rect 5302 3782 5354 3834
rect 5366 3782 5418 3834
rect 5430 3782 5482 3834
rect 13622 3782 13674 3834
rect 13686 3782 13738 3834
rect 13750 3782 13802 3834
rect 13814 3782 13866 3834
rect 13878 3782 13930 3834
rect 22070 3782 22122 3834
rect 22134 3782 22186 3834
rect 22198 3782 22250 3834
rect 22262 3782 22314 3834
rect 22326 3782 22378 3834
rect 30518 3782 30570 3834
rect 30582 3782 30634 3834
rect 30646 3782 30698 3834
rect 30710 3782 30762 3834
rect 30774 3782 30826 3834
rect 3792 3680 3844 3732
rect 21640 3680 21692 3732
rect 24584 3723 24636 3732
rect 24584 3689 24593 3723
rect 24593 3689 24627 3723
rect 24627 3689 24636 3723
rect 24584 3680 24636 3689
rect 11980 3612 12032 3664
rect 15660 3612 15712 3664
rect 23664 3655 23716 3664
rect 23664 3621 23673 3655
rect 23673 3621 23707 3655
rect 23707 3621 23716 3655
rect 27252 3680 27304 3732
rect 29644 3723 29696 3732
rect 29644 3689 29653 3723
rect 29653 3689 29687 3723
rect 29687 3689 29696 3723
rect 29644 3680 29696 3689
rect 31576 3723 31628 3732
rect 23664 3612 23716 3621
rect 5080 3587 5132 3596
rect 5080 3553 5089 3587
rect 5089 3553 5123 3587
rect 5123 3553 5132 3587
rect 5080 3544 5132 3553
rect 12164 3544 12216 3596
rect 12808 3544 12860 3596
rect 6828 3476 6880 3528
rect 11704 3476 11756 3528
rect 12716 3519 12768 3528
rect 12716 3485 12725 3519
rect 12725 3485 12759 3519
rect 12759 3485 12768 3519
rect 12716 3476 12768 3485
rect 12532 3451 12584 3460
rect 12532 3417 12541 3451
rect 12541 3417 12575 3451
rect 12575 3417 12584 3451
rect 12532 3408 12584 3417
rect 12348 3340 12400 3392
rect 23756 3476 23808 3528
rect 31576 3689 31585 3723
rect 31585 3689 31619 3723
rect 31619 3689 31628 3723
rect 31576 3680 31628 3689
rect 22560 3451 22612 3460
rect 22560 3417 22569 3451
rect 22569 3417 22603 3451
rect 22603 3417 22612 3451
rect 22560 3408 22612 3417
rect 23388 3408 23440 3460
rect 24400 3451 24452 3460
rect 24400 3417 24409 3451
rect 24409 3417 24443 3451
rect 24443 3417 24452 3451
rect 24400 3408 24452 3417
rect 30748 3476 30800 3528
rect 31668 3519 31720 3528
rect 31668 3485 31677 3519
rect 31677 3485 31711 3519
rect 31711 3485 31720 3519
rect 31668 3476 31720 3485
rect 33876 3476 33928 3528
rect 30932 3340 30984 3392
rect 9398 3238 9450 3290
rect 9462 3238 9514 3290
rect 9526 3238 9578 3290
rect 9590 3238 9642 3290
rect 9654 3238 9706 3290
rect 17846 3238 17898 3290
rect 17910 3238 17962 3290
rect 17974 3238 18026 3290
rect 18038 3238 18090 3290
rect 18102 3238 18154 3290
rect 26294 3238 26346 3290
rect 26358 3238 26410 3290
rect 26422 3238 26474 3290
rect 26486 3238 26538 3290
rect 26550 3238 26602 3290
rect 12532 3179 12584 3188
rect 12532 3145 12541 3179
rect 12541 3145 12575 3179
rect 12575 3145 12584 3179
rect 12532 3136 12584 3145
rect 23756 3179 23808 3188
rect 23756 3145 23765 3179
rect 23765 3145 23799 3179
rect 23799 3145 23808 3179
rect 23756 3136 23808 3145
rect 30748 3179 30800 3188
rect 30748 3145 30757 3179
rect 30757 3145 30791 3179
rect 30791 3145 30800 3179
rect 30748 3136 30800 3145
rect 24400 3068 24452 3120
rect 12164 3043 12216 3052
rect 12164 3009 12173 3043
rect 12173 3009 12207 3043
rect 12207 3009 12216 3043
rect 12164 3000 12216 3009
rect 12624 3000 12676 3052
rect 24584 3000 24636 3052
rect 30932 3043 30984 3052
rect 30932 3009 30941 3043
rect 30941 3009 30975 3043
rect 30975 3009 30984 3043
rect 30932 3000 30984 3009
rect 1768 2839 1820 2848
rect 1768 2805 1777 2839
rect 1777 2805 1811 2839
rect 1811 2805 1820 2839
rect 1768 2796 1820 2805
rect 13544 2796 13596 2848
rect 23388 2796 23440 2848
rect 5174 2694 5226 2746
rect 5238 2694 5290 2746
rect 5302 2694 5354 2746
rect 5366 2694 5418 2746
rect 5430 2694 5482 2746
rect 13622 2694 13674 2746
rect 13686 2694 13738 2746
rect 13750 2694 13802 2746
rect 13814 2694 13866 2746
rect 13878 2694 13930 2746
rect 22070 2694 22122 2746
rect 22134 2694 22186 2746
rect 22198 2694 22250 2746
rect 22262 2694 22314 2746
rect 22326 2694 22378 2746
rect 30518 2694 30570 2746
rect 30582 2694 30634 2746
rect 30646 2694 30698 2746
rect 30710 2694 30762 2746
rect 30774 2694 30826 2746
rect 3148 2592 3200 2644
rect 15384 2592 15436 2644
rect 3884 2524 3936 2576
rect 5080 2524 5132 2576
rect 6828 2567 6880 2576
rect 6828 2533 6837 2567
rect 6837 2533 6871 2567
rect 6871 2533 6880 2567
rect 6828 2524 6880 2533
rect 1768 2388 1820 2440
rect 4252 2388 4304 2440
rect 6920 2388 6972 2440
rect 9220 2388 9272 2440
rect 23664 2456 23716 2508
rect 33968 2456 34020 2508
rect 21640 2388 21692 2440
rect 29644 2388 29696 2440
rect 31576 2388 31628 2440
rect 22560 2320 22612 2372
rect 14188 2252 14240 2304
rect 21640 2252 21692 2304
rect 29092 2252 29144 2304
rect 34060 2295 34112 2304
rect 34060 2261 34069 2295
rect 34069 2261 34103 2295
rect 34103 2261 34112 2295
rect 34060 2252 34112 2261
rect 9398 2150 9450 2202
rect 9462 2150 9514 2202
rect 9526 2150 9578 2202
rect 9590 2150 9642 2202
rect 9654 2150 9706 2202
rect 17846 2150 17898 2202
rect 17910 2150 17962 2202
rect 17974 2150 18026 2202
rect 18038 2150 18090 2202
rect 18102 2150 18154 2202
rect 26294 2150 26346 2202
rect 26358 2150 26410 2202
rect 26422 2150 26474 2202
rect 26486 2150 26538 2202
rect 26550 2150 26602 2202
<< metal2 >>
rect 3606 19200 3662 20000
rect 10782 19200 10838 20000
rect 17958 19200 18014 20000
rect 18064 19230 18276 19258
rect 1398 17368 1454 17377
rect 3620 17338 3648 19200
rect 9398 17436 9706 17445
rect 9398 17434 9404 17436
rect 9460 17434 9484 17436
rect 9540 17434 9564 17436
rect 9620 17434 9644 17436
rect 9700 17434 9706 17436
rect 9460 17382 9462 17434
rect 9642 17382 9644 17434
rect 9398 17380 9404 17382
rect 9460 17380 9484 17382
rect 9540 17380 9564 17382
rect 9620 17380 9644 17382
rect 9700 17380 9706 17382
rect 9398 17371 9706 17380
rect 10796 17338 10824 19200
rect 17972 19122 18000 19200
rect 18064 19122 18092 19230
rect 17972 19094 18092 19122
rect 17846 17436 18154 17445
rect 17846 17434 17852 17436
rect 17908 17434 17932 17436
rect 17988 17434 18012 17436
rect 18068 17434 18092 17436
rect 18148 17434 18154 17436
rect 17908 17382 17910 17434
rect 18090 17382 18092 17434
rect 17846 17380 17852 17382
rect 17908 17380 17932 17382
rect 17988 17380 18012 17382
rect 18068 17380 18092 17382
rect 18148 17380 18154 17382
rect 17846 17371 18154 17380
rect 18248 17338 18276 19230
rect 25134 19200 25190 20000
rect 32310 19200 32366 20000
rect 25148 17338 25176 19200
rect 26294 17436 26602 17445
rect 26294 17434 26300 17436
rect 26356 17434 26380 17436
rect 26436 17434 26460 17436
rect 26516 17434 26540 17436
rect 26596 17434 26602 17436
rect 26356 17382 26358 17434
rect 26538 17382 26540 17434
rect 26294 17380 26300 17382
rect 26356 17380 26380 17382
rect 26436 17380 26460 17382
rect 26516 17380 26540 17382
rect 26596 17380 26602 17382
rect 26294 17371 26602 17380
rect 32324 17338 32352 19200
rect 34058 18592 34114 18601
rect 34058 18527 34114 18536
rect 34072 17338 34100 18527
rect 1398 17303 1454 17312
rect 3608 17332 3660 17338
rect 1412 17202 1440 17303
rect 3608 17274 3660 17280
rect 10784 17332 10836 17338
rect 10784 17274 10836 17280
rect 18236 17332 18288 17338
rect 18236 17274 18288 17280
rect 25136 17332 25188 17338
rect 25136 17274 25188 17280
rect 32312 17332 32364 17338
rect 32312 17274 32364 17280
rect 34060 17332 34112 17338
rect 34060 17274 34112 17280
rect 1400 17196 1452 17202
rect 1400 17138 1452 17144
rect 6828 17196 6880 17202
rect 6828 17138 6880 17144
rect 11520 17196 11572 17202
rect 11520 17138 11572 17144
rect 18328 17196 18380 17202
rect 18328 17138 18380 17144
rect 25504 17196 25556 17202
rect 25504 17138 25556 17144
rect 29920 17196 29972 17202
rect 29920 17138 29972 17144
rect 33324 17196 33376 17202
rect 33324 17138 33376 17144
rect 1412 16794 1440 17138
rect 5174 16892 5482 16901
rect 5174 16890 5180 16892
rect 5236 16890 5260 16892
rect 5316 16890 5340 16892
rect 5396 16890 5420 16892
rect 5476 16890 5482 16892
rect 5236 16838 5238 16890
rect 5418 16838 5420 16890
rect 5174 16836 5180 16838
rect 5236 16836 5260 16838
rect 5316 16836 5340 16838
rect 5396 16836 5420 16838
rect 5476 16836 5482 16838
rect 5174 16827 5482 16836
rect 1400 16788 1452 16794
rect 1400 16730 1452 16736
rect 6552 16584 6604 16590
rect 6840 16574 6868 17138
rect 6552 16526 6604 16532
rect 6748 16546 6868 16574
rect 6460 16040 6512 16046
rect 6460 15982 6512 15988
rect 5174 15804 5482 15813
rect 5174 15802 5180 15804
rect 5236 15802 5260 15804
rect 5316 15802 5340 15804
rect 5396 15802 5420 15804
rect 5476 15802 5482 15804
rect 5236 15750 5238 15802
rect 5418 15750 5420 15802
rect 5174 15748 5180 15750
rect 5236 15748 5260 15750
rect 5316 15748 5340 15750
rect 5396 15748 5420 15750
rect 5476 15748 5482 15750
rect 5174 15739 5482 15748
rect 5174 14716 5482 14725
rect 5174 14714 5180 14716
rect 5236 14714 5260 14716
rect 5316 14714 5340 14716
rect 5396 14714 5420 14716
rect 5476 14714 5482 14716
rect 5236 14662 5238 14714
rect 5418 14662 5420 14714
rect 5174 14660 5180 14662
rect 5236 14660 5260 14662
rect 5316 14660 5340 14662
rect 5396 14660 5420 14662
rect 5476 14660 5482 14662
rect 5174 14651 5482 14660
rect 5908 14408 5960 14414
rect 5908 14350 5960 14356
rect 5172 14272 5224 14278
rect 5172 14214 5224 14220
rect 5184 13938 5212 14214
rect 5172 13932 5224 13938
rect 5172 13874 5224 13880
rect 4436 13728 4488 13734
rect 4436 13670 4488 13676
rect 4448 13258 4476 13670
rect 5174 13628 5482 13637
rect 5174 13626 5180 13628
rect 5236 13626 5260 13628
rect 5316 13626 5340 13628
rect 5396 13626 5420 13628
rect 5476 13626 5482 13628
rect 5236 13574 5238 13626
rect 5418 13574 5420 13626
rect 5174 13572 5180 13574
rect 5236 13572 5260 13574
rect 5316 13572 5340 13574
rect 5396 13572 5420 13574
rect 5476 13572 5482 13574
rect 5174 13563 5482 13572
rect 5920 13530 5948 14350
rect 6472 13530 6500 15982
rect 6564 15706 6592 16526
rect 6552 15700 6604 15706
rect 6552 15642 6604 15648
rect 6644 15564 6696 15570
rect 6644 15506 6696 15512
rect 6656 14822 6684 15506
rect 6748 15366 6776 16546
rect 7012 16448 7064 16454
rect 7012 16390 7064 16396
rect 6920 16244 6972 16250
rect 6920 16186 6972 16192
rect 6828 15496 6880 15502
rect 6828 15438 6880 15444
rect 6736 15360 6788 15366
rect 6736 15302 6788 15308
rect 6644 14816 6696 14822
rect 6644 14758 6696 14764
rect 6656 14482 6684 14758
rect 6644 14476 6696 14482
rect 6644 14418 6696 14424
rect 6656 13954 6684 14418
rect 6748 14414 6776 15302
rect 6736 14408 6788 14414
rect 6736 14350 6788 14356
rect 6656 13926 6776 13954
rect 6748 13870 6776 13926
rect 6736 13864 6788 13870
rect 6736 13806 6788 13812
rect 5908 13524 5960 13530
rect 5908 13466 5960 13472
rect 6460 13524 6512 13530
rect 6460 13466 6512 13472
rect 4436 13252 4488 13258
rect 4436 13194 4488 13200
rect 6368 13252 6420 13258
rect 6368 13194 6420 13200
rect 6380 12986 6408 13194
rect 6368 12980 6420 12986
rect 6368 12922 6420 12928
rect 1400 12776 1452 12782
rect 1400 12718 1452 12724
rect 6368 12776 6420 12782
rect 6368 12718 6420 12724
rect 1412 12481 1440 12718
rect 5174 12540 5482 12549
rect 5174 12538 5180 12540
rect 5236 12538 5260 12540
rect 5316 12538 5340 12540
rect 5396 12538 5420 12540
rect 5476 12538 5482 12540
rect 5236 12486 5238 12538
rect 5418 12486 5420 12538
rect 5174 12484 5180 12486
rect 5236 12484 5260 12486
rect 5316 12484 5340 12486
rect 5396 12484 5420 12486
rect 5476 12484 5482 12486
rect 1398 12472 1454 12481
rect 5174 12475 5482 12484
rect 1398 12407 1400 12416
rect 1452 12407 1454 12416
rect 1400 12378 1452 12384
rect 6000 12096 6052 12102
rect 6000 12038 6052 12044
rect 5724 11552 5776 11558
rect 5724 11494 5776 11500
rect 5174 11452 5482 11461
rect 5174 11450 5180 11452
rect 5236 11450 5260 11452
rect 5316 11450 5340 11452
rect 5396 11450 5420 11452
rect 5476 11450 5482 11452
rect 5236 11398 5238 11450
rect 5418 11398 5420 11450
rect 5174 11396 5180 11398
rect 5236 11396 5260 11398
rect 5316 11396 5340 11398
rect 5396 11396 5420 11398
rect 5476 11396 5482 11398
rect 5174 11387 5482 11396
rect 3884 10668 3936 10674
rect 3884 10610 3936 10616
rect 3896 10470 3924 10610
rect 3884 10464 3936 10470
rect 3884 10406 3936 10412
rect 4804 10464 4856 10470
rect 4804 10406 4856 10412
rect 3608 9376 3660 9382
rect 3608 9318 3660 9324
rect 1400 7880 1452 7886
rect 1400 7822 1452 7828
rect 1412 7585 1440 7822
rect 1398 7576 1454 7585
rect 1398 7511 1400 7520
rect 1452 7511 1454 7520
rect 1400 7482 1452 7488
rect 3620 7410 3648 9318
rect 3608 7404 3660 7410
rect 3608 7346 3660 7352
rect 3792 4072 3844 4078
rect 3792 4014 3844 4020
rect 3804 3738 3832 4014
rect 3792 3732 3844 3738
rect 3792 3674 3844 3680
rect 1768 2848 1820 2854
rect 1768 2790 1820 2796
rect 1780 2446 1808 2790
rect 3146 2680 3202 2689
rect 3146 2615 3148 2624
rect 3200 2615 3202 2624
rect 3148 2586 3200 2592
rect 3896 2582 3924 10406
rect 4816 10062 4844 10406
rect 5174 10364 5482 10373
rect 5174 10362 5180 10364
rect 5236 10362 5260 10364
rect 5316 10362 5340 10364
rect 5396 10362 5420 10364
rect 5476 10362 5482 10364
rect 5236 10310 5238 10362
rect 5418 10310 5420 10362
rect 5174 10308 5180 10310
rect 5236 10308 5260 10310
rect 5316 10308 5340 10310
rect 5396 10308 5420 10310
rect 5476 10308 5482 10310
rect 5174 10299 5482 10308
rect 4804 10056 4856 10062
rect 4804 9998 4856 10004
rect 4816 9738 4844 9998
rect 4988 9920 5040 9926
rect 4988 9862 5040 9868
rect 4816 9722 4936 9738
rect 4816 9716 4948 9722
rect 4816 9710 4896 9716
rect 4252 9512 4304 9518
rect 4252 9454 4304 9460
rect 4264 9178 4292 9454
rect 4252 9172 4304 9178
rect 4252 9114 4304 9120
rect 4816 6798 4844 9710
rect 4896 9658 4948 9664
rect 5000 9654 5028 9862
rect 4988 9648 5040 9654
rect 4988 9590 5040 9596
rect 5540 9444 5592 9450
rect 5540 9386 5592 9392
rect 5174 9276 5482 9285
rect 5174 9274 5180 9276
rect 5236 9274 5260 9276
rect 5316 9274 5340 9276
rect 5396 9274 5420 9276
rect 5476 9274 5482 9276
rect 5236 9222 5238 9274
rect 5418 9222 5420 9274
rect 5174 9220 5180 9222
rect 5236 9220 5260 9222
rect 5316 9220 5340 9222
rect 5396 9220 5420 9222
rect 5476 9220 5482 9222
rect 5174 9211 5482 9220
rect 5174 8188 5482 8197
rect 5174 8186 5180 8188
rect 5236 8186 5260 8188
rect 5316 8186 5340 8188
rect 5396 8186 5420 8188
rect 5476 8186 5482 8188
rect 5236 8134 5238 8186
rect 5418 8134 5420 8186
rect 5174 8132 5180 8134
rect 5236 8132 5260 8134
rect 5316 8132 5340 8134
rect 5396 8132 5420 8134
rect 5476 8132 5482 8134
rect 5174 8123 5482 8132
rect 4896 7472 4948 7478
rect 4896 7414 4948 7420
rect 4908 6866 4936 7414
rect 5174 7100 5482 7109
rect 5174 7098 5180 7100
rect 5236 7098 5260 7100
rect 5316 7098 5340 7100
rect 5396 7098 5420 7100
rect 5476 7098 5482 7100
rect 5236 7046 5238 7098
rect 5418 7046 5420 7098
rect 5174 7044 5180 7046
rect 5236 7044 5260 7046
rect 5316 7044 5340 7046
rect 5396 7044 5420 7046
rect 5476 7044 5482 7046
rect 5174 7035 5482 7044
rect 5552 7002 5580 9386
rect 5736 8090 5764 11494
rect 6012 10674 6040 12038
rect 6380 11762 6408 12718
rect 6368 11756 6420 11762
rect 6368 11698 6420 11704
rect 6380 11354 6408 11698
rect 6368 11348 6420 11354
rect 6368 11290 6420 11296
rect 6000 10668 6052 10674
rect 6000 10610 6052 10616
rect 6472 9654 6500 13466
rect 6748 11626 6776 13806
rect 6840 12850 6868 15438
rect 6932 15434 6960 16186
rect 7024 16182 7052 16390
rect 9398 16348 9706 16357
rect 9398 16346 9404 16348
rect 9460 16346 9484 16348
rect 9540 16346 9564 16348
rect 9620 16346 9644 16348
rect 9700 16346 9706 16348
rect 9460 16294 9462 16346
rect 9642 16294 9644 16346
rect 9398 16292 9404 16294
rect 9460 16292 9484 16294
rect 9540 16292 9564 16294
rect 9620 16292 9644 16294
rect 9700 16292 9706 16294
rect 9398 16283 9706 16292
rect 11532 16250 11560 17138
rect 13622 16892 13930 16901
rect 13622 16890 13628 16892
rect 13684 16890 13708 16892
rect 13764 16890 13788 16892
rect 13844 16890 13868 16892
rect 13924 16890 13930 16892
rect 13684 16838 13686 16890
rect 13866 16838 13868 16890
rect 13622 16836 13628 16838
rect 13684 16836 13708 16838
rect 13764 16836 13788 16838
rect 13844 16836 13868 16838
rect 13924 16836 13930 16838
rect 13622 16827 13930 16836
rect 17846 16348 18154 16357
rect 17846 16346 17852 16348
rect 17908 16346 17932 16348
rect 17988 16346 18012 16348
rect 18068 16346 18092 16348
rect 18148 16346 18154 16348
rect 17908 16294 17910 16346
rect 18090 16294 18092 16346
rect 17846 16292 17852 16294
rect 17908 16292 17932 16294
rect 17988 16292 18012 16294
rect 18068 16292 18092 16294
rect 18148 16292 18154 16294
rect 17846 16283 18154 16292
rect 11520 16244 11572 16250
rect 11520 16186 11572 16192
rect 7012 16176 7064 16182
rect 7012 16118 7064 16124
rect 8024 16176 8076 16182
rect 8024 16118 8076 16124
rect 8036 15706 8064 16118
rect 17776 16108 17828 16114
rect 17776 16050 17828 16056
rect 13452 16040 13504 16046
rect 13452 15982 13504 15988
rect 13464 15706 13492 15982
rect 14372 15904 14424 15910
rect 14372 15846 14424 15852
rect 13622 15804 13930 15813
rect 13622 15802 13628 15804
rect 13684 15802 13708 15804
rect 13764 15802 13788 15804
rect 13844 15802 13868 15804
rect 13924 15802 13930 15804
rect 13684 15750 13686 15802
rect 13866 15750 13868 15802
rect 13622 15748 13628 15750
rect 13684 15748 13708 15750
rect 13764 15748 13788 15750
rect 13844 15748 13868 15750
rect 13924 15748 13930 15750
rect 13622 15739 13930 15748
rect 8024 15700 8076 15706
rect 8024 15642 8076 15648
rect 13452 15700 13504 15706
rect 13452 15642 13504 15648
rect 6920 15428 6972 15434
rect 6920 15370 6972 15376
rect 9398 15260 9706 15269
rect 9398 15258 9404 15260
rect 9460 15258 9484 15260
rect 9540 15258 9564 15260
rect 9620 15258 9644 15260
rect 9700 15258 9706 15260
rect 9460 15206 9462 15258
rect 9642 15206 9644 15258
rect 9398 15204 9404 15206
rect 9460 15204 9484 15206
rect 9540 15204 9564 15206
rect 9620 15204 9644 15206
rect 9700 15204 9706 15206
rect 9398 15195 9706 15204
rect 12440 14272 12492 14278
rect 12440 14214 12492 14220
rect 9398 14172 9706 14181
rect 9398 14170 9404 14172
rect 9460 14170 9484 14172
rect 9540 14170 9564 14172
rect 9620 14170 9644 14172
rect 9700 14170 9706 14172
rect 9460 14118 9462 14170
rect 9642 14118 9644 14170
rect 9398 14116 9404 14118
rect 9460 14116 9484 14118
rect 9540 14116 9564 14118
rect 9620 14116 9644 14118
rect 9700 14116 9706 14118
rect 9398 14107 9706 14116
rect 9398 13084 9706 13093
rect 9398 13082 9404 13084
rect 9460 13082 9484 13084
rect 9540 13082 9564 13084
rect 9620 13082 9644 13084
rect 9700 13082 9706 13084
rect 9460 13030 9462 13082
rect 9642 13030 9644 13082
rect 9398 13028 9404 13030
rect 9460 13028 9484 13030
rect 9540 13028 9564 13030
rect 9620 13028 9644 13030
rect 9700 13028 9706 13030
rect 9398 13019 9706 13028
rect 6828 12844 6880 12850
rect 6828 12786 6880 12792
rect 6840 12442 6868 12786
rect 12452 12646 12480 14214
rect 13464 12986 13492 15642
rect 14384 15570 14412 15846
rect 14372 15564 14424 15570
rect 14372 15506 14424 15512
rect 15384 15428 15436 15434
rect 15384 15370 15436 15376
rect 15396 15162 15424 15370
rect 17788 15162 17816 16050
rect 18340 16046 18368 17138
rect 20076 17060 20128 17066
rect 20076 17002 20128 17008
rect 18328 16040 18380 16046
rect 18328 15982 18380 15988
rect 18340 15706 18368 15982
rect 18328 15700 18380 15706
rect 18328 15642 18380 15648
rect 19340 15428 19392 15434
rect 19340 15370 19392 15376
rect 17846 15260 18154 15269
rect 17846 15258 17852 15260
rect 17908 15258 17932 15260
rect 17988 15258 18012 15260
rect 18068 15258 18092 15260
rect 18148 15258 18154 15260
rect 17908 15206 17910 15258
rect 18090 15206 18092 15258
rect 17846 15204 17852 15206
rect 17908 15204 17932 15206
rect 17988 15204 18012 15206
rect 18068 15204 18092 15206
rect 18148 15204 18154 15206
rect 17846 15195 18154 15204
rect 15384 15156 15436 15162
rect 15384 15098 15436 15104
rect 17776 15156 17828 15162
rect 17776 15098 17828 15104
rect 14280 15020 14332 15026
rect 14280 14962 14332 14968
rect 13622 14716 13930 14725
rect 13622 14714 13628 14716
rect 13684 14714 13708 14716
rect 13764 14714 13788 14716
rect 13844 14714 13868 14716
rect 13924 14714 13930 14716
rect 13684 14662 13686 14714
rect 13866 14662 13868 14714
rect 13622 14660 13628 14662
rect 13684 14660 13708 14662
rect 13764 14660 13788 14662
rect 13844 14660 13868 14662
rect 13924 14660 13930 14662
rect 13622 14651 13930 14660
rect 13622 13628 13930 13637
rect 13622 13626 13628 13628
rect 13684 13626 13708 13628
rect 13764 13626 13788 13628
rect 13844 13626 13868 13628
rect 13924 13626 13930 13628
rect 13684 13574 13686 13626
rect 13866 13574 13868 13626
rect 13622 13572 13628 13574
rect 13684 13572 13708 13574
rect 13764 13572 13788 13574
rect 13844 13572 13868 13574
rect 13924 13572 13930 13574
rect 13622 13563 13930 13572
rect 14292 13326 14320 14962
rect 19352 14890 19380 15370
rect 19340 14884 19392 14890
rect 19340 14826 19392 14832
rect 17846 14172 18154 14181
rect 17846 14170 17852 14172
rect 17908 14170 17932 14172
rect 17988 14170 18012 14172
rect 18068 14170 18092 14172
rect 18148 14170 18154 14172
rect 17908 14118 17910 14170
rect 18090 14118 18092 14170
rect 17846 14116 17852 14118
rect 17908 14116 17932 14118
rect 17988 14116 18012 14118
rect 18068 14116 18092 14118
rect 18148 14116 18154 14118
rect 17846 14107 18154 14116
rect 20088 13530 20116 17002
rect 22070 16892 22378 16901
rect 22070 16890 22076 16892
rect 22132 16890 22156 16892
rect 22212 16890 22236 16892
rect 22292 16890 22316 16892
rect 22372 16890 22378 16892
rect 22132 16838 22134 16890
rect 22314 16838 22316 16890
rect 22070 16836 22076 16838
rect 22132 16836 22156 16838
rect 22212 16836 22236 16838
rect 22292 16836 22316 16838
rect 22372 16836 22378 16838
rect 22070 16827 22378 16836
rect 25516 16182 25544 17138
rect 26294 16348 26602 16357
rect 26294 16346 26300 16348
rect 26356 16346 26380 16348
rect 26436 16346 26460 16348
rect 26516 16346 26540 16348
rect 26596 16346 26602 16348
rect 26356 16294 26358 16346
rect 26538 16294 26540 16346
rect 26294 16292 26300 16294
rect 26356 16292 26380 16294
rect 26436 16292 26460 16294
rect 26516 16292 26540 16294
rect 26596 16292 26602 16294
rect 26294 16283 26602 16292
rect 29932 16250 29960 17138
rect 33336 16998 33364 17138
rect 33324 16992 33376 16998
rect 33324 16934 33376 16940
rect 30518 16892 30826 16901
rect 30518 16890 30524 16892
rect 30580 16890 30604 16892
rect 30660 16890 30684 16892
rect 30740 16890 30764 16892
rect 30820 16890 30826 16892
rect 30580 16838 30582 16890
rect 30762 16838 30764 16890
rect 30518 16836 30524 16838
rect 30580 16836 30604 16838
rect 30660 16836 30684 16838
rect 30740 16836 30764 16838
rect 30820 16836 30826 16838
rect 30518 16827 30826 16836
rect 31392 16584 31444 16590
rect 31392 16526 31444 16532
rect 29920 16244 29972 16250
rect 29920 16186 29972 16192
rect 22468 16176 22520 16182
rect 22468 16118 22520 16124
rect 25504 16176 25556 16182
rect 25504 16118 25556 16124
rect 21916 16108 21968 16114
rect 21916 16050 21968 16056
rect 20628 15904 20680 15910
rect 20628 15846 20680 15852
rect 21180 15904 21232 15910
rect 21180 15846 21232 15852
rect 20640 15570 20668 15846
rect 20628 15564 20680 15570
rect 20628 15506 20680 15512
rect 20352 15496 20404 15502
rect 20352 15438 20404 15444
rect 20076 13524 20128 13530
rect 20076 13466 20128 13472
rect 14280 13320 14332 13326
rect 14280 13262 14332 13268
rect 19248 13320 19300 13326
rect 19248 13262 19300 13268
rect 14188 13184 14240 13190
rect 14188 13126 14240 13132
rect 12900 12980 12952 12986
rect 12900 12922 12952 12928
rect 13452 12980 13504 12986
rect 13452 12922 13504 12928
rect 12440 12640 12492 12646
rect 12440 12582 12492 12588
rect 6828 12436 6880 12442
rect 6828 12378 6880 12384
rect 9398 11996 9706 12005
rect 9398 11994 9404 11996
rect 9460 11994 9484 11996
rect 9540 11994 9564 11996
rect 9620 11994 9644 11996
rect 9700 11994 9706 11996
rect 9460 11942 9462 11994
rect 9642 11942 9644 11994
rect 9398 11940 9404 11942
rect 9460 11940 9484 11942
rect 9540 11940 9564 11942
rect 9620 11940 9644 11942
rect 9700 11940 9706 11942
rect 9398 11931 9706 11940
rect 6736 11620 6788 11626
rect 6736 11562 6788 11568
rect 12912 11354 12940 12922
rect 14200 12918 14228 13126
rect 14188 12912 14240 12918
rect 14188 12854 14240 12860
rect 14292 12782 14320 13262
rect 17846 13084 18154 13093
rect 17846 13082 17852 13084
rect 17908 13082 17932 13084
rect 17988 13082 18012 13084
rect 18068 13082 18092 13084
rect 18148 13082 18154 13084
rect 17908 13030 17910 13082
rect 18090 13030 18092 13082
rect 17846 13028 17852 13030
rect 17908 13028 17932 13030
rect 17988 13028 18012 13030
rect 18068 13028 18092 13030
rect 18148 13028 18154 13030
rect 17846 13019 18154 13028
rect 15292 12980 15344 12986
rect 15292 12922 15344 12928
rect 14280 12776 14332 12782
rect 14280 12718 14332 12724
rect 15304 12646 15332 12922
rect 15292 12640 15344 12646
rect 15292 12582 15344 12588
rect 13622 12540 13930 12549
rect 13622 12538 13628 12540
rect 13684 12538 13708 12540
rect 13764 12538 13788 12540
rect 13844 12538 13868 12540
rect 13924 12538 13930 12540
rect 13684 12486 13686 12538
rect 13866 12486 13868 12538
rect 13622 12484 13628 12486
rect 13684 12484 13708 12486
rect 13764 12484 13788 12486
rect 13844 12484 13868 12486
rect 13924 12484 13930 12486
rect 13622 12475 13930 12484
rect 17846 11996 18154 12005
rect 17846 11994 17852 11996
rect 17908 11994 17932 11996
rect 17988 11994 18012 11996
rect 18068 11994 18092 11996
rect 18148 11994 18154 11996
rect 17908 11942 17910 11994
rect 18090 11942 18092 11994
rect 17846 11940 17852 11942
rect 17908 11940 17932 11942
rect 17988 11940 18012 11942
rect 18068 11940 18092 11942
rect 18148 11940 18154 11942
rect 17846 11931 18154 11940
rect 13622 11452 13930 11461
rect 13622 11450 13628 11452
rect 13684 11450 13708 11452
rect 13764 11450 13788 11452
rect 13844 11450 13868 11452
rect 13924 11450 13930 11452
rect 13684 11398 13686 11450
rect 13866 11398 13868 11450
rect 13622 11396 13628 11398
rect 13684 11396 13708 11398
rect 13764 11396 13788 11398
rect 13844 11396 13868 11398
rect 13924 11396 13930 11398
rect 13622 11387 13930 11396
rect 11244 11348 11296 11354
rect 11244 11290 11296 11296
rect 12900 11348 12952 11354
rect 12900 11290 12952 11296
rect 9398 10908 9706 10917
rect 9398 10906 9404 10908
rect 9460 10906 9484 10908
rect 9540 10906 9564 10908
rect 9620 10906 9644 10908
rect 9700 10906 9706 10908
rect 9460 10854 9462 10906
rect 9642 10854 9644 10906
rect 9398 10852 9404 10854
rect 9460 10852 9484 10854
rect 9540 10852 9564 10854
rect 9620 10852 9644 10854
rect 9700 10852 9706 10854
rect 9398 10843 9706 10852
rect 11256 10266 11284 11290
rect 12624 11212 12676 11218
rect 12624 11154 12676 11160
rect 11244 10260 11296 10266
rect 11244 10202 11296 10208
rect 9398 9820 9706 9829
rect 9398 9818 9404 9820
rect 9460 9818 9484 9820
rect 9540 9818 9564 9820
rect 9620 9818 9644 9820
rect 9700 9818 9706 9820
rect 9460 9766 9462 9818
rect 9642 9766 9644 9818
rect 9398 9764 9404 9766
rect 9460 9764 9484 9766
rect 9540 9764 9564 9766
rect 9620 9764 9644 9766
rect 9700 9764 9706 9766
rect 9398 9755 9706 9764
rect 6460 9648 6512 9654
rect 6460 9590 6512 9596
rect 6472 9450 6500 9590
rect 12256 9580 12308 9586
rect 12256 9522 12308 9528
rect 6460 9444 6512 9450
rect 6460 9386 6512 9392
rect 11796 9376 11848 9382
rect 11796 9318 11848 9324
rect 10876 9172 10928 9178
rect 10876 9114 10928 9120
rect 9398 8732 9706 8741
rect 9398 8730 9404 8732
rect 9460 8730 9484 8732
rect 9540 8730 9564 8732
rect 9620 8730 9644 8732
rect 9700 8730 9706 8732
rect 9460 8678 9462 8730
rect 9642 8678 9644 8730
rect 9398 8676 9404 8678
rect 9460 8676 9484 8678
rect 9540 8676 9564 8678
rect 9620 8676 9644 8678
rect 9700 8676 9706 8678
rect 9398 8667 9706 8676
rect 10888 8090 10916 9114
rect 11808 8974 11836 9318
rect 11796 8968 11848 8974
rect 11796 8910 11848 8916
rect 11808 8498 11836 8910
rect 11796 8492 11848 8498
rect 11796 8434 11848 8440
rect 5724 8084 5776 8090
rect 5724 8026 5776 8032
rect 10876 8084 10928 8090
rect 10876 8026 10928 8032
rect 11808 7954 11836 8434
rect 11980 8424 12032 8430
rect 11980 8366 12032 8372
rect 11796 7948 11848 7954
rect 11796 7890 11848 7896
rect 10968 7880 11020 7886
rect 10968 7822 11020 7828
rect 11704 7880 11756 7886
rect 11704 7822 11756 7828
rect 9398 7644 9706 7653
rect 9398 7642 9404 7644
rect 9460 7642 9484 7644
rect 9540 7642 9564 7644
rect 9620 7642 9644 7644
rect 9700 7642 9706 7644
rect 9460 7590 9462 7642
rect 9642 7590 9644 7642
rect 9398 7588 9404 7590
rect 9460 7588 9484 7590
rect 9540 7588 9564 7590
rect 9620 7588 9644 7590
rect 9700 7588 9706 7590
rect 9398 7579 9706 7588
rect 10980 7546 11008 7822
rect 10968 7540 11020 7546
rect 10968 7482 11020 7488
rect 5632 7336 5684 7342
rect 5632 7278 5684 7284
rect 5540 6996 5592 7002
rect 5540 6938 5592 6944
rect 5644 6934 5672 7278
rect 6184 7200 6236 7206
rect 6184 7142 6236 7148
rect 5632 6928 5684 6934
rect 5632 6870 5684 6876
rect 4896 6860 4948 6866
rect 4896 6802 4948 6808
rect 5540 6860 5592 6866
rect 5540 6802 5592 6808
rect 4804 6792 4856 6798
rect 4804 6734 4856 6740
rect 4816 6458 4844 6734
rect 5552 6662 5580 6802
rect 5540 6656 5592 6662
rect 5540 6598 5592 6604
rect 4804 6452 4856 6458
rect 4804 6394 4856 6400
rect 4816 5710 4844 6394
rect 5174 6012 5482 6021
rect 5174 6010 5180 6012
rect 5236 6010 5260 6012
rect 5316 6010 5340 6012
rect 5396 6010 5420 6012
rect 5476 6010 5482 6012
rect 5236 5958 5238 6010
rect 5418 5958 5420 6010
rect 5174 5956 5180 5958
rect 5236 5956 5260 5958
rect 5316 5956 5340 5958
rect 5396 5956 5420 5958
rect 5476 5956 5482 5958
rect 5174 5947 5482 5956
rect 4804 5704 4856 5710
rect 4804 5646 4856 5652
rect 4528 5568 4580 5574
rect 4528 5510 4580 5516
rect 4540 4214 4568 5510
rect 5174 4924 5482 4933
rect 5174 4922 5180 4924
rect 5236 4922 5260 4924
rect 5316 4922 5340 4924
rect 5396 4922 5420 4924
rect 5476 4922 5482 4924
rect 5236 4870 5238 4922
rect 5418 4870 5420 4922
rect 5174 4868 5180 4870
rect 5236 4868 5260 4870
rect 5316 4868 5340 4870
rect 5396 4868 5420 4870
rect 5476 4868 5482 4870
rect 5174 4859 5482 4868
rect 4528 4208 4580 4214
rect 4528 4150 4580 4156
rect 5552 4010 5580 6598
rect 6196 5710 6224 7142
rect 9398 6556 9706 6565
rect 9398 6554 9404 6556
rect 9460 6554 9484 6556
rect 9540 6554 9564 6556
rect 9620 6554 9644 6556
rect 9700 6554 9706 6556
rect 9460 6502 9462 6554
rect 9642 6502 9644 6554
rect 9398 6500 9404 6502
rect 9460 6500 9484 6502
rect 9540 6500 9564 6502
rect 9620 6500 9644 6502
rect 9700 6500 9706 6502
rect 9398 6491 9706 6500
rect 11716 5778 11744 7822
rect 11796 7812 11848 7818
rect 11796 7754 11848 7760
rect 11808 6798 11836 7754
rect 11992 6798 12020 8366
rect 12268 7002 12296 9522
rect 12636 8974 12664 11154
rect 12716 11076 12768 11082
rect 12716 11018 12768 11024
rect 13268 11076 13320 11082
rect 13268 11018 13320 11024
rect 14372 11076 14424 11082
rect 14372 11018 14424 11024
rect 12728 10810 12756 11018
rect 12716 10804 12768 10810
rect 12716 10746 12768 10752
rect 12808 10668 12860 10674
rect 12808 10610 12860 10616
rect 12820 9722 12848 10610
rect 13280 10266 13308 11018
rect 13622 10364 13930 10373
rect 13622 10362 13628 10364
rect 13684 10362 13708 10364
rect 13764 10362 13788 10364
rect 13844 10362 13868 10364
rect 13924 10362 13930 10364
rect 13684 10310 13686 10362
rect 13866 10310 13868 10362
rect 13622 10308 13628 10310
rect 13684 10308 13708 10310
rect 13764 10308 13788 10310
rect 13844 10308 13868 10310
rect 13924 10308 13930 10310
rect 13622 10299 13930 10308
rect 13268 10260 13320 10266
rect 13268 10202 13320 10208
rect 14280 10056 14332 10062
rect 14280 9998 14332 10004
rect 13636 9920 13688 9926
rect 13636 9862 13688 9868
rect 12808 9716 12860 9722
rect 12808 9658 12860 9664
rect 13648 9586 13676 9862
rect 13636 9580 13688 9586
rect 13636 9522 13688 9528
rect 12716 9512 12768 9518
rect 12716 9454 12768 9460
rect 12728 9042 12756 9454
rect 13622 9276 13930 9285
rect 13622 9274 13628 9276
rect 13684 9274 13708 9276
rect 13764 9274 13788 9276
rect 13844 9274 13868 9276
rect 13924 9274 13930 9276
rect 13684 9222 13686 9274
rect 13866 9222 13868 9274
rect 13622 9220 13628 9222
rect 13684 9220 13708 9222
rect 13764 9220 13788 9222
rect 13844 9220 13868 9222
rect 13924 9220 13930 9222
rect 13622 9211 13930 9220
rect 12716 9036 12768 9042
rect 12716 8978 12768 8984
rect 12624 8968 12676 8974
rect 12624 8910 12676 8916
rect 12636 8498 12664 8910
rect 12624 8492 12676 8498
rect 12624 8434 12676 8440
rect 12636 8090 12664 8434
rect 12624 8084 12676 8090
rect 12624 8026 12676 8032
rect 12348 7744 12400 7750
rect 12348 7686 12400 7692
rect 12360 7410 12388 7686
rect 12348 7404 12400 7410
rect 12348 7346 12400 7352
rect 12532 7404 12584 7410
rect 12532 7346 12584 7352
rect 12624 7404 12676 7410
rect 12624 7346 12676 7352
rect 12360 7002 12388 7346
rect 12256 6996 12308 7002
rect 12256 6938 12308 6944
rect 12348 6996 12400 7002
rect 12348 6938 12400 6944
rect 11796 6792 11848 6798
rect 11796 6734 11848 6740
rect 11980 6792 12032 6798
rect 11980 6734 12032 6740
rect 11704 5772 11756 5778
rect 11704 5714 11756 5720
rect 6184 5704 6236 5710
rect 6184 5646 6236 5652
rect 6276 5636 6328 5642
rect 6276 5578 6328 5584
rect 6288 5522 6316 5578
rect 6288 5494 6408 5522
rect 6380 4554 6408 5494
rect 9398 5468 9706 5477
rect 9398 5466 9404 5468
rect 9460 5466 9484 5468
rect 9540 5466 9564 5468
rect 9620 5466 9644 5468
rect 9700 5466 9706 5468
rect 9460 5414 9462 5466
rect 9642 5414 9644 5466
rect 9398 5412 9404 5414
rect 9460 5412 9484 5414
rect 9540 5412 9564 5414
rect 9620 5412 9644 5414
rect 9700 5412 9706 5414
rect 9398 5403 9706 5412
rect 6368 4548 6420 4554
rect 6368 4490 6420 4496
rect 6380 4078 6408 4490
rect 11520 4480 11572 4486
rect 11520 4422 11572 4428
rect 9398 4380 9706 4389
rect 9398 4378 9404 4380
rect 9460 4378 9484 4380
rect 9540 4378 9564 4380
rect 9620 4378 9644 4380
rect 9700 4378 9706 4380
rect 9460 4326 9462 4378
rect 9642 4326 9644 4378
rect 9398 4324 9404 4326
rect 9460 4324 9484 4326
rect 9540 4324 9564 4326
rect 9620 4324 9644 4326
rect 9700 4324 9706 4326
rect 9398 4315 9706 4324
rect 11532 4146 11560 4422
rect 11520 4140 11572 4146
rect 11520 4082 11572 4088
rect 11808 4078 11836 6734
rect 11992 4146 12020 6734
rect 12268 6458 12296 6938
rect 12348 6860 12400 6866
rect 12348 6802 12400 6808
rect 12256 6452 12308 6458
rect 12256 6394 12308 6400
rect 12164 5568 12216 5574
rect 12164 5510 12216 5516
rect 12176 4146 12204 5510
rect 12360 5370 12388 6802
rect 12544 6322 12572 7346
rect 12532 6316 12584 6322
rect 12532 6258 12584 6264
rect 12440 6180 12492 6186
rect 12440 6122 12492 6128
rect 12452 5710 12480 6122
rect 12440 5704 12492 5710
rect 12440 5646 12492 5652
rect 12348 5364 12400 5370
rect 12348 5306 12400 5312
rect 11980 4140 12032 4146
rect 11980 4082 12032 4088
rect 12164 4140 12216 4146
rect 12164 4082 12216 4088
rect 6368 4072 6420 4078
rect 6368 4014 6420 4020
rect 11796 4072 11848 4078
rect 11796 4014 11848 4020
rect 5540 4004 5592 4010
rect 5540 3946 5592 3952
rect 11704 3936 11756 3942
rect 11704 3878 11756 3884
rect 5174 3836 5482 3845
rect 5174 3834 5180 3836
rect 5236 3834 5260 3836
rect 5316 3834 5340 3836
rect 5396 3834 5420 3836
rect 5476 3834 5482 3836
rect 5236 3782 5238 3834
rect 5418 3782 5420 3834
rect 5174 3780 5180 3782
rect 5236 3780 5260 3782
rect 5316 3780 5340 3782
rect 5396 3780 5420 3782
rect 5476 3780 5482 3782
rect 5174 3771 5482 3780
rect 5080 3596 5132 3602
rect 5080 3538 5132 3544
rect 5092 2582 5120 3538
rect 11716 3534 11744 3878
rect 11992 3670 12020 4082
rect 12176 3942 12204 4082
rect 12164 3936 12216 3942
rect 12164 3878 12216 3884
rect 11980 3664 12032 3670
rect 11980 3606 12032 3612
rect 12164 3596 12216 3602
rect 12164 3538 12216 3544
rect 6828 3528 6880 3534
rect 6828 3470 6880 3476
rect 11704 3528 11756 3534
rect 11704 3470 11756 3476
rect 5174 2748 5482 2757
rect 5174 2746 5180 2748
rect 5236 2746 5260 2748
rect 5316 2746 5340 2748
rect 5396 2746 5420 2748
rect 5476 2746 5482 2748
rect 5236 2694 5238 2746
rect 5418 2694 5420 2746
rect 5174 2692 5180 2694
rect 5236 2692 5260 2694
rect 5316 2692 5340 2694
rect 5396 2692 5420 2694
rect 5476 2692 5482 2694
rect 5174 2683 5482 2692
rect 6840 2582 6868 3470
rect 9398 3292 9706 3301
rect 9398 3290 9404 3292
rect 9460 3290 9484 3292
rect 9540 3290 9564 3292
rect 9620 3290 9644 3292
rect 9700 3290 9706 3292
rect 9460 3238 9462 3290
rect 9642 3238 9644 3290
rect 9398 3236 9404 3238
rect 9460 3236 9484 3238
rect 9540 3236 9564 3238
rect 9620 3236 9644 3238
rect 9700 3236 9706 3238
rect 9398 3227 9706 3236
rect 12176 3058 12204 3538
rect 12360 3398 12388 5306
rect 12452 5234 12480 5646
rect 12440 5228 12492 5234
rect 12440 5170 12492 5176
rect 12544 5166 12572 6258
rect 12532 5160 12584 5166
rect 12532 5102 12584 5108
rect 12544 4758 12572 5102
rect 12532 4752 12584 4758
rect 12532 4694 12584 4700
rect 12636 4690 12664 7346
rect 12728 7274 12756 8978
rect 14292 8634 14320 9998
rect 14384 9994 14412 11018
rect 17846 10908 18154 10917
rect 17846 10906 17852 10908
rect 17908 10906 17932 10908
rect 17988 10906 18012 10908
rect 18068 10906 18092 10908
rect 18148 10906 18154 10908
rect 17908 10854 17910 10906
rect 18090 10854 18092 10906
rect 17846 10852 17852 10854
rect 17908 10852 17932 10854
rect 17988 10852 18012 10854
rect 18068 10852 18092 10854
rect 18148 10852 18154 10854
rect 17846 10843 18154 10852
rect 19260 10810 19288 13262
rect 20088 12782 20116 13466
rect 20260 12980 20312 12986
rect 20260 12922 20312 12928
rect 20076 12776 20128 12782
rect 20076 12718 20128 12724
rect 19248 10804 19300 10810
rect 19248 10746 19300 10752
rect 17684 10668 17736 10674
rect 17684 10610 17736 10616
rect 17696 10130 17724 10610
rect 20088 10266 20116 12718
rect 20272 12102 20300 12922
rect 20260 12096 20312 12102
rect 20260 12038 20312 12044
rect 20364 10674 20392 15438
rect 21192 14958 21220 15846
rect 21928 15162 21956 16050
rect 22070 15804 22378 15813
rect 22070 15802 22076 15804
rect 22132 15802 22156 15804
rect 22212 15802 22236 15804
rect 22292 15802 22316 15804
rect 22372 15802 22378 15804
rect 22132 15750 22134 15802
rect 22314 15750 22316 15802
rect 22070 15748 22076 15750
rect 22132 15748 22156 15750
rect 22212 15748 22236 15750
rect 22292 15748 22316 15750
rect 22372 15748 22378 15750
rect 22070 15739 22378 15748
rect 22480 15706 22508 16118
rect 29092 15904 29144 15910
rect 29092 15846 29144 15852
rect 22468 15700 22520 15706
rect 22468 15642 22520 15648
rect 26294 15260 26602 15269
rect 26294 15258 26300 15260
rect 26356 15258 26380 15260
rect 26436 15258 26460 15260
rect 26516 15258 26540 15260
rect 26596 15258 26602 15260
rect 26356 15206 26358 15258
rect 26538 15206 26540 15258
rect 26294 15204 26300 15206
rect 26356 15204 26380 15206
rect 26436 15204 26460 15206
rect 26516 15204 26540 15206
rect 26596 15204 26602 15206
rect 26294 15195 26602 15204
rect 21916 15156 21968 15162
rect 21916 15098 21968 15104
rect 24860 15088 24912 15094
rect 24860 15030 24912 15036
rect 21180 14952 21232 14958
rect 21180 14894 21232 14900
rect 20720 13184 20772 13190
rect 20720 13126 20772 13132
rect 20732 12646 20760 13126
rect 21192 12986 21220 14894
rect 22070 14716 22378 14725
rect 22070 14714 22076 14716
rect 22132 14714 22156 14716
rect 22212 14714 22236 14716
rect 22292 14714 22316 14716
rect 22372 14714 22378 14716
rect 22132 14662 22134 14714
rect 22314 14662 22316 14714
rect 22070 14660 22076 14662
rect 22132 14660 22156 14662
rect 22212 14660 22236 14662
rect 22292 14660 22316 14662
rect 22372 14660 22378 14662
rect 22070 14651 22378 14660
rect 22070 13628 22378 13637
rect 22070 13626 22076 13628
rect 22132 13626 22156 13628
rect 22212 13626 22236 13628
rect 22292 13626 22316 13628
rect 22372 13626 22378 13628
rect 22132 13574 22134 13626
rect 22314 13574 22316 13626
rect 22070 13572 22076 13574
rect 22132 13572 22156 13574
rect 22212 13572 22236 13574
rect 22292 13572 22316 13574
rect 22372 13572 22378 13574
rect 22070 13563 22378 13572
rect 24872 13530 24900 15030
rect 29104 14958 29132 15846
rect 29932 15162 29960 16186
rect 30518 15804 30826 15813
rect 30518 15802 30524 15804
rect 30580 15802 30604 15804
rect 30660 15802 30684 15804
rect 30740 15802 30764 15804
rect 30820 15802 30826 15804
rect 30580 15750 30582 15802
rect 30762 15750 30764 15802
rect 30518 15748 30524 15750
rect 30580 15748 30604 15750
rect 30660 15748 30684 15750
rect 30740 15748 30764 15750
rect 30820 15748 30826 15750
rect 30518 15739 30826 15748
rect 29920 15156 29972 15162
rect 29920 15098 29972 15104
rect 28080 14952 28132 14958
rect 28080 14894 28132 14900
rect 29092 14952 29144 14958
rect 29092 14894 29144 14900
rect 26294 14172 26602 14181
rect 26294 14170 26300 14172
rect 26356 14170 26380 14172
rect 26436 14170 26460 14172
rect 26516 14170 26540 14172
rect 26596 14170 26602 14172
rect 26356 14118 26358 14170
rect 26538 14118 26540 14170
rect 26294 14116 26300 14118
rect 26356 14116 26380 14118
rect 26436 14116 26460 14118
rect 26516 14116 26540 14118
rect 26596 14116 26602 14118
rect 26294 14107 26602 14116
rect 28092 13938 28120 14894
rect 29644 14816 29696 14822
rect 29644 14758 29696 14764
rect 29000 14000 29052 14006
rect 29000 13942 29052 13948
rect 28080 13932 28132 13938
rect 28080 13874 28132 13880
rect 24860 13524 24912 13530
rect 24860 13466 24912 13472
rect 26294 13084 26602 13093
rect 26294 13082 26300 13084
rect 26356 13082 26380 13084
rect 26436 13082 26460 13084
rect 26516 13082 26540 13084
rect 26596 13082 26602 13084
rect 26356 13030 26358 13082
rect 26538 13030 26540 13082
rect 26294 13028 26300 13030
rect 26356 13028 26380 13030
rect 26436 13028 26460 13030
rect 26516 13028 26540 13030
rect 26596 13028 26602 13030
rect 26294 13019 26602 13028
rect 21180 12980 21232 12986
rect 21180 12922 21232 12928
rect 20812 12844 20864 12850
rect 20812 12786 20864 12792
rect 27896 12844 27948 12850
rect 27896 12786 27948 12792
rect 20720 12640 20772 12646
rect 20720 12582 20772 12588
rect 20732 11762 20760 12582
rect 20824 12442 20852 12786
rect 21088 12776 21140 12782
rect 21088 12718 21140 12724
rect 20812 12436 20864 12442
rect 20812 12378 20864 12384
rect 20720 11756 20772 11762
rect 20720 11698 20772 11704
rect 20732 11286 20760 11698
rect 21100 11558 21128 12718
rect 22836 12640 22888 12646
rect 22836 12582 22888 12588
rect 22070 12540 22378 12549
rect 22070 12538 22076 12540
rect 22132 12538 22156 12540
rect 22212 12538 22236 12540
rect 22292 12538 22316 12540
rect 22372 12538 22378 12540
rect 22132 12486 22134 12538
rect 22314 12486 22316 12538
rect 22070 12484 22076 12486
rect 22132 12484 22156 12486
rect 22212 12484 22236 12486
rect 22292 12484 22316 12486
rect 22372 12484 22378 12486
rect 22070 12475 22378 12484
rect 21272 12300 21324 12306
rect 21272 12242 21324 12248
rect 21284 11626 21312 12242
rect 21640 12164 21692 12170
rect 21640 12106 21692 12112
rect 21272 11620 21324 11626
rect 21272 11562 21324 11568
rect 21088 11552 21140 11558
rect 21088 11494 21140 11500
rect 21272 11348 21324 11354
rect 21272 11290 21324 11296
rect 20720 11280 20772 11286
rect 20720 11222 20772 11228
rect 20352 10668 20404 10674
rect 20352 10610 20404 10616
rect 20076 10260 20128 10266
rect 20076 10202 20128 10208
rect 21284 10130 21312 11290
rect 17684 10124 17736 10130
rect 17684 10066 17736 10072
rect 21272 10124 21324 10130
rect 21272 10066 21324 10072
rect 20996 10056 21048 10062
rect 20996 9998 21048 10004
rect 14372 9988 14424 9994
rect 14372 9930 14424 9936
rect 14384 9722 14412 9930
rect 15384 9920 15436 9926
rect 15384 9862 15436 9868
rect 14372 9716 14424 9722
rect 14372 9658 14424 9664
rect 14280 8628 14332 8634
rect 14280 8570 14332 8576
rect 13544 8492 13596 8498
rect 13544 8434 13596 8440
rect 12716 7268 12768 7274
rect 12716 7210 12768 7216
rect 12808 5228 12860 5234
rect 12808 5170 12860 5176
rect 12440 4684 12492 4690
rect 12440 4626 12492 4632
rect 12624 4684 12676 4690
rect 12624 4626 12676 4632
rect 12452 4146 12480 4626
rect 12820 4622 12848 5170
rect 12808 4616 12860 4622
rect 12808 4558 12860 4564
rect 12820 4282 12848 4558
rect 12808 4276 12860 4282
rect 12808 4218 12860 4224
rect 12624 4208 12676 4214
rect 12624 4150 12676 4156
rect 12440 4140 12492 4146
rect 12440 4082 12492 4088
rect 12532 3460 12584 3466
rect 12532 3402 12584 3408
rect 12348 3392 12400 3398
rect 12348 3334 12400 3340
rect 12544 3194 12572 3402
rect 12532 3188 12584 3194
rect 12532 3130 12584 3136
rect 12636 3058 12664 4150
rect 12808 4140 12860 4146
rect 12808 4082 12860 4088
rect 12716 4004 12768 4010
rect 12716 3946 12768 3952
rect 12728 3534 12756 3946
rect 12820 3602 12848 4082
rect 13556 4026 13584 8434
rect 13622 8188 13930 8197
rect 13622 8186 13628 8188
rect 13684 8186 13708 8188
rect 13764 8186 13788 8188
rect 13844 8186 13868 8188
rect 13924 8186 13930 8188
rect 13684 8134 13686 8186
rect 13866 8134 13868 8186
rect 13622 8132 13628 8134
rect 13684 8132 13708 8134
rect 13764 8132 13788 8134
rect 13844 8132 13868 8134
rect 13924 8132 13930 8134
rect 13622 8123 13930 8132
rect 14292 7410 14320 8570
rect 14280 7404 14332 7410
rect 14280 7346 14332 7352
rect 14740 7404 14792 7410
rect 14740 7346 14792 7352
rect 13622 7100 13930 7109
rect 13622 7098 13628 7100
rect 13684 7098 13708 7100
rect 13764 7098 13788 7100
rect 13844 7098 13868 7100
rect 13924 7098 13930 7100
rect 13684 7046 13686 7098
rect 13866 7046 13868 7098
rect 13622 7044 13628 7046
rect 13684 7044 13708 7046
rect 13764 7044 13788 7046
rect 13844 7044 13868 7046
rect 13924 7044 13930 7046
rect 13622 7035 13930 7044
rect 13622 6012 13930 6021
rect 13622 6010 13628 6012
rect 13684 6010 13708 6012
rect 13764 6010 13788 6012
rect 13844 6010 13868 6012
rect 13924 6010 13930 6012
rect 13684 5958 13686 6010
rect 13866 5958 13868 6010
rect 13622 5956 13628 5958
rect 13684 5956 13708 5958
rect 13764 5956 13788 5958
rect 13844 5956 13868 5958
rect 13924 5956 13930 5958
rect 13622 5947 13930 5956
rect 13622 4924 13930 4933
rect 13622 4922 13628 4924
rect 13684 4922 13708 4924
rect 13764 4922 13788 4924
rect 13844 4922 13868 4924
rect 13924 4922 13930 4924
rect 13684 4870 13686 4922
rect 13866 4870 13868 4922
rect 13622 4868 13628 4870
rect 13684 4868 13708 4870
rect 13764 4868 13788 4870
rect 13844 4868 13868 4870
rect 13924 4868 13930 4870
rect 13622 4859 13930 4868
rect 13820 4072 13872 4078
rect 13556 4020 13820 4026
rect 13556 4014 13872 4020
rect 13556 3998 13860 4014
rect 12808 3596 12860 3602
rect 12808 3538 12860 3544
rect 12716 3528 12768 3534
rect 12716 3470 12768 3476
rect 12164 3052 12216 3058
rect 12164 2994 12216 3000
rect 12624 3052 12676 3058
rect 12624 2994 12676 3000
rect 13556 2854 13584 3998
rect 14752 3942 14780 7346
rect 14740 3936 14792 3942
rect 14740 3878 14792 3884
rect 13622 3836 13930 3845
rect 13622 3834 13628 3836
rect 13684 3834 13708 3836
rect 13764 3834 13788 3836
rect 13844 3834 13868 3836
rect 13924 3834 13930 3836
rect 13684 3782 13686 3834
rect 13866 3782 13868 3834
rect 13622 3780 13628 3782
rect 13684 3780 13708 3782
rect 13764 3780 13788 3782
rect 13844 3780 13868 3782
rect 13924 3780 13930 3782
rect 13622 3771 13930 3780
rect 13544 2848 13596 2854
rect 13544 2790 13596 2796
rect 13622 2748 13930 2757
rect 13622 2746 13628 2748
rect 13684 2746 13708 2748
rect 13764 2746 13788 2748
rect 13844 2746 13868 2748
rect 13924 2746 13930 2748
rect 13684 2694 13686 2746
rect 13866 2694 13868 2746
rect 13622 2692 13628 2694
rect 13684 2692 13708 2694
rect 13764 2692 13788 2694
rect 13844 2692 13868 2694
rect 13924 2692 13930 2694
rect 13622 2683 13930 2692
rect 15396 2650 15424 9862
rect 17846 9820 18154 9829
rect 17846 9818 17852 9820
rect 17908 9818 17932 9820
rect 17988 9818 18012 9820
rect 18068 9818 18092 9820
rect 18148 9818 18154 9820
rect 17908 9766 17910 9818
rect 18090 9766 18092 9818
rect 17846 9764 17852 9766
rect 17908 9764 17932 9766
rect 17988 9764 18012 9766
rect 18068 9764 18092 9766
rect 18148 9764 18154 9766
rect 17846 9755 18154 9764
rect 17846 8732 18154 8741
rect 17846 8730 17852 8732
rect 17908 8730 17932 8732
rect 17988 8730 18012 8732
rect 18068 8730 18092 8732
rect 18148 8730 18154 8732
rect 17908 8678 17910 8730
rect 18090 8678 18092 8730
rect 17846 8676 17852 8678
rect 17908 8676 17932 8678
rect 17988 8676 18012 8678
rect 18068 8676 18092 8678
rect 18148 8676 18154 8678
rect 17846 8667 18154 8676
rect 20260 7948 20312 7954
rect 20260 7890 20312 7896
rect 19340 7880 19392 7886
rect 19340 7822 19392 7828
rect 19800 7880 19852 7886
rect 19800 7822 19852 7828
rect 17846 7644 18154 7653
rect 17846 7642 17852 7644
rect 17908 7642 17932 7644
rect 17988 7642 18012 7644
rect 18068 7642 18092 7644
rect 18148 7642 18154 7644
rect 17908 7590 17910 7642
rect 18090 7590 18092 7642
rect 17846 7588 17852 7590
rect 17908 7588 17932 7590
rect 17988 7588 18012 7590
rect 18068 7588 18092 7590
rect 18148 7588 18154 7590
rect 17846 7579 18154 7588
rect 17846 6556 18154 6565
rect 17846 6554 17852 6556
rect 17908 6554 17932 6556
rect 17988 6554 18012 6556
rect 18068 6554 18092 6556
rect 18148 6554 18154 6556
rect 17908 6502 17910 6554
rect 18090 6502 18092 6554
rect 17846 6500 17852 6502
rect 17908 6500 17932 6502
rect 17988 6500 18012 6502
rect 18068 6500 18092 6502
rect 18148 6500 18154 6502
rect 17846 6491 18154 6500
rect 17846 5468 18154 5477
rect 17846 5466 17852 5468
rect 17908 5466 17932 5468
rect 17988 5466 18012 5468
rect 18068 5466 18092 5468
rect 18148 5466 18154 5468
rect 17908 5414 17910 5466
rect 18090 5414 18092 5466
rect 17846 5412 17852 5414
rect 17908 5412 17932 5414
rect 17988 5412 18012 5414
rect 18068 5412 18092 5414
rect 18148 5412 18154 5414
rect 17846 5403 18154 5412
rect 19352 4690 19380 7822
rect 19812 7274 19840 7822
rect 19800 7268 19852 7274
rect 19800 7210 19852 7216
rect 20272 7002 20300 7890
rect 20812 7880 20864 7886
rect 20812 7822 20864 7828
rect 20352 7268 20404 7274
rect 20352 7210 20404 7216
rect 20260 6996 20312 7002
rect 20260 6938 20312 6944
rect 20272 6798 20300 6938
rect 20168 6792 20220 6798
rect 20168 6734 20220 6740
rect 20260 6792 20312 6798
rect 20260 6734 20312 6740
rect 19616 5228 19668 5234
rect 19616 5170 19668 5176
rect 19628 4826 19656 5170
rect 19616 4820 19668 4826
rect 19616 4762 19668 4768
rect 19340 4684 19392 4690
rect 19340 4626 19392 4632
rect 20180 4622 20208 6734
rect 20364 6662 20392 7210
rect 20824 7206 20852 7822
rect 21008 7818 21036 9998
rect 21284 9042 21312 10066
rect 21272 9036 21324 9042
rect 21272 8978 21324 8984
rect 20996 7812 21048 7818
rect 20996 7754 21048 7760
rect 20812 7200 20864 7206
rect 20812 7142 20864 7148
rect 20824 7002 20852 7142
rect 20812 6996 20864 7002
rect 20812 6938 20864 6944
rect 20352 6656 20404 6662
rect 20352 6598 20404 6604
rect 17132 4616 17184 4622
rect 17132 4558 17184 4564
rect 20168 4616 20220 4622
rect 20168 4558 20220 4564
rect 15660 4548 15712 4554
rect 15660 4490 15712 4496
rect 15672 4010 15700 4490
rect 17144 4078 17172 4558
rect 17846 4380 18154 4389
rect 17846 4378 17852 4380
rect 17908 4378 17932 4380
rect 17988 4378 18012 4380
rect 18068 4378 18092 4380
rect 18148 4378 18154 4380
rect 17908 4326 17910 4378
rect 18090 4326 18092 4378
rect 17846 4324 17852 4326
rect 17908 4324 17932 4326
rect 17988 4324 18012 4326
rect 18068 4324 18092 4326
rect 18148 4324 18154 4326
rect 17846 4315 18154 4324
rect 17132 4072 17184 4078
rect 17132 4014 17184 4020
rect 15660 4004 15712 4010
rect 15660 3946 15712 3952
rect 15672 3670 15700 3946
rect 21652 3738 21680 12106
rect 22070 11452 22378 11461
rect 22070 11450 22076 11452
rect 22132 11450 22156 11452
rect 22212 11450 22236 11452
rect 22292 11450 22316 11452
rect 22372 11450 22378 11452
rect 22132 11398 22134 11450
rect 22314 11398 22316 11450
rect 22070 11396 22076 11398
rect 22132 11396 22156 11398
rect 22212 11396 22236 11398
rect 22292 11396 22316 11398
rect 22372 11396 22378 11398
rect 22070 11387 22378 11396
rect 22070 10364 22378 10373
rect 22070 10362 22076 10364
rect 22132 10362 22156 10364
rect 22212 10362 22236 10364
rect 22292 10362 22316 10364
rect 22372 10362 22378 10364
rect 22132 10310 22134 10362
rect 22314 10310 22316 10362
rect 22070 10308 22076 10310
rect 22132 10308 22156 10310
rect 22212 10308 22236 10310
rect 22292 10308 22316 10310
rect 22372 10308 22378 10310
rect 22070 10299 22378 10308
rect 22070 9276 22378 9285
rect 22070 9274 22076 9276
rect 22132 9274 22156 9276
rect 22212 9274 22236 9276
rect 22292 9274 22316 9276
rect 22372 9274 22378 9276
rect 22132 9222 22134 9274
rect 22314 9222 22316 9274
rect 22070 9220 22076 9222
rect 22132 9220 22156 9222
rect 22212 9220 22236 9222
rect 22292 9220 22316 9222
rect 22372 9220 22378 9222
rect 22070 9211 22378 9220
rect 21732 9036 21784 9042
rect 21732 8978 21784 8984
rect 21744 5302 21772 8978
rect 22848 8974 22876 12582
rect 27908 12238 27936 12786
rect 28092 12434 28120 13874
rect 28356 13864 28408 13870
rect 28356 13806 28408 13812
rect 28368 13530 28396 13806
rect 28356 13524 28408 13530
rect 28356 13466 28408 13472
rect 29012 12986 29040 13942
rect 29000 12980 29052 12986
rect 29000 12922 29052 12928
rect 28000 12406 28120 12434
rect 27896 12232 27948 12238
rect 27896 12174 27948 12180
rect 26294 11996 26602 12005
rect 26294 11994 26300 11996
rect 26356 11994 26380 11996
rect 26436 11994 26460 11996
rect 26516 11994 26540 11996
rect 26596 11994 26602 11996
rect 26356 11942 26358 11994
rect 26538 11942 26540 11994
rect 26294 11940 26300 11942
rect 26356 11940 26380 11942
rect 26436 11940 26460 11942
rect 26516 11940 26540 11942
rect 26596 11940 26602 11942
rect 26294 11931 26602 11940
rect 27908 11354 27936 12174
rect 27896 11348 27948 11354
rect 27896 11290 27948 11296
rect 27908 11150 27936 11290
rect 27896 11144 27948 11150
rect 27896 11086 27948 11092
rect 26294 10908 26602 10917
rect 26294 10906 26300 10908
rect 26356 10906 26380 10908
rect 26436 10906 26460 10908
rect 26516 10906 26540 10908
rect 26596 10906 26602 10908
rect 26356 10854 26358 10906
rect 26538 10854 26540 10906
rect 26294 10852 26300 10854
rect 26356 10852 26380 10854
rect 26436 10852 26460 10854
rect 26516 10852 26540 10854
rect 26596 10852 26602 10854
rect 26294 10843 26602 10852
rect 27804 10668 27856 10674
rect 27804 10610 27856 10616
rect 26294 9820 26602 9829
rect 26294 9818 26300 9820
rect 26356 9818 26380 9820
rect 26436 9818 26460 9820
rect 26516 9818 26540 9820
rect 26596 9818 26602 9820
rect 26356 9766 26358 9818
rect 26538 9766 26540 9818
rect 26294 9764 26300 9766
rect 26356 9764 26380 9766
rect 26436 9764 26460 9766
rect 26516 9764 26540 9766
rect 26596 9764 26602 9766
rect 26294 9755 26602 9764
rect 21916 8968 21968 8974
rect 21916 8910 21968 8916
rect 22836 8968 22888 8974
rect 22836 8910 22888 8916
rect 26700 8968 26752 8974
rect 26700 8910 26752 8916
rect 21928 7954 21956 8910
rect 26294 8732 26602 8741
rect 26294 8730 26300 8732
rect 26356 8730 26380 8732
rect 26436 8730 26460 8732
rect 26516 8730 26540 8732
rect 26596 8730 26602 8732
rect 26356 8678 26358 8730
rect 26538 8678 26540 8730
rect 26294 8676 26300 8678
rect 26356 8676 26380 8678
rect 26436 8676 26460 8678
rect 26516 8676 26540 8678
rect 26596 8676 26602 8678
rect 26294 8667 26602 8676
rect 22070 8188 22378 8197
rect 22070 8186 22076 8188
rect 22132 8186 22156 8188
rect 22212 8186 22236 8188
rect 22292 8186 22316 8188
rect 22372 8186 22378 8188
rect 22132 8134 22134 8186
rect 22314 8134 22316 8186
rect 22070 8132 22076 8134
rect 22132 8132 22156 8134
rect 22212 8132 22236 8134
rect 22292 8132 22316 8134
rect 22372 8132 22378 8134
rect 22070 8123 22378 8132
rect 26712 8022 26740 8910
rect 27816 8498 27844 10610
rect 27908 9178 27936 11086
rect 28000 10674 28028 12406
rect 29000 11076 29052 11082
rect 29000 11018 29052 11024
rect 29012 10742 29040 11018
rect 29000 10736 29052 10742
rect 29000 10678 29052 10684
rect 27988 10668 28040 10674
rect 27988 10610 28040 10616
rect 27896 9172 27948 9178
rect 27896 9114 27948 9120
rect 28724 8832 28776 8838
rect 28724 8774 28776 8780
rect 28736 8566 28764 8774
rect 28724 8560 28776 8566
rect 28724 8502 28776 8508
rect 27804 8492 27856 8498
rect 27804 8434 27856 8440
rect 28080 8424 28132 8430
rect 28080 8366 28132 8372
rect 27344 8288 27396 8294
rect 27344 8230 27396 8236
rect 26700 8016 26752 8022
rect 26700 7958 26752 7964
rect 21916 7948 21968 7954
rect 21916 7890 21968 7896
rect 24768 7744 24820 7750
rect 24768 7686 24820 7692
rect 22070 7100 22378 7109
rect 22070 7098 22076 7100
rect 22132 7098 22156 7100
rect 22212 7098 22236 7100
rect 22292 7098 22316 7100
rect 22372 7098 22378 7100
rect 22132 7046 22134 7098
rect 22314 7046 22316 7098
rect 22070 7044 22076 7046
rect 22132 7044 22156 7046
rect 22212 7044 22236 7046
rect 22292 7044 22316 7046
rect 22372 7044 22378 7046
rect 22070 7035 22378 7044
rect 23204 6656 23256 6662
rect 23204 6598 23256 6604
rect 22070 6012 22378 6021
rect 22070 6010 22076 6012
rect 22132 6010 22156 6012
rect 22212 6010 22236 6012
rect 22292 6010 22316 6012
rect 22372 6010 22378 6012
rect 22132 5958 22134 6010
rect 22314 5958 22316 6010
rect 22070 5956 22076 5958
rect 22132 5956 22156 5958
rect 22212 5956 22236 5958
rect 22292 5956 22316 5958
rect 22372 5956 22378 5958
rect 22070 5947 22378 5956
rect 21732 5296 21784 5302
rect 21732 5238 21784 5244
rect 23216 5234 23244 6598
rect 24780 6322 24808 7686
rect 26294 7644 26602 7653
rect 26294 7642 26300 7644
rect 26356 7642 26380 7644
rect 26436 7642 26460 7644
rect 26516 7642 26540 7644
rect 26596 7642 26602 7644
rect 26356 7590 26358 7642
rect 26538 7590 26540 7642
rect 26294 7588 26300 7590
rect 26356 7588 26380 7590
rect 26436 7588 26460 7590
rect 26516 7588 26540 7590
rect 26596 7588 26602 7590
rect 26294 7579 26602 7588
rect 26712 7546 26740 7958
rect 27356 7546 27384 8230
rect 28092 8090 28120 8366
rect 28080 8084 28132 8090
rect 28080 8026 28132 8032
rect 27712 7880 27764 7886
rect 27712 7822 27764 7828
rect 27724 7546 27752 7822
rect 26700 7540 26752 7546
rect 26700 7482 26752 7488
rect 27344 7540 27396 7546
rect 27344 7482 27396 7488
rect 27712 7540 27764 7546
rect 27712 7482 27764 7488
rect 26712 7342 26740 7482
rect 26700 7336 26752 7342
rect 26700 7278 26752 7284
rect 27252 7336 27304 7342
rect 27252 7278 27304 7284
rect 26294 6556 26602 6565
rect 26294 6554 26300 6556
rect 26356 6554 26380 6556
rect 26436 6554 26460 6556
rect 26516 6554 26540 6556
rect 26596 6554 26602 6556
rect 26356 6502 26358 6554
rect 26538 6502 26540 6554
rect 26294 6500 26300 6502
rect 26356 6500 26380 6502
rect 26436 6500 26460 6502
rect 26516 6500 26540 6502
rect 26596 6500 26602 6502
rect 26294 6491 26602 6500
rect 24768 6316 24820 6322
rect 24768 6258 24820 6264
rect 26294 5468 26602 5477
rect 26294 5466 26300 5468
rect 26356 5466 26380 5468
rect 26436 5466 26460 5468
rect 26516 5466 26540 5468
rect 26596 5466 26602 5468
rect 26356 5414 26358 5466
rect 26538 5414 26540 5466
rect 26294 5412 26300 5414
rect 26356 5412 26380 5414
rect 26436 5412 26460 5414
rect 26516 5412 26540 5414
rect 26596 5412 26602 5414
rect 26294 5403 26602 5412
rect 23204 5228 23256 5234
rect 23204 5170 23256 5176
rect 24584 5024 24636 5030
rect 24584 4966 24636 4972
rect 22070 4924 22378 4933
rect 22070 4922 22076 4924
rect 22132 4922 22156 4924
rect 22212 4922 22236 4924
rect 22292 4922 22316 4924
rect 22372 4922 22378 4924
rect 22132 4870 22134 4922
rect 22314 4870 22316 4922
rect 22070 4868 22076 4870
rect 22132 4868 22156 4870
rect 22212 4868 22236 4870
rect 22292 4868 22316 4870
rect 22372 4868 22378 4870
rect 22070 4859 22378 4868
rect 24596 3942 24624 4966
rect 26294 4380 26602 4389
rect 26294 4378 26300 4380
rect 26356 4378 26380 4380
rect 26436 4378 26460 4380
rect 26516 4378 26540 4380
rect 26596 4378 26602 4380
rect 26356 4326 26358 4378
rect 26538 4326 26540 4378
rect 26294 4324 26300 4326
rect 26356 4324 26380 4326
rect 26436 4324 26460 4326
rect 26516 4324 26540 4326
rect 26596 4324 26602 4326
rect 26294 4315 26602 4324
rect 24584 3936 24636 3942
rect 24584 3878 24636 3884
rect 22070 3836 22378 3845
rect 22070 3834 22076 3836
rect 22132 3834 22156 3836
rect 22212 3834 22236 3836
rect 22292 3834 22316 3836
rect 22372 3834 22378 3836
rect 22132 3782 22134 3834
rect 22314 3782 22316 3834
rect 22070 3780 22076 3782
rect 22132 3780 22156 3782
rect 22212 3780 22236 3782
rect 22292 3780 22316 3782
rect 22372 3780 22378 3782
rect 22070 3771 22378 3780
rect 24596 3738 24624 3878
rect 27264 3738 27292 7278
rect 29552 5296 29604 5302
rect 29552 5238 29604 5244
rect 29564 4690 29592 5238
rect 29552 4684 29604 4690
rect 29552 4626 29604 4632
rect 29656 3738 29684 14758
rect 30518 14716 30826 14725
rect 30518 14714 30524 14716
rect 30580 14714 30604 14716
rect 30660 14714 30684 14716
rect 30740 14714 30764 14716
rect 30820 14714 30826 14716
rect 30580 14662 30582 14714
rect 30762 14662 30764 14714
rect 30518 14660 30524 14662
rect 30580 14660 30604 14662
rect 30660 14660 30684 14662
rect 30740 14660 30764 14662
rect 30820 14660 30826 14662
rect 30518 14651 30826 14660
rect 31404 14074 31432 16526
rect 31392 14068 31444 14074
rect 31392 14010 31444 14016
rect 30518 13628 30826 13637
rect 30518 13626 30524 13628
rect 30580 13626 30604 13628
rect 30660 13626 30684 13628
rect 30740 13626 30764 13628
rect 30820 13626 30826 13628
rect 30580 13574 30582 13626
rect 30762 13574 30764 13626
rect 30518 13572 30524 13574
rect 30580 13572 30604 13574
rect 30660 13572 30684 13574
rect 30740 13572 30764 13574
rect 30820 13572 30826 13574
rect 30518 13563 30826 13572
rect 30380 13456 30432 13462
rect 30380 13398 30432 13404
rect 30392 13190 30420 13398
rect 31404 13326 31432 14010
rect 31484 13932 31536 13938
rect 31484 13874 31536 13880
rect 31496 13394 31524 13874
rect 31484 13388 31536 13394
rect 31484 13330 31536 13336
rect 31392 13320 31444 13326
rect 31392 13262 31444 13268
rect 30380 13184 30432 13190
rect 30380 13126 30432 13132
rect 30392 11082 30420 13126
rect 30518 12540 30826 12549
rect 30518 12538 30524 12540
rect 30580 12538 30604 12540
rect 30660 12538 30684 12540
rect 30740 12538 30764 12540
rect 30820 12538 30826 12540
rect 30580 12486 30582 12538
rect 30762 12486 30764 12538
rect 30518 12484 30524 12486
rect 30580 12484 30604 12486
rect 30660 12484 30684 12486
rect 30740 12484 30764 12486
rect 30820 12484 30826 12486
rect 30518 12475 30826 12484
rect 31496 12434 31524 13330
rect 31404 12406 31524 12434
rect 30518 11452 30826 11461
rect 30518 11450 30524 11452
rect 30580 11450 30604 11452
rect 30660 11450 30684 11452
rect 30740 11450 30764 11452
rect 30820 11450 30826 11452
rect 30580 11398 30582 11450
rect 30762 11398 30764 11450
rect 30518 11396 30524 11398
rect 30580 11396 30604 11398
rect 30660 11396 30684 11398
rect 30740 11396 30764 11398
rect 30820 11396 30826 11398
rect 30518 11387 30826 11396
rect 31404 11082 31432 12406
rect 33336 12102 33364 16934
rect 34060 16448 34112 16454
rect 34060 16390 34112 16396
rect 34072 16153 34100 16390
rect 34058 16144 34114 16153
rect 34058 16079 34114 16088
rect 34060 13728 34112 13734
rect 34058 13696 34060 13705
rect 34112 13696 34114 13705
rect 34058 13631 34114 13640
rect 33324 12096 33376 12102
rect 33324 12038 33376 12044
rect 31484 11756 31536 11762
rect 31484 11698 31536 11704
rect 31496 11082 31524 11698
rect 34060 11552 34112 11558
rect 34060 11494 34112 11500
rect 34072 11257 34100 11494
rect 34058 11248 34114 11257
rect 34058 11183 34114 11192
rect 30380 11076 30432 11082
rect 30380 11018 30432 11024
rect 31392 11076 31444 11082
rect 31392 11018 31444 11024
rect 31484 11076 31536 11082
rect 31484 11018 31536 11024
rect 29736 11008 29788 11014
rect 29736 10950 29788 10956
rect 29748 10606 29776 10950
rect 29736 10600 29788 10606
rect 29736 10542 29788 10548
rect 30392 8022 30420 11018
rect 31404 10810 31432 11018
rect 31392 10804 31444 10810
rect 31392 10746 31444 10752
rect 30518 10364 30826 10373
rect 30518 10362 30524 10364
rect 30580 10362 30604 10364
rect 30660 10362 30684 10364
rect 30740 10362 30764 10364
rect 30820 10362 30826 10364
rect 30580 10310 30582 10362
rect 30762 10310 30764 10362
rect 30518 10308 30524 10310
rect 30580 10308 30604 10310
rect 30660 10308 30684 10310
rect 30740 10308 30764 10310
rect 30820 10308 30826 10310
rect 30518 10299 30826 10308
rect 30518 9276 30826 9285
rect 30518 9274 30524 9276
rect 30580 9274 30604 9276
rect 30660 9274 30684 9276
rect 30740 9274 30764 9276
rect 30820 9274 30826 9276
rect 30580 9222 30582 9274
rect 30762 9222 30764 9274
rect 30518 9220 30524 9222
rect 30580 9220 30604 9222
rect 30660 9220 30684 9222
rect 30740 9220 30764 9222
rect 30820 9220 30826 9222
rect 30518 9211 30826 9220
rect 31496 8362 31524 11018
rect 33876 8968 33928 8974
rect 33876 8910 33928 8916
rect 31484 8356 31536 8362
rect 31484 8298 31536 8304
rect 30518 8188 30826 8197
rect 30518 8186 30524 8188
rect 30580 8186 30604 8188
rect 30660 8186 30684 8188
rect 30740 8186 30764 8188
rect 30820 8186 30826 8188
rect 30580 8134 30582 8186
rect 30762 8134 30764 8186
rect 30518 8132 30524 8134
rect 30580 8132 30604 8134
rect 30660 8132 30684 8134
rect 30740 8132 30764 8134
rect 30820 8132 30826 8134
rect 30518 8123 30826 8132
rect 33888 8090 33916 8910
rect 34060 8832 34112 8838
rect 34058 8800 34060 8809
rect 34112 8800 34114 8809
rect 34058 8735 34114 8744
rect 33876 8084 33928 8090
rect 33876 8026 33928 8032
rect 30380 8016 30432 8022
rect 30380 7958 30432 7964
rect 31668 7880 31720 7886
rect 31668 7822 31720 7828
rect 30518 7100 30826 7109
rect 30518 7098 30524 7100
rect 30580 7098 30604 7100
rect 30660 7098 30684 7100
rect 30740 7098 30764 7100
rect 30820 7098 30826 7100
rect 30580 7046 30582 7098
rect 30762 7046 30764 7098
rect 30518 7044 30524 7046
rect 30580 7044 30604 7046
rect 30660 7044 30684 7046
rect 30740 7044 30764 7046
rect 30820 7044 30826 7046
rect 30518 7035 30826 7044
rect 31680 6730 31708 7822
rect 32128 7812 32180 7818
rect 32128 7754 32180 7760
rect 31668 6724 31720 6730
rect 31668 6666 31720 6672
rect 30564 6656 30616 6662
rect 30564 6598 30616 6604
rect 30576 6322 30604 6598
rect 30564 6316 30616 6322
rect 30564 6258 30616 6264
rect 32140 6254 32168 7754
rect 33140 6792 33192 6798
rect 33140 6734 33192 6740
rect 33152 6458 33180 6734
rect 34060 6656 34112 6662
rect 34060 6598 34112 6604
rect 33140 6452 33192 6458
rect 33140 6394 33192 6400
rect 34072 6361 34100 6598
rect 34058 6352 34114 6361
rect 34058 6287 34114 6296
rect 32128 6248 32180 6254
rect 32128 6190 32180 6196
rect 29828 6112 29880 6118
rect 29828 6054 29880 6060
rect 29840 4622 29868 6054
rect 30518 6012 30826 6021
rect 30518 6010 30524 6012
rect 30580 6010 30604 6012
rect 30660 6010 30684 6012
rect 30740 6010 30764 6012
rect 30820 6010 30826 6012
rect 30580 5958 30582 6010
rect 30762 5958 30764 6010
rect 30518 5956 30524 5958
rect 30580 5956 30604 5958
rect 30660 5956 30684 5958
rect 30740 5956 30764 5958
rect 30820 5956 30826 5958
rect 30518 5947 30826 5956
rect 32140 5302 32168 6190
rect 32128 5296 32180 5302
rect 32128 5238 32180 5244
rect 30518 4924 30826 4933
rect 30518 4922 30524 4924
rect 30580 4922 30604 4924
rect 30660 4922 30684 4924
rect 30740 4922 30764 4924
rect 30820 4922 30826 4924
rect 30580 4870 30582 4922
rect 30762 4870 30764 4922
rect 30518 4868 30524 4870
rect 30580 4868 30604 4870
rect 30660 4868 30684 4870
rect 30740 4868 30764 4870
rect 30820 4868 30826 4870
rect 30518 4859 30826 4868
rect 29828 4616 29880 4622
rect 29828 4558 29880 4564
rect 31576 4480 31628 4486
rect 31576 4422 31628 4428
rect 30518 3836 30826 3845
rect 30518 3834 30524 3836
rect 30580 3834 30604 3836
rect 30660 3834 30684 3836
rect 30740 3834 30764 3836
rect 30820 3834 30826 3836
rect 30580 3782 30582 3834
rect 30762 3782 30764 3834
rect 30518 3780 30524 3782
rect 30580 3780 30604 3782
rect 30660 3780 30684 3782
rect 30740 3780 30764 3782
rect 30820 3780 30826 3782
rect 30518 3771 30826 3780
rect 31588 3738 31616 4422
rect 33876 4140 33928 4146
rect 33876 4082 33928 4088
rect 31668 3936 31720 3942
rect 31668 3878 31720 3884
rect 21640 3732 21692 3738
rect 21640 3674 21692 3680
rect 24584 3732 24636 3738
rect 24584 3674 24636 3680
rect 27252 3732 27304 3738
rect 27252 3674 27304 3680
rect 29644 3732 29696 3738
rect 29644 3674 29696 3680
rect 31576 3732 31628 3738
rect 31576 3674 31628 3680
rect 15660 3664 15712 3670
rect 15660 3606 15712 3612
rect 17846 3292 18154 3301
rect 17846 3290 17852 3292
rect 17908 3290 17932 3292
rect 17988 3290 18012 3292
rect 18068 3290 18092 3292
rect 18148 3290 18154 3292
rect 17908 3238 17910 3290
rect 18090 3238 18092 3290
rect 17846 3236 17852 3238
rect 17908 3236 17932 3238
rect 17988 3236 18012 3238
rect 18068 3236 18092 3238
rect 18148 3236 18154 3238
rect 17846 3227 18154 3236
rect 15384 2644 15436 2650
rect 15384 2586 15436 2592
rect 3884 2576 3936 2582
rect 3884 2518 3936 2524
rect 5080 2576 5132 2582
rect 5080 2518 5132 2524
rect 6828 2576 6880 2582
rect 6828 2518 6880 2524
rect 21652 2446 21680 3674
rect 23664 3664 23716 3670
rect 23664 3606 23716 3612
rect 22560 3460 22612 3466
rect 22560 3402 22612 3408
rect 23388 3460 23440 3466
rect 23388 3402 23440 3408
rect 22070 2748 22378 2757
rect 22070 2746 22076 2748
rect 22132 2746 22156 2748
rect 22212 2746 22236 2748
rect 22292 2746 22316 2748
rect 22372 2746 22378 2748
rect 22132 2694 22134 2746
rect 22314 2694 22316 2746
rect 22070 2692 22076 2694
rect 22132 2692 22156 2694
rect 22212 2692 22236 2694
rect 22292 2692 22316 2694
rect 22372 2692 22378 2694
rect 22070 2683 22378 2692
rect 1768 2440 1820 2446
rect 1768 2382 1820 2388
rect 4252 2440 4304 2446
rect 6920 2440 6972 2446
rect 4252 2382 4304 2388
rect 6748 2388 6920 2394
rect 6748 2382 6972 2388
rect 9220 2440 9272 2446
rect 9220 2382 9272 2388
rect 21640 2440 21692 2446
rect 21640 2382 21692 2388
rect 1780 800 1808 2382
rect 4264 800 4292 2382
rect 6748 2366 6960 2382
rect 6748 800 6776 2366
rect 9232 800 9260 2382
rect 22572 2378 22600 3402
rect 23400 2854 23428 3402
rect 23388 2848 23440 2854
rect 23388 2790 23440 2796
rect 23676 2514 23704 3606
rect 23756 3528 23808 3534
rect 23756 3470 23808 3476
rect 23768 3194 23796 3470
rect 24400 3460 24452 3466
rect 24400 3402 24452 3408
rect 23756 3188 23808 3194
rect 23756 3130 23808 3136
rect 24412 3126 24440 3402
rect 24400 3120 24452 3126
rect 24400 3062 24452 3068
rect 24596 3058 24624 3674
rect 26294 3292 26602 3301
rect 26294 3290 26300 3292
rect 26356 3290 26380 3292
rect 26436 3290 26460 3292
rect 26516 3290 26540 3292
rect 26596 3290 26602 3292
rect 26356 3238 26358 3290
rect 26538 3238 26540 3290
rect 26294 3236 26300 3238
rect 26356 3236 26380 3238
rect 26436 3236 26460 3238
rect 26516 3236 26540 3238
rect 26596 3236 26602 3238
rect 26294 3227 26602 3236
rect 24584 3052 24636 3058
rect 24584 2994 24636 3000
rect 23664 2508 23716 2514
rect 23664 2450 23716 2456
rect 29656 2446 29684 3674
rect 30748 3528 30800 3534
rect 30748 3470 30800 3476
rect 30760 3194 30788 3470
rect 30932 3392 30984 3398
rect 30932 3334 30984 3340
rect 30748 3188 30800 3194
rect 30748 3130 30800 3136
rect 30944 3058 30972 3334
rect 30932 3052 30984 3058
rect 30932 2994 30984 3000
rect 30518 2748 30826 2757
rect 30518 2746 30524 2748
rect 30580 2746 30604 2748
rect 30660 2746 30684 2748
rect 30740 2746 30764 2748
rect 30820 2746 30826 2748
rect 30580 2694 30582 2746
rect 30762 2694 30764 2746
rect 30518 2692 30524 2694
rect 30580 2692 30604 2694
rect 30660 2692 30684 2694
rect 30740 2692 30764 2694
rect 30820 2692 30826 2694
rect 30518 2683 30826 2692
rect 31588 2446 31616 3674
rect 31680 3534 31708 3878
rect 33888 3534 33916 4082
rect 34060 3936 34112 3942
rect 34058 3904 34060 3913
rect 34112 3904 34114 3913
rect 34058 3839 34114 3848
rect 31668 3528 31720 3534
rect 31668 3470 31720 3476
rect 33876 3528 33928 3534
rect 33876 3470 33928 3476
rect 33968 2508 34020 2514
rect 33968 2450 34020 2456
rect 29644 2440 29696 2446
rect 29644 2382 29696 2388
rect 31576 2440 31628 2446
rect 31576 2382 31628 2388
rect 22560 2372 22612 2378
rect 22560 2314 22612 2320
rect 14188 2304 14240 2310
rect 14188 2246 14240 2252
rect 21640 2304 21692 2310
rect 21640 2246 21692 2252
rect 29092 2304 29144 2310
rect 29092 2246 29144 2252
rect 9398 2204 9706 2213
rect 9398 2202 9404 2204
rect 9460 2202 9484 2204
rect 9540 2202 9564 2204
rect 9620 2202 9644 2204
rect 9700 2202 9706 2204
rect 9460 2150 9462 2202
rect 9642 2150 9644 2202
rect 9398 2148 9404 2150
rect 9460 2148 9484 2150
rect 9540 2148 9564 2150
rect 9620 2148 9644 2150
rect 9700 2148 9706 2150
rect 9398 2139 9706 2148
rect 14200 800 14228 2246
rect 17846 2204 18154 2213
rect 17846 2202 17852 2204
rect 17908 2202 17932 2204
rect 17988 2202 18012 2204
rect 18068 2202 18092 2204
rect 18148 2202 18154 2204
rect 17908 2150 17910 2202
rect 18090 2150 18092 2202
rect 17846 2148 17852 2150
rect 17908 2148 17932 2150
rect 17988 2148 18012 2150
rect 18068 2148 18092 2150
rect 18148 2148 18154 2150
rect 17846 2139 18154 2148
rect 21652 800 21680 2246
rect 26294 2204 26602 2213
rect 26294 2202 26300 2204
rect 26356 2202 26380 2204
rect 26436 2202 26460 2204
rect 26516 2202 26540 2204
rect 26596 2202 26602 2204
rect 26356 2150 26358 2202
rect 26538 2150 26540 2202
rect 26294 2148 26300 2150
rect 26356 2148 26380 2150
rect 26436 2148 26460 2150
rect 26516 2148 26540 2150
rect 26596 2148 26602 2150
rect 26294 2139 26602 2148
rect 29104 800 29132 2246
rect 33980 1306 34008 2450
rect 34060 2304 34112 2310
rect 34060 2246 34112 2252
rect 34072 1465 34100 2246
rect 34058 1456 34114 1465
rect 34058 1391 34114 1400
rect 33980 1278 34100 1306
rect 34072 800 34100 1278
rect 1766 0 1822 800
rect 4250 0 4306 800
rect 6734 0 6790 800
rect 9218 0 9274 800
rect 11702 0 11758 800
rect 14186 0 14242 800
rect 16670 0 16726 800
rect 19154 0 19210 800
rect 21638 0 21694 800
rect 24122 0 24178 800
rect 26606 0 26662 800
rect 29090 0 29146 800
rect 31574 0 31630 800
rect 34058 0 34114 800
<< via2 >>
rect 1398 17312 1454 17368
rect 9404 17434 9460 17436
rect 9484 17434 9540 17436
rect 9564 17434 9620 17436
rect 9644 17434 9700 17436
rect 9404 17382 9450 17434
rect 9450 17382 9460 17434
rect 9484 17382 9514 17434
rect 9514 17382 9526 17434
rect 9526 17382 9540 17434
rect 9564 17382 9578 17434
rect 9578 17382 9590 17434
rect 9590 17382 9620 17434
rect 9644 17382 9654 17434
rect 9654 17382 9700 17434
rect 9404 17380 9460 17382
rect 9484 17380 9540 17382
rect 9564 17380 9620 17382
rect 9644 17380 9700 17382
rect 17852 17434 17908 17436
rect 17932 17434 17988 17436
rect 18012 17434 18068 17436
rect 18092 17434 18148 17436
rect 17852 17382 17898 17434
rect 17898 17382 17908 17434
rect 17932 17382 17962 17434
rect 17962 17382 17974 17434
rect 17974 17382 17988 17434
rect 18012 17382 18026 17434
rect 18026 17382 18038 17434
rect 18038 17382 18068 17434
rect 18092 17382 18102 17434
rect 18102 17382 18148 17434
rect 17852 17380 17908 17382
rect 17932 17380 17988 17382
rect 18012 17380 18068 17382
rect 18092 17380 18148 17382
rect 26300 17434 26356 17436
rect 26380 17434 26436 17436
rect 26460 17434 26516 17436
rect 26540 17434 26596 17436
rect 26300 17382 26346 17434
rect 26346 17382 26356 17434
rect 26380 17382 26410 17434
rect 26410 17382 26422 17434
rect 26422 17382 26436 17434
rect 26460 17382 26474 17434
rect 26474 17382 26486 17434
rect 26486 17382 26516 17434
rect 26540 17382 26550 17434
rect 26550 17382 26596 17434
rect 26300 17380 26356 17382
rect 26380 17380 26436 17382
rect 26460 17380 26516 17382
rect 26540 17380 26596 17382
rect 34058 18536 34114 18592
rect 5180 16890 5236 16892
rect 5260 16890 5316 16892
rect 5340 16890 5396 16892
rect 5420 16890 5476 16892
rect 5180 16838 5226 16890
rect 5226 16838 5236 16890
rect 5260 16838 5290 16890
rect 5290 16838 5302 16890
rect 5302 16838 5316 16890
rect 5340 16838 5354 16890
rect 5354 16838 5366 16890
rect 5366 16838 5396 16890
rect 5420 16838 5430 16890
rect 5430 16838 5476 16890
rect 5180 16836 5236 16838
rect 5260 16836 5316 16838
rect 5340 16836 5396 16838
rect 5420 16836 5476 16838
rect 5180 15802 5236 15804
rect 5260 15802 5316 15804
rect 5340 15802 5396 15804
rect 5420 15802 5476 15804
rect 5180 15750 5226 15802
rect 5226 15750 5236 15802
rect 5260 15750 5290 15802
rect 5290 15750 5302 15802
rect 5302 15750 5316 15802
rect 5340 15750 5354 15802
rect 5354 15750 5366 15802
rect 5366 15750 5396 15802
rect 5420 15750 5430 15802
rect 5430 15750 5476 15802
rect 5180 15748 5236 15750
rect 5260 15748 5316 15750
rect 5340 15748 5396 15750
rect 5420 15748 5476 15750
rect 5180 14714 5236 14716
rect 5260 14714 5316 14716
rect 5340 14714 5396 14716
rect 5420 14714 5476 14716
rect 5180 14662 5226 14714
rect 5226 14662 5236 14714
rect 5260 14662 5290 14714
rect 5290 14662 5302 14714
rect 5302 14662 5316 14714
rect 5340 14662 5354 14714
rect 5354 14662 5366 14714
rect 5366 14662 5396 14714
rect 5420 14662 5430 14714
rect 5430 14662 5476 14714
rect 5180 14660 5236 14662
rect 5260 14660 5316 14662
rect 5340 14660 5396 14662
rect 5420 14660 5476 14662
rect 5180 13626 5236 13628
rect 5260 13626 5316 13628
rect 5340 13626 5396 13628
rect 5420 13626 5476 13628
rect 5180 13574 5226 13626
rect 5226 13574 5236 13626
rect 5260 13574 5290 13626
rect 5290 13574 5302 13626
rect 5302 13574 5316 13626
rect 5340 13574 5354 13626
rect 5354 13574 5366 13626
rect 5366 13574 5396 13626
rect 5420 13574 5430 13626
rect 5430 13574 5476 13626
rect 5180 13572 5236 13574
rect 5260 13572 5316 13574
rect 5340 13572 5396 13574
rect 5420 13572 5476 13574
rect 5180 12538 5236 12540
rect 5260 12538 5316 12540
rect 5340 12538 5396 12540
rect 5420 12538 5476 12540
rect 5180 12486 5226 12538
rect 5226 12486 5236 12538
rect 5260 12486 5290 12538
rect 5290 12486 5302 12538
rect 5302 12486 5316 12538
rect 5340 12486 5354 12538
rect 5354 12486 5366 12538
rect 5366 12486 5396 12538
rect 5420 12486 5430 12538
rect 5430 12486 5476 12538
rect 5180 12484 5236 12486
rect 5260 12484 5316 12486
rect 5340 12484 5396 12486
rect 5420 12484 5476 12486
rect 1398 12436 1454 12472
rect 1398 12416 1400 12436
rect 1400 12416 1452 12436
rect 1452 12416 1454 12436
rect 5180 11450 5236 11452
rect 5260 11450 5316 11452
rect 5340 11450 5396 11452
rect 5420 11450 5476 11452
rect 5180 11398 5226 11450
rect 5226 11398 5236 11450
rect 5260 11398 5290 11450
rect 5290 11398 5302 11450
rect 5302 11398 5316 11450
rect 5340 11398 5354 11450
rect 5354 11398 5366 11450
rect 5366 11398 5396 11450
rect 5420 11398 5430 11450
rect 5430 11398 5476 11450
rect 5180 11396 5236 11398
rect 5260 11396 5316 11398
rect 5340 11396 5396 11398
rect 5420 11396 5476 11398
rect 1398 7540 1454 7576
rect 1398 7520 1400 7540
rect 1400 7520 1452 7540
rect 1452 7520 1454 7540
rect 3146 2644 3202 2680
rect 3146 2624 3148 2644
rect 3148 2624 3200 2644
rect 3200 2624 3202 2644
rect 5180 10362 5236 10364
rect 5260 10362 5316 10364
rect 5340 10362 5396 10364
rect 5420 10362 5476 10364
rect 5180 10310 5226 10362
rect 5226 10310 5236 10362
rect 5260 10310 5290 10362
rect 5290 10310 5302 10362
rect 5302 10310 5316 10362
rect 5340 10310 5354 10362
rect 5354 10310 5366 10362
rect 5366 10310 5396 10362
rect 5420 10310 5430 10362
rect 5430 10310 5476 10362
rect 5180 10308 5236 10310
rect 5260 10308 5316 10310
rect 5340 10308 5396 10310
rect 5420 10308 5476 10310
rect 5180 9274 5236 9276
rect 5260 9274 5316 9276
rect 5340 9274 5396 9276
rect 5420 9274 5476 9276
rect 5180 9222 5226 9274
rect 5226 9222 5236 9274
rect 5260 9222 5290 9274
rect 5290 9222 5302 9274
rect 5302 9222 5316 9274
rect 5340 9222 5354 9274
rect 5354 9222 5366 9274
rect 5366 9222 5396 9274
rect 5420 9222 5430 9274
rect 5430 9222 5476 9274
rect 5180 9220 5236 9222
rect 5260 9220 5316 9222
rect 5340 9220 5396 9222
rect 5420 9220 5476 9222
rect 5180 8186 5236 8188
rect 5260 8186 5316 8188
rect 5340 8186 5396 8188
rect 5420 8186 5476 8188
rect 5180 8134 5226 8186
rect 5226 8134 5236 8186
rect 5260 8134 5290 8186
rect 5290 8134 5302 8186
rect 5302 8134 5316 8186
rect 5340 8134 5354 8186
rect 5354 8134 5366 8186
rect 5366 8134 5396 8186
rect 5420 8134 5430 8186
rect 5430 8134 5476 8186
rect 5180 8132 5236 8134
rect 5260 8132 5316 8134
rect 5340 8132 5396 8134
rect 5420 8132 5476 8134
rect 5180 7098 5236 7100
rect 5260 7098 5316 7100
rect 5340 7098 5396 7100
rect 5420 7098 5476 7100
rect 5180 7046 5226 7098
rect 5226 7046 5236 7098
rect 5260 7046 5290 7098
rect 5290 7046 5302 7098
rect 5302 7046 5316 7098
rect 5340 7046 5354 7098
rect 5354 7046 5366 7098
rect 5366 7046 5396 7098
rect 5420 7046 5430 7098
rect 5430 7046 5476 7098
rect 5180 7044 5236 7046
rect 5260 7044 5316 7046
rect 5340 7044 5396 7046
rect 5420 7044 5476 7046
rect 9404 16346 9460 16348
rect 9484 16346 9540 16348
rect 9564 16346 9620 16348
rect 9644 16346 9700 16348
rect 9404 16294 9450 16346
rect 9450 16294 9460 16346
rect 9484 16294 9514 16346
rect 9514 16294 9526 16346
rect 9526 16294 9540 16346
rect 9564 16294 9578 16346
rect 9578 16294 9590 16346
rect 9590 16294 9620 16346
rect 9644 16294 9654 16346
rect 9654 16294 9700 16346
rect 9404 16292 9460 16294
rect 9484 16292 9540 16294
rect 9564 16292 9620 16294
rect 9644 16292 9700 16294
rect 13628 16890 13684 16892
rect 13708 16890 13764 16892
rect 13788 16890 13844 16892
rect 13868 16890 13924 16892
rect 13628 16838 13674 16890
rect 13674 16838 13684 16890
rect 13708 16838 13738 16890
rect 13738 16838 13750 16890
rect 13750 16838 13764 16890
rect 13788 16838 13802 16890
rect 13802 16838 13814 16890
rect 13814 16838 13844 16890
rect 13868 16838 13878 16890
rect 13878 16838 13924 16890
rect 13628 16836 13684 16838
rect 13708 16836 13764 16838
rect 13788 16836 13844 16838
rect 13868 16836 13924 16838
rect 17852 16346 17908 16348
rect 17932 16346 17988 16348
rect 18012 16346 18068 16348
rect 18092 16346 18148 16348
rect 17852 16294 17898 16346
rect 17898 16294 17908 16346
rect 17932 16294 17962 16346
rect 17962 16294 17974 16346
rect 17974 16294 17988 16346
rect 18012 16294 18026 16346
rect 18026 16294 18038 16346
rect 18038 16294 18068 16346
rect 18092 16294 18102 16346
rect 18102 16294 18148 16346
rect 17852 16292 17908 16294
rect 17932 16292 17988 16294
rect 18012 16292 18068 16294
rect 18092 16292 18148 16294
rect 13628 15802 13684 15804
rect 13708 15802 13764 15804
rect 13788 15802 13844 15804
rect 13868 15802 13924 15804
rect 13628 15750 13674 15802
rect 13674 15750 13684 15802
rect 13708 15750 13738 15802
rect 13738 15750 13750 15802
rect 13750 15750 13764 15802
rect 13788 15750 13802 15802
rect 13802 15750 13814 15802
rect 13814 15750 13844 15802
rect 13868 15750 13878 15802
rect 13878 15750 13924 15802
rect 13628 15748 13684 15750
rect 13708 15748 13764 15750
rect 13788 15748 13844 15750
rect 13868 15748 13924 15750
rect 9404 15258 9460 15260
rect 9484 15258 9540 15260
rect 9564 15258 9620 15260
rect 9644 15258 9700 15260
rect 9404 15206 9450 15258
rect 9450 15206 9460 15258
rect 9484 15206 9514 15258
rect 9514 15206 9526 15258
rect 9526 15206 9540 15258
rect 9564 15206 9578 15258
rect 9578 15206 9590 15258
rect 9590 15206 9620 15258
rect 9644 15206 9654 15258
rect 9654 15206 9700 15258
rect 9404 15204 9460 15206
rect 9484 15204 9540 15206
rect 9564 15204 9620 15206
rect 9644 15204 9700 15206
rect 9404 14170 9460 14172
rect 9484 14170 9540 14172
rect 9564 14170 9620 14172
rect 9644 14170 9700 14172
rect 9404 14118 9450 14170
rect 9450 14118 9460 14170
rect 9484 14118 9514 14170
rect 9514 14118 9526 14170
rect 9526 14118 9540 14170
rect 9564 14118 9578 14170
rect 9578 14118 9590 14170
rect 9590 14118 9620 14170
rect 9644 14118 9654 14170
rect 9654 14118 9700 14170
rect 9404 14116 9460 14118
rect 9484 14116 9540 14118
rect 9564 14116 9620 14118
rect 9644 14116 9700 14118
rect 9404 13082 9460 13084
rect 9484 13082 9540 13084
rect 9564 13082 9620 13084
rect 9644 13082 9700 13084
rect 9404 13030 9450 13082
rect 9450 13030 9460 13082
rect 9484 13030 9514 13082
rect 9514 13030 9526 13082
rect 9526 13030 9540 13082
rect 9564 13030 9578 13082
rect 9578 13030 9590 13082
rect 9590 13030 9620 13082
rect 9644 13030 9654 13082
rect 9654 13030 9700 13082
rect 9404 13028 9460 13030
rect 9484 13028 9540 13030
rect 9564 13028 9620 13030
rect 9644 13028 9700 13030
rect 17852 15258 17908 15260
rect 17932 15258 17988 15260
rect 18012 15258 18068 15260
rect 18092 15258 18148 15260
rect 17852 15206 17898 15258
rect 17898 15206 17908 15258
rect 17932 15206 17962 15258
rect 17962 15206 17974 15258
rect 17974 15206 17988 15258
rect 18012 15206 18026 15258
rect 18026 15206 18038 15258
rect 18038 15206 18068 15258
rect 18092 15206 18102 15258
rect 18102 15206 18148 15258
rect 17852 15204 17908 15206
rect 17932 15204 17988 15206
rect 18012 15204 18068 15206
rect 18092 15204 18148 15206
rect 13628 14714 13684 14716
rect 13708 14714 13764 14716
rect 13788 14714 13844 14716
rect 13868 14714 13924 14716
rect 13628 14662 13674 14714
rect 13674 14662 13684 14714
rect 13708 14662 13738 14714
rect 13738 14662 13750 14714
rect 13750 14662 13764 14714
rect 13788 14662 13802 14714
rect 13802 14662 13814 14714
rect 13814 14662 13844 14714
rect 13868 14662 13878 14714
rect 13878 14662 13924 14714
rect 13628 14660 13684 14662
rect 13708 14660 13764 14662
rect 13788 14660 13844 14662
rect 13868 14660 13924 14662
rect 13628 13626 13684 13628
rect 13708 13626 13764 13628
rect 13788 13626 13844 13628
rect 13868 13626 13924 13628
rect 13628 13574 13674 13626
rect 13674 13574 13684 13626
rect 13708 13574 13738 13626
rect 13738 13574 13750 13626
rect 13750 13574 13764 13626
rect 13788 13574 13802 13626
rect 13802 13574 13814 13626
rect 13814 13574 13844 13626
rect 13868 13574 13878 13626
rect 13878 13574 13924 13626
rect 13628 13572 13684 13574
rect 13708 13572 13764 13574
rect 13788 13572 13844 13574
rect 13868 13572 13924 13574
rect 17852 14170 17908 14172
rect 17932 14170 17988 14172
rect 18012 14170 18068 14172
rect 18092 14170 18148 14172
rect 17852 14118 17898 14170
rect 17898 14118 17908 14170
rect 17932 14118 17962 14170
rect 17962 14118 17974 14170
rect 17974 14118 17988 14170
rect 18012 14118 18026 14170
rect 18026 14118 18038 14170
rect 18038 14118 18068 14170
rect 18092 14118 18102 14170
rect 18102 14118 18148 14170
rect 17852 14116 17908 14118
rect 17932 14116 17988 14118
rect 18012 14116 18068 14118
rect 18092 14116 18148 14118
rect 22076 16890 22132 16892
rect 22156 16890 22212 16892
rect 22236 16890 22292 16892
rect 22316 16890 22372 16892
rect 22076 16838 22122 16890
rect 22122 16838 22132 16890
rect 22156 16838 22186 16890
rect 22186 16838 22198 16890
rect 22198 16838 22212 16890
rect 22236 16838 22250 16890
rect 22250 16838 22262 16890
rect 22262 16838 22292 16890
rect 22316 16838 22326 16890
rect 22326 16838 22372 16890
rect 22076 16836 22132 16838
rect 22156 16836 22212 16838
rect 22236 16836 22292 16838
rect 22316 16836 22372 16838
rect 26300 16346 26356 16348
rect 26380 16346 26436 16348
rect 26460 16346 26516 16348
rect 26540 16346 26596 16348
rect 26300 16294 26346 16346
rect 26346 16294 26356 16346
rect 26380 16294 26410 16346
rect 26410 16294 26422 16346
rect 26422 16294 26436 16346
rect 26460 16294 26474 16346
rect 26474 16294 26486 16346
rect 26486 16294 26516 16346
rect 26540 16294 26550 16346
rect 26550 16294 26596 16346
rect 26300 16292 26356 16294
rect 26380 16292 26436 16294
rect 26460 16292 26516 16294
rect 26540 16292 26596 16294
rect 30524 16890 30580 16892
rect 30604 16890 30660 16892
rect 30684 16890 30740 16892
rect 30764 16890 30820 16892
rect 30524 16838 30570 16890
rect 30570 16838 30580 16890
rect 30604 16838 30634 16890
rect 30634 16838 30646 16890
rect 30646 16838 30660 16890
rect 30684 16838 30698 16890
rect 30698 16838 30710 16890
rect 30710 16838 30740 16890
rect 30764 16838 30774 16890
rect 30774 16838 30820 16890
rect 30524 16836 30580 16838
rect 30604 16836 30660 16838
rect 30684 16836 30740 16838
rect 30764 16836 30820 16838
rect 9404 11994 9460 11996
rect 9484 11994 9540 11996
rect 9564 11994 9620 11996
rect 9644 11994 9700 11996
rect 9404 11942 9450 11994
rect 9450 11942 9460 11994
rect 9484 11942 9514 11994
rect 9514 11942 9526 11994
rect 9526 11942 9540 11994
rect 9564 11942 9578 11994
rect 9578 11942 9590 11994
rect 9590 11942 9620 11994
rect 9644 11942 9654 11994
rect 9654 11942 9700 11994
rect 9404 11940 9460 11942
rect 9484 11940 9540 11942
rect 9564 11940 9620 11942
rect 9644 11940 9700 11942
rect 17852 13082 17908 13084
rect 17932 13082 17988 13084
rect 18012 13082 18068 13084
rect 18092 13082 18148 13084
rect 17852 13030 17898 13082
rect 17898 13030 17908 13082
rect 17932 13030 17962 13082
rect 17962 13030 17974 13082
rect 17974 13030 17988 13082
rect 18012 13030 18026 13082
rect 18026 13030 18038 13082
rect 18038 13030 18068 13082
rect 18092 13030 18102 13082
rect 18102 13030 18148 13082
rect 17852 13028 17908 13030
rect 17932 13028 17988 13030
rect 18012 13028 18068 13030
rect 18092 13028 18148 13030
rect 13628 12538 13684 12540
rect 13708 12538 13764 12540
rect 13788 12538 13844 12540
rect 13868 12538 13924 12540
rect 13628 12486 13674 12538
rect 13674 12486 13684 12538
rect 13708 12486 13738 12538
rect 13738 12486 13750 12538
rect 13750 12486 13764 12538
rect 13788 12486 13802 12538
rect 13802 12486 13814 12538
rect 13814 12486 13844 12538
rect 13868 12486 13878 12538
rect 13878 12486 13924 12538
rect 13628 12484 13684 12486
rect 13708 12484 13764 12486
rect 13788 12484 13844 12486
rect 13868 12484 13924 12486
rect 17852 11994 17908 11996
rect 17932 11994 17988 11996
rect 18012 11994 18068 11996
rect 18092 11994 18148 11996
rect 17852 11942 17898 11994
rect 17898 11942 17908 11994
rect 17932 11942 17962 11994
rect 17962 11942 17974 11994
rect 17974 11942 17988 11994
rect 18012 11942 18026 11994
rect 18026 11942 18038 11994
rect 18038 11942 18068 11994
rect 18092 11942 18102 11994
rect 18102 11942 18148 11994
rect 17852 11940 17908 11942
rect 17932 11940 17988 11942
rect 18012 11940 18068 11942
rect 18092 11940 18148 11942
rect 13628 11450 13684 11452
rect 13708 11450 13764 11452
rect 13788 11450 13844 11452
rect 13868 11450 13924 11452
rect 13628 11398 13674 11450
rect 13674 11398 13684 11450
rect 13708 11398 13738 11450
rect 13738 11398 13750 11450
rect 13750 11398 13764 11450
rect 13788 11398 13802 11450
rect 13802 11398 13814 11450
rect 13814 11398 13844 11450
rect 13868 11398 13878 11450
rect 13878 11398 13924 11450
rect 13628 11396 13684 11398
rect 13708 11396 13764 11398
rect 13788 11396 13844 11398
rect 13868 11396 13924 11398
rect 9404 10906 9460 10908
rect 9484 10906 9540 10908
rect 9564 10906 9620 10908
rect 9644 10906 9700 10908
rect 9404 10854 9450 10906
rect 9450 10854 9460 10906
rect 9484 10854 9514 10906
rect 9514 10854 9526 10906
rect 9526 10854 9540 10906
rect 9564 10854 9578 10906
rect 9578 10854 9590 10906
rect 9590 10854 9620 10906
rect 9644 10854 9654 10906
rect 9654 10854 9700 10906
rect 9404 10852 9460 10854
rect 9484 10852 9540 10854
rect 9564 10852 9620 10854
rect 9644 10852 9700 10854
rect 9404 9818 9460 9820
rect 9484 9818 9540 9820
rect 9564 9818 9620 9820
rect 9644 9818 9700 9820
rect 9404 9766 9450 9818
rect 9450 9766 9460 9818
rect 9484 9766 9514 9818
rect 9514 9766 9526 9818
rect 9526 9766 9540 9818
rect 9564 9766 9578 9818
rect 9578 9766 9590 9818
rect 9590 9766 9620 9818
rect 9644 9766 9654 9818
rect 9654 9766 9700 9818
rect 9404 9764 9460 9766
rect 9484 9764 9540 9766
rect 9564 9764 9620 9766
rect 9644 9764 9700 9766
rect 9404 8730 9460 8732
rect 9484 8730 9540 8732
rect 9564 8730 9620 8732
rect 9644 8730 9700 8732
rect 9404 8678 9450 8730
rect 9450 8678 9460 8730
rect 9484 8678 9514 8730
rect 9514 8678 9526 8730
rect 9526 8678 9540 8730
rect 9564 8678 9578 8730
rect 9578 8678 9590 8730
rect 9590 8678 9620 8730
rect 9644 8678 9654 8730
rect 9654 8678 9700 8730
rect 9404 8676 9460 8678
rect 9484 8676 9540 8678
rect 9564 8676 9620 8678
rect 9644 8676 9700 8678
rect 9404 7642 9460 7644
rect 9484 7642 9540 7644
rect 9564 7642 9620 7644
rect 9644 7642 9700 7644
rect 9404 7590 9450 7642
rect 9450 7590 9460 7642
rect 9484 7590 9514 7642
rect 9514 7590 9526 7642
rect 9526 7590 9540 7642
rect 9564 7590 9578 7642
rect 9578 7590 9590 7642
rect 9590 7590 9620 7642
rect 9644 7590 9654 7642
rect 9654 7590 9700 7642
rect 9404 7588 9460 7590
rect 9484 7588 9540 7590
rect 9564 7588 9620 7590
rect 9644 7588 9700 7590
rect 5180 6010 5236 6012
rect 5260 6010 5316 6012
rect 5340 6010 5396 6012
rect 5420 6010 5476 6012
rect 5180 5958 5226 6010
rect 5226 5958 5236 6010
rect 5260 5958 5290 6010
rect 5290 5958 5302 6010
rect 5302 5958 5316 6010
rect 5340 5958 5354 6010
rect 5354 5958 5366 6010
rect 5366 5958 5396 6010
rect 5420 5958 5430 6010
rect 5430 5958 5476 6010
rect 5180 5956 5236 5958
rect 5260 5956 5316 5958
rect 5340 5956 5396 5958
rect 5420 5956 5476 5958
rect 5180 4922 5236 4924
rect 5260 4922 5316 4924
rect 5340 4922 5396 4924
rect 5420 4922 5476 4924
rect 5180 4870 5226 4922
rect 5226 4870 5236 4922
rect 5260 4870 5290 4922
rect 5290 4870 5302 4922
rect 5302 4870 5316 4922
rect 5340 4870 5354 4922
rect 5354 4870 5366 4922
rect 5366 4870 5396 4922
rect 5420 4870 5430 4922
rect 5430 4870 5476 4922
rect 5180 4868 5236 4870
rect 5260 4868 5316 4870
rect 5340 4868 5396 4870
rect 5420 4868 5476 4870
rect 9404 6554 9460 6556
rect 9484 6554 9540 6556
rect 9564 6554 9620 6556
rect 9644 6554 9700 6556
rect 9404 6502 9450 6554
rect 9450 6502 9460 6554
rect 9484 6502 9514 6554
rect 9514 6502 9526 6554
rect 9526 6502 9540 6554
rect 9564 6502 9578 6554
rect 9578 6502 9590 6554
rect 9590 6502 9620 6554
rect 9644 6502 9654 6554
rect 9654 6502 9700 6554
rect 9404 6500 9460 6502
rect 9484 6500 9540 6502
rect 9564 6500 9620 6502
rect 9644 6500 9700 6502
rect 13628 10362 13684 10364
rect 13708 10362 13764 10364
rect 13788 10362 13844 10364
rect 13868 10362 13924 10364
rect 13628 10310 13674 10362
rect 13674 10310 13684 10362
rect 13708 10310 13738 10362
rect 13738 10310 13750 10362
rect 13750 10310 13764 10362
rect 13788 10310 13802 10362
rect 13802 10310 13814 10362
rect 13814 10310 13844 10362
rect 13868 10310 13878 10362
rect 13878 10310 13924 10362
rect 13628 10308 13684 10310
rect 13708 10308 13764 10310
rect 13788 10308 13844 10310
rect 13868 10308 13924 10310
rect 13628 9274 13684 9276
rect 13708 9274 13764 9276
rect 13788 9274 13844 9276
rect 13868 9274 13924 9276
rect 13628 9222 13674 9274
rect 13674 9222 13684 9274
rect 13708 9222 13738 9274
rect 13738 9222 13750 9274
rect 13750 9222 13764 9274
rect 13788 9222 13802 9274
rect 13802 9222 13814 9274
rect 13814 9222 13844 9274
rect 13868 9222 13878 9274
rect 13878 9222 13924 9274
rect 13628 9220 13684 9222
rect 13708 9220 13764 9222
rect 13788 9220 13844 9222
rect 13868 9220 13924 9222
rect 9404 5466 9460 5468
rect 9484 5466 9540 5468
rect 9564 5466 9620 5468
rect 9644 5466 9700 5468
rect 9404 5414 9450 5466
rect 9450 5414 9460 5466
rect 9484 5414 9514 5466
rect 9514 5414 9526 5466
rect 9526 5414 9540 5466
rect 9564 5414 9578 5466
rect 9578 5414 9590 5466
rect 9590 5414 9620 5466
rect 9644 5414 9654 5466
rect 9654 5414 9700 5466
rect 9404 5412 9460 5414
rect 9484 5412 9540 5414
rect 9564 5412 9620 5414
rect 9644 5412 9700 5414
rect 9404 4378 9460 4380
rect 9484 4378 9540 4380
rect 9564 4378 9620 4380
rect 9644 4378 9700 4380
rect 9404 4326 9450 4378
rect 9450 4326 9460 4378
rect 9484 4326 9514 4378
rect 9514 4326 9526 4378
rect 9526 4326 9540 4378
rect 9564 4326 9578 4378
rect 9578 4326 9590 4378
rect 9590 4326 9620 4378
rect 9644 4326 9654 4378
rect 9654 4326 9700 4378
rect 9404 4324 9460 4326
rect 9484 4324 9540 4326
rect 9564 4324 9620 4326
rect 9644 4324 9700 4326
rect 5180 3834 5236 3836
rect 5260 3834 5316 3836
rect 5340 3834 5396 3836
rect 5420 3834 5476 3836
rect 5180 3782 5226 3834
rect 5226 3782 5236 3834
rect 5260 3782 5290 3834
rect 5290 3782 5302 3834
rect 5302 3782 5316 3834
rect 5340 3782 5354 3834
rect 5354 3782 5366 3834
rect 5366 3782 5396 3834
rect 5420 3782 5430 3834
rect 5430 3782 5476 3834
rect 5180 3780 5236 3782
rect 5260 3780 5316 3782
rect 5340 3780 5396 3782
rect 5420 3780 5476 3782
rect 5180 2746 5236 2748
rect 5260 2746 5316 2748
rect 5340 2746 5396 2748
rect 5420 2746 5476 2748
rect 5180 2694 5226 2746
rect 5226 2694 5236 2746
rect 5260 2694 5290 2746
rect 5290 2694 5302 2746
rect 5302 2694 5316 2746
rect 5340 2694 5354 2746
rect 5354 2694 5366 2746
rect 5366 2694 5396 2746
rect 5420 2694 5430 2746
rect 5430 2694 5476 2746
rect 5180 2692 5236 2694
rect 5260 2692 5316 2694
rect 5340 2692 5396 2694
rect 5420 2692 5476 2694
rect 9404 3290 9460 3292
rect 9484 3290 9540 3292
rect 9564 3290 9620 3292
rect 9644 3290 9700 3292
rect 9404 3238 9450 3290
rect 9450 3238 9460 3290
rect 9484 3238 9514 3290
rect 9514 3238 9526 3290
rect 9526 3238 9540 3290
rect 9564 3238 9578 3290
rect 9578 3238 9590 3290
rect 9590 3238 9620 3290
rect 9644 3238 9654 3290
rect 9654 3238 9700 3290
rect 9404 3236 9460 3238
rect 9484 3236 9540 3238
rect 9564 3236 9620 3238
rect 9644 3236 9700 3238
rect 17852 10906 17908 10908
rect 17932 10906 17988 10908
rect 18012 10906 18068 10908
rect 18092 10906 18148 10908
rect 17852 10854 17898 10906
rect 17898 10854 17908 10906
rect 17932 10854 17962 10906
rect 17962 10854 17974 10906
rect 17974 10854 17988 10906
rect 18012 10854 18026 10906
rect 18026 10854 18038 10906
rect 18038 10854 18068 10906
rect 18092 10854 18102 10906
rect 18102 10854 18148 10906
rect 17852 10852 17908 10854
rect 17932 10852 17988 10854
rect 18012 10852 18068 10854
rect 18092 10852 18148 10854
rect 22076 15802 22132 15804
rect 22156 15802 22212 15804
rect 22236 15802 22292 15804
rect 22316 15802 22372 15804
rect 22076 15750 22122 15802
rect 22122 15750 22132 15802
rect 22156 15750 22186 15802
rect 22186 15750 22198 15802
rect 22198 15750 22212 15802
rect 22236 15750 22250 15802
rect 22250 15750 22262 15802
rect 22262 15750 22292 15802
rect 22316 15750 22326 15802
rect 22326 15750 22372 15802
rect 22076 15748 22132 15750
rect 22156 15748 22212 15750
rect 22236 15748 22292 15750
rect 22316 15748 22372 15750
rect 26300 15258 26356 15260
rect 26380 15258 26436 15260
rect 26460 15258 26516 15260
rect 26540 15258 26596 15260
rect 26300 15206 26346 15258
rect 26346 15206 26356 15258
rect 26380 15206 26410 15258
rect 26410 15206 26422 15258
rect 26422 15206 26436 15258
rect 26460 15206 26474 15258
rect 26474 15206 26486 15258
rect 26486 15206 26516 15258
rect 26540 15206 26550 15258
rect 26550 15206 26596 15258
rect 26300 15204 26356 15206
rect 26380 15204 26436 15206
rect 26460 15204 26516 15206
rect 26540 15204 26596 15206
rect 22076 14714 22132 14716
rect 22156 14714 22212 14716
rect 22236 14714 22292 14716
rect 22316 14714 22372 14716
rect 22076 14662 22122 14714
rect 22122 14662 22132 14714
rect 22156 14662 22186 14714
rect 22186 14662 22198 14714
rect 22198 14662 22212 14714
rect 22236 14662 22250 14714
rect 22250 14662 22262 14714
rect 22262 14662 22292 14714
rect 22316 14662 22326 14714
rect 22326 14662 22372 14714
rect 22076 14660 22132 14662
rect 22156 14660 22212 14662
rect 22236 14660 22292 14662
rect 22316 14660 22372 14662
rect 22076 13626 22132 13628
rect 22156 13626 22212 13628
rect 22236 13626 22292 13628
rect 22316 13626 22372 13628
rect 22076 13574 22122 13626
rect 22122 13574 22132 13626
rect 22156 13574 22186 13626
rect 22186 13574 22198 13626
rect 22198 13574 22212 13626
rect 22236 13574 22250 13626
rect 22250 13574 22262 13626
rect 22262 13574 22292 13626
rect 22316 13574 22326 13626
rect 22326 13574 22372 13626
rect 22076 13572 22132 13574
rect 22156 13572 22212 13574
rect 22236 13572 22292 13574
rect 22316 13572 22372 13574
rect 30524 15802 30580 15804
rect 30604 15802 30660 15804
rect 30684 15802 30740 15804
rect 30764 15802 30820 15804
rect 30524 15750 30570 15802
rect 30570 15750 30580 15802
rect 30604 15750 30634 15802
rect 30634 15750 30646 15802
rect 30646 15750 30660 15802
rect 30684 15750 30698 15802
rect 30698 15750 30710 15802
rect 30710 15750 30740 15802
rect 30764 15750 30774 15802
rect 30774 15750 30820 15802
rect 30524 15748 30580 15750
rect 30604 15748 30660 15750
rect 30684 15748 30740 15750
rect 30764 15748 30820 15750
rect 26300 14170 26356 14172
rect 26380 14170 26436 14172
rect 26460 14170 26516 14172
rect 26540 14170 26596 14172
rect 26300 14118 26346 14170
rect 26346 14118 26356 14170
rect 26380 14118 26410 14170
rect 26410 14118 26422 14170
rect 26422 14118 26436 14170
rect 26460 14118 26474 14170
rect 26474 14118 26486 14170
rect 26486 14118 26516 14170
rect 26540 14118 26550 14170
rect 26550 14118 26596 14170
rect 26300 14116 26356 14118
rect 26380 14116 26436 14118
rect 26460 14116 26516 14118
rect 26540 14116 26596 14118
rect 26300 13082 26356 13084
rect 26380 13082 26436 13084
rect 26460 13082 26516 13084
rect 26540 13082 26596 13084
rect 26300 13030 26346 13082
rect 26346 13030 26356 13082
rect 26380 13030 26410 13082
rect 26410 13030 26422 13082
rect 26422 13030 26436 13082
rect 26460 13030 26474 13082
rect 26474 13030 26486 13082
rect 26486 13030 26516 13082
rect 26540 13030 26550 13082
rect 26550 13030 26596 13082
rect 26300 13028 26356 13030
rect 26380 13028 26436 13030
rect 26460 13028 26516 13030
rect 26540 13028 26596 13030
rect 22076 12538 22132 12540
rect 22156 12538 22212 12540
rect 22236 12538 22292 12540
rect 22316 12538 22372 12540
rect 22076 12486 22122 12538
rect 22122 12486 22132 12538
rect 22156 12486 22186 12538
rect 22186 12486 22198 12538
rect 22198 12486 22212 12538
rect 22236 12486 22250 12538
rect 22250 12486 22262 12538
rect 22262 12486 22292 12538
rect 22316 12486 22326 12538
rect 22326 12486 22372 12538
rect 22076 12484 22132 12486
rect 22156 12484 22212 12486
rect 22236 12484 22292 12486
rect 22316 12484 22372 12486
rect 13628 8186 13684 8188
rect 13708 8186 13764 8188
rect 13788 8186 13844 8188
rect 13868 8186 13924 8188
rect 13628 8134 13674 8186
rect 13674 8134 13684 8186
rect 13708 8134 13738 8186
rect 13738 8134 13750 8186
rect 13750 8134 13764 8186
rect 13788 8134 13802 8186
rect 13802 8134 13814 8186
rect 13814 8134 13844 8186
rect 13868 8134 13878 8186
rect 13878 8134 13924 8186
rect 13628 8132 13684 8134
rect 13708 8132 13764 8134
rect 13788 8132 13844 8134
rect 13868 8132 13924 8134
rect 13628 7098 13684 7100
rect 13708 7098 13764 7100
rect 13788 7098 13844 7100
rect 13868 7098 13924 7100
rect 13628 7046 13674 7098
rect 13674 7046 13684 7098
rect 13708 7046 13738 7098
rect 13738 7046 13750 7098
rect 13750 7046 13764 7098
rect 13788 7046 13802 7098
rect 13802 7046 13814 7098
rect 13814 7046 13844 7098
rect 13868 7046 13878 7098
rect 13878 7046 13924 7098
rect 13628 7044 13684 7046
rect 13708 7044 13764 7046
rect 13788 7044 13844 7046
rect 13868 7044 13924 7046
rect 13628 6010 13684 6012
rect 13708 6010 13764 6012
rect 13788 6010 13844 6012
rect 13868 6010 13924 6012
rect 13628 5958 13674 6010
rect 13674 5958 13684 6010
rect 13708 5958 13738 6010
rect 13738 5958 13750 6010
rect 13750 5958 13764 6010
rect 13788 5958 13802 6010
rect 13802 5958 13814 6010
rect 13814 5958 13844 6010
rect 13868 5958 13878 6010
rect 13878 5958 13924 6010
rect 13628 5956 13684 5958
rect 13708 5956 13764 5958
rect 13788 5956 13844 5958
rect 13868 5956 13924 5958
rect 13628 4922 13684 4924
rect 13708 4922 13764 4924
rect 13788 4922 13844 4924
rect 13868 4922 13924 4924
rect 13628 4870 13674 4922
rect 13674 4870 13684 4922
rect 13708 4870 13738 4922
rect 13738 4870 13750 4922
rect 13750 4870 13764 4922
rect 13788 4870 13802 4922
rect 13802 4870 13814 4922
rect 13814 4870 13844 4922
rect 13868 4870 13878 4922
rect 13878 4870 13924 4922
rect 13628 4868 13684 4870
rect 13708 4868 13764 4870
rect 13788 4868 13844 4870
rect 13868 4868 13924 4870
rect 13628 3834 13684 3836
rect 13708 3834 13764 3836
rect 13788 3834 13844 3836
rect 13868 3834 13924 3836
rect 13628 3782 13674 3834
rect 13674 3782 13684 3834
rect 13708 3782 13738 3834
rect 13738 3782 13750 3834
rect 13750 3782 13764 3834
rect 13788 3782 13802 3834
rect 13802 3782 13814 3834
rect 13814 3782 13844 3834
rect 13868 3782 13878 3834
rect 13878 3782 13924 3834
rect 13628 3780 13684 3782
rect 13708 3780 13764 3782
rect 13788 3780 13844 3782
rect 13868 3780 13924 3782
rect 13628 2746 13684 2748
rect 13708 2746 13764 2748
rect 13788 2746 13844 2748
rect 13868 2746 13924 2748
rect 13628 2694 13674 2746
rect 13674 2694 13684 2746
rect 13708 2694 13738 2746
rect 13738 2694 13750 2746
rect 13750 2694 13764 2746
rect 13788 2694 13802 2746
rect 13802 2694 13814 2746
rect 13814 2694 13844 2746
rect 13868 2694 13878 2746
rect 13878 2694 13924 2746
rect 13628 2692 13684 2694
rect 13708 2692 13764 2694
rect 13788 2692 13844 2694
rect 13868 2692 13924 2694
rect 17852 9818 17908 9820
rect 17932 9818 17988 9820
rect 18012 9818 18068 9820
rect 18092 9818 18148 9820
rect 17852 9766 17898 9818
rect 17898 9766 17908 9818
rect 17932 9766 17962 9818
rect 17962 9766 17974 9818
rect 17974 9766 17988 9818
rect 18012 9766 18026 9818
rect 18026 9766 18038 9818
rect 18038 9766 18068 9818
rect 18092 9766 18102 9818
rect 18102 9766 18148 9818
rect 17852 9764 17908 9766
rect 17932 9764 17988 9766
rect 18012 9764 18068 9766
rect 18092 9764 18148 9766
rect 17852 8730 17908 8732
rect 17932 8730 17988 8732
rect 18012 8730 18068 8732
rect 18092 8730 18148 8732
rect 17852 8678 17898 8730
rect 17898 8678 17908 8730
rect 17932 8678 17962 8730
rect 17962 8678 17974 8730
rect 17974 8678 17988 8730
rect 18012 8678 18026 8730
rect 18026 8678 18038 8730
rect 18038 8678 18068 8730
rect 18092 8678 18102 8730
rect 18102 8678 18148 8730
rect 17852 8676 17908 8678
rect 17932 8676 17988 8678
rect 18012 8676 18068 8678
rect 18092 8676 18148 8678
rect 17852 7642 17908 7644
rect 17932 7642 17988 7644
rect 18012 7642 18068 7644
rect 18092 7642 18148 7644
rect 17852 7590 17898 7642
rect 17898 7590 17908 7642
rect 17932 7590 17962 7642
rect 17962 7590 17974 7642
rect 17974 7590 17988 7642
rect 18012 7590 18026 7642
rect 18026 7590 18038 7642
rect 18038 7590 18068 7642
rect 18092 7590 18102 7642
rect 18102 7590 18148 7642
rect 17852 7588 17908 7590
rect 17932 7588 17988 7590
rect 18012 7588 18068 7590
rect 18092 7588 18148 7590
rect 17852 6554 17908 6556
rect 17932 6554 17988 6556
rect 18012 6554 18068 6556
rect 18092 6554 18148 6556
rect 17852 6502 17898 6554
rect 17898 6502 17908 6554
rect 17932 6502 17962 6554
rect 17962 6502 17974 6554
rect 17974 6502 17988 6554
rect 18012 6502 18026 6554
rect 18026 6502 18038 6554
rect 18038 6502 18068 6554
rect 18092 6502 18102 6554
rect 18102 6502 18148 6554
rect 17852 6500 17908 6502
rect 17932 6500 17988 6502
rect 18012 6500 18068 6502
rect 18092 6500 18148 6502
rect 17852 5466 17908 5468
rect 17932 5466 17988 5468
rect 18012 5466 18068 5468
rect 18092 5466 18148 5468
rect 17852 5414 17898 5466
rect 17898 5414 17908 5466
rect 17932 5414 17962 5466
rect 17962 5414 17974 5466
rect 17974 5414 17988 5466
rect 18012 5414 18026 5466
rect 18026 5414 18038 5466
rect 18038 5414 18068 5466
rect 18092 5414 18102 5466
rect 18102 5414 18148 5466
rect 17852 5412 17908 5414
rect 17932 5412 17988 5414
rect 18012 5412 18068 5414
rect 18092 5412 18148 5414
rect 17852 4378 17908 4380
rect 17932 4378 17988 4380
rect 18012 4378 18068 4380
rect 18092 4378 18148 4380
rect 17852 4326 17898 4378
rect 17898 4326 17908 4378
rect 17932 4326 17962 4378
rect 17962 4326 17974 4378
rect 17974 4326 17988 4378
rect 18012 4326 18026 4378
rect 18026 4326 18038 4378
rect 18038 4326 18068 4378
rect 18092 4326 18102 4378
rect 18102 4326 18148 4378
rect 17852 4324 17908 4326
rect 17932 4324 17988 4326
rect 18012 4324 18068 4326
rect 18092 4324 18148 4326
rect 22076 11450 22132 11452
rect 22156 11450 22212 11452
rect 22236 11450 22292 11452
rect 22316 11450 22372 11452
rect 22076 11398 22122 11450
rect 22122 11398 22132 11450
rect 22156 11398 22186 11450
rect 22186 11398 22198 11450
rect 22198 11398 22212 11450
rect 22236 11398 22250 11450
rect 22250 11398 22262 11450
rect 22262 11398 22292 11450
rect 22316 11398 22326 11450
rect 22326 11398 22372 11450
rect 22076 11396 22132 11398
rect 22156 11396 22212 11398
rect 22236 11396 22292 11398
rect 22316 11396 22372 11398
rect 22076 10362 22132 10364
rect 22156 10362 22212 10364
rect 22236 10362 22292 10364
rect 22316 10362 22372 10364
rect 22076 10310 22122 10362
rect 22122 10310 22132 10362
rect 22156 10310 22186 10362
rect 22186 10310 22198 10362
rect 22198 10310 22212 10362
rect 22236 10310 22250 10362
rect 22250 10310 22262 10362
rect 22262 10310 22292 10362
rect 22316 10310 22326 10362
rect 22326 10310 22372 10362
rect 22076 10308 22132 10310
rect 22156 10308 22212 10310
rect 22236 10308 22292 10310
rect 22316 10308 22372 10310
rect 22076 9274 22132 9276
rect 22156 9274 22212 9276
rect 22236 9274 22292 9276
rect 22316 9274 22372 9276
rect 22076 9222 22122 9274
rect 22122 9222 22132 9274
rect 22156 9222 22186 9274
rect 22186 9222 22198 9274
rect 22198 9222 22212 9274
rect 22236 9222 22250 9274
rect 22250 9222 22262 9274
rect 22262 9222 22292 9274
rect 22316 9222 22326 9274
rect 22326 9222 22372 9274
rect 22076 9220 22132 9222
rect 22156 9220 22212 9222
rect 22236 9220 22292 9222
rect 22316 9220 22372 9222
rect 26300 11994 26356 11996
rect 26380 11994 26436 11996
rect 26460 11994 26516 11996
rect 26540 11994 26596 11996
rect 26300 11942 26346 11994
rect 26346 11942 26356 11994
rect 26380 11942 26410 11994
rect 26410 11942 26422 11994
rect 26422 11942 26436 11994
rect 26460 11942 26474 11994
rect 26474 11942 26486 11994
rect 26486 11942 26516 11994
rect 26540 11942 26550 11994
rect 26550 11942 26596 11994
rect 26300 11940 26356 11942
rect 26380 11940 26436 11942
rect 26460 11940 26516 11942
rect 26540 11940 26596 11942
rect 26300 10906 26356 10908
rect 26380 10906 26436 10908
rect 26460 10906 26516 10908
rect 26540 10906 26596 10908
rect 26300 10854 26346 10906
rect 26346 10854 26356 10906
rect 26380 10854 26410 10906
rect 26410 10854 26422 10906
rect 26422 10854 26436 10906
rect 26460 10854 26474 10906
rect 26474 10854 26486 10906
rect 26486 10854 26516 10906
rect 26540 10854 26550 10906
rect 26550 10854 26596 10906
rect 26300 10852 26356 10854
rect 26380 10852 26436 10854
rect 26460 10852 26516 10854
rect 26540 10852 26596 10854
rect 26300 9818 26356 9820
rect 26380 9818 26436 9820
rect 26460 9818 26516 9820
rect 26540 9818 26596 9820
rect 26300 9766 26346 9818
rect 26346 9766 26356 9818
rect 26380 9766 26410 9818
rect 26410 9766 26422 9818
rect 26422 9766 26436 9818
rect 26460 9766 26474 9818
rect 26474 9766 26486 9818
rect 26486 9766 26516 9818
rect 26540 9766 26550 9818
rect 26550 9766 26596 9818
rect 26300 9764 26356 9766
rect 26380 9764 26436 9766
rect 26460 9764 26516 9766
rect 26540 9764 26596 9766
rect 26300 8730 26356 8732
rect 26380 8730 26436 8732
rect 26460 8730 26516 8732
rect 26540 8730 26596 8732
rect 26300 8678 26346 8730
rect 26346 8678 26356 8730
rect 26380 8678 26410 8730
rect 26410 8678 26422 8730
rect 26422 8678 26436 8730
rect 26460 8678 26474 8730
rect 26474 8678 26486 8730
rect 26486 8678 26516 8730
rect 26540 8678 26550 8730
rect 26550 8678 26596 8730
rect 26300 8676 26356 8678
rect 26380 8676 26436 8678
rect 26460 8676 26516 8678
rect 26540 8676 26596 8678
rect 22076 8186 22132 8188
rect 22156 8186 22212 8188
rect 22236 8186 22292 8188
rect 22316 8186 22372 8188
rect 22076 8134 22122 8186
rect 22122 8134 22132 8186
rect 22156 8134 22186 8186
rect 22186 8134 22198 8186
rect 22198 8134 22212 8186
rect 22236 8134 22250 8186
rect 22250 8134 22262 8186
rect 22262 8134 22292 8186
rect 22316 8134 22326 8186
rect 22326 8134 22372 8186
rect 22076 8132 22132 8134
rect 22156 8132 22212 8134
rect 22236 8132 22292 8134
rect 22316 8132 22372 8134
rect 22076 7098 22132 7100
rect 22156 7098 22212 7100
rect 22236 7098 22292 7100
rect 22316 7098 22372 7100
rect 22076 7046 22122 7098
rect 22122 7046 22132 7098
rect 22156 7046 22186 7098
rect 22186 7046 22198 7098
rect 22198 7046 22212 7098
rect 22236 7046 22250 7098
rect 22250 7046 22262 7098
rect 22262 7046 22292 7098
rect 22316 7046 22326 7098
rect 22326 7046 22372 7098
rect 22076 7044 22132 7046
rect 22156 7044 22212 7046
rect 22236 7044 22292 7046
rect 22316 7044 22372 7046
rect 22076 6010 22132 6012
rect 22156 6010 22212 6012
rect 22236 6010 22292 6012
rect 22316 6010 22372 6012
rect 22076 5958 22122 6010
rect 22122 5958 22132 6010
rect 22156 5958 22186 6010
rect 22186 5958 22198 6010
rect 22198 5958 22212 6010
rect 22236 5958 22250 6010
rect 22250 5958 22262 6010
rect 22262 5958 22292 6010
rect 22316 5958 22326 6010
rect 22326 5958 22372 6010
rect 22076 5956 22132 5958
rect 22156 5956 22212 5958
rect 22236 5956 22292 5958
rect 22316 5956 22372 5958
rect 26300 7642 26356 7644
rect 26380 7642 26436 7644
rect 26460 7642 26516 7644
rect 26540 7642 26596 7644
rect 26300 7590 26346 7642
rect 26346 7590 26356 7642
rect 26380 7590 26410 7642
rect 26410 7590 26422 7642
rect 26422 7590 26436 7642
rect 26460 7590 26474 7642
rect 26474 7590 26486 7642
rect 26486 7590 26516 7642
rect 26540 7590 26550 7642
rect 26550 7590 26596 7642
rect 26300 7588 26356 7590
rect 26380 7588 26436 7590
rect 26460 7588 26516 7590
rect 26540 7588 26596 7590
rect 26300 6554 26356 6556
rect 26380 6554 26436 6556
rect 26460 6554 26516 6556
rect 26540 6554 26596 6556
rect 26300 6502 26346 6554
rect 26346 6502 26356 6554
rect 26380 6502 26410 6554
rect 26410 6502 26422 6554
rect 26422 6502 26436 6554
rect 26460 6502 26474 6554
rect 26474 6502 26486 6554
rect 26486 6502 26516 6554
rect 26540 6502 26550 6554
rect 26550 6502 26596 6554
rect 26300 6500 26356 6502
rect 26380 6500 26436 6502
rect 26460 6500 26516 6502
rect 26540 6500 26596 6502
rect 26300 5466 26356 5468
rect 26380 5466 26436 5468
rect 26460 5466 26516 5468
rect 26540 5466 26596 5468
rect 26300 5414 26346 5466
rect 26346 5414 26356 5466
rect 26380 5414 26410 5466
rect 26410 5414 26422 5466
rect 26422 5414 26436 5466
rect 26460 5414 26474 5466
rect 26474 5414 26486 5466
rect 26486 5414 26516 5466
rect 26540 5414 26550 5466
rect 26550 5414 26596 5466
rect 26300 5412 26356 5414
rect 26380 5412 26436 5414
rect 26460 5412 26516 5414
rect 26540 5412 26596 5414
rect 22076 4922 22132 4924
rect 22156 4922 22212 4924
rect 22236 4922 22292 4924
rect 22316 4922 22372 4924
rect 22076 4870 22122 4922
rect 22122 4870 22132 4922
rect 22156 4870 22186 4922
rect 22186 4870 22198 4922
rect 22198 4870 22212 4922
rect 22236 4870 22250 4922
rect 22250 4870 22262 4922
rect 22262 4870 22292 4922
rect 22316 4870 22326 4922
rect 22326 4870 22372 4922
rect 22076 4868 22132 4870
rect 22156 4868 22212 4870
rect 22236 4868 22292 4870
rect 22316 4868 22372 4870
rect 26300 4378 26356 4380
rect 26380 4378 26436 4380
rect 26460 4378 26516 4380
rect 26540 4378 26596 4380
rect 26300 4326 26346 4378
rect 26346 4326 26356 4378
rect 26380 4326 26410 4378
rect 26410 4326 26422 4378
rect 26422 4326 26436 4378
rect 26460 4326 26474 4378
rect 26474 4326 26486 4378
rect 26486 4326 26516 4378
rect 26540 4326 26550 4378
rect 26550 4326 26596 4378
rect 26300 4324 26356 4326
rect 26380 4324 26436 4326
rect 26460 4324 26516 4326
rect 26540 4324 26596 4326
rect 22076 3834 22132 3836
rect 22156 3834 22212 3836
rect 22236 3834 22292 3836
rect 22316 3834 22372 3836
rect 22076 3782 22122 3834
rect 22122 3782 22132 3834
rect 22156 3782 22186 3834
rect 22186 3782 22198 3834
rect 22198 3782 22212 3834
rect 22236 3782 22250 3834
rect 22250 3782 22262 3834
rect 22262 3782 22292 3834
rect 22316 3782 22326 3834
rect 22326 3782 22372 3834
rect 22076 3780 22132 3782
rect 22156 3780 22212 3782
rect 22236 3780 22292 3782
rect 22316 3780 22372 3782
rect 30524 14714 30580 14716
rect 30604 14714 30660 14716
rect 30684 14714 30740 14716
rect 30764 14714 30820 14716
rect 30524 14662 30570 14714
rect 30570 14662 30580 14714
rect 30604 14662 30634 14714
rect 30634 14662 30646 14714
rect 30646 14662 30660 14714
rect 30684 14662 30698 14714
rect 30698 14662 30710 14714
rect 30710 14662 30740 14714
rect 30764 14662 30774 14714
rect 30774 14662 30820 14714
rect 30524 14660 30580 14662
rect 30604 14660 30660 14662
rect 30684 14660 30740 14662
rect 30764 14660 30820 14662
rect 30524 13626 30580 13628
rect 30604 13626 30660 13628
rect 30684 13626 30740 13628
rect 30764 13626 30820 13628
rect 30524 13574 30570 13626
rect 30570 13574 30580 13626
rect 30604 13574 30634 13626
rect 30634 13574 30646 13626
rect 30646 13574 30660 13626
rect 30684 13574 30698 13626
rect 30698 13574 30710 13626
rect 30710 13574 30740 13626
rect 30764 13574 30774 13626
rect 30774 13574 30820 13626
rect 30524 13572 30580 13574
rect 30604 13572 30660 13574
rect 30684 13572 30740 13574
rect 30764 13572 30820 13574
rect 30524 12538 30580 12540
rect 30604 12538 30660 12540
rect 30684 12538 30740 12540
rect 30764 12538 30820 12540
rect 30524 12486 30570 12538
rect 30570 12486 30580 12538
rect 30604 12486 30634 12538
rect 30634 12486 30646 12538
rect 30646 12486 30660 12538
rect 30684 12486 30698 12538
rect 30698 12486 30710 12538
rect 30710 12486 30740 12538
rect 30764 12486 30774 12538
rect 30774 12486 30820 12538
rect 30524 12484 30580 12486
rect 30604 12484 30660 12486
rect 30684 12484 30740 12486
rect 30764 12484 30820 12486
rect 30524 11450 30580 11452
rect 30604 11450 30660 11452
rect 30684 11450 30740 11452
rect 30764 11450 30820 11452
rect 30524 11398 30570 11450
rect 30570 11398 30580 11450
rect 30604 11398 30634 11450
rect 30634 11398 30646 11450
rect 30646 11398 30660 11450
rect 30684 11398 30698 11450
rect 30698 11398 30710 11450
rect 30710 11398 30740 11450
rect 30764 11398 30774 11450
rect 30774 11398 30820 11450
rect 30524 11396 30580 11398
rect 30604 11396 30660 11398
rect 30684 11396 30740 11398
rect 30764 11396 30820 11398
rect 34058 16088 34114 16144
rect 34058 13676 34060 13696
rect 34060 13676 34112 13696
rect 34112 13676 34114 13696
rect 34058 13640 34114 13676
rect 34058 11192 34114 11248
rect 30524 10362 30580 10364
rect 30604 10362 30660 10364
rect 30684 10362 30740 10364
rect 30764 10362 30820 10364
rect 30524 10310 30570 10362
rect 30570 10310 30580 10362
rect 30604 10310 30634 10362
rect 30634 10310 30646 10362
rect 30646 10310 30660 10362
rect 30684 10310 30698 10362
rect 30698 10310 30710 10362
rect 30710 10310 30740 10362
rect 30764 10310 30774 10362
rect 30774 10310 30820 10362
rect 30524 10308 30580 10310
rect 30604 10308 30660 10310
rect 30684 10308 30740 10310
rect 30764 10308 30820 10310
rect 30524 9274 30580 9276
rect 30604 9274 30660 9276
rect 30684 9274 30740 9276
rect 30764 9274 30820 9276
rect 30524 9222 30570 9274
rect 30570 9222 30580 9274
rect 30604 9222 30634 9274
rect 30634 9222 30646 9274
rect 30646 9222 30660 9274
rect 30684 9222 30698 9274
rect 30698 9222 30710 9274
rect 30710 9222 30740 9274
rect 30764 9222 30774 9274
rect 30774 9222 30820 9274
rect 30524 9220 30580 9222
rect 30604 9220 30660 9222
rect 30684 9220 30740 9222
rect 30764 9220 30820 9222
rect 30524 8186 30580 8188
rect 30604 8186 30660 8188
rect 30684 8186 30740 8188
rect 30764 8186 30820 8188
rect 30524 8134 30570 8186
rect 30570 8134 30580 8186
rect 30604 8134 30634 8186
rect 30634 8134 30646 8186
rect 30646 8134 30660 8186
rect 30684 8134 30698 8186
rect 30698 8134 30710 8186
rect 30710 8134 30740 8186
rect 30764 8134 30774 8186
rect 30774 8134 30820 8186
rect 30524 8132 30580 8134
rect 30604 8132 30660 8134
rect 30684 8132 30740 8134
rect 30764 8132 30820 8134
rect 34058 8780 34060 8800
rect 34060 8780 34112 8800
rect 34112 8780 34114 8800
rect 34058 8744 34114 8780
rect 30524 7098 30580 7100
rect 30604 7098 30660 7100
rect 30684 7098 30740 7100
rect 30764 7098 30820 7100
rect 30524 7046 30570 7098
rect 30570 7046 30580 7098
rect 30604 7046 30634 7098
rect 30634 7046 30646 7098
rect 30646 7046 30660 7098
rect 30684 7046 30698 7098
rect 30698 7046 30710 7098
rect 30710 7046 30740 7098
rect 30764 7046 30774 7098
rect 30774 7046 30820 7098
rect 30524 7044 30580 7046
rect 30604 7044 30660 7046
rect 30684 7044 30740 7046
rect 30764 7044 30820 7046
rect 34058 6296 34114 6352
rect 30524 6010 30580 6012
rect 30604 6010 30660 6012
rect 30684 6010 30740 6012
rect 30764 6010 30820 6012
rect 30524 5958 30570 6010
rect 30570 5958 30580 6010
rect 30604 5958 30634 6010
rect 30634 5958 30646 6010
rect 30646 5958 30660 6010
rect 30684 5958 30698 6010
rect 30698 5958 30710 6010
rect 30710 5958 30740 6010
rect 30764 5958 30774 6010
rect 30774 5958 30820 6010
rect 30524 5956 30580 5958
rect 30604 5956 30660 5958
rect 30684 5956 30740 5958
rect 30764 5956 30820 5958
rect 30524 4922 30580 4924
rect 30604 4922 30660 4924
rect 30684 4922 30740 4924
rect 30764 4922 30820 4924
rect 30524 4870 30570 4922
rect 30570 4870 30580 4922
rect 30604 4870 30634 4922
rect 30634 4870 30646 4922
rect 30646 4870 30660 4922
rect 30684 4870 30698 4922
rect 30698 4870 30710 4922
rect 30710 4870 30740 4922
rect 30764 4870 30774 4922
rect 30774 4870 30820 4922
rect 30524 4868 30580 4870
rect 30604 4868 30660 4870
rect 30684 4868 30740 4870
rect 30764 4868 30820 4870
rect 30524 3834 30580 3836
rect 30604 3834 30660 3836
rect 30684 3834 30740 3836
rect 30764 3834 30820 3836
rect 30524 3782 30570 3834
rect 30570 3782 30580 3834
rect 30604 3782 30634 3834
rect 30634 3782 30646 3834
rect 30646 3782 30660 3834
rect 30684 3782 30698 3834
rect 30698 3782 30710 3834
rect 30710 3782 30740 3834
rect 30764 3782 30774 3834
rect 30774 3782 30820 3834
rect 30524 3780 30580 3782
rect 30604 3780 30660 3782
rect 30684 3780 30740 3782
rect 30764 3780 30820 3782
rect 17852 3290 17908 3292
rect 17932 3290 17988 3292
rect 18012 3290 18068 3292
rect 18092 3290 18148 3292
rect 17852 3238 17898 3290
rect 17898 3238 17908 3290
rect 17932 3238 17962 3290
rect 17962 3238 17974 3290
rect 17974 3238 17988 3290
rect 18012 3238 18026 3290
rect 18026 3238 18038 3290
rect 18038 3238 18068 3290
rect 18092 3238 18102 3290
rect 18102 3238 18148 3290
rect 17852 3236 17908 3238
rect 17932 3236 17988 3238
rect 18012 3236 18068 3238
rect 18092 3236 18148 3238
rect 22076 2746 22132 2748
rect 22156 2746 22212 2748
rect 22236 2746 22292 2748
rect 22316 2746 22372 2748
rect 22076 2694 22122 2746
rect 22122 2694 22132 2746
rect 22156 2694 22186 2746
rect 22186 2694 22198 2746
rect 22198 2694 22212 2746
rect 22236 2694 22250 2746
rect 22250 2694 22262 2746
rect 22262 2694 22292 2746
rect 22316 2694 22326 2746
rect 22326 2694 22372 2746
rect 22076 2692 22132 2694
rect 22156 2692 22212 2694
rect 22236 2692 22292 2694
rect 22316 2692 22372 2694
rect 26300 3290 26356 3292
rect 26380 3290 26436 3292
rect 26460 3290 26516 3292
rect 26540 3290 26596 3292
rect 26300 3238 26346 3290
rect 26346 3238 26356 3290
rect 26380 3238 26410 3290
rect 26410 3238 26422 3290
rect 26422 3238 26436 3290
rect 26460 3238 26474 3290
rect 26474 3238 26486 3290
rect 26486 3238 26516 3290
rect 26540 3238 26550 3290
rect 26550 3238 26596 3290
rect 26300 3236 26356 3238
rect 26380 3236 26436 3238
rect 26460 3236 26516 3238
rect 26540 3236 26596 3238
rect 30524 2746 30580 2748
rect 30604 2746 30660 2748
rect 30684 2746 30740 2748
rect 30764 2746 30820 2748
rect 30524 2694 30570 2746
rect 30570 2694 30580 2746
rect 30604 2694 30634 2746
rect 30634 2694 30646 2746
rect 30646 2694 30660 2746
rect 30684 2694 30698 2746
rect 30698 2694 30710 2746
rect 30710 2694 30740 2746
rect 30764 2694 30774 2746
rect 30774 2694 30820 2746
rect 30524 2692 30580 2694
rect 30604 2692 30660 2694
rect 30684 2692 30740 2694
rect 30764 2692 30820 2694
rect 34058 3884 34060 3904
rect 34060 3884 34112 3904
rect 34112 3884 34114 3904
rect 34058 3848 34114 3884
rect 9404 2202 9460 2204
rect 9484 2202 9540 2204
rect 9564 2202 9620 2204
rect 9644 2202 9700 2204
rect 9404 2150 9450 2202
rect 9450 2150 9460 2202
rect 9484 2150 9514 2202
rect 9514 2150 9526 2202
rect 9526 2150 9540 2202
rect 9564 2150 9578 2202
rect 9578 2150 9590 2202
rect 9590 2150 9620 2202
rect 9644 2150 9654 2202
rect 9654 2150 9700 2202
rect 9404 2148 9460 2150
rect 9484 2148 9540 2150
rect 9564 2148 9620 2150
rect 9644 2148 9700 2150
rect 17852 2202 17908 2204
rect 17932 2202 17988 2204
rect 18012 2202 18068 2204
rect 18092 2202 18148 2204
rect 17852 2150 17898 2202
rect 17898 2150 17908 2202
rect 17932 2150 17962 2202
rect 17962 2150 17974 2202
rect 17974 2150 17988 2202
rect 18012 2150 18026 2202
rect 18026 2150 18038 2202
rect 18038 2150 18068 2202
rect 18092 2150 18102 2202
rect 18102 2150 18148 2202
rect 17852 2148 17908 2150
rect 17932 2148 17988 2150
rect 18012 2148 18068 2150
rect 18092 2148 18148 2150
rect 26300 2202 26356 2204
rect 26380 2202 26436 2204
rect 26460 2202 26516 2204
rect 26540 2202 26596 2204
rect 26300 2150 26346 2202
rect 26346 2150 26356 2202
rect 26380 2150 26410 2202
rect 26410 2150 26422 2202
rect 26422 2150 26436 2202
rect 26460 2150 26474 2202
rect 26474 2150 26486 2202
rect 26486 2150 26516 2202
rect 26540 2150 26550 2202
rect 26550 2150 26596 2202
rect 26300 2148 26356 2150
rect 26380 2148 26436 2150
rect 26460 2148 26516 2150
rect 26540 2148 26596 2150
rect 34058 1400 34114 1456
<< metal3 >>
rect 34053 18594 34119 18597
rect 35200 18594 36000 18624
rect 34053 18592 36000 18594
rect 34053 18536 34058 18592
rect 34114 18536 36000 18592
rect 34053 18534 36000 18536
rect 34053 18531 34119 18534
rect 35200 18504 36000 18534
rect 9394 17440 9710 17441
rect 0 17370 800 17400
rect 9394 17376 9400 17440
rect 9464 17376 9480 17440
rect 9544 17376 9560 17440
rect 9624 17376 9640 17440
rect 9704 17376 9710 17440
rect 9394 17375 9710 17376
rect 17842 17440 18158 17441
rect 17842 17376 17848 17440
rect 17912 17376 17928 17440
rect 17992 17376 18008 17440
rect 18072 17376 18088 17440
rect 18152 17376 18158 17440
rect 17842 17375 18158 17376
rect 26290 17440 26606 17441
rect 26290 17376 26296 17440
rect 26360 17376 26376 17440
rect 26440 17376 26456 17440
rect 26520 17376 26536 17440
rect 26600 17376 26606 17440
rect 26290 17375 26606 17376
rect 1393 17370 1459 17373
rect 0 17368 1459 17370
rect 0 17312 1398 17368
rect 1454 17312 1459 17368
rect 0 17310 1459 17312
rect 0 17280 800 17310
rect 1393 17307 1459 17310
rect 5170 16896 5486 16897
rect 5170 16832 5176 16896
rect 5240 16832 5256 16896
rect 5320 16832 5336 16896
rect 5400 16832 5416 16896
rect 5480 16832 5486 16896
rect 5170 16831 5486 16832
rect 13618 16896 13934 16897
rect 13618 16832 13624 16896
rect 13688 16832 13704 16896
rect 13768 16832 13784 16896
rect 13848 16832 13864 16896
rect 13928 16832 13934 16896
rect 13618 16831 13934 16832
rect 22066 16896 22382 16897
rect 22066 16832 22072 16896
rect 22136 16832 22152 16896
rect 22216 16832 22232 16896
rect 22296 16832 22312 16896
rect 22376 16832 22382 16896
rect 22066 16831 22382 16832
rect 30514 16896 30830 16897
rect 30514 16832 30520 16896
rect 30584 16832 30600 16896
rect 30664 16832 30680 16896
rect 30744 16832 30760 16896
rect 30824 16832 30830 16896
rect 30514 16831 30830 16832
rect 9394 16352 9710 16353
rect 9394 16288 9400 16352
rect 9464 16288 9480 16352
rect 9544 16288 9560 16352
rect 9624 16288 9640 16352
rect 9704 16288 9710 16352
rect 9394 16287 9710 16288
rect 17842 16352 18158 16353
rect 17842 16288 17848 16352
rect 17912 16288 17928 16352
rect 17992 16288 18008 16352
rect 18072 16288 18088 16352
rect 18152 16288 18158 16352
rect 17842 16287 18158 16288
rect 26290 16352 26606 16353
rect 26290 16288 26296 16352
rect 26360 16288 26376 16352
rect 26440 16288 26456 16352
rect 26520 16288 26536 16352
rect 26600 16288 26606 16352
rect 26290 16287 26606 16288
rect 34053 16146 34119 16149
rect 35200 16146 36000 16176
rect 34053 16144 36000 16146
rect 34053 16088 34058 16144
rect 34114 16088 36000 16144
rect 34053 16086 36000 16088
rect 34053 16083 34119 16086
rect 35200 16056 36000 16086
rect 5170 15808 5486 15809
rect 5170 15744 5176 15808
rect 5240 15744 5256 15808
rect 5320 15744 5336 15808
rect 5400 15744 5416 15808
rect 5480 15744 5486 15808
rect 5170 15743 5486 15744
rect 13618 15808 13934 15809
rect 13618 15744 13624 15808
rect 13688 15744 13704 15808
rect 13768 15744 13784 15808
rect 13848 15744 13864 15808
rect 13928 15744 13934 15808
rect 13618 15743 13934 15744
rect 22066 15808 22382 15809
rect 22066 15744 22072 15808
rect 22136 15744 22152 15808
rect 22216 15744 22232 15808
rect 22296 15744 22312 15808
rect 22376 15744 22382 15808
rect 22066 15743 22382 15744
rect 30514 15808 30830 15809
rect 30514 15744 30520 15808
rect 30584 15744 30600 15808
rect 30664 15744 30680 15808
rect 30744 15744 30760 15808
rect 30824 15744 30830 15808
rect 30514 15743 30830 15744
rect 9394 15264 9710 15265
rect 9394 15200 9400 15264
rect 9464 15200 9480 15264
rect 9544 15200 9560 15264
rect 9624 15200 9640 15264
rect 9704 15200 9710 15264
rect 9394 15199 9710 15200
rect 17842 15264 18158 15265
rect 17842 15200 17848 15264
rect 17912 15200 17928 15264
rect 17992 15200 18008 15264
rect 18072 15200 18088 15264
rect 18152 15200 18158 15264
rect 17842 15199 18158 15200
rect 26290 15264 26606 15265
rect 26290 15200 26296 15264
rect 26360 15200 26376 15264
rect 26440 15200 26456 15264
rect 26520 15200 26536 15264
rect 26600 15200 26606 15264
rect 26290 15199 26606 15200
rect 5170 14720 5486 14721
rect 5170 14656 5176 14720
rect 5240 14656 5256 14720
rect 5320 14656 5336 14720
rect 5400 14656 5416 14720
rect 5480 14656 5486 14720
rect 5170 14655 5486 14656
rect 13618 14720 13934 14721
rect 13618 14656 13624 14720
rect 13688 14656 13704 14720
rect 13768 14656 13784 14720
rect 13848 14656 13864 14720
rect 13928 14656 13934 14720
rect 13618 14655 13934 14656
rect 22066 14720 22382 14721
rect 22066 14656 22072 14720
rect 22136 14656 22152 14720
rect 22216 14656 22232 14720
rect 22296 14656 22312 14720
rect 22376 14656 22382 14720
rect 22066 14655 22382 14656
rect 30514 14720 30830 14721
rect 30514 14656 30520 14720
rect 30584 14656 30600 14720
rect 30664 14656 30680 14720
rect 30744 14656 30760 14720
rect 30824 14656 30830 14720
rect 30514 14655 30830 14656
rect 9394 14176 9710 14177
rect 9394 14112 9400 14176
rect 9464 14112 9480 14176
rect 9544 14112 9560 14176
rect 9624 14112 9640 14176
rect 9704 14112 9710 14176
rect 9394 14111 9710 14112
rect 17842 14176 18158 14177
rect 17842 14112 17848 14176
rect 17912 14112 17928 14176
rect 17992 14112 18008 14176
rect 18072 14112 18088 14176
rect 18152 14112 18158 14176
rect 17842 14111 18158 14112
rect 26290 14176 26606 14177
rect 26290 14112 26296 14176
rect 26360 14112 26376 14176
rect 26440 14112 26456 14176
rect 26520 14112 26536 14176
rect 26600 14112 26606 14176
rect 26290 14111 26606 14112
rect 34053 13698 34119 13701
rect 35200 13698 36000 13728
rect 34053 13696 36000 13698
rect 34053 13640 34058 13696
rect 34114 13640 36000 13696
rect 34053 13638 36000 13640
rect 34053 13635 34119 13638
rect 5170 13632 5486 13633
rect 5170 13568 5176 13632
rect 5240 13568 5256 13632
rect 5320 13568 5336 13632
rect 5400 13568 5416 13632
rect 5480 13568 5486 13632
rect 5170 13567 5486 13568
rect 13618 13632 13934 13633
rect 13618 13568 13624 13632
rect 13688 13568 13704 13632
rect 13768 13568 13784 13632
rect 13848 13568 13864 13632
rect 13928 13568 13934 13632
rect 13618 13567 13934 13568
rect 22066 13632 22382 13633
rect 22066 13568 22072 13632
rect 22136 13568 22152 13632
rect 22216 13568 22232 13632
rect 22296 13568 22312 13632
rect 22376 13568 22382 13632
rect 22066 13567 22382 13568
rect 30514 13632 30830 13633
rect 30514 13568 30520 13632
rect 30584 13568 30600 13632
rect 30664 13568 30680 13632
rect 30744 13568 30760 13632
rect 30824 13568 30830 13632
rect 35200 13608 36000 13638
rect 30514 13567 30830 13568
rect 9394 13088 9710 13089
rect 9394 13024 9400 13088
rect 9464 13024 9480 13088
rect 9544 13024 9560 13088
rect 9624 13024 9640 13088
rect 9704 13024 9710 13088
rect 9394 13023 9710 13024
rect 17842 13088 18158 13089
rect 17842 13024 17848 13088
rect 17912 13024 17928 13088
rect 17992 13024 18008 13088
rect 18072 13024 18088 13088
rect 18152 13024 18158 13088
rect 17842 13023 18158 13024
rect 26290 13088 26606 13089
rect 26290 13024 26296 13088
rect 26360 13024 26376 13088
rect 26440 13024 26456 13088
rect 26520 13024 26536 13088
rect 26600 13024 26606 13088
rect 26290 13023 26606 13024
rect 5170 12544 5486 12545
rect 0 12474 800 12504
rect 5170 12480 5176 12544
rect 5240 12480 5256 12544
rect 5320 12480 5336 12544
rect 5400 12480 5416 12544
rect 5480 12480 5486 12544
rect 5170 12479 5486 12480
rect 13618 12544 13934 12545
rect 13618 12480 13624 12544
rect 13688 12480 13704 12544
rect 13768 12480 13784 12544
rect 13848 12480 13864 12544
rect 13928 12480 13934 12544
rect 13618 12479 13934 12480
rect 22066 12544 22382 12545
rect 22066 12480 22072 12544
rect 22136 12480 22152 12544
rect 22216 12480 22232 12544
rect 22296 12480 22312 12544
rect 22376 12480 22382 12544
rect 22066 12479 22382 12480
rect 30514 12544 30830 12545
rect 30514 12480 30520 12544
rect 30584 12480 30600 12544
rect 30664 12480 30680 12544
rect 30744 12480 30760 12544
rect 30824 12480 30830 12544
rect 30514 12479 30830 12480
rect 1393 12474 1459 12477
rect 0 12472 1459 12474
rect 0 12416 1398 12472
rect 1454 12416 1459 12472
rect 0 12414 1459 12416
rect 0 12384 800 12414
rect 1393 12411 1459 12414
rect 9394 12000 9710 12001
rect 9394 11936 9400 12000
rect 9464 11936 9480 12000
rect 9544 11936 9560 12000
rect 9624 11936 9640 12000
rect 9704 11936 9710 12000
rect 9394 11935 9710 11936
rect 17842 12000 18158 12001
rect 17842 11936 17848 12000
rect 17912 11936 17928 12000
rect 17992 11936 18008 12000
rect 18072 11936 18088 12000
rect 18152 11936 18158 12000
rect 17842 11935 18158 11936
rect 26290 12000 26606 12001
rect 26290 11936 26296 12000
rect 26360 11936 26376 12000
rect 26440 11936 26456 12000
rect 26520 11936 26536 12000
rect 26600 11936 26606 12000
rect 26290 11935 26606 11936
rect 5170 11456 5486 11457
rect 5170 11392 5176 11456
rect 5240 11392 5256 11456
rect 5320 11392 5336 11456
rect 5400 11392 5416 11456
rect 5480 11392 5486 11456
rect 5170 11391 5486 11392
rect 13618 11456 13934 11457
rect 13618 11392 13624 11456
rect 13688 11392 13704 11456
rect 13768 11392 13784 11456
rect 13848 11392 13864 11456
rect 13928 11392 13934 11456
rect 13618 11391 13934 11392
rect 22066 11456 22382 11457
rect 22066 11392 22072 11456
rect 22136 11392 22152 11456
rect 22216 11392 22232 11456
rect 22296 11392 22312 11456
rect 22376 11392 22382 11456
rect 22066 11391 22382 11392
rect 30514 11456 30830 11457
rect 30514 11392 30520 11456
rect 30584 11392 30600 11456
rect 30664 11392 30680 11456
rect 30744 11392 30760 11456
rect 30824 11392 30830 11456
rect 30514 11391 30830 11392
rect 34053 11250 34119 11253
rect 35200 11250 36000 11280
rect 34053 11248 36000 11250
rect 34053 11192 34058 11248
rect 34114 11192 36000 11248
rect 34053 11190 36000 11192
rect 34053 11187 34119 11190
rect 35200 11160 36000 11190
rect 9394 10912 9710 10913
rect 9394 10848 9400 10912
rect 9464 10848 9480 10912
rect 9544 10848 9560 10912
rect 9624 10848 9640 10912
rect 9704 10848 9710 10912
rect 9394 10847 9710 10848
rect 17842 10912 18158 10913
rect 17842 10848 17848 10912
rect 17912 10848 17928 10912
rect 17992 10848 18008 10912
rect 18072 10848 18088 10912
rect 18152 10848 18158 10912
rect 17842 10847 18158 10848
rect 26290 10912 26606 10913
rect 26290 10848 26296 10912
rect 26360 10848 26376 10912
rect 26440 10848 26456 10912
rect 26520 10848 26536 10912
rect 26600 10848 26606 10912
rect 26290 10847 26606 10848
rect 5170 10368 5486 10369
rect 5170 10304 5176 10368
rect 5240 10304 5256 10368
rect 5320 10304 5336 10368
rect 5400 10304 5416 10368
rect 5480 10304 5486 10368
rect 5170 10303 5486 10304
rect 13618 10368 13934 10369
rect 13618 10304 13624 10368
rect 13688 10304 13704 10368
rect 13768 10304 13784 10368
rect 13848 10304 13864 10368
rect 13928 10304 13934 10368
rect 13618 10303 13934 10304
rect 22066 10368 22382 10369
rect 22066 10304 22072 10368
rect 22136 10304 22152 10368
rect 22216 10304 22232 10368
rect 22296 10304 22312 10368
rect 22376 10304 22382 10368
rect 22066 10303 22382 10304
rect 30514 10368 30830 10369
rect 30514 10304 30520 10368
rect 30584 10304 30600 10368
rect 30664 10304 30680 10368
rect 30744 10304 30760 10368
rect 30824 10304 30830 10368
rect 30514 10303 30830 10304
rect 9394 9824 9710 9825
rect 9394 9760 9400 9824
rect 9464 9760 9480 9824
rect 9544 9760 9560 9824
rect 9624 9760 9640 9824
rect 9704 9760 9710 9824
rect 9394 9759 9710 9760
rect 17842 9824 18158 9825
rect 17842 9760 17848 9824
rect 17912 9760 17928 9824
rect 17992 9760 18008 9824
rect 18072 9760 18088 9824
rect 18152 9760 18158 9824
rect 17842 9759 18158 9760
rect 26290 9824 26606 9825
rect 26290 9760 26296 9824
rect 26360 9760 26376 9824
rect 26440 9760 26456 9824
rect 26520 9760 26536 9824
rect 26600 9760 26606 9824
rect 26290 9759 26606 9760
rect 5170 9280 5486 9281
rect 5170 9216 5176 9280
rect 5240 9216 5256 9280
rect 5320 9216 5336 9280
rect 5400 9216 5416 9280
rect 5480 9216 5486 9280
rect 5170 9215 5486 9216
rect 13618 9280 13934 9281
rect 13618 9216 13624 9280
rect 13688 9216 13704 9280
rect 13768 9216 13784 9280
rect 13848 9216 13864 9280
rect 13928 9216 13934 9280
rect 13618 9215 13934 9216
rect 22066 9280 22382 9281
rect 22066 9216 22072 9280
rect 22136 9216 22152 9280
rect 22216 9216 22232 9280
rect 22296 9216 22312 9280
rect 22376 9216 22382 9280
rect 22066 9215 22382 9216
rect 30514 9280 30830 9281
rect 30514 9216 30520 9280
rect 30584 9216 30600 9280
rect 30664 9216 30680 9280
rect 30744 9216 30760 9280
rect 30824 9216 30830 9280
rect 30514 9215 30830 9216
rect 34053 8802 34119 8805
rect 35200 8802 36000 8832
rect 34053 8800 36000 8802
rect 34053 8744 34058 8800
rect 34114 8744 36000 8800
rect 34053 8742 36000 8744
rect 34053 8739 34119 8742
rect 9394 8736 9710 8737
rect 9394 8672 9400 8736
rect 9464 8672 9480 8736
rect 9544 8672 9560 8736
rect 9624 8672 9640 8736
rect 9704 8672 9710 8736
rect 9394 8671 9710 8672
rect 17842 8736 18158 8737
rect 17842 8672 17848 8736
rect 17912 8672 17928 8736
rect 17992 8672 18008 8736
rect 18072 8672 18088 8736
rect 18152 8672 18158 8736
rect 17842 8671 18158 8672
rect 26290 8736 26606 8737
rect 26290 8672 26296 8736
rect 26360 8672 26376 8736
rect 26440 8672 26456 8736
rect 26520 8672 26536 8736
rect 26600 8672 26606 8736
rect 35200 8712 36000 8742
rect 26290 8671 26606 8672
rect 5170 8192 5486 8193
rect 5170 8128 5176 8192
rect 5240 8128 5256 8192
rect 5320 8128 5336 8192
rect 5400 8128 5416 8192
rect 5480 8128 5486 8192
rect 5170 8127 5486 8128
rect 13618 8192 13934 8193
rect 13618 8128 13624 8192
rect 13688 8128 13704 8192
rect 13768 8128 13784 8192
rect 13848 8128 13864 8192
rect 13928 8128 13934 8192
rect 13618 8127 13934 8128
rect 22066 8192 22382 8193
rect 22066 8128 22072 8192
rect 22136 8128 22152 8192
rect 22216 8128 22232 8192
rect 22296 8128 22312 8192
rect 22376 8128 22382 8192
rect 22066 8127 22382 8128
rect 30514 8192 30830 8193
rect 30514 8128 30520 8192
rect 30584 8128 30600 8192
rect 30664 8128 30680 8192
rect 30744 8128 30760 8192
rect 30824 8128 30830 8192
rect 30514 8127 30830 8128
rect 9394 7648 9710 7649
rect 0 7578 800 7608
rect 9394 7584 9400 7648
rect 9464 7584 9480 7648
rect 9544 7584 9560 7648
rect 9624 7584 9640 7648
rect 9704 7584 9710 7648
rect 9394 7583 9710 7584
rect 17842 7648 18158 7649
rect 17842 7584 17848 7648
rect 17912 7584 17928 7648
rect 17992 7584 18008 7648
rect 18072 7584 18088 7648
rect 18152 7584 18158 7648
rect 17842 7583 18158 7584
rect 26290 7648 26606 7649
rect 26290 7584 26296 7648
rect 26360 7584 26376 7648
rect 26440 7584 26456 7648
rect 26520 7584 26536 7648
rect 26600 7584 26606 7648
rect 26290 7583 26606 7584
rect 1393 7578 1459 7581
rect 0 7576 1459 7578
rect 0 7520 1398 7576
rect 1454 7520 1459 7576
rect 0 7518 1459 7520
rect 0 7488 800 7518
rect 1393 7515 1459 7518
rect 5170 7104 5486 7105
rect 5170 7040 5176 7104
rect 5240 7040 5256 7104
rect 5320 7040 5336 7104
rect 5400 7040 5416 7104
rect 5480 7040 5486 7104
rect 5170 7039 5486 7040
rect 13618 7104 13934 7105
rect 13618 7040 13624 7104
rect 13688 7040 13704 7104
rect 13768 7040 13784 7104
rect 13848 7040 13864 7104
rect 13928 7040 13934 7104
rect 13618 7039 13934 7040
rect 22066 7104 22382 7105
rect 22066 7040 22072 7104
rect 22136 7040 22152 7104
rect 22216 7040 22232 7104
rect 22296 7040 22312 7104
rect 22376 7040 22382 7104
rect 22066 7039 22382 7040
rect 30514 7104 30830 7105
rect 30514 7040 30520 7104
rect 30584 7040 30600 7104
rect 30664 7040 30680 7104
rect 30744 7040 30760 7104
rect 30824 7040 30830 7104
rect 30514 7039 30830 7040
rect 9394 6560 9710 6561
rect 9394 6496 9400 6560
rect 9464 6496 9480 6560
rect 9544 6496 9560 6560
rect 9624 6496 9640 6560
rect 9704 6496 9710 6560
rect 9394 6495 9710 6496
rect 17842 6560 18158 6561
rect 17842 6496 17848 6560
rect 17912 6496 17928 6560
rect 17992 6496 18008 6560
rect 18072 6496 18088 6560
rect 18152 6496 18158 6560
rect 17842 6495 18158 6496
rect 26290 6560 26606 6561
rect 26290 6496 26296 6560
rect 26360 6496 26376 6560
rect 26440 6496 26456 6560
rect 26520 6496 26536 6560
rect 26600 6496 26606 6560
rect 26290 6495 26606 6496
rect 34053 6354 34119 6357
rect 35200 6354 36000 6384
rect 34053 6352 36000 6354
rect 34053 6296 34058 6352
rect 34114 6296 36000 6352
rect 34053 6294 36000 6296
rect 34053 6291 34119 6294
rect 35200 6264 36000 6294
rect 5170 6016 5486 6017
rect 5170 5952 5176 6016
rect 5240 5952 5256 6016
rect 5320 5952 5336 6016
rect 5400 5952 5416 6016
rect 5480 5952 5486 6016
rect 5170 5951 5486 5952
rect 13618 6016 13934 6017
rect 13618 5952 13624 6016
rect 13688 5952 13704 6016
rect 13768 5952 13784 6016
rect 13848 5952 13864 6016
rect 13928 5952 13934 6016
rect 13618 5951 13934 5952
rect 22066 6016 22382 6017
rect 22066 5952 22072 6016
rect 22136 5952 22152 6016
rect 22216 5952 22232 6016
rect 22296 5952 22312 6016
rect 22376 5952 22382 6016
rect 22066 5951 22382 5952
rect 30514 6016 30830 6017
rect 30514 5952 30520 6016
rect 30584 5952 30600 6016
rect 30664 5952 30680 6016
rect 30744 5952 30760 6016
rect 30824 5952 30830 6016
rect 30514 5951 30830 5952
rect 9394 5472 9710 5473
rect 9394 5408 9400 5472
rect 9464 5408 9480 5472
rect 9544 5408 9560 5472
rect 9624 5408 9640 5472
rect 9704 5408 9710 5472
rect 9394 5407 9710 5408
rect 17842 5472 18158 5473
rect 17842 5408 17848 5472
rect 17912 5408 17928 5472
rect 17992 5408 18008 5472
rect 18072 5408 18088 5472
rect 18152 5408 18158 5472
rect 17842 5407 18158 5408
rect 26290 5472 26606 5473
rect 26290 5408 26296 5472
rect 26360 5408 26376 5472
rect 26440 5408 26456 5472
rect 26520 5408 26536 5472
rect 26600 5408 26606 5472
rect 26290 5407 26606 5408
rect 5170 4928 5486 4929
rect 5170 4864 5176 4928
rect 5240 4864 5256 4928
rect 5320 4864 5336 4928
rect 5400 4864 5416 4928
rect 5480 4864 5486 4928
rect 5170 4863 5486 4864
rect 13618 4928 13934 4929
rect 13618 4864 13624 4928
rect 13688 4864 13704 4928
rect 13768 4864 13784 4928
rect 13848 4864 13864 4928
rect 13928 4864 13934 4928
rect 13618 4863 13934 4864
rect 22066 4928 22382 4929
rect 22066 4864 22072 4928
rect 22136 4864 22152 4928
rect 22216 4864 22232 4928
rect 22296 4864 22312 4928
rect 22376 4864 22382 4928
rect 22066 4863 22382 4864
rect 30514 4928 30830 4929
rect 30514 4864 30520 4928
rect 30584 4864 30600 4928
rect 30664 4864 30680 4928
rect 30744 4864 30760 4928
rect 30824 4864 30830 4928
rect 30514 4863 30830 4864
rect 9394 4384 9710 4385
rect 9394 4320 9400 4384
rect 9464 4320 9480 4384
rect 9544 4320 9560 4384
rect 9624 4320 9640 4384
rect 9704 4320 9710 4384
rect 9394 4319 9710 4320
rect 17842 4384 18158 4385
rect 17842 4320 17848 4384
rect 17912 4320 17928 4384
rect 17992 4320 18008 4384
rect 18072 4320 18088 4384
rect 18152 4320 18158 4384
rect 17842 4319 18158 4320
rect 26290 4384 26606 4385
rect 26290 4320 26296 4384
rect 26360 4320 26376 4384
rect 26440 4320 26456 4384
rect 26520 4320 26536 4384
rect 26600 4320 26606 4384
rect 26290 4319 26606 4320
rect 34053 3906 34119 3909
rect 35200 3906 36000 3936
rect 34053 3904 36000 3906
rect 34053 3848 34058 3904
rect 34114 3848 36000 3904
rect 34053 3846 36000 3848
rect 34053 3843 34119 3846
rect 5170 3840 5486 3841
rect 5170 3776 5176 3840
rect 5240 3776 5256 3840
rect 5320 3776 5336 3840
rect 5400 3776 5416 3840
rect 5480 3776 5486 3840
rect 5170 3775 5486 3776
rect 13618 3840 13934 3841
rect 13618 3776 13624 3840
rect 13688 3776 13704 3840
rect 13768 3776 13784 3840
rect 13848 3776 13864 3840
rect 13928 3776 13934 3840
rect 13618 3775 13934 3776
rect 22066 3840 22382 3841
rect 22066 3776 22072 3840
rect 22136 3776 22152 3840
rect 22216 3776 22232 3840
rect 22296 3776 22312 3840
rect 22376 3776 22382 3840
rect 22066 3775 22382 3776
rect 30514 3840 30830 3841
rect 30514 3776 30520 3840
rect 30584 3776 30600 3840
rect 30664 3776 30680 3840
rect 30744 3776 30760 3840
rect 30824 3776 30830 3840
rect 35200 3816 36000 3846
rect 30514 3775 30830 3776
rect 9394 3296 9710 3297
rect 9394 3232 9400 3296
rect 9464 3232 9480 3296
rect 9544 3232 9560 3296
rect 9624 3232 9640 3296
rect 9704 3232 9710 3296
rect 9394 3231 9710 3232
rect 17842 3296 18158 3297
rect 17842 3232 17848 3296
rect 17912 3232 17928 3296
rect 17992 3232 18008 3296
rect 18072 3232 18088 3296
rect 18152 3232 18158 3296
rect 17842 3231 18158 3232
rect 26290 3296 26606 3297
rect 26290 3232 26296 3296
rect 26360 3232 26376 3296
rect 26440 3232 26456 3296
rect 26520 3232 26536 3296
rect 26600 3232 26606 3296
rect 26290 3231 26606 3232
rect 5170 2752 5486 2753
rect 0 2682 800 2712
rect 5170 2688 5176 2752
rect 5240 2688 5256 2752
rect 5320 2688 5336 2752
rect 5400 2688 5416 2752
rect 5480 2688 5486 2752
rect 5170 2687 5486 2688
rect 13618 2752 13934 2753
rect 13618 2688 13624 2752
rect 13688 2688 13704 2752
rect 13768 2688 13784 2752
rect 13848 2688 13864 2752
rect 13928 2688 13934 2752
rect 13618 2687 13934 2688
rect 22066 2752 22382 2753
rect 22066 2688 22072 2752
rect 22136 2688 22152 2752
rect 22216 2688 22232 2752
rect 22296 2688 22312 2752
rect 22376 2688 22382 2752
rect 22066 2687 22382 2688
rect 30514 2752 30830 2753
rect 30514 2688 30520 2752
rect 30584 2688 30600 2752
rect 30664 2688 30680 2752
rect 30744 2688 30760 2752
rect 30824 2688 30830 2752
rect 30514 2687 30830 2688
rect 3141 2682 3207 2685
rect 0 2680 3207 2682
rect 0 2624 3146 2680
rect 3202 2624 3207 2680
rect 0 2622 3207 2624
rect 0 2592 800 2622
rect 3141 2619 3207 2622
rect 9394 2208 9710 2209
rect 9394 2144 9400 2208
rect 9464 2144 9480 2208
rect 9544 2144 9560 2208
rect 9624 2144 9640 2208
rect 9704 2144 9710 2208
rect 9394 2143 9710 2144
rect 17842 2208 18158 2209
rect 17842 2144 17848 2208
rect 17912 2144 17928 2208
rect 17992 2144 18008 2208
rect 18072 2144 18088 2208
rect 18152 2144 18158 2208
rect 17842 2143 18158 2144
rect 26290 2208 26606 2209
rect 26290 2144 26296 2208
rect 26360 2144 26376 2208
rect 26440 2144 26456 2208
rect 26520 2144 26536 2208
rect 26600 2144 26606 2208
rect 26290 2143 26606 2144
rect 34053 1458 34119 1461
rect 35200 1458 36000 1488
rect 34053 1456 36000 1458
rect 34053 1400 34058 1456
rect 34114 1400 36000 1456
rect 34053 1398 36000 1400
rect 34053 1395 34119 1398
rect 35200 1368 36000 1398
<< via3 >>
rect 9400 17436 9464 17440
rect 9400 17380 9404 17436
rect 9404 17380 9460 17436
rect 9460 17380 9464 17436
rect 9400 17376 9464 17380
rect 9480 17436 9544 17440
rect 9480 17380 9484 17436
rect 9484 17380 9540 17436
rect 9540 17380 9544 17436
rect 9480 17376 9544 17380
rect 9560 17436 9624 17440
rect 9560 17380 9564 17436
rect 9564 17380 9620 17436
rect 9620 17380 9624 17436
rect 9560 17376 9624 17380
rect 9640 17436 9704 17440
rect 9640 17380 9644 17436
rect 9644 17380 9700 17436
rect 9700 17380 9704 17436
rect 9640 17376 9704 17380
rect 17848 17436 17912 17440
rect 17848 17380 17852 17436
rect 17852 17380 17908 17436
rect 17908 17380 17912 17436
rect 17848 17376 17912 17380
rect 17928 17436 17992 17440
rect 17928 17380 17932 17436
rect 17932 17380 17988 17436
rect 17988 17380 17992 17436
rect 17928 17376 17992 17380
rect 18008 17436 18072 17440
rect 18008 17380 18012 17436
rect 18012 17380 18068 17436
rect 18068 17380 18072 17436
rect 18008 17376 18072 17380
rect 18088 17436 18152 17440
rect 18088 17380 18092 17436
rect 18092 17380 18148 17436
rect 18148 17380 18152 17436
rect 18088 17376 18152 17380
rect 26296 17436 26360 17440
rect 26296 17380 26300 17436
rect 26300 17380 26356 17436
rect 26356 17380 26360 17436
rect 26296 17376 26360 17380
rect 26376 17436 26440 17440
rect 26376 17380 26380 17436
rect 26380 17380 26436 17436
rect 26436 17380 26440 17436
rect 26376 17376 26440 17380
rect 26456 17436 26520 17440
rect 26456 17380 26460 17436
rect 26460 17380 26516 17436
rect 26516 17380 26520 17436
rect 26456 17376 26520 17380
rect 26536 17436 26600 17440
rect 26536 17380 26540 17436
rect 26540 17380 26596 17436
rect 26596 17380 26600 17436
rect 26536 17376 26600 17380
rect 5176 16892 5240 16896
rect 5176 16836 5180 16892
rect 5180 16836 5236 16892
rect 5236 16836 5240 16892
rect 5176 16832 5240 16836
rect 5256 16892 5320 16896
rect 5256 16836 5260 16892
rect 5260 16836 5316 16892
rect 5316 16836 5320 16892
rect 5256 16832 5320 16836
rect 5336 16892 5400 16896
rect 5336 16836 5340 16892
rect 5340 16836 5396 16892
rect 5396 16836 5400 16892
rect 5336 16832 5400 16836
rect 5416 16892 5480 16896
rect 5416 16836 5420 16892
rect 5420 16836 5476 16892
rect 5476 16836 5480 16892
rect 5416 16832 5480 16836
rect 13624 16892 13688 16896
rect 13624 16836 13628 16892
rect 13628 16836 13684 16892
rect 13684 16836 13688 16892
rect 13624 16832 13688 16836
rect 13704 16892 13768 16896
rect 13704 16836 13708 16892
rect 13708 16836 13764 16892
rect 13764 16836 13768 16892
rect 13704 16832 13768 16836
rect 13784 16892 13848 16896
rect 13784 16836 13788 16892
rect 13788 16836 13844 16892
rect 13844 16836 13848 16892
rect 13784 16832 13848 16836
rect 13864 16892 13928 16896
rect 13864 16836 13868 16892
rect 13868 16836 13924 16892
rect 13924 16836 13928 16892
rect 13864 16832 13928 16836
rect 22072 16892 22136 16896
rect 22072 16836 22076 16892
rect 22076 16836 22132 16892
rect 22132 16836 22136 16892
rect 22072 16832 22136 16836
rect 22152 16892 22216 16896
rect 22152 16836 22156 16892
rect 22156 16836 22212 16892
rect 22212 16836 22216 16892
rect 22152 16832 22216 16836
rect 22232 16892 22296 16896
rect 22232 16836 22236 16892
rect 22236 16836 22292 16892
rect 22292 16836 22296 16892
rect 22232 16832 22296 16836
rect 22312 16892 22376 16896
rect 22312 16836 22316 16892
rect 22316 16836 22372 16892
rect 22372 16836 22376 16892
rect 22312 16832 22376 16836
rect 30520 16892 30584 16896
rect 30520 16836 30524 16892
rect 30524 16836 30580 16892
rect 30580 16836 30584 16892
rect 30520 16832 30584 16836
rect 30600 16892 30664 16896
rect 30600 16836 30604 16892
rect 30604 16836 30660 16892
rect 30660 16836 30664 16892
rect 30600 16832 30664 16836
rect 30680 16892 30744 16896
rect 30680 16836 30684 16892
rect 30684 16836 30740 16892
rect 30740 16836 30744 16892
rect 30680 16832 30744 16836
rect 30760 16892 30824 16896
rect 30760 16836 30764 16892
rect 30764 16836 30820 16892
rect 30820 16836 30824 16892
rect 30760 16832 30824 16836
rect 9400 16348 9464 16352
rect 9400 16292 9404 16348
rect 9404 16292 9460 16348
rect 9460 16292 9464 16348
rect 9400 16288 9464 16292
rect 9480 16348 9544 16352
rect 9480 16292 9484 16348
rect 9484 16292 9540 16348
rect 9540 16292 9544 16348
rect 9480 16288 9544 16292
rect 9560 16348 9624 16352
rect 9560 16292 9564 16348
rect 9564 16292 9620 16348
rect 9620 16292 9624 16348
rect 9560 16288 9624 16292
rect 9640 16348 9704 16352
rect 9640 16292 9644 16348
rect 9644 16292 9700 16348
rect 9700 16292 9704 16348
rect 9640 16288 9704 16292
rect 17848 16348 17912 16352
rect 17848 16292 17852 16348
rect 17852 16292 17908 16348
rect 17908 16292 17912 16348
rect 17848 16288 17912 16292
rect 17928 16348 17992 16352
rect 17928 16292 17932 16348
rect 17932 16292 17988 16348
rect 17988 16292 17992 16348
rect 17928 16288 17992 16292
rect 18008 16348 18072 16352
rect 18008 16292 18012 16348
rect 18012 16292 18068 16348
rect 18068 16292 18072 16348
rect 18008 16288 18072 16292
rect 18088 16348 18152 16352
rect 18088 16292 18092 16348
rect 18092 16292 18148 16348
rect 18148 16292 18152 16348
rect 18088 16288 18152 16292
rect 26296 16348 26360 16352
rect 26296 16292 26300 16348
rect 26300 16292 26356 16348
rect 26356 16292 26360 16348
rect 26296 16288 26360 16292
rect 26376 16348 26440 16352
rect 26376 16292 26380 16348
rect 26380 16292 26436 16348
rect 26436 16292 26440 16348
rect 26376 16288 26440 16292
rect 26456 16348 26520 16352
rect 26456 16292 26460 16348
rect 26460 16292 26516 16348
rect 26516 16292 26520 16348
rect 26456 16288 26520 16292
rect 26536 16348 26600 16352
rect 26536 16292 26540 16348
rect 26540 16292 26596 16348
rect 26596 16292 26600 16348
rect 26536 16288 26600 16292
rect 5176 15804 5240 15808
rect 5176 15748 5180 15804
rect 5180 15748 5236 15804
rect 5236 15748 5240 15804
rect 5176 15744 5240 15748
rect 5256 15804 5320 15808
rect 5256 15748 5260 15804
rect 5260 15748 5316 15804
rect 5316 15748 5320 15804
rect 5256 15744 5320 15748
rect 5336 15804 5400 15808
rect 5336 15748 5340 15804
rect 5340 15748 5396 15804
rect 5396 15748 5400 15804
rect 5336 15744 5400 15748
rect 5416 15804 5480 15808
rect 5416 15748 5420 15804
rect 5420 15748 5476 15804
rect 5476 15748 5480 15804
rect 5416 15744 5480 15748
rect 13624 15804 13688 15808
rect 13624 15748 13628 15804
rect 13628 15748 13684 15804
rect 13684 15748 13688 15804
rect 13624 15744 13688 15748
rect 13704 15804 13768 15808
rect 13704 15748 13708 15804
rect 13708 15748 13764 15804
rect 13764 15748 13768 15804
rect 13704 15744 13768 15748
rect 13784 15804 13848 15808
rect 13784 15748 13788 15804
rect 13788 15748 13844 15804
rect 13844 15748 13848 15804
rect 13784 15744 13848 15748
rect 13864 15804 13928 15808
rect 13864 15748 13868 15804
rect 13868 15748 13924 15804
rect 13924 15748 13928 15804
rect 13864 15744 13928 15748
rect 22072 15804 22136 15808
rect 22072 15748 22076 15804
rect 22076 15748 22132 15804
rect 22132 15748 22136 15804
rect 22072 15744 22136 15748
rect 22152 15804 22216 15808
rect 22152 15748 22156 15804
rect 22156 15748 22212 15804
rect 22212 15748 22216 15804
rect 22152 15744 22216 15748
rect 22232 15804 22296 15808
rect 22232 15748 22236 15804
rect 22236 15748 22292 15804
rect 22292 15748 22296 15804
rect 22232 15744 22296 15748
rect 22312 15804 22376 15808
rect 22312 15748 22316 15804
rect 22316 15748 22372 15804
rect 22372 15748 22376 15804
rect 22312 15744 22376 15748
rect 30520 15804 30584 15808
rect 30520 15748 30524 15804
rect 30524 15748 30580 15804
rect 30580 15748 30584 15804
rect 30520 15744 30584 15748
rect 30600 15804 30664 15808
rect 30600 15748 30604 15804
rect 30604 15748 30660 15804
rect 30660 15748 30664 15804
rect 30600 15744 30664 15748
rect 30680 15804 30744 15808
rect 30680 15748 30684 15804
rect 30684 15748 30740 15804
rect 30740 15748 30744 15804
rect 30680 15744 30744 15748
rect 30760 15804 30824 15808
rect 30760 15748 30764 15804
rect 30764 15748 30820 15804
rect 30820 15748 30824 15804
rect 30760 15744 30824 15748
rect 9400 15260 9464 15264
rect 9400 15204 9404 15260
rect 9404 15204 9460 15260
rect 9460 15204 9464 15260
rect 9400 15200 9464 15204
rect 9480 15260 9544 15264
rect 9480 15204 9484 15260
rect 9484 15204 9540 15260
rect 9540 15204 9544 15260
rect 9480 15200 9544 15204
rect 9560 15260 9624 15264
rect 9560 15204 9564 15260
rect 9564 15204 9620 15260
rect 9620 15204 9624 15260
rect 9560 15200 9624 15204
rect 9640 15260 9704 15264
rect 9640 15204 9644 15260
rect 9644 15204 9700 15260
rect 9700 15204 9704 15260
rect 9640 15200 9704 15204
rect 17848 15260 17912 15264
rect 17848 15204 17852 15260
rect 17852 15204 17908 15260
rect 17908 15204 17912 15260
rect 17848 15200 17912 15204
rect 17928 15260 17992 15264
rect 17928 15204 17932 15260
rect 17932 15204 17988 15260
rect 17988 15204 17992 15260
rect 17928 15200 17992 15204
rect 18008 15260 18072 15264
rect 18008 15204 18012 15260
rect 18012 15204 18068 15260
rect 18068 15204 18072 15260
rect 18008 15200 18072 15204
rect 18088 15260 18152 15264
rect 18088 15204 18092 15260
rect 18092 15204 18148 15260
rect 18148 15204 18152 15260
rect 18088 15200 18152 15204
rect 26296 15260 26360 15264
rect 26296 15204 26300 15260
rect 26300 15204 26356 15260
rect 26356 15204 26360 15260
rect 26296 15200 26360 15204
rect 26376 15260 26440 15264
rect 26376 15204 26380 15260
rect 26380 15204 26436 15260
rect 26436 15204 26440 15260
rect 26376 15200 26440 15204
rect 26456 15260 26520 15264
rect 26456 15204 26460 15260
rect 26460 15204 26516 15260
rect 26516 15204 26520 15260
rect 26456 15200 26520 15204
rect 26536 15260 26600 15264
rect 26536 15204 26540 15260
rect 26540 15204 26596 15260
rect 26596 15204 26600 15260
rect 26536 15200 26600 15204
rect 5176 14716 5240 14720
rect 5176 14660 5180 14716
rect 5180 14660 5236 14716
rect 5236 14660 5240 14716
rect 5176 14656 5240 14660
rect 5256 14716 5320 14720
rect 5256 14660 5260 14716
rect 5260 14660 5316 14716
rect 5316 14660 5320 14716
rect 5256 14656 5320 14660
rect 5336 14716 5400 14720
rect 5336 14660 5340 14716
rect 5340 14660 5396 14716
rect 5396 14660 5400 14716
rect 5336 14656 5400 14660
rect 5416 14716 5480 14720
rect 5416 14660 5420 14716
rect 5420 14660 5476 14716
rect 5476 14660 5480 14716
rect 5416 14656 5480 14660
rect 13624 14716 13688 14720
rect 13624 14660 13628 14716
rect 13628 14660 13684 14716
rect 13684 14660 13688 14716
rect 13624 14656 13688 14660
rect 13704 14716 13768 14720
rect 13704 14660 13708 14716
rect 13708 14660 13764 14716
rect 13764 14660 13768 14716
rect 13704 14656 13768 14660
rect 13784 14716 13848 14720
rect 13784 14660 13788 14716
rect 13788 14660 13844 14716
rect 13844 14660 13848 14716
rect 13784 14656 13848 14660
rect 13864 14716 13928 14720
rect 13864 14660 13868 14716
rect 13868 14660 13924 14716
rect 13924 14660 13928 14716
rect 13864 14656 13928 14660
rect 22072 14716 22136 14720
rect 22072 14660 22076 14716
rect 22076 14660 22132 14716
rect 22132 14660 22136 14716
rect 22072 14656 22136 14660
rect 22152 14716 22216 14720
rect 22152 14660 22156 14716
rect 22156 14660 22212 14716
rect 22212 14660 22216 14716
rect 22152 14656 22216 14660
rect 22232 14716 22296 14720
rect 22232 14660 22236 14716
rect 22236 14660 22292 14716
rect 22292 14660 22296 14716
rect 22232 14656 22296 14660
rect 22312 14716 22376 14720
rect 22312 14660 22316 14716
rect 22316 14660 22372 14716
rect 22372 14660 22376 14716
rect 22312 14656 22376 14660
rect 30520 14716 30584 14720
rect 30520 14660 30524 14716
rect 30524 14660 30580 14716
rect 30580 14660 30584 14716
rect 30520 14656 30584 14660
rect 30600 14716 30664 14720
rect 30600 14660 30604 14716
rect 30604 14660 30660 14716
rect 30660 14660 30664 14716
rect 30600 14656 30664 14660
rect 30680 14716 30744 14720
rect 30680 14660 30684 14716
rect 30684 14660 30740 14716
rect 30740 14660 30744 14716
rect 30680 14656 30744 14660
rect 30760 14716 30824 14720
rect 30760 14660 30764 14716
rect 30764 14660 30820 14716
rect 30820 14660 30824 14716
rect 30760 14656 30824 14660
rect 9400 14172 9464 14176
rect 9400 14116 9404 14172
rect 9404 14116 9460 14172
rect 9460 14116 9464 14172
rect 9400 14112 9464 14116
rect 9480 14172 9544 14176
rect 9480 14116 9484 14172
rect 9484 14116 9540 14172
rect 9540 14116 9544 14172
rect 9480 14112 9544 14116
rect 9560 14172 9624 14176
rect 9560 14116 9564 14172
rect 9564 14116 9620 14172
rect 9620 14116 9624 14172
rect 9560 14112 9624 14116
rect 9640 14172 9704 14176
rect 9640 14116 9644 14172
rect 9644 14116 9700 14172
rect 9700 14116 9704 14172
rect 9640 14112 9704 14116
rect 17848 14172 17912 14176
rect 17848 14116 17852 14172
rect 17852 14116 17908 14172
rect 17908 14116 17912 14172
rect 17848 14112 17912 14116
rect 17928 14172 17992 14176
rect 17928 14116 17932 14172
rect 17932 14116 17988 14172
rect 17988 14116 17992 14172
rect 17928 14112 17992 14116
rect 18008 14172 18072 14176
rect 18008 14116 18012 14172
rect 18012 14116 18068 14172
rect 18068 14116 18072 14172
rect 18008 14112 18072 14116
rect 18088 14172 18152 14176
rect 18088 14116 18092 14172
rect 18092 14116 18148 14172
rect 18148 14116 18152 14172
rect 18088 14112 18152 14116
rect 26296 14172 26360 14176
rect 26296 14116 26300 14172
rect 26300 14116 26356 14172
rect 26356 14116 26360 14172
rect 26296 14112 26360 14116
rect 26376 14172 26440 14176
rect 26376 14116 26380 14172
rect 26380 14116 26436 14172
rect 26436 14116 26440 14172
rect 26376 14112 26440 14116
rect 26456 14172 26520 14176
rect 26456 14116 26460 14172
rect 26460 14116 26516 14172
rect 26516 14116 26520 14172
rect 26456 14112 26520 14116
rect 26536 14172 26600 14176
rect 26536 14116 26540 14172
rect 26540 14116 26596 14172
rect 26596 14116 26600 14172
rect 26536 14112 26600 14116
rect 5176 13628 5240 13632
rect 5176 13572 5180 13628
rect 5180 13572 5236 13628
rect 5236 13572 5240 13628
rect 5176 13568 5240 13572
rect 5256 13628 5320 13632
rect 5256 13572 5260 13628
rect 5260 13572 5316 13628
rect 5316 13572 5320 13628
rect 5256 13568 5320 13572
rect 5336 13628 5400 13632
rect 5336 13572 5340 13628
rect 5340 13572 5396 13628
rect 5396 13572 5400 13628
rect 5336 13568 5400 13572
rect 5416 13628 5480 13632
rect 5416 13572 5420 13628
rect 5420 13572 5476 13628
rect 5476 13572 5480 13628
rect 5416 13568 5480 13572
rect 13624 13628 13688 13632
rect 13624 13572 13628 13628
rect 13628 13572 13684 13628
rect 13684 13572 13688 13628
rect 13624 13568 13688 13572
rect 13704 13628 13768 13632
rect 13704 13572 13708 13628
rect 13708 13572 13764 13628
rect 13764 13572 13768 13628
rect 13704 13568 13768 13572
rect 13784 13628 13848 13632
rect 13784 13572 13788 13628
rect 13788 13572 13844 13628
rect 13844 13572 13848 13628
rect 13784 13568 13848 13572
rect 13864 13628 13928 13632
rect 13864 13572 13868 13628
rect 13868 13572 13924 13628
rect 13924 13572 13928 13628
rect 13864 13568 13928 13572
rect 22072 13628 22136 13632
rect 22072 13572 22076 13628
rect 22076 13572 22132 13628
rect 22132 13572 22136 13628
rect 22072 13568 22136 13572
rect 22152 13628 22216 13632
rect 22152 13572 22156 13628
rect 22156 13572 22212 13628
rect 22212 13572 22216 13628
rect 22152 13568 22216 13572
rect 22232 13628 22296 13632
rect 22232 13572 22236 13628
rect 22236 13572 22292 13628
rect 22292 13572 22296 13628
rect 22232 13568 22296 13572
rect 22312 13628 22376 13632
rect 22312 13572 22316 13628
rect 22316 13572 22372 13628
rect 22372 13572 22376 13628
rect 22312 13568 22376 13572
rect 30520 13628 30584 13632
rect 30520 13572 30524 13628
rect 30524 13572 30580 13628
rect 30580 13572 30584 13628
rect 30520 13568 30584 13572
rect 30600 13628 30664 13632
rect 30600 13572 30604 13628
rect 30604 13572 30660 13628
rect 30660 13572 30664 13628
rect 30600 13568 30664 13572
rect 30680 13628 30744 13632
rect 30680 13572 30684 13628
rect 30684 13572 30740 13628
rect 30740 13572 30744 13628
rect 30680 13568 30744 13572
rect 30760 13628 30824 13632
rect 30760 13572 30764 13628
rect 30764 13572 30820 13628
rect 30820 13572 30824 13628
rect 30760 13568 30824 13572
rect 9400 13084 9464 13088
rect 9400 13028 9404 13084
rect 9404 13028 9460 13084
rect 9460 13028 9464 13084
rect 9400 13024 9464 13028
rect 9480 13084 9544 13088
rect 9480 13028 9484 13084
rect 9484 13028 9540 13084
rect 9540 13028 9544 13084
rect 9480 13024 9544 13028
rect 9560 13084 9624 13088
rect 9560 13028 9564 13084
rect 9564 13028 9620 13084
rect 9620 13028 9624 13084
rect 9560 13024 9624 13028
rect 9640 13084 9704 13088
rect 9640 13028 9644 13084
rect 9644 13028 9700 13084
rect 9700 13028 9704 13084
rect 9640 13024 9704 13028
rect 17848 13084 17912 13088
rect 17848 13028 17852 13084
rect 17852 13028 17908 13084
rect 17908 13028 17912 13084
rect 17848 13024 17912 13028
rect 17928 13084 17992 13088
rect 17928 13028 17932 13084
rect 17932 13028 17988 13084
rect 17988 13028 17992 13084
rect 17928 13024 17992 13028
rect 18008 13084 18072 13088
rect 18008 13028 18012 13084
rect 18012 13028 18068 13084
rect 18068 13028 18072 13084
rect 18008 13024 18072 13028
rect 18088 13084 18152 13088
rect 18088 13028 18092 13084
rect 18092 13028 18148 13084
rect 18148 13028 18152 13084
rect 18088 13024 18152 13028
rect 26296 13084 26360 13088
rect 26296 13028 26300 13084
rect 26300 13028 26356 13084
rect 26356 13028 26360 13084
rect 26296 13024 26360 13028
rect 26376 13084 26440 13088
rect 26376 13028 26380 13084
rect 26380 13028 26436 13084
rect 26436 13028 26440 13084
rect 26376 13024 26440 13028
rect 26456 13084 26520 13088
rect 26456 13028 26460 13084
rect 26460 13028 26516 13084
rect 26516 13028 26520 13084
rect 26456 13024 26520 13028
rect 26536 13084 26600 13088
rect 26536 13028 26540 13084
rect 26540 13028 26596 13084
rect 26596 13028 26600 13084
rect 26536 13024 26600 13028
rect 5176 12540 5240 12544
rect 5176 12484 5180 12540
rect 5180 12484 5236 12540
rect 5236 12484 5240 12540
rect 5176 12480 5240 12484
rect 5256 12540 5320 12544
rect 5256 12484 5260 12540
rect 5260 12484 5316 12540
rect 5316 12484 5320 12540
rect 5256 12480 5320 12484
rect 5336 12540 5400 12544
rect 5336 12484 5340 12540
rect 5340 12484 5396 12540
rect 5396 12484 5400 12540
rect 5336 12480 5400 12484
rect 5416 12540 5480 12544
rect 5416 12484 5420 12540
rect 5420 12484 5476 12540
rect 5476 12484 5480 12540
rect 5416 12480 5480 12484
rect 13624 12540 13688 12544
rect 13624 12484 13628 12540
rect 13628 12484 13684 12540
rect 13684 12484 13688 12540
rect 13624 12480 13688 12484
rect 13704 12540 13768 12544
rect 13704 12484 13708 12540
rect 13708 12484 13764 12540
rect 13764 12484 13768 12540
rect 13704 12480 13768 12484
rect 13784 12540 13848 12544
rect 13784 12484 13788 12540
rect 13788 12484 13844 12540
rect 13844 12484 13848 12540
rect 13784 12480 13848 12484
rect 13864 12540 13928 12544
rect 13864 12484 13868 12540
rect 13868 12484 13924 12540
rect 13924 12484 13928 12540
rect 13864 12480 13928 12484
rect 22072 12540 22136 12544
rect 22072 12484 22076 12540
rect 22076 12484 22132 12540
rect 22132 12484 22136 12540
rect 22072 12480 22136 12484
rect 22152 12540 22216 12544
rect 22152 12484 22156 12540
rect 22156 12484 22212 12540
rect 22212 12484 22216 12540
rect 22152 12480 22216 12484
rect 22232 12540 22296 12544
rect 22232 12484 22236 12540
rect 22236 12484 22292 12540
rect 22292 12484 22296 12540
rect 22232 12480 22296 12484
rect 22312 12540 22376 12544
rect 22312 12484 22316 12540
rect 22316 12484 22372 12540
rect 22372 12484 22376 12540
rect 22312 12480 22376 12484
rect 30520 12540 30584 12544
rect 30520 12484 30524 12540
rect 30524 12484 30580 12540
rect 30580 12484 30584 12540
rect 30520 12480 30584 12484
rect 30600 12540 30664 12544
rect 30600 12484 30604 12540
rect 30604 12484 30660 12540
rect 30660 12484 30664 12540
rect 30600 12480 30664 12484
rect 30680 12540 30744 12544
rect 30680 12484 30684 12540
rect 30684 12484 30740 12540
rect 30740 12484 30744 12540
rect 30680 12480 30744 12484
rect 30760 12540 30824 12544
rect 30760 12484 30764 12540
rect 30764 12484 30820 12540
rect 30820 12484 30824 12540
rect 30760 12480 30824 12484
rect 9400 11996 9464 12000
rect 9400 11940 9404 11996
rect 9404 11940 9460 11996
rect 9460 11940 9464 11996
rect 9400 11936 9464 11940
rect 9480 11996 9544 12000
rect 9480 11940 9484 11996
rect 9484 11940 9540 11996
rect 9540 11940 9544 11996
rect 9480 11936 9544 11940
rect 9560 11996 9624 12000
rect 9560 11940 9564 11996
rect 9564 11940 9620 11996
rect 9620 11940 9624 11996
rect 9560 11936 9624 11940
rect 9640 11996 9704 12000
rect 9640 11940 9644 11996
rect 9644 11940 9700 11996
rect 9700 11940 9704 11996
rect 9640 11936 9704 11940
rect 17848 11996 17912 12000
rect 17848 11940 17852 11996
rect 17852 11940 17908 11996
rect 17908 11940 17912 11996
rect 17848 11936 17912 11940
rect 17928 11996 17992 12000
rect 17928 11940 17932 11996
rect 17932 11940 17988 11996
rect 17988 11940 17992 11996
rect 17928 11936 17992 11940
rect 18008 11996 18072 12000
rect 18008 11940 18012 11996
rect 18012 11940 18068 11996
rect 18068 11940 18072 11996
rect 18008 11936 18072 11940
rect 18088 11996 18152 12000
rect 18088 11940 18092 11996
rect 18092 11940 18148 11996
rect 18148 11940 18152 11996
rect 18088 11936 18152 11940
rect 26296 11996 26360 12000
rect 26296 11940 26300 11996
rect 26300 11940 26356 11996
rect 26356 11940 26360 11996
rect 26296 11936 26360 11940
rect 26376 11996 26440 12000
rect 26376 11940 26380 11996
rect 26380 11940 26436 11996
rect 26436 11940 26440 11996
rect 26376 11936 26440 11940
rect 26456 11996 26520 12000
rect 26456 11940 26460 11996
rect 26460 11940 26516 11996
rect 26516 11940 26520 11996
rect 26456 11936 26520 11940
rect 26536 11996 26600 12000
rect 26536 11940 26540 11996
rect 26540 11940 26596 11996
rect 26596 11940 26600 11996
rect 26536 11936 26600 11940
rect 5176 11452 5240 11456
rect 5176 11396 5180 11452
rect 5180 11396 5236 11452
rect 5236 11396 5240 11452
rect 5176 11392 5240 11396
rect 5256 11452 5320 11456
rect 5256 11396 5260 11452
rect 5260 11396 5316 11452
rect 5316 11396 5320 11452
rect 5256 11392 5320 11396
rect 5336 11452 5400 11456
rect 5336 11396 5340 11452
rect 5340 11396 5396 11452
rect 5396 11396 5400 11452
rect 5336 11392 5400 11396
rect 5416 11452 5480 11456
rect 5416 11396 5420 11452
rect 5420 11396 5476 11452
rect 5476 11396 5480 11452
rect 5416 11392 5480 11396
rect 13624 11452 13688 11456
rect 13624 11396 13628 11452
rect 13628 11396 13684 11452
rect 13684 11396 13688 11452
rect 13624 11392 13688 11396
rect 13704 11452 13768 11456
rect 13704 11396 13708 11452
rect 13708 11396 13764 11452
rect 13764 11396 13768 11452
rect 13704 11392 13768 11396
rect 13784 11452 13848 11456
rect 13784 11396 13788 11452
rect 13788 11396 13844 11452
rect 13844 11396 13848 11452
rect 13784 11392 13848 11396
rect 13864 11452 13928 11456
rect 13864 11396 13868 11452
rect 13868 11396 13924 11452
rect 13924 11396 13928 11452
rect 13864 11392 13928 11396
rect 22072 11452 22136 11456
rect 22072 11396 22076 11452
rect 22076 11396 22132 11452
rect 22132 11396 22136 11452
rect 22072 11392 22136 11396
rect 22152 11452 22216 11456
rect 22152 11396 22156 11452
rect 22156 11396 22212 11452
rect 22212 11396 22216 11452
rect 22152 11392 22216 11396
rect 22232 11452 22296 11456
rect 22232 11396 22236 11452
rect 22236 11396 22292 11452
rect 22292 11396 22296 11452
rect 22232 11392 22296 11396
rect 22312 11452 22376 11456
rect 22312 11396 22316 11452
rect 22316 11396 22372 11452
rect 22372 11396 22376 11452
rect 22312 11392 22376 11396
rect 30520 11452 30584 11456
rect 30520 11396 30524 11452
rect 30524 11396 30580 11452
rect 30580 11396 30584 11452
rect 30520 11392 30584 11396
rect 30600 11452 30664 11456
rect 30600 11396 30604 11452
rect 30604 11396 30660 11452
rect 30660 11396 30664 11452
rect 30600 11392 30664 11396
rect 30680 11452 30744 11456
rect 30680 11396 30684 11452
rect 30684 11396 30740 11452
rect 30740 11396 30744 11452
rect 30680 11392 30744 11396
rect 30760 11452 30824 11456
rect 30760 11396 30764 11452
rect 30764 11396 30820 11452
rect 30820 11396 30824 11452
rect 30760 11392 30824 11396
rect 9400 10908 9464 10912
rect 9400 10852 9404 10908
rect 9404 10852 9460 10908
rect 9460 10852 9464 10908
rect 9400 10848 9464 10852
rect 9480 10908 9544 10912
rect 9480 10852 9484 10908
rect 9484 10852 9540 10908
rect 9540 10852 9544 10908
rect 9480 10848 9544 10852
rect 9560 10908 9624 10912
rect 9560 10852 9564 10908
rect 9564 10852 9620 10908
rect 9620 10852 9624 10908
rect 9560 10848 9624 10852
rect 9640 10908 9704 10912
rect 9640 10852 9644 10908
rect 9644 10852 9700 10908
rect 9700 10852 9704 10908
rect 9640 10848 9704 10852
rect 17848 10908 17912 10912
rect 17848 10852 17852 10908
rect 17852 10852 17908 10908
rect 17908 10852 17912 10908
rect 17848 10848 17912 10852
rect 17928 10908 17992 10912
rect 17928 10852 17932 10908
rect 17932 10852 17988 10908
rect 17988 10852 17992 10908
rect 17928 10848 17992 10852
rect 18008 10908 18072 10912
rect 18008 10852 18012 10908
rect 18012 10852 18068 10908
rect 18068 10852 18072 10908
rect 18008 10848 18072 10852
rect 18088 10908 18152 10912
rect 18088 10852 18092 10908
rect 18092 10852 18148 10908
rect 18148 10852 18152 10908
rect 18088 10848 18152 10852
rect 26296 10908 26360 10912
rect 26296 10852 26300 10908
rect 26300 10852 26356 10908
rect 26356 10852 26360 10908
rect 26296 10848 26360 10852
rect 26376 10908 26440 10912
rect 26376 10852 26380 10908
rect 26380 10852 26436 10908
rect 26436 10852 26440 10908
rect 26376 10848 26440 10852
rect 26456 10908 26520 10912
rect 26456 10852 26460 10908
rect 26460 10852 26516 10908
rect 26516 10852 26520 10908
rect 26456 10848 26520 10852
rect 26536 10908 26600 10912
rect 26536 10852 26540 10908
rect 26540 10852 26596 10908
rect 26596 10852 26600 10908
rect 26536 10848 26600 10852
rect 5176 10364 5240 10368
rect 5176 10308 5180 10364
rect 5180 10308 5236 10364
rect 5236 10308 5240 10364
rect 5176 10304 5240 10308
rect 5256 10364 5320 10368
rect 5256 10308 5260 10364
rect 5260 10308 5316 10364
rect 5316 10308 5320 10364
rect 5256 10304 5320 10308
rect 5336 10364 5400 10368
rect 5336 10308 5340 10364
rect 5340 10308 5396 10364
rect 5396 10308 5400 10364
rect 5336 10304 5400 10308
rect 5416 10364 5480 10368
rect 5416 10308 5420 10364
rect 5420 10308 5476 10364
rect 5476 10308 5480 10364
rect 5416 10304 5480 10308
rect 13624 10364 13688 10368
rect 13624 10308 13628 10364
rect 13628 10308 13684 10364
rect 13684 10308 13688 10364
rect 13624 10304 13688 10308
rect 13704 10364 13768 10368
rect 13704 10308 13708 10364
rect 13708 10308 13764 10364
rect 13764 10308 13768 10364
rect 13704 10304 13768 10308
rect 13784 10364 13848 10368
rect 13784 10308 13788 10364
rect 13788 10308 13844 10364
rect 13844 10308 13848 10364
rect 13784 10304 13848 10308
rect 13864 10364 13928 10368
rect 13864 10308 13868 10364
rect 13868 10308 13924 10364
rect 13924 10308 13928 10364
rect 13864 10304 13928 10308
rect 22072 10364 22136 10368
rect 22072 10308 22076 10364
rect 22076 10308 22132 10364
rect 22132 10308 22136 10364
rect 22072 10304 22136 10308
rect 22152 10364 22216 10368
rect 22152 10308 22156 10364
rect 22156 10308 22212 10364
rect 22212 10308 22216 10364
rect 22152 10304 22216 10308
rect 22232 10364 22296 10368
rect 22232 10308 22236 10364
rect 22236 10308 22292 10364
rect 22292 10308 22296 10364
rect 22232 10304 22296 10308
rect 22312 10364 22376 10368
rect 22312 10308 22316 10364
rect 22316 10308 22372 10364
rect 22372 10308 22376 10364
rect 22312 10304 22376 10308
rect 30520 10364 30584 10368
rect 30520 10308 30524 10364
rect 30524 10308 30580 10364
rect 30580 10308 30584 10364
rect 30520 10304 30584 10308
rect 30600 10364 30664 10368
rect 30600 10308 30604 10364
rect 30604 10308 30660 10364
rect 30660 10308 30664 10364
rect 30600 10304 30664 10308
rect 30680 10364 30744 10368
rect 30680 10308 30684 10364
rect 30684 10308 30740 10364
rect 30740 10308 30744 10364
rect 30680 10304 30744 10308
rect 30760 10364 30824 10368
rect 30760 10308 30764 10364
rect 30764 10308 30820 10364
rect 30820 10308 30824 10364
rect 30760 10304 30824 10308
rect 9400 9820 9464 9824
rect 9400 9764 9404 9820
rect 9404 9764 9460 9820
rect 9460 9764 9464 9820
rect 9400 9760 9464 9764
rect 9480 9820 9544 9824
rect 9480 9764 9484 9820
rect 9484 9764 9540 9820
rect 9540 9764 9544 9820
rect 9480 9760 9544 9764
rect 9560 9820 9624 9824
rect 9560 9764 9564 9820
rect 9564 9764 9620 9820
rect 9620 9764 9624 9820
rect 9560 9760 9624 9764
rect 9640 9820 9704 9824
rect 9640 9764 9644 9820
rect 9644 9764 9700 9820
rect 9700 9764 9704 9820
rect 9640 9760 9704 9764
rect 17848 9820 17912 9824
rect 17848 9764 17852 9820
rect 17852 9764 17908 9820
rect 17908 9764 17912 9820
rect 17848 9760 17912 9764
rect 17928 9820 17992 9824
rect 17928 9764 17932 9820
rect 17932 9764 17988 9820
rect 17988 9764 17992 9820
rect 17928 9760 17992 9764
rect 18008 9820 18072 9824
rect 18008 9764 18012 9820
rect 18012 9764 18068 9820
rect 18068 9764 18072 9820
rect 18008 9760 18072 9764
rect 18088 9820 18152 9824
rect 18088 9764 18092 9820
rect 18092 9764 18148 9820
rect 18148 9764 18152 9820
rect 18088 9760 18152 9764
rect 26296 9820 26360 9824
rect 26296 9764 26300 9820
rect 26300 9764 26356 9820
rect 26356 9764 26360 9820
rect 26296 9760 26360 9764
rect 26376 9820 26440 9824
rect 26376 9764 26380 9820
rect 26380 9764 26436 9820
rect 26436 9764 26440 9820
rect 26376 9760 26440 9764
rect 26456 9820 26520 9824
rect 26456 9764 26460 9820
rect 26460 9764 26516 9820
rect 26516 9764 26520 9820
rect 26456 9760 26520 9764
rect 26536 9820 26600 9824
rect 26536 9764 26540 9820
rect 26540 9764 26596 9820
rect 26596 9764 26600 9820
rect 26536 9760 26600 9764
rect 5176 9276 5240 9280
rect 5176 9220 5180 9276
rect 5180 9220 5236 9276
rect 5236 9220 5240 9276
rect 5176 9216 5240 9220
rect 5256 9276 5320 9280
rect 5256 9220 5260 9276
rect 5260 9220 5316 9276
rect 5316 9220 5320 9276
rect 5256 9216 5320 9220
rect 5336 9276 5400 9280
rect 5336 9220 5340 9276
rect 5340 9220 5396 9276
rect 5396 9220 5400 9276
rect 5336 9216 5400 9220
rect 5416 9276 5480 9280
rect 5416 9220 5420 9276
rect 5420 9220 5476 9276
rect 5476 9220 5480 9276
rect 5416 9216 5480 9220
rect 13624 9276 13688 9280
rect 13624 9220 13628 9276
rect 13628 9220 13684 9276
rect 13684 9220 13688 9276
rect 13624 9216 13688 9220
rect 13704 9276 13768 9280
rect 13704 9220 13708 9276
rect 13708 9220 13764 9276
rect 13764 9220 13768 9276
rect 13704 9216 13768 9220
rect 13784 9276 13848 9280
rect 13784 9220 13788 9276
rect 13788 9220 13844 9276
rect 13844 9220 13848 9276
rect 13784 9216 13848 9220
rect 13864 9276 13928 9280
rect 13864 9220 13868 9276
rect 13868 9220 13924 9276
rect 13924 9220 13928 9276
rect 13864 9216 13928 9220
rect 22072 9276 22136 9280
rect 22072 9220 22076 9276
rect 22076 9220 22132 9276
rect 22132 9220 22136 9276
rect 22072 9216 22136 9220
rect 22152 9276 22216 9280
rect 22152 9220 22156 9276
rect 22156 9220 22212 9276
rect 22212 9220 22216 9276
rect 22152 9216 22216 9220
rect 22232 9276 22296 9280
rect 22232 9220 22236 9276
rect 22236 9220 22292 9276
rect 22292 9220 22296 9276
rect 22232 9216 22296 9220
rect 22312 9276 22376 9280
rect 22312 9220 22316 9276
rect 22316 9220 22372 9276
rect 22372 9220 22376 9276
rect 22312 9216 22376 9220
rect 30520 9276 30584 9280
rect 30520 9220 30524 9276
rect 30524 9220 30580 9276
rect 30580 9220 30584 9276
rect 30520 9216 30584 9220
rect 30600 9276 30664 9280
rect 30600 9220 30604 9276
rect 30604 9220 30660 9276
rect 30660 9220 30664 9276
rect 30600 9216 30664 9220
rect 30680 9276 30744 9280
rect 30680 9220 30684 9276
rect 30684 9220 30740 9276
rect 30740 9220 30744 9276
rect 30680 9216 30744 9220
rect 30760 9276 30824 9280
rect 30760 9220 30764 9276
rect 30764 9220 30820 9276
rect 30820 9220 30824 9276
rect 30760 9216 30824 9220
rect 9400 8732 9464 8736
rect 9400 8676 9404 8732
rect 9404 8676 9460 8732
rect 9460 8676 9464 8732
rect 9400 8672 9464 8676
rect 9480 8732 9544 8736
rect 9480 8676 9484 8732
rect 9484 8676 9540 8732
rect 9540 8676 9544 8732
rect 9480 8672 9544 8676
rect 9560 8732 9624 8736
rect 9560 8676 9564 8732
rect 9564 8676 9620 8732
rect 9620 8676 9624 8732
rect 9560 8672 9624 8676
rect 9640 8732 9704 8736
rect 9640 8676 9644 8732
rect 9644 8676 9700 8732
rect 9700 8676 9704 8732
rect 9640 8672 9704 8676
rect 17848 8732 17912 8736
rect 17848 8676 17852 8732
rect 17852 8676 17908 8732
rect 17908 8676 17912 8732
rect 17848 8672 17912 8676
rect 17928 8732 17992 8736
rect 17928 8676 17932 8732
rect 17932 8676 17988 8732
rect 17988 8676 17992 8732
rect 17928 8672 17992 8676
rect 18008 8732 18072 8736
rect 18008 8676 18012 8732
rect 18012 8676 18068 8732
rect 18068 8676 18072 8732
rect 18008 8672 18072 8676
rect 18088 8732 18152 8736
rect 18088 8676 18092 8732
rect 18092 8676 18148 8732
rect 18148 8676 18152 8732
rect 18088 8672 18152 8676
rect 26296 8732 26360 8736
rect 26296 8676 26300 8732
rect 26300 8676 26356 8732
rect 26356 8676 26360 8732
rect 26296 8672 26360 8676
rect 26376 8732 26440 8736
rect 26376 8676 26380 8732
rect 26380 8676 26436 8732
rect 26436 8676 26440 8732
rect 26376 8672 26440 8676
rect 26456 8732 26520 8736
rect 26456 8676 26460 8732
rect 26460 8676 26516 8732
rect 26516 8676 26520 8732
rect 26456 8672 26520 8676
rect 26536 8732 26600 8736
rect 26536 8676 26540 8732
rect 26540 8676 26596 8732
rect 26596 8676 26600 8732
rect 26536 8672 26600 8676
rect 5176 8188 5240 8192
rect 5176 8132 5180 8188
rect 5180 8132 5236 8188
rect 5236 8132 5240 8188
rect 5176 8128 5240 8132
rect 5256 8188 5320 8192
rect 5256 8132 5260 8188
rect 5260 8132 5316 8188
rect 5316 8132 5320 8188
rect 5256 8128 5320 8132
rect 5336 8188 5400 8192
rect 5336 8132 5340 8188
rect 5340 8132 5396 8188
rect 5396 8132 5400 8188
rect 5336 8128 5400 8132
rect 5416 8188 5480 8192
rect 5416 8132 5420 8188
rect 5420 8132 5476 8188
rect 5476 8132 5480 8188
rect 5416 8128 5480 8132
rect 13624 8188 13688 8192
rect 13624 8132 13628 8188
rect 13628 8132 13684 8188
rect 13684 8132 13688 8188
rect 13624 8128 13688 8132
rect 13704 8188 13768 8192
rect 13704 8132 13708 8188
rect 13708 8132 13764 8188
rect 13764 8132 13768 8188
rect 13704 8128 13768 8132
rect 13784 8188 13848 8192
rect 13784 8132 13788 8188
rect 13788 8132 13844 8188
rect 13844 8132 13848 8188
rect 13784 8128 13848 8132
rect 13864 8188 13928 8192
rect 13864 8132 13868 8188
rect 13868 8132 13924 8188
rect 13924 8132 13928 8188
rect 13864 8128 13928 8132
rect 22072 8188 22136 8192
rect 22072 8132 22076 8188
rect 22076 8132 22132 8188
rect 22132 8132 22136 8188
rect 22072 8128 22136 8132
rect 22152 8188 22216 8192
rect 22152 8132 22156 8188
rect 22156 8132 22212 8188
rect 22212 8132 22216 8188
rect 22152 8128 22216 8132
rect 22232 8188 22296 8192
rect 22232 8132 22236 8188
rect 22236 8132 22292 8188
rect 22292 8132 22296 8188
rect 22232 8128 22296 8132
rect 22312 8188 22376 8192
rect 22312 8132 22316 8188
rect 22316 8132 22372 8188
rect 22372 8132 22376 8188
rect 22312 8128 22376 8132
rect 30520 8188 30584 8192
rect 30520 8132 30524 8188
rect 30524 8132 30580 8188
rect 30580 8132 30584 8188
rect 30520 8128 30584 8132
rect 30600 8188 30664 8192
rect 30600 8132 30604 8188
rect 30604 8132 30660 8188
rect 30660 8132 30664 8188
rect 30600 8128 30664 8132
rect 30680 8188 30744 8192
rect 30680 8132 30684 8188
rect 30684 8132 30740 8188
rect 30740 8132 30744 8188
rect 30680 8128 30744 8132
rect 30760 8188 30824 8192
rect 30760 8132 30764 8188
rect 30764 8132 30820 8188
rect 30820 8132 30824 8188
rect 30760 8128 30824 8132
rect 9400 7644 9464 7648
rect 9400 7588 9404 7644
rect 9404 7588 9460 7644
rect 9460 7588 9464 7644
rect 9400 7584 9464 7588
rect 9480 7644 9544 7648
rect 9480 7588 9484 7644
rect 9484 7588 9540 7644
rect 9540 7588 9544 7644
rect 9480 7584 9544 7588
rect 9560 7644 9624 7648
rect 9560 7588 9564 7644
rect 9564 7588 9620 7644
rect 9620 7588 9624 7644
rect 9560 7584 9624 7588
rect 9640 7644 9704 7648
rect 9640 7588 9644 7644
rect 9644 7588 9700 7644
rect 9700 7588 9704 7644
rect 9640 7584 9704 7588
rect 17848 7644 17912 7648
rect 17848 7588 17852 7644
rect 17852 7588 17908 7644
rect 17908 7588 17912 7644
rect 17848 7584 17912 7588
rect 17928 7644 17992 7648
rect 17928 7588 17932 7644
rect 17932 7588 17988 7644
rect 17988 7588 17992 7644
rect 17928 7584 17992 7588
rect 18008 7644 18072 7648
rect 18008 7588 18012 7644
rect 18012 7588 18068 7644
rect 18068 7588 18072 7644
rect 18008 7584 18072 7588
rect 18088 7644 18152 7648
rect 18088 7588 18092 7644
rect 18092 7588 18148 7644
rect 18148 7588 18152 7644
rect 18088 7584 18152 7588
rect 26296 7644 26360 7648
rect 26296 7588 26300 7644
rect 26300 7588 26356 7644
rect 26356 7588 26360 7644
rect 26296 7584 26360 7588
rect 26376 7644 26440 7648
rect 26376 7588 26380 7644
rect 26380 7588 26436 7644
rect 26436 7588 26440 7644
rect 26376 7584 26440 7588
rect 26456 7644 26520 7648
rect 26456 7588 26460 7644
rect 26460 7588 26516 7644
rect 26516 7588 26520 7644
rect 26456 7584 26520 7588
rect 26536 7644 26600 7648
rect 26536 7588 26540 7644
rect 26540 7588 26596 7644
rect 26596 7588 26600 7644
rect 26536 7584 26600 7588
rect 5176 7100 5240 7104
rect 5176 7044 5180 7100
rect 5180 7044 5236 7100
rect 5236 7044 5240 7100
rect 5176 7040 5240 7044
rect 5256 7100 5320 7104
rect 5256 7044 5260 7100
rect 5260 7044 5316 7100
rect 5316 7044 5320 7100
rect 5256 7040 5320 7044
rect 5336 7100 5400 7104
rect 5336 7044 5340 7100
rect 5340 7044 5396 7100
rect 5396 7044 5400 7100
rect 5336 7040 5400 7044
rect 5416 7100 5480 7104
rect 5416 7044 5420 7100
rect 5420 7044 5476 7100
rect 5476 7044 5480 7100
rect 5416 7040 5480 7044
rect 13624 7100 13688 7104
rect 13624 7044 13628 7100
rect 13628 7044 13684 7100
rect 13684 7044 13688 7100
rect 13624 7040 13688 7044
rect 13704 7100 13768 7104
rect 13704 7044 13708 7100
rect 13708 7044 13764 7100
rect 13764 7044 13768 7100
rect 13704 7040 13768 7044
rect 13784 7100 13848 7104
rect 13784 7044 13788 7100
rect 13788 7044 13844 7100
rect 13844 7044 13848 7100
rect 13784 7040 13848 7044
rect 13864 7100 13928 7104
rect 13864 7044 13868 7100
rect 13868 7044 13924 7100
rect 13924 7044 13928 7100
rect 13864 7040 13928 7044
rect 22072 7100 22136 7104
rect 22072 7044 22076 7100
rect 22076 7044 22132 7100
rect 22132 7044 22136 7100
rect 22072 7040 22136 7044
rect 22152 7100 22216 7104
rect 22152 7044 22156 7100
rect 22156 7044 22212 7100
rect 22212 7044 22216 7100
rect 22152 7040 22216 7044
rect 22232 7100 22296 7104
rect 22232 7044 22236 7100
rect 22236 7044 22292 7100
rect 22292 7044 22296 7100
rect 22232 7040 22296 7044
rect 22312 7100 22376 7104
rect 22312 7044 22316 7100
rect 22316 7044 22372 7100
rect 22372 7044 22376 7100
rect 22312 7040 22376 7044
rect 30520 7100 30584 7104
rect 30520 7044 30524 7100
rect 30524 7044 30580 7100
rect 30580 7044 30584 7100
rect 30520 7040 30584 7044
rect 30600 7100 30664 7104
rect 30600 7044 30604 7100
rect 30604 7044 30660 7100
rect 30660 7044 30664 7100
rect 30600 7040 30664 7044
rect 30680 7100 30744 7104
rect 30680 7044 30684 7100
rect 30684 7044 30740 7100
rect 30740 7044 30744 7100
rect 30680 7040 30744 7044
rect 30760 7100 30824 7104
rect 30760 7044 30764 7100
rect 30764 7044 30820 7100
rect 30820 7044 30824 7100
rect 30760 7040 30824 7044
rect 9400 6556 9464 6560
rect 9400 6500 9404 6556
rect 9404 6500 9460 6556
rect 9460 6500 9464 6556
rect 9400 6496 9464 6500
rect 9480 6556 9544 6560
rect 9480 6500 9484 6556
rect 9484 6500 9540 6556
rect 9540 6500 9544 6556
rect 9480 6496 9544 6500
rect 9560 6556 9624 6560
rect 9560 6500 9564 6556
rect 9564 6500 9620 6556
rect 9620 6500 9624 6556
rect 9560 6496 9624 6500
rect 9640 6556 9704 6560
rect 9640 6500 9644 6556
rect 9644 6500 9700 6556
rect 9700 6500 9704 6556
rect 9640 6496 9704 6500
rect 17848 6556 17912 6560
rect 17848 6500 17852 6556
rect 17852 6500 17908 6556
rect 17908 6500 17912 6556
rect 17848 6496 17912 6500
rect 17928 6556 17992 6560
rect 17928 6500 17932 6556
rect 17932 6500 17988 6556
rect 17988 6500 17992 6556
rect 17928 6496 17992 6500
rect 18008 6556 18072 6560
rect 18008 6500 18012 6556
rect 18012 6500 18068 6556
rect 18068 6500 18072 6556
rect 18008 6496 18072 6500
rect 18088 6556 18152 6560
rect 18088 6500 18092 6556
rect 18092 6500 18148 6556
rect 18148 6500 18152 6556
rect 18088 6496 18152 6500
rect 26296 6556 26360 6560
rect 26296 6500 26300 6556
rect 26300 6500 26356 6556
rect 26356 6500 26360 6556
rect 26296 6496 26360 6500
rect 26376 6556 26440 6560
rect 26376 6500 26380 6556
rect 26380 6500 26436 6556
rect 26436 6500 26440 6556
rect 26376 6496 26440 6500
rect 26456 6556 26520 6560
rect 26456 6500 26460 6556
rect 26460 6500 26516 6556
rect 26516 6500 26520 6556
rect 26456 6496 26520 6500
rect 26536 6556 26600 6560
rect 26536 6500 26540 6556
rect 26540 6500 26596 6556
rect 26596 6500 26600 6556
rect 26536 6496 26600 6500
rect 5176 6012 5240 6016
rect 5176 5956 5180 6012
rect 5180 5956 5236 6012
rect 5236 5956 5240 6012
rect 5176 5952 5240 5956
rect 5256 6012 5320 6016
rect 5256 5956 5260 6012
rect 5260 5956 5316 6012
rect 5316 5956 5320 6012
rect 5256 5952 5320 5956
rect 5336 6012 5400 6016
rect 5336 5956 5340 6012
rect 5340 5956 5396 6012
rect 5396 5956 5400 6012
rect 5336 5952 5400 5956
rect 5416 6012 5480 6016
rect 5416 5956 5420 6012
rect 5420 5956 5476 6012
rect 5476 5956 5480 6012
rect 5416 5952 5480 5956
rect 13624 6012 13688 6016
rect 13624 5956 13628 6012
rect 13628 5956 13684 6012
rect 13684 5956 13688 6012
rect 13624 5952 13688 5956
rect 13704 6012 13768 6016
rect 13704 5956 13708 6012
rect 13708 5956 13764 6012
rect 13764 5956 13768 6012
rect 13704 5952 13768 5956
rect 13784 6012 13848 6016
rect 13784 5956 13788 6012
rect 13788 5956 13844 6012
rect 13844 5956 13848 6012
rect 13784 5952 13848 5956
rect 13864 6012 13928 6016
rect 13864 5956 13868 6012
rect 13868 5956 13924 6012
rect 13924 5956 13928 6012
rect 13864 5952 13928 5956
rect 22072 6012 22136 6016
rect 22072 5956 22076 6012
rect 22076 5956 22132 6012
rect 22132 5956 22136 6012
rect 22072 5952 22136 5956
rect 22152 6012 22216 6016
rect 22152 5956 22156 6012
rect 22156 5956 22212 6012
rect 22212 5956 22216 6012
rect 22152 5952 22216 5956
rect 22232 6012 22296 6016
rect 22232 5956 22236 6012
rect 22236 5956 22292 6012
rect 22292 5956 22296 6012
rect 22232 5952 22296 5956
rect 22312 6012 22376 6016
rect 22312 5956 22316 6012
rect 22316 5956 22372 6012
rect 22372 5956 22376 6012
rect 22312 5952 22376 5956
rect 30520 6012 30584 6016
rect 30520 5956 30524 6012
rect 30524 5956 30580 6012
rect 30580 5956 30584 6012
rect 30520 5952 30584 5956
rect 30600 6012 30664 6016
rect 30600 5956 30604 6012
rect 30604 5956 30660 6012
rect 30660 5956 30664 6012
rect 30600 5952 30664 5956
rect 30680 6012 30744 6016
rect 30680 5956 30684 6012
rect 30684 5956 30740 6012
rect 30740 5956 30744 6012
rect 30680 5952 30744 5956
rect 30760 6012 30824 6016
rect 30760 5956 30764 6012
rect 30764 5956 30820 6012
rect 30820 5956 30824 6012
rect 30760 5952 30824 5956
rect 9400 5468 9464 5472
rect 9400 5412 9404 5468
rect 9404 5412 9460 5468
rect 9460 5412 9464 5468
rect 9400 5408 9464 5412
rect 9480 5468 9544 5472
rect 9480 5412 9484 5468
rect 9484 5412 9540 5468
rect 9540 5412 9544 5468
rect 9480 5408 9544 5412
rect 9560 5468 9624 5472
rect 9560 5412 9564 5468
rect 9564 5412 9620 5468
rect 9620 5412 9624 5468
rect 9560 5408 9624 5412
rect 9640 5468 9704 5472
rect 9640 5412 9644 5468
rect 9644 5412 9700 5468
rect 9700 5412 9704 5468
rect 9640 5408 9704 5412
rect 17848 5468 17912 5472
rect 17848 5412 17852 5468
rect 17852 5412 17908 5468
rect 17908 5412 17912 5468
rect 17848 5408 17912 5412
rect 17928 5468 17992 5472
rect 17928 5412 17932 5468
rect 17932 5412 17988 5468
rect 17988 5412 17992 5468
rect 17928 5408 17992 5412
rect 18008 5468 18072 5472
rect 18008 5412 18012 5468
rect 18012 5412 18068 5468
rect 18068 5412 18072 5468
rect 18008 5408 18072 5412
rect 18088 5468 18152 5472
rect 18088 5412 18092 5468
rect 18092 5412 18148 5468
rect 18148 5412 18152 5468
rect 18088 5408 18152 5412
rect 26296 5468 26360 5472
rect 26296 5412 26300 5468
rect 26300 5412 26356 5468
rect 26356 5412 26360 5468
rect 26296 5408 26360 5412
rect 26376 5468 26440 5472
rect 26376 5412 26380 5468
rect 26380 5412 26436 5468
rect 26436 5412 26440 5468
rect 26376 5408 26440 5412
rect 26456 5468 26520 5472
rect 26456 5412 26460 5468
rect 26460 5412 26516 5468
rect 26516 5412 26520 5468
rect 26456 5408 26520 5412
rect 26536 5468 26600 5472
rect 26536 5412 26540 5468
rect 26540 5412 26596 5468
rect 26596 5412 26600 5468
rect 26536 5408 26600 5412
rect 5176 4924 5240 4928
rect 5176 4868 5180 4924
rect 5180 4868 5236 4924
rect 5236 4868 5240 4924
rect 5176 4864 5240 4868
rect 5256 4924 5320 4928
rect 5256 4868 5260 4924
rect 5260 4868 5316 4924
rect 5316 4868 5320 4924
rect 5256 4864 5320 4868
rect 5336 4924 5400 4928
rect 5336 4868 5340 4924
rect 5340 4868 5396 4924
rect 5396 4868 5400 4924
rect 5336 4864 5400 4868
rect 5416 4924 5480 4928
rect 5416 4868 5420 4924
rect 5420 4868 5476 4924
rect 5476 4868 5480 4924
rect 5416 4864 5480 4868
rect 13624 4924 13688 4928
rect 13624 4868 13628 4924
rect 13628 4868 13684 4924
rect 13684 4868 13688 4924
rect 13624 4864 13688 4868
rect 13704 4924 13768 4928
rect 13704 4868 13708 4924
rect 13708 4868 13764 4924
rect 13764 4868 13768 4924
rect 13704 4864 13768 4868
rect 13784 4924 13848 4928
rect 13784 4868 13788 4924
rect 13788 4868 13844 4924
rect 13844 4868 13848 4924
rect 13784 4864 13848 4868
rect 13864 4924 13928 4928
rect 13864 4868 13868 4924
rect 13868 4868 13924 4924
rect 13924 4868 13928 4924
rect 13864 4864 13928 4868
rect 22072 4924 22136 4928
rect 22072 4868 22076 4924
rect 22076 4868 22132 4924
rect 22132 4868 22136 4924
rect 22072 4864 22136 4868
rect 22152 4924 22216 4928
rect 22152 4868 22156 4924
rect 22156 4868 22212 4924
rect 22212 4868 22216 4924
rect 22152 4864 22216 4868
rect 22232 4924 22296 4928
rect 22232 4868 22236 4924
rect 22236 4868 22292 4924
rect 22292 4868 22296 4924
rect 22232 4864 22296 4868
rect 22312 4924 22376 4928
rect 22312 4868 22316 4924
rect 22316 4868 22372 4924
rect 22372 4868 22376 4924
rect 22312 4864 22376 4868
rect 30520 4924 30584 4928
rect 30520 4868 30524 4924
rect 30524 4868 30580 4924
rect 30580 4868 30584 4924
rect 30520 4864 30584 4868
rect 30600 4924 30664 4928
rect 30600 4868 30604 4924
rect 30604 4868 30660 4924
rect 30660 4868 30664 4924
rect 30600 4864 30664 4868
rect 30680 4924 30744 4928
rect 30680 4868 30684 4924
rect 30684 4868 30740 4924
rect 30740 4868 30744 4924
rect 30680 4864 30744 4868
rect 30760 4924 30824 4928
rect 30760 4868 30764 4924
rect 30764 4868 30820 4924
rect 30820 4868 30824 4924
rect 30760 4864 30824 4868
rect 9400 4380 9464 4384
rect 9400 4324 9404 4380
rect 9404 4324 9460 4380
rect 9460 4324 9464 4380
rect 9400 4320 9464 4324
rect 9480 4380 9544 4384
rect 9480 4324 9484 4380
rect 9484 4324 9540 4380
rect 9540 4324 9544 4380
rect 9480 4320 9544 4324
rect 9560 4380 9624 4384
rect 9560 4324 9564 4380
rect 9564 4324 9620 4380
rect 9620 4324 9624 4380
rect 9560 4320 9624 4324
rect 9640 4380 9704 4384
rect 9640 4324 9644 4380
rect 9644 4324 9700 4380
rect 9700 4324 9704 4380
rect 9640 4320 9704 4324
rect 17848 4380 17912 4384
rect 17848 4324 17852 4380
rect 17852 4324 17908 4380
rect 17908 4324 17912 4380
rect 17848 4320 17912 4324
rect 17928 4380 17992 4384
rect 17928 4324 17932 4380
rect 17932 4324 17988 4380
rect 17988 4324 17992 4380
rect 17928 4320 17992 4324
rect 18008 4380 18072 4384
rect 18008 4324 18012 4380
rect 18012 4324 18068 4380
rect 18068 4324 18072 4380
rect 18008 4320 18072 4324
rect 18088 4380 18152 4384
rect 18088 4324 18092 4380
rect 18092 4324 18148 4380
rect 18148 4324 18152 4380
rect 18088 4320 18152 4324
rect 26296 4380 26360 4384
rect 26296 4324 26300 4380
rect 26300 4324 26356 4380
rect 26356 4324 26360 4380
rect 26296 4320 26360 4324
rect 26376 4380 26440 4384
rect 26376 4324 26380 4380
rect 26380 4324 26436 4380
rect 26436 4324 26440 4380
rect 26376 4320 26440 4324
rect 26456 4380 26520 4384
rect 26456 4324 26460 4380
rect 26460 4324 26516 4380
rect 26516 4324 26520 4380
rect 26456 4320 26520 4324
rect 26536 4380 26600 4384
rect 26536 4324 26540 4380
rect 26540 4324 26596 4380
rect 26596 4324 26600 4380
rect 26536 4320 26600 4324
rect 5176 3836 5240 3840
rect 5176 3780 5180 3836
rect 5180 3780 5236 3836
rect 5236 3780 5240 3836
rect 5176 3776 5240 3780
rect 5256 3836 5320 3840
rect 5256 3780 5260 3836
rect 5260 3780 5316 3836
rect 5316 3780 5320 3836
rect 5256 3776 5320 3780
rect 5336 3836 5400 3840
rect 5336 3780 5340 3836
rect 5340 3780 5396 3836
rect 5396 3780 5400 3836
rect 5336 3776 5400 3780
rect 5416 3836 5480 3840
rect 5416 3780 5420 3836
rect 5420 3780 5476 3836
rect 5476 3780 5480 3836
rect 5416 3776 5480 3780
rect 13624 3836 13688 3840
rect 13624 3780 13628 3836
rect 13628 3780 13684 3836
rect 13684 3780 13688 3836
rect 13624 3776 13688 3780
rect 13704 3836 13768 3840
rect 13704 3780 13708 3836
rect 13708 3780 13764 3836
rect 13764 3780 13768 3836
rect 13704 3776 13768 3780
rect 13784 3836 13848 3840
rect 13784 3780 13788 3836
rect 13788 3780 13844 3836
rect 13844 3780 13848 3836
rect 13784 3776 13848 3780
rect 13864 3836 13928 3840
rect 13864 3780 13868 3836
rect 13868 3780 13924 3836
rect 13924 3780 13928 3836
rect 13864 3776 13928 3780
rect 22072 3836 22136 3840
rect 22072 3780 22076 3836
rect 22076 3780 22132 3836
rect 22132 3780 22136 3836
rect 22072 3776 22136 3780
rect 22152 3836 22216 3840
rect 22152 3780 22156 3836
rect 22156 3780 22212 3836
rect 22212 3780 22216 3836
rect 22152 3776 22216 3780
rect 22232 3836 22296 3840
rect 22232 3780 22236 3836
rect 22236 3780 22292 3836
rect 22292 3780 22296 3836
rect 22232 3776 22296 3780
rect 22312 3836 22376 3840
rect 22312 3780 22316 3836
rect 22316 3780 22372 3836
rect 22372 3780 22376 3836
rect 22312 3776 22376 3780
rect 30520 3836 30584 3840
rect 30520 3780 30524 3836
rect 30524 3780 30580 3836
rect 30580 3780 30584 3836
rect 30520 3776 30584 3780
rect 30600 3836 30664 3840
rect 30600 3780 30604 3836
rect 30604 3780 30660 3836
rect 30660 3780 30664 3836
rect 30600 3776 30664 3780
rect 30680 3836 30744 3840
rect 30680 3780 30684 3836
rect 30684 3780 30740 3836
rect 30740 3780 30744 3836
rect 30680 3776 30744 3780
rect 30760 3836 30824 3840
rect 30760 3780 30764 3836
rect 30764 3780 30820 3836
rect 30820 3780 30824 3836
rect 30760 3776 30824 3780
rect 9400 3292 9464 3296
rect 9400 3236 9404 3292
rect 9404 3236 9460 3292
rect 9460 3236 9464 3292
rect 9400 3232 9464 3236
rect 9480 3292 9544 3296
rect 9480 3236 9484 3292
rect 9484 3236 9540 3292
rect 9540 3236 9544 3292
rect 9480 3232 9544 3236
rect 9560 3292 9624 3296
rect 9560 3236 9564 3292
rect 9564 3236 9620 3292
rect 9620 3236 9624 3292
rect 9560 3232 9624 3236
rect 9640 3292 9704 3296
rect 9640 3236 9644 3292
rect 9644 3236 9700 3292
rect 9700 3236 9704 3292
rect 9640 3232 9704 3236
rect 17848 3292 17912 3296
rect 17848 3236 17852 3292
rect 17852 3236 17908 3292
rect 17908 3236 17912 3292
rect 17848 3232 17912 3236
rect 17928 3292 17992 3296
rect 17928 3236 17932 3292
rect 17932 3236 17988 3292
rect 17988 3236 17992 3292
rect 17928 3232 17992 3236
rect 18008 3292 18072 3296
rect 18008 3236 18012 3292
rect 18012 3236 18068 3292
rect 18068 3236 18072 3292
rect 18008 3232 18072 3236
rect 18088 3292 18152 3296
rect 18088 3236 18092 3292
rect 18092 3236 18148 3292
rect 18148 3236 18152 3292
rect 18088 3232 18152 3236
rect 26296 3292 26360 3296
rect 26296 3236 26300 3292
rect 26300 3236 26356 3292
rect 26356 3236 26360 3292
rect 26296 3232 26360 3236
rect 26376 3292 26440 3296
rect 26376 3236 26380 3292
rect 26380 3236 26436 3292
rect 26436 3236 26440 3292
rect 26376 3232 26440 3236
rect 26456 3292 26520 3296
rect 26456 3236 26460 3292
rect 26460 3236 26516 3292
rect 26516 3236 26520 3292
rect 26456 3232 26520 3236
rect 26536 3292 26600 3296
rect 26536 3236 26540 3292
rect 26540 3236 26596 3292
rect 26596 3236 26600 3292
rect 26536 3232 26600 3236
rect 5176 2748 5240 2752
rect 5176 2692 5180 2748
rect 5180 2692 5236 2748
rect 5236 2692 5240 2748
rect 5176 2688 5240 2692
rect 5256 2748 5320 2752
rect 5256 2692 5260 2748
rect 5260 2692 5316 2748
rect 5316 2692 5320 2748
rect 5256 2688 5320 2692
rect 5336 2748 5400 2752
rect 5336 2692 5340 2748
rect 5340 2692 5396 2748
rect 5396 2692 5400 2748
rect 5336 2688 5400 2692
rect 5416 2748 5480 2752
rect 5416 2692 5420 2748
rect 5420 2692 5476 2748
rect 5476 2692 5480 2748
rect 5416 2688 5480 2692
rect 13624 2748 13688 2752
rect 13624 2692 13628 2748
rect 13628 2692 13684 2748
rect 13684 2692 13688 2748
rect 13624 2688 13688 2692
rect 13704 2748 13768 2752
rect 13704 2692 13708 2748
rect 13708 2692 13764 2748
rect 13764 2692 13768 2748
rect 13704 2688 13768 2692
rect 13784 2748 13848 2752
rect 13784 2692 13788 2748
rect 13788 2692 13844 2748
rect 13844 2692 13848 2748
rect 13784 2688 13848 2692
rect 13864 2748 13928 2752
rect 13864 2692 13868 2748
rect 13868 2692 13924 2748
rect 13924 2692 13928 2748
rect 13864 2688 13928 2692
rect 22072 2748 22136 2752
rect 22072 2692 22076 2748
rect 22076 2692 22132 2748
rect 22132 2692 22136 2748
rect 22072 2688 22136 2692
rect 22152 2748 22216 2752
rect 22152 2692 22156 2748
rect 22156 2692 22212 2748
rect 22212 2692 22216 2748
rect 22152 2688 22216 2692
rect 22232 2748 22296 2752
rect 22232 2692 22236 2748
rect 22236 2692 22292 2748
rect 22292 2692 22296 2748
rect 22232 2688 22296 2692
rect 22312 2748 22376 2752
rect 22312 2692 22316 2748
rect 22316 2692 22372 2748
rect 22372 2692 22376 2748
rect 22312 2688 22376 2692
rect 30520 2748 30584 2752
rect 30520 2692 30524 2748
rect 30524 2692 30580 2748
rect 30580 2692 30584 2748
rect 30520 2688 30584 2692
rect 30600 2748 30664 2752
rect 30600 2692 30604 2748
rect 30604 2692 30660 2748
rect 30660 2692 30664 2748
rect 30600 2688 30664 2692
rect 30680 2748 30744 2752
rect 30680 2692 30684 2748
rect 30684 2692 30740 2748
rect 30740 2692 30744 2748
rect 30680 2688 30744 2692
rect 30760 2748 30824 2752
rect 30760 2692 30764 2748
rect 30764 2692 30820 2748
rect 30820 2692 30824 2748
rect 30760 2688 30824 2692
rect 9400 2204 9464 2208
rect 9400 2148 9404 2204
rect 9404 2148 9460 2204
rect 9460 2148 9464 2204
rect 9400 2144 9464 2148
rect 9480 2204 9544 2208
rect 9480 2148 9484 2204
rect 9484 2148 9540 2204
rect 9540 2148 9544 2204
rect 9480 2144 9544 2148
rect 9560 2204 9624 2208
rect 9560 2148 9564 2204
rect 9564 2148 9620 2204
rect 9620 2148 9624 2204
rect 9560 2144 9624 2148
rect 9640 2204 9704 2208
rect 9640 2148 9644 2204
rect 9644 2148 9700 2204
rect 9700 2148 9704 2204
rect 9640 2144 9704 2148
rect 17848 2204 17912 2208
rect 17848 2148 17852 2204
rect 17852 2148 17908 2204
rect 17908 2148 17912 2204
rect 17848 2144 17912 2148
rect 17928 2204 17992 2208
rect 17928 2148 17932 2204
rect 17932 2148 17988 2204
rect 17988 2148 17992 2204
rect 17928 2144 17992 2148
rect 18008 2204 18072 2208
rect 18008 2148 18012 2204
rect 18012 2148 18068 2204
rect 18068 2148 18072 2204
rect 18008 2144 18072 2148
rect 18088 2204 18152 2208
rect 18088 2148 18092 2204
rect 18092 2148 18148 2204
rect 18148 2148 18152 2204
rect 18088 2144 18152 2148
rect 26296 2204 26360 2208
rect 26296 2148 26300 2204
rect 26300 2148 26356 2204
rect 26356 2148 26360 2204
rect 26296 2144 26360 2148
rect 26376 2204 26440 2208
rect 26376 2148 26380 2204
rect 26380 2148 26436 2204
rect 26436 2148 26440 2204
rect 26376 2144 26440 2148
rect 26456 2204 26520 2208
rect 26456 2148 26460 2204
rect 26460 2148 26516 2204
rect 26516 2148 26520 2204
rect 26456 2144 26520 2148
rect 26536 2204 26600 2208
rect 26536 2148 26540 2204
rect 26540 2148 26596 2204
rect 26596 2148 26600 2204
rect 26536 2144 26600 2148
<< metal4 >>
rect 5168 16896 5488 17456
rect 5168 16832 5176 16896
rect 5240 16832 5256 16896
rect 5320 16832 5336 16896
rect 5400 16832 5416 16896
rect 5480 16832 5488 16896
rect 5168 15808 5488 16832
rect 5168 15744 5176 15808
rect 5240 15744 5256 15808
rect 5320 15744 5336 15808
rect 5400 15744 5416 15808
rect 5480 15744 5488 15808
rect 5168 14720 5488 15744
rect 5168 14656 5176 14720
rect 5240 14656 5256 14720
rect 5320 14656 5336 14720
rect 5400 14656 5416 14720
rect 5480 14656 5488 14720
rect 5168 13632 5488 14656
rect 5168 13568 5176 13632
rect 5240 13568 5256 13632
rect 5320 13568 5336 13632
rect 5400 13568 5416 13632
rect 5480 13568 5488 13632
rect 5168 12544 5488 13568
rect 5168 12480 5176 12544
rect 5240 12480 5256 12544
rect 5320 12480 5336 12544
rect 5400 12480 5416 12544
rect 5480 12480 5488 12544
rect 5168 11456 5488 12480
rect 5168 11392 5176 11456
rect 5240 11392 5256 11456
rect 5320 11392 5336 11456
rect 5400 11392 5416 11456
rect 5480 11392 5488 11456
rect 5168 10368 5488 11392
rect 5168 10304 5176 10368
rect 5240 10304 5256 10368
rect 5320 10304 5336 10368
rect 5400 10304 5416 10368
rect 5480 10304 5488 10368
rect 5168 9280 5488 10304
rect 5168 9216 5176 9280
rect 5240 9216 5256 9280
rect 5320 9216 5336 9280
rect 5400 9216 5416 9280
rect 5480 9216 5488 9280
rect 5168 8192 5488 9216
rect 5168 8128 5176 8192
rect 5240 8128 5256 8192
rect 5320 8128 5336 8192
rect 5400 8128 5416 8192
rect 5480 8128 5488 8192
rect 5168 7104 5488 8128
rect 5168 7040 5176 7104
rect 5240 7040 5256 7104
rect 5320 7040 5336 7104
rect 5400 7040 5416 7104
rect 5480 7040 5488 7104
rect 5168 6016 5488 7040
rect 5168 5952 5176 6016
rect 5240 5952 5256 6016
rect 5320 5952 5336 6016
rect 5400 5952 5416 6016
rect 5480 5952 5488 6016
rect 5168 4928 5488 5952
rect 5168 4864 5176 4928
rect 5240 4864 5256 4928
rect 5320 4864 5336 4928
rect 5400 4864 5416 4928
rect 5480 4864 5488 4928
rect 5168 3840 5488 4864
rect 5168 3776 5176 3840
rect 5240 3776 5256 3840
rect 5320 3776 5336 3840
rect 5400 3776 5416 3840
rect 5480 3776 5488 3840
rect 5168 2752 5488 3776
rect 5168 2688 5176 2752
rect 5240 2688 5256 2752
rect 5320 2688 5336 2752
rect 5400 2688 5416 2752
rect 5480 2688 5488 2752
rect 5168 2128 5488 2688
rect 9392 17440 9712 17456
rect 9392 17376 9400 17440
rect 9464 17376 9480 17440
rect 9544 17376 9560 17440
rect 9624 17376 9640 17440
rect 9704 17376 9712 17440
rect 9392 16352 9712 17376
rect 9392 16288 9400 16352
rect 9464 16288 9480 16352
rect 9544 16288 9560 16352
rect 9624 16288 9640 16352
rect 9704 16288 9712 16352
rect 9392 15264 9712 16288
rect 9392 15200 9400 15264
rect 9464 15200 9480 15264
rect 9544 15200 9560 15264
rect 9624 15200 9640 15264
rect 9704 15200 9712 15264
rect 9392 14176 9712 15200
rect 9392 14112 9400 14176
rect 9464 14112 9480 14176
rect 9544 14112 9560 14176
rect 9624 14112 9640 14176
rect 9704 14112 9712 14176
rect 9392 13088 9712 14112
rect 9392 13024 9400 13088
rect 9464 13024 9480 13088
rect 9544 13024 9560 13088
rect 9624 13024 9640 13088
rect 9704 13024 9712 13088
rect 9392 12000 9712 13024
rect 9392 11936 9400 12000
rect 9464 11936 9480 12000
rect 9544 11936 9560 12000
rect 9624 11936 9640 12000
rect 9704 11936 9712 12000
rect 9392 10912 9712 11936
rect 9392 10848 9400 10912
rect 9464 10848 9480 10912
rect 9544 10848 9560 10912
rect 9624 10848 9640 10912
rect 9704 10848 9712 10912
rect 9392 9824 9712 10848
rect 9392 9760 9400 9824
rect 9464 9760 9480 9824
rect 9544 9760 9560 9824
rect 9624 9760 9640 9824
rect 9704 9760 9712 9824
rect 9392 8736 9712 9760
rect 9392 8672 9400 8736
rect 9464 8672 9480 8736
rect 9544 8672 9560 8736
rect 9624 8672 9640 8736
rect 9704 8672 9712 8736
rect 9392 7648 9712 8672
rect 9392 7584 9400 7648
rect 9464 7584 9480 7648
rect 9544 7584 9560 7648
rect 9624 7584 9640 7648
rect 9704 7584 9712 7648
rect 9392 6560 9712 7584
rect 9392 6496 9400 6560
rect 9464 6496 9480 6560
rect 9544 6496 9560 6560
rect 9624 6496 9640 6560
rect 9704 6496 9712 6560
rect 9392 5472 9712 6496
rect 9392 5408 9400 5472
rect 9464 5408 9480 5472
rect 9544 5408 9560 5472
rect 9624 5408 9640 5472
rect 9704 5408 9712 5472
rect 9392 4384 9712 5408
rect 9392 4320 9400 4384
rect 9464 4320 9480 4384
rect 9544 4320 9560 4384
rect 9624 4320 9640 4384
rect 9704 4320 9712 4384
rect 9392 3296 9712 4320
rect 9392 3232 9400 3296
rect 9464 3232 9480 3296
rect 9544 3232 9560 3296
rect 9624 3232 9640 3296
rect 9704 3232 9712 3296
rect 9392 2208 9712 3232
rect 9392 2144 9400 2208
rect 9464 2144 9480 2208
rect 9544 2144 9560 2208
rect 9624 2144 9640 2208
rect 9704 2144 9712 2208
rect 9392 2128 9712 2144
rect 13616 16896 13936 17456
rect 13616 16832 13624 16896
rect 13688 16832 13704 16896
rect 13768 16832 13784 16896
rect 13848 16832 13864 16896
rect 13928 16832 13936 16896
rect 13616 15808 13936 16832
rect 13616 15744 13624 15808
rect 13688 15744 13704 15808
rect 13768 15744 13784 15808
rect 13848 15744 13864 15808
rect 13928 15744 13936 15808
rect 13616 14720 13936 15744
rect 13616 14656 13624 14720
rect 13688 14656 13704 14720
rect 13768 14656 13784 14720
rect 13848 14656 13864 14720
rect 13928 14656 13936 14720
rect 13616 13632 13936 14656
rect 13616 13568 13624 13632
rect 13688 13568 13704 13632
rect 13768 13568 13784 13632
rect 13848 13568 13864 13632
rect 13928 13568 13936 13632
rect 13616 12544 13936 13568
rect 13616 12480 13624 12544
rect 13688 12480 13704 12544
rect 13768 12480 13784 12544
rect 13848 12480 13864 12544
rect 13928 12480 13936 12544
rect 13616 11456 13936 12480
rect 13616 11392 13624 11456
rect 13688 11392 13704 11456
rect 13768 11392 13784 11456
rect 13848 11392 13864 11456
rect 13928 11392 13936 11456
rect 13616 10368 13936 11392
rect 13616 10304 13624 10368
rect 13688 10304 13704 10368
rect 13768 10304 13784 10368
rect 13848 10304 13864 10368
rect 13928 10304 13936 10368
rect 13616 9280 13936 10304
rect 13616 9216 13624 9280
rect 13688 9216 13704 9280
rect 13768 9216 13784 9280
rect 13848 9216 13864 9280
rect 13928 9216 13936 9280
rect 13616 8192 13936 9216
rect 13616 8128 13624 8192
rect 13688 8128 13704 8192
rect 13768 8128 13784 8192
rect 13848 8128 13864 8192
rect 13928 8128 13936 8192
rect 13616 7104 13936 8128
rect 13616 7040 13624 7104
rect 13688 7040 13704 7104
rect 13768 7040 13784 7104
rect 13848 7040 13864 7104
rect 13928 7040 13936 7104
rect 13616 6016 13936 7040
rect 13616 5952 13624 6016
rect 13688 5952 13704 6016
rect 13768 5952 13784 6016
rect 13848 5952 13864 6016
rect 13928 5952 13936 6016
rect 13616 4928 13936 5952
rect 13616 4864 13624 4928
rect 13688 4864 13704 4928
rect 13768 4864 13784 4928
rect 13848 4864 13864 4928
rect 13928 4864 13936 4928
rect 13616 3840 13936 4864
rect 13616 3776 13624 3840
rect 13688 3776 13704 3840
rect 13768 3776 13784 3840
rect 13848 3776 13864 3840
rect 13928 3776 13936 3840
rect 13616 2752 13936 3776
rect 13616 2688 13624 2752
rect 13688 2688 13704 2752
rect 13768 2688 13784 2752
rect 13848 2688 13864 2752
rect 13928 2688 13936 2752
rect 13616 2128 13936 2688
rect 17840 17440 18160 17456
rect 17840 17376 17848 17440
rect 17912 17376 17928 17440
rect 17992 17376 18008 17440
rect 18072 17376 18088 17440
rect 18152 17376 18160 17440
rect 17840 16352 18160 17376
rect 17840 16288 17848 16352
rect 17912 16288 17928 16352
rect 17992 16288 18008 16352
rect 18072 16288 18088 16352
rect 18152 16288 18160 16352
rect 17840 15264 18160 16288
rect 17840 15200 17848 15264
rect 17912 15200 17928 15264
rect 17992 15200 18008 15264
rect 18072 15200 18088 15264
rect 18152 15200 18160 15264
rect 17840 14176 18160 15200
rect 17840 14112 17848 14176
rect 17912 14112 17928 14176
rect 17992 14112 18008 14176
rect 18072 14112 18088 14176
rect 18152 14112 18160 14176
rect 17840 13088 18160 14112
rect 17840 13024 17848 13088
rect 17912 13024 17928 13088
rect 17992 13024 18008 13088
rect 18072 13024 18088 13088
rect 18152 13024 18160 13088
rect 17840 12000 18160 13024
rect 17840 11936 17848 12000
rect 17912 11936 17928 12000
rect 17992 11936 18008 12000
rect 18072 11936 18088 12000
rect 18152 11936 18160 12000
rect 17840 10912 18160 11936
rect 17840 10848 17848 10912
rect 17912 10848 17928 10912
rect 17992 10848 18008 10912
rect 18072 10848 18088 10912
rect 18152 10848 18160 10912
rect 17840 9824 18160 10848
rect 17840 9760 17848 9824
rect 17912 9760 17928 9824
rect 17992 9760 18008 9824
rect 18072 9760 18088 9824
rect 18152 9760 18160 9824
rect 17840 8736 18160 9760
rect 17840 8672 17848 8736
rect 17912 8672 17928 8736
rect 17992 8672 18008 8736
rect 18072 8672 18088 8736
rect 18152 8672 18160 8736
rect 17840 7648 18160 8672
rect 17840 7584 17848 7648
rect 17912 7584 17928 7648
rect 17992 7584 18008 7648
rect 18072 7584 18088 7648
rect 18152 7584 18160 7648
rect 17840 6560 18160 7584
rect 17840 6496 17848 6560
rect 17912 6496 17928 6560
rect 17992 6496 18008 6560
rect 18072 6496 18088 6560
rect 18152 6496 18160 6560
rect 17840 5472 18160 6496
rect 17840 5408 17848 5472
rect 17912 5408 17928 5472
rect 17992 5408 18008 5472
rect 18072 5408 18088 5472
rect 18152 5408 18160 5472
rect 17840 4384 18160 5408
rect 17840 4320 17848 4384
rect 17912 4320 17928 4384
rect 17992 4320 18008 4384
rect 18072 4320 18088 4384
rect 18152 4320 18160 4384
rect 17840 3296 18160 4320
rect 17840 3232 17848 3296
rect 17912 3232 17928 3296
rect 17992 3232 18008 3296
rect 18072 3232 18088 3296
rect 18152 3232 18160 3296
rect 17840 2208 18160 3232
rect 17840 2144 17848 2208
rect 17912 2144 17928 2208
rect 17992 2144 18008 2208
rect 18072 2144 18088 2208
rect 18152 2144 18160 2208
rect 17840 2128 18160 2144
rect 22064 16896 22384 17456
rect 22064 16832 22072 16896
rect 22136 16832 22152 16896
rect 22216 16832 22232 16896
rect 22296 16832 22312 16896
rect 22376 16832 22384 16896
rect 22064 15808 22384 16832
rect 22064 15744 22072 15808
rect 22136 15744 22152 15808
rect 22216 15744 22232 15808
rect 22296 15744 22312 15808
rect 22376 15744 22384 15808
rect 22064 14720 22384 15744
rect 22064 14656 22072 14720
rect 22136 14656 22152 14720
rect 22216 14656 22232 14720
rect 22296 14656 22312 14720
rect 22376 14656 22384 14720
rect 22064 13632 22384 14656
rect 22064 13568 22072 13632
rect 22136 13568 22152 13632
rect 22216 13568 22232 13632
rect 22296 13568 22312 13632
rect 22376 13568 22384 13632
rect 22064 12544 22384 13568
rect 22064 12480 22072 12544
rect 22136 12480 22152 12544
rect 22216 12480 22232 12544
rect 22296 12480 22312 12544
rect 22376 12480 22384 12544
rect 22064 11456 22384 12480
rect 22064 11392 22072 11456
rect 22136 11392 22152 11456
rect 22216 11392 22232 11456
rect 22296 11392 22312 11456
rect 22376 11392 22384 11456
rect 22064 10368 22384 11392
rect 22064 10304 22072 10368
rect 22136 10304 22152 10368
rect 22216 10304 22232 10368
rect 22296 10304 22312 10368
rect 22376 10304 22384 10368
rect 22064 9280 22384 10304
rect 22064 9216 22072 9280
rect 22136 9216 22152 9280
rect 22216 9216 22232 9280
rect 22296 9216 22312 9280
rect 22376 9216 22384 9280
rect 22064 8192 22384 9216
rect 22064 8128 22072 8192
rect 22136 8128 22152 8192
rect 22216 8128 22232 8192
rect 22296 8128 22312 8192
rect 22376 8128 22384 8192
rect 22064 7104 22384 8128
rect 22064 7040 22072 7104
rect 22136 7040 22152 7104
rect 22216 7040 22232 7104
rect 22296 7040 22312 7104
rect 22376 7040 22384 7104
rect 22064 6016 22384 7040
rect 22064 5952 22072 6016
rect 22136 5952 22152 6016
rect 22216 5952 22232 6016
rect 22296 5952 22312 6016
rect 22376 5952 22384 6016
rect 22064 4928 22384 5952
rect 22064 4864 22072 4928
rect 22136 4864 22152 4928
rect 22216 4864 22232 4928
rect 22296 4864 22312 4928
rect 22376 4864 22384 4928
rect 22064 3840 22384 4864
rect 22064 3776 22072 3840
rect 22136 3776 22152 3840
rect 22216 3776 22232 3840
rect 22296 3776 22312 3840
rect 22376 3776 22384 3840
rect 22064 2752 22384 3776
rect 22064 2688 22072 2752
rect 22136 2688 22152 2752
rect 22216 2688 22232 2752
rect 22296 2688 22312 2752
rect 22376 2688 22384 2752
rect 22064 2128 22384 2688
rect 26288 17440 26608 17456
rect 26288 17376 26296 17440
rect 26360 17376 26376 17440
rect 26440 17376 26456 17440
rect 26520 17376 26536 17440
rect 26600 17376 26608 17440
rect 26288 16352 26608 17376
rect 26288 16288 26296 16352
rect 26360 16288 26376 16352
rect 26440 16288 26456 16352
rect 26520 16288 26536 16352
rect 26600 16288 26608 16352
rect 26288 15264 26608 16288
rect 26288 15200 26296 15264
rect 26360 15200 26376 15264
rect 26440 15200 26456 15264
rect 26520 15200 26536 15264
rect 26600 15200 26608 15264
rect 26288 14176 26608 15200
rect 26288 14112 26296 14176
rect 26360 14112 26376 14176
rect 26440 14112 26456 14176
rect 26520 14112 26536 14176
rect 26600 14112 26608 14176
rect 26288 13088 26608 14112
rect 26288 13024 26296 13088
rect 26360 13024 26376 13088
rect 26440 13024 26456 13088
rect 26520 13024 26536 13088
rect 26600 13024 26608 13088
rect 26288 12000 26608 13024
rect 26288 11936 26296 12000
rect 26360 11936 26376 12000
rect 26440 11936 26456 12000
rect 26520 11936 26536 12000
rect 26600 11936 26608 12000
rect 26288 10912 26608 11936
rect 26288 10848 26296 10912
rect 26360 10848 26376 10912
rect 26440 10848 26456 10912
rect 26520 10848 26536 10912
rect 26600 10848 26608 10912
rect 26288 9824 26608 10848
rect 26288 9760 26296 9824
rect 26360 9760 26376 9824
rect 26440 9760 26456 9824
rect 26520 9760 26536 9824
rect 26600 9760 26608 9824
rect 26288 8736 26608 9760
rect 26288 8672 26296 8736
rect 26360 8672 26376 8736
rect 26440 8672 26456 8736
rect 26520 8672 26536 8736
rect 26600 8672 26608 8736
rect 26288 7648 26608 8672
rect 26288 7584 26296 7648
rect 26360 7584 26376 7648
rect 26440 7584 26456 7648
rect 26520 7584 26536 7648
rect 26600 7584 26608 7648
rect 26288 6560 26608 7584
rect 26288 6496 26296 6560
rect 26360 6496 26376 6560
rect 26440 6496 26456 6560
rect 26520 6496 26536 6560
rect 26600 6496 26608 6560
rect 26288 5472 26608 6496
rect 26288 5408 26296 5472
rect 26360 5408 26376 5472
rect 26440 5408 26456 5472
rect 26520 5408 26536 5472
rect 26600 5408 26608 5472
rect 26288 4384 26608 5408
rect 26288 4320 26296 4384
rect 26360 4320 26376 4384
rect 26440 4320 26456 4384
rect 26520 4320 26536 4384
rect 26600 4320 26608 4384
rect 26288 3296 26608 4320
rect 26288 3232 26296 3296
rect 26360 3232 26376 3296
rect 26440 3232 26456 3296
rect 26520 3232 26536 3296
rect 26600 3232 26608 3296
rect 26288 2208 26608 3232
rect 26288 2144 26296 2208
rect 26360 2144 26376 2208
rect 26440 2144 26456 2208
rect 26520 2144 26536 2208
rect 26600 2144 26608 2208
rect 26288 2128 26608 2144
rect 30512 16896 30832 17456
rect 30512 16832 30520 16896
rect 30584 16832 30600 16896
rect 30664 16832 30680 16896
rect 30744 16832 30760 16896
rect 30824 16832 30832 16896
rect 30512 15808 30832 16832
rect 30512 15744 30520 15808
rect 30584 15744 30600 15808
rect 30664 15744 30680 15808
rect 30744 15744 30760 15808
rect 30824 15744 30832 15808
rect 30512 14720 30832 15744
rect 30512 14656 30520 14720
rect 30584 14656 30600 14720
rect 30664 14656 30680 14720
rect 30744 14656 30760 14720
rect 30824 14656 30832 14720
rect 30512 13632 30832 14656
rect 30512 13568 30520 13632
rect 30584 13568 30600 13632
rect 30664 13568 30680 13632
rect 30744 13568 30760 13632
rect 30824 13568 30832 13632
rect 30512 12544 30832 13568
rect 30512 12480 30520 12544
rect 30584 12480 30600 12544
rect 30664 12480 30680 12544
rect 30744 12480 30760 12544
rect 30824 12480 30832 12544
rect 30512 11456 30832 12480
rect 30512 11392 30520 11456
rect 30584 11392 30600 11456
rect 30664 11392 30680 11456
rect 30744 11392 30760 11456
rect 30824 11392 30832 11456
rect 30512 10368 30832 11392
rect 30512 10304 30520 10368
rect 30584 10304 30600 10368
rect 30664 10304 30680 10368
rect 30744 10304 30760 10368
rect 30824 10304 30832 10368
rect 30512 9280 30832 10304
rect 30512 9216 30520 9280
rect 30584 9216 30600 9280
rect 30664 9216 30680 9280
rect 30744 9216 30760 9280
rect 30824 9216 30832 9280
rect 30512 8192 30832 9216
rect 30512 8128 30520 8192
rect 30584 8128 30600 8192
rect 30664 8128 30680 8192
rect 30744 8128 30760 8192
rect 30824 8128 30832 8192
rect 30512 7104 30832 8128
rect 30512 7040 30520 7104
rect 30584 7040 30600 7104
rect 30664 7040 30680 7104
rect 30744 7040 30760 7104
rect 30824 7040 30832 7104
rect 30512 6016 30832 7040
rect 30512 5952 30520 6016
rect 30584 5952 30600 6016
rect 30664 5952 30680 6016
rect 30744 5952 30760 6016
rect 30824 5952 30832 6016
rect 30512 4928 30832 5952
rect 30512 4864 30520 4928
rect 30584 4864 30600 4928
rect 30664 4864 30680 4928
rect 30744 4864 30760 4928
rect 30824 4864 30832 4928
rect 30512 3840 30832 4864
rect 30512 3776 30520 3840
rect 30584 3776 30600 3840
rect 30664 3776 30680 3840
rect 30744 3776 30760 3840
rect 30824 3776 30832 3840
rect 30512 2752 30832 3776
rect 30512 2688 30520 2752
rect 30584 2688 30600 2752
rect 30664 2688 30680 2752
rect 30744 2688 30760 2752
rect 30824 2688 30832 2752
rect 30512 2128 30832 2688
use sky130_fd_sc_hd__diode_2  ANTENNA__073__S dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 26312 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__075__S
timestamp 1649977179
transform 1 0 30452 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__077__S
timestamp 1649977179
transform 1 0 30452 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__081__A
timestamp 1649977179
transform 1 0 5704 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__081__B_N
timestamp 1649977179
transform 1 0 5980 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__082__A1
timestamp 1649977179
transform 1 0 20148 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__082__S
timestamp 1649977179
transform -1 0 20700 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__084__A0
timestamp 1649977179
transform 1 0 7176 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__084__S
timestamp 1649977179
transform 1 0 6808 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__086__S
timestamp 1649977179
transform 1 0 7268 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__088__A
timestamp 1649977179
transform 1 0 21804 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__088__B
timestamp 1649977179
transform -1 0 20884 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__088__C_N
timestamp 1649977179
transform 1 0 20148 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__089__A0
timestamp 1649977179
transform 1 0 21804 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__133__A
timestamp 1649977179
transform 1 0 3864 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__134__A
timestamp 1649977179
transform 1 0 5152 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__135__A
timestamp 1649977179
transform 1 0 4876 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__136__A
timestamp 1649977179
transform 1 0 13248 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__137__A
timestamp 1649977179
transform 1 0 5520 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__138__A
timestamp 1649977179
transform -1 0 22448 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__139__A
timestamp 1649977179
transform 1 0 5980 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__145__A
timestamp 1649977179
transform -1 0 29256 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__146__A
timestamp 1649977179
transform 1 0 27876 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__147__A
timestamp 1649977179
transform 1 0 28060 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__150__CLK
timestamp 1649977179
transform -1 0 5888 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__151__CLK
timestamp 1649977179
transform 1 0 5428 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__152__CLK
timestamp 1649977179
transform 1 0 11132 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__153__CLK
timestamp 1649977179
transform 1 0 6348 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__156__CLK
timestamp 1649977179
transform 1 0 13432 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__157__CLK
timestamp 1649977179
transform 1 0 8924 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__158__CLK
timestamp 1649977179
transform 1 0 6348 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__159__CLK
timestamp 1649977179
transform 1 0 12788 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_clk_A
timestamp 1649977179
transform -1 0 15548 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input1_A
timestamp 1649977179
transform -1 0 1564 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input2_A
timestamp 1649977179
transform -1 0 1564 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input3_A
timestamp 1649977179
transform -1 0 1564 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input4_A
timestamp 1649977179
transform -1 0 10120 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input5_A
timestamp 1649977179
transform -1 0 5152 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input6_A
timestamp 1649977179
transform -1 0 7636 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input7_A
timestamp 1649977179
transform -1 0 1840 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output12_A
timestamp 1649977179
transform 1 0 30268 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output18_A
timestamp 1649977179
transform 1 0 33304 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 1380 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 1748 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 2208 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24
timestamp 1649977179
transform 1 0 3312 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 3772 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38
timestamp 1649977179
transform 1 0 4600 0 1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44
timestamp 1649977179
transform 1 0 5152 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_57
timestamp 1649977179
transform 1 0 6348 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61
timestamp 1649977179
transform 1 0 6716 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_65
timestamp 1649977179
transform 1 0 7084 0 1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71
timestamp 1649977179
transform 1 0 7636 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_83
timestamp 1649977179
transform 1 0 8740 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_85
timestamp 1649977179
transform 1 0 8924 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_92
timestamp 1649977179
transform 1 0 9568 0 1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98
timestamp 1649977179
transform 1 0 10120 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_110 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 11224 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113
timestamp 1649977179
transform 1 0 11500 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_125
timestamp 1649977179
transform 1 0 12604 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_137 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 13708 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_141
timestamp 1649977179
transform 1 0 14076 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_147
timestamp 1649977179
transform 1 0 14628 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_159 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 15732 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_167
timestamp 1649977179
transform 1 0 16468 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_169
timestamp 1649977179
transform 1 0 16652 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_181
timestamp 1649977179
transform 1 0 17756 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_193
timestamp 1649977179
transform 1 0 18860 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_197
timestamp 1649977179
transform 1 0 19228 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_209
timestamp 1649977179
transform 1 0 20332 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_221
timestamp 1649977179
transform 1 0 21436 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_229
timestamp 1649977179
transform 1 0 22172 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_241
timestamp 1649977179
transform 1 0 23276 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_249
timestamp 1649977179
transform 1 0 24012 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_253
timestamp 1649977179
transform 1 0 24380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_265
timestamp 1649977179
transform 1 0 25484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_277
timestamp 1649977179
transform 1 0 26588 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_281
timestamp 1649977179
transform 1 0 26956 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_293
timestamp 1649977179
transform 1 0 28060 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_305
timestamp 1649977179
transform 1 0 29164 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_313
timestamp 1649977179
transform 1 0 29900 0 1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_319
timestamp 1649977179
transform 1 0 30452 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_331
timestamp 1649977179
transform 1 0 31556 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_335
timestamp 1649977179
transform 1 0 31924 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_337
timestamp 1649977179
transform 1 0 32108 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_352
timestamp 1649977179
transform 1 0 33488 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_360
timestamp 1649977179
transform 1 0 34224 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_1_3
timestamp 1649977179
transform 1 0 1380 0 -1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_1_8
timestamp 1649977179
transform 1 0 1840 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_20
timestamp 1649977179
transform 1 0 2944 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_32
timestamp 1649977179
transform 1 0 4048 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_44
timestamp 1649977179
transform 1 0 5152 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_57
timestamp 1649977179
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_69
timestamp 1649977179
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_81
timestamp 1649977179
transform 1 0 8556 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_93
timestamp 1649977179
transform 1 0 9660 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_105
timestamp 1649977179
transform 1 0 10764 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_111
timestamp 1649977179
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_1_113
timestamp 1649977179
transform 1 0 11500 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_119
timestamp 1649977179
transform 1 0 12052 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_125
timestamp 1649977179
transform 1 0 12604 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_137
timestamp 1649977179
transform 1 0 13708 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_149
timestamp 1649977179
transform 1 0 14812 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_161
timestamp 1649977179
transform 1 0 15916 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_167
timestamp 1649977179
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_169
timestamp 1649977179
transform 1 0 16652 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_181
timestamp 1649977179
transform 1 0 17756 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_193
timestamp 1649977179
transform 1 0 18860 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_205
timestamp 1649977179
transform 1 0 19964 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_217
timestamp 1649977179
transform 1 0 21068 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_223
timestamp 1649977179
transform 1 0 21620 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_225
timestamp 1649977179
transform 1 0 21804 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_1_237
timestamp 1649977179
transform 1 0 22908 0 -1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_1_247
timestamp 1649977179
transform 1 0 23828 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_259
timestamp 1649977179
transform 1 0 24932 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_271
timestamp 1649977179
transform 1 0 26036 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_279
timestamp 1649977179
transform 1 0 26772 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_281
timestamp 1649977179
transform 1 0 26956 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_293
timestamp 1649977179
transform 1 0 28060 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_305
timestamp 1649977179
transform 1 0 29164 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_317
timestamp 1649977179
transform 1 0 30268 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_321
timestamp 1649977179
transform 1 0 30636 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_325
timestamp 1649977179
transform 1 0 31004 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_1_333
timestamp 1649977179
transform 1 0 31740 0 -1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_1_337
timestamp 1649977179
transform 1 0 32108 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_349
timestamp 1649977179
transform 1 0 33212 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_1_361
timestamp 1649977179
transform 1 0 34316 0 -1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3
timestamp 1649977179
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_15
timestamp 1649977179
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp 1649977179
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_29
timestamp 1649977179
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_41
timestamp 1649977179
transform 1 0 4876 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_49
timestamp 1649977179
transform 1 0 5612 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_61
timestamp 1649977179
transform 1 0 6716 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_73
timestamp 1649977179
transform 1 0 7820 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_2_81
timestamp 1649977179
transform 1 0 8556 0 1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_2_85
timestamp 1649977179
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_97
timestamp 1649977179
transform 1 0 10028 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_109
timestamp 1649977179
transform 1 0 11132 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_121
timestamp 1649977179
transform 1 0 12236 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_129
timestamp 1649977179
transform 1 0 12972 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_2_137
timestamp 1649977179
transform 1 0 13708 0 1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_2_141
timestamp 1649977179
transform 1 0 14076 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_153
timestamp 1649977179
transform 1 0 15180 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_165
timestamp 1649977179
transform 1 0 16284 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_177
timestamp 1649977179
transform 1 0 17388 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_189
timestamp 1649977179
transform 1 0 18492 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_195
timestamp 1649977179
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_197
timestamp 1649977179
transform 1 0 19228 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_209
timestamp 1649977179
transform 1 0 20332 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_2_221
timestamp 1649977179
transform 1 0 21436 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_2_227
timestamp 1649977179
transform 1 0 21988 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_238
timestamp 1649977179
transform 1 0 23000 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_244
timestamp 1649977179
transform 1 0 23552 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_248
timestamp 1649977179
transform 1 0 23920 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_2_258
timestamp 1649977179
transform 1 0 24840 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_270
timestamp 1649977179
transform 1 0 25944 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_282
timestamp 1649977179
transform 1 0 27048 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_294
timestamp 1649977179
transform 1 0 28152 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_301
timestamp 1649977179
transform 1 0 28796 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_307
timestamp 1649977179
transform 1 0 29348 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_309
timestamp 1649977179
transform 1 0 29532 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_322
timestamp 1649977179
transform 1 0 30728 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_326
timestamp 1649977179
transform 1 0 31096 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_333
timestamp 1649977179
transform 1 0 31740 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_345
timestamp 1649977179
transform 1 0 32844 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_357
timestamp 1649977179
transform 1 0 33948 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_363
timestamp 1649977179
transform 1 0 34500 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3
timestamp 1649977179
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_15
timestamp 1649977179
transform 1 0 2484 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_3_23
timestamp 1649977179
transform 1 0 3220 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_46
timestamp 1649977179
transform 1 0 5336 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_52
timestamp 1649977179
transform 1 0 5888 0 -1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_3_57
timestamp 1649977179
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_69
timestamp 1649977179
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_81
timestamp 1649977179
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_93
timestamp 1649977179
transform 1 0 9660 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_105
timestamp 1649977179
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_111
timestamp 1649977179
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_116
timestamp 1649977179
transform 1 0 11776 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_132
timestamp 1649977179
transform 1 0 13248 0 -1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_3_139
timestamp 1649977179
transform 1 0 13892 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_151
timestamp 1649977179
transform 1 0 14996 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_161
timestamp 1649977179
transform 1 0 15916 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_167
timestamp 1649977179
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_169
timestamp 1649977179
transform 1 0 16652 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_181
timestamp 1649977179
transform 1 0 17756 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_193
timestamp 1649977179
transform 1 0 18860 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_205
timestamp 1649977179
transform 1 0 19964 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_217
timestamp 1649977179
transform 1 0 21068 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_223
timestamp 1649977179
transform 1 0 21620 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_225
timestamp 1649977179
transform 1 0 21804 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_237
timestamp 1649977179
transform 1 0 22908 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_249
timestamp 1649977179
transform 1 0 24012 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_261
timestamp 1649977179
transform 1 0 25116 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_273
timestamp 1649977179
transform 1 0 26220 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_279
timestamp 1649977179
transform 1 0 26772 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_281
timestamp 1649977179
transform 1 0 26956 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_293
timestamp 1649977179
transform 1 0 28060 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_305
timestamp 1649977179
transform 1 0 29164 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_317
timestamp 1649977179
transform 1 0 30268 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_329
timestamp 1649977179
transform 1 0 31372 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_335
timestamp 1649977179
transform 1 0 31924 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_337
timestamp 1649977179
transform 1 0 32108 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_349
timestamp 1649977179
transform 1 0 33212 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_355
timestamp 1649977179
transform 1 0 33764 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_360
timestamp 1649977179
transform 1 0 34224 0 -1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3
timestamp 1649977179
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_15
timestamp 1649977179
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 1649977179
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_29
timestamp 1649977179
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_41
timestamp 1649977179
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_53
timestamp 1649977179
transform 1 0 5980 0 1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_4_60
timestamp 1649977179
transform 1 0 6624 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_72
timestamp 1649977179
transform 1 0 7728 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_85
timestamp 1649977179
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_97
timestamp 1649977179
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_109
timestamp 1649977179
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_121
timestamp 1649977179
transform 1 0 12236 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_127
timestamp 1649977179
transform 1 0 12788 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_139
timestamp 1649977179
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_141
timestamp 1649977179
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_153
timestamp 1649977179
transform 1 0 15180 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_165
timestamp 1649977179
transform 1 0 16284 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_177
timestamp 1649977179
transform 1 0 17388 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_185
timestamp 1649977179
transform 1 0 18124 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_4_190
timestamp 1649977179
transform 1 0 18584 0 1 4352
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_4_202
timestamp 1649977179
transform 1 0 19688 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_214
timestamp 1649977179
transform 1 0 20792 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_226
timestamp 1649977179
transform 1 0 21896 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_238
timestamp 1649977179
transform 1 0 23000 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_4_250
timestamp 1649977179
transform 1 0 24104 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_4_253
timestamp 1649977179
transform 1 0 24380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_265
timestamp 1649977179
transform 1 0 25484 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_277
timestamp 1649977179
transform 1 0 26588 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_289
timestamp 1649977179
transform 1 0 27692 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_301
timestamp 1649977179
transform 1 0 28796 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_307
timestamp 1649977179
transform 1 0 29348 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_321
timestamp 1649977179
transform 1 0 30636 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_333
timestamp 1649977179
transform 1 0 31740 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_345
timestamp 1649977179
transform 1 0 32844 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_357
timestamp 1649977179
transform 1 0 33948 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_363
timestamp 1649977179
transform 1 0 34500 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3
timestamp 1649977179
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_15
timestamp 1649977179
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_27
timestamp 1649977179
transform 1 0 3588 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_39
timestamp 1649977179
transform 1 0 4692 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_51
timestamp 1649977179
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_55
timestamp 1649977179
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_57
timestamp 1649977179
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_69
timestamp 1649977179
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_81
timestamp 1649977179
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_93
timestamp 1649977179
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_105
timestamp 1649977179
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_111
timestamp 1649977179
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_113
timestamp 1649977179
transform 1 0 11500 0 -1 5440
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_5_124
timestamp 1649977179
transform 1 0 12512 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_136
timestamp 1649977179
transform 1 0 13616 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_148
timestamp 1649977179
transform 1 0 14720 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_160
timestamp 1649977179
transform 1 0 15824 0 -1 5440
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_5_169
timestamp 1649977179
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_181
timestamp 1649977179
transform 1 0 17756 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_193
timestamp 1649977179
transform 1 0 18860 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_199
timestamp 1649977179
transform 1 0 19412 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_204
timestamp 1649977179
transform 1 0 19872 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_5_212
timestamp 1649977179
transform 1 0 20608 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_225
timestamp 1649977179
transform 1 0 21804 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_249
timestamp 1649977179
transform 1 0 24012 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_261
timestamp 1649977179
transform 1 0 25116 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_273
timestamp 1649977179
transform 1 0 26220 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_279
timestamp 1649977179
transform 1 0 26772 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_281
timestamp 1649977179
transform 1 0 26956 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_293
timestamp 1649977179
transform 1 0 28060 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_305
timestamp 1649977179
transform 1 0 29164 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_317
timestamp 1649977179
transform 1 0 30268 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_329
timestamp 1649977179
transform 1 0 31372 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_335
timestamp 1649977179
transform 1 0 31924 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_337
timestamp 1649977179
transform 1 0 32108 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_349
timestamp 1649977179
transform 1 0 33212 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_5_361
timestamp 1649977179
transform 1 0 34316 0 -1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3
timestamp 1649977179
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_15
timestamp 1649977179
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1649977179
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_29
timestamp 1649977179
transform 1 0 3772 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_6_40
timestamp 1649977179
transform 1 0 4784 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_6_46
timestamp 1649977179
transform 1 0 5336 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_52
timestamp 1649977179
transform 1 0 5888 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_58
timestamp 1649977179
transform 1 0 6440 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_70
timestamp 1649977179
transform 1 0 7544 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_6_82
timestamp 1649977179
transform 1 0 8648 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_85
timestamp 1649977179
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_97
timestamp 1649977179
transform 1 0 10028 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_105
timestamp 1649977179
transform 1 0 10764 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_116
timestamp 1649977179
transform 1 0 11776 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_128
timestamp 1649977179
transform 1 0 12880 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_141
timestamp 1649977179
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_153
timestamp 1649977179
transform 1 0 15180 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_165
timestamp 1649977179
transform 1 0 16284 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_177
timestamp 1649977179
transform 1 0 17388 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_189
timestamp 1649977179
transform 1 0 18492 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_195
timestamp 1649977179
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_197
timestamp 1649977179
transform 1 0 19228 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_209
timestamp 1649977179
transform 1 0 20332 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_221
timestamp 1649977179
transform 1 0 21436 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_233
timestamp 1649977179
transform 1 0 22540 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_245
timestamp 1649977179
transform 1 0 23644 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_251
timestamp 1649977179
transform 1 0 24196 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_253
timestamp 1649977179
transform 1 0 24380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_265
timestamp 1649977179
transform 1 0 25484 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_277
timestamp 1649977179
transform 1 0 26588 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_289
timestamp 1649977179
transform 1 0 27692 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_301
timestamp 1649977179
transform 1 0 28796 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_307
timestamp 1649977179
transform 1 0 29348 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_309
timestamp 1649977179
transform 1 0 29532 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_321
timestamp 1649977179
transform 1 0 30636 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_333
timestamp 1649977179
transform 1 0 31740 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_345
timestamp 1649977179
transform 1 0 32844 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_357
timestamp 1649977179
transform 1 0 33948 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_363
timestamp 1649977179
transform 1 0 34500 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3
timestamp 1649977179
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_15
timestamp 1649977179
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_27
timestamp 1649977179
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_7_39
timestamp 1649977179
transform 1 0 4692 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_7_43
timestamp 1649977179
transform 1 0 5060 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp 1649977179
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_57
timestamp 1649977179
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_69
timestamp 1649977179
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_81
timestamp 1649977179
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_93
timestamp 1649977179
transform 1 0 9660 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_105
timestamp 1649977179
transform 1 0 10764 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_111
timestamp 1649977179
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_113
timestamp 1649977179
transform 1 0 11500 0 -1 6528
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_7_126
timestamp 1649977179
transform 1 0 12696 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_138
timestamp 1649977179
transform 1 0 13800 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_150
timestamp 1649977179
transform 1 0 14904 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_162
timestamp 1649977179
transform 1 0 16008 0 -1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_7_169
timestamp 1649977179
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_181
timestamp 1649977179
transform 1 0 17756 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_193
timestamp 1649977179
transform 1 0 18860 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_205
timestamp 1649977179
transform 1 0 19964 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_217
timestamp 1649977179
transform 1 0 21068 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_223
timestamp 1649977179
transform 1 0 21620 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_225
timestamp 1649977179
transform 1 0 21804 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_237
timestamp 1649977179
transform 1 0 22908 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_249
timestamp 1649977179
transform 1 0 24012 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_261
timestamp 1649977179
transform 1 0 25116 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_273
timestamp 1649977179
transform 1 0 26220 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_279
timestamp 1649977179
transform 1 0 26772 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_281
timestamp 1649977179
transform 1 0 26956 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_296
timestamp 1649977179
transform 1 0 28336 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_308
timestamp 1649977179
transform 1 0 29440 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_320
timestamp 1649977179
transform 1 0 30544 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_332
timestamp 1649977179
transform 1 0 31648 0 -1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_7_349
timestamp 1649977179
transform 1 0 33212 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_7_361
timestamp 1649977179
transform 1 0 34316 0 -1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3
timestamp 1649977179
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_15
timestamp 1649977179
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 1649977179
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_29
timestamp 1649977179
transform 1 0 3772 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_37
timestamp 1649977179
transform 1 0 4508 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_8_41
timestamp 1649977179
transform 1 0 4876 0 1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_8_49
timestamp 1649977179
transform 1 0 5612 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_61
timestamp 1649977179
transform 1 0 6716 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_73
timestamp 1649977179
transform 1 0 7820 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_8_81
timestamp 1649977179
transform 1 0 8556 0 1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_8_85
timestamp 1649977179
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_97
timestamp 1649977179
transform 1 0 10028 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_109
timestamp 1649977179
transform 1 0 11132 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_115
timestamp 1649977179
transform 1 0 11684 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_122
timestamp 1649977179
transform 1 0 12328 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_134
timestamp 1649977179
transform 1 0 13432 0 1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_8_141
timestamp 1649977179
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_153
timestamp 1649977179
transform 1 0 15180 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_165
timestamp 1649977179
transform 1 0 16284 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_177
timestamp 1649977179
transform 1 0 17388 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_189
timestamp 1649977179
transform 1 0 18492 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_195
timestamp 1649977179
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_197
timestamp 1649977179
transform 1 0 19228 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_8_208
timestamp 1649977179
transform 1 0 20240 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_217
timestamp 1649977179
transform 1 0 21068 0 1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_8_224
timestamp 1649977179
transform 1 0 21712 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_236
timestamp 1649977179
transform 1 0 22816 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_248
timestamp 1649977179
transform 1 0 23920 0 1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_8_253
timestamp 1649977179
transform 1 0 24380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_265
timestamp 1649977179
transform 1 0 25484 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_277
timestamp 1649977179
transform 1 0 26588 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_289
timestamp 1649977179
transform 1 0 27692 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_301
timestamp 1649977179
transform 1 0 28796 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_307
timestamp 1649977179
transform 1 0 29348 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_309
timestamp 1649977179
transform 1 0 29532 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_317
timestamp 1649977179
transform 1 0 30268 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_321
timestamp 1649977179
transform 1 0 30636 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_333
timestamp 1649977179
transform 1 0 31740 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_345
timestamp 1649977179
transform 1 0 32844 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_8_353
timestamp 1649977179
transform 1 0 33580 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_8_360
timestamp 1649977179
transform 1 0 34224 0 1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_9_5
timestamp 1649977179
transform 1 0 1564 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_17
timestamp 1649977179
transform 1 0 2668 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_25
timestamp 1649977179
transform 1 0 3404 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_9_47
timestamp 1649977179
transform 1 0 5428 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_55
timestamp 1649977179
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_57
timestamp 1649977179
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_69
timestamp 1649977179
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_81
timestamp 1649977179
transform 1 0 8556 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_93
timestamp 1649977179
transform 1 0 9660 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_105
timestamp 1649977179
transform 1 0 10764 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_111
timestamp 1649977179
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_9_113
timestamp 1649977179
transform 1 0 11500 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_119
timestamp 1649977179
transform 1 0 12052 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_127
timestamp 1649977179
transform 1 0 12788 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_139
timestamp 1649977179
transform 1 0 13892 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_145
timestamp 1649977179
transform 1 0 14444 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_149
timestamp 1649977179
transform 1 0 14812 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_161
timestamp 1649977179
transform 1 0 15916 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_167
timestamp 1649977179
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_169
timestamp 1649977179
transform 1 0 16652 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_181
timestamp 1649977179
transform 1 0 17756 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_193
timestamp 1649977179
transform 1 0 18860 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_205
timestamp 1649977179
transform 1 0 19964 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_217
timestamp 1649977179
transform 1 0 21068 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_223
timestamp 1649977179
transform 1 0 21620 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_225
timestamp 1649977179
transform 1 0 21804 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_237
timestamp 1649977179
transform 1 0 22908 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_249
timestamp 1649977179
transform 1 0 24012 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_261
timestamp 1649977179
transform 1 0 25116 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_9_273
timestamp 1649977179
transform 1 0 26220 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_276
timestamp 1649977179
transform 1 0 26496 0 -1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_9_290
timestamp 1649977179
transform 1 0 27784 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_302
timestamp 1649977179
transform 1 0 28888 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_314
timestamp 1649977179
transform 1 0 29992 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_326
timestamp 1649977179
transform 1 0 31096 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_334
timestamp 1649977179
transform 1 0 31832 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_337
timestamp 1649977179
transform 1 0 32108 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_349
timestamp 1649977179
transform 1 0 33212 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_361
timestamp 1649977179
transform 1 0 34316 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_10_7
timestamp 1649977179
transform 1 0 1748 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_19
timestamp 1649977179
transform 1 0 2852 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 1649977179
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_29
timestamp 1649977179
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_41
timestamp 1649977179
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_53
timestamp 1649977179
transform 1 0 5980 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_65
timestamp 1649977179
transform 1 0 7084 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_77
timestamp 1649977179
transform 1 0 8188 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_83
timestamp 1649977179
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_85
timestamp 1649977179
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_97
timestamp 1649977179
transform 1 0 10028 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_10_108
timestamp 1649977179
transform 1 0 11040 0 1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_10_119
timestamp 1649977179
transform 1 0 12052 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_131
timestamp 1649977179
transform 1 0 13156 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_139
timestamp 1649977179
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_141
timestamp 1649977179
transform 1 0 14076 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_153
timestamp 1649977179
transform 1 0 15180 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_165
timestamp 1649977179
transform 1 0 16284 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_177
timestamp 1649977179
transform 1 0 17388 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_189
timestamp 1649977179
transform 1 0 18492 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_195
timestamp 1649977179
transform 1 0 19044 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_197
timestamp 1649977179
transform 1 0 19228 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_201
timestamp 1649977179
transform 1 0 19596 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_206
timestamp 1649977179
transform 1 0 20056 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_221
timestamp 1649977179
transform 1 0 21436 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_225
timestamp 1649977179
transform 1 0 21804 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_231
timestamp 1649977179
transform 1 0 22356 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_243
timestamp 1649977179
transform 1 0 23460 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_251
timestamp 1649977179
transform 1 0 24196 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_253
timestamp 1649977179
transform 1 0 24380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_265
timestamp 1649977179
transform 1 0 25484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_277
timestamp 1649977179
transform 1 0 26588 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_283
timestamp 1649977179
transform 1 0 27140 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_287
timestamp 1649977179
transform 1 0 27508 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_299
timestamp 1649977179
transform 1 0 28612 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_307
timestamp 1649977179
transform 1 0 29348 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_309
timestamp 1649977179
transform 1 0 29532 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_321
timestamp 1649977179
transform 1 0 30636 0 1 7616
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_10_341
timestamp 1649977179
transform 1 0 32476 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_353
timestamp 1649977179
transform 1 0 33580 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_10_361
timestamp 1649977179
transform 1 0 34316 0 1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3
timestamp 1649977179
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_15
timestamp 1649977179
transform 1 0 2484 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_27
timestamp 1649977179
transform 1 0 3588 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_39
timestamp 1649977179
transform 1 0 4692 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_51
timestamp 1649977179
transform 1 0 5796 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_55
timestamp 1649977179
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_57
timestamp 1649977179
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_69
timestamp 1649977179
transform 1 0 7452 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_81
timestamp 1649977179
transform 1 0 8556 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_93
timestamp 1649977179
transform 1 0 9660 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_105
timestamp 1649977179
transform 1 0 10764 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_111
timestamp 1649977179
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_11_113
timestamp 1649977179
transform 1 0 11500 0 -1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_11_126
timestamp 1649977179
transform 1 0 12696 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_138
timestamp 1649977179
transform 1 0 13800 0 -1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_11_145
timestamp 1649977179
transform 1 0 14444 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_157
timestamp 1649977179
transform 1 0 15548 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_11_165
timestamp 1649977179
transform 1 0 16284 0 -1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_11_169
timestamp 1649977179
transform 1 0 16652 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_181
timestamp 1649977179
transform 1 0 17756 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_193
timestamp 1649977179
transform 1 0 18860 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_205
timestamp 1649977179
transform 1 0 19964 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_217
timestamp 1649977179
transform 1 0 21068 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_223
timestamp 1649977179
transform 1 0 21620 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_225
timestamp 1649977179
transform 1 0 21804 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_237
timestamp 1649977179
transform 1 0 22908 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_249
timestamp 1649977179
transform 1 0 24012 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_261
timestamp 1649977179
transform 1 0 25116 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_273
timestamp 1649977179
transform 1 0 26220 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_279
timestamp 1649977179
transform 1 0 26772 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_281
timestamp 1649977179
transform 1 0 26956 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_289
timestamp 1649977179
transform 1 0 27692 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_310
timestamp 1649977179
transform 1 0 29624 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_322
timestamp 1649977179
transform 1 0 30728 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_11_334
timestamp 1649977179
transform 1 0 31832 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_337
timestamp 1649977179
transform 1 0 32108 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_349
timestamp 1649977179
transform 1 0 33212 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_11_361
timestamp 1649977179
transform 1 0 34316 0 -1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3
timestamp 1649977179
transform 1 0 1380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_15
timestamp 1649977179
transform 1 0 2484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_27
timestamp 1649977179
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_29
timestamp 1649977179
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_41
timestamp 1649977179
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_53
timestamp 1649977179
transform 1 0 5980 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_65
timestamp 1649977179
transform 1 0 7084 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_77
timestamp 1649977179
transform 1 0 8188 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_83
timestamp 1649977179
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_85
timestamp 1649977179
transform 1 0 8924 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_97
timestamp 1649977179
transform 1 0 10028 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_109
timestamp 1649977179
transform 1 0 11132 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_128
timestamp 1649977179
transform 1 0 12880 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_141
timestamp 1649977179
transform 1 0 14076 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_153
timestamp 1649977179
transform 1 0 15180 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_165
timestamp 1649977179
transform 1 0 16284 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_177
timestamp 1649977179
transform 1 0 17388 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_189
timestamp 1649977179
transform 1 0 18492 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_195
timestamp 1649977179
transform 1 0 19044 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_197
timestamp 1649977179
transform 1 0 19228 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_209
timestamp 1649977179
transform 1 0 20332 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_12_221
timestamp 1649977179
transform 1 0 21436 0 1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_12_237
timestamp 1649977179
transform 1 0 22908 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_12_249
timestamp 1649977179
transform 1 0 24012 0 1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_12_253
timestamp 1649977179
transform 1 0 24380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_265
timestamp 1649977179
transform 1 0 25484 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_277
timestamp 1649977179
transform 1 0 26588 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_289
timestamp 1649977179
transform 1 0 27692 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_295
timestamp 1649977179
transform 1 0 28244 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_12_302
timestamp 1649977179
transform 1 0 28888 0 1 8704
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_12_309
timestamp 1649977179
transform 1 0 29532 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_321
timestamp 1649977179
transform 1 0 30636 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_333
timestamp 1649977179
transform 1 0 31740 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_345
timestamp 1649977179
transform 1 0 32844 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_12_353
timestamp 1649977179
transform 1 0 33580 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_12_360
timestamp 1649977179
transform 1 0 34224 0 1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3
timestamp 1649977179
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_15
timestamp 1649977179
transform 1 0 2484 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_27
timestamp 1649977179
transform 1 0 3588 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_51
timestamp 1649977179
transform 1 0 5796 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_55
timestamp 1649977179
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_59
timestamp 1649977179
transform 1 0 6532 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_71
timestamp 1649977179
transform 1 0 7636 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_83
timestamp 1649977179
transform 1 0 8740 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_95
timestamp 1649977179
transform 1 0 9844 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_107
timestamp 1649977179
transform 1 0 10948 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_111
timestamp 1649977179
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_113
timestamp 1649977179
transform 1 0 11500 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_125
timestamp 1649977179
transform 1 0 12604 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_13_133
timestamp 1649977179
transform 1 0 13340 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_139
timestamp 1649977179
transform 1 0 13892 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_151
timestamp 1649977179
transform 1 0 14996 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_163
timestamp 1649977179
transform 1 0 16100 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_167
timestamp 1649977179
transform 1 0 16468 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_169
timestamp 1649977179
transform 1 0 16652 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_181
timestamp 1649977179
transform 1 0 17756 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_193
timestamp 1649977179
transform 1 0 18860 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_205
timestamp 1649977179
transform 1 0 19964 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_217
timestamp 1649977179
transform 1 0 21068 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_223
timestamp 1649977179
transform 1 0 21620 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_225
timestamp 1649977179
transform 1 0 21804 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_237
timestamp 1649977179
transform 1 0 22908 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_249
timestamp 1649977179
transform 1 0 24012 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_261
timestamp 1649977179
transform 1 0 25116 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_273
timestamp 1649977179
transform 1 0 26220 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_279
timestamp 1649977179
transform 1 0 26772 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_281
timestamp 1649977179
transform 1 0 26956 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_293
timestamp 1649977179
transform 1 0 28060 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_305
timestamp 1649977179
transform 1 0 29164 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_317
timestamp 1649977179
transform 1 0 30268 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_329
timestamp 1649977179
transform 1 0 31372 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_335
timestamp 1649977179
transform 1 0 31924 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_337
timestamp 1649977179
transform 1 0 32108 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_349
timestamp 1649977179
transform 1 0 33212 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_361
timestamp 1649977179
transform 1 0 34316 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_14_3
timestamp 1649977179
transform 1 0 1380 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_15
timestamp 1649977179
transform 1 0 2484 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_27
timestamp 1649977179
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_29
timestamp 1649977179
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_44
timestamp 1649977179
transform 1 0 5152 0 1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_14_50
timestamp 1649977179
transform 1 0 5704 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_62
timestamp 1649977179
transform 1 0 6808 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_74
timestamp 1649977179
transform 1 0 7912 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_82
timestamp 1649977179
transform 1 0 8648 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_85
timestamp 1649977179
transform 1 0 8924 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_97
timestamp 1649977179
transform 1 0 10028 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_14_121
timestamp 1649977179
transform 1 0 12236 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_129
timestamp 1649977179
transform 1 0 12972 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_136
timestamp 1649977179
transform 1 0 13616 0 1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_14_141
timestamp 1649977179
transform 1 0 14076 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_14_153
timestamp 1649977179
transform 1 0 15180 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_157
timestamp 1649977179
transform 1 0 15548 0 1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_14_181
timestamp 1649977179
transform 1 0 17756 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_14_193
timestamp 1649977179
transform 1 0 18860 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_14_197
timestamp 1649977179
transform 1 0 19228 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_14_205
timestamp 1649977179
transform 1 0 19964 0 1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_14_220
timestamp 1649977179
transform 1 0 21344 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_232
timestamp 1649977179
transform 1 0 22448 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_244
timestamp 1649977179
transform 1 0 23552 0 1 9792
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_14_253
timestamp 1649977179
transform 1 0 24380 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_265
timestamp 1649977179
transform 1 0 25484 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_277
timestamp 1649977179
transform 1 0 26588 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_289
timestamp 1649977179
transform 1 0 27692 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_301
timestamp 1649977179
transform 1 0 28796 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_307
timestamp 1649977179
transform 1 0 29348 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_309
timestamp 1649977179
transform 1 0 29532 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_321
timestamp 1649977179
transform 1 0 30636 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_333
timestamp 1649977179
transform 1 0 31740 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_345
timestamp 1649977179
transform 1 0 32844 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_357
timestamp 1649977179
transform 1 0 33948 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_363
timestamp 1649977179
transform 1 0 34500 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_3
timestamp 1649977179
transform 1 0 1380 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_15
timestamp 1649977179
transform 1 0 2484 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_15_27
timestamp 1649977179
transform 1 0 3588 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_15_32
timestamp 1649977179
transform 1 0 4048 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_15_40
timestamp 1649977179
transform 1 0 4784 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_52
timestamp 1649977179
transform 1 0 5888 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_15_57
timestamp 1649977179
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_69
timestamp 1649977179
transform 1 0 7452 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_81
timestamp 1649977179
transform 1 0 8556 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_93
timestamp 1649977179
transform 1 0 9660 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_105
timestamp 1649977179
transform 1 0 10764 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_111
timestamp 1649977179
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_113
timestamp 1649977179
transform 1 0 11500 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_128
timestamp 1649977179
transform 1 0 12880 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_15_134
timestamp 1649977179
transform 1 0 13432 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_146
timestamp 1649977179
transform 1 0 14536 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_158
timestamp 1649977179
transform 1 0 15640 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_166
timestamp 1649977179
transform 1 0 16376 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_15_169
timestamp 1649977179
transform 1 0 16652 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_181
timestamp 1649977179
transform 1 0 17756 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_185
timestamp 1649977179
transform 1 0 18124 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_206
timestamp 1649977179
transform 1 0 20056 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_218
timestamp 1649977179
transform 1 0 21160 0 -1 10880
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_15_225
timestamp 1649977179
transform 1 0 21804 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_237
timestamp 1649977179
transform 1 0 22908 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_249
timestamp 1649977179
transform 1 0 24012 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_261
timestamp 1649977179
transform 1 0 25116 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_273
timestamp 1649977179
transform 1 0 26220 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_279
timestamp 1649977179
transform 1 0 26772 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_281
timestamp 1649977179
transform 1 0 26956 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_15_289
timestamp 1649977179
transform 1 0 27692 0 -1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_15_312
timestamp 1649977179
transform 1 0 29808 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_324
timestamp 1649977179
transform 1 0 30912 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_337
timestamp 1649977179
transform 1 0 32108 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_349
timestamp 1649977179
transform 1 0 33212 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_15_361
timestamp 1649977179
transform 1 0 34316 0 -1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_16_3
timestamp 1649977179
transform 1 0 1380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_15
timestamp 1649977179
transform 1 0 2484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_27
timestamp 1649977179
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_29
timestamp 1649977179
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_41
timestamp 1649977179
transform 1 0 4876 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_55
timestamp 1649977179
transform 1 0 6164 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_67
timestamp 1649977179
transform 1 0 7268 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_79
timestamp 1649977179
transform 1 0 8372 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_83
timestamp 1649977179
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_85
timestamp 1649977179
transform 1 0 8924 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_97
timestamp 1649977179
transform 1 0 10028 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_111
timestamp 1649977179
transform 1 0 11316 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_136
timestamp 1649977179
transform 1 0 13616 0 1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_16_141
timestamp 1649977179
transform 1 0 14076 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_153
timestamp 1649977179
transform 1 0 15180 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_165
timestamp 1649977179
transform 1 0 16284 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_177
timestamp 1649977179
transform 1 0 17388 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_189
timestamp 1649977179
transform 1 0 18492 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_195
timestamp 1649977179
transform 1 0 19044 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_197
timestamp 1649977179
transform 1 0 19228 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_211
timestamp 1649977179
transform 1 0 20516 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_223
timestamp 1649977179
transform 1 0 21620 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_235
timestamp 1649977179
transform 1 0 22724 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_247
timestamp 1649977179
transform 1 0 23828 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_251
timestamp 1649977179
transform 1 0 24196 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_253
timestamp 1649977179
transform 1 0 24380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_265
timestamp 1649977179
transform 1 0 25484 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_277
timestamp 1649977179
transform 1 0 26588 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_16_289
timestamp 1649977179
transform 1 0 27692 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_293
timestamp 1649977179
transform 1 0 28060 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_16_300
timestamp 1649977179
transform 1 0 28704 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_309
timestamp 1649977179
transform 1 0 29532 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_314
timestamp 1649977179
transform 1 0 29992 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_318
timestamp 1649977179
transform 1 0 30360 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_321
timestamp 1649977179
transform 1 0 30636 0 1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_16_334
timestamp 1649977179
transform 1 0 31832 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_346
timestamp 1649977179
transform 1 0 32936 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_358
timestamp 1649977179
transform 1 0 34040 0 1 10880
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_17_3
timestamp 1649977179
transform 1 0 1380 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_15
timestamp 1649977179
transform 1 0 2484 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_27
timestamp 1649977179
transform 1 0 3588 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_39
timestamp 1649977179
transform 1 0 4692 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_17_47
timestamp 1649977179
transform 1 0 5428 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_17_52
timestamp 1649977179
transform 1 0 5888 0 -1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_17_64
timestamp 1649977179
transform 1 0 6992 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_76
timestamp 1649977179
transform 1 0 8096 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_88
timestamp 1649977179
transform 1 0 9200 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_100
timestamp 1649977179
transform 1 0 10304 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_113
timestamp 1649977179
transform 1 0 11500 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_125
timestamp 1649977179
transform 1 0 12604 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_137
timestamp 1649977179
transform 1 0 13708 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_149
timestamp 1649977179
transform 1 0 14812 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_161
timestamp 1649977179
transform 1 0 15916 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_167
timestamp 1649977179
transform 1 0 16468 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_169
timestamp 1649977179
transform 1 0 16652 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_181
timestamp 1649977179
transform 1 0 17756 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_193
timestamp 1649977179
transform 1 0 18860 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_205
timestamp 1649977179
transform 1 0 19964 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_17_213
timestamp 1649977179
transform 1 0 20700 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_17_221
timestamp 1649977179
transform 1 0 21436 0 -1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_17_225
timestamp 1649977179
transform 1 0 21804 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_237
timestamp 1649977179
transform 1 0 22908 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_249
timestamp 1649977179
transform 1 0 24012 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_261
timestamp 1649977179
transform 1 0 25116 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_273
timestamp 1649977179
transform 1 0 26220 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_279
timestamp 1649977179
transform 1 0 26772 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_281
timestamp 1649977179
transform 1 0 26956 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_293
timestamp 1649977179
transform 1 0 28060 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_305
timestamp 1649977179
transform 1 0 29164 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_317
timestamp 1649977179
transform 1 0 30268 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_329
timestamp 1649977179
transform 1 0 31372 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_335
timestamp 1649977179
transform 1 0 31924 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_337
timestamp 1649977179
transform 1 0 32108 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_349
timestamp 1649977179
transform 1 0 33212 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_355
timestamp 1649977179
transform 1 0 33764 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_360
timestamp 1649977179
transform 1 0 34224 0 -1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_18_5
timestamp 1649977179
transform 1 0 1564 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_17
timestamp 1649977179
transform 1 0 2668 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_18_25
timestamp 1649977179
transform 1 0 3404 0 1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_18_29
timestamp 1649977179
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_41
timestamp 1649977179
transform 1 0 4876 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_55
timestamp 1649977179
transform 1 0 6164 0 1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_18_63
timestamp 1649977179
transform 1 0 6900 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_75
timestamp 1649977179
transform 1 0 8004 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_83
timestamp 1649977179
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_85
timestamp 1649977179
transform 1 0 8924 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_97
timestamp 1649977179
transform 1 0 10028 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_109
timestamp 1649977179
transform 1 0 11132 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_121
timestamp 1649977179
transform 1 0 12236 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_133
timestamp 1649977179
transform 1 0 13340 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_139
timestamp 1649977179
transform 1 0 13892 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_141
timestamp 1649977179
transform 1 0 14076 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_153
timestamp 1649977179
transform 1 0 15180 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_165
timestamp 1649977179
transform 1 0 16284 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_177
timestamp 1649977179
transform 1 0 17388 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_189
timestamp 1649977179
transform 1 0 18492 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_195
timestamp 1649977179
transform 1 0 19044 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_197
timestamp 1649977179
transform 1 0 19228 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_205
timestamp 1649977179
transform 1 0 19964 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_209
timestamp 1649977179
transform 1 0 20332 0 1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_18_222
timestamp 1649977179
transform 1 0 21528 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_234
timestamp 1649977179
transform 1 0 22632 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_246
timestamp 1649977179
transform 1 0 23736 0 1 11968
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_18_253
timestamp 1649977179
transform 1 0 24380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_265
timestamp 1649977179
transform 1 0 25484 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_277
timestamp 1649977179
transform 1 0 26588 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_289
timestamp 1649977179
transform 1 0 27692 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_301
timestamp 1649977179
transform 1 0 28796 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_307
timestamp 1649977179
transform 1 0 29348 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_309
timestamp 1649977179
transform 1 0 29532 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_321
timestamp 1649977179
transform 1 0 30636 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_333
timestamp 1649977179
transform 1 0 31740 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_345
timestamp 1649977179
transform 1 0 32844 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_357
timestamp 1649977179
transform 1 0 33948 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_363
timestamp 1649977179
transform 1 0 34500 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_13
timestamp 1649977179
transform 1 0 2300 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_25
timestamp 1649977179
transform 1 0 3404 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_37
timestamp 1649977179
transform 1 0 4508 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_49
timestamp 1649977179
transform 1 0 5612 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_55
timestamp 1649977179
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_60
timestamp 1649977179
transform 1 0 6624 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_72
timestamp 1649977179
transform 1 0 7728 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_84
timestamp 1649977179
transform 1 0 8832 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_96
timestamp 1649977179
transform 1 0 9936 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_108
timestamp 1649977179
transform 1 0 11040 0 -1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_19_113
timestamp 1649977179
transform 1 0 11500 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_19_125
timestamp 1649977179
transform 1 0 12604 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_129
timestamp 1649977179
transform 1 0 12972 0 -1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_19_154
timestamp 1649977179
transform 1 0 15272 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_19_166
timestamp 1649977179
transform 1 0 16376 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_19_169
timestamp 1649977179
transform 1 0 16652 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_181
timestamp 1649977179
transform 1 0 17756 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_193
timestamp 1649977179
transform 1 0 18860 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_19_204
timestamp 1649977179
transform 1 0 19872 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_212
timestamp 1649977179
transform 1 0 20608 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_220
timestamp 1649977179
transform 1 0 21344 0 -1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_19_227
timestamp 1649977179
transform 1 0 21988 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_239
timestamp 1649977179
transform 1 0 23092 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_251
timestamp 1649977179
transform 1 0 24196 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_263
timestamp 1649977179
transform 1 0 25300 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_275
timestamp 1649977179
transform 1 0 26404 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_279
timestamp 1649977179
transform 1 0 26772 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_281
timestamp 1649977179
transform 1 0 26956 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_293
timestamp 1649977179
transform 1 0 28060 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_300
timestamp 1649977179
transform 1 0 28704 0 -1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_19_306
timestamp 1649977179
transform 1 0 29256 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_318
timestamp 1649977179
transform 1 0 30360 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_330
timestamp 1649977179
transform 1 0 31464 0 -1 13056
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_19_337
timestamp 1649977179
transform 1 0 32108 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_349
timestamp 1649977179
transform 1 0 33212 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_19_361
timestamp 1649977179
transform 1 0 34316 0 -1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_20_3
timestamp 1649977179
transform 1 0 1380 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_15
timestamp 1649977179
transform 1 0 2484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_27
timestamp 1649977179
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_29
timestamp 1649977179
transform 1 0 3772 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_53
timestamp 1649977179
transform 1 0 5980 0 1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_20_59
timestamp 1649977179
transform 1 0 6532 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_71
timestamp 1649977179
transform 1 0 7636 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_83
timestamp 1649977179
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_85
timestamp 1649977179
transform 1 0 8924 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_97
timestamp 1649977179
transform 1 0 10028 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_109
timestamp 1649977179
transform 1 0 11132 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_121
timestamp 1649977179
transform 1 0 12236 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_133
timestamp 1649977179
transform 1 0 13340 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_139
timestamp 1649977179
transform 1 0 13892 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_144
timestamp 1649977179
transform 1 0 14352 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_156
timestamp 1649977179
transform 1 0 15456 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_168
timestamp 1649977179
transform 1 0 16560 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_180
timestamp 1649977179
transform 1 0 17664 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_192
timestamp 1649977179
transform 1 0 18768 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_197
timestamp 1649977179
transform 1 0 19228 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_205
timestamp 1649977179
transform 1 0 19964 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_209
timestamp 1649977179
transform 1 0 20332 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_215
timestamp 1649977179
transform 1 0 20884 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_20_226
timestamp 1649977179
transform 1 0 21896 0 1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_20_232
timestamp 1649977179
transform 1 0 22448 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_244
timestamp 1649977179
transform 1 0 23552 0 1 13056
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_20_253
timestamp 1649977179
transform 1 0 24380 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_265
timestamp 1649977179
transform 1 0 25484 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_277
timestamp 1649977179
transform 1 0 26588 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_289
timestamp 1649977179
transform 1 0 27692 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_301
timestamp 1649977179
transform 1 0 28796 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_307
timestamp 1649977179
transform 1 0 29348 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_309
timestamp 1649977179
transform 1 0 29532 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_314
timestamp 1649977179
transform 1 0 29992 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_318
timestamp 1649977179
transform 1 0 30360 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_321
timestamp 1649977179
transform 1 0 30636 0 1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_20_334
timestamp 1649977179
transform 1 0 31832 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_346
timestamp 1649977179
transform 1 0 32936 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_358
timestamp 1649977179
transform 1 0 34040 0 1 13056
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_21_3
timestamp 1649977179
transform 1 0 1380 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_15
timestamp 1649977179
transform 1 0 2484 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_27
timestamp 1649977179
transform 1 0 3588 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_21_39
timestamp 1649977179
transform 1 0 4692 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_21_45
timestamp 1649977179
transform 1 0 5244 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_21_53
timestamp 1649977179
transform 1 0 5980 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_21_57
timestamp 1649977179
transform 1 0 6348 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_61
timestamp 1649977179
transform 1 0 6716 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_64
timestamp 1649977179
transform 1 0 6992 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_76
timestamp 1649977179
transform 1 0 8096 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_88
timestamp 1649977179
transform 1 0 9200 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_100
timestamp 1649977179
transform 1 0 10304 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_113
timestamp 1649977179
transform 1 0 11500 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_125
timestamp 1649977179
transform 1 0 12604 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_137
timestamp 1649977179
transform 1 0 13708 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_149
timestamp 1649977179
transform 1 0 14812 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_161
timestamp 1649977179
transform 1 0 15916 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_167
timestamp 1649977179
transform 1 0 16468 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_169
timestamp 1649977179
transform 1 0 16652 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_181
timestamp 1649977179
transform 1 0 17756 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_193
timestamp 1649977179
transform 1 0 18860 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_205
timestamp 1649977179
transform 1 0 19964 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_217
timestamp 1649977179
transform 1 0 21068 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_223
timestamp 1649977179
transform 1 0 21620 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_225
timestamp 1649977179
transform 1 0 21804 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_237
timestamp 1649977179
transform 1 0 22908 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_249
timestamp 1649977179
transform 1 0 24012 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_261
timestamp 1649977179
transform 1 0 25116 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_273
timestamp 1649977179
transform 1 0 26220 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_279
timestamp 1649977179
transform 1 0 26772 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_281
timestamp 1649977179
transform 1 0 26956 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_313
timestamp 1649977179
transform 1 0 29900 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_325
timestamp 1649977179
transform 1 0 31004 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_21_333
timestamp 1649977179
transform 1 0 31740 0 -1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_21_337
timestamp 1649977179
transform 1 0 32108 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_349
timestamp 1649977179
transform 1 0 33212 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_355
timestamp 1649977179
transform 1 0 33764 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_360
timestamp 1649977179
transform 1 0 34224 0 -1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_22_3
timestamp 1649977179
transform 1 0 1380 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_15
timestamp 1649977179
transform 1 0 2484 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_27
timestamp 1649977179
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_29
timestamp 1649977179
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_41
timestamp 1649977179
transform 1 0 4876 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_62
timestamp 1649977179
transform 1 0 6808 0 1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_22_68
timestamp 1649977179
transform 1 0 7360 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_80
timestamp 1649977179
transform 1 0 8464 0 1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_22_85
timestamp 1649977179
transform 1 0 8924 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_97
timestamp 1649977179
transform 1 0 10028 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_109
timestamp 1649977179
transform 1 0 11132 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_121
timestamp 1649977179
transform 1 0 12236 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_133
timestamp 1649977179
transform 1 0 13340 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_139
timestamp 1649977179
transform 1 0 13892 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_141
timestamp 1649977179
transform 1 0 14076 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_153
timestamp 1649977179
transform 1 0 15180 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_165
timestamp 1649977179
transform 1 0 16284 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_177
timestamp 1649977179
transform 1 0 17388 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_189
timestamp 1649977179
transform 1 0 18492 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_195
timestamp 1649977179
transform 1 0 19044 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_197
timestamp 1649977179
transform 1 0 19228 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_209
timestamp 1649977179
transform 1 0 20332 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_221
timestamp 1649977179
transform 1 0 21436 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_233
timestamp 1649977179
transform 1 0 22540 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_245
timestamp 1649977179
transform 1 0 23644 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_251
timestamp 1649977179
transform 1 0 24196 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_253
timestamp 1649977179
transform 1 0 24380 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_265
timestamp 1649977179
transform 1 0 25484 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_277
timestamp 1649977179
transform 1 0 26588 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_289
timestamp 1649977179
transform 1 0 27692 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_301
timestamp 1649977179
transform 1 0 28796 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_307
timestamp 1649977179
transform 1 0 29348 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_309
timestamp 1649977179
transform 1 0 29532 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_321
timestamp 1649977179
transform 1 0 30636 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_333
timestamp 1649977179
transform 1 0 31740 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_345
timestamp 1649977179
transform 1 0 32844 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_357
timestamp 1649977179
transform 1 0 33948 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_363
timestamp 1649977179
transform 1 0 34500 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_3
timestamp 1649977179
transform 1 0 1380 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_15
timestamp 1649977179
transform 1 0 2484 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_27
timestamp 1649977179
transform 1 0 3588 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_39
timestamp 1649977179
transform 1 0 4692 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_51
timestamp 1649977179
transform 1 0 5796 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_55
timestamp 1649977179
transform 1 0 6164 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_57
timestamp 1649977179
transform 1 0 6348 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_65
timestamp 1649977179
transform 1 0 7084 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_23_69
timestamp 1649977179
transform 1 0 7452 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_81
timestamp 1649977179
transform 1 0 8556 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_93
timestamp 1649977179
transform 1 0 9660 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_105
timestamp 1649977179
transform 1 0 10764 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_111
timestamp 1649977179
transform 1 0 11316 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_113
timestamp 1649977179
transform 1 0 11500 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_125
timestamp 1649977179
transform 1 0 12604 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_137
timestamp 1649977179
transform 1 0 13708 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_23_146
timestamp 1649977179
transform 1 0 14536 0 -1 15232
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_23_155
timestamp 1649977179
transform 1 0 15364 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_23_167
timestamp 1649977179
transform 1 0 16468 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_169
timestamp 1649977179
transform 1 0 16652 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_181
timestamp 1649977179
transform 1 0 17756 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_193
timestamp 1649977179
transform 1 0 18860 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_205
timestamp 1649977179
transform 1 0 19964 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_23_220
timestamp 1649977179
transform 1 0 21344 0 -1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_23_227
timestamp 1649977179
transform 1 0 21988 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_239
timestamp 1649977179
transform 1 0 23092 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_251
timestamp 1649977179
transform 1 0 24196 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_263
timestamp 1649977179
transform 1 0 25300 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_275
timestamp 1649977179
transform 1 0 26404 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_279
timestamp 1649977179
transform 1 0 26772 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_281
timestamp 1649977179
transform 1 0 26956 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_23_293
timestamp 1649977179
transform 1 0 28060 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_314
timestamp 1649977179
transform 1 0 29992 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_326
timestamp 1649977179
transform 1 0 31096 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_334
timestamp 1649977179
transform 1 0 31832 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_23_337
timestamp 1649977179
transform 1 0 32108 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_349
timestamp 1649977179
transform 1 0 33212 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_23_361
timestamp 1649977179
transform 1 0 34316 0 -1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_24_3
timestamp 1649977179
transform 1 0 1380 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_15
timestamp 1649977179
transform 1 0 2484 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_27
timestamp 1649977179
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_29
timestamp 1649977179
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_41
timestamp 1649977179
transform 1 0 4876 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_53
timestamp 1649977179
transform 1 0 5980 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_57
timestamp 1649977179
transform 1 0 6348 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_24_67
timestamp 1649977179
transform 1 0 7268 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_24_76
timestamp 1649977179
transform 1 0 8096 0 1 15232
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_24_85
timestamp 1649977179
transform 1 0 8924 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_97
timestamp 1649977179
transform 1 0 10028 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_109
timestamp 1649977179
transform 1 0 11132 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_121
timestamp 1649977179
transform 1 0 12236 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_133
timestamp 1649977179
transform 1 0 13340 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_136
timestamp 1649977179
transform 1 0 13616 0 1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_24_161
timestamp 1649977179
transform 1 0 15916 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_173
timestamp 1649977179
transform 1 0 17020 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_185
timestamp 1649977179
transform 1 0 18124 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_24_193
timestamp 1649977179
transform 1 0 18860 0 1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_24_197
timestamp 1649977179
transform 1 0 19228 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_229
timestamp 1649977179
transform 1 0 22172 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_241
timestamp 1649977179
transform 1 0 23276 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_24_249
timestamp 1649977179
transform 1 0 24012 0 1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_24_253
timestamp 1649977179
transform 1 0 24380 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_265
timestamp 1649977179
transform 1 0 25484 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_277
timestamp 1649977179
transform 1 0 26588 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_289
timestamp 1649977179
transform 1 0 27692 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_301
timestamp 1649977179
transform 1 0 28796 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_307
timestamp 1649977179
transform 1 0 29348 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_309
timestamp 1649977179
transform 1 0 29532 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_321
timestamp 1649977179
transform 1 0 30636 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_333
timestamp 1649977179
transform 1 0 31740 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_345
timestamp 1649977179
transform 1 0 32844 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_357
timestamp 1649977179
transform 1 0 33948 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_363
timestamp 1649977179
transform 1 0 34500 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_3
timestamp 1649977179
transform 1 0 1380 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_15
timestamp 1649977179
transform 1 0 2484 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_27
timestamp 1649977179
transform 1 0 3588 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_39
timestamp 1649977179
transform 1 0 4692 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_51
timestamp 1649977179
transform 1 0 5796 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_55
timestamp 1649977179
transform 1 0 6164 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_57
timestamp 1649977179
transform 1 0 6348 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_81
timestamp 1649977179
transform 1 0 8556 0 -1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_25_87
timestamp 1649977179
transform 1 0 9108 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_99
timestamp 1649977179
transform 1 0 10212 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_25_111
timestamp 1649977179
transform 1 0 11316 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_113
timestamp 1649977179
transform 1 0 11500 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_125
timestamp 1649977179
transform 1 0 12604 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_137
timestamp 1649977179
transform 1 0 13708 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_25_149
timestamp 1649977179
transform 1 0 14812 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_25_154
timestamp 1649977179
transform 1 0 15272 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_25_166
timestamp 1649977179
transform 1 0 16376 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_25_169
timestamp 1649977179
transform 1 0 16652 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_181
timestamp 1649977179
transform 1 0 17756 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_193
timestamp 1649977179
transform 1 0 18860 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_205
timestamp 1649977179
transform 1 0 19964 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_213
timestamp 1649977179
transform 1 0 20700 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_25_217
timestamp 1649977179
transform 1 0 21068 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_223
timestamp 1649977179
transform 1 0 21620 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_234
timestamp 1649977179
transform 1 0 22632 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_246
timestamp 1649977179
transform 1 0 23736 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_258
timestamp 1649977179
transform 1 0 24840 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_270
timestamp 1649977179
transform 1 0 25944 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_278
timestamp 1649977179
transform 1 0 26680 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_25_281
timestamp 1649977179
transform 1 0 26956 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_289
timestamp 1649977179
transform 1 0 27692 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_300
timestamp 1649977179
transform 1 0 28704 0 -1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_25_307
timestamp 1649977179
transform 1 0 29348 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_319
timestamp 1649977179
transform 1 0 30452 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_331
timestamp 1649977179
transform 1 0 31556 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_335
timestamp 1649977179
transform 1 0 31924 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_337
timestamp 1649977179
transform 1 0 32108 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_349
timestamp 1649977179
transform 1 0 33212 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_25_361
timestamp 1649977179
transform 1 0 34316 0 -1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_26_5
timestamp 1649977179
transform 1 0 1564 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_17
timestamp 1649977179
transform 1 0 2668 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_26_25
timestamp 1649977179
transform 1 0 3404 0 1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_26_29
timestamp 1649977179
transform 1 0 3772 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_41
timestamp 1649977179
transform 1 0 4876 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_53
timestamp 1649977179
transform 1 0 5980 0 1 16320
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_26_62
timestamp 1649977179
transform 1 0 6808 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_74
timestamp 1649977179
transform 1 0 7912 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_82
timestamp 1649977179
transform 1 0 8648 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_26_85
timestamp 1649977179
transform 1 0 8924 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_97
timestamp 1649977179
transform 1 0 10028 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_109
timestamp 1649977179
transform 1 0 11132 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_121
timestamp 1649977179
transform 1 0 12236 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_133
timestamp 1649977179
transform 1 0 13340 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_139
timestamp 1649977179
transform 1 0 13892 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_141
timestamp 1649977179
transform 1 0 14076 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_153
timestamp 1649977179
transform 1 0 15180 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_165
timestamp 1649977179
transform 1 0 16284 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_177
timestamp 1649977179
transform 1 0 17388 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_189
timestamp 1649977179
transform 1 0 18492 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_195
timestamp 1649977179
transform 1 0 19044 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_197
timestamp 1649977179
transform 1 0 19228 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_209
timestamp 1649977179
transform 1 0 20332 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_221
timestamp 1649977179
transform 1 0 21436 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_233
timestamp 1649977179
transform 1 0 22540 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_245
timestamp 1649977179
transform 1 0 23644 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_251
timestamp 1649977179
transform 1 0 24196 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_253
timestamp 1649977179
transform 1 0 24380 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_265
timestamp 1649977179
transform 1 0 25484 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_277
timestamp 1649977179
transform 1 0 26588 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_289
timestamp 1649977179
transform 1 0 27692 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_301
timestamp 1649977179
transform 1 0 28796 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_307
timestamp 1649977179
transform 1 0 29348 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_309
timestamp 1649977179
transform 1 0 29532 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_321
timestamp 1649977179
transform 1 0 30636 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_333
timestamp 1649977179
transform 1 0 31740 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_345
timestamp 1649977179
transform 1 0 32844 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_26_353
timestamp 1649977179
transform 1 0 33580 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_26_360
timestamp 1649977179
transform 1 0 34224 0 1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_27_13
timestamp 1649977179
transform 1 0 2300 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_27_25
timestamp 1649977179
transform 1 0 3404 0 -1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_27_33
timestamp 1649977179
transform 1 0 4140 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_45
timestamp 1649977179
transform 1 0 5244 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_27_53
timestamp 1649977179
transform 1 0 5980 0 -1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_27_57
timestamp 1649977179
transform 1 0 6348 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_69
timestamp 1649977179
transform 1 0 7452 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_27_81
timestamp 1649977179
transform 1 0 8556 0 -1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_27_85
timestamp 1649977179
transform 1 0 8924 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_97
timestamp 1649977179
transform 1 0 10028 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_27_109
timestamp 1649977179
transform 1 0 11132 0 -1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_27_117
timestamp 1649977179
transform 1 0 11868 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_129
timestamp 1649977179
transform 1 0 12972 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_27_137
timestamp 1649977179
transform 1 0 13708 0 -1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_27_141
timestamp 1649977179
transform 1 0 14076 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_153
timestamp 1649977179
transform 1 0 15180 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_27_165
timestamp 1649977179
transform 1 0 16284 0 -1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_27_169
timestamp 1649977179
transform 1 0 16652 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_27_181
timestamp 1649977179
transform 1 0 17756 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_27_188
timestamp 1649977179
transform 1 0 18400 0 -1 17408
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_27_197
timestamp 1649977179
transform 1 0 19228 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_209
timestamp 1649977179
transform 1 0 20332 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_27_221
timestamp 1649977179
transform 1 0 21436 0 -1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_27_225
timestamp 1649977179
transform 1 0 21804 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_237
timestamp 1649977179
transform 1 0 22908 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_27_249
timestamp 1649977179
transform 1 0 24012 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_27_253
timestamp 1649977179
transform 1 0 24380 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_261
timestamp 1649977179
transform 1 0 25116 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_266
timestamp 1649977179
transform 1 0 25576 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_27_278
timestamp 1649977179
transform 1 0 26680 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_27_281
timestamp 1649977179
transform 1 0 26956 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_293
timestamp 1649977179
transform 1 0 28060 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_27_305
timestamp 1649977179
transform 1 0 29164 0 -1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_27_309
timestamp 1649977179
transform 1 0 29532 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_321
timestamp 1649977179
transform 1 0 30636 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_27_333
timestamp 1649977179
transform 1 0 31740 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_27_337
timestamp 1649977179
transform 1 0 32108 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_27_344
timestamp 1649977179
transform 1 0 32752 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_27_352
timestamp 1649977179
transform 1 0 33488 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_360
timestamp 1649977179
transform 1 0 34224 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1649977179
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1649977179
transform -1 0 34868 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1649977179
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1649977179
transform -1 0 34868 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1649977179
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1649977179
transform -1 0 34868 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1649977179
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1649977179
transform -1 0 34868 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1649977179
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1649977179
transform -1 0 34868 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1649977179
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1649977179
transform -1 0 34868 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1649977179
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1649977179
transform -1 0 34868 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1649977179
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1649977179
transform -1 0 34868 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1649977179
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1649977179
transform -1 0 34868 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1649977179
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1649977179
transform -1 0 34868 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1649977179
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1649977179
transform -1 0 34868 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1649977179
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1649977179
transform -1 0 34868 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1649977179
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1649977179
transform -1 0 34868 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1649977179
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1649977179
transform -1 0 34868 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1649977179
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1649977179
transform -1 0 34868 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1649977179
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1649977179
transform -1 0 34868 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1649977179
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1649977179
transform -1 0 34868 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1649977179
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1649977179
transform -1 0 34868 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1649977179
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1649977179
transform -1 0 34868 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1649977179
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1649977179
transform -1 0 34868 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1649977179
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1649977179
transform -1 0 34868 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1649977179
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1649977179
transform -1 0 34868 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1649977179
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1649977179
transform -1 0 34868 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1649977179
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1649977179
transform -1 0 34868 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1649977179
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1649977179
transform -1 0 34868 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1649977179
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1649977179
transform -1 0 34868 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1649977179
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1649977179
transform -1 0 34868 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1649977179
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1649977179
transform -1 0 34868 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_56 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_57
timestamp 1649977179
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_58
timestamp 1649977179
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_59
timestamp 1649977179
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_60
timestamp 1649977179
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_61
timestamp 1649977179
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_62
timestamp 1649977179
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_63
timestamp 1649977179
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_64
timestamp 1649977179
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_65
timestamp 1649977179
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_66
timestamp 1649977179
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_67
timestamp 1649977179
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_68
timestamp 1649977179
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_69
timestamp 1649977179
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_70
timestamp 1649977179
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_71
timestamp 1649977179
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_72
timestamp 1649977179
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_73
timestamp 1649977179
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_74
timestamp 1649977179
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_75
timestamp 1649977179
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_76
timestamp 1649977179
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_77
timestamp 1649977179
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_78
timestamp 1649977179
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_79
timestamp 1649977179
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_80
timestamp 1649977179
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_81
timestamp 1649977179
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_82
timestamp 1649977179
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_83
timestamp 1649977179
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_84
timestamp 1649977179
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_85
timestamp 1649977179
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_86
timestamp 1649977179
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_87
timestamp 1649977179
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_88
timestamp 1649977179
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_89
timestamp 1649977179
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_90
timestamp 1649977179
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_91
timestamp 1649977179
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_92
timestamp 1649977179
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_93
timestamp 1649977179
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_94
timestamp 1649977179
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_95
timestamp 1649977179
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_96
timestamp 1649977179
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_97
timestamp 1649977179
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_98
timestamp 1649977179
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_99
timestamp 1649977179
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_100
timestamp 1649977179
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_101
timestamp 1649977179
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_102
timestamp 1649977179
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_103
timestamp 1649977179
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_104
timestamp 1649977179
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_105
timestamp 1649977179
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_106
timestamp 1649977179
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_107
timestamp 1649977179
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_108
timestamp 1649977179
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_109
timestamp 1649977179
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_110
timestamp 1649977179
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_111
timestamp 1649977179
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_112
timestamp 1649977179
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_113
timestamp 1649977179
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_114
timestamp 1649977179
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_115
timestamp 1649977179
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_116
timestamp 1649977179
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_117
timestamp 1649977179
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_118
timestamp 1649977179
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_119
timestamp 1649977179
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_120
timestamp 1649977179
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_121
timestamp 1649977179
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_122
timestamp 1649977179
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_123
timestamp 1649977179
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_124
timestamp 1649977179
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_125
timestamp 1649977179
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_126
timestamp 1649977179
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_127
timestamp 1649977179
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_128
timestamp 1649977179
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_129
timestamp 1649977179
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130
timestamp 1649977179
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 1649977179
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 1649977179
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 1649977179
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 1649977179
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1649977179
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1649977179
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1649977179
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1649977179
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1649977179
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1649977179
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1649977179
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1649977179
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1649977179
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1649977179
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1649977179
transform 1 0 32016 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1649977179
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1649977179
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1649977179
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1649977179
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1649977179
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1649977179
transform 1 0 29440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1649977179
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1649977179
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1649977179
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1649977179
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1649977179
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1649977179
transform 1 0 32016 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1649977179
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1649977179
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1649977179
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1649977179
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1649977179
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1649977179
transform 1 0 29440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1649977179
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1649977179
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1649977179
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1649977179
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1649977179
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1649977179
transform 1 0 32016 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1649977179
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1649977179
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1649977179
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1649977179
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1649977179
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1649977179
transform 1 0 29440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1649977179
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1649977179
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1649977179
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1649977179
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1649977179
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1649977179
transform 1 0 32016 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1649977179
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1649977179
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1649977179
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1649977179
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1649977179
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1649977179
transform 1 0 29440 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1649977179
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1649977179
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1649977179
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1649977179
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1649977179
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1649977179
transform 1 0 32016 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1649977179
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1649977179
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1649977179
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1649977179
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1649977179
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1649977179
transform 1 0 29440 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1649977179
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1649977179
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1649977179
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1649977179
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1649977179
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1649977179
transform 1 0 32016 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1649977179
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1649977179
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1649977179
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1649977179
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1649977179
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1649977179
transform 1 0 29440 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1649977179
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1649977179
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1649977179
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1649977179
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1649977179
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1649977179
transform 1 0 32016 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1649977179
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1649977179
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1649977179
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1649977179
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1649977179
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1649977179
transform 1 0 29440 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1649977179
transform 1 0 3680 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1649977179
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1649977179
transform 1 0 8832 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1649977179
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1649977179
transform 1 0 13984 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1649977179
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1649977179
transform 1 0 19136 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1649977179
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1649977179
transform 1 0 24288 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1649977179
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1649977179
transform 1 0 29440 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1649977179
transform 1 0 32016 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__and3b_1  _071_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 23184 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _072_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 23644 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _073_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 27784 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _074_
timestamp 1649977179
transform -1 0 27508 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _075_
timestamp 1649977179
transform 1 0 31004 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _076_
timestamp 1649977179
transform 1 0 29716 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _077_
timestamp 1649977179
transform 1 0 31004 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _078_
timestamp 1649977179
transform 1 0 29716 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _079_
timestamp 1649977179
transform -1 0 23000 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _080_
timestamp 1649977179
transform 1 0 21712 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_2  _081_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 6348 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _082_
timestamp 1649977179
transform 1 0 20700 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _083_
timestamp 1649977179
transform 1 0 19596 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _084_
timestamp 1649977179
transform 1 0 5980 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _085_
timestamp 1649977179
transform 1 0 4968 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _086_
timestamp 1649977179
transform 1 0 6440 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _087_
timestamp 1649977179
transform -1 0 6808 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_2  _088_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 20700 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _089_
timestamp 1649977179
transform 1 0 20516 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _090_
timestamp 1649977179
transform 1 0 14996 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _091_
timestamp 1649977179
transform 1 0 21804 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _092_
timestamp 1649977179
transform 1 0 20792 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _093_
timestamp 1649977179
transform -1 0 28704 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _094_
timestamp 1649977179
transform 1 0 29072 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _095_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 31740 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _096_
timestamp 1649977179
transform 1 0 30728 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _097_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 11776 0 1 5440
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _098_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 6256 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _099_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 12236 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_2  _100_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 12328 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _101_
timestamp 1649977179
transform 1 0 11776 0 -1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__and2b_1  _102_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 15364 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _103_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 18308 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _104_
timestamp 1649977179
transform -1 0 20240 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _105_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 5980 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _106_
timestamp 1649977179
transform -1 0 14444 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _107_
timestamp 1649977179
transform 1 0 14536 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _108_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 21160 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__nand2b_2  _109_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 12236 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__or3b_1  _110_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 11408 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _111_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 19688 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _112_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 12696 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _113_
timestamp 1649977179
transform -1 0 13892 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _114_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 4968 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _115_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 12144 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _116_
timestamp 1649977179
transform -1 0 11776 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _117_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 12328 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _118_
timestamp 1649977179
transform 1 0 13616 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__o2111ai_2  _119_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 12144 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__o31ai_1  _120_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 12328 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _121_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 13064 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__o22a_1  _122_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 12144 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _123_
timestamp 1649977179
transform -1 0 11040 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _124_
timestamp 1649977179
transform 1 0 21896 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _125_
timestamp 1649977179
transform -1 0 28336 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _126_
timestamp 1649977179
transform 1 0 21436 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _127_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 20608 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _128_
timestamp 1649977179
transform -1 0 30636 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _129_
timestamp 1649977179
transform 1 0 24380 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _130_
timestamp 1649977179
transform -1 0 28796 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _131_
timestamp 1649977179
transform 1 0 19228 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _132_
timestamp 1649977179
transform 1 0 19504 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _133_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 4416 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _134_
timestamp 1649977179
transform -1 0 4784 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _135_
timestamp 1649977179
transform 1 0 4600 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _136_
timestamp 1649977179
transform -1 0 12880 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _137_
timestamp 1649977179
transform 1 0 4876 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _138_
timestamp 1649977179
transform 1 0 21620 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _139_
timestamp 1649977179
transform -1 0 6900 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _140_
timestamp 1649977179
transform 1 0 15088 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _141_
timestamp 1649977179
transform 1 0 14260 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _142_
timestamp 1649977179
transform -1 0 8096 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _143_
timestamp 1649977179
transform -1 0 6624 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _144_
timestamp 1649977179
transform -1 0 14352 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _145_
timestamp 1649977179
transform 1 0 28428 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _146_
timestamp 1649977179
transform 1 0 28428 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _147_
timestamp 1649977179
transform 1 0 28612 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__dlxtn_1  _148_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 29532 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _149_
timestamp 1649977179
transform 1 0 22908 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__dfrtp_1  _150_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 3496 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _151_
timestamp 1649977179
transform 1 0 3588 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _152_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 13616 0 1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _153_
timestamp 1649977179
transform 1 0 3956 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _154_
timestamp 1649977179
transform 1 0 28152 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _155_
timestamp 1649977179
transform 1 0 20332 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _156_
timestamp 1649977179
transform 1 0 14076 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _157_
timestamp 1649977179
transform 1 0 6716 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _158_
timestamp 1649977179
transform 1 0 4140 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _159_
timestamp 1649977179
transform -1 0 15272 0 -1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _160_
timestamp 1649977179
transform 1 0 28060 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _161_
timestamp 1649977179
transform 1 0 27968 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _162_
timestamp 1649977179
transform 1 0 27784 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dlxtp_1  _163_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 30728 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _164_
timestamp 1649977179
transform 1 0 19412 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _165_
timestamp 1649977179
transform 1 0 31372 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_2  _166_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 21712 0 1 8704
box -38 -48 1234 592
use sky130_fd_sc_hd__dlxtn_1  _167_
timestamp 1649977179
transform -1 0 21344 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _168_
timestamp 1649977179
transform 1 0 32108 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 15916 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_clk
timestamp 1649977179
transform -1 0 12236 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_clk
timestamp 1649977179
transform 1 0 18216 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__buf_2  input1
timestamp 1649977179
transform 1 0 1380 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input2
timestamp 1649977179
transform 1 0 1380 0 -1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input3
timestamp 1649977179
transform 1 0 1380 0 -1 17408
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1649977179
transform -1 0 9568 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1649977179
transform -1 0 4600 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1649977179
transform 1 0 6808 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input7
timestamp 1649977179
transform 1 0 1840 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output8
timestamp 1649977179
transform 1 0 33856 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output9
timestamp 1649977179
transform 1 0 33856 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output10
timestamp 1649977179
transform -1 0 14628 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output11
timestamp 1649977179
transform 1 0 21804 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output12
timestamp 1649977179
transform -1 0 29900 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output13
timestamp 1649977179
transform 1 0 33856 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output14
timestamp 1649977179
transform 1 0 33856 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output15
timestamp 1649977179
transform 1 0 33856 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output16
timestamp 1649977179
transform 1 0 11500 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output17
timestamp 1649977179
transform -1 0 4140 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output18
timestamp 1649977179
transform 1 0 33856 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output19
timestamp 1649977179
transform 1 0 32384 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output20
timestamp 1649977179
transform -1 0 25576 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output21
timestamp 1649977179
transform -1 0 18400 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output22
timestamp 1649977179
transform 1 0 33856 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output23
timestamp 1649977179
transform 1 0 33856 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  repeater24
timestamp 1649977179
transform 1 0 20240 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  rlbp_25 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 33212 0 1 2176
box -38 -48 314 592
<< labels >>
flabel metal3 s 0 7488 800 7608 0 FreeSans 480 0 0 0 ce_d1
port 0 nsew signal input
flabel metal3 s 0 12384 800 12504 0 FreeSans 480 0 0 0 ce_d2
port 1 nsew signal input
flabel metal3 s 0 17280 800 17400 0 FreeSans 480 0 0 0 ce_d3
port 2 nsew signal input
flabel metal3 s 0 2592 800 2712 0 FreeSans 480 0 0 0 clk
port 3 nsew signal input
flabel metal3 s 35200 1368 36000 1488 0 FreeSans 480 0 0 0 control_signals[0]
port 4 nsew signal tristate
flabel metal3 s 35200 3816 36000 3936 0 FreeSans 480 0 0 0 control_signals[1]
port 5 nsew signal tristate
flabel metal2 s 11702 0 11758 800 0 FreeSans 224 90 0 0 d[0]
port 6 nsew signal input
flabel metal2 s 19154 0 19210 800 0 FreeSans 224 90 0 0 d[1]
port 7 nsew signal input
flabel metal2 s 26606 0 26662 800 0 FreeSans 224 90 0 0 d[2]
port 8 nsew signal input
flabel metal2 s 31574 0 31630 800 0 FreeSans 224 90 0 0 d[3]
port 9 nsew signal input
flabel metal2 s 9218 0 9274 800 0 FreeSans 224 90 0 0 data_in
port 10 nsew signal input
flabel metal2 s 14186 0 14242 800 0 FreeSans 224 90 0 0 data_out[0]
port 11 nsew signal tristate
flabel metal2 s 21638 0 21694 800 0 FreeSans 224 90 0 0 data_out[1]
port 12 nsew signal tristate
flabel metal2 s 29090 0 29146 800 0 FreeSans 224 90 0 0 data_out[2]
port 13 nsew signal tristate
flabel metal2 s 34058 0 34114 800 0 FreeSans 224 90 0 0 data_out[3]
port 14 nsew signal tristate
flabel metal2 s 16670 0 16726 800 0 FreeSans 224 90 0 0 data_sel[0]
port 15 nsew signal input
flabel metal2 s 24122 0 24178 800 0 FreeSans 224 90 0 0 data_sel[1]
port 16 nsew signal input
flabel metal2 s 4250 0 4306 800 0 FreeSans 224 90 0 0 gpio_start
port 17 nsew signal input
flabel metal2 s 6734 0 6790 800 0 FreeSans 224 90 0 0 logic_analyzer_start
port 18 nsew signal input
flabel metal3 s 35200 16056 36000 16176 0 FreeSans 480 0 0 0 q1_1
port 19 nsew signal tristate
flabel metal3 s 35200 13608 36000 13728 0 FreeSans 480 0 0 0 q1_2
port 20 nsew signal tristate
flabel metal3 s 35200 11160 36000 11280 0 FreeSans 480 0 0 0 q1_3
port 21 nsew signal tristate
flabel metal2 s 10782 19200 10838 20000 0 FreeSans 224 90 0 0 q2_1
port 22 nsew signal tristate
flabel metal2 s 3606 19200 3662 20000 0 FreeSans 224 90 0 0 q2_2
port 23 nsew signal tristate
flabel metal3 s 35200 18504 36000 18624 0 FreeSans 480 0 0 0 q2_3
port 24 nsew signal tristate
flabel metal2 s 32310 19200 32366 20000 0 FreeSans 224 90 0 0 q3_1
port 25 nsew signal tristate
flabel metal2 s 25134 19200 25190 20000 0 FreeSans 224 90 0 0 q3_2
port 26 nsew signal tristate
flabel metal2 s 17958 19200 18014 20000 0 FreeSans 224 90 0 0 q3_3
port 27 nsew signal tristate
flabel metal2 s 1766 0 1822 800 0 FreeSans 224 90 0 0 reset
port 28 nsew signal input
flabel metal3 s 35200 6264 36000 6384 0 FreeSans 480 0 0 0 reset_fsm
port 29 nsew signal tristate
flabel metal3 s 35200 8712 36000 8832 0 FreeSans 480 0 0 0 rlbp_done
port 30 nsew signal tristate
flabel metal4 s 5168 2128 5488 17456 0 FreeSans 1920 90 0 0 vccd1
port 31 nsew power bidirectional
flabel metal4 s 13616 2128 13936 17456 0 FreeSans 1920 90 0 0 vccd1
port 31 nsew power bidirectional
flabel metal4 s 22064 2128 22384 17456 0 FreeSans 1920 90 0 0 vccd1
port 31 nsew power bidirectional
flabel metal4 s 30512 2128 30832 17456 0 FreeSans 1920 90 0 0 vccd1
port 31 nsew power bidirectional
flabel metal4 s 9392 2128 9712 17456 0 FreeSans 1920 90 0 0 vssd1
port 32 nsew ground bidirectional
flabel metal4 s 17840 2128 18160 17456 0 FreeSans 1920 90 0 0 vssd1
port 32 nsew ground bidirectional
flabel metal4 s 26288 2128 26608 17456 0 FreeSans 1920 90 0 0 vssd1
port 32 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 36000 20000
<< end >>
