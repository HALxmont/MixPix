magic
tech sky130B
magscale 1 2
timestamp 1662148786
<< obsli1 >>
rect 1104 2159 34868 17425
<< obsm1 >>
rect 1104 2128 34868 17456
<< metal2 >>
rect 3606 19200 3662 20000
rect 10782 19200 10838 20000
rect 17958 19200 18014 20000
rect 25134 19200 25190 20000
rect 32310 19200 32366 20000
rect 1766 0 1822 800
rect 4250 0 4306 800
rect 6734 0 6790 800
rect 9218 0 9274 800
rect 11702 0 11758 800
rect 14186 0 14242 800
rect 16670 0 16726 800
rect 19154 0 19210 800
rect 21638 0 21694 800
rect 24122 0 24178 800
rect 26606 0 26662 800
rect 29090 0 29146 800
rect 31574 0 31630 800
rect 34058 0 34114 800
<< obsm2 >>
rect 1398 19144 3550 19258
rect 3718 19144 10726 19258
rect 10894 19144 17902 19258
rect 18070 19144 25078 19258
rect 25246 19144 32254 19258
rect 32422 19144 34114 19258
rect 1398 856 34114 19144
rect 1398 800 1710 856
rect 1878 800 4194 856
rect 4362 800 6678 856
rect 6846 800 9162 856
rect 9330 800 11646 856
rect 11814 800 14130 856
rect 14298 800 16614 856
rect 16782 800 19098 856
rect 19266 800 21582 856
rect 21750 800 24066 856
rect 24234 800 26550 856
rect 26718 800 29034 856
rect 29202 800 31518 856
rect 31686 800 34002 856
<< metal3 >>
rect 35200 18504 36000 18624
rect 0 17280 800 17400
rect 35200 16056 36000 16176
rect 35200 13608 36000 13728
rect 0 12384 800 12504
rect 35200 11160 36000 11280
rect 35200 8712 36000 8832
rect 0 7488 800 7608
rect 35200 6264 36000 6384
rect 35200 3816 36000 3936
rect 0 2592 800 2712
rect 35200 1368 36000 1488
<< obsm3 >>
rect 800 18424 35120 18597
rect 800 17480 35200 18424
rect 880 17200 35200 17480
rect 800 16256 35200 17200
rect 800 15976 35120 16256
rect 800 13808 35200 15976
rect 800 13528 35120 13808
rect 800 12584 35200 13528
rect 880 12304 35200 12584
rect 800 11360 35200 12304
rect 800 11080 35120 11360
rect 800 8912 35200 11080
rect 800 8632 35120 8912
rect 800 7688 35200 8632
rect 880 7408 35200 7688
rect 800 6464 35200 7408
rect 800 6184 35120 6464
rect 800 4016 35200 6184
rect 800 3736 35120 4016
rect 800 2792 35200 3736
rect 880 2512 35200 2792
rect 800 1568 35200 2512
rect 800 1395 35120 1568
<< metal4 >>
rect 5168 2128 5488 17456
rect 9392 2128 9712 17456
rect 13616 2128 13936 17456
rect 17840 2128 18160 17456
rect 22064 2128 22384 17456
rect 26288 2128 26608 17456
rect 30512 2128 30832 17456
<< labels >>
rlabel metal3 s 0 7488 800 7608 6 ce_d1
port 1 nsew signal input
rlabel metal3 s 0 12384 800 12504 6 ce_d2
port 2 nsew signal input
rlabel metal3 s 0 17280 800 17400 6 ce_d3
port 3 nsew signal input
rlabel metal3 s 0 2592 800 2712 6 clk
port 4 nsew signal input
rlabel metal3 s 35200 1368 36000 1488 6 control_signals[0]
port 5 nsew signal output
rlabel metal3 s 35200 3816 36000 3936 6 control_signals[1]
port 6 nsew signal output
rlabel metal2 s 11702 0 11758 800 6 d[0]
port 7 nsew signal input
rlabel metal2 s 19154 0 19210 800 6 d[1]
port 8 nsew signal input
rlabel metal2 s 26606 0 26662 800 6 d[2]
port 9 nsew signal input
rlabel metal2 s 31574 0 31630 800 6 d[3]
port 10 nsew signal input
rlabel metal2 s 9218 0 9274 800 6 data_in
port 11 nsew signal input
rlabel metal2 s 14186 0 14242 800 6 data_out[0]
port 12 nsew signal output
rlabel metal2 s 21638 0 21694 800 6 data_out[1]
port 13 nsew signal output
rlabel metal2 s 29090 0 29146 800 6 data_out[2]
port 14 nsew signal output
rlabel metal2 s 34058 0 34114 800 6 data_out[3]
port 15 nsew signal output
rlabel metal2 s 16670 0 16726 800 6 data_sel[0]
port 16 nsew signal input
rlabel metal2 s 24122 0 24178 800 6 data_sel[1]
port 17 nsew signal input
rlabel metal2 s 4250 0 4306 800 6 gpio_start
port 18 nsew signal input
rlabel metal2 s 6734 0 6790 800 6 logic_analyzer_start
port 19 nsew signal input
rlabel metal3 s 35200 16056 36000 16176 6 q1_1
port 20 nsew signal output
rlabel metal3 s 35200 13608 36000 13728 6 q1_2
port 21 nsew signal output
rlabel metal3 s 35200 11160 36000 11280 6 q1_3
port 22 nsew signal output
rlabel metal2 s 10782 19200 10838 20000 6 q2_1
port 23 nsew signal output
rlabel metal2 s 3606 19200 3662 20000 6 q2_2
port 24 nsew signal output
rlabel metal3 s 35200 18504 36000 18624 6 q2_3
port 25 nsew signal output
rlabel metal2 s 32310 19200 32366 20000 6 q3_1
port 26 nsew signal output
rlabel metal2 s 25134 19200 25190 20000 6 q3_2
port 27 nsew signal output
rlabel metal2 s 17958 19200 18014 20000 6 q3_3
port 28 nsew signal output
rlabel metal2 s 1766 0 1822 800 6 reset
port 29 nsew signal input
rlabel metal3 s 35200 6264 36000 6384 6 reset_fsm
port 30 nsew signal output
rlabel metal3 s 35200 8712 36000 8832 6 rlbp_done
port 31 nsew signal output
rlabel metal4 s 5168 2128 5488 17456 6 vccd1
port 32 nsew power bidirectional
rlabel metal4 s 13616 2128 13936 17456 6 vccd1
port 32 nsew power bidirectional
rlabel metal4 s 22064 2128 22384 17456 6 vccd1
port 32 nsew power bidirectional
rlabel metal4 s 30512 2128 30832 17456 6 vccd1
port 32 nsew power bidirectional
rlabel metal4 s 9392 2128 9712 17456 6 vssd1
port 33 nsew ground bidirectional
rlabel metal4 s 17840 2128 18160 17456 6 vssd1
port 33 nsew ground bidirectional
rlabel metal4 s 26288 2128 26608 17456 6 vssd1
port 33 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 36000 20000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 702856
string GDS_FILE /home/mxmont/Documents/Universidad/IC-UBB/MixPix/CARAVEL_WRAPPER/MixPix/openlane/rlbp/runs/22_09_02_15_58/results/signoff/rlbp.magic.gds
string GDS_START 253776
<< end >>

