magic
tech sky130B
magscale 1 2
timestamp 1667009656
<< metal1 >>
rect 30374 702992 30380 703044
rect 30432 703032 30438 703044
rect 31570 703032 31576 703044
rect 30432 703004 31576 703032
rect 30432 702992 30438 703004
rect 31570 702992 31576 703004
rect 31628 702992 31634 703044
rect 405734 702992 405740 703044
rect 405792 703032 405798 703044
rect 407022 703032 407028 703044
rect 405792 703004 407028 703032
rect 405792 702992 405798 703004
rect 407022 702992 407028 703004
rect 407080 702992 407086 703044
rect 425054 702992 425060 703044
rect 425112 703032 425118 703044
rect 426342 703032 426348 703044
rect 425112 703004 426348 703032
rect 425112 702992 425118 703004
rect 426342 702992 426348 703004
rect 426400 702992 426406 703044
rect 436094 702992 436100 703044
rect 436152 703032 436158 703044
rect 437290 703032 437296 703044
rect 436152 703004 437296 703032
rect 436152 702992 436158 703004
rect 437290 702992 437296 703004
rect 437348 702992 437354 703044
rect 455414 702992 455420 703044
rect 455472 703032 455478 703044
rect 456610 703032 456616 703044
rect 455472 703004 456616 703032
rect 455472 702992 455478 703004
rect 456610 702992 456616 703004
rect 456668 702992 456674 703044
rect 544378 702448 544384 702500
rect 544436 702488 544442 702500
rect 580166 702488 580172 702500
rect 544436 702460 580172 702488
rect 544436 702448 544442 702460
rect 580166 702448 580172 702460
rect 580224 702448 580230 702500
rect 3418 701020 3424 701072
rect 3476 701060 3482 701072
rect 131114 701060 131120 701072
rect 3476 701032 131120 701060
rect 3476 701020 3482 701032
rect 131114 701020 131120 701032
rect 131172 701020 131178 701072
rect 88242 700680 88248 700732
rect 88300 700720 88306 700732
rect 102778 700720 102784 700732
rect 88300 700692 102784 700720
rect 88300 700680 88306 700692
rect 102778 700680 102784 700692
rect 102836 700680 102842 700732
rect 65702 700612 65708 700664
rect 65760 700652 65766 700664
rect 79318 700652 79324 700664
rect 65760 700624 79324 700652
rect 65760 700612 65766 700624
rect 79318 700612 79324 700624
rect 79376 700612 79382 700664
rect 80514 700612 80520 700664
rect 80572 700652 80578 700664
rect 88978 700652 88984 700664
rect 80572 700624 88984 700652
rect 80572 700612 80578 700624
rect 88978 700612 88984 700624
rect 89036 700612 89042 700664
rect 95970 700612 95976 700664
rect 96028 700652 96034 700664
rect 122834 700652 122840 700664
rect 96028 700624 122840 700652
rect 96028 700612 96034 700624
rect 122834 700612 122840 700624
rect 122892 700612 122898 700664
rect 4522 700544 4528 700596
rect 4580 700584 4586 700596
rect 26878 700584 26884 700596
rect 4580 700556 26884 700584
rect 4580 700544 4586 700556
rect 26878 700544 26884 700556
rect 26936 700544 26942 700596
rect 46382 700544 46388 700596
rect 46440 700584 46446 700596
rect 98730 700584 98736 700596
rect 46440 700556 98736 700584
rect 46440 700544 46446 700556
rect 98730 700544 98736 700556
rect 98788 700544 98794 700596
rect 179046 700544 179052 700596
rect 179104 700584 179110 700596
rect 189534 700584 189540 700596
rect 179104 700556 189540 700584
rect 179104 700544 179110 700556
rect 189534 700544 189540 700556
rect 189592 700544 189598 700596
rect 19978 700476 19984 700528
rect 20036 700516 20042 700528
rect 48958 700516 48964 700528
rect 20036 700488 48964 700516
rect 20036 700476 20042 700488
rect 48958 700476 48964 700488
rect 49016 700476 49022 700528
rect 54110 700476 54116 700528
rect 54168 700516 54174 700528
rect 117958 700516 117964 700528
rect 54168 700488 117964 700516
rect 54168 700476 54174 700488
rect 117958 700476 117964 700488
rect 118016 700476 118022 700528
rect 133966 700476 133972 700528
rect 134024 700516 134030 700528
rect 149698 700516 149704 700528
rect 134024 700488 149704 700516
rect 134024 700476 134030 700488
rect 149698 700476 149704 700488
rect 149756 700476 149762 700528
rect 168098 700476 168104 700528
rect 168156 700516 168162 700528
rect 191834 700516 191840 700528
rect 168156 700488 191840 700516
rect 168156 700476 168162 700488
rect 191834 700476 191840 700488
rect 191892 700476 191898 700528
rect 23842 700408 23848 700460
rect 23900 700448 23906 700460
rect 109034 700448 109040 700460
rect 23900 700420 109040 700448
rect 23900 700408 23906 700420
rect 109034 700408 109040 700420
rect 109092 700408 109098 700460
rect 117222 700408 117228 700460
rect 117280 700448 117286 700460
rect 137830 700448 137836 700460
rect 117280 700420 137836 700448
rect 117280 700408 117286 700420
rect 137830 700408 137836 700420
rect 137888 700408 137894 700460
rect 164234 700408 164240 700460
rect 164292 700448 164298 700460
rect 193214 700448 193220 700460
rect 164292 700420 193220 700448
rect 164292 700408 164298 700420
rect 193214 700408 193220 700420
rect 193272 700408 193278 700460
rect 542998 700408 543004 700460
rect 543056 700448 543062 700460
rect 574462 700448 574468 700460
rect 543056 700420 574468 700448
rect 543056 700408 543062 700420
rect 574462 700408 574468 700420
rect 574520 700408 574526 700460
rect 12250 700340 12256 700392
rect 12308 700380 12314 700392
rect 100110 700380 100116 700392
rect 12308 700352 100116 700380
rect 12308 700340 12314 700352
rect 100110 700340 100116 700352
rect 100168 700340 100174 700392
rect 115842 700340 115848 700392
rect 115900 700380 115906 700392
rect 141694 700380 141700 700392
rect 115900 700352 141700 700380
rect 115900 700340 115906 700352
rect 141694 700340 141700 700352
rect 141752 700340 141758 700392
rect 175826 700340 175832 700392
rect 175884 700380 175890 700392
rect 189442 700380 189448 700392
rect 175884 700352 189448 700380
rect 175884 700340 175890 700352
rect 189442 700340 189448 700352
rect 189500 700340 189506 700392
rect 189718 700340 189724 700392
rect 189776 700380 189782 700392
rect 244090 700380 244096 700392
rect 189776 700352 244096 700380
rect 189776 700340 189782 700352
rect 244090 700340 244096 700352
rect 244148 700340 244154 700392
rect 514018 700340 514024 700392
rect 514076 700380 514082 700392
rect 566734 700380 566740 700392
rect 514076 700352 566740 700380
rect 514076 700340 514082 700352
rect 566734 700340 566740 700352
rect 566792 700340 566798 700392
rect 658 700272 664 700324
rect 716 700312 722 700324
rect 100018 700312 100024 700324
rect 716 700284 100024 700312
rect 716 700272 722 700284
rect 100018 700272 100024 700284
rect 100076 700272 100082 700324
rect 120718 700272 120724 700324
rect 120776 700312 120782 700324
rect 198366 700312 198372 700324
rect 120776 700284 198372 700312
rect 120776 700272 120782 700284
rect 198366 700272 198372 700284
rect 198424 700272 198430 700324
rect 239398 700272 239404 700324
rect 239456 700312 239462 700324
rect 555142 700312 555148 700324
rect 239456 700284 555148 700312
rect 239456 700272 239462 700284
rect 555142 700272 555148 700284
rect 555200 700272 555206 700324
rect 190638 699728 190644 699780
rect 190696 699768 190702 699780
rect 195974 699768 195980 699780
rect 190696 699740 195980 699768
rect 190696 699728 190702 699740
rect 195974 699728 195980 699740
rect 196032 699728 196038 699780
rect 42518 699660 42524 699712
rect 42576 699700 42582 699712
rect 43438 699700 43444 699712
rect 42576 699672 43444 699700
rect 42576 699660 42582 699672
rect 43438 699660 43444 699672
rect 43496 699660 43502 699712
rect 144178 699660 144184 699712
rect 144236 699700 144242 699712
rect 144914 699700 144920 699712
rect 144236 699672 144920 699700
rect 144236 699660 144242 699672
rect 144914 699660 144920 699672
rect 144972 699660 144978 699712
rect 192478 699660 192484 699712
rect 192536 699700 192542 699712
rect 194502 699700 194508 699712
rect 192536 699672 194508 699700
rect 192536 699660 192542 699672
rect 194502 699660 194508 699672
rect 194560 699660 194566 699712
rect 260098 699660 260104 699712
rect 260156 699700 260162 699712
rect 262766 699700 262772 699712
rect 260156 699672 262772 699700
rect 260156 699660 260162 699672
rect 262766 699660 262772 699672
rect 262824 699660 262830 699712
rect 305638 699660 305644 699712
rect 305696 699700 305702 699712
rect 308490 699700 308496 699712
rect 305696 699672 308496 699700
rect 305696 699660 305702 699672
rect 308490 699660 308496 699672
rect 308548 699660 308554 699712
rect 309778 699660 309784 699712
rect 309836 699700 309842 699712
rect 312354 699700 312360 699712
rect 309836 699672 312360 699700
rect 309836 699660 309842 699672
rect 312354 699660 312360 699672
rect 312412 699660 312418 699712
rect 313918 699660 313924 699712
rect 313976 699700 313982 699712
rect 316218 699700 316224 699712
rect 313976 699672 316224 699700
rect 313976 699660 313982 699672
rect 316218 699660 316224 699672
rect 316276 699660 316282 699712
rect 327718 699660 327724 699712
rect 327776 699700 327782 699712
rect 331030 699700 331036 699712
rect 327776 699672 331036 699700
rect 327776 699660 327782 699672
rect 331030 699660 331036 699672
rect 331088 699660 331094 699712
rect 359458 699660 359464 699712
rect 359516 699700 359522 699712
rect 361942 699700 361948 699712
rect 359516 699672 361948 699700
rect 359516 699660 359522 699672
rect 361942 699660 361948 699672
rect 362000 699660 362006 699712
rect 377398 699660 377404 699712
rect 377456 699700 377462 699712
rect 380618 699700 380624 699712
rect 377456 699672 380624 699700
rect 377456 699660 377462 699672
rect 380618 699660 380624 699672
rect 380676 699660 380682 699712
rect 381538 699660 381544 699712
rect 381596 699700 381602 699712
rect 384482 699700 384488 699712
rect 381596 699672 384488 699700
rect 381596 699660 381602 699672
rect 384482 699660 384488 699672
rect 384540 699660 384546 699712
rect 428458 699660 428464 699712
rect 428516 699700 428522 699712
rect 430206 699700 430212 699712
rect 428516 699672 430212 699700
rect 428516 699660 428522 699672
rect 430206 699660 430212 699672
rect 430264 699660 430270 699712
rect 431218 699660 431224 699712
rect 431276 699700 431282 699712
rect 434070 699700 434076 699712
rect 431276 699672 434076 699700
rect 431276 699660 431282 699672
rect 434070 699660 434076 699672
rect 434128 699660 434134 699712
rect 476758 699660 476764 699712
rect 476816 699700 476822 699712
rect 479150 699700 479156 699712
rect 476816 699672 479156 699700
rect 476816 699660 476822 699672
rect 479150 699660 479156 699672
rect 479208 699660 479214 699712
rect 548518 699660 548524 699712
rect 548576 699700 548582 699712
rect 551278 699700 551284 699712
rect 548576 699672 551284 699700
rect 548576 699660 548582 699672
rect 551278 699660 551284 699672
rect 551336 699660 551342 699712
rect 558178 699660 558184 699712
rect 558236 699700 558242 699712
rect 559006 699700 559012 699712
rect 558236 699672 559012 699700
rect 558236 699660 558242 699672
rect 559006 699660 559012 699672
rect 559064 699660 559070 699712
rect 16114 698912 16120 698964
rect 16172 698952 16178 698964
rect 62758 698952 62764 698964
rect 16172 698924 62764 698952
rect 16172 698912 16178 698924
rect 62758 698912 62764 698924
rect 62816 698912 62822 698964
rect 199378 698300 199384 698352
rect 199436 698340 199442 698352
rect 580166 698340 580172 698352
rect 199436 698312 580172 698340
rect 199436 698300 199442 698312
rect 580166 698300 580172 698312
rect 580224 698300 580230 698352
rect 67634 697552 67640 697604
rect 67692 697592 67698 697604
rect 68922 697592 68928 697604
rect 67692 697564 68928 697592
rect 67692 697552 67698 697564
rect 68922 697552 68928 697564
rect 68980 697552 68986 697604
rect 531314 697552 531320 697604
rect 531372 697592 531378 697604
rect 532602 697592 532608 697604
rect 531372 697564 532608 697592
rect 531372 697552 531378 697564
rect 532602 697552 532608 697564
rect 532660 697552 532666 697604
rect 3050 696940 3056 696992
rect 3108 696980 3114 696992
rect 98638 696980 98644 696992
rect 3108 696952 98644 696980
rect 3108 696940 3114 696952
rect 98638 696940 98644 696952
rect 98696 696940 98702 696992
rect 299474 696600 299480 696652
rect 299532 696640 299538 696652
rect 300762 696640 300768 696652
rect 299532 696612 300768 696640
rect 299532 696600 299538 696612
rect 300762 696600 300768 696612
rect 300820 696600 300826 696652
rect 511994 696600 512000 696652
rect 512052 696640 512058 696652
rect 513282 696640 513288 696652
rect 512052 696612 513288 696640
rect 512052 696600 512058 696612
rect 513282 696600 513288 696612
rect 513340 696600 513346 696652
rect 559558 694152 559564 694204
rect 559616 694192 559622 694204
rect 580166 694192 580172 694204
rect 559616 694164 580172 694192
rect 559616 694152 559622 694164
rect 580166 694152 580172 694164
rect 580224 694152 580230 694204
rect 552658 690004 552664 690056
rect 552716 690044 552722 690056
rect 580166 690044 580172 690056
rect 552716 690016 580172 690044
rect 552716 690004 552722 690016
rect 580166 690004 580172 690016
rect 580224 690004 580230 690056
rect 3418 688644 3424 688696
rect 3476 688684 3482 688696
rect 14458 688684 14464 688696
rect 3476 688656 14464 688684
rect 3476 688644 3482 688656
rect 14458 688644 14464 688656
rect 14516 688644 14522 688696
rect 556798 685856 556804 685908
rect 556856 685896 556862 685908
rect 579798 685896 579804 685908
rect 556856 685868 579804 685896
rect 556856 685856 556862 685868
rect 579798 685856 579804 685868
rect 579856 685856 579862 685908
rect 3142 684496 3148 684548
rect 3200 684536 3206 684548
rect 93118 684536 93124 684548
rect 3200 684508 93124 684536
rect 3200 684496 3206 684508
rect 93118 684496 93124 684508
rect 93176 684496 93182 684548
rect 552750 681708 552756 681760
rect 552808 681748 552814 681760
rect 580166 681748 580172 681760
rect 552808 681720 580172 681748
rect 552808 681708 552814 681720
rect 580166 681708 580172 681720
rect 580224 681708 580230 681760
rect 3418 680348 3424 680400
rect 3476 680388 3482 680400
rect 104158 680388 104164 680400
rect 3476 680360 104164 680388
rect 3476 680348 3482 680360
rect 104158 680348 104164 680360
rect 104216 680348 104222 680400
rect 566458 677560 566464 677612
rect 566516 677600 566522 677612
rect 580166 677600 580172 677612
rect 566516 677572 580172 677600
rect 566516 677560 566522 677572
rect 580166 677560 580172 677572
rect 580224 677560 580230 677612
rect 3418 676200 3424 676252
rect 3476 676240 3482 676252
rect 93302 676240 93308 676252
rect 3476 676212 93308 676240
rect 3476 676200 3482 676212
rect 93302 676200 93308 676212
rect 93360 676200 93366 676252
rect 200758 673480 200764 673532
rect 200816 673520 200822 673532
rect 580166 673520 580172 673532
rect 200816 673492 580172 673520
rect 200816 673480 200822 673492
rect 580166 673480 580172 673492
rect 580224 673480 580230 673532
rect 548610 669332 548616 669384
rect 548668 669372 548674 669384
rect 580166 669372 580172 669384
rect 548668 669344 580172 669372
rect 548668 669332 548674 669344
rect 580166 669332 580172 669344
rect 580224 669332 580230 669384
rect 3234 663756 3240 663808
rect 3292 663796 3298 663808
rect 112438 663796 112444 663808
rect 3292 663768 112444 663796
rect 3292 663756 3298 663768
rect 112438 663756 112444 663768
rect 112496 663756 112502 663808
rect 3418 661036 3424 661088
rect 3476 661076 3482 661088
rect 86218 661076 86224 661088
rect 3476 661048 86224 661076
rect 3476 661036 3482 661048
rect 86218 661036 86224 661048
rect 86276 661036 86282 661088
rect 541618 661036 541624 661088
rect 541676 661076 541682 661088
rect 580166 661076 580172 661088
rect 541676 661048 580172 661076
rect 541676 661036 541682 661048
rect 580166 661036 580172 661048
rect 580224 661036 580230 661088
rect 124306 658248 124312 658300
rect 124364 658288 124370 658300
rect 580166 658288 580172 658300
rect 124364 658260 580172 658288
rect 124364 658248 124370 658260
rect 580166 658248 580172 658260
rect 580224 658248 580230 658300
rect 566550 654100 566556 654152
rect 566608 654140 566614 654152
rect 580166 654140 580172 654152
rect 566608 654112 580172 654140
rect 566608 654100 566614 654112
rect 580166 654100 580172 654112
rect 580224 654100 580230 654152
rect 3050 652740 3056 652792
rect 3108 652780 3114 652792
rect 108298 652780 108304 652792
rect 3108 652752 108304 652780
rect 3108 652740 3114 652752
rect 108298 652740 108304 652752
rect 108356 652740 108362 652792
rect 179322 645872 179328 645924
rect 179380 645912 179386 645924
rect 580166 645912 580172 645924
rect 179380 645884 580172 645912
rect 179380 645872 179386 645884
rect 580166 645872 580172 645884
rect 580224 645872 580230 645924
rect 3418 644444 3424 644496
rect 3476 644484 3482 644496
rect 89070 644484 89076 644496
rect 3476 644456 89076 644484
rect 3476 644444 3482 644456
rect 89070 644444 89076 644456
rect 89128 644444 89134 644496
rect 558270 641724 558276 641776
rect 558328 641764 558334 641776
rect 580166 641764 580172 641776
rect 558328 641736 580172 641764
rect 558328 641724 558334 641736
rect 580166 641724 580172 641736
rect 580224 641724 580230 641776
rect 3142 640296 3148 640348
rect 3200 640336 3206 640348
rect 94498 640336 94504 640348
rect 3200 640308 94504 640336
rect 3200 640296 3206 640308
rect 94498 640296 94504 640308
rect 94556 640296 94562 640348
rect 3142 636216 3148 636268
rect 3200 636256 3206 636268
rect 13078 636256 13084 636268
rect 3200 636228 13084 636256
rect 3200 636216 3206 636228
rect 13078 636216 13084 636228
rect 13136 636216 13142 636268
rect 3418 632068 3424 632120
rect 3476 632108 3482 632120
rect 90358 632108 90364 632120
rect 3476 632080 90364 632108
rect 3476 632068 3482 632080
rect 90358 632068 90364 632080
rect 90416 632068 90422 632120
rect 570598 625132 570604 625184
rect 570656 625172 570662 625184
rect 580166 625172 580172 625184
rect 570656 625144 580172 625172
rect 570656 625132 570662 625144
rect 580166 625132 580172 625144
rect 580224 625132 580230 625184
rect 3234 623772 3240 623824
rect 3292 623812 3298 623824
rect 102870 623812 102876 623824
rect 3292 623784 102876 623812
rect 3292 623772 3298 623784
rect 102870 623772 102876 623784
rect 102928 623772 102934 623824
rect 3418 620984 3424 621036
rect 3476 621024 3482 621036
rect 104250 621024 104256 621036
rect 3476 620996 104256 621024
rect 3476 620984 3482 620996
rect 104250 620984 104256 620996
rect 104308 620984 104314 621036
rect 576118 620984 576124 621036
rect 576176 621024 576182 621036
rect 579798 621024 579804 621036
rect 576176 620996 579804 621024
rect 576176 620984 576182 620996
rect 579798 620984 579804 620996
rect 579856 620984 579862 621036
rect 3142 616836 3148 616888
rect 3200 616876 3206 616888
rect 21358 616876 21364 616888
rect 3200 616848 21364 616876
rect 3200 616836 3206 616848
rect 21358 616836 21364 616848
rect 21416 616836 21422 616888
rect 3142 612756 3148 612808
rect 3200 612796 3206 612808
rect 64138 612796 64144 612808
rect 3200 612768 64144 612796
rect 3200 612756 3206 612768
rect 64138 612756 64144 612768
rect 64196 612756 64202 612808
rect 120074 605820 120080 605872
rect 120132 605860 120138 605872
rect 580166 605860 580172 605872
rect 120132 605832 580172 605860
rect 120132 605820 120138 605832
rect 580166 605820 580172 605832
rect 580224 605820 580230 605872
rect 3050 604460 3056 604512
rect 3108 604500 3114 604512
rect 104342 604500 104348 604512
rect 3108 604472 104348 604500
rect 3108 604460 3114 604472
rect 104342 604460 104348 604472
rect 104400 604460 104406 604512
rect 560938 601672 560944 601724
rect 560996 601712 561002 601724
rect 580166 601712 580172 601724
rect 560996 601684 580172 601712
rect 560996 601672 561002 601684
rect 580166 601672 580172 601684
rect 580224 601672 580230 601724
rect 3510 600312 3516 600364
rect 3568 600352 3574 600364
rect 115934 600352 115940 600364
rect 3568 600324 115940 600352
rect 3568 600312 3574 600324
rect 115934 600312 115940 600324
rect 115992 600312 115998 600364
rect 3050 596164 3056 596216
rect 3108 596204 3114 596216
rect 104894 596204 104900 596216
rect 3108 596176 104900 596204
rect 3108 596164 3114 596176
rect 104894 596164 104900 596176
rect 104952 596164 104958 596216
rect 3142 592016 3148 592068
rect 3200 592056 3206 592068
rect 80698 592056 80704 592068
rect 3200 592028 80704 592056
rect 3200 592016 3206 592028
rect 80698 592016 80704 592028
rect 80756 592016 80762 592068
rect 574738 589296 574744 589348
rect 574796 589336 574802 589348
rect 580166 589336 580172 589348
rect 574796 589308 580172 589336
rect 574796 589296 574802 589308
rect 580166 589296 580172 589308
rect 580224 589296 580230 589348
rect 3234 587868 3240 587920
rect 3292 587908 3298 587920
rect 180794 587908 180800 587920
rect 3292 587880 180800 587908
rect 3292 587868 3298 587880
rect 180794 587868 180800 587880
rect 180852 587868 180858 587920
rect 3142 583720 3148 583772
rect 3200 583760 3206 583772
rect 84838 583760 84844 583772
rect 3200 583732 84844 583760
rect 3200 583720 3206 583732
rect 84838 583720 84844 583732
rect 84896 583720 84902 583772
rect 3326 581000 3332 581052
rect 3384 581040 3390 581052
rect 90450 581040 90456 581052
rect 3384 581012 90456 581040
rect 3384 581000 3390 581012
rect 90450 581000 90456 581012
rect 90508 581000 90514 581052
rect 3510 576852 3516 576904
rect 3568 576892 3574 576904
rect 80790 576892 80796 576904
rect 3568 576864 80796 576892
rect 3568 576852 3574 576864
rect 80790 576852 80796 576864
rect 80848 576852 80854 576904
rect 2866 568556 2872 568608
rect 2924 568596 2930 568608
rect 94590 568596 94596 568608
rect 2924 568568 94596 568596
rect 2924 568556 2930 568568
rect 94590 568556 94596 568568
rect 94648 568556 94654 568608
rect 562318 568556 562324 568608
rect 562376 568596 562382 568608
rect 580166 568596 580172 568608
rect 562376 568568 580172 568596
rect 562376 568556 562382 568568
rect 580166 568556 580172 568568
rect 580224 568556 580230 568608
rect 130378 565836 130384 565888
rect 130436 565876 130442 565888
rect 580166 565876 580172 565888
rect 130436 565848 580172 565876
rect 130436 565836 130442 565848
rect 580166 565836 580172 565848
rect 580224 565836 580230 565888
rect 3050 560260 3056 560312
rect 3108 560300 3114 560312
rect 106918 560300 106924 560312
rect 3108 560272 106924 560300
rect 3108 560260 3114 560272
rect 106918 560260 106924 560272
rect 106976 560260 106982 560312
rect 3050 556180 3056 556232
rect 3108 556220 3114 556232
rect 97258 556220 97264 556232
rect 3108 556192 97264 556220
rect 3108 556180 3114 556192
rect 97258 556180 97264 556192
rect 97316 556180 97322 556232
rect 576210 553392 576216 553444
rect 576268 553432 576274 553444
rect 580166 553432 580172 553444
rect 576268 553404 580172 553432
rect 576268 553392 576274 553404
rect 580166 553392 580172 553404
rect 580224 553392 580230 553444
rect 3510 552032 3516 552084
rect 3568 552072 3574 552084
rect 84930 552072 84936 552084
rect 3568 552044 84936 552072
rect 3568 552032 3574 552044
rect 84930 552032 84936 552044
rect 84988 552032 84994 552084
rect 571978 549244 571984 549296
rect 572036 549284 572042 549296
rect 580166 549284 580172 549296
rect 572036 549256 580172 549284
rect 572036 549244 572042 549256
rect 580166 549244 580172 549256
rect 580224 549244 580230 549296
rect 3050 547884 3056 547936
rect 3108 547924 3114 547936
rect 98822 547924 98828 547936
rect 3108 547896 98828 547924
rect 3108 547884 3114 547896
rect 98822 547884 98828 547896
rect 98880 547884 98886 547936
rect 558362 545096 558368 545148
rect 558420 545136 558426 545148
rect 579890 545136 579896 545148
rect 558420 545108 579896 545136
rect 558420 545096 558426 545108
rect 579890 545096 579896 545108
rect 579948 545096 579954 545148
rect 3142 543736 3148 543788
rect 3200 543776 3206 543788
rect 110506 543776 110512 543788
rect 3200 543748 110512 543776
rect 3200 543736 3206 543748
rect 110506 543736 110512 543748
rect 110564 543736 110570 543788
rect 3510 540948 3516 541000
rect 3568 540988 3574 541000
rect 94682 540988 94688 541000
rect 3568 540960 94688 540988
rect 3568 540948 3574 540960
rect 94682 540948 94688 540960
rect 94740 540948 94746 541000
rect 565078 540948 565084 541000
rect 565136 540988 565142 541000
rect 580166 540988 580172 541000
rect 565136 540960 580172 540988
rect 565136 540948 565142 540960
rect 580166 540948 580172 540960
rect 580224 540948 580230 541000
rect 3326 536800 3332 536852
rect 3384 536840 3390 536852
rect 97350 536840 97356 536852
rect 3384 536812 97356 536840
rect 3384 536800 3390 536812
rect 97350 536800 97356 536812
rect 97408 536800 97414 536852
rect 120166 536800 120172 536852
rect 120224 536840 120230 536852
rect 580166 536840 580172 536852
rect 120224 536812 580172 536840
rect 120224 536800 120230 536812
rect 580166 536800 580172 536812
rect 580224 536800 580230 536852
rect 3326 532720 3332 532772
rect 3384 532760 3390 532772
rect 167086 532760 167092 532772
rect 3384 532732 167092 532760
rect 3384 532720 3390 532732
rect 167086 532720 167092 532732
rect 167144 532720 167150 532772
rect 577498 529048 577504 529100
rect 577556 529088 577562 529100
rect 579798 529088 579804 529100
rect 577556 529060 579804 529088
rect 577556 529048 577562 529060
rect 579798 529048 579804 529060
rect 579856 529048 579862 529100
rect 3510 528572 3516 528624
rect 3568 528612 3574 528624
rect 95878 528612 95884 528624
rect 3568 528584 95884 528612
rect 3568 528572 3574 528584
rect 95878 528572 95884 528584
rect 95936 528572 95942 528624
rect 3510 524424 3516 524476
rect 3568 524464 3574 524476
rect 86310 524464 86316 524476
rect 3568 524436 86316 524464
rect 3568 524424 3574 524436
rect 86310 524424 86316 524436
rect 86368 524424 86374 524476
rect 555418 524424 555424 524476
rect 555476 524464 555482 524476
rect 580166 524464 580172 524476
rect 555476 524436 580172 524464
rect 555476 524424 555482 524436
rect 580166 524424 580172 524436
rect 580224 524424 580230 524476
rect 2866 520276 2872 520328
rect 2924 520316 2930 520328
rect 115198 520316 115204 520328
rect 2924 520288 115204 520316
rect 2924 520276 2930 520288
rect 115198 520276 115204 520288
rect 115256 520276 115262 520328
rect 189810 520276 189816 520328
rect 189868 520316 189874 520328
rect 580166 520316 580172 520328
rect 189868 520288 580172 520316
rect 189868 520276 189874 520288
rect 580166 520276 580172 520288
rect 580224 520276 580230 520328
rect 2958 516128 2964 516180
rect 3016 516168 3022 516180
rect 97442 516168 97448 516180
rect 3016 516140 97448 516168
rect 3016 516128 3022 516140
rect 97442 516128 97448 516140
rect 97500 516128 97506 516180
rect 3050 511980 3056 512032
rect 3108 512020 3114 512032
rect 108390 512020 108396 512032
rect 3108 511992 108396 512020
rect 3108 511980 3114 511992
rect 108390 511980 108396 511992
rect 108448 511980 108454 512032
rect 574830 509260 574836 509312
rect 574888 509300 574894 509312
rect 580166 509300 580172 509312
rect 574888 509272 580172 509300
rect 574888 509260 574894 509272
rect 580166 509260 580172 509272
rect 580224 509260 580230 509312
rect 3510 507832 3516 507884
rect 3568 507872 3574 507884
rect 95970 507872 95976 507884
rect 3568 507844 95976 507872
rect 3568 507832 3574 507844
rect 95970 507832 95976 507844
rect 96028 507832 96034 507884
rect 138658 507832 138664 507884
rect 138716 507872 138722 507884
rect 144178 507872 144184 507884
rect 138716 507844 144184 507872
rect 138716 507832 138722 507844
rect 144178 507832 144184 507844
rect 144236 507832 144242 507884
rect 554038 505112 554044 505164
rect 554096 505152 554102 505164
rect 580074 505152 580080 505164
rect 554096 505124 580080 505152
rect 554096 505112 554102 505124
rect 580074 505112 580080 505124
rect 580132 505112 580138 505164
rect 3050 503684 3056 503736
rect 3108 503724 3114 503736
rect 127158 503724 127164 503736
rect 3108 503696 127164 503724
rect 3108 503684 3114 503696
rect 127158 503684 127164 503696
rect 127216 503684 127222 503736
rect 576302 500964 576308 501016
rect 576360 501004 576366 501016
rect 580074 501004 580080 501016
rect 576360 500976 580080 501004
rect 576360 500964 576366 500976
rect 580074 500964 580080 500976
rect 580132 500964 580138 501016
rect 3326 496816 3332 496868
rect 3384 496856 3390 496868
rect 108482 496856 108488 496868
rect 3384 496828 108488 496856
rect 3384 496816 3390 496828
rect 108482 496816 108488 496828
rect 108540 496816 108546 496868
rect 554130 496816 554136 496868
rect 554188 496856 554194 496868
rect 579890 496856 579896 496868
rect 554188 496828 579896 496856
rect 554188 496816 554194 496828
rect 579890 496816 579896 496828
rect 579948 496816 579954 496868
rect 3510 492668 3516 492720
rect 3568 492708 3574 492720
rect 90542 492708 90548 492720
rect 3568 492680 90548 492708
rect 3568 492668 3574 492680
rect 90542 492668 90548 492680
rect 90600 492668 90606 492720
rect 574922 492668 574928 492720
rect 574980 492708 574986 492720
rect 580166 492708 580172 492720
rect 574980 492680 580172 492708
rect 574980 492668 574986 492680
rect 580166 492668 580172 492680
rect 580224 492668 580230 492720
rect 3326 488520 3332 488572
rect 3384 488560 3390 488572
rect 111058 488560 111064 488572
rect 3384 488532 111064 488560
rect 3384 488520 3390 488532
rect 111058 488520 111064 488532
rect 111116 488520 111122 488572
rect 566642 488520 566648 488572
rect 566700 488560 566706 488572
rect 580166 488560 580172 488572
rect 566700 488532 580172 488560
rect 566700 488520 566706 488532
rect 580166 488520 580172 488532
rect 580224 488520 580230 488572
rect 3510 484372 3516 484424
rect 3568 484412 3574 484424
rect 104434 484412 104440 484424
rect 3568 484384 104440 484412
rect 3568 484372 3574 484384
rect 104434 484372 104440 484384
rect 104492 484372 104498 484424
rect 215938 484372 215944 484424
rect 215996 484412 216002 484424
rect 580166 484412 580172 484424
rect 215996 484384 580172 484412
rect 215996 484372 216002 484384
rect 580166 484372 580172 484384
rect 580224 484372 580230 484424
rect 3510 480224 3516 480276
rect 3568 480264 3574 480276
rect 101398 480264 101404 480276
rect 3568 480236 101404 480264
rect 3568 480224 3574 480236
rect 101398 480224 101404 480236
rect 101456 480224 101462 480276
rect 561030 480224 561036 480276
rect 561088 480264 561094 480276
rect 580166 480264 580172 480276
rect 561088 480236 580172 480264
rect 561088 480224 561094 480236
rect 580166 480224 580172 480236
rect 580224 480224 580230 480276
rect 2866 476076 2872 476128
rect 2924 476116 2930 476128
rect 102962 476116 102968 476128
rect 2924 476088 102968 476116
rect 2924 476076 2930 476088
rect 102962 476076 102968 476088
rect 103020 476076 103026 476128
rect 567838 476076 567844 476128
rect 567896 476116 567902 476128
rect 580166 476116 580172 476128
rect 567896 476088 580172 476116
rect 567896 476076 567902 476088
rect 580166 476076 580172 476088
rect 580224 476076 580230 476128
rect 561122 473356 561128 473408
rect 561180 473396 561186 473408
rect 580166 473396 580172 473408
rect 561180 473368 580172 473396
rect 561180 473356 561186 473368
rect 580166 473356 580172 473368
rect 580224 473356 580230 473408
rect 2866 471996 2872 472048
rect 2924 472036 2930 472048
rect 87598 472036 87604 472048
rect 2924 472008 87604 472036
rect 2924 471996 2930 472008
rect 87598 471996 87604 472008
rect 87656 471996 87662 472048
rect 128354 469820 128360 469872
rect 128412 469860 128418 469872
rect 147674 469860 147680 469872
rect 128412 469832 147680 469860
rect 128412 469820 128418 469832
rect 147674 469820 147680 469832
rect 147732 469820 147738 469872
rect 2958 467848 2964 467900
rect 3016 467888 3022 467900
rect 100202 467888 100208 467900
rect 3016 467860 100208 467888
rect 3016 467848 3022 467860
rect 100202 467848 100208 467860
rect 100260 467848 100266 467900
rect 3510 465060 3516 465112
rect 3568 465100 3574 465112
rect 93210 465100 93216 465112
rect 3568 465072 93216 465100
rect 3568 465060 3574 465072
rect 93210 465060 93216 465072
rect 93268 465060 93274 465112
rect 573358 465060 573364 465112
rect 573416 465100 573422 465112
rect 580166 465100 580172 465112
rect 573416 465072 580172 465100
rect 573416 465060 573422 465072
rect 580166 465060 580172 465072
rect 580224 465060 580230 465112
rect 3510 460912 3516 460964
rect 3568 460952 3574 460964
rect 113818 460952 113824 460964
rect 3568 460924 113824 460952
rect 3568 460912 3574 460924
rect 113818 460912 113824 460924
rect 113876 460912 113882 460964
rect 556890 460912 556896 460964
rect 556948 460952 556954 460964
rect 580074 460952 580080 460964
rect 556948 460924 580080 460952
rect 556948 460912 556954 460924
rect 580074 460912 580080 460924
rect 580132 460912 580138 460964
rect 3234 456764 3240 456816
rect 3292 456804 3298 456816
rect 105538 456804 105544 456816
rect 3292 456776 105544 456804
rect 3292 456764 3298 456776
rect 105538 456764 105544 456776
rect 105596 456764 105602 456816
rect 119982 456764 119988 456816
rect 120040 456804 120046 456816
rect 580074 456804 580080 456816
rect 120040 456776 580080 456804
rect 120040 456764 120046 456776
rect 580074 456764 580080 456776
rect 580132 456764 580138 456816
rect 3326 452616 3332 452668
rect 3384 452656 3390 452668
rect 126238 452656 126244 452668
rect 3384 452628 126244 452656
rect 3384 452616 3390 452628
rect 126238 452616 126244 452628
rect 126296 452616 126302 452668
rect 3326 448536 3332 448588
rect 3384 448576 3390 448588
rect 120810 448576 120816 448588
rect 3384 448548 120816 448576
rect 3384 448536 3390 448548
rect 120810 448536 120816 448548
rect 120868 448536 120874 448588
rect 563698 448536 563704 448588
rect 563756 448576 563762 448588
rect 579706 448576 579712 448588
rect 563756 448548 579712 448576
rect 563756 448536 563762 448548
rect 579706 448536 579712 448548
rect 579764 448536 579770 448588
rect 3510 444388 3516 444440
rect 3568 444428 3574 444440
rect 109126 444428 109132 444440
rect 3568 444400 109132 444428
rect 3568 444388 3574 444400
rect 109126 444388 109132 444400
rect 109184 444388 109190 444440
rect 570690 444388 570696 444440
rect 570748 444428 570754 444440
rect 580166 444428 580172 444440
rect 570748 444400 580172 444428
rect 570748 444388 570754 444400
rect 580166 444388 580172 444400
rect 580224 444388 580230 444440
rect 3326 440240 3332 440292
rect 3384 440280 3390 440292
rect 119338 440280 119344 440292
rect 3384 440252 119344 440280
rect 3384 440240 3390 440252
rect 119338 440240 119344 440252
rect 119396 440240 119402 440292
rect 572070 440240 572076 440292
rect 572128 440280 572134 440292
rect 580166 440280 580172 440292
rect 572128 440252 580172 440280
rect 572128 440240 572134 440252
rect 580166 440240 580172 440252
rect 580224 440240 580230 440292
rect 3510 436092 3516 436144
rect 3568 436132 3574 436144
rect 183646 436132 183652 436144
rect 3568 436104 183652 436132
rect 3568 436092 3574 436104
rect 183646 436092 183652 436104
rect 183704 436092 183710 436144
rect 567930 436092 567936 436144
rect 567988 436132 567994 436144
rect 579614 436132 579620 436144
rect 567988 436104 579620 436132
rect 567988 436092 567994 436104
rect 579614 436092 579620 436104
rect 579672 436092 579678 436144
rect 3510 431944 3516 431996
rect 3568 431984 3574 431996
rect 93394 431984 93400 431996
rect 3568 431956 93400 431984
rect 3568 431944 3574 431956
rect 93394 431944 93400 431956
rect 93452 431944 93458 431996
rect 563790 431944 563796 431996
rect 563848 431984 563854 431996
rect 580166 431984 580172 431996
rect 563848 431956 580172 431984
rect 563848 431944 563854 431956
rect 580166 431944 580172 431956
rect 580224 431944 580230 431996
rect 563882 429156 563888 429208
rect 563940 429196 563946 429208
rect 579982 429196 579988 429208
rect 563940 429168 579988 429196
rect 563940 429156 563946 429168
rect 579982 429156 579988 429168
rect 580040 429156 580046 429208
rect 2866 427796 2872 427848
rect 2924 427836 2930 427848
rect 108574 427836 108580 427848
rect 2924 427808 108580 427836
rect 2924 427796 2930 427808
rect 108574 427796 108580 427808
rect 108632 427796 108638 427848
rect 577590 425076 577596 425128
rect 577648 425116 577654 425128
rect 579614 425116 579620 425128
rect 577648 425088 579620 425116
rect 577648 425076 577654 425088
rect 579614 425076 579620 425088
rect 579672 425076 579678 425128
rect 3510 416780 3516 416832
rect 3568 416820 3574 416832
rect 112530 416820 112536 416832
rect 3568 416792 112536 416820
rect 3568 416780 3574 416792
rect 112530 416780 112536 416792
rect 112588 416780 112594 416832
rect 3510 412632 3516 412684
rect 3568 412672 3574 412684
rect 118050 412672 118056 412684
rect 3568 412644 118056 412672
rect 3568 412632 3574 412644
rect 118050 412632 118056 412644
rect 118108 412632 118114 412684
rect 572162 412632 572168 412684
rect 572220 412672 572226 412684
rect 580166 412672 580172 412684
rect 572220 412644 580172 412672
rect 572220 412632 572226 412644
rect 580166 412632 580172 412644
rect 580224 412632 580230 412684
rect 3510 408484 3516 408536
rect 3568 408524 3574 408536
rect 104986 408524 104992 408536
rect 3568 408496 104992 408524
rect 3568 408484 3574 408496
rect 104986 408484 104992 408496
rect 105044 408484 105050 408536
rect 149698 407736 149704 407788
rect 149756 407776 149762 407788
rect 182266 407776 182272 407788
rect 149756 407748 182272 407776
rect 149756 407736 149762 407748
rect 182266 407736 182272 407748
rect 182324 407736 182330 407788
rect 552842 404336 552848 404388
rect 552900 404376 552906 404388
rect 580166 404376 580172 404388
rect 552900 404348 580172 404376
rect 552900 404336 552906 404348
rect 580166 404336 580172 404348
rect 580224 404336 580230 404388
rect 3234 400188 3240 400240
rect 3292 400228 3298 400240
rect 184934 400228 184940 400240
rect 3292 400200 184940 400228
rect 3292 400188 3298 400200
rect 184934 400188 184940 400200
rect 184992 400188 184998 400240
rect 191742 400188 191748 400240
rect 191800 400228 191806 400240
rect 580166 400228 580172 400240
rect 191800 400200 580172 400228
rect 191800 400188 191806 400200
rect 580166 400188 580172 400200
rect 580224 400188 580230 400240
rect 3602 396040 3608 396092
rect 3660 396080 3666 396092
rect 79410 396080 79416 396092
rect 3660 396052 79416 396080
rect 3660 396040 3666 396052
rect 79410 396040 79416 396052
rect 79468 396040 79474 396092
rect 569218 391960 569224 392012
rect 569276 392000 569282 392012
rect 580166 392000 580172 392012
rect 569276 391972 580172 392000
rect 569276 391960 569282 391972
rect 580166 391960 580172 391972
rect 580224 391960 580230 392012
rect 2958 387812 2964 387864
rect 3016 387852 3022 387864
rect 87690 387852 87696 387864
rect 3016 387824 87696 387852
rect 3016 387812 3022 387824
rect 87690 387812 87696 387824
rect 87748 387812 87754 387864
rect 121270 385024 121276 385076
rect 121328 385064 121334 385076
rect 579798 385064 579804 385076
rect 121328 385036 579804 385064
rect 121328 385024 121334 385036
rect 579798 385024 579804 385036
rect 579856 385024 579862 385076
rect 3142 383664 3148 383716
rect 3200 383704 3206 383716
rect 94774 383704 94780 383716
rect 3200 383676 94780 383704
rect 3200 383664 3206 383676
rect 94774 383664 94780 383676
rect 94832 383664 94838 383716
rect 196618 380876 196624 380928
rect 196676 380916 196682 380928
rect 579982 380916 579988 380928
rect 196676 380888 579988 380916
rect 196676 380876 196682 380888
rect 579982 380876 579988 380888
rect 580040 380876 580046 380928
rect 3326 379516 3332 379568
rect 3384 379556 3390 379568
rect 107010 379556 107016 379568
rect 3384 379528 107016 379556
rect 3384 379516 3390 379528
rect 107010 379516 107016 379528
rect 107068 379516 107074 379568
rect 3326 376728 3332 376780
rect 3384 376768 3390 376780
rect 90634 376768 90640 376780
rect 3384 376740 90640 376768
rect 3384 376728 3390 376740
rect 90634 376728 90640 376740
rect 90692 376728 90698 376780
rect 569310 376728 569316 376780
rect 569368 376768 569374 376780
rect 580166 376768 580172 376780
rect 569368 376740 580172 376768
rect 569368 376728 569374 376740
rect 580166 376728 580172 376740
rect 580224 376728 580230 376780
rect 3326 372580 3332 372632
rect 3384 372620 3390 372632
rect 194594 372620 194600 372632
rect 3384 372592 194600 372620
rect 3384 372580 3390 372592
rect 194594 372580 194600 372592
rect 194652 372580 194658 372632
rect 556982 372580 556988 372632
rect 557040 372620 557046 372632
rect 580166 372620 580172 372632
rect 557040 372592 580172 372620
rect 557040 372580 557046 372592
rect 580166 372580 580172 372592
rect 580224 372580 580230 372632
rect 3326 368500 3332 368552
rect 3384 368540 3390 368552
rect 97534 368540 97540 368552
rect 3384 368512 97540 368540
rect 3384 368500 3390 368512
rect 97534 368500 97540 368512
rect 97592 368500 97598 368552
rect 559650 368500 559656 368552
rect 559708 368540 559714 368552
rect 580166 368540 580172 368552
rect 559708 368512 580172 368540
rect 559708 368500 559714 368512
rect 580166 368500 580172 368512
rect 580224 368500 580230 368552
rect 3326 364488 3332 364540
rect 3384 364528 3390 364540
rect 7558 364528 7564 364540
rect 3384 364500 7564 364528
rect 3384 364488 3390 364500
rect 7558 364488 7564 364500
rect 7616 364488 7622 364540
rect 191098 364352 191104 364404
rect 191156 364392 191162 364404
rect 579614 364392 579620 364404
rect 191156 364364 579620 364392
rect 191156 364352 191162 364364
rect 579614 364352 579620 364364
rect 579672 364352 579678 364404
rect 3326 360204 3332 360256
rect 3384 360244 3390 360256
rect 103054 360244 103060 360256
rect 3384 360216 103060 360244
rect 3384 360204 3390 360216
rect 103054 360204 103060 360216
rect 103112 360204 103118 360256
rect 561214 360204 561220 360256
rect 561272 360244 561278 360256
rect 579614 360244 579620 360256
rect 561272 360216 579620 360244
rect 561272 360204 561278 360216
rect 579614 360204 579620 360216
rect 579672 360204 579678 360256
rect 3326 356056 3332 356108
rect 3384 356096 3390 356108
rect 98914 356096 98920 356108
rect 3384 356068 98920 356096
rect 3384 356056 3390 356068
rect 98914 356056 98920 356068
rect 98972 356056 98978 356108
rect 192570 356056 192576 356108
rect 192628 356096 192634 356108
rect 580166 356096 580172 356108
rect 192628 356068 580172 356096
rect 192628 356056 192634 356068
rect 580166 356056 580172 356068
rect 580224 356056 580230 356108
rect 563974 353268 563980 353320
rect 564032 353308 564038 353320
rect 579614 353308 579620 353320
rect 564032 353280 579620 353308
rect 564032 353268 564038 353280
rect 579614 353268 579620 353280
rect 579672 353268 579678 353320
rect 3234 351908 3240 351960
rect 3292 351948 3298 351960
rect 96062 351948 96068 351960
rect 3292 351920 96068 351948
rect 3292 351908 3298 351920
rect 96062 351908 96068 351920
rect 96120 351908 96126 351960
rect 194502 349120 194508 349172
rect 194560 349160 194566 349172
rect 580166 349160 580172 349172
rect 194560 349132 580172 349160
rect 194560 349120 194566 349132
rect 580166 349120 580172 349132
rect 580224 349120 580230 349172
rect 3142 347760 3148 347812
rect 3200 347800 3206 347812
rect 120902 347800 120908 347812
rect 3200 347772 120908 347800
rect 3200 347760 3206 347772
rect 120902 347760 120908 347772
rect 120960 347760 120966 347812
rect 558454 345040 558460 345092
rect 558512 345080 558518 345092
rect 580166 345080 580172 345092
rect 558512 345052 580172 345080
rect 558512 345040 558518 345052
rect 580166 345040 580172 345052
rect 580224 345040 580230 345092
rect 3326 343612 3332 343664
rect 3384 343652 3390 343664
rect 107102 343652 107108 343664
rect 3384 343624 107108 343652
rect 3384 343612 3390 343624
rect 107102 343612 107108 343624
rect 107160 343612 107166 343664
rect 575014 340892 575020 340944
rect 575072 340932 575078 340944
rect 580166 340932 580172 340944
rect 575072 340904 580172 340932
rect 575072 340892 575078 340904
rect 580166 340892 580172 340904
rect 580224 340892 580230 340944
rect 3142 339464 3148 339516
rect 3200 339504 3206 339516
rect 113910 339504 113916 339516
rect 3200 339476 113916 339504
rect 3200 339464 3206 339476
rect 113910 339464 113916 339476
rect 113968 339464 113974 339516
rect 128446 336744 128452 336796
rect 128504 336784 128510 336796
rect 579982 336784 579988 336796
rect 128504 336756 579988 336784
rect 128504 336744 128510 336756
rect 579982 336744 579988 336756
rect 580040 336744 580046 336796
rect 171042 335996 171048 336048
rect 171100 336036 171106 336048
rect 359458 336036 359464 336048
rect 171100 336008 359464 336036
rect 171100 335996 171106 336008
rect 359458 335996 359464 336008
rect 359516 335996 359522 336048
rect 3326 335316 3332 335368
rect 3384 335356 3390 335368
rect 103146 335356 103152 335368
rect 3384 335328 103152 335356
rect 3384 335316 3390 335328
rect 103146 335316 103152 335328
rect 103204 335316 103210 335368
rect 3326 332596 3332 332648
rect 3384 332636 3390 332648
rect 101490 332636 101496 332648
rect 3384 332608 101496 332636
rect 3384 332596 3390 332608
rect 101490 332596 101496 332608
rect 101548 332596 101554 332648
rect 572254 332596 572260 332648
rect 572312 332636 572318 332648
rect 579982 332636 579988 332648
rect 572312 332608 579988 332636
rect 572312 332596 572318 332608
rect 579982 332596 579988 332608
rect 580040 332596 580046 332648
rect 3326 328448 3332 328500
rect 3384 328488 3390 328500
rect 99006 328488 99012 328500
rect 3384 328460 99012 328488
rect 3384 328448 3390 328460
rect 99006 328448 99012 328460
rect 99064 328448 99070 328500
rect 3326 324300 3332 324352
rect 3384 324340 3390 324352
rect 96154 324340 96160 324352
rect 3384 324312 96160 324340
rect 3384 324300 3390 324312
rect 96154 324300 96160 324312
rect 96212 324300 96218 324352
rect 3142 320152 3148 320204
rect 3200 320192 3206 320204
rect 125686 320192 125692 320204
rect 3200 320164 125692 320192
rect 3200 320152 3206 320164
rect 125686 320152 125692 320164
rect 125744 320152 125750 320204
rect 575106 320152 575112 320204
rect 575164 320192 575170 320204
rect 579614 320192 579620 320204
rect 575164 320164 579620 320192
rect 575164 320152 575170 320164
rect 579614 320152 579620 320164
rect 579672 320152 579678 320204
rect 3326 316004 3332 316056
rect 3384 316044 3390 316056
rect 119430 316044 119436 316056
rect 3384 316016 119436 316044
rect 3384 316004 3390 316016
rect 119430 316004 119436 316016
rect 119488 316004 119494 316056
rect 566734 316004 566740 316056
rect 566792 316044 566798 316056
rect 579614 316044 579620 316056
rect 566792 316016 579620 316044
rect 566792 316004 566798 316016
rect 579614 316004 579620 316016
rect 579672 316004 579678 316056
rect 577682 313284 577688 313336
rect 577740 313324 577746 313336
rect 580626 313324 580632 313336
rect 577740 313296 580632 313324
rect 577740 313284 577746 313296
rect 580626 313284 580632 313296
rect 580684 313284 580690 313336
rect 555510 309136 555516 309188
rect 555568 309176 555574 309188
rect 580166 309176 580172 309188
rect 555568 309148 580172 309176
rect 555568 309136 555574 309148
rect 580166 309136 580172 309148
rect 580224 309136 580230 309188
rect 3326 307776 3332 307828
rect 3384 307816 3390 307828
rect 107194 307816 107200 307828
rect 3384 307788 107200 307816
rect 3384 307776 3390 307788
rect 107194 307776 107200 307788
rect 107252 307776 107258 307828
rect 572346 304988 572352 305040
rect 572404 305028 572410 305040
rect 579614 305028 579620 305040
rect 572404 305000 579620 305028
rect 572404 304988 572410 305000
rect 579614 304988 579620 305000
rect 579672 304988 579678 305040
rect 3050 303628 3056 303680
rect 3108 303668 3114 303680
rect 104618 303668 104624 303680
rect 3108 303640 104624 303668
rect 3108 303628 3114 303640
rect 104618 303628 104624 303640
rect 104676 303628 104682 303680
rect 577774 300840 577780 300892
rect 577832 300880 577838 300892
rect 580626 300880 580632 300892
rect 577832 300852 580632 300880
rect 577832 300840 577838 300852
rect 580626 300840 580632 300852
rect 580684 300840 580690 300892
rect 3142 299480 3148 299532
rect 3200 299520 3206 299532
rect 104066 299520 104072 299532
rect 3200 299492 104072 299520
rect 3200 299480 3206 299492
rect 104066 299480 104072 299492
rect 104124 299480 104130 299532
rect 180058 296692 180064 296744
rect 180116 296732 180122 296744
rect 580166 296732 580172 296744
rect 180116 296704 580172 296732
rect 180116 296692 180122 296704
rect 580166 296692 580172 296704
rect 580224 296692 580230 296744
rect 3326 295332 3332 295384
rect 3384 295372 3390 295384
rect 10318 295372 10324 295384
rect 3384 295344 10324 295372
rect 3384 295332 3390 295344
rect 10318 295332 10324 295344
rect 10376 295332 10382 295384
rect 569402 292544 569408 292596
rect 569460 292584 569466 292596
rect 579982 292584 579988 292596
rect 569460 292556 579988 292584
rect 569460 292544 569466 292556
rect 579982 292544 579988 292556
rect 580040 292544 580046 292596
rect 3142 291184 3148 291236
rect 3200 291224 3206 291236
rect 122098 291224 122104 291236
rect 3200 291196 122104 291224
rect 3200 291184 3206 291196
rect 122098 291184 122104 291196
rect 122156 291184 122162 291236
rect 561306 288396 561312 288448
rect 561364 288436 561370 288448
rect 579982 288436 579988 288448
rect 561364 288408 579988 288436
rect 561364 288396 561370 288408
rect 579982 288396 579988 288408
rect 580040 288396 580046 288448
rect 3326 287036 3332 287088
rect 3384 287076 3390 287088
rect 108666 287076 108672 287088
rect 3384 287048 108672 287076
rect 3384 287036 3390 287048
rect 108666 287036 108672 287048
rect 108724 287036 108730 287088
rect 3326 284316 3332 284368
rect 3384 284356 3390 284368
rect 101582 284356 101588 284368
rect 3384 284328 101588 284356
rect 3384 284316 3390 284328
rect 101582 284316 101588 284328
rect 101640 284316 101646 284368
rect 3326 280168 3332 280220
rect 3384 280208 3390 280220
rect 99098 280208 99104 280220
rect 3384 280180 99104 280208
rect 3384 280168 3390 280180
rect 99098 280168 99104 280180
rect 99156 280168 99162 280220
rect 558546 280168 558552 280220
rect 558604 280208 558610 280220
rect 580166 280208 580172 280220
rect 558604 280180 580172 280208
rect 558604 280168 558610 280180
rect 580166 280168 580172 280180
rect 580224 280168 580230 280220
rect 13078 277992 13084 278044
rect 13136 278032 13142 278044
rect 174538 278032 174544 278044
rect 13136 278004 174544 278032
rect 13136 277992 13142 278004
rect 174538 277992 174544 278004
rect 174596 277992 174602 278044
rect 564066 276020 564072 276072
rect 564124 276060 564130 276072
rect 580166 276060 580172 276072
rect 564124 276032 580172 276060
rect 564124 276020 564130 276032
rect 580166 276020 580172 276032
rect 580224 276020 580230 276072
rect 124858 275272 124864 275324
rect 124916 275312 124922 275324
rect 396074 275312 396080 275324
rect 124916 275284 396080 275312
rect 124916 275272 124922 275284
rect 396074 275272 396080 275284
rect 396132 275272 396138 275324
rect 14458 273912 14464 273964
rect 14516 273952 14522 273964
rect 109218 273952 109224 273964
rect 14516 273924 109224 273952
rect 14516 273912 14522 273924
rect 109218 273912 109224 273924
rect 109276 273912 109282 273964
rect 109218 273232 109224 273284
rect 109276 273272 109282 273284
rect 110230 273272 110236 273284
rect 109276 273244 110236 273272
rect 109276 273232 109282 273244
rect 110230 273232 110236 273244
rect 110288 273272 110294 273284
rect 133874 273272 133880 273284
rect 110288 273244 133880 273272
rect 110288 273232 110294 273244
rect 133874 273232 133880 273244
rect 133932 273232 133938 273284
rect 575198 273232 575204 273284
rect 575256 273272 575262 273284
rect 580166 273272 580172 273284
rect 575256 273244 580172 273272
rect 575256 273232 575262 273244
rect 580166 273232 580172 273244
rect 580224 273232 580230 273284
rect 3142 271872 3148 271924
rect 3200 271912 3206 271924
rect 145558 271912 145564 271924
rect 3200 271884 145564 271912
rect 3200 271872 3206 271884
rect 145558 271872 145564 271884
rect 145616 271872 145622 271924
rect 7558 271124 7564 271176
rect 7616 271164 7622 271176
rect 165614 271164 165620 271176
rect 7616 271136 165620 271164
rect 7616 271124 7622 271136
rect 165614 271124 165620 271136
rect 165672 271124 165678 271176
rect 148962 269832 148968 269884
rect 149020 269872 149026 269884
rect 288434 269872 288440 269884
rect 149020 269844 288440 269872
rect 149020 269832 149026 269844
rect 288434 269832 288440 269844
rect 288492 269832 288498 269884
rect 10318 269764 10324 269816
rect 10376 269804 10382 269816
rect 161474 269804 161480 269816
rect 10376 269776 161480 269804
rect 10376 269764 10382 269776
rect 161474 269764 161480 269776
rect 161532 269764 161538 269816
rect 79410 268336 79416 268388
rect 79468 268376 79474 268388
rect 156046 268376 156052 268388
rect 79468 268348 156052 268376
rect 79468 268336 79474 268348
rect 156046 268336 156052 268348
rect 156104 268336 156110 268388
rect 153102 267044 153108 267096
rect 153160 267084 153166 267096
rect 199378 267084 199384 267096
rect 153160 267056 199384 267084
rect 153160 267044 153166 267056
rect 199378 267044 199384 267056
rect 199436 267044 199442 267096
rect 21358 266976 21364 267028
rect 21416 267016 21422 267028
rect 115382 267016 115388 267028
rect 21416 266988 115388 267016
rect 21416 266976 21422 266988
rect 115382 266976 115388 266988
rect 115440 266976 115446 267028
rect 191650 266976 191656 267028
rect 191708 267016 191714 267028
rect 440234 267016 440240 267028
rect 191708 266988 440240 267016
rect 191708 266976 191714 266988
rect 440234 266976 440240 266988
rect 440292 266976 440298 267028
rect 155678 266364 155684 266416
rect 155736 266404 155742 266416
rect 190546 266404 190552 266416
rect 155736 266376 190552 266404
rect 155736 266364 155742 266376
rect 190546 266364 190552 266376
rect 190604 266404 190610 266416
rect 191650 266404 191656 266416
rect 190604 266376 191656 266404
rect 190604 266364 190610 266376
rect 191650 266364 191656 266376
rect 191708 266364 191714 266416
rect 145558 265820 145564 265872
rect 145616 265860 145622 265872
rect 169754 265860 169760 265872
rect 145616 265832 169760 265860
rect 145616 265820 145622 265832
rect 169754 265820 169760 265832
rect 169812 265820 169818 265872
rect 155954 265752 155960 265804
rect 156012 265792 156018 265804
rect 190454 265792 190460 265804
rect 156012 265764 190460 265792
rect 156012 265752 156018 265764
rect 190454 265752 190460 265764
rect 190512 265752 190518 265804
rect 151814 265684 151820 265736
rect 151872 265724 151878 265736
rect 196066 265724 196072 265736
rect 151872 265696 196072 265724
rect 151872 265684 151878 265696
rect 196066 265684 196072 265696
rect 196124 265684 196130 265736
rect 67634 265616 67640 265668
rect 67692 265656 67698 265668
rect 173066 265656 173072 265668
rect 67692 265628 173072 265656
rect 67692 265616 67698 265628
rect 173066 265616 173072 265628
rect 173124 265616 173130 265668
rect 179322 265140 179328 265192
rect 179380 265180 179386 265192
rect 197538 265180 197544 265192
rect 179380 265152 197544 265180
rect 179380 265140 179386 265152
rect 197538 265140 197544 265152
rect 197596 265140 197602 265192
rect 174538 265072 174544 265124
rect 174596 265112 174602 265124
rect 193490 265112 193496 265124
rect 174596 265084 193496 265112
rect 174596 265072 174602 265084
rect 193490 265072 193496 265084
rect 193548 265072 193554 265124
rect 162762 265004 162768 265056
rect 162820 265044 162826 265056
rect 193306 265044 193312 265056
rect 162820 265016 193312 265044
rect 162820 265004 162826 265016
rect 193306 265004 193312 265016
rect 193364 265044 193370 265056
rect 196618 265044 196624 265056
rect 193364 265016 196624 265044
rect 193364 265004 193370 265016
rect 196618 265004 196624 265016
rect 196676 265004 196682 265056
rect 112530 264936 112536 264988
rect 112588 264976 112594 264988
rect 115750 264976 115756 264988
rect 112588 264948 115756 264976
rect 112588 264936 112594 264948
rect 115750 264936 115756 264948
rect 115808 264976 115814 264988
rect 146754 264976 146760 264988
rect 115808 264948 146760 264976
rect 115808 264936 115814 264948
rect 146754 264936 146760 264948
rect 146812 264936 146818 264988
rect 161474 264936 161480 264988
rect 161532 264976 161538 264988
rect 194778 264976 194784 264988
rect 161532 264948 194784 264976
rect 161532 264936 161538 264948
rect 194778 264936 194784 264948
rect 194836 264936 194842 264988
rect 566826 264936 566832 264988
rect 566884 264976 566890 264988
rect 580166 264976 580172 264988
rect 566884 264948 580172 264976
rect 566884 264936 566890 264948
rect 580166 264936 580172 264948
rect 580224 264936 580230 264988
rect 146202 264256 146208 264308
rect 146260 264296 146266 264308
rect 180058 264296 180064 264308
rect 146260 264268 180064 264296
rect 146260 264256 146266 264268
rect 180058 264256 180064 264268
rect 180116 264256 180122 264308
rect 34514 264188 34520 264240
rect 34572 264228 34578 264240
rect 118694 264228 118700 264240
rect 34572 264200 118700 264228
rect 34572 264188 34578 264200
rect 118694 264188 118700 264200
rect 118752 264188 118758 264240
rect 192570 264228 192576 264240
rect 151786 264200 192576 264228
rect 115014 264052 115020 264104
rect 115072 264092 115078 264104
rect 148962 264092 148968 264104
rect 115072 264064 148968 264092
rect 115072 264052 115078 264064
rect 148962 264052 148968 264064
rect 149020 264052 149026 264104
rect 115566 263984 115572 264036
rect 115624 264024 115630 264036
rect 135438 264024 135444 264036
rect 115624 263996 135444 264024
rect 115624 263984 115630 263996
rect 135438 263984 135444 263996
rect 135496 263984 135502 264036
rect 112714 263916 112720 263968
rect 112772 263956 112778 263968
rect 138658 263956 138664 263968
rect 112772 263928 138664 263956
rect 112772 263916 112778 263928
rect 138658 263916 138664 263928
rect 138716 263916 138722 263968
rect 117682 263848 117688 263900
rect 117740 263888 117746 263900
rect 145374 263888 145380 263900
rect 117740 263860 145380 263888
rect 117740 263848 117746 263860
rect 145374 263848 145380 263860
rect 145432 263888 145438 263900
rect 151786 263888 151814 264200
rect 192570 264188 192576 264200
rect 192628 264188 192634 264240
rect 195054 264188 195060 264240
rect 195112 264228 195118 264240
rect 215938 264228 215944 264240
rect 195112 264200 215944 264228
rect 195112 264188 195118 264200
rect 215938 264188 215944 264200
rect 215996 264188 216002 264240
rect 145432 263860 151814 263888
rect 145432 263848 145438 263860
rect 117130 263780 117136 263832
rect 117188 263820 117194 263832
rect 146202 263820 146208 263832
rect 117188 263792 146208 263820
rect 117188 263780 117194 263792
rect 146202 263780 146208 263792
rect 146260 263780 146266 263832
rect 120994 263712 121000 263764
rect 121052 263752 121058 263764
rect 151998 263752 152004 263764
rect 121052 263724 152004 263752
rect 121052 263712 121058 263724
rect 151998 263712 152004 263724
rect 152056 263752 152062 263764
rect 153102 263752 153108 263764
rect 152056 263724 153108 263752
rect 152056 263712 152062 263724
rect 153102 263712 153108 263724
rect 153160 263712 153166 263764
rect 118694 263644 118700 263696
rect 118752 263684 118758 263696
rect 119062 263684 119068 263696
rect 118752 263656 119068 263684
rect 118752 263644 118758 263656
rect 119062 263644 119068 263656
rect 119120 263684 119126 263696
rect 152550 263684 152556 263696
rect 119120 263656 152556 263684
rect 119120 263644 119126 263656
rect 152550 263644 152556 263656
rect 152608 263644 152614 263696
rect 185486 263644 185492 263696
rect 185544 263684 185550 263696
rect 194686 263684 194692 263696
rect 185544 263656 194692 263684
rect 185544 263644 185550 263656
rect 194686 263644 194692 263656
rect 194744 263684 194750 263696
rect 195054 263684 195060 263696
rect 194744 263656 195060 263684
rect 194744 263644 194750 263656
rect 195054 263644 195060 263656
rect 195112 263644 195118 263696
rect 3326 263576 3332 263628
rect 3384 263616 3390 263628
rect 107286 263616 107292 263628
rect 3384 263588 107292 263616
rect 3384 263576 3390 263588
rect 107286 263576 107292 263588
rect 107344 263576 107350 263628
rect 113910 263576 113916 263628
rect 113968 263616 113974 263628
rect 115566 263616 115572 263628
rect 113968 263588 115572 263616
rect 113968 263576 113974 263588
rect 115566 263576 115572 263588
rect 115624 263576 115630 263628
rect 159818 263576 159824 263628
rect 159876 263616 159882 263628
rect 194962 263616 194968 263628
rect 159876 263588 194968 263616
rect 159876 263576 159882 263588
rect 194962 263576 194968 263588
rect 195020 263616 195026 263628
rect 200758 263616 200764 263628
rect 195020 263588 200764 263616
rect 195020 263576 195026 263588
rect 200758 263576 200764 263588
rect 200816 263576 200822 263628
rect 113910 263168 113916 263220
rect 113968 263208 113974 263220
rect 143534 263208 143540 263220
rect 113968 263180 143540 263208
rect 113968 263168 113974 263180
rect 143534 263168 143540 263180
rect 143592 263168 143598 263220
rect 160646 263168 160652 263220
rect 160704 263208 160710 263220
rect 193398 263208 193404 263220
rect 160704 263180 193404 263208
rect 160704 263168 160710 263180
rect 193398 263168 193404 263180
rect 193456 263168 193462 263220
rect 111610 263100 111616 263152
rect 111668 263140 111674 263152
rect 141786 263140 141792 263152
rect 111668 263112 141792 263140
rect 111668 263100 111674 263112
rect 141786 263100 141792 263112
rect 141844 263100 141850 263152
rect 169662 263100 169668 263152
rect 169720 263140 169726 263152
rect 198918 263140 198924 263152
rect 169720 263112 198924 263140
rect 169720 263100 169726 263112
rect 198918 263100 198924 263112
rect 198976 263100 198982 263152
rect 112530 263032 112536 263084
rect 112588 263072 112594 263084
rect 131298 263072 131304 263084
rect 112588 263044 131304 263072
rect 112588 263032 112594 263044
rect 131298 263032 131304 263044
rect 131356 263072 131362 263084
rect 131356 263044 132494 263072
rect 131356 263032 131362 263044
rect 126238 262964 126244 263016
rect 126296 263004 126302 263016
rect 127894 263004 127900 263016
rect 126296 262976 127900 263004
rect 126296 262964 126302 262976
rect 127894 262964 127900 262976
rect 127952 262964 127958 263016
rect 132466 263004 132494 263044
rect 157242 263032 157248 263084
rect 157300 263072 157306 263084
rect 182174 263072 182180 263084
rect 157300 263044 182180 263072
rect 157300 263032 157306 263044
rect 182174 263032 182180 263044
rect 182232 263072 182238 263084
rect 183462 263072 183468 263084
rect 182232 263044 183468 263072
rect 182232 263032 182238 263044
rect 183462 263032 183468 263044
rect 183520 263032 183526 263084
rect 198734 263032 198740 263084
rect 198792 263072 198798 263084
rect 285674 263072 285680 263084
rect 198792 263044 285680 263072
rect 198792 263032 198798 263044
rect 285674 263032 285680 263044
rect 285732 263032 285738 263084
rect 327074 263004 327080 263016
rect 132466 262976 327080 263004
rect 327074 262964 327080 262976
rect 327132 262964 327138 263016
rect 122098 262896 122104 262948
rect 122156 262936 122162 262948
rect 188154 262936 188160 262948
rect 122156 262908 188160 262936
rect 122156 262896 122162 262908
rect 188154 262896 188160 262908
rect 188212 262896 188218 262948
rect 444374 262936 444380 262948
rect 198476 262908 444380 262936
rect 38654 262828 38660 262880
rect 38712 262868 38718 262880
rect 38712 262840 161474 262868
rect 38712 262828 38718 262840
rect 117038 262760 117044 262812
rect 117096 262800 117102 262812
rect 150066 262800 150072 262812
rect 117096 262772 150072 262800
rect 117096 262760 117102 262772
rect 150066 262760 150072 262772
rect 150124 262760 150130 262812
rect 161446 262800 161474 262840
rect 183462 262828 183468 262880
rect 183520 262868 183526 262880
rect 192570 262868 192576 262880
rect 183520 262840 192576 262868
rect 183520 262828 183526 262840
rect 192570 262828 192576 262840
rect 192628 262828 192634 262880
rect 164418 262800 164424 262812
rect 161446 262772 164424 262800
rect 164418 262760 164424 262772
rect 164476 262800 164482 262812
rect 197814 262800 197820 262812
rect 164476 262772 197820 262800
rect 164476 262760 164482 262772
rect 197814 262760 197820 262772
rect 197872 262760 197878 262812
rect 114278 262692 114284 262744
rect 114336 262732 114342 262744
rect 133506 262732 133512 262744
rect 114336 262704 133512 262732
rect 114336 262692 114342 262704
rect 133506 262692 133512 262704
rect 133564 262692 133570 262744
rect 183462 262692 183468 262744
rect 183520 262732 183526 262744
rect 198366 262732 198372 262744
rect 183520 262704 198372 262732
rect 183520 262692 183526 262704
rect 198366 262692 198372 262704
rect 198424 262692 198430 262744
rect 198476 262676 198504 262908
rect 444374 262896 444380 262908
rect 444432 262896 444438 262948
rect 198918 262828 198924 262880
rect 198976 262868 198982 262880
rect 199562 262868 199568 262880
rect 198976 262840 199568 262868
rect 198976 262828 198982 262840
rect 199562 262828 199568 262840
rect 199620 262868 199626 262880
rect 467834 262868 467840 262880
rect 199620 262840 467840 262868
rect 199620 262828 199626 262840
rect 467834 262828 467840 262840
rect 467892 262828 467898 262880
rect 116946 262624 116952 262676
rect 117004 262664 117010 262676
rect 140130 262664 140136 262676
rect 117004 262636 140136 262664
rect 117004 262624 117010 262636
rect 140130 262624 140136 262636
rect 140188 262624 140194 262676
rect 177206 262624 177212 262676
rect 177264 262664 177270 262676
rect 198458 262664 198464 262676
rect 177264 262636 198464 262664
rect 177264 262624 177270 262636
rect 198458 262624 198464 262636
rect 198516 262624 198522 262676
rect 112898 262556 112904 262608
rect 112956 262596 112962 262608
rect 139394 262596 139400 262608
rect 112956 262568 139400 262596
rect 112956 262556 112962 262568
rect 139394 262556 139400 262568
rect 139452 262556 139458 262608
rect 165522 262556 165528 262608
rect 165580 262596 165586 262608
rect 192110 262596 192116 262608
rect 165580 262568 192116 262596
rect 165580 262556 165586 262568
rect 192110 262556 192116 262568
rect 192168 262556 192174 262608
rect 119890 262488 119896 262540
rect 119948 262528 119954 262540
rect 147674 262528 147680 262540
rect 119948 262500 147680 262528
rect 119948 262488 119954 262500
rect 147674 262488 147680 262500
rect 147732 262488 147738 262540
rect 172238 262488 172244 262540
rect 172296 262528 172302 262540
rect 198734 262528 198740 262540
rect 172296 262500 198740 262528
rect 172296 262488 172302 262500
rect 198734 262488 198740 262500
rect 198792 262528 198798 262540
rect 199194 262528 199200 262540
rect 198792 262500 199200 262528
rect 198792 262488 198798 262500
rect 199194 262488 199200 262500
rect 199252 262488 199258 262540
rect 114094 262420 114100 262472
rect 114152 262460 114158 262472
rect 142614 262460 142620 262472
rect 114152 262432 142620 262460
rect 114152 262420 114158 262432
rect 142614 262420 142620 262432
rect 142672 262420 142678 262472
rect 168926 262420 168932 262472
rect 168984 262460 168990 262472
rect 196618 262460 196624 262472
rect 168984 262432 196624 262460
rect 168984 262420 168990 262432
rect 196618 262420 196624 262432
rect 196676 262420 196682 262472
rect 115290 262352 115296 262404
rect 115348 262392 115354 262404
rect 115348 262364 125594 262392
rect 115348 262352 115354 262364
rect 125566 262324 125594 262364
rect 126974 262352 126980 262404
rect 127032 262392 127038 262404
rect 135254 262392 135260 262404
rect 127032 262364 135260 262392
rect 127032 262352 127038 262364
rect 135254 262352 135260 262364
rect 135312 262352 135318 262404
rect 179874 262352 179880 262404
rect 179932 262392 179938 262404
rect 190638 262392 190644 262404
rect 179932 262364 190644 262392
rect 179932 262352 179938 262364
rect 190638 262352 190644 262364
rect 190696 262352 190702 262404
rect 127710 262324 127716 262336
rect 125566 262296 127716 262324
rect 127710 262284 127716 262296
rect 127768 262284 127774 262336
rect 132770 262324 132776 262336
rect 127820 262296 132776 262324
rect 116854 262216 116860 262268
rect 116912 262256 116918 262268
rect 125226 262256 125232 262268
rect 116912 262228 125232 262256
rect 116912 262216 116918 262228
rect 125226 262216 125232 262228
rect 125284 262216 125290 262268
rect 127820 262256 127848 262296
rect 132770 262284 132776 262296
rect 132828 262284 132834 262336
rect 135438 262284 135444 262336
rect 135496 262324 135502 262336
rect 137646 262324 137652 262336
rect 135496 262296 137652 262324
rect 135496 262284 135502 262296
rect 137646 262284 137652 262296
rect 137704 262284 137710 262336
rect 187602 262284 187608 262336
rect 187660 262324 187666 262336
rect 211154 262324 211160 262336
rect 187660 262296 211160 262324
rect 187660 262284 187666 262296
rect 211154 262284 211160 262296
rect 211212 262284 211218 262336
rect 125336 262228 127848 262256
rect 119706 262148 119712 262200
rect 119764 262188 119770 262200
rect 125336 262188 125364 262228
rect 127894 262216 127900 262268
rect 127952 262256 127958 262268
rect 136818 262256 136824 262268
rect 127952 262228 136824 262256
rect 127952 262216 127958 262228
rect 136818 262216 136824 262228
rect 136876 262216 136882 262268
rect 177942 262216 177948 262268
rect 178000 262256 178006 262268
rect 192202 262256 192208 262268
rect 178000 262228 192208 262256
rect 178000 262216 178006 262228
rect 192202 262216 192208 262228
rect 192260 262216 192266 262268
rect 119764 262160 125364 262188
rect 119764 262148 119770 262160
rect 53098 260992 53104 261044
rect 53156 261032 53162 261044
rect 179874 261032 179880 261044
rect 53156 261004 179880 261032
rect 53156 260992 53162 261004
rect 179874 260992 179880 261004
rect 179932 260992 179938 261044
rect 182082 260992 182088 261044
rect 182140 261032 182146 261044
rect 197446 261032 197452 261044
rect 182140 261004 197452 261032
rect 182140 260992 182146 261004
rect 197446 260992 197452 261004
rect 197504 260992 197510 261044
rect 114370 260924 114376 260976
rect 114428 260964 114434 260976
rect 189074 260964 189080 260976
rect 114428 260936 189080 260964
rect 114428 260924 114434 260936
rect 189074 260924 189080 260936
rect 189132 260924 189138 260976
rect 176378 260856 176384 260908
rect 176436 260896 176442 260908
rect 192754 260896 192760 260908
rect 176436 260868 192760 260896
rect 176436 260856 176442 260868
rect 192754 260856 192760 260868
rect 192812 260856 192818 260908
rect 577866 260856 577872 260908
rect 577924 260896 577930 260908
rect 580718 260896 580724 260908
rect 577924 260868 580724 260896
rect 577924 260856 577930 260868
rect 580718 260856 580724 260868
rect 580776 260856 580782 260908
rect 118602 260788 118608 260840
rect 118660 260828 118666 260840
rect 122834 260828 122840 260840
rect 118660 260800 122840 260828
rect 118660 260788 118666 260800
rect 122834 260788 122840 260800
rect 122892 260788 122898 260840
rect 118666 260324 132494 260352
rect 114002 260176 114008 260228
rect 114060 260216 114066 260228
rect 118666 260216 118694 260324
rect 126238 260216 126244 260228
rect 114060 260188 118694 260216
rect 123312 260188 126244 260216
rect 114060 260176 114066 260188
rect 111242 260108 111248 260160
rect 111300 260148 111306 260160
rect 123312 260148 123340 260188
rect 126238 260176 126244 260188
rect 126296 260176 126302 260228
rect 128446 260176 128452 260228
rect 128504 260216 128510 260228
rect 129688 260216 129694 260228
rect 128504 260188 129694 260216
rect 128504 260176 128510 260188
rect 129688 260176 129694 260188
rect 129746 260176 129752 260228
rect 132466 260216 132494 260324
rect 158162 260312 158168 260364
rect 158220 260352 158226 260364
rect 191190 260352 191196 260364
rect 158220 260324 191196 260352
rect 158220 260312 158226 260324
rect 191190 260312 191196 260324
rect 191248 260312 191254 260364
rect 156046 260244 156052 260296
rect 156104 260284 156110 260296
rect 190730 260284 190736 260296
rect 156104 260256 190736 260284
rect 156104 260244 156110 260256
rect 190730 260244 190736 260256
rect 190788 260244 190794 260296
rect 144592 260216 144598 260228
rect 132466 260188 144598 260216
rect 144592 260176 144598 260188
rect 144650 260176 144656 260228
rect 161152 260176 161158 260228
rect 161210 260216 161216 260228
rect 196434 260216 196440 260228
rect 161210 260188 196440 260216
rect 161210 260176 161216 260188
rect 196434 260176 196440 260188
rect 196492 260176 196498 260228
rect 127204 260148 127210 260160
rect 111300 260120 123340 260148
rect 123404 260120 127210 260148
rect 111300 260108 111306 260120
rect 116670 260040 116676 260092
rect 116728 260080 116734 260092
rect 123404 260080 123432 260120
rect 127204 260108 127210 260120
rect 127262 260108 127268 260160
rect 128464 260148 128492 260176
rect 128326 260120 128492 260148
rect 116728 260052 123432 260080
rect 116728 260040 116734 260052
rect 117866 259972 117872 260024
rect 117924 260012 117930 260024
rect 128326 260012 128354 260120
rect 158668 260108 158674 260160
rect 158726 260148 158732 260160
rect 193674 260148 193680 260160
rect 158726 260120 193680 260148
rect 158726 260108 158732 260120
rect 193674 260108 193680 260120
rect 193732 260108 193738 260160
rect 149560 260080 149566 260092
rect 117924 259984 128354 260012
rect 132466 260052 149566 260080
rect 117924 259972 117930 259984
rect 124030 259904 124036 259956
rect 124088 259944 124094 259956
rect 132466 259944 132494 260052
rect 149560 260040 149566 260052
rect 149618 260040 149624 260092
rect 182680 260040 182686 260092
rect 182738 260080 182744 260092
rect 195054 260080 195060 260092
rect 182738 260052 195060 260080
rect 182738 260040 182744 260052
rect 195054 260040 195060 260052
rect 195112 260040 195118 260092
rect 181346 259972 181352 260024
rect 181404 260012 181410 260024
rect 197906 260012 197912 260024
rect 181404 259984 197912 260012
rect 181404 259972 181410 259984
rect 197906 259972 197912 259984
rect 197964 259972 197970 260024
rect 124088 259916 132494 259944
rect 124088 259904 124094 259916
rect 168098 259904 168104 259956
rect 168156 259944 168162 259956
rect 192662 259944 192668 259956
rect 168156 259916 192668 259944
rect 168156 259904 168162 259916
rect 192662 259904 192668 259916
rect 192720 259904 192726 259956
rect 112622 259836 112628 259888
rect 112680 259876 112686 259888
rect 126054 259876 126060 259888
rect 112680 259848 126060 259876
rect 112680 259836 112686 259848
rect 126054 259836 126060 259848
rect 126112 259836 126118 259888
rect 169754 259836 169760 259888
rect 169812 259876 169818 259888
rect 170950 259876 170956 259888
rect 169812 259848 170956 259876
rect 169812 259836 169818 259848
rect 170950 259836 170956 259848
rect 171008 259876 171014 259888
rect 196250 259876 196256 259888
rect 171008 259848 196256 259876
rect 171008 259836 171014 259848
rect 196250 259836 196256 259848
rect 196308 259836 196314 259888
rect 112346 259768 112352 259820
rect 112404 259808 112410 259820
rect 128354 259808 128360 259820
rect 112404 259780 128360 259808
rect 112404 259768 112410 259780
rect 128354 259768 128360 259780
rect 128412 259768 128418 259820
rect 166442 259768 166448 259820
rect 166500 259808 166506 259820
rect 196342 259808 196348 259820
rect 166500 259780 196348 259808
rect 166500 259768 166506 259780
rect 196342 259768 196348 259780
rect 196400 259768 196406 259820
rect 111150 259700 111156 259752
rect 111208 259740 111214 259752
rect 131114 259740 131120 259752
rect 111208 259712 131120 259740
rect 111208 259700 111214 259712
rect 131114 259700 131120 259712
rect 131172 259740 131178 259752
rect 131850 259740 131856 259752
rect 131172 259712 131856 259740
rect 131172 259700 131178 259712
rect 131850 259700 131856 259712
rect 131908 259700 131914 259752
rect 163958 259700 163964 259752
rect 164016 259740 164022 259752
rect 193766 259740 193772 259752
rect 164016 259712 193772 259740
rect 164016 259700 164022 259712
rect 193766 259700 193772 259712
rect 193824 259700 193830 259752
rect 113634 259632 113640 259684
rect 113692 259672 113698 259684
rect 135990 259672 135996 259684
rect 113692 259644 135996 259672
rect 113692 259632 113698 259644
rect 135990 259632 135996 259644
rect 136048 259632 136054 259684
rect 184658 259632 184664 259684
rect 184716 259672 184722 259684
rect 196158 259672 196164 259684
rect 184716 259644 196164 259672
rect 184716 259632 184722 259644
rect 196158 259632 196164 259644
rect 196216 259632 196222 259684
rect 115106 259564 115112 259616
rect 115164 259604 115170 259616
rect 123570 259604 123576 259616
rect 115164 259576 123576 259604
rect 115164 259564 115170 259576
rect 123570 259564 123576 259576
rect 123628 259604 123634 259616
rect 124858 259604 124864 259616
rect 123628 259576 124864 259604
rect 123628 259564 123634 259576
rect 124858 259564 124864 259576
rect 124916 259564 124922 259616
rect 178862 259564 178868 259616
rect 178920 259604 178926 259616
rect 198918 259604 198924 259616
rect 178920 259576 198924 259604
rect 178920 259564 178926 259576
rect 198918 259564 198924 259576
rect 198976 259564 198982 259616
rect 118326 259496 118332 259548
rect 118384 259536 118390 259548
rect 150894 259536 150900 259548
rect 118384 259508 150900 259536
rect 118384 259496 118390 259508
rect 150894 259496 150900 259508
rect 150952 259496 150958 259548
rect 175366 259496 175372 259548
rect 175424 259536 175430 259548
rect 189626 259536 189632 259548
rect 175424 259508 189632 259536
rect 175424 259496 175430 259508
rect 189626 259496 189632 259508
rect 189684 259496 189690 259548
rect 3050 259428 3056 259480
rect 3108 259468 3114 259480
rect 101674 259468 101680 259480
rect 3108 259440 101680 259468
rect 3108 259428 3114 259440
rect 101674 259428 101680 259440
rect 101732 259428 101738 259480
rect 119246 259428 119252 259480
rect 119304 259468 119310 259480
rect 124398 259468 124404 259480
rect 119304 259440 124404 259468
rect 119304 259428 119310 259440
rect 124398 259428 124404 259440
rect 124456 259428 124462 259480
rect 173802 259428 173808 259480
rect 173860 259468 173866 259480
rect 194870 259468 194876 259480
rect 173860 259440 194876 259468
rect 173860 259428 173866 259440
rect 194870 259428 194876 259440
rect 194928 259428 194934 259480
rect 116762 259292 116768 259344
rect 116820 259332 116826 259344
rect 124030 259332 124036 259344
rect 116820 259304 124036 259332
rect 116820 259292 116826 259304
rect 124030 259292 124036 259304
rect 124088 259292 124094 259344
rect 120074 259224 120080 259276
rect 120132 259264 120138 259276
rect 121270 259264 121276 259276
rect 120132 259236 121276 259264
rect 120132 259224 120138 259236
rect 121270 259224 121276 259236
rect 121328 259224 121334 259276
rect 120442 258748 120448 258800
rect 120500 258788 120506 258800
rect 120994 258788 121000 258800
rect 120500 258760 121000 258788
rect 120500 258748 120506 258760
rect 120994 258748 121000 258760
rect 121052 258748 121058 258800
rect 3142 255280 3148 255332
rect 3200 255320 3206 255332
rect 117406 255320 117412 255332
rect 3200 255292 117412 255320
rect 3200 255280 3206 255292
rect 117406 255280 117412 255292
rect 117464 255280 117470 255332
rect 120166 253376 120172 253428
rect 120224 253376 120230 253428
rect 120074 253172 120080 253224
rect 120132 253212 120138 253224
rect 120184 253212 120212 253376
rect 120132 253184 120212 253212
rect 120132 253172 120138 253184
rect 192754 252560 192760 252612
rect 192812 252600 192818 252612
rect 196526 252600 196532 252612
rect 192812 252572 196532 252600
rect 192812 252560 192818 252572
rect 196526 252560 196532 252572
rect 196584 252600 196590 252612
rect 579798 252600 579804 252612
rect 196584 252572 579804 252600
rect 196584 252560 196590 252572
rect 579798 252560 579804 252572
rect 579856 252560 579862 252612
rect 3142 251200 3148 251252
rect 3200 251240 3206 251252
rect 119522 251240 119528 251252
rect 3200 251212 119528 251240
rect 3200 251200 3206 251212
rect 119522 251200 119528 251212
rect 119580 251200 119586 251252
rect 191282 248412 191288 248464
rect 191340 248452 191346 248464
rect 579798 248452 579804 248464
rect 191340 248424 579804 248452
rect 191340 248412 191346 248424
rect 579798 248412 579804 248424
rect 579856 248412 579862 248464
rect 3326 247052 3332 247104
rect 3384 247092 3390 247104
rect 96522 247092 96528 247104
rect 3384 247064 96528 247092
rect 3384 247052 3390 247064
rect 96522 247052 96528 247064
rect 96580 247052 96586 247104
rect 190086 244264 190092 244316
rect 190144 244304 190150 244316
rect 580166 244304 580172 244316
rect 190144 244276 580172 244304
rect 190144 244264 190150 244276
rect 580166 244264 580172 244276
rect 580224 244264 580230 244316
rect 3142 242904 3148 242956
rect 3200 242944 3206 242956
rect 119614 242944 119620 242956
rect 3200 242916 119620 242944
rect 3200 242904 3206 242916
rect 119614 242904 119620 242916
rect 119672 242904 119678 242956
rect 3326 240048 3332 240100
rect 3384 240088 3390 240100
rect 53098 240088 53104 240100
rect 3384 240060 53104 240088
rect 3384 240048 3390 240060
rect 53098 240048 53104 240060
rect 53156 240048 53162 240100
rect 191650 237396 191656 237448
rect 191708 237436 191714 237448
rect 580166 237436 580172 237448
rect 191708 237408 580172 237436
rect 191708 237396 191714 237408
rect 580166 237396 580172 237408
rect 580224 237396 580230 237448
rect 3326 235968 3332 236020
rect 3384 236008 3390 236020
rect 109678 236008 109684 236020
rect 3384 235980 109684 236008
rect 3384 235968 3390 235980
rect 109678 235968 109684 235980
rect 109736 235968 109742 236020
rect 3326 231820 3332 231872
rect 3384 231860 3390 231872
rect 112990 231860 112996 231872
rect 3384 231832 112996 231860
rect 3384 231820 3390 231832
rect 112990 231820 112996 231832
rect 113048 231820 113054 231872
rect 3326 227740 3332 227792
rect 3384 227780 3390 227792
rect 92474 227780 92480 227792
rect 3384 227752 92480 227780
rect 3384 227740 3390 227752
rect 92474 227740 92480 227752
rect 92532 227740 92538 227792
rect 3326 223592 3332 223644
rect 3384 223632 3390 223644
rect 120626 223632 120632 223644
rect 3384 223604 120632 223632
rect 3384 223592 3390 223604
rect 120626 223592 120632 223604
rect 120684 223592 120690 223644
rect 208394 220804 208400 220856
rect 208452 220844 208458 220856
rect 580166 220844 580172 220856
rect 208452 220816 580172 220844
rect 208452 220804 208458 220816
rect 580166 220804 580172 220816
rect 580224 220804 580230 220856
rect 3234 220736 3240 220788
rect 3292 220776 3298 220788
rect 114370 220776 114376 220788
rect 3292 220748 114376 220776
rect 3292 220736 3298 220748
rect 114370 220736 114376 220748
rect 114428 220736 114434 220788
rect 191190 217268 191196 217320
rect 191248 217308 191254 217320
rect 580166 217308 580172 217320
rect 191248 217280 580172 217308
rect 191248 217268 191254 217280
rect 580166 217268 580172 217280
rect 580224 217268 580230 217320
rect 3326 215296 3332 215348
rect 3384 215336 3390 215348
rect 96430 215336 96436 215348
rect 3384 215308 96436 215336
rect 3384 215296 3390 215308
rect 96430 215296 96436 215308
rect 96488 215336 96494 215348
rect 119154 215336 119160 215348
rect 96488 215308 119160 215336
rect 96488 215296 96494 215308
rect 119154 215296 119160 215308
rect 119212 215296 119218 215348
rect 190454 208904 190460 208956
rect 190512 208944 190518 208956
rect 190822 208944 190828 208956
rect 190512 208916 190828 208944
rect 190512 208904 190518 208916
rect 190822 208904 190828 208916
rect 190880 208904 190886 208956
rect 202782 206252 202788 206304
rect 202840 206292 202846 206304
rect 580626 206292 580632 206304
rect 202840 206264 580632 206292
rect 202840 206252 202846 206264
rect 580626 206252 580632 206264
rect 580684 206252 580690 206304
rect 191374 205640 191380 205692
rect 191432 205680 191438 205692
rect 201678 205680 201684 205692
rect 191432 205652 201684 205680
rect 191432 205640 191438 205652
rect 201678 205640 201684 205652
rect 201736 205680 201742 205692
rect 202782 205680 202788 205692
rect 201736 205652 202788 205680
rect 201736 205640 201742 205652
rect 202782 205640 202788 205652
rect 202840 205640 202846 205692
rect 576394 205572 576400 205624
rect 576452 205612 576458 205624
rect 579982 205612 579988 205624
rect 576452 205584 579988 205612
rect 576452 205572 576458 205584
rect 579982 205572 579988 205584
rect 580040 205572 580046 205624
rect 115934 202784 115940 202836
rect 115992 202824 115998 202836
rect 116578 202824 116584 202836
rect 115992 202796 116584 202824
rect 115992 202784 115998 202796
rect 116578 202784 116584 202796
rect 116636 202784 116642 202836
rect 96982 201560 96988 201612
rect 97040 201600 97046 201612
rect 116578 201600 116584 201612
rect 97040 201572 116584 201600
rect 97040 201560 97046 201572
rect 116578 201560 116584 201572
rect 116636 201560 116642 201612
rect 96338 201492 96344 201544
rect 96396 201532 96402 201544
rect 117406 201532 117412 201544
rect 96396 201504 117412 201532
rect 96396 201492 96402 201504
rect 117406 201492 117412 201504
rect 117464 201532 117470 201544
rect 117774 201532 117780 201544
rect 117464 201504 117780 201532
rect 117464 201492 117470 201504
rect 117774 201492 117780 201504
rect 117832 201492 117838 201544
rect 211062 200880 211068 200932
rect 211120 200920 211126 200932
rect 474734 200920 474740 200932
rect 211120 200892 474740 200920
rect 211120 200880 211126 200892
rect 474734 200880 474740 200892
rect 474792 200880 474798 200932
rect 191742 200812 191748 200864
rect 191800 200852 191806 200864
rect 204530 200852 204536 200864
rect 191800 200824 204536 200852
rect 191800 200812 191806 200824
rect 204530 200812 204536 200824
rect 204588 200812 204594 200864
rect 220998 200812 221004 200864
rect 221056 200852 221062 200864
rect 531314 200852 531320 200864
rect 221056 200824 531320 200852
rect 221056 200812 221062 200824
rect 531314 200812 531320 200824
rect 531372 200812 531378 200864
rect 3510 200744 3516 200796
rect 3568 200784 3574 200796
rect 92474 200784 92480 200796
rect 3568 200756 92480 200784
rect 3568 200744 3574 200756
rect 92474 200744 92480 200756
rect 92532 200744 92538 200796
rect 113818 200744 113824 200796
rect 113876 200784 113882 200796
rect 580718 200784 580724 200796
rect 113876 200756 153148 200784
rect 113876 200744 113882 200756
rect 115198 200676 115204 200728
rect 115256 200716 115262 200728
rect 115256 200688 150618 200716
rect 115256 200676 115262 200688
rect 119614 200608 119620 200660
rect 119672 200648 119678 200660
rect 131850 200648 131856 200660
rect 119672 200620 131856 200648
rect 119672 200608 119678 200620
rect 131850 200608 131856 200620
rect 131908 200608 131914 200660
rect 124186 200416 141786 200444
rect 119430 200200 119436 200252
rect 119488 200240 119494 200252
rect 122834 200240 122840 200252
rect 119488 200212 122840 200240
rect 119488 200200 119494 200212
rect 122834 200200 122840 200212
rect 122892 200200 122898 200252
rect 92474 200132 92480 200184
rect 92532 200172 92538 200184
rect 93670 200172 93676 200184
rect 92532 200144 93676 200172
rect 92532 200132 92538 200144
rect 93670 200132 93676 200144
rect 93728 200172 93734 200184
rect 124186 200172 124214 200416
rect 132034 200336 132040 200388
rect 132092 200376 132098 200388
rect 132092 200348 137554 200376
rect 132092 200336 132098 200348
rect 124858 200200 124864 200252
rect 124916 200240 124922 200252
rect 124916 200212 136082 200240
rect 124916 200200 124922 200212
rect 93728 200144 124214 200172
rect 93728 200132 93734 200144
rect 131942 199928 131948 199980
rect 132000 199968 132006 199980
rect 132000 199940 134104 199968
rect 132000 199928 132006 199940
rect 128538 199860 128544 199912
rect 128596 199900 128602 199912
rect 131758 199900 131764 199912
rect 128596 199872 131764 199900
rect 128596 199860 128602 199872
rect 131758 199860 131764 199872
rect 131816 199860 131822 199912
rect 132218 199860 132224 199912
rect 132276 199900 132282 199912
rect 132816 199900 132822 199912
rect 132276 199872 132822 199900
rect 132276 199860 132282 199872
rect 132816 199860 132822 199872
rect 132874 199860 132880 199912
rect 133920 199860 133926 199912
rect 133978 199860 133984 199912
rect 117958 199792 117964 199844
rect 118016 199832 118022 199844
rect 124858 199832 124864 199844
rect 118016 199804 124864 199832
rect 118016 199792 118022 199804
rect 124858 199792 124864 199804
rect 124916 199792 124922 199844
rect 124950 199792 124956 199844
rect 125008 199832 125014 199844
rect 133276 199832 133282 199844
rect 125008 199804 133138 199832
rect 125008 199792 125014 199804
rect 133110 199776 133138 199804
rect 133248 199792 133282 199832
rect 133334 199792 133340 199844
rect 133644 199832 133650 199844
rect 133616 199792 133650 199832
rect 133702 199792 133708 199844
rect 133736 199792 133742 199844
rect 133794 199792 133800 199844
rect 110322 199724 110328 199776
rect 110380 199764 110386 199776
rect 110380 199736 122834 199764
rect 110380 199724 110386 199736
rect 88978 199588 88984 199640
rect 89036 199628 89042 199640
rect 108114 199628 108120 199640
rect 89036 199600 108120 199628
rect 89036 199588 89042 199600
rect 108114 199588 108120 199600
rect 108172 199588 108178 199640
rect 122806 199628 122834 199736
rect 132126 199724 132132 199776
rect 132184 199764 132190 199776
rect 132494 199764 132500 199776
rect 132184 199736 132500 199764
rect 132184 199724 132190 199736
rect 132494 199724 132500 199736
rect 132552 199724 132558 199776
rect 133000 199724 133006 199776
rect 133058 199724 133064 199776
rect 133092 199724 133098 199776
rect 133150 199724 133156 199776
rect 125502 199656 125508 199708
rect 125560 199696 125566 199708
rect 131666 199696 131672 199708
rect 125560 199668 131672 199696
rect 125560 199656 125566 199668
rect 131666 199656 131672 199668
rect 131724 199656 131730 199708
rect 122806 199600 131114 199628
rect 75914 199520 75920 199572
rect 75972 199560 75978 199572
rect 108206 199560 108212 199572
rect 75972 199532 108212 199560
rect 75972 199520 75978 199532
rect 108206 199520 108212 199532
rect 108264 199520 108270 199572
rect 118050 199520 118056 199572
rect 118108 199560 118114 199572
rect 124306 199560 124312 199572
rect 118108 199532 124312 199560
rect 118108 199520 118114 199532
rect 124306 199520 124312 199532
rect 124364 199560 124370 199572
rect 125502 199560 125508 199572
rect 124364 199532 125508 199560
rect 124364 199520 124370 199532
rect 125502 199520 125508 199532
rect 125560 199520 125566 199572
rect 71774 199452 71780 199504
rect 71832 199492 71838 199504
rect 131086 199492 131114 199600
rect 132218 199588 132224 199640
rect 132276 199628 132282 199640
rect 132770 199628 132776 199640
rect 132276 199600 132776 199628
rect 132276 199588 132282 199600
rect 132770 199588 132776 199600
rect 132828 199588 132834 199640
rect 131758 199520 131764 199572
rect 131816 199560 131822 199572
rect 133018 199560 133046 199724
rect 133248 199640 133276 199792
rect 133368 199724 133374 199776
rect 133426 199724 133432 199776
rect 133230 199588 133236 199640
rect 133288 199588 133294 199640
rect 131816 199532 133046 199560
rect 133386 199560 133414 199724
rect 133616 199640 133644 199792
rect 133754 199640 133782 199792
rect 133598 199588 133604 199640
rect 133656 199588 133662 199640
rect 133690 199588 133696 199640
rect 133748 199600 133782 199640
rect 133938 199628 133966 199860
rect 134076 199696 134104 199940
rect 134306 199940 134702 199968
rect 134306 199912 134334 199940
rect 134288 199860 134294 199912
rect 134346 199860 134352 199912
rect 134472 199900 134478 199912
rect 134444 199860 134478 199900
rect 134530 199860 134536 199912
rect 134564 199860 134570 199912
rect 134622 199860 134628 199912
rect 134444 199708 134472 199860
rect 134582 199708 134610 199860
rect 134334 199696 134340 199708
rect 134076 199668 134340 199696
rect 134334 199656 134340 199668
rect 134392 199656 134398 199708
rect 134426 199656 134432 199708
rect 134484 199656 134490 199708
rect 134518 199656 134524 199708
rect 134576 199668 134610 199708
rect 134576 199656 134582 199668
rect 134058 199628 134064 199640
rect 133938 199600 134064 199628
rect 133748 199588 133754 199600
rect 134058 199588 134064 199600
rect 134116 199588 134122 199640
rect 134242 199588 134248 199640
rect 134300 199628 134306 199640
rect 134674 199628 134702 199940
rect 136054 199912 136082 200212
rect 136698 200076 137416 200104
rect 136698 199912 136726 200076
rect 134840 199860 134846 199912
rect 134898 199860 134904 199912
rect 135116 199860 135122 199912
rect 135174 199860 135180 199912
rect 135300 199860 135306 199912
rect 135358 199860 135364 199912
rect 135392 199860 135398 199912
rect 135450 199860 135456 199912
rect 135484 199860 135490 199912
rect 135542 199860 135548 199912
rect 135668 199860 135674 199912
rect 135726 199860 135732 199912
rect 135760 199860 135766 199912
rect 135818 199860 135824 199912
rect 136036 199860 136042 199912
rect 136094 199860 136100 199912
rect 136404 199860 136410 199912
rect 136462 199860 136468 199912
rect 136588 199860 136594 199912
rect 136646 199860 136652 199912
rect 136680 199860 136686 199912
rect 136738 199860 136744 199912
rect 136772 199860 136778 199912
rect 136830 199860 136836 199912
rect 136864 199860 136870 199912
rect 136922 199860 136928 199912
rect 137140 199860 137146 199912
rect 137198 199860 137204 199912
rect 134858 199776 134886 199860
rect 134794 199724 134800 199776
rect 134852 199736 134886 199776
rect 134852 199724 134858 199736
rect 134932 199724 134938 199776
rect 134990 199724 134996 199776
rect 134950 199640 134978 199724
rect 134300 199600 134702 199628
rect 134300 199588 134306 199600
rect 134886 199588 134892 199640
rect 134944 199600 134978 199640
rect 134944 199588 134950 199600
rect 134334 199560 134340 199572
rect 133386 199532 134340 199560
rect 131816 199520 131822 199532
rect 134334 199520 134340 199532
rect 134392 199520 134398 199572
rect 134978 199520 134984 199572
rect 135036 199560 135042 199572
rect 135134 199560 135162 199860
rect 135318 199832 135346 199860
rect 135272 199804 135346 199832
rect 135272 199572 135300 199804
rect 135410 199776 135438 199860
rect 135346 199724 135352 199776
rect 135404 199736 135438 199776
rect 135404 199724 135410 199736
rect 135502 199708 135530 199860
rect 135686 199832 135714 199860
rect 135438 199656 135444 199708
rect 135496 199668 135530 199708
rect 135640 199804 135714 199832
rect 135496 199656 135502 199668
rect 135640 199628 135668 199804
rect 135778 199764 135806 199860
rect 135944 199792 135950 199844
rect 136002 199832 136008 199844
rect 136002 199804 136128 199832
rect 136002 199792 136008 199804
rect 135732 199736 135806 199764
rect 135732 199708 135760 199736
rect 135714 199656 135720 199708
rect 135772 199656 135778 199708
rect 135990 199696 135996 199708
rect 135824 199668 135996 199696
rect 135824 199628 135852 199668
rect 135990 199656 135996 199668
rect 136048 199656 136054 199708
rect 135640 199600 135852 199628
rect 135898 199588 135904 199640
rect 135956 199628 135962 199640
rect 136100 199628 136128 199804
rect 135956 199600 136128 199628
rect 136422 199640 136450 199860
rect 136606 199776 136634 199860
rect 136606 199736 136640 199776
rect 136634 199724 136640 199736
rect 136692 199724 136698 199776
rect 136422 199600 136456 199640
rect 135956 199588 135962 199600
rect 136450 199588 136456 199600
rect 136508 199588 136514 199640
rect 136790 199572 136818 199860
rect 136882 199696 136910 199860
rect 136882 199668 136956 199696
rect 136928 199572 136956 199668
rect 135036 199532 135162 199560
rect 135036 199520 135042 199532
rect 135254 199520 135260 199572
rect 135312 199520 135318 199572
rect 135622 199520 135628 199572
rect 135680 199560 135686 199572
rect 135806 199560 135812 199572
rect 135680 199532 135812 199560
rect 135680 199520 135686 199532
rect 135806 199520 135812 199532
rect 135864 199520 135870 199572
rect 136790 199532 136824 199572
rect 136818 199520 136824 199532
rect 136876 199520 136882 199572
rect 136910 199520 136916 199572
rect 136968 199520 136974 199572
rect 137002 199520 137008 199572
rect 137060 199560 137066 199572
rect 137158 199560 137186 199860
rect 137388 199640 137416 200076
rect 137526 199844 137554 200348
rect 138722 199940 139486 199968
rect 138722 199912 138750 199940
rect 137600 199860 137606 199912
rect 137658 199860 137664 199912
rect 137784 199860 137790 199912
rect 137842 199860 137848 199912
rect 137968 199900 137974 199912
rect 137940 199860 137974 199900
rect 138026 199900 138032 199912
rect 138612 199900 138618 199912
rect 138026 199872 138073 199900
rect 138026 199860 138032 199872
rect 138584 199860 138618 199900
rect 138670 199860 138676 199912
rect 138704 199860 138710 199912
rect 138762 199860 138768 199912
rect 139072 199860 139078 199912
rect 139130 199860 139136 199912
rect 137508 199792 137514 199844
rect 137566 199792 137572 199844
rect 137618 199708 137646 199860
rect 137802 199764 137830 199860
rect 137940 199776 137968 199860
rect 137554 199656 137560 199708
rect 137612 199668 137646 199708
rect 137756 199736 137830 199764
rect 137612 199656 137618 199668
rect 137370 199588 137376 199640
rect 137428 199588 137434 199640
rect 137756 199572 137784 199736
rect 137922 199724 137928 199776
rect 137980 199724 137986 199776
rect 138152 199724 138158 199776
rect 138210 199724 138216 199776
rect 138336 199724 138342 199776
rect 138394 199764 138400 199776
rect 138394 199724 138428 199764
rect 137830 199656 137836 199708
rect 137888 199696 137894 199708
rect 138170 199696 138198 199724
rect 137888 199668 138198 199696
rect 137888 199656 137894 199668
rect 138400 199572 138428 199724
rect 138584 199628 138612 199860
rect 138888 199832 138894 199844
rect 138676 199804 138894 199832
rect 138676 199776 138704 199804
rect 138888 199792 138894 199804
rect 138946 199792 138952 199844
rect 139090 199832 139118 199860
rect 139044 199804 139118 199832
rect 138658 199724 138664 199776
rect 138716 199724 138722 199776
rect 138750 199656 138756 199708
rect 138808 199696 138814 199708
rect 138934 199696 138940 199708
rect 138808 199668 138940 199696
rect 138808 199656 138814 199668
rect 138934 199656 138940 199668
rect 138992 199656 138998 199708
rect 139044 199640 139072 199804
rect 139164 199792 139170 199844
rect 139222 199792 139228 199844
rect 139348 199792 139354 199844
rect 139406 199792 139412 199844
rect 139182 199764 139210 199792
rect 139136 199736 139210 199764
rect 139136 199708 139164 199736
rect 139118 199656 139124 199708
rect 139176 199656 139182 199708
rect 139210 199656 139216 199708
rect 139268 199696 139274 199708
rect 139366 199696 139394 199792
rect 139268 199668 139394 199696
rect 139268 199656 139274 199668
rect 138842 199628 138848 199640
rect 138584 199600 138848 199628
rect 138842 199588 138848 199600
rect 138900 199588 138906 199640
rect 139026 199588 139032 199640
rect 139084 199588 139090 199640
rect 139302 199588 139308 199640
rect 139360 199628 139366 199640
rect 139458 199628 139486 199940
rect 139992 199860 139998 199912
rect 140050 199860 140056 199912
rect 140820 199900 140826 199912
rect 140378 199872 140826 199900
rect 139624 199832 139630 199844
rect 139596 199792 139630 199832
rect 139682 199792 139688 199844
rect 139596 199708 139624 199792
rect 140010 199708 140038 199860
rect 140176 199792 140182 199844
rect 140234 199792 140240 199844
rect 139578 199656 139584 199708
rect 139636 199656 139642 199708
rect 139946 199656 139952 199708
rect 140004 199668 140038 199708
rect 140004 199656 140010 199668
rect 140194 199640 140222 199792
rect 139360 199600 139486 199628
rect 139360 199588 139366 199600
rect 140130 199588 140136 199640
rect 140188 199600 140222 199640
rect 140188 199588 140194 199600
rect 140378 199572 140406 199872
rect 140820 199860 140826 199872
rect 140878 199860 140884 199912
rect 141096 199860 141102 199912
rect 141154 199860 141160 199912
rect 141372 199860 141378 199912
rect 141430 199860 141436 199912
rect 140452 199792 140458 199844
rect 140510 199832 140516 199844
rect 140510 199804 140636 199832
rect 140510 199792 140516 199804
rect 140498 199656 140504 199708
rect 140556 199656 140562 199708
rect 137060 199532 137186 199560
rect 137060 199520 137066 199532
rect 137738 199520 137744 199572
rect 137796 199520 137802 199572
rect 138382 199520 138388 199572
rect 138440 199520 138446 199572
rect 140314 199520 140320 199572
rect 140372 199532 140406 199572
rect 140372 199520 140378 199532
rect 71832 199464 128354 199492
rect 131086 199464 133184 199492
rect 71832 199452 71838 199464
rect 3418 199384 3424 199436
rect 3476 199424 3482 199436
rect 108758 199424 108764 199436
rect 3476 199396 108764 199424
rect 3476 199384 3482 199396
rect 108758 199384 108764 199396
rect 108816 199424 108822 199436
rect 108816 199396 113174 199424
rect 108816 199384 108822 199396
rect 113146 199288 113174 199396
rect 119338 199384 119344 199436
rect 119396 199424 119402 199436
rect 126790 199424 126796 199436
rect 119396 199396 126796 199424
rect 119396 199384 119402 199396
rect 126790 199384 126796 199396
rect 126848 199384 126854 199436
rect 128326 199424 128354 199464
rect 131206 199424 131212 199436
rect 128326 199396 131212 199424
rect 131206 199384 131212 199396
rect 131264 199424 131270 199436
rect 132218 199424 132224 199436
rect 131264 199396 132224 199424
rect 131264 199384 131270 199396
rect 132218 199384 132224 199396
rect 132276 199384 132282 199436
rect 133156 199424 133184 199464
rect 140222 199452 140228 199504
rect 140280 199492 140286 199504
rect 140516 199492 140544 199656
rect 140608 199504 140636 199804
rect 141114 199696 141142 199860
rect 140700 199668 141142 199696
rect 140700 199572 140728 199668
rect 141390 199628 141418 199860
rect 141758 199844 141786 200416
rect 142172 200008 143350 200036
rect 142016 199860 142022 199912
rect 142074 199860 142080 199912
rect 141464 199792 141470 199844
rect 141522 199792 141528 199844
rect 141740 199792 141746 199844
rect 141798 199792 141804 199844
rect 141924 199792 141930 199844
rect 141982 199792 141988 199844
rect 140884 199600 141418 199628
rect 141482 199628 141510 199792
rect 141482 199600 141740 199628
rect 140682 199520 140688 199572
rect 140740 199520 140746 199572
rect 140280 199464 140544 199492
rect 140280 199452 140286 199464
rect 140590 199452 140596 199504
rect 140648 199452 140654 199504
rect 140884 199492 140912 199600
rect 141712 199504 141740 199600
rect 141942 199504 141970 199792
rect 142034 199560 142062 199860
rect 142172 199640 142200 200008
rect 142356 199940 142982 199968
rect 142356 199640 142384 199940
rect 142568 199900 142574 199912
rect 142540 199860 142574 199900
rect 142626 199860 142632 199912
rect 142660 199860 142666 199912
rect 142718 199860 142724 199912
rect 142752 199860 142758 199912
rect 142810 199900 142816 199912
rect 142810 199872 142890 199900
rect 142810 199860 142816 199872
rect 142540 199708 142568 199860
rect 142522 199656 142528 199708
rect 142580 199656 142586 199708
rect 142678 199696 142706 199860
rect 142862 199764 142890 199872
rect 142954 199844 142982 199940
rect 143322 199912 143350 200008
rect 143782 200008 146662 200036
rect 143304 199860 143310 199912
rect 143362 199860 143368 199912
rect 143580 199860 143586 199912
rect 143638 199900 143644 199912
rect 143638 199872 143718 199900
rect 143638 199860 143644 199872
rect 142936 199792 142942 199844
rect 142994 199792 143000 199844
rect 143276 199804 143534 199832
rect 142862 199736 142936 199764
rect 142678 199668 142844 199696
rect 142816 199640 142844 199668
rect 142154 199588 142160 199640
rect 142212 199588 142218 199640
rect 142338 199588 142344 199640
rect 142396 199588 142402 199640
rect 142798 199588 142804 199640
rect 142856 199588 142862 199640
rect 142614 199560 142620 199572
rect 142034 199532 142620 199560
rect 142614 199520 142620 199532
rect 142672 199520 142678 199572
rect 142706 199520 142712 199572
rect 142764 199560 142770 199572
rect 142908 199560 142936 199736
rect 143120 199724 143126 199776
rect 143178 199764 143184 199776
rect 143178 199724 143212 199764
rect 142982 199656 142988 199708
rect 143040 199696 143046 199708
rect 143040 199668 143120 199696
rect 143040 199656 143046 199668
rect 143092 199640 143120 199668
rect 143184 199640 143212 199724
rect 143074 199588 143080 199640
rect 143132 199588 143138 199640
rect 143166 199588 143172 199640
rect 143224 199588 143230 199640
rect 142764 199532 142936 199560
rect 142764 199520 142770 199532
rect 143276 199504 143304 199804
rect 143506 199776 143534 199804
rect 143488 199724 143494 199776
rect 143546 199724 143552 199776
rect 143396 199656 143402 199708
rect 143454 199696 143460 199708
rect 143454 199656 143488 199696
rect 141418 199492 141424 199504
rect 140884 199464 141424 199492
rect 141418 199452 141424 199464
rect 141476 199452 141482 199504
rect 141694 199452 141700 199504
rect 141752 199452 141758 199504
rect 141878 199452 141884 199504
rect 141936 199464 141970 199504
rect 141936 199452 141942 199464
rect 143258 199452 143264 199504
rect 143316 199452 143322 199504
rect 143350 199452 143356 199504
rect 143408 199492 143414 199504
rect 143460 199492 143488 199656
rect 143534 199588 143540 199640
rect 143592 199628 143598 199640
rect 143690 199628 143718 199872
rect 143782 199844 143810 200008
rect 144132 199860 144138 199912
rect 144190 199860 144196 199912
rect 144408 199860 144414 199912
rect 144466 199860 144472 199912
rect 144868 199860 144874 199912
rect 144926 199860 144932 199912
rect 144960 199860 144966 199912
rect 145018 199860 145024 199912
rect 145144 199860 145150 199912
rect 145202 199860 145208 199912
rect 145236 199860 145242 199912
rect 145294 199860 145300 199912
rect 145328 199860 145334 199912
rect 145386 199860 145392 199912
rect 145420 199860 145426 199912
rect 145478 199860 145484 199912
rect 145512 199860 145518 199912
rect 145570 199900 145576 199912
rect 145570 199860 145604 199900
rect 145696 199860 145702 199912
rect 145754 199860 145760 199912
rect 145880 199900 145886 199912
rect 145852 199860 145886 199900
rect 145938 199860 145944 199912
rect 145972 199860 145978 199912
rect 146030 199860 146036 199912
rect 146064 199860 146070 199912
rect 146122 199860 146128 199912
rect 146248 199900 146254 199912
rect 146220 199860 146254 199900
rect 146306 199860 146312 199912
rect 146340 199860 146346 199912
rect 146398 199860 146404 199912
rect 146432 199860 146438 199912
rect 146490 199860 146496 199912
rect 146524 199860 146530 199912
rect 146582 199860 146588 199912
rect 143764 199792 143770 199844
rect 143822 199792 143828 199844
rect 143856 199724 143862 199776
rect 143914 199724 143920 199776
rect 143592 199600 143718 199628
rect 143592 199588 143598 199600
rect 143874 199572 143902 199724
rect 143874 199532 143908 199572
rect 143902 199520 143908 199532
rect 143960 199520 143966 199572
rect 144150 199560 144178 199860
rect 144426 199832 144454 199860
rect 144776 199832 144782 199844
rect 144426 199804 144500 199832
rect 144362 199724 144368 199776
rect 144420 199724 144426 199776
rect 144270 199588 144276 199640
rect 144328 199628 144334 199640
rect 144380 199628 144408 199724
rect 144328 199600 144408 199628
rect 144328 199588 144334 199600
rect 144472 199572 144500 199804
rect 144564 199804 144782 199832
rect 144362 199560 144368 199572
rect 144150 199532 144368 199560
rect 144362 199520 144368 199532
rect 144420 199520 144426 199572
rect 144454 199520 144460 199572
rect 144512 199520 144518 199572
rect 144564 199560 144592 199804
rect 144776 199792 144782 199804
rect 144834 199792 144840 199844
rect 144886 199764 144914 199860
rect 144840 199736 144914 199764
rect 144840 199708 144868 199736
rect 144978 199708 145006 199860
rect 145162 199832 145190 199860
rect 144822 199656 144828 199708
rect 144880 199656 144886 199708
rect 144914 199656 144920 199708
rect 144972 199668 145006 199708
rect 145116 199804 145190 199832
rect 144972 199656 144978 199668
rect 145006 199560 145012 199572
rect 144564 199532 145012 199560
rect 145006 199520 145012 199532
rect 145064 199520 145070 199572
rect 143408 199464 143488 199492
rect 143408 199452 143414 199464
rect 143810 199452 143816 199504
rect 143868 199492 143874 199504
rect 145116 199492 145144 199804
rect 145254 199776 145282 199860
rect 145190 199724 145196 199776
rect 145248 199736 145282 199776
rect 145248 199724 145254 199736
rect 145346 199640 145374 199860
rect 145438 199696 145466 199860
rect 145576 199708 145604 199860
rect 145714 199708 145742 199860
rect 145438 199668 145512 199696
rect 145346 199600 145380 199640
rect 145374 199588 145380 199600
rect 145432 199588 145438 199640
rect 145282 199520 145288 199572
rect 145340 199560 145346 199572
rect 145484 199560 145512 199668
rect 145558 199656 145564 199708
rect 145616 199656 145622 199708
rect 145650 199656 145656 199708
rect 145708 199668 145742 199708
rect 145708 199656 145714 199668
rect 145852 199640 145880 199860
rect 145990 199832 146018 199860
rect 145944 199804 146018 199832
rect 145944 199640 145972 199804
rect 146082 199708 146110 199860
rect 146220 199776 146248 199860
rect 146358 199832 146386 199860
rect 146312 199804 146386 199832
rect 146312 199776 146340 199804
rect 146450 199776 146478 199860
rect 146202 199724 146208 199776
rect 146260 199724 146266 199776
rect 146294 199724 146300 199776
rect 146352 199724 146358 199776
rect 146386 199724 146392 199776
rect 146444 199736 146478 199776
rect 146444 199724 146450 199736
rect 146018 199656 146024 199708
rect 146076 199668 146110 199708
rect 146076 199656 146082 199668
rect 145834 199588 145840 199640
rect 145892 199588 145898 199640
rect 145926 199588 145932 199640
rect 145984 199588 145990 199640
rect 146542 199572 146570 199860
rect 145340 199532 145512 199560
rect 145340 199520 145346 199532
rect 146478 199520 146484 199572
rect 146536 199532 146570 199572
rect 146536 199520 146542 199532
rect 143868 199464 145144 199492
rect 146634 199492 146662 200008
rect 146772 199940 147766 199968
rect 146772 199572 146800 199940
rect 147738 199912 147766 199940
rect 148612 199940 150388 199968
rect 147076 199860 147082 199912
rect 147134 199860 147140 199912
rect 147536 199860 147542 199912
rect 147594 199860 147600 199912
rect 147720 199860 147726 199912
rect 147778 199860 147784 199912
rect 147904 199860 147910 199912
rect 147962 199860 147968 199912
rect 147996 199860 148002 199912
rect 148054 199860 148060 199912
rect 148364 199860 148370 199912
rect 148422 199860 148428 199912
rect 146754 199520 146760 199572
rect 146812 199520 146818 199572
rect 146846 199492 146852 199504
rect 146634 199464 146852 199492
rect 143868 199452 143874 199464
rect 146846 199452 146852 199464
rect 146904 199452 146910 199504
rect 147094 199492 147122 199860
rect 147554 199832 147582 199860
rect 147554 199804 147720 199832
rect 147692 199640 147720 199804
rect 147766 199724 147772 199776
rect 147824 199764 147830 199776
rect 147922 199764 147950 199860
rect 147824 199736 147950 199764
rect 147824 199724 147830 199736
rect 147674 199588 147680 199640
rect 147732 199588 147738 199640
rect 148014 199628 148042 199860
rect 148382 199640 148410 199860
rect 148612 199640 148640 199940
rect 148732 199860 148738 199912
rect 148790 199860 148796 199912
rect 149008 199900 149014 199912
rect 148980 199860 149014 199900
rect 149066 199900 149072 199912
rect 149066 199872 149113 199900
rect 149066 199860 149072 199872
rect 149744 199860 149750 199912
rect 149802 199900 149808 199912
rect 149802 199872 150296 199900
rect 149802 199860 149808 199872
rect 148134 199628 148140 199640
rect 148014 199600 148140 199628
rect 148134 199588 148140 199600
rect 148192 199588 148198 199640
rect 148382 199600 148416 199640
rect 148410 199588 148416 199600
rect 148468 199588 148474 199640
rect 148594 199588 148600 199640
rect 148652 199588 148658 199640
rect 148750 199628 148778 199860
rect 148870 199628 148876 199640
rect 148750 199600 148876 199628
rect 148870 199588 148876 199600
rect 148928 199588 148934 199640
rect 148980 199560 149008 199860
rect 149284 199792 149290 199844
rect 149342 199792 149348 199844
rect 149376 199792 149382 199844
rect 149434 199832 149440 199844
rect 149434 199804 149928 199832
rect 149434 199792 149440 199804
rect 149302 199640 149330 199792
rect 149422 199656 149428 199708
rect 149480 199656 149486 199708
rect 149302 199600 149336 199640
rect 149330 199588 149336 199600
rect 149388 199588 149394 199640
rect 149440 199560 149468 199656
rect 149606 199560 149612 199572
rect 148980 199532 149376 199560
rect 149440 199532 149612 199560
rect 149348 199504 149376 199532
rect 149606 199520 149612 199532
rect 149664 199520 149670 199572
rect 149900 199504 149928 199804
rect 150020 199724 150026 199776
rect 150078 199724 150084 199776
rect 150038 199504 150066 199724
rect 147398 199492 147404 199504
rect 147094 199464 147404 199492
rect 147398 199452 147404 199464
rect 147456 199452 147462 199504
rect 149330 199452 149336 199504
rect 149388 199452 149394 199504
rect 149882 199452 149888 199504
rect 149940 199452 149946 199504
rect 149974 199452 149980 199504
rect 150032 199464 150066 199504
rect 150268 199492 150296 199872
rect 150360 199572 150388 199940
rect 150480 199832 150486 199844
rect 150452 199792 150486 199832
rect 150538 199792 150544 199844
rect 150452 199572 150480 199792
rect 150342 199520 150348 199572
rect 150400 199520 150406 199572
rect 150434 199520 150440 199572
rect 150492 199520 150498 199572
rect 150590 199560 150618 200688
rect 151234 199940 152274 199968
rect 151032 199832 151038 199844
rect 150820 199804 151038 199832
rect 150820 199628 150848 199804
rect 151032 199792 151038 199804
rect 151090 199792 151096 199844
rect 150986 199628 150992 199640
rect 150820 199600 150992 199628
rect 150986 199588 150992 199600
rect 151044 199588 151050 199640
rect 151234 199628 151262 199940
rect 152246 199912 152274 199940
rect 151676 199860 151682 199912
rect 151734 199900 151740 199912
rect 151734 199872 151906 199900
rect 151734 199860 151740 199872
rect 151400 199832 151406 199844
rect 151188 199600 151262 199628
rect 151372 199792 151406 199832
rect 151458 199792 151464 199844
rect 151492 199792 151498 199844
rect 151550 199792 151556 199844
rect 150590 199532 150848 199560
rect 150268 199464 150756 199492
rect 150032 199452 150038 199464
rect 150728 199436 150756 199464
rect 147950 199424 147956 199436
rect 133156 199396 147956 199424
rect 147950 199384 147956 199396
rect 148008 199384 148014 199436
rect 148502 199384 148508 199436
rect 148560 199424 148566 199436
rect 150526 199424 150532 199436
rect 148560 199396 150532 199424
rect 148560 199384 148566 199396
rect 150526 199384 150532 199396
rect 150584 199384 150590 199436
rect 150710 199384 150716 199436
rect 150768 199384 150774 199436
rect 119430 199316 119436 199368
rect 119488 199356 119494 199368
rect 121914 199356 121920 199368
rect 119488 199328 121920 199356
rect 119488 199316 119494 199328
rect 121914 199316 121920 199328
rect 121972 199356 121978 199368
rect 148962 199356 148968 199368
rect 121972 199328 148968 199356
rect 121972 199316 121978 199328
rect 148962 199316 148968 199328
rect 149020 199316 149026 199368
rect 149348 199328 149560 199356
rect 140498 199288 140504 199300
rect 113146 199260 140504 199288
rect 140498 199248 140504 199260
rect 140556 199248 140562 199300
rect 144086 199248 144092 199300
rect 144144 199288 144150 199300
rect 149348 199288 149376 199328
rect 144144 199260 149376 199288
rect 149532 199288 149560 199328
rect 150342 199316 150348 199368
rect 150400 199356 150406 199368
rect 150820 199356 150848 199532
rect 150400 199328 150848 199356
rect 151188 199356 151216 199600
rect 151372 199504 151400 199792
rect 151510 199708 151538 199792
rect 151878 199764 151906 199872
rect 151952 199860 151958 199912
rect 152010 199860 152016 199912
rect 152228 199860 152234 199912
rect 152286 199860 152292 199912
rect 152320 199860 152326 199912
rect 152378 199860 152384 199912
rect 152504 199860 152510 199912
rect 152562 199860 152568 199912
rect 152596 199860 152602 199912
rect 152654 199860 152660 199912
rect 152688 199860 152694 199912
rect 152746 199860 152752 199912
rect 152872 199860 152878 199912
rect 152930 199860 152936 199912
rect 151970 199832 151998 199860
rect 152338 199832 152366 199860
rect 151970 199804 152228 199832
rect 151878 199736 152136 199764
rect 151446 199656 151452 199708
rect 151504 199668 151538 199708
rect 151504 199656 151510 199668
rect 151722 199588 151728 199640
rect 151780 199628 151786 199640
rect 152108 199628 152136 199736
rect 151780 199600 152136 199628
rect 152200 199628 152228 199804
rect 152292 199804 152366 199832
rect 152292 199708 152320 199804
rect 152522 199776 152550 199860
rect 152458 199724 152464 199776
rect 152516 199736 152550 199776
rect 152516 199724 152522 199736
rect 152274 199656 152280 199708
rect 152332 199656 152338 199708
rect 152614 199640 152642 199860
rect 152366 199628 152372 199640
rect 152200 199600 152372 199628
rect 151780 199588 151786 199600
rect 152366 199588 152372 199600
rect 152424 199588 152430 199640
rect 152550 199588 152556 199640
rect 152608 199600 152642 199640
rect 152608 199588 152614 199600
rect 151906 199520 151912 199572
rect 151964 199560 151970 199572
rect 152706 199560 152734 199860
rect 152890 199640 152918 199860
rect 152826 199588 152832 199640
rect 152884 199600 152918 199640
rect 152884 199588 152890 199600
rect 151964 199532 152734 199560
rect 153120 199560 153148 200756
rect 154500 200756 180794 200784
rect 154500 199968 154528 200756
rect 178218 200716 178224 200728
rect 156064 200688 178224 200716
rect 156064 200308 156092 200688
rect 178218 200676 178224 200688
rect 178276 200676 178282 200728
rect 180766 200716 180794 200756
rect 181916 200756 580724 200784
rect 181916 200728 181944 200756
rect 580718 200744 580724 200756
rect 580776 200744 580782 200796
rect 180766 200688 181852 200716
rect 163010 200620 175734 200648
rect 155972 200280 156092 200308
rect 162826 200280 162946 200308
rect 155190 200212 155908 200240
rect 155190 200104 155218 200212
rect 155880 200172 155908 200212
rect 155972 200172 156000 200280
rect 155880 200144 156000 200172
rect 162826 200104 162854 200280
rect 153810 199940 154022 199968
rect 153810 199912 153838 199940
rect 153424 199860 153430 199912
rect 153482 199900 153488 199912
rect 153608 199900 153614 199912
rect 153482 199860 153516 199900
rect 153332 199792 153338 199844
rect 153390 199792 153396 199844
rect 153350 199640 153378 199792
rect 153488 199640 153516 199860
rect 153580 199860 153614 199900
rect 153666 199860 153672 199912
rect 153700 199860 153706 199912
rect 153758 199860 153764 199912
rect 153792 199860 153798 199912
rect 153850 199860 153856 199912
rect 153884 199860 153890 199912
rect 153942 199860 153948 199912
rect 153580 199708 153608 199860
rect 153718 199776 153746 199860
rect 153718 199736 153752 199776
rect 153746 199724 153752 199736
rect 153804 199724 153810 199776
rect 153562 199656 153568 199708
rect 153620 199656 153626 199708
rect 153902 199696 153930 199860
rect 153672 199668 153930 199696
rect 153286 199588 153292 199640
rect 153344 199600 153378 199640
rect 153344 199588 153350 199600
rect 153470 199588 153476 199640
rect 153528 199588 153534 199640
rect 153378 199560 153384 199572
rect 153120 199532 153384 199560
rect 151964 199520 151970 199532
rect 153378 199520 153384 199532
rect 153436 199520 153442 199572
rect 153672 199504 153700 199668
rect 153838 199588 153844 199640
rect 153896 199628 153902 199640
rect 153994 199628 154022 199940
rect 154224 199940 154528 199968
rect 154638 200076 155218 200104
rect 156984 200076 162854 200104
rect 154068 199860 154074 199912
rect 154126 199860 154132 199912
rect 153896 199600 154022 199628
rect 153896 199588 153902 199600
rect 153930 199520 153936 199572
rect 153988 199560 153994 199572
rect 154086 199560 154114 199860
rect 154224 199628 154252 199940
rect 154638 199912 154666 200076
rect 155098 199940 155402 199968
rect 154344 199860 154350 199912
rect 154402 199860 154408 199912
rect 154436 199860 154442 199912
rect 154494 199860 154500 199912
rect 154528 199860 154534 199912
rect 154586 199860 154592 199912
rect 154620 199860 154626 199912
rect 154678 199860 154684 199912
rect 154988 199860 154994 199912
rect 155046 199860 155052 199912
rect 154362 199708 154390 199860
rect 154298 199656 154304 199708
rect 154356 199668 154390 199708
rect 154454 199708 154482 199860
rect 154546 199764 154574 199860
rect 154546 199736 154620 199764
rect 154592 199708 154620 199736
rect 154454 199668 154488 199708
rect 154356 199656 154362 199668
rect 154482 199656 154488 199668
rect 154540 199656 154546 199708
rect 154574 199656 154580 199708
rect 154632 199656 154638 199708
rect 154850 199628 154856 199640
rect 154224 199600 154856 199628
rect 154850 199588 154856 199600
rect 154908 199588 154914 199640
rect 153988 199532 154114 199560
rect 153988 199520 153994 199532
rect 154758 199520 154764 199572
rect 154816 199560 154822 199572
rect 155006 199560 155034 199860
rect 154816 199532 155034 199560
rect 154816 199520 154822 199532
rect 151354 199452 151360 199504
rect 151412 199452 151418 199504
rect 151998 199452 152004 199504
rect 152056 199492 152062 199504
rect 152366 199492 152372 199504
rect 152056 199464 152372 199492
rect 152056 199452 152062 199464
rect 152366 199452 152372 199464
rect 152424 199452 152430 199504
rect 153654 199452 153660 199504
rect 153712 199452 153718 199504
rect 152642 199384 152648 199436
rect 152700 199424 152706 199436
rect 155098 199424 155126 199940
rect 155374 199912 155402 199940
rect 155558 199940 155770 199968
rect 155558 199912 155586 199940
rect 155264 199860 155270 199912
rect 155322 199860 155328 199912
rect 155356 199860 155362 199912
rect 155414 199860 155420 199912
rect 155448 199860 155454 199912
rect 155506 199860 155512 199912
rect 155540 199860 155546 199912
rect 155598 199860 155604 199912
rect 155632 199860 155638 199912
rect 155690 199860 155696 199912
rect 155282 199776 155310 199860
rect 155466 199776 155494 199860
rect 155282 199736 155316 199776
rect 155310 199724 155316 199736
rect 155368 199724 155374 199776
rect 155402 199724 155408 199776
rect 155460 199736 155494 199776
rect 155460 199724 155466 199736
rect 155650 199708 155678 199860
rect 155586 199656 155592 199708
rect 155644 199668 155678 199708
rect 155644 199656 155650 199668
rect 155494 199588 155500 199640
rect 155552 199628 155558 199640
rect 155742 199628 155770 199940
rect 156386 199940 156598 199968
rect 155908 199860 155914 199912
rect 155966 199860 155972 199912
rect 155552 199600 155770 199628
rect 155552 199588 155558 199600
rect 155926 199572 155954 199860
rect 155862 199520 155868 199572
rect 155920 199532 155954 199572
rect 155920 199520 155926 199532
rect 152700 199396 155126 199424
rect 156386 199436 156414 199940
rect 156570 199912 156598 199940
rect 156460 199860 156466 199912
rect 156518 199860 156524 199912
rect 156552 199860 156558 199912
rect 156610 199860 156616 199912
rect 156736 199860 156742 199912
rect 156794 199860 156800 199912
rect 156478 199776 156506 199860
rect 156478 199736 156512 199776
rect 156506 199724 156512 199736
rect 156564 199724 156570 199776
rect 156754 199640 156782 199860
rect 156984 199640 157012 200076
rect 160066 200008 161934 200036
rect 158502 199940 158852 199968
rect 158502 199912 158530 199940
rect 157104 199860 157110 199912
rect 157162 199860 157168 199912
rect 157196 199860 157202 199912
rect 157254 199860 157260 199912
rect 157380 199860 157386 199912
rect 157438 199860 157444 199912
rect 157564 199860 157570 199912
rect 157622 199860 157628 199912
rect 157748 199860 157754 199912
rect 157806 199900 157812 199912
rect 157932 199900 157938 199912
rect 157806 199860 157840 199900
rect 157122 199708 157150 199860
rect 157214 199764 157242 199860
rect 157214 199736 157288 199764
rect 157122 199668 157156 199708
rect 157150 199656 157156 199668
rect 157208 199656 157214 199708
rect 157260 199640 157288 199736
rect 156754 199600 156788 199640
rect 156782 199588 156788 199600
rect 156840 199588 156846 199640
rect 156966 199588 156972 199640
rect 157024 199588 157030 199640
rect 157242 199588 157248 199640
rect 157300 199588 157306 199640
rect 157398 199572 157426 199860
rect 157582 199640 157610 199860
rect 157812 199776 157840 199860
rect 157904 199860 157938 199900
rect 157990 199860 157996 199912
rect 158024 199860 158030 199912
rect 158082 199860 158088 199912
rect 158116 199860 158122 199912
rect 158174 199860 158180 199912
rect 158208 199860 158214 199912
rect 158266 199860 158272 199912
rect 158300 199860 158306 199912
rect 158358 199860 158364 199912
rect 158484 199860 158490 199912
rect 158542 199860 158548 199912
rect 158668 199860 158674 199912
rect 158726 199860 158732 199912
rect 157904 199776 157932 199860
rect 158042 199832 158070 199860
rect 157996 199804 158070 199832
rect 157794 199724 157800 199776
rect 157852 199724 157858 199776
rect 157886 199724 157892 199776
rect 157944 199724 157950 199776
rect 157996 199708 158024 199804
rect 158134 199776 158162 199860
rect 158070 199724 158076 199776
rect 158128 199736 158162 199776
rect 158226 199764 158254 199860
rect 158318 199832 158346 199860
rect 158318 199804 158484 199832
rect 158226 199736 158300 199764
rect 158128 199724 158134 199736
rect 157978 199656 157984 199708
rect 158036 199656 158042 199708
rect 157582 199600 157616 199640
rect 157610 199588 157616 199600
rect 157668 199588 157674 199640
rect 158162 199588 158168 199640
rect 158220 199628 158226 199640
rect 158272 199628 158300 199736
rect 158220 199600 158300 199628
rect 158220 199588 158226 199600
rect 157398 199532 157432 199572
rect 157426 199520 157432 199532
rect 157484 199520 157490 199572
rect 158254 199520 158260 199572
rect 158312 199560 158318 199572
rect 158456 199560 158484 199804
rect 158312 199532 158484 199560
rect 158312 199520 158318 199532
rect 156386 199396 156420 199436
rect 152700 199384 152706 199396
rect 156414 199384 156420 199396
rect 156472 199384 156478 199436
rect 158686 199424 158714 199860
rect 158824 199560 158852 199940
rect 160066 199912 160094 200008
rect 160802 199940 161750 199968
rect 160802 199912 160830 199940
rect 158944 199860 158950 199912
rect 159002 199900 159008 199912
rect 159128 199900 159134 199912
rect 159002 199860 159036 199900
rect 159008 199776 159036 199860
rect 159100 199860 159134 199900
rect 159186 199860 159192 199912
rect 159220 199860 159226 199912
rect 159278 199860 159284 199912
rect 159680 199860 159686 199912
rect 159738 199860 159744 199912
rect 159864 199860 159870 199912
rect 159922 199860 159928 199912
rect 160048 199860 160054 199912
rect 160106 199860 160112 199912
rect 160692 199860 160698 199912
rect 160750 199860 160756 199912
rect 160784 199860 160790 199912
rect 160842 199860 160848 199912
rect 160876 199860 160882 199912
rect 160934 199860 160940 199912
rect 161060 199860 161066 199912
rect 161118 199860 161124 199912
rect 161152 199860 161158 199912
rect 161210 199860 161216 199912
rect 161428 199860 161434 199912
rect 161486 199860 161492 199912
rect 159100 199776 159128 199860
rect 158990 199724 158996 199776
rect 159048 199724 159054 199776
rect 159082 199724 159088 199776
rect 159140 199724 159146 199776
rect 159238 199628 159266 199860
rect 159358 199628 159364 199640
rect 159238 199600 159364 199628
rect 159358 199588 159364 199600
rect 159416 199588 159422 199640
rect 158824 199532 158944 199560
rect 158806 199424 158812 199436
rect 158686 199396 158812 199424
rect 158806 199384 158812 199396
rect 158864 199384 158870 199436
rect 152366 199356 152372 199368
rect 151188 199328 152372 199356
rect 150400 199316 150406 199328
rect 152366 199316 152372 199328
rect 152424 199316 152430 199368
rect 153746 199316 153752 199368
rect 153804 199356 153810 199368
rect 153804 199328 154114 199356
rect 153804 199316 153810 199328
rect 149532 199260 153884 199288
rect 144144 199248 144150 199260
rect 132218 199180 132224 199232
rect 132276 199220 132282 199232
rect 153102 199220 153108 199232
rect 132276 199192 153108 199220
rect 132276 199180 132282 199192
rect 153102 199180 153108 199192
rect 153160 199180 153166 199232
rect 119522 199112 119528 199164
rect 119580 199152 119586 199164
rect 122926 199152 122932 199164
rect 119580 199124 122932 199152
rect 119580 199112 119586 199124
rect 122926 199112 122932 199124
rect 122984 199152 122990 199164
rect 143994 199152 144000 199164
rect 122984 199124 144000 199152
rect 122984 199112 122990 199124
rect 143994 199112 144000 199124
rect 144052 199112 144058 199164
rect 145650 199112 145656 199164
rect 145708 199152 145714 199164
rect 147858 199152 147864 199164
rect 145708 199124 147864 199152
rect 145708 199112 145714 199124
rect 147858 199112 147864 199124
rect 147916 199112 147922 199164
rect 147950 199112 147956 199164
rect 148008 199152 148014 199164
rect 148008 199124 149422 199152
rect 148008 199112 148014 199124
rect 119154 199044 119160 199096
rect 119212 199084 119218 199096
rect 148502 199084 148508 199096
rect 119212 199056 148508 199084
rect 119212 199044 119218 199056
rect 148502 199044 148508 199056
rect 148560 199044 148566 199096
rect 108114 198976 108120 199028
rect 108172 199016 108178 199028
rect 108942 199016 108948 199028
rect 108172 198988 108948 199016
rect 108172 198976 108178 198988
rect 108942 198976 108948 198988
rect 109000 199016 109006 199028
rect 142154 199016 142160 199028
rect 109000 198988 142160 199016
rect 109000 198976 109006 198988
rect 142154 198976 142160 198988
rect 142212 198976 142218 199028
rect 108206 198908 108212 198960
rect 108264 198948 108270 198960
rect 108850 198948 108856 198960
rect 108264 198920 108856 198948
rect 108264 198908 108270 198920
rect 108850 198908 108856 198920
rect 108908 198948 108914 198960
rect 142246 198948 142252 198960
rect 108908 198920 142252 198948
rect 108908 198908 108914 198920
rect 142246 198908 142252 198920
rect 142304 198908 142310 198960
rect 149394 198948 149422 199124
rect 149514 199112 149520 199164
rect 149572 199152 149578 199164
rect 149882 199152 149888 199164
rect 149572 199124 149888 199152
rect 149572 199112 149578 199124
rect 149882 199112 149888 199124
rect 149940 199112 149946 199164
rect 153856 199016 153884 199260
rect 154086 199084 154114 199328
rect 154390 199180 154396 199232
rect 154448 199220 154454 199232
rect 158916 199220 158944 199532
rect 159542 199384 159548 199436
rect 159600 199424 159606 199436
rect 159698 199424 159726 199860
rect 159882 199696 159910 199860
rect 160324 199832 160330 199844
rect 159836 199668 159910 199696
rect 160296 199792 160330 199832
rect 160382 199792 160388 199844
rect 160416 199792 160422 199844
rect 160474 199792 160480 199844
rect 159836 199640 159864 199668
rect 160296 199640 160324 199792
rect 159818 199588 159824 199640
rect 159876 199588 159882 199640
rect 160278 199588 160284 199640
rect 160336 199588 160342 199640
rect 160434 199560 160462 199792
rect 160710 199776 160738 199860
rect 160710 199736 160744 199776
rect 160738 199724 160744 199736
rect 160796 199724 160802 199776
rect 160894 199696 160922 199860
rect 160848 199668 160922 199696
rect 161078 199708 161106 199860
rect 161170 199776 161198 199860
rect 161336 199792 161342 199844
rect 161394 199792 161400 199844
rect 161170 199736 161204 199776
rect 161198 199724 161204 199736
rect 161256 199724 161262 199776
rect 161354 199708 161382 199792
rect 161078 199668 161112 199708
rect 160848 199572 160876 199668
rect 161106 199656 161112 199668
rect 161164 199656 161170 199708
rect 161290 199656 161296 199708
rect 161348 199668 161382 199708
rect 161348 199656 161354 199668
rect 161446 199640 161474 199860
rect 161612 199792 161618 199844
rect 161670 199792 161676 199844
rect 161382 199588 161388 199640
rect 161440 199600 161474 199640
rect 161440 199588 161446 199600
rect 159600 199396 159726 199424
rect 160112 199532 160462 199560
rect 160112 199424 160140 199532
rect 160830 199520 160836 199572
rect 160888 199520 160894 199572
rect 161630 199492 161658 199792
rect 160664 199464 161658 199492
rect 160370 199424 160376 199436
rect 160112 199396 160376 199424
rect 159600 199384 159606 199396
rect 160370 199384 160376 199396
rect 160428 199384 160434 199436
rect 160186 199316 160192 199368
rect 160244 199356 160250 199368
rect 160664 199356 160692 199464
rect 161722 199436 161750 199940
rect 161796 199860 161802 199912
rect 161854 199860 161860 199912
rect 161658 199384 161664 199436
rect 161716 199396 161750 199436
rect 161716 199384 161722 199396
rect 160244 199328 160692 199356
rect 160244 199316 160250 199328
rect 160922 199316 160928 199368
rect 160980 199356 160986 199368
rect 161814 199356 161842 199860
rect 161906 199560 161934 200008
rect 162090 199940 162394 199968
rect 162090 199628 162118 199940
rect 162366 199912 162394 199940
rect 162164 199860 162170 199912
rect 162222 199900 162228 199912
rect 162222 199872 162302 199900
rect 162222 199860 162228 199872
rect 162274 199696 162302 199872
rect 162348 199860 162354 199912
rect 162406 199860 162412 199912
rect 162440 199860 162446 199912
rect 162498 199860 162504 199912
rect 162532 199860 162538 199912
rect 162590 199900 162596 199912
rect 162590 199872 162854 199900
rect 162590 199860 162596 199872
rect 162458 199776 162486 199860
rect 162624 199832 162630 199844
rect 162394 199724 162400 199776
rect 162452 199736 162486 199776
rect 162596 199792 162630 199832
rect 162682 199792 162688 199844
rect 162452 199724 162458 199736
rect 162596 199708 162624 199792
rect 162486 199696 162492 199708
rect 162274 199668 162492 199696
rect 162486 199656 162492 199668
rect 162544 199656 162550 199708
rect 162578 199656 162584 199708
rect 162636 199656 162642 199708
rect 162210 199628 162216 199640
rect 162090 199600 162216 199628
rect 162210 199588 162216 199600
rect 162268 199588 162274 199640
rect 162118 199560 162124 199572
rect 161906 199532 162124 199560
rect 162118 199520 162124 199532
rect 162176 199520 162182 199572
rect 162826 199436 162854 199872
rect 162918 199492 162946 200280
rect 163010 199912 163038 200620
rect 175706 200512 175734 200620
rect 177850 200608 177856 200660
rect 177908 200648 177914 200660
rect 178034 200648 178040 200660
rect 177908 200620 178040 200648
rect 177908 200608 177914 200620
rect 178034 200608 178040 200620
rect 178092 200608 178098 200660
rect 181824 200648 181852 200688
rect 181898 200676 181904 200728
rect 181956 200676 181962 200728
rect 182818 200676 182824 200728
rect 182876 200716 182882 200728
rect 428458 200716 428464 200728
rect 182876 200688 428464 200716
rect 182876 200676 182882 200688
rect 428458 200676 428464 200688
rect 428516 200676 428522 200728
rect 191282 200648 191288 200660
rect 181824 200620 191288 200648
rect 191282 200608 191288 200620
rect 191340 200608 191346 200660
rect 177758 200540 177764 200592
rect 177816 200580 177822 200592
rect 179138 200580 179144 200592
rect 177816 200552 179144 200580
rect 177816 200540 177822 200552
rect 179138 200540 179144 200552
rect 179196 200540 179202 200592
rect 191742 200580 191748 200592
rect 186286 200552 191748 200580
rect 177942 200512 177948 200524
rect 175706 200484 177948 200512
rect 177942 200472 177948 200484
rect 178000 200472 178006 200524
rect 178586 200444 178592 200456
rect 174970 200416 178592 200444
rect 164206 200348 165614 200376
rect 164206 199968 164234 200348
rect 165586 200172 165614 200348
rect 165586 200144 166994 200172
rect 166966 200104 166994 200144
rect 166966 200076 168374 200104
rect 168346 200036 168374 200076
rect 168346 200008 171962 200036
rect 163654 199940 164234 199968
rect 164390 199940 164970 199968
rect 162992 199860 162998 199912
rect 163050 199860 163056 199912
rect 163084 199860 163090 199912
rect 163142 199860 163148 199912
rect 163176 199860 163182 199912
rect 163234 199860 163240 199912
rect 163360 199860 163366 199912
rect 163418 199860 163424 199912
rect 163452 199860 163458 199912
rect 163510 199860 163516 199912
rect 163102 199708 163130 199860
rect 163038 199656 163044 199708
rect 163096 199668 163130 199708
rect 163096 199656 163102 199668
rect 163194 199572 163222 199860
rect 163378 199832 163406 199860
rect 163332 199804 163406 199832
rect 163332 199640 163360 199804
rect 163470 199708 163498 199860
rect 163406 199656 163412 199708
rect 163464 199668 163498 199708
rect 163464 199656 163470 199668
rect 163314 199588 163320 199640
rect 163372 199588 163378 199640
rect 163130 199520 163136 199572
rect 163188 199532 163222 199572
rect 163654 199572 163682 199940
rect 163728 199860 163734 199912
rect 163786 199860 163792 199912
rect 164004 199860 164010 199912
rect 164062 199900 164068 199912
rect 164062 199860 164096 199900
rect 164280 199860 164286 199912
rect 164338 199860 164344 199912
rect 163746 199764 163774 199860
rect 163958 199764 163964 199776
rect 163746 199736 163964 199764
rect 163958 199724 163964 199736
rect 164016 199724 164022 199776
rect 163654 199532 163688 199572
rect 163188 199520 163194 199532
rect 163682 199520 163688 199532
rect 163740 199520 163746 199572
rect 164068 199492 164096 199860
rect 164298 199708 164326 199860
rect 164234 199656 164240 199708
rect 164292 199668 164326 199708
rect 164292 199656 164298 199668
rect 164234 199492 164240 199504
rect 162918 199464 164240 199492
rect 164234 199452 164240 199464
rect 164292 199452 164298 199504
rect 164390 199492 164418 199940
rect 164942 199912 164970 199940
rect 170094 199940 170444 199968
rect 170094 199912 170122 199940
rect 164464 199860 164470 199912
rect 164522 199860 164528 199912
rect 164648 199860 164654 199912
rect 164706 199860 164712 199912
rect 164924 199860 164930 199912
rect 164982 199860 164988 199912
rect 165200 199900 165206 199912
rect 165172 199860 165206 199900
rect 165258 199860 165264 199912
rect 165476 199900 165482 199912
rect 165310 199872 165482 199900
rect 164482 199776 164510 199860
rect 164482 199736 164516 199776
rect 164510 199724 164516 199736
rect 164568 199724 164574 199776
rect 164666 199628 164694 199860
rect 165172 199640 165200 199860
rect 165310 199640 165338 199872
rect 165476 199860 165482 199872
rect 165534 199860 165540 199912
rect 165752 199860 165758 199912
rect 165810 199860 165816 199912
rect 165936 199860 165942 199912
rect 165994 199860 166000 199912
rect 166028 199860 166034 199912
rect 166086 199860 166092 199912
rect 166212 199900 166218 199912
rect 166184 199860 166218 199900
rect 166270 199860 166276 199912
rect 166304 199860 166310 199912
rect 166362 199860 166368 199912
rect 166396 199860 166402 199912
rect 166454 199860 166460 199912
rect 166580 199860 166586 199912
rect 166638 199860 166644 199912
rect 166856 199860 166862 199912
rect 166914 199860 166920 199912
rect 166948 199860 166954 199912
rect 167006 199860 167012 199912
rect 167132 199860 167138 199912
rect 167190 199860 167196 199912
rect 167684 199860 167690 199912
rect 167742 199860 167748 199912
rect 168052 199860 168058 199912
rect 168110 199860 168116 199912
rect 168144 199860 168150 199912
rect 168202 199860 168208 199912
rect 168328 199860 168334 199912
rect 168386 199860 168392 199912
rect 168420 199860 168426 199912
rect 168478 199860 168484 199912
rect 168512 199860 168518 199912
rect 168570 199860 168576 199912
rect 168604 199860 168610 199912
rect 168662 199860 168668 199912
rect 168880 199860 168886 199912
rect 168938 199860 168944 199912
rect 168972 199860 168978 199912
rect 169030 199860 169036 199912
rect 169064 199860 169070 199912
rect 169122 199860 169128 199912
rect 169616 199860 169622 199912
rect 169674 199860 169680 199912
rect 169800 199860 169806 199912
rect 169858 199860 169864 199912
rect 169892 199860 169898 199912
rect 169950 199860 169956 199912
rect 169984 199860 169990 199912
rect 170042 199860 170048 199912
rect 170076 199860 170082 199912
rect 170134 199860 170140 199912
rect 170168 199860 170174 199912
rect 170226 199860 170232 199912
rect 165062 199628 165068 199640
rect 164666 199600 165068 199628
rect 165062 199588 165068 199600
rect 165120 199588 165126 199640
rect 165154 199588 165160 199640
rect 165212 199588 165218 199640
rect 165246 199588 165252 199640
rect 165304 199600 165338 199640
rect 165770 199640 165798 199860
rect 165770 199600 165804 199640
rect 165304 199588 165310 199600
rect 165798 199588 165804 199600
rect 165856 199588 165862 199640
rect 165954 199504 165982 199860
rect 166046 199560 166074 199860
rect 166184 199640 166212 199860
rect 166322 199832 166350 199860
rect 166276 199804 166350 199832
rect 166276 199776 166304 199804
rect 166414 199776 166442 199860
rect 166258 199724 166264 199776
rect 166316 199724 166322 199776
rect 166350 199724 166356 199776
rect 166408 199736 166442 199776
rect 166408 199724 166414 199736
rect 166598 199640 166626 199860
rect 166874 199832 166902 199860
rect 166166 199588 166172 199640
rect 166224 199588 166230 199640
rect 166534 199588 166540 199640
rect 166592 199600 166626 199640
rect 166828 199804 166902 199832
rect 166592 199588 166598 199600
rect 166828 199572 166856 199804
rect 166966 199776 166994 199860
rect 166902 199724 166908 199776
rect 166960 199736 166994 199776
rect 166960 199724 166966 199736
rect 167150 199696 167178 199860
rect 167592 199832 167598 199844
rect 167564 199792 167598 199832
rect 167650 199792 167656 199844
rect 167150 199668 167408 199696
rect 167380 199572 167408 199668
rect 167564 199640 167592 199792
rect 167546 199588 167552 199640
rect 167604 199588 167610 199640
rect 167702 199628 167730 199860
rect 168070 199696 168098 199860
rect 168162 199776 168190 199860
rect 168346 199832 168374 199860
rect 168300 199804 168374 199832
rect 168300 199776 168328 199804
rect 168162 199736 168196 199776
rect 168190 199724 168196 199736
rect 168248 199724 168254 199776
rect 168282 199724 168288 199776
rect 168340 199724 168346 199776
rect 168438 199708 168466 199860
rect 168530 199764 168558 199860
rect 168622 199832 168650 199860
rect 168622 199804 168696 199832
rect 168530 199736 168604 199764
rect 168070 199668 168144 199696
rect 168438 199668 168472 199708
rect 168006 199628 168012 199640
rect 167702 199600 168012 199628
rect 168006 199588 168012 199600
rect 168064 199588 168070 199640
rect 166718 199560 166724 199572
rect 166046 199532 166724 199560
rect 166718 199520 166724 199532
rect 166776 199520 166782 199572
rect 166810 199520 166816 199572
rect 166868 199520 166874 199572
rect 167362 199520 167368 199572
rect 167420 199520 167426 199572
rect 167730 199520 167736 199572
rect 167788 199560 167794 199572
rect 168116 199560 168144 199668
rect 168466 199656 168472 199668
rect 168524 199656 168530 199708
rect 168576 199572 168604 199736
rect 168668 199640 168696 199804
rect 168650 199588 168656 199640
rect 168708 199588 168714 199640
rect 168742 199588 168748 199640
rect 168800 199628 168806 199640
rect 168898 199628 168926 199860
rect 168800 199600 168926 199628
rect 168800 199588 168806 199600
rect 167788 199532 168144 199560
rect 167788 199520 167794 199532
rect 168558 199520 168564 199572
rect 168616 199520 168622 199572
rect 168834 199520 168840 199572
rect 168892 199560 168898 199572
rect 168990 199560 169018 199860
rect 168892 199532 169018 199560
rect 168892 199520 168898 199532
rect 169082 199504 169110 199860
rect 169634 199708 169662 199860
rect 169818 199776 169846 199860
rect 169754 199724 169760 199776
rect 169812 199736 169846 199776
rect 169812 199724 169818 199736
rect 169910 199708 169938 199860
rect 169634 199668 169668 199708
rect 169662 199656 169668 199668
rect 169720 199656 169726 199708
rect 169846 199656 169852 199708
rect 169904 199668 169938 199708
rect 169904 199656 169910 199668
rect 169570 199588 169576 199640
rect 169628 199628 169634 199640
rect 170002 199628 170030 199860
rect 170186 199776 170214 199860
rect 170122 199724 170128 199776
rect 170180 199736 170214 199776
rect 170180 199724 170186 199736
rect 169628 199600 170030 199628
rect 169628 199588 169634 199600
rect 170416 199504 170444 199940
rect 170646 199940 171640 199968
rect 170646 199912 170674 199940
rect 170628 199860 170634 199912
rect 170686 199860 170692 199912
rect 170812 199900 170818 199912
rect 170784 199860 170818 199900
rect 170870 199860 170876 199912
rect 170996 199860 171002 199912
rect 171054 199860 171060 199912
rect 171088 199860 171094 199912
rect 171146 199860 171152 199912
rect 171180 199860 171186 199912
rect 171238 199900 171244 199912
rect 171238 199872 171318 199900
rect 171238 199860 171244 199872
rect 170784 199776 170812 199860
rect 171014 199776 171042 199860
rect 171106 199832 171134 199860
rect 171106 199804 171180 199832
rect 171152 199776 171180 199804
rect 170766 199724 170772 199776
rect 170824 199724 170830 199776
rect 171014 199736 171048 199776
rect 171042 199724 171048 199736
rect 171100 199724 171106 199776
rect 171134 199724 171140 199776
rect 171192 199724 171198 199776
rect 171290 199504 171318 199872
rect 164786 199492 164792 199504
rect 164390 199464 164792 199492
rect 164786 199452 164792 199464
rect 164844 199452 164850 199504
rect 165954 199464 165988 199504
rect 165982 199452 165988 199464
rect 166040 199452 166046 199504
rect 169082 199464 169116 199504
rect 169110 199452 169116 199464
rect 169168 199452 169174 199504
rect 170398 199452 170404 199504
rect 170456 199452 170462 199504
rect 171290 199464 171324 199504
rect 171318 199452 171324 199464
rect 171376 199452 171382 199504
rect 171612 199436 171640 199940
rect 171934 199912 171962 200008
rect 172118 200008 174906 200036
rect 172118 199912 172146 200008
rect 172716 199940 173710 199968
rect 171732 199860 171738 199912
rect 171790 199860 171796 199912
rect 171916 199860 171922 199912
rect 171974 199860 171980 199912
rect 172100 199860 172106 199912
rect 172158 199860 172164 199912
rect 172284 199860 172290 199912
rect 172342 199860 172348 199912
rect 171750 199640 171778 199860
rect 171750 199600 171784 199640
rect 171778 199588 171784 199600
rect 171836 199588 171842 199640
rect 171934 199492 171962 199860
rect 172054 199588 172060 199640
rect 172112 199628 172118 199640
rect 172302 199628 172330 199860
rect 172112 199600 172330 199628
rect 172112 199588 172118 199600
rect 172514 199492 172520 199504
rect 171934 199464 172520 199492
rect 172514 199452 172520 199464
rect 172572 199452 172578 199504
rect 162026 199384 162032 199436
rect 162084 199424 162090 199436
rect 162302 199424 162308 199436
rect 162084 199396 162308 199424
rect 162084 199384 162090 199396
rect 162302 199384 162308 199396
rect 162360 199384 162366 199436
rect 162826 199396 162860 199436
rect 162854 199384 162860 199396
rect 162912 199384 162918 199436
rect 165890 199384 165896 199436
rect 165948 199424 165954 199436
rect 167914 199424 167920 199436
rect 165948 199396 167920 199424
rect 165948 199384 165954 199396
rect 167914 199384 167920 199396
rect 167972 199384 167978 199436
rect 168374 199384 168380 199436
rect 168432 199424 168438 199436
rect 168432 199396 171548 199424
rect 168432 199384 168438 199396
rect 167086 199356 167092 199368
rect 160980 199328 161750 199356
rect 161814 199328 167092 199356
rect 160980 199316 160986 199328
rect 161198 199248 161204 199300
rect 161256 199288 161262 199300
rect 161474 199288 161480 199300
rect 161256 199260 161480 199288
rect 161256 199248 161262 199260
rect 161474 199248 161480 199260
rect 161532 199248 161538 199300
rect 161722 199288 161750 199328
rect 167086 199316 167092 199328
rect 167144 199316 167150 199368
rect 167362 199316 167368 199368
rect 167420 199356 167426 199368
rect 167730 199356 167736 199368
rect 167420 199328 167736 199356
rect 167420 199316 167426 199328
rect 167730 199316 167736 199328
rect 167788 199316 167794 199368
rect 170214 199316 170220 199368
rect 170272 199356 170278 199368
rect 170582 199356 170588 199368
rect 170272 199328 170588 199356
rect 170272 199316 170278 199328
rect 170582 199316 170588 199328
rect 170640 199316 170646 199368
rect 171520 199356 171548 199396
rect 171594 199384 171600 199436
rect 171652 199384 171658 199436
rect 172716 199356 172744 199940
rect 173682 199912 173710 199940
rect 172836 199860 172842 199912
rect 172894 199860 172900 199912
rect 172928 199860 172934 199912
rect 172986 199860 172992 199912
rect 173020 199860 173026 199912
rect 173078 199860 173084 199912
rect 173296 199900 173302 199912
rect 173268 199860 173302 199900
rect 173354 199860 173360 199912
rect 173388 199860 173394 199912
rect 173446 199860 173452 199912
rect 173480 199860 173486 199912
rect 173538 199860 173544 199912
rect 173572 199860 173578 199912
rect 173630 199860 173636 199912
rect 173664 199860 173670 199912
rect 173722 199860 173728 199912
rect 173756 199860 173762 199912
rect 173814 199860 173820 199912
rect 173848 199860 173854 199912
rect 173906 199900 173912 199912
rect 173906 199872 173986 199900
rect 173906 199860 173912 199872
rect 172854 199776 172882 199860
rect 172790 199724 172796 199776
rect 172848 199736 172882 199776
rect 172848 199724 172854 199736
rect 172946 199560 172974 199860
rect 172900 199532 172974 199560
rect 172900 199424 172928 199532
rect 173038 199504 173066 199860
rect 173268 199776 173296 199860
rect 173406 199776 173434 199860
rect 173250 199724 173256 199776
rect 173308 199724 173314 199776
rect 173342 199724 173348 199776
rect 173400 199736 173434 199776
rect 173498 199776 173526 199860
rect 173590 199832 173618 199860
rect 173590 199804 173664 199832
rect 173636 199776 173664 199804
rect 173498 199736 173532 199776
rect 173400 199724 173406 199736
rect 173526 199724 173532 199736
rect 173584 199724 173590 199776
rect 173618 199724 173624 199776
rect 173676 199724 173682 199776
rect 173774 199696 173802 199860
rect 173360 199668 173802 199696
rect 173360 199560 173388 199668
rect 173710 199560 173716 199572
rect 173360 199532 173716 199560
rect 173710 199520 173716 199532
rect 173768 199520 173774 199572
rect 173958 199504 173986 199872
rect 174584 199860 174590 199912
rect 174642 199860 174648 199912
rect 174602 199640 174630 199860
rect 174602 199600 174636 199640
rect 174630 199588 174636 199600
rect 174688 199588 174694 199640
rect 174878 199560 174906 200008
rect 174970 199912 174998 200416
rect 178586 200404 178592 200416
rect 178644 200404 178650 200456
rect 186286 200376 186314 200552
rect 191742 200540 191748 200552
rect 191800 200540 191806 200592
rect 194502 200404 194508 200456
rect 194560 200444 194566 200456
rect 200114 200444 200120 200456
rect 194560 200416 200120 200444
rect 194560 200404 194566 200416
rect 200114 200404 200120 200416
rect 200172 200404 200178 200456
rect 176902 200348 186314 200376
rect 176902 200240 176930 200348
rect 190454 200336 190460 200388
rect 190512 200376 190518 200388
rect 191650 200376 191656 200388
rect 190512 200348 191656 200376
rect 190512 200336 190518 200348
rect 191650 200336 191656 200348
rect 191708 200376 191714 200388
rect 214098 200376 214104 200388
rect 191708 200348 214104 200376
rect 191708 200336 191714 200348
rect 214098 200336 214104 200348
rect 214156 200336 214162 200388
rect 177850 200308 177856 200320
rect 175614 200212 176930 200240
rect 177592 200280 177856 200308
rect 175614 199912 175642 200212
rect 177592 200172 177620 200280
rect 177850 200268 177856 200280
rect 177908 200268 177914 200320
rect 179046 200268 179052 200320
rect 179104 200308 179110 200320
rect 209958 200308 209964 200320
rect 179104 200280 209964 200308
rect 179104 200268 179110 200280
rect 209958 200268 209964 200280
rect 210016 200308 210022 200320
rect 211062 200308 211068 200320
rect 210016 200280 211068 200308
rect 210016 200268 210022 200280
rect 211062 200268 211068 200280
rect 211120 200268 211126 200320
rect 220998 200240 221004 200252
rect 175798 200144 177620 200172
rect 177868 200212 221004 200240
rect 175798 199912 175826 200144
rect 177868 200036 177896 200212
rect 220998 200200 221004 200212
rect 221056 200200 221062 200252
rect 177942 200132 177948 200184
rect 178000 200172 178006 200184
rect 188982 200172 188988 200184
rect 178000 200144 188988 200172
rect 178000 200132 178006 200144
rect 188982 200132 188988 200144
rect 189040 200172 189046 200184
rect 580166 200172 580172 200184
rect 189040 200144 580172 200172
rect 189040 200132 189046 200144
rect 580166 200132 580172 200144
rect 580224 200132 580230 200184
rect 179046 200104 179052 200116
rect 178006 200076 179052 200104
rect 178006 200048 178034 200076
rect 179046 200064 179052 200076
rect 179104 200064 179110 200116
rect 179230 200064 179236 200116
rect 179288 200104 179294 200116
rect 182910 200104 182916 200116
rect 179288 200076 182916 200104
rect 179288 200064 179294 200076
rect 182910 200064 182916 200076
rect 182968 200064 182974 200116
rect 175982 200008 177896 200036
rect 174952 199860 174958 199912
rect 175010 199860 175016 199912
rect 175504 199860 175510 199912
rect 175562 199860 175568 199912
rect 175596 199860 175602 199912
rect 175654 199860 175660 199912
rect 175688 199860 175694 199912
rect 175746 199860 175752 199912
rect 175780 199860 175786 199912
rect 175838 199860 175844 199912
rect 175522 199832 175550 199860
rect 175476 199804 175550 199832
rect 175706 199832 175734 199860
rect 175706 199804 175872 199832
rect 175476 199628 175504 199804
rect 175642 199656 175648 199708
rect 175700 199696 175706 199708
rect 175844 199696 175872 199804
rect 175700 199668 175872 199696
rect 175700 199656 175706 199668
rect 175550 199628 175556 199640
rect 175476 199600 175556 199628
rect 175550 199588 175556 199600
rect 175608 199588 175614 199640
rect 175982 199560 176010 200008
rect 177942 199996 177948 200048
rect 178000 200008 178034 200048
rect 178000 199996 178006 200008
rect 177758 199928 177764 199980
rect 177816 199968 177822 199980
rect 181898 199968 181904 199980
rect 177816 199940 181904 199968
rect 177816 199928 177822 199940
rect 181898 199928 181904 199940
rect 181956 199928 181962 199980
rect 176056 199860 176062 199912
rect 176114 199860 176120 199912
rect 176424 199860 176430 199912
rect 176482 199860 176488 199912
rect 176516 199860 176522 199912
rect 176574 199860 176580 199912
rect 176976 199860 176982 199912
rect 177034 199860 177040 199912
rect 177252 199860 177258 199912
rect 177310 199860 177316 199912
rect 177436 199860 177442 199912
rect 177494 199900 177500 199912
rect 181806 199900 181812 199912
rect 177494 199872 181812 199900
rect 177494 199860 177500 199872
rect 181806 199860 181812 199872
rect 181864 199860 181870 199912
rect 176074 199708 176102 199860
rect 176148 199792 176154 199844
rect 176206 199832 176212 199844
rect 176206 199792 176240 199832
rect 176074 199668 176108 199708
rect 176102 199656 176108 199668
rect 176160 199656 176166 199708
rect 174878 199532 176010 199560
rect 172974 199452 172980 199504
rect 173032 199464 173066 199504
rect 173032 199452 173038 199464
rect 173894 199452 173900 199504
rect 173952 199464 173986 199504
rect 173952 199452 173958 199464
rect 176102 199452 176108 199504
rect 176160 199492 176166 199504
rect 176212 199492 176240 199792
rect 176442 199696 176470 199860
rect 176160 199464 176240 199492
rect 176304 199668 176470 199696
rect 176160 199452 176166 199464
rect 174446 199424 174452 199436
rect 172900 199396 174452 199424
rect 174446 199384 174452 199396
rect 174504 199384 174510 199436
rect 172974 199356 172980 199368
rect 171520 199328 172980 199356
rect 172974 199316 172980 199328
rect 173032 199316 173038 199368
rect 174906 199288 174912 199300
rect 161722 199260 174912 199288
rect 174906 199248 174912 199260
rect 174964 199248 174970 199300
rect 176304 199288 176332 199668
rect 176534 199628 176562 199860
rect 176994 199776 177022 199860
rect 176994 199736 177028 199776
rect 177022 199724 177028 199736
rect 177080 199724 177086 199776
rect 177270 199764 177298 199860
rect 177942 199764 177948 199776
rect 177270 199736 177948 199764
rect 177942 199724 177948 199736
rect 178000 199724 178006 199776
rect 180978 199764 180984 199776
rect 180444 199736 180984 199764
rect 176838 199628 176844 199640
rect 176534 199600 176844 199628
rect 176838 199588 176844 199600
rect 176896 199588 176902 199640
rect 177298 199588 177304 199640
rect 177356 199628 177362 199640
rect 179506 199628 179512 199640
rect 177356 199600 179512 199628
rect 177356 199588 177362 199600
rect 179506 199588 179512 199600
rect 179564 199628 179570 199640
rect 180334 199628 180340 199640
rect 179564 199600 180340 199628
rect 179564 199588 179570 199600
rect 180334 199588 180340 199600
rect 180392 199588 180398 199640
rect 176654 199520 176660 199572
rect 176712 199560 176718 199572
rect 180444 199560 180472 199736
rect 180978 199724 180984 199736
rect 181036 199764 181042 199776
rect 303614 199764 303620 199776
rect 181036 199736 303620 199764
rect 181036 199724 181042 199736
rect 303614 199724 303620 199736
rect 303672 199724 303678 199776
rect 180702 199656 180708 199708
rect 180760 199696 180766 199708
rect 191098 199696 191104 199708
rect 180760 199668 191104 199696
rect 180760 199656 180766 199668
rect 191098 199656 191104 199668
rect 191156 199656 191162 199708
rect 218422 199656 218428 199708
rect 218480 199696 218486 199708
rect 402974 199696 402980 199708
rect 218480 199668 402980 199696
rect 218480 199656 218486 199668
rect 402974 199656 402980 199668
rect 403032 199656 403038 199708
rect 180518 199588 180524 199640
rect 180576 199628 180582 199640
rect 180576 199600 180840 199628
rect 180576 199588 180582 199600
rect 176712 199532 180472 199560
rect 180812 199560 180840 199600
rect 184934 199588 184940 199640
rect 184992 199628 184998 199640
rect 186222 199628 186228 199640
rect 184992 199600 186228 199628
rect 184992 199588 184998 199600
rect 186222 199588 186228 199600
rect 186280 199628 186286 199640
rect 448514 199628 448520 199640
rect 186280 199600 448520 199628
rect 186280 199588 186286 199600
rect 448514 199588 448520 199600
rect 448572 199588 448578 199640
rect 528554 199560 528560 199572
rect 180812 199532 528560 199560
rect 176712 199520 176718 199532
rect 528554 199520 528560 199532
rect 528612 199520 528618 199572
rect 176838 199452 176844 199504
rect 176896 199492 176902 199504
rect 539594 199492 539600 199504
rect 176896 199464 539600 199492
rect 176896 199452 176902 199464
rect 539594 199452 539600 199464
rect 539652 199452 539658 199504
rect 176378 199384 176384 199436
rect 176436 199384 176442 199436
rect 176470 199384 176476 199436
rect 176528 199424 176534 199436
rect 177298 199424 177304 199436
rect 176528 199396 177304 199424
rect 176528 199384 176534 199396
rect 177298 199384 177304 199396
rect 177356 199384 177362 199436
rect 177666 199384 177672 199436
rect 177724 199424 177730 199436
rect 582466 199424 582472 199436
rect 177724 199396 582472 199424
rect 177724 199384 177730 199396
rect 582466 199384 582472 199396
rect 582524 199384 582530 199436
rect 176396 199356 176424 199384
rect 179230 199356 179236 199368
rect 176396 199328 179236 199356
rect 179230 199316 179236 199328
rect 179288 199316 179294 199368
rect 176378 199288 176384 199300
rect 176304 199260 176384 199288
rect 176378 199248 176384 199260
rect 176436 199248 176442 199300
rect 192478 199288 192484 199300
rect 176626 199260 192484 199288
rect 154448 199192 158944 199220
rect 154448 199180 154454 199192
rect 160646 199180 160652 199232
rect 160704 199220 160710 199232
rect 160704 199192 169754 199220
rect 160704 199180 160710 199192
rect 161014 199112 161020 199164
rect 161072 199152 161078 199164
rect 161474 199152 161480 199164
rect 161072 199124 161480 199152
rect 161072 199112 161078 199124
rect 161474 199112 161480 199124
rect 161532 199112 161538 199164
rect 161566 199112 161572 199164
rect 161624 199152 161630 199164
rect 162118 199152 162124 199164
rect 161624 199124 162124 199152
rect 161624 199112 161630 199124
rect 162118 199112 162124 199124
rect 162176 199112 162182 199164
rect 169726 199152 169754 199192
rect 170950 199180 170956 199232
rect 171008 199220 171014 199232
rect 176626 199220 176654 199260
rect 192478 199248 192484 199260
rect 192536 199248 192542 199300
rect 171008 199192 176654 199220
rect 171008 199180 171014 199192
rect 177206 199180 177212 199232
rect 177264 199220 177270 199232
rect 185394 199220 185400 199232
rect 177264 199192 185400 199220
rect 177264 199180 177270 199192
rect 185394 199180 185400 199192
rect 185452 199180 185458 199232
rect 184934 199152 184940 199164
rect 169726 199124 184940 199152
rect 184934 199112 184940 199124
rect 184992 199112 184998 199164
rect 179690 199084 179696 199096
rect 154086 199056 179696 199084
rect 179690 199044 179696 199056
rect 179748 199084 179754 199096
rect 180702 199084 180708 199096
rect 179748 199056 180708 199084
rect 179748 199044 179754 199056
rect 180702 199044 180708 199056
rect 180760 199044 180766 199096
rect 165430 199016 165436 199028
rect 153856 198988 165436 199016
rect 165430 198976 165436 198988
rect 165488 198976 165494 199028
rect 190454 199016 190460 199028
rect 165816 198988 190460 199016
rect 156874 198948 156880 198960
rect 149394 198920 156880 198948
rect 156874 198908 156880 198920
rect 156932 198908 156938 198960
rect 156966 198908 156972 198960
rect 157024 198948 157030 198960
rect 163682 198948 163688 198960
rect 157024 198920 163688 198948
rect 157024 198908 157030 198920
rect 163682 198908 163688 198920
rect 163740 198908 163746 198960
rect 165338 198908 165344 198960
rect 165396 198948 165402 198960
rect 165816 198948 165844 198988
rect 190454 198976 190460 198988
rect 190512 198976 190518 199028
rect 165396 198920 165844 198948
rect 165396 198908 165402 198920
rect 167086 198908 167092 198960
rect 167144 198948 167150 198960
rect 188890 198948 188896 198960
rect 167144 198920 188896 198948
rect 167144 198908 167150 198920
rect 188890 198908 188896 198920
rect 188948 198948 188954 198960
rect 190086 198948 190092 198960
rect 188948 198920 190092 198948
rect 188948 198908 188954 198920
rect 190086 198908 190092 198920
rect 190144 198908 190150 198960
rect 105998 198840 106004 198892
rect 106056 198880 106062 198892
rect 120718 198880 120724 198892
rect 106056 198852 120724 198880
rect 106056 198840 106062 198852
rect 120718 198840 120724 198852
rect 120776 198840 120782 198892
rect 120994 198840 121000 198892
rect 121052 198880 121058 198892
rect 121052 198852 144914 198880
rect 121052 198840 121058 198852
rect 3510 198772 3516 198824
rect 3568 198812 3574 198824
rect 119430 198812 119436 198824
rect 3568 198784 119436 198812
rect 3568 198772 3574 198784
rect 119430 198772 119436 198784
rect 119488 198772 119494 198824
rect 120810 198772 120816 198824
rect 120868 198812 120874 198824
rect 124214 198812 124220 198824
rect 120868 198784 124220 198812
rect 120868 198772 120874 198784
rect 124214 198772 124220 198784
rect 124272 198812 124278 198824
rect 142062 198812 142068 198824
rect 124272 198784 142068 198812
rect 124272 198772 124278 198784
rect 142062 198772 142068 198784
rect 142120 198772 142126 198824
rect 117958 198704 117964 198756
rect 118016 198744 118022 198756
rect 118694 198744 118700 198756
rect 118016 198716 118700 198744
rect 118016 198704 118022 198716
rect 118694 198704 118700 198716
rect 118752 198704 118758 198756
rect 120902 198704 120908 198756
rect 120960 198744 120966 198756
rect 131298 198744 131304 198756
rect 120960 198716 131304 198744
rect 120960 198704 120966 198716
rect 131298 198704 131304 198716
rect 131356 198744 131362 198756
rect 132402 198744 132408 198756
rect 131356 198716 132408 198744
rect 131356 198704 131362 198716
rect 132402 198704 132408 198716
rect 132460 198704 132466 198756
rect 132494 198704 132500 198756
rect 132552 198744 132558 198756
rect 137002 198744 137008 198756
rect 132552 198716 137008 198744
rect 132552 198704 132558 198716
rect 137002 198704 137008 198716
rect 137060 198704 137066 198756
rect 120718 198636 120724 198688
rect 120776 198676 120782 198688
rect 133046 198676 133052 198688
rect 120776 198648 133052 198676
rect 120776 198636 120782 198648
rect 133046 198636 133052 198648
rect 133104 198636 133110 198688
rect 126882 198568 126888 198620
rect 126940 198608 126946 198620
rect 130930 198608 130936 198620
rect 126940 198580 130936 198608
rect 126940 198568 126946 198580
rect 130930 198568 130936 198580
rect 130988 198568 130994 198620
rect 144886 198608 144914 198852
rect 151262 198840 151268 198892
rect 151320 198880 151326 198892
rect 154574 198880 154580 198892
rect 151320 198852 154580 198880
rect 151320 198840 151326 198852
rect 154574 198840 154580 198852
rect 154632 198840 154638 198892
rect 160922 198840 160928 198892
rect 160980 198880 160986 198892
rect 166534 198880 166540 198892
rect 160980 198852 166540 198880
rect 160980 198840 160986 198852
rect 166534 198840 166540 198852
rect 166592 198840 166598 198892
rect 167914 198840 167920 198892
rect 167972 198880 167978 198892
rect 194502 198880 194508 198892
rect 167972 198852 194508 198880
rect 167972 198840 167978 198852
rect 194502 198840 194508 198852
rect 194560 198840 194566 198892
rect 146386 198772 146392 198824
rect 146444 198812 146450 198824
rect 146846 198812 146852 198824
rect 146444 198784 146852 198812
rect 146444 198772 146450 198784
rect 146846 198772 146852 198784
rect 146904 198772 146910 198824
rect 149422 198772 149428 198824
rect 149480 198812 149486 198824
rect 161842 198812 161848 198824
rect 149480 198784 161848 198812
rect 149480 198772 149486 198784
rect 161842 198772 161848 198784
rect 161900 198812 161906 198824
rect 165338 198812 165344 198824
rect 161900 198784 165344 198812
rect 161900 198772 161906 198784
rect 165338 198772 165344 198784
rect 165396 198772 165402 198824
rect 165430 198772 165436 198824
rect 165488 198812 165494 198824
rect 170950 198812 170956 198824
rect 165488 198784 170956 198812
rect 165488 198772 165494 198784
rect 170950 198772 170956 198784
rect 171008 198772 171014 198824
rect 171042 198772 171048 198824
rect 171100 198812 171106 198824
rect 218054 198812 218060 198824
rect 171100 198784 218060 198812
rect 171100 198772 171106 198784
rect 218054 198772 218060 198784
rect 218112 198812 218118 198824
rect 218422 198812 218428 198824
rect 218112 198784 218428 198812
rect 218112 198772 218118 198784
rect 218422 198772 218428 198784
rect 218480 198772 218486 198824
rect 147674 198704 147680 198756
rect 147732 198744 147738 198756
rect 153102 198744 153108 198756
rect 147732 198716 153108 198744
rect 147732 198704 147738 198716
rect 153102 198704 153108 198716
rect 153160 198704 153166 198756
rect 153838 198704 153844 198756
rect 153896 198744 153902 198756
rect 154022 198744 154028 198756
rect 153896 198716 154028 198744
rect 153896 198704 153902 198716
rect 154022 198704 154028 198716
rect 154080 198704 154086 198756
rect 157794 198704 157800 198756
rect 157852 198744 157858 198756
rect 158438 198744 158444 198756
rect 157852 198716 158444 198744
rect 157852 198704 157858 198716
rect 158438 198704 158444 198716
rect 158496 198704 158502 198756
rect 176470 198744 176476 198756
rect 168346 198716 176476 198744
rect 148962 198636 148968 198688
rect 149020 198676 149026 198688
rect 154390 198676 154396 198688
rect 149020 198648 154396 198676
rect 149020 198636 149026 198648
rect 154390 198636 154396 198648
rect 154448 198636 154454 198688
rect 160738 198636 160744 198688
rect 160796 198676 160802 198688
rect 165614 198676 165620 198688
rect 160796 198648 165620 198676
rect 160796 198636 160802 198648
rect 165614 198636 165620 198648
rect 165672 198636 165678 198688
rect 149422 198608 149428 198620
rect 144886 198580 149428 198608
rect 149422 198568 149428 198580
rect 149480 198568 149486 198620
rect 149882 198568 149888 198620
rect 149940 198608 149946 198620
rect 168346 198608 168374 198716
rect 176470 198704 176476 198716
rect 176528 198704 176534 198756
rect 176930 198704 176936 198756
rect 176988 198744 176994 198756
rect 177114 198744 177120 198756
rect 176988 198716 177120 198744
rect 176988 198704 176994 198716
rect 177114 198704 177120 198716
rect 177172 198704 177178 198756
rect 182910 198704 182916 198756
rect 182968 198744 182974 198756
rect 185578 198744 185584 198756
rect 182968 198716 185584 198744
rect 182968 198704 182974 198716
rect 185578 198704 185584 198716
rect 185636 198744 185642 198756
rect 189718 198744 189724 198756
rect 185636 198716 189724 198744
rect 185636 198704 185642 198716
rect 189718 198704 189724 198716
rect 189776 198704 189782 198756
rect 168466 198636 168472 198688
rect 168524 198676 168530 198688
rect 168742 198676 168748 198688
rect 168524 198648 168748 198676
rect 168524 198636 168530 198648
rect 168742 198636 168748 198648
rect 168800 198636 168806 198688
rect 169294 198636 169300 198688
rect 169352 198676 169358 198688
rect 194594 198676 194600 198688
rect 169352 198648 194600 198676
rect 169352 198636 169358 198648
rect 194594 198636 194600 198648
rect 194652 198636 194658 198688
rect 149940 198580 168374 198608
rect 149940 198568 149946 198580
rect 172514 198568 172520 198620
rect 172572 198608 172578 198620
rect 177482 198608 177488 198620
rect 172572 198580 177488 198608
rect 172572 198568 172578 198580
rect 177482 198568 177488 198580
rect 177540 198568 177546 198620
rect 190822 198608 190828 198620
rect 180904 198580 190828 198608
rect 129182 198500 129188 198552
rect 129240 198540 129246 198552
rect 140958 198540 140964 198552
rect 129240 198512 140964 198540
rect 129240 198500 129246 198512
rect 140958 198500 140964 198512
rect 141016 198500 141022 198552
rect 142246 198500 142252 198552
rect 142304 198540 142310 198552
rect 147030 198540 147036 198552
rect 142304 198512 147036 198540
rect 142304 198500 142310 198512
rect 147030 198500 147036 198512
rect 147088 198500 147094 198552
rect 151446 198500 151452 198552
rect 151504 198540 151510 198552
rect 151504 198512 170628 198540
rect 151504 198500 151510 198512
rect 125502 198432 125508 198484
rect 125560 198472 125566 198484
rect 138014 198472 138020 198484
rect 125560 198444 138020 198472
rect 125560 198432 125566 198444
rect 138014 198432 138020 198444
rect 138072 198432 138078 198484
rect 153010 198432 153016 198484
rect 153068 198472 153074 198484
rect 161014 198472 161020 198484
rect 153068 198444 161020 198472
rect 153068 198432 153074 198444
rect 161014 198432 161020 198444
rect 161072 198432 161078 198484
rect 163222 198432 163228 198484
rect 163280 198472 163286 198484
rect 163280 198444 167914 198472
rect 163280 198432 163286 198444
rect 128170 198364 128176 198416
rect 128228 198404 128234 198416
rect 141234 198404 141240 198416
rect 128228 198376 141240 198404
rect 128228 198364 128234 198376
rect 141234 198364 141240 198376
rect 141292 198364 141298 198416
rect 151078 198364 151084 198416
rect 151136 198404 151142 198416
rect 154850 198404 154856 198416
rect 151136 198376 154856 198404
rect 151136 198364 151142 198376
rect 154850 198364 154856 198376
rect 154908 198364 154914 198416
rect 159818 198364 159824 198416
rect 159876 198404 159882 198416
rect 166534 198404 166540 198416
rect 159876 198376 166540 198404
rect 159876 198364 159882 198376
rect 166534 198364 166540 198376
rect 166592 198364 166598 198416
rect 166902 198364 166908 198416
rect 166960 198404 166966 198416
rect 167730 198404 167736 198416
rect 166960 198376 167736 198404
rect 166960 198364 166966 198376
rect 167730 198364 167736 198376
rect 167788 198364 167794 198416
rect 167886 198404 167914 198444
rect 169754 198432 169760 198484
rect 169812 198472 169818 198484
rect 170030 198472 170036 198484
rect 169812 198444 170036 198472
rect 169812 198432 169818 198444
rect 170030 198432 170036 198444
rect 170088 198432 170094 198484
rect 170600 198472 170628 198512
rect 170674 198500 170680 198552
rect 170732 198540 170738 198552
rect 171686 198540 171692 198552
rect 170732 198512 171692 198540
rect 170732 198500 170738 198512
rect 171686 198500 171692 198512
rect 171744 198500 171750 198552
rect 171962 198500 171968 198552
rect 172020 198540 172026 198552
rect 180904 198540 180932 198580
rect 190822 198568 190828 198580
rect 190880 198608 190886 198620
rect 191742 198608 191748 198620
rect 190880 198580 191748 198608
rect 190880 198568 190886 198580
rect 191742 198568 191748 198580
rect 191800 198568 191806 198620
rect 172020 198512 180932 198540
rect 172020 198500 172026 198512
rect 185394 198500 185400 198552
rect 185452 198540 185458 198552
rect 191374 198540 191380 198552
rect 185452 198512 191380 198540
rect 185452 198500 185458 198512
rect 191374 198500 191380 198512
rect 191432 198500 191438 198552
rect 172422 198472 172428 198484
rect 170600 198444 172428 198472
rect 172422 198432 172428 198444
rect 172480 198432 172486 198484
rect 172790 198432 172796 198484
rect 172848 198472 172854 198484
rect 173066 198472 173072 198484
rect 172848 198444 173072 198472
rect 172848 198432 172854 198444
rect 173066 198432 173072 198444
rect 173124 198432 173130 198484
rect 175550 198432 175556 198484
rect 175608 198472 175614 198484
rect 175918 198472 175924 198484
rect 175608 198444 175924 198472
rect 175608 198432 175614 198444
rect 175918 198432 175924 198444
rect 175976 198432 175982 198484
rect 176010 198432 176016 198484
rect 176068 198472 176074 198484
rect 176654 198472 176660 198484
rect 176068 198444 176660 198472
rect 176068 198432 176074 198444
rect 176654 198432 176660 198444
rect 176712 198432 176718 198484
rect 176746 198432 176752 198484
rect 176804 198472 176810 198484
rect 189534 198472 189540 198484
rect 176804 198444 189540 198472
rect 176804 198432 176810 198444
rect 189534 198432 189540 198444
rect 189592 198432 189598 198484
rect 167886 198376 176746 198404
rect 129642 198296 129648 198348
rect 129700 198336 129706 198348
rect 140866 198336 140872 198348
rect 129700 198308 140872 198336
rect 129700 198296 129706 198308
rect 140866 198296 140872 198308
rect 140924 198296 140930 198348
rect 142890 198296 142896 198348
rect 142948 198336 142954 198348
rect 143902 198336 143908 198348
rect 142948 198308 143908 198336
rect 142948 198296 142954 198308
rect 143902 198296 143908 198308
rect 143960 198296 143966 198348
rect 163866 198296 163872 198348
rect 163924 198336 163930 198348
rect 165614 198336 165620 198348
rect 163924 198308 165620 198336
rect 163924 198296 163930 198308
rect 165614 198296 165620 198308
rect 165672 198296 165678 198348
rect 166718 198296 166724 198348
rect 166776 198336 166782 198348
rect 172514 198336 172520 198348
rect 166776 198308 172520 198336
rect 166776 198296 166782 198308
rect 172514 198296 172520 198308
rect 172572 198296 172578 198348
rect 176010 198336 176016 198348
rect 172624 198308 176016 198336
rect 126514 198228 126520 198280
rect 126572 198268 126578 198280
rect 134150 198268 134156 198280
rect 126572 198240 134156 198268
rect 126572 198228 126578 198240
rect 134150 198228 134156 198240
rect 134208 198228 134214 198280
rect 137094 198228 137100 198280
rect 137152 198268 137158 198280
rect 137646 198268 137652 198280
rect 137152 198240 137652 198268
rect 137152 198228 137158 198240
rect 137646 198228 137652 198240
rect 137704 198228 137710 198280
rect 140958 198228 140964 198280
rect 141016 198268 141022 198280
rect 141878 198268 141884 198280
rect 141016 198240 141884 198268
rect 141016 198228 141022 198240
rect 141878 198228 141884 198240
rect 141936 198228 141942 198280
rect 158162 198228 158168 198280
rect 158220 198268 158226 198280
rect 159450 198268 159456 198280
rect 158220 198240 159456 198268
rect 158220 198228 158226 198240
rect 159450 198228 159456 198240
rect 159508 198228 159514 198280
rect 168558 198228 168564 198280
rect 168616 198268 168622 198280
rect 171778 198268 171784 198280
rect 168616 198240 171784 198268
rect 168616 198228 168622 198240
rect 171778 198228 171784 198240
rect 171836 198228 171842 198280
rect 172422 198228 172428 198280
rect 172480 198268 172486 198280
rect 172624 198268 172652 198308
rect 176010 198296 176016 198308
rect 176068 198296 176074 198348
rect 176718 198336 176746 198376
rect 177390 198336 177396 198348
rect 176718 198308 177396 198336
rect 177390 198296 177396 198308
rect 177448 198296 177454 198348
rect 172480 198240 172652 198268
rect 172480 198228 172486 198240
rect 173066 198228 173072 198280
rect 173124 198268 173130 198280
rect 177758 198268 177764 198280
rect 173124 198240 177764 198268
rect 173124 198228 173130 198240
rect 177758 198228 177764 198240
rect 177816 198228 177822 198280
rect 193214 198228 193220 198280
rect 193272 198268 193278 198280
rect 204346 198268 204352 198280
rect 193272 198240 204352 198268
rect 193272 198228 193278 198240
rect 204346 198228 204352 198240
rect 204404 198228 204410 198280
rect 100662 198160 100668 198212
rect 100720 198200 100726 198212
rect 129734 198200 129740 198212
rect 100720 198172 129740 198200
rect 100720 198160 100726 198172
rect 129734 198160 129740 198172
rect 129792 198160 129798 198212
rect 137278 198160 137284 198212
rect 137336 198200 137342 198212
rect 139670 198200 139676 198212
rect 137336 198172 139676 198200
rect 137336 198160 137342 198172
rect 139670 198160 139676 198172
rect 139728 198160 139734 198212
rect 140038 198160 140044 198212
rect 140096 198200 140102 198212
rect 140314 198200 140320 198212
rect 140096 198172 140320 198200
rect 140096 198160 140102 198172
rect 140314 198160 140320 198172
rect 140372 198160 140378 198212
rect 142338 198160 142344 198212
rect 142396 198200 142402 198212
rect 143442 198200 143448 198212
rect 142396 198172 143448 198200
rect 142396 198160 142402 198172
rect 143442 198160 143448 198172
rect 143500 198160 143506 198212
rect 159818 198160 159824 198212
rect 159876 198200 159882 198212
rect 160922 198200 160928 198212
rect 159876 198172 160928 198200
rect 159876 198160 159882 198172
rect 160922 198160 160928 198172
rect 160980 198160 160986 198212
rect 161290 198160 161296 198212
rect 161348 198200 161354 198212
rect 163682 198200 163688 198212
rect 161348 198172 163688 198200
rect 161348 198160 161354 198172
rect 163682 198160 163688 198172
rect 163740 198160 163746 198212
rect 166902 198160 166908 198212
rect 166960 198200 166966 198212
rect 180794 198200 180800 198212
rect 166960 198172 180800 198200
rect 166960 198160 166966 198172
rect 180794 198160 180800 198172
rect 180852 198160 180858 198212
rect 181070 198160 181076 198212
rect 181128 198200 181134 198212
rect 196066 198200 196072 198212
rect 181128 198172 196072 198200
rect 181128 198160 181134 198172
rect 196066 198160 196072 198172
rect 196124 198200 196130 198212
rect 201586 198200 201592 198212
rect 196124 198172 201592 198200
rect 196124 198160 196130 198172
rect 201586 198160 201592 198172
rect 201644 198160 201650 198212
rect 114462 198092 114468 198144
rect 114520 198132 114526 198144
rect 128446 198132 128452 198144
rect 114520 198104 128452 198132
rect 114520 198092 114526 198104
rect 128446 198092 128452 198104
rect 128504 198132 128510 198144
rect 129642 198132 129648 198144
rect 128504 198104 129648 198132
rect 128504 198092 128510 198104
rect 129642 198092 129648 198104
rect 129700 198092 129706 198144
rect 141878 198092 141884 198144
rect 141936 198132 141942 198144
rect 150802 198132 150808 198144
rect 141936 198104 150808 198132
rect 141936 198092 141942 198104
rect 150802 198092 150808 198104
rect 150860 198092 150866 198144
rect 159450 198092 159456 198144
rect 159508 198132 159514 198144
rect 159726 198132 159732 198144
rect 159508 198104 159732 198132
rect 159508 198092 159514 198104
rect 159726 198092 159732 198104
rect 159784 198092 159790 198144
rect 164694 198092 164700 198144
rect 164752 198132 164758 198144
rect 184934 198132 184940 198144
rect 164752 198104 184940 198132
rect 164752 198092 164758 198104
rect 184934 198092 184940 198104
rect 184992 198092 184998 198144
rect 194594 198092 194600 198144
rect 194652 198132 194658 198144
rect 212534 198132 212540 198144
rect 194652 198104 212540 198132
rect 194652 198092 194658 198104
rect 212534 198092 212540 198104
rect 212592 198092 212598 198144
rect 100570 198024 100576 198076
rect 100628 198064 100634 198076
rect 131942 198064 131948 198076
rect 100628 198036 131948 198064
rect 100628 198024 100634 198036
rect 131942 198024 131948 198036
rect 132000 198024 132006 198076
rect 132954 198024 132960 198076
rect 133012 198064 133018 198076
rect 133230 198064 133236 198076
rect 133012 198036 133236 198064
rect 133012 198024 133018 198036
rect 133230 198024 133236 198036
rect 133288 198024 133294 198076
rect 139854 198064 139860 198076
rect 137986 198036 139860 198064
rect 62758 197956 62764 198008
rect 62816 197996 62822 198008
rect 99190 197996 99196 198008
rect 62816 197968 99196 197996
rect 62816 197956 62822 197968
rect 99190 197956 99196 197968
rect 99248 197996 99254 198008
rect 133506 197996 133512 198008
rect 99248 197968 133512 197996
rect 99248 197956 99254 197968
rect 133506 197956 133512 197968
rect 133564 197956 133570 198008
rect 137986 197996 138014 198036
rect 139854 198024 139860 198036
rect 139912 198024 139918 198076
rect 140682 198024 140688 198076
rect 140740 198064 140746 198076
rect 141694 198064 141700 198076
rect 140740 198036 141700 198064
rect 140740 198024 140746 198036
rect 141694 198024 141700 198036
rect 141752 198024 141758 198076
rect 144730 198024 144736 198076
rect 144788 198064 144794 198076
rect 145006 198064 145012 198076
rect 144788 198036 145012 198064
rect 144788 198024 144794 198036
rect 145006 198024 145012 198036
rect 145064 198024 145070 198076
rect 156874 198024 156880 198076
rect 156932 198064 156938 198076
rect 180150 198064 180156 198076
rect 156932 198036 180156 198064
rect 156932 198024 156938 198036
rect 180150 198024 180156 198036
rect 180208 198024 180214 198076
rect 191742 198024 191748 198076
rect 191800 198064 191806 198076
rect 211430 198064 211436 198076
rect 191800 198036 211436 198064
rect 191800 198024 191806 198036
rect 211430 198024 211436 198036
rect 211488 198024 211494 198076
rect 137526 197968 138014 197996
rect 127986 197888 127992 197940
rect 128044 197928 128050 197940
rect 131758 197928 131764 197940
rect 128044 197900 131764 197928
rect 128044 197888 128050 197900
rect 131758 197888 131764 197900
rect 131816 197888 131822 197940
rect 135346 197928 135352 197940
rect 131868 197900 135352 197928
rect 127802 197820 127808 197872
rect 127860 197860 127866 197872
rect 131868 197860 131896 197900
rect 135346 197888 135352 197900
rect 135404 197888 135410 197940
rect 137526 197860 137554 197968
rect 138382 197956 138388 198008
rect 138440 197996 138446 198008
rect 139302 197996 139308 198008
rect 138440 197968 139308 197996
rect 138440 197956 138446 197968
rect 139302 197956 139308 197968
rect 139360 197956 139366 198008
rect 139946 197956 139952 198008
rect 140004 197996 140010 198008
rect 141050 197996 141056 198008
rect 140004 197968 141056 197996
rect 140004 197956 140010 197968
rect 141050 197956 141056 197968
rect 141108 197956 141114 198008
rect 142062 197956 142068 198008
rect 142120 197996 142126 198008
rect 142120 197968 142844 197996
rect 142120 197956 142126 197968
rect 139762 197888 139768 197940
rect 139820 197928 139826 197940
rect 140774 197928 140780 197940
rect 139820 197900 140780 197928
rect 139820 197888 139826 197900
rect 140774 197888 140780 197900
rect 140832 197888 140838 197940
rect 127860 197832 131896 197860
rect 133156 197832 137554 197860
rect 127860 197820 127866 197832
rect 125686 197616 125692 197668
rect 125744 197656 125750 197668
rect 133156 197656 133184 197832
rect 139578 197820 139584 197872
rect 139636 197860 139642 197872
rect 139946 197860 139952 197872
rect 139636 197832 139952 197860
rect 139636 197820 139642 197832
rect 139946 197820 139952 197832
rect 140004 197820 140010 197872
rect 140314 197820 140320 197872
rect 140372 197860 140378 197872
rect 142816 197860 142844 197968
rect 154850 197956 154856 198008
rect 154908 197996 154914 198008
rect 165062 197996 165068 198008
rect 154908 197968 165068 197996
rect 154908 197956 154914 197968
rect 165062 197956 165068 197968
rect 165120 197956 165126 198008
rect 166902 197996 166908 198008
rect 166184 197968 166908 197996
rect 144270 197888 144276 197940
rect 144328 197928 144334 197940
rect 145282 197928 145288 197940
rect 144328 197900 145288 197928
rect 144328 197888 144334 197900
rect 145282 197888 145288 197900
rect 145340 197888 145346 197940
rect 150710 197888 150716 197940
rect 150768 197928 150774 197940
rect 151630 197928 151636 197940
rect 150768 197900 151636 197928
rect 150768 197888 150774 197900
rect 151630 197888 151636 197900
rect 151688 197888 151694 197940
rect 146110 197860 146116 197872
rect 140372 197832 142568 197860
rect 142816 197832 146116 197860
rect 140372 197820 140378 197832
rect 125744 197628 133184 197656
rect 133248 197764 133874 197792
rect 125744 197616 125750 197628
rect 132126 197548 132132 197600
rect 132184 197588 132190 197600
rect 133248 197588 133276 197764
rect 133846 197656 133874 197764
rect 140774 197752 140780 197804
rect 140832 197792 140838 197804
rect 141142 197792 141148 197804
rect 140832 197764 141148 197792
rect 140832 197752 140838 197764
rect 141142 197752 141148 197764
rect 141200 197752 141206 197804
rect 141510 197752 141516 197804
rect 141568 197792 141574 197804
rect 142062 197792 142068 197804
rect 141568 197764 142068 197792
rect 141568 197752 141574 197764
rect 142062 197752 142068 197764
rect 142120 197752 142126 197804
rect 142540 197792 142568 197832
rect 146110 197820 146116 197832
rect 146168 197820 146174 197872
rect 161474 197820 161480 197872
rect 161532 197860 161538 197872
rect 166184 197860 166212 197968
rect 166902 197956 166908 197968
rect 166960 197956 166966 198008
rect 168650 197956 168656 198008
rect 168708 197996 168714 198008
rect 168708 197968 173894 197996
rect 168708 197956 168714 197968
rect 167086 197888 167092 197940
rect 167144 197928 167150 197940
rect 169754 197928 169760 197940
rect 167144 197900 169760 197928
rect 167144 197888 167150 197900
rect 169754 197888 169760 197900
rect 169812 197888 169818 197940
rect 173158 197888 173164 197940
rect 173216 197928 173222 197940
rect 173342 197928 173348 197940
rect 173216 197900 173348 197928
rect 173216 197888 173222 197900
rect 173342 197888 173348 197900
rect 173400 197888 173406 197940
rect 173866 197928 173894 197968
rect 174538 197956 174544 198008
rect 174596 197996 174602 198008
rect 174814 197996 174820 198008
rect 174596 197968 174820 197996
rect 174596 197956 174602 197968
rect 174814 197956 174820 197968
rect 174872 197956 174878 198008
rect 177942 197956 177948 198008
rect 178000 197996 178006 198008
rect 178218 197996 178224 198008
rect 178000 197968 178224 197996
rect 178000 197956 178006 197968
rect 178218 197956 178224 197968
rect 178276 197956 178282 198008
rect 180702 197956 180708 198008
rect 180760 197996 180766 198008
rect 582558 197996 582564 198008
rect 180760 197968 582564 197996
rect 180760 197956 180766 197968
rect 582558 197956 582564 197968
rect 582616 197956 582622 198008
rect 182174 197928 182180 197940
rect 173866 197900 182180 197928
rect 182174 197888 182180 197900
rect 182232 197888 182238 197940
rect 161532 197832 166212 197860
rect 161532 197820 161538 197832
rect 166534 197820 166540 197872
rect 166592 197860 166598 197872
rect 168190 197860 168196 197872
rect 166592 197832 168196 197860
rect 166592 197820 166598 197832
rect 168190 197820 168196 197832
rect 168248 197820 168254 197872
rect 172698 197820 172704 197872
rect 172756 197860 172762 197872
rect 177574 197860 177580 197872
rect 172756 197832 177580 197860
rect 172756 197820 172762 197832
rect 177574 197820 177580 197832
rect 177632 197820 177638 197872
rect 177850 197820 177856 197872
rect 177908 197860 177914 197872
rect 186406 197860 186412 197872
rect 177908 197832 186412 197860
rect 177908 197820 177914 197832
rect 186406 197820 186412 197832
rect 186464 197820 186470 197872
rect 145282 197792 145288 197804
rect 142540 197764 145288 197792
rect 145282 197752 145288 197764
rect 145340 197752 145346 197804
rect 158254 197752 158260 197804
rect 158312 197792 158318 197804
rect 166718 197792 166724 197804
rect 158312 197764 166724 197792
rect 158312 197752 158318 197764
rect 166718 197752 166724 197764
rect 166776 197752 166782 197804
rect 172514 197752 172520 197804
rect 172572 197792 172578 197804
rect 174538 197792 174544 197804
rect 172572 197764 174544 197792
rect 172572 197752 172578 197764
rect 174538 197752 174544 197764
rect 174596 197752 174602 197804
rect 177666 197752 177672 197804
rect 177724 197792 177730 197804
rect 186314 197792 186320 197804
rect 177724 197764 186320 197792
rect 177724 197752 177730 197764
rect 186314 197752 186320 197764
rect 186372 197752 186378 197804
rect 136726 197684 136732 197736
rect 136784 197724 136790 197736
rect 148226 197724 148232 197736
rect 136784 197696 148232 197724
rect 136784 197684 136790 197696
rect 148226 197684 148232 197696
rect 148284 197684 148290 197736
rect 159358 197684 159364 197736
rect 159416 197724 159422 197736
rect 165890 197724 165896 197736
rect 159416 197696 165896 197724
rect 159416 197684 159422 197696
rect 165890 197684 165896 197696
rect 165948 197684 165954 197736
rect 171778 197684 171784 197736
rect 171836 197724 171842 197736
rect 182082 197724 182088 197736
rect 171836 197696 182088 197724
rect 171836 197684 171842 197696
rect 182082 197684 182088 197696
rect 182140 197684 182146 197736
rect 140038 197656 140044 197668
rect 133846 197628 140044 197656
rect 140038 197616 140044 197628
rect 140096 197616 140102 197668
rect 140682 197616 140688 197668
rect 140740 197656 140746 197668
rect 142246 197656 142252 197668
rect 140740 197628 142252 197656
rect 140740 197616 140746 197628
rect 142246 197616 142252 197628
rect 142304 197616 142310 197668
rect 145006 197616 145012 197668
rect 145064 197656 145070 197668
rect 146386 197656 146392 197668
rect 145064 197628 146392 197656
rect 145064 197616 145070 197628
rect 146386 197616 146392 197628
rect 146444 197616 146450 197668
rect 165614 197616 165620 197668
rect 165672 197656 165678 197668
rect 177758 197656 177764 197668
rect 165672 197628 177764 197656
rect 165672 197616 165678 197628
rect 177758 197616 177764 197628
rect 177816 197616 177822 197668
rect 132184 197560 133276 197588
rect 132184 197548 132190 197560
rect 137094 197548 137100 197600
rect 137152 197588 137158 197600
rect 173066 197588 173072 197600
rect 137152 197560 173072 197588
rect 137152 197548 137158 197560
rect 173066 197548 173072 197560
rect 173124 197548 173130 197600
rect 174722 197548 174728 197600
rect 174780 197588 174786 197600
rect 174906 197588 174912 197600
rect 174780 197560 174912 197588
rect 174780 197548 174786 197560
rect 174906 197548 174912 197560
rect 174964 197548 174970 197600
rect 175274 197548 175280 197600
rect 175332 197588 175338 197600
rect 182634 197588 182640 197600
rect 175332 197560 182640 197588
rect 175332 197548 175338 197560
rect 182634 197548 182640 197560
rect 182692 197548 182698 197600
rect 126606 197480 126612 197532
rect 126664 197520 126670 197532
rect 137278 197520 137284 197532
rect 126664 197492 137284 197520
rect 126664 197480 126670 197492
rect 137278 197480 137284 197492
rect 137336 197480 137342 197532
rect 146570 197520 146576 197532
rect 142264 197492 146576 197520
rect 95694 197412 95700 197464
rect 95752 197452 95758 197464
rect 109126 197452 109132 197464
rect 95752 197424 109132 197452
rect 95752 197412 95758 197424
rect 109126 197412 109132 197424
rect 109184 197412 109190 197464
rect 119982 197412 119988 197464
rect 120040 197452 120046 197464
rect 125594 197452 125600 197464
rect 120040 197424 125600 197452
rect 120040 197412 120046 197424
rect 125594 197412 125600 197424
rect 125652 197452 125658 197464
rect 126882 197452 126888 197464
rect 125652 197424 126888 197452
rect 125652 197412 125658 197424
rect 126882 197412 126888 197424
rect 126940 197412 126946 197464
rect 94682 197344 94688 197396
rect 94740 197384 94746 197396
rect 99282 197384 99288 197396
rect 94740 197356 99288 197384
rect 94740 197344 94746 197356
rect 99282 197344 99288 197356
rect 99340 197384 99346 197396
rect 128354 197384 128360 197396
rect 99340 197356 128360 197384
rect 99340 197344 99346 197356
rect 128354 197344 128360 197356
rect 128412 197344 128418 197396
rect 133138 197344 133144 197396
rect 133196 197384 133202 197396
rect 133874 197384 133880 197396
rect 133196 197356 133880 197384
rect 133196 197344 133202 197356
rect 133874 197344 133880 197356
rect 133932 197384 133938 197396
rect 137094 197384 137100 197396
rect 133932 197356 137100 197384
rect 133932 197344 133938 197356
rect 137094 197344 137100 197356
rect 137152 197344 137158 197396
rect 139486 197344 139492 197396
rect 139544 197384 139550 197396
rect 140314 197384 140320 197396
rect 139544 197356 140320 197384
rect 139544 197344 139550 197356
rect 140314 197344 140320 197356
rect 140372 197344 140378 197396
rect 142264 197384 142292 197492
rect 146570 197480 146576 197492
rect 146628 197480 146634 197532
rect 155034 197480 155040 197532
rect 155092 197520 155098 197532
rect 155092 197492 163820 197520
rect 155092 197480 155098 197492
rect 144178 197412 144184 197464
rect 144236 197452 144242 197464
rect 144638 197452 144644 197464
rect 144236 197424 144644 197452
rect 144236 197412 144242 197424
rect 144638 197412 144644 197424
rect 144696 197412 144702 197464
rect 146386 197412 146392 197464
rect 146444 197452 146450 197464
rect 147674 197452 147680 197464
rect 146444 197424 147680 197452
rect 146444 197412 146450 197424
rect 147674 197412 147680 197424
rect 147732 197412 147738 197464
rect 140424 197356 142292 197384
rect 133966 197276 133972 197328
rect 134024 197316 134030 197328
rect 134334 197316 134340 197328
rect 134024 197288 134340 197316
rect 134024 197276 134030 197288
rect 134334 197276 134340 197288
rect 134392 197276 134398 197328
rect 139302 197276 139308 197328
rect 139360 197316 139366 197328
rect 140424 197316 140452 197356
rect 142982 197344 142988 197396
rect 143040 197384 143046 197396
rect 145190 197384 145196 197396
rect 143040 197356 145196 197384
rect 143040 197344 143046 197356
rect 145190 197344 145196 197356
rect 145248 197344 145254 197396
rect 139360 197288 140452 197316
rect 139360 197276 139366 197288
rect 141510 197276 141516 197328
rect 141568 197316 141574 197328
rect 144822 197316 144828 197328
rect 141568 197288 144828 197316
rect 141568 197276 141574 197288
rect 144822 197276 144828 197288
rect 144880 197276 144886 197328
rect 108574 197208 108580 197260
rect 108632 197248 108638 197260
rect 156598 197248 156604 197260
rect 108632 197220 156604 197248
rect 108632 197208 108638 197220
rect 156598 197208 156604 197220
rect 156656 197248 156662 197260
rect 156874 197248 156880 197260
rect 156656 197220 156880 197248
rect 156656 197208 156662 197220
rect 156874 197208 156880 197220
rect 156932 197208 156938 197260
rect 163792 197192 163820 197492
rect 168190 197480 168196 197532
rect 168248 197520 168254 197532
rect 168834 197520 168840 197532
rect 168248 197492 168840 197520
rect 168248 197480 168254 197492
rect 168834 197480 168840 197492
rect 168892 197480 168898 197532
rect 164234 197412 164240 197464
rect 164292 197452 164298 197464
rect 172054 197452 172060 197464
rect 164292 197424 172060 197452
rect 164292 197412 164298 197424
rect 172054 197412 172060 197424
rect 172112 197412 172118 197464
rect 165338 197344 165344 197396
rect 165396 197384 165402 197396
rect 173434 197384 173440 197396
rect 165396 197356 173440 197384
rect 165396 197344 165402 197356
rect 173434 197344 173440 197356
rect 173492 197344 173498 197396
rect 165062 197276 165068 197328
rect 165120 197316 165126 197328
rect 167086 197316 167092 197328
rect 165120 197288 167092 197316
rect 165120 197276 165126 197288
rect 167086 197276 167092 197288
rect 167144 197276 167150 197328
rect 169938 197276 169944 197328
rect 169996 197316 170002 197328
rect 170674 197316 170680 197328
rect 169996 197288 170680 197316
rect 169996 197276 170002 197288
rect 170674 197276 170680 197288
rect 170732 197316 170738 197328
rect 175182 197316 175188 197328
rect 170732 197288 175188 197316
rect 170732 197276 170738 197288
rect 175182 197276 175188 197288
rect 175240 197276 175246 197328
rect 175458 197276 175464 197328
rect 175516 197316 175522 197328
rect 189074 197316 189080 197328
rect 175516 197288 189080 197316
rect 175516 197276 175522 197288
rect 189074 197276 189080 197288
rect 189132 197276 189138 197328
rect 167270 197208 167276 197260
rect 167328 197248 167334 197260
rect 175918 197248 175924 197260
rect 167328 197220 175924 197248
rect 167328 197208 167334 197220
rect 175918 197208 175924 197220
rect 175976 197208 175982 197260
rect 176562 197208 176568 197260
rect 176620 197248 176626 197260
rect 185670 197248 185676 197260
rect 176620 197220 185676 197248
rect 176620 197208 176626 197220
rect 185670 197208 185676 197220
rect 185728 197208 185734 197260
rect 111058 197140 111064 197192
rect 111116 197180 111122 197192
rect 158162 197180 158168 197192
rect 111116 197152 158168 197180
rect 111116 197140 111122 197152
rect 158162 197140 158168 197152
rect 158220 197140 158226 197192
rect 163774 197140 163780 197192
rect 163832 197140 163838 197192
rect 186498 197180 186504 197192
rect 163976 197152 186504 197180
rect 109126 197072 109132 197124
rect 109184 197112 109190 197124
rect 144270 197112 144276 197124
rect 109184 197084 144276 197112
rect 109184 197072 109190 197084
rect 144270 197072 144276 197084
rect 144328 197072 144334 197124
rect 146202 197072 146208 197124
rect 146260 197112 146266 197124
rect 149054 197112 149060 197124
rect 146260 197084 149060 197112
rect 146260 197072 146266 197084
rect 149054 197072 149060 197084
rect 149112 197072 149118 197124
rect 130654 197004 130660 197056
rect 130712 197044 130718 197056
rect 141878 197044 141884 197056
rect 130712 197016 141884 197044
rect 130712 197004 130718 197016
rect 141878 197004 141884 197016
rect 141936 197004 141942 197056
rect 145650 197044 145656 197056
rect 142724 197016 145656 197044
rect 133966 196936 133972 196988
rect 134024 196976 134030 196988
rect 142724 196976 142752 197016
rect 145650 197004 145656 197016
rect 145708 197004 145714 197056
rect 159082 197004 159088 197056
rect 159140 197044 159146 197056
rect 163976 197044 164004 197152
rect 186498 197140 186504 197152
rect 186556 197140 186562 197192
rect 164878 197072 164884 197124
rect 164936 197112 164942 197124
rect 192478 197112 192484 197124
rect 164936 197084 192484 197112
rect 164936 197072 164942 197084
rect 192478 197072 192484 197084
rect 192536 197072 192542 197124
rect 159140 197016 164004 197044
rect 159140 197004 159146 197016
rect 171134 197004 171140 197056
rect 171192 197044 171198 197056
rect 200758 197044 200764 197056
rect 171192 197016 200764 197044
rect 171192 197004 171198 197016
rect 200758 197004 200764 197016
rect 200816 197004 200822 197056
rect 152826 196976 152832 196988
rect 134024 196948 142752 196976
rect 142816 196948 152832 196976
rect 134024 196936 134030 196948
rect 125410 196868 125416 196920
rect 125468 196908 125474 196920
rect 142816 196908 142844 196948
rect 152826 196936 152832 196948
rect 152884 196936 152890 196988
rect 166074 196936 166080 196988
rect 166132 196976 166138 196988
rect 200298 196976 200304 196988
rect 166132 196948 200304 196976
rect 166132 196936 166138 196948
rect 200298 196936 200304 196948
rect 200356 196936 200362 196988
rect 125468 196880 142844 196908
rect 125468 196868 125474 196880
rect 162762 196868 162768 196920
rect 162820 196908 162826 196920
rect 168558 196908 168564 196920
rect 162820 196880 168564 196908
rect 162820 196868 162826 196880
rect 168558 196868 168564 196880
rect 168616 196868 168622 196920
rect 168742 196868 168748 196920
rect 168800 196908 168806 196920
rect 169110 196908 169116 196920
rect 168800 196880 169116 196908
rect 168800 196868 168806 196880
rect 169110 196868 169116 196880
rect 169168 196868 169174 196920
rect 170398 196868 170404 196920
rect 170456 196908 170462 196920
rect 204714 196908 204720 196920
rect 170456 196880 204720 196908
rect 170456 196868 170462 196880
rect 204714 196868 204720 196880
rect 204772 196868 204778 196920
rect 104802 196800 104808 196852
rect 104860 196840 104866 196852
rect 138566 196840 138572 196852
rect 104860 196812 138572 196840
rect 104860 196800 104866 196812
rect 138566 196800 138572 196812
rect 138624 196800 138630 196852
rect 151906 196840 151912 196852
rect 139780 196812 151912 196840
rect 117958 196732 117964 196784
rect 118016 196772 118022 196784
rect 139780 196772 139808 196812
rect 151906 196800 151912 196812
rect 151964 196800 151970 196852
rect 152274 196800 152280 196852
rect 152332 196840 152338 196852
rect 153010 196840 153016 196852
rect 152332 196812 153016 196840
rect 152332 196800 152338 196812
rect 153010 196800 153016 196812
rect 153068 196800 153074 196852
rect 169018 196800 169024 196852
rect 169076 196840 169082 196852
rect 169294 196840 169300 196852
rect 169076 196812 169300 196840
rect 169076 196800 169082 196812
rect 169294 196800 169300 196812
rect 169352 196800 169358 196852
rect 169570 196800 169576 196852
rect 169628 196840 169634 196852
rect 169628 196812 173894 196840
rect 169628 196800 169634 196812
rect 118016 196744 139808 196772
rect 118016 196732 118022 196744
rect 141326 196732 141332 196784
rect 141384 196772 141390 196784
rect 142798 196772 142804 196784
rect 141384 196744 142804 196772
rect 141384 196732 141390 196744
rect 142798 196732 142804 196744
rect 142856 196732 142862 196784
rect 159174 196772 159180 196784
rect 147646 196744 159180 196772
rect 97718 196664 97724 196716
rect 97776 196704 97782 196716
rect 109034 196704 109040 196716
rect 97776 196676 109040 196704
rect 97776 196664 97782 196676
rect 109034 196664 109040 196676
rect 109092 196664 109098 196716
rect 117774 196664 117780 196716
rect 117832 196704 117838 196716
rect 147646 196704 147674 196744
rect 159174 196732 159180 196744
rect 159232 196772 159238 196784
rect 171778 196772 171784 196784
rect 159232 196744 171784 196772
rect 159232 196732 159238 196744
rect 171778 196732 171784 196744
rect 171836 196732 171842 196784
rect 171962 196732 171968 196784
rect 172020 196772 172026 196784
rect 173250 196772 173256 196784
rect 172020 196744 173256 196772
rect 172020 196732 172026 196744
rect 173250 196732 173256 196744
rect 173308 196732 173314 196784
rect 117832 196676 147674 196704
rect 117832 196664 117838 196676
rect 149790 196664 149796 196716
rect 149848 196704 149854 196716
rect 150066 196704 150072 196716
rect 149848 196676 150072 196704
rect 149848 196664 149854 196676
rect 150066 196664 150072 196676
rect 150124 196664 150130 196716
rect 150802 196664 150808 196716
rect 150860 196704 150866 196716
rect 153470 196704 153476 196716
rect 150860 196676 153476 196704
rect 150860 196664 150866 196676
rect 153470 196664 153476 196676
rect 153528 196664 153534 196716
rect 164234 196664 164240 196716
rect 164292 196704 164298 196716
rect 164510 196704 164516 196716
rect 164292 196676 164516 196704
rect 164292 196664 164298 196676
rect 164510 196664 164516 196676
rect 164568 196664 164574 196716
rect 166350 196664 166356 196716
rect 166408 196704 166414 196716
rect 166902 196704 166908 196716
rect 166408 196676 166908 196704
rect 166408 196664 166414 196676
rect 166902 196664 166908 196676
rect 166960 196664 166966 196716
rect 169846 196664 169852 196716
rect 169904 196704 169910 196716
rect 170674 196704 170680 196716
rect 169904 196676 170680 196704
rect 169904 196664 169910 196676
rect 170674 196664 170680 196676
rect 170732 196664 170738 196716
rect 173866 196704 173894 196812
rect 178402 196800 178408 196852
rect 178460 196840 178466 196852
rect 214190 196840 214196 196852
rect 178460 196812 214196 196840
rect 178460 196800 178466 196812
rect 214190 196800 214196 196812
rect 214248 196800 214254 196852
rect 178586 196732 178592 196784
rect 178644 196772 178650 196784
rect 213914 196772 213920 196784
rect 178644 196744 213920 196772
rect 178644 196732 178650 196744
rect 213914 196732 213920 196744
rect 213972 196732 213978 196784
rect 174538 196704 174544 196716
rect 173866 196676 174544 196704
rect 174538 196664 174544 196676
rect 174596 196664 174602 196716
rect 175182 196664 175188 196716
rect 175240 196704 175246 196716
rect 214006 196704 214012 196716
rect 175240 196676 214012 196704
rect 175240 196664 175246 196676
rect 214006 196664 214012 196676
rect 214064 196664 214070 196716
rect 102042 196596 102048 196648
rect 102100 196636 102106 196648
rect 135438 196636 135444 196648
rect 102100 196608 135444 196636
rect 102100 196596 102106 196608
rect 135438 196596 135444 196608
rect 135496 196596 135502 196648
rect 137462 196596 137468 196648
rect 137520 196636 137526 196648
rect 138566 196636 138572 196648
rect 137520 196608 138572 196636
rect 137520 196596 137526 196608
rect 138566 196596 138572 196608
rect 138624 196596 138630 196648
rect 146938 196596 146944 196648
rect 146996 196636 147002 196648
rect 149146 196636 149152 196648
rect 146996 196608 149152 196636
rect 146996 196596 147002 196608
rect 149146 196596 149152 196608
rect 149204 196596 149210 196648
rect 151630 196596 151636 196648
rect 151688 196636 151694 196648
rect 192754 196636 192760 196648
rect 151688 196608 192760 196636
rect 151688 196596 151694 196608
rect 192754 196596 192760 196608
rect 192812 196596 192818 196648
rect 145374 196528 145380 196580
rect 145432 196568 145438 196580
rect 145742 196568 145748 196580
rect 145432 196540 145748 196568
rect 145432 196528 145438 196540
rect 145742 196528 145748 196540
rect 145800 196528 145806 196580
rect 164510 196528 164516 196580
rect 164568 196568 164574 196580
rect 165154 196568 165160 196580
rect 164568 196540 165160 196568
rect 164568 196528 164574 196540
rect 165154 196528 165160 196540
rect 165212 196528 165218 196580
rect 165246 196528 165252 196580
rect 165304 196568 165310 196580
rect 165522 196568 165528 196580
rect 165304 196540 165528 196568
rect 165304 196528 165310 196540
rect 165522 196528 165528 196540
rect 165580 196528 165586 196580
rect 165890 196528 165896 196580
rect 165948 196568 165954 196580
rect 170398 196568 170404 196580
rect 165948 196540 170404 196568
rect 165948 196528 165954 196540
rect 170398 196528 170404 196540
rect 170456 196528 170462 196580
rect 171318 196528 171324 196580
rect 171376 196568 171382 196580
rect 171870 196568 171876 196580
rect 171376 196540 171876 196568
rect 171376 196528 171382 196540
rect 171870 196528 171876 196540
rect 171928 196528 171934 196580
rect 132218 196460 132224 196512
rect 132276 196500 132282 196512
rect 134978 196500 134984 196512
rect 132276 196472 134984 196500
rect 132276 196460 132282 196472
rect 134978 196460 134984 196472
rect 135036 196460 135042 196512
rect 137462 196460 137468 196512
rect 137520 196500 137526 196512
rect 144086 196500 144092 196512
rect 137520 196472 144092 196500
rect 137520 196460 137526 196472
rect 144086 196460 144092 196472
rect 144144 196460 144150 196512
rect 148502 196460 148508 196512
rect 148560 196500 148566 196512
rect 154114 196500 154120 196512
rect 148560 196472 154120 196500
rect 148560 196460 148566 196472
rect 154114 196460 154120 196472
rect 154172 196460 154178 196512
rect 168558 196460 168564 196512
rect 168616 196500 168622 196512
rect 169202 196500 169208 196512
rect 168616 196472 169208 196500
rect 168616 196460 168622 196472
rect 169202 196460 169208 196472
rect 169260 196460 169266 196512
rect 174170 196460 174176 196512
rect 174228 196500 174234 196512
rect 178218 196500 178224 196512
rect 174228 196472 178224 196500
rect 174228 196460 174234 196472
rect 178218 196460 178224 196472
rect 178276 196460 178282 196512
rect 107010 196392 107016 196444
rect 107068 196432 107074 196444
rect 107068 196404 157334 196432
rect 107068 196392 107074 196404
rect 131758 196324 131764 196376
rect 131816 196364 131822 196376
rect 139302 196364 139308 196376
rect 131816 196336 139308 196364
rect 131816 196324 131822 196336
rect 139302 196324 139308 196336
rect 139360 196324 139366 196376
rect 140038 196324 140044 196376
rect 140096 196364 140102 196376
rect 141786 196364 141792 196376
rect 140096 196336 141792 196364
rect 140096 196324 140102 196336
rect 141786 196324 141792 196336
rect 141844 196324 141850 196376
rect 142522 196324 142528 196376
rect 142580 196364 142586 196376
rect 143074 196364 143080 196376
rect 142580 196336 143080 196364
rect 142580 196324 142586 196336
rect 143074 196324 143080 196336
rect 143132 196324 143138 196376
rect 157306 196364 157334 196404
rect 170582 196364 170588 196376
rect 157306 196336 170588 196364
rect 170582 196324 170588 196336
rect 170640 196364 170646 196376
rect 176562 196364 176568 196376
rect 170640 196336 176568 196364
rect 170640 196324 170646 196336
rect 176562 196324 176568 196336
rect 176620 196324 176626 196376
rect 168098 196256 168104 196308
rect 168156 196296 168162 196308
rect 169202 196296 169208 196308
rect 168156 196268 169208 196296
rect 168156 196256 168162 196268
rect 169202 196256 169208 196268
rect 169260 196256 169266 196308
rect 134978 196188 134984 196240
rect 135036 196228 135042 196240
rect 135806 196228 135812 196240
rect 135036 196200 135812 196228
rect 135036 196188 135042 196200
rect 135806 196188 135812 196200
rect 135864 196188 135870 196240
rect 135990 196188 135996 196240
rect 136048 196228 136054 196240
rect 136174 196228 136180 196240
rect 136048 196200 136180 196228
rect 136048 196188 136054 196200
rect 136174 196188 136180 196200
rect 136232 196188 136238 196240
rect 144822 196188 144828 196240
rect 144880 196228 144886 196240
rect 145558 196228 145564 196240
rect 144880 196200 145564 196228
rect 144880 196188 144886 196200
rect 145558 196188 145564 196200
rect 145616 196188 145622 196240
rect 152550 196188 152556 196240
rect 152608 196228 152614 196240
rect 152734 196228 152740 196240
rect 152608 196200 152740 196228
rect 152608 196188 152614 196200
rect 152734 196188 152740 196200
rect 152792 196188 152798 196240
rect 167178 196188 167184 196240
rect 167236 196228 167242 196240
rect 167638 196228 167644 196240
rect 167236 196200 167644 196228
rect 167236 196188 167242 196200
rect 167638 196188 167644 196200
rect 167696 196188 167702 196240
rect 171226 196188 171232 196240
rect 171284 196228 171290 196240
rect 172238 196228 172244 196240
rect 171284 196200 172244 196228
rect 171284 196188 171290 196200
rect 172238 196188 172244 196200
rect 172296 196188 172302 196240
rect 134886 196120 134892 196172
rect 134944 196160 134950 196172
rect 135622 196160 135628 196172
rect 134944 196132 135628 196160
rect 134944 196120 134950 196132
rect 135622 196120 135628 196132
rect 135680 196120 135686 196172
rect 156598 196120 156604 196172
rect 156656 196160 156662 196172
rect 159542 196160 159548 196172
rect 156656 196132 159548 196160
rect 156656 196120 156662 196132
rect 159542 196120 159548 196132
rect 159600 196120 159606 196172
rect 175274 196120 175280 196172
rect 175332 196160 175338 196172
rect 176378 196160 176384 196172
rect 175332 196132 176384 196160
rect 175332 196120 175338 196132
rect 176378 196120 176384 196132
rect 176436 196120 176442 196172
rect 3602 196052 3608 196104
rect 3660 196092 3666 196104
rect 124398 196092 124404 196104
rect 3660 196064 124404 196092
rect 3660 196052 3666 196064
rect 124398 196052 124404 196064
rect 124456 196092 124462 196104
rect 125410 196092 125416 196104
rect 124456 196064 125416 196092
rect 124456 196052 124462 196064
rect 125410 196052 125416 196064
rect 125468 196052 125474 196104
rect 136174 196052 136180 196104
rect 136232 196092 136238 196104
rect 138198 196092 138204 196104
rect 136232 196064 138204 196092
rect 136232 196052 136238 196064
rect 138198 196052 138204 196064
rect 138256 196052 138262 196104
rect 143810 196092 143816 196104
rect 138308 196064 143816 196092
rect 3510 195984 3516 196036
rect 3568 196024 3574 196036
rect 128354 196024 128360 196036
rect 3568 195996 128360 196024
rect 3568 195984 3574 195996
rect 128354 195984 128360 195996
rect 128412 196024 128418 196036
rect 133966 196024 133972 196036
rect 128412 195996 133972 196024
rect 128412 195984 128418 195996
rect 133966 195984 133972 195996
rect 134024 195984 134030 196036
rect 135806 195984 135812 196036
rect 135864 196024 135870 196036
rect 136542 196024 136548 196036
rect 135864 195996 136548 196024
rect 135864 195984 135870 195996
rect 136542 195984 136548 195996
rect 136600 195984 136606 196036
rect 136910 195984 136916 196036
rect 136968 196024 136974 196036
rect 137094 196024 137100 196036
rect 136968 195996 137100 196024
rect 136968 195984 136974 195996
rect 137094 195984 137100 195996
rect 137152 195984 137158 196036
rect 138106 195984 138112 196036
rect 138164 196024 138170 196036
rect 138308 196024 138336 196064
rect 143810 196052 143816 196064
rect 143868 196052 143874 196104
rect 157794 196052 157800 196104
rect 157852 196092 157858 196104
rect 158346 196092 158352 196104
rect 157852 196064 158352 196092
rect 157852 196052 157858 196064
rect 158346 196052 158352 196064
rect 158404 196052 158410 196104
rect 175458 196052 175464 196104
rect 175516 196092 175522 196104
rect 176286 196092 176292 196104
rect 175516 196064 176292 196092
rect 175516 196052 175522 196064
rect 176286 196052 176292 196064
rect 176344 196052 176350 196104
rect 204438 196052 204444 196104
rect 204496 196092 204502 196104
rect 204714 196092 204720 196104
rect 204496 196064 204720 196092
rect 204496 196052 204502 196064
rect 204714 196052 204720 196064
rect 204772 196092 204778 196104
rect 580166 196092 580172 196104
rect 204772 196064 580172 196092
rect 204772 196052 204778 196064
rect 580166 196052 580172 196064
rect 580224 196052 580230 196104
rect 138164 195996 138336 196024
rect 138164 195984 138170 195996
rect 145558 195984 145564 196036
rect 145616 196024 145622 196036
rect 146294 196024 146300 196036
rect 145616 195996 146300 196024
rect 145616 195984 145622 195996
rect 146294 195984 146300 195996
rect 146352 195984 146358 196036
rect 147766 195984 147772 196036
rect 147824 196024 147830 196036
rect 148042 196024 148048 196036
rect 147824 195996 148048 196024
rect 147824 195984 147830 195996
rect 148042 195984 148048 195996
rect 148100 195984 148106 196036
rect 156966 195984 156972 196036
rect 157024 196024 157030 196036
rect 157242 196024 157248 196036
rect 157024 195996 157248 196024
rect 157024 195984 157030 195996
rect 157242 195984 157248 195996
rect 157300 195984 157306 196036
rect 161842 195984 161848 196036
rect 161900 196024 161906 196036
rect 162118 196024 162124 196036
rect 161900 195996 162124 196024
rect 161900 195984 161906 195996
rect 162118 195984 162124 195996
rect 162176 195984 162182 196036
rect 173986 195984 173992 196036
rect 174044 196024 174050 196036
rect 174998 196024 175004 196036
rect 174044 195996 175004 196024
rect 174044 195984 174050 195996
rect 174998 195984 175004 195996
rect 175056 195984 175062 196036
rect 175734 195984 175740 196036
rect 175792 196024 175798 196036
rect 176010 196024 176016 196036
rect 175792 195996 176016 196024
rect 175792 195984 175798 195996
rect 176010 195984 176016 195996
rect 176068 195984 176074 196036
rect 176746 195984 176752 196036
rect 176804 196024 176810 196036
rect 177298 196024 177304 196036
rect 176804 195996 177304 196024
rect 176804 195984 176810 195996
rect 177298 195984 177304 195996
rect 177356 195984 177362 196036
rect 186498 195984 186504 196036
rect 186556 196024 186562 196036
rect 187510 196024 187516 196036
rect 186556 195996 187516 196024
rect 186556 195984 186562 195996
rect 187510 195984 187516 195996
rect 187568 196024 187574 196036
rect 580626 196024 580632 196036
rect 187568 195996 580632 196024
rect 187568 195984 187574 195996
rect 580626 195984 580632 195996
rect 580684 195984 580690 196036
rect 130378 195916 130384 195968
rect 130436 195956 130442 195968
rect 132310 195956 132316 195968
rect 130436 195928 132316 195956
rect 130436 195916 130442 195928
rect 132310 195916 132316 195928
rect 132368 195956 132374 195968
rect 580258 195956 580264 195968
rect 132368 195928 580264 195956
rect 132368 195916 132374 195928
rect 580258 195916 580264 195928
rect 580316 195916 580322 195968
rect 109862 195848 109868 195900
rect 109920 195888 109926 195900
rect 142338 195888 142344 195900
rect 109920 195860 142344 195888
rect 109920 195848 109926 195860
rect 142338 195848 142344 195860
rect 142396 195888 142402 195900
rect 577682 195888 577688 195900
rect 142396 195860 577688 195888
rect 142396 195848 142402 195860
rect 577682 195848 577688 195860
rect 577740 195848 577746 195900
rect 104526 195780 104532 195832
rect 104584 195820 104590 195832
rect 138106 195820 138112 195832
rect 104584 195792 138112 195820
rect 104584 195780 104590 195792
rect 138106 195780 138112 195792
rect 138164 195780 138170 195832
rect 141970 195780 141976 195832
rect 142028 195820 142034 195832
rect 327718 195820 327724 195832
rect 142028 195792 327724 195820
rect 142028 195780 142034 195792
rect 327718 195780 327724 195792
rect 327776 195780 327782 195832
rect 104434 195712 104440 195764
rect 104492 195752 104498 195764
rect 176930 195752 176936 195764
rect 104492 195724 176936 195752
rect 104492 195712 104498 195724
rect 176930 195712 176936 195724
rect 176988 195712 176994 195764
rect 102962 195644 102968 195696
rect 103020 195684 103026 195696
rect 103020 195656 157334 195684
rect 103020 195644 103026 195656
rect 133046 195576 133052 195628
rect 133104 195616 133110 195628
rect 142798 195616 142804 195628
rect 133104 195588 142804 195616
rect 133104 195576 133110 195588
rect 142798 195576 142804 195588
rect 142856 195576 142862 195628
rect 154206 195576 154212 195628
rect 154264 195616 154270 195628
rect 155402 195616 155408 195628
rect 154264 195588 155408 195616
rect 154264 195576 154270 195588
rect 155402 195576 155408 195588
rect 155460 195576 155466 195628
rect 98822 195508 98828 195560
rect 98880 195548 98886 195560
rect 152550 195548 152556 195560
rect 98880 195520 152556 195548
rect 98880 195508 98886 195520
rect 152550 195508 152556 195520
rect 152608 195508 152614 195560
rect 97810 195440 97816 195492
rect 97868 195480 97874 195492
rect 152458 195480 152464 195492
rect 97868 195452 152464 195480
rect 97868 195440 97874 195452
rect 152458 195440 152464 195452
rect 152516 195440 152522 195492
rect 157306 195480 157334 195656
rect 160002 195644 160008 195696
rect 160060 195684 160066 195696
rect 160186 195684 160192 195696
rect 160060 195656 160192 195684
rect 160060 195644 160066 195656
rect 160186 195644 160192 195656
rect 160244 195644 160250 195696
rect 163590 195644 163596 195696
rect 163648 195684 163654 195696
rect 163648 195656 170352 195684
rect 163648 195644 163654 195656
rect 167270 195576 167276 195628
rect 167328 195616 167334 195628
rect 167822 195616 167828 195628
rect 167328 195588 167828 195616
rect 167328 195576 167334 195588
rect 167822 195576 167828 195588
rect 167880 195576 167886 195628
rect 160370 195508 160376 195560
rect 160428 195548 160434 195560
rect 161658 195548 161664 195560
rect 160428 195520 161664 195548
rect 160428 195508 160434 195520
rect 161658 195508 161664 195520
rect 161716 195508 161722 195560
rect 164142 195508 164148 195560
rect 164200 195548 164206 195560
rect 170324 195548 170352 195656
rect 170766 195644 170772 195696
rect 170824 195684 170830 195696
rect 193582 195684 193588 195696
rect 170824 195656 193588 195684
rect 170824 195644 170830 195656
rect 193582 195644 193588 195656
rect 193640 195644 193646 195696
rect 170490 195576 170496 195628
rect 170548 195616 170554 195628
rect 172882 195616 172888 195628
rect 170548 195588 172888 195616
rect 170548 195576 170554 195588
rect 172882 195576 172888 195588
rect 172940 195616 172946 195628
rect 193214 195616 193220 195628
rect 172940 195588 193220 195616
rect 172940 195576 172946 195588
rect 193214 195576 193220 195588
rect 193272 195576 193278 195628
rect 197998 195548 198004 195560
rect 164200 195520 168328 195548
rect 170324 195520 198004 195548
rect 164200 195508 164206 195520
rect 168300 195480 168328 195520
rect 197998 195508 198004 195520
rect 198056 195508 198062 195560
rect 157306 195452 164234 195480
rect 168300 195452 173894 195480
rect 96246 195372 96252 195424
rect 96304 195412 96310 195424
rect 155954 195412 155960 195424
rect 96304 195384 155960 195412
rect 96304 195372 96310 195384
rect 155954 195372 155960 195384
rect 156012 195372 156018 195424
rect 164206 195412 164234 195452
rect 170950 195412 170956 195424
rect 164206 195384 170956 195412
rect 170950 195372 170956 195384
rect 171008 195372 171014 195424
rect 173866 195412 173894 195452
rect 175826 195440 175832 195492
rect 175884 195480 175890 195492
rect 176286 195480 176292 195492
rect 175884 195452 176292 195480
rect 175884 195440 175890 195452
rect 176286 195440 176292 195452
rect 176344 195440 176350 195492
rect 176930 195440 176936 195492
rect 176988 195480 176994 195492
rect 178034 195480 178040 195492
rect 176988 195452 178040 195480
rect 176988 195440 176994 195452
rect 178034 195440 178040 195452
rect 178092 195480 178098 195492
rect 214282 195480 214288 195492
rect 178092 195452 214288 195480
rect 178092 195440 178098 195452
rect 214282 195440 214288 195452
rect 214340 195440 214346 195492
rect 204254 195412 204260 195424
rect 173866 195384 204260 195412
rect 204254 195372 204260 195384
rect 204312 195372 204318 195424
rect 3418 195304 3424 195356
rect 3476 195344 3482 195356
rect 3476 195316 157334 195344
rect 3476 195304 3482 195316
rect 120166 195236 120172 195288
rect 120224 195276 120230 195288
rect 121454 195276 121460 195288
rect 120224 195248 121460 195276
rect 120224 195236 120230 195248
rect 121454 195236 121460 195248
rect 121512 195236 121518 195288
rect 126330 195236 126336 195288
rect 126388 195276 126394 195288
rect 133046 195276 133052 195288
rect 126388 195248 133052 195276
rect 126388 195236 126394 195248
rect 133046 195236 133052 195248
rect 133104 195236 133110 195288
rect 138658 195236 138664 195288
rect 138716 195276 138722 195288
rect 140774 195276 140780 195288
rect 138716 195248 140780 195276
rect 138716 195236 138722 195248
rect 140774 195236 140780 195248
rect 140832 195236 140838 195288
rect 157306 195276 157334 195316
rect 160370 195304 160376 195356
rect 160428 195344 160434 195356
rect 160554 195344 160560 195356
rect 160428 195316 160560 195344
rect 160428 195304 160434 195316
rect 160554 195304 160560 195316
rect 160612 195304 160618 195356
rect 177298 195304 177304 195356
rect 177356 195344 177362 195356
rect 214558 195344 214564 195356
rect 177356 195316 214564 195344
rect 177356 195304 177362 195316
rect 214558 195304 214564 195316
rect 214616 195304 214622 195356
rect 167638 195276 167644 195288
rect 157306 195248 167644 195276
rect 167638 195236 167644 195248
rect 167696 195236 167702 195288
rect 200758 195236 200764 195288
rect 200816 195276 200822 195288
rect 214374 195276 214380 195288
rect 200816 195248 214380 195276
rect 200816 195236 200822 195248
rect 214374 195236 214380 195248
rect 214432 195276 214438 195288
rect 580810 195276 580816 195288
rect 214432 195248 580816 195276
rect 214432 195236 214438 195248
rect 580810 195236 580816 195248
rect 580868 195236 580874 195288
rect 111702 195168 111708 195220
rect 111760 195208 111766 195220
rect 143258 195208 143264 195220
rect 111760 195180 143264 195208
rect 111760 195168 111766 195180
rect 143258 195168 143264 195180
rect 143316 195168 143322 195220
rect 192018 195208 192024 195220
rect 167196 195180 192024 195208
rect 124122 195100 124128 195152
rect 124180 195140 124186 195152
rect 134978 195140 134984 195152
rect 124180 195112 134984 195140
rect 124180 195100 124186 195112
rect 134978 195100 134984 195112
rect 135036 195100 135042 195152
rect 152458 195100 152464 195152
rect 152516 195140 152522 195152
rect 156598 195140 156604 195152
rect 152516 195112 156604 195140
rect 152516 195100 152522 195112
rect 156598 195100 156604 195112
rect 156656 195100 156662 195152
rect 156690 195032 156696 195084
rect 156748 195072 156754 195084
rect 167196 195072 167224 195180
rect 192018 195168 192024 195180
rect 192076 195168 192082 195220
rect 168282 195100 168288 195152
rect 168340 195140 168346 195152
rect 175182 195140 175188 195152
rect 168340 195112 175188 195140
rect 168340 195100 168346 195112
rect 175182 195100 175188 195112
rect 175240 195100 175246 195152
rect 156748 195044 167224 195072
rect 156748 195032 156754 195044
rect 167730 195032 167736 195084
rect 167788 195072 167794 195084
rect 178678 195072 178684 195084
rect 167788 195044 178684 195072
rect 167788 195032 167794 195044
rect 178678 195032 178684 195044
rect 178736 195032 178742 195084
rect 142798 194964 142804 195016
rect 142856 195004 142862 195016
rect 149330 195004 149336 195016
rect 142856 194976 149336 195004
rect 142856 194964 142862 194976
rect 149330 194964 149336 194976
rect 149388 195004 149394 195016
rect 206278 195004 206284 195016
rect 149388 194976 206284 195004
rect 149388 194964 149394 194976
rect 206278 194964 206284 194976
rect 206336 194964 206342 195016
rect 108390 194896 108396 194948
rect 108448 194936 108454 194948
rect 108448 194908 157334 194936
rect 108448 194896 108454 194908
rect 157306 194868 157334 194908
rect 175182 194896 175188 194948
rect 175240 194936 175246 194948
rect 180058 194936 180064 194948
rect 175240 194908 180064 194936
rect 175240 194896 175246 194908
rect 180058 194896 180064 194908
rect 180116 194896 180122 194948
rect 174906 194868 174912 194880
rect 157306 194840 174912 194868
rect 174906 194828 174912 194840
rect 174964 194868 174970 194880
rect 177298 194868 177304 194880
rect 174964 194840 177304 194868
rect 174964 194828 174970 194840
rect 177298 194828 177304 194840
rect 177356 194828 177362 194880
rect 132034 194760 132040 194812
rect 132092 194800 132098 194812
rect 134518 194800 134524 194812
rect 132092 194772 134524 194800
rect 132092 194760 132098 194772
rect 134518 194760 134524 194772
rect 134576 194760 134582 194812
rect 152550 194760 152556 194812
rect 152608 194800 152614 194812
rect 157610 194800 157616 194812
rect 152608 194772 157616 194800
rect 152608 194760 152614 194772
rect 157610 194760 157616 194772
rect 157668 194800 157674 194812
rect 160738 194800 160744 194812
rect 157668 194772 160744 194800
rect 157668 194760 157674 194772
rect 160738 194760 160744 194772
rect 160796 194760 160802 194812
rect 139854 194556 139860 194608
rect 139912 194596 139918 194608
rect 142430 194596 142436 194608
rect 139912 194568 142436 194596
rect 139912 194556 139918 194568
rect 142430 194556 142436 194568
rect 142488 194556 142494 194608
rect 114830 194488 114836 194540
rect 114888 194528 114894 194540
rect 149238 194528 149244 194540
rect 114888 194500 149244 194528
rect 114888 194488 114894 194500
rect 149238 194488 149244 194500
rect 149296 194488 149302 194540
rect 149790 194488 149796 194540
rect 149848 194528 149854 194540
rect 152734 194528 152740 194540
rect 149848 194500 152740 194528
rect 149848 194488 149854 194500
rect 152734 194488 152740 194500
rect 152792 194528 152798 194540
rect 578970 194528 578976 194540
rect 152792 194500 578976 194528
rect 152792 194488 152798 194500
rect 578970 194488 578976 194500
rect 579028 194488 579034 194540
rect 107102 194420 107108 194472
rect 107160 194460 107166 194472
rect 114462 194460 114468 194472
rect 107160 194432 114468 194460
rect 107160 194420 107166 194432
rect 114462 194420 114468 194432
rect 114520 194420 114526 194472
rect 122098 194420 122104 194472
rect 122156 194460 122162 194472
rect 141510 194460 141516 194472
rect 122156 194432 141516 194460
rect 122156 194420 122162 194432
rect 141510 194420 141516 194432
rect 141568 194420 141574 194472
rect 142614 194420 142620 194472
rect 142672 194460 142678 194472
rect 567838 194460 567844 194472
rect 142672 194432 567844 194460
rect 142672 194420 142678 194432
rect 567838 194420 567844 194432
rect 567896 194420 567902 194472
rect 107470 194352 107476 194404
rect 107528 194392 107534 194404
rect 118694 194392 118700 194404
rect 107528 194364 118700 194392
rect 107528 194352 107534 194364
rect 118694 194352 118700 194364
rect 118752 194352 118758 194404
rect 139946 194352 139952 194404
rect 140004 194392 140010 194404
rect 564066 194392 564072 194404
rect 140004 194364 564072 194392
rect 140004 194352 140010 194364
rect 564066 194352 564072 194364
rect 564124 194352 564130 194404
rect 104250 194284 104256 194336
rect 104308 194324 104314 194336
rect 177114 194324 177120 194336
rect 104308 194296 177120 194324
rect 104308 194284 104314 194296
rect 177114 194284 177120 194296
rect 177172 194284 177178 194336
rect 107194 194216 107200 194268
rect 107252 194256 107258 194268
rect 161934 194256 161940 194268
rect 107252 194228 161940 194256
rect 107252 194216 107258 194228
rect 161934 194216 161940 194228
rect 161992 194216 161998 194268
rect 174354 194216 174360 194268
rect 174412 194256 174418 194268
rect 192294 194256 192300 194268
rect 174412 194228 192300 194256
rect 174412 194216 174418 194228
rect 192294 194216 192300 194228
rect 192352 194216 192358 194268
rect 108666 194148 108672 194200
rect 108724 194188 108730 194200
rect 163314 194188 163320 194200
rect 108724 194160 163320 194188
rect 108724 194148 108730 194160
rect 163314 194148 163320 194160
rect 163372 194188 163378 194200
rect 163590 194188 163596 194200
rect 163372 194160 163596 194188
rect 163372 194148 163378 194160
rect 163590 194148 163596 194160
rect 163648 194148 163654 194200
rect 174078 194148 174084 194200
rect 174136 194188 174142 194200
rect 175090 194188 175096 194200
rect 174136 194160 175096 194188
rect 174136 194148 174142 194160
rect 175090 194148 175096 194160
rect 175148 194148 175154 194200
rect 176470 194148 176476 194200
rect 176528 194188 176534 194200
rect 198826 194188 198832 194200
rect 176528 194160 198832 194188
rect 176528 194148 176534 194160
rect 198826 194148 198832 194160
rect 198884 194148 198890 194200
rect 107010 194080 107016 194132
rect 107068 194120 107074 194132
rect 139946 194120 139952 194132
rect 107068 194092 139952 194120
rect 107068 194080 107074 194092
rect 139946 194080 139952 194092
rect 140004 194080 140010 194132
rect 157702 194080 157708 194132
rect 157760 194120 157766 194132
rect 158438 194120 158444 194132
rect 157760 194092 158444 194120
rect 157760 194080 157766 194092
rect 158438 194080 158444 194092
rect 158496 194080 158502 194132
rect 158714 194080 158720 194132
rect 158772 194120 158778 194132
rect 185762 194120 185768 194132
rect 158772 194092 185768 194120
rect 158772 194080 158778 194092
rect 185762 194080 185768 194092
rect 185820 194080 185826 194132
rect 189534 194080 189540 194132
rect 189592 194120 189598 194132
rect 189592 194092 190454 194120
rect 189592 194080 189598 194092
rect 104710 194012 104716 194064
rect 104768 194052 104774 194064
rect 135070 194052 135076 194064
rect 104768 194024 135076 194052
rect 104768 194012 104774 194024
rect 135070 194012 135076 194024
rect 135128 194012 135134 194064
rect 162394 194012 162400 194064
rect 162452 194052 162458 194064
rect 189718 194052 189724 194064
rect 162452 194024 189724 194052
rect 162452 194012 162458 194024
rect 189718 194012 189724 194024
rect 189776 194012 189782 194064
rect 190426 194052 190454 194092
rect 209866 194052 209872 194064
rect 190426 194024 209872 194052
rect 209866 194012 209872 194024
rect 209924 194012 209930 194064
rect 95602 193944 95608 193996
rect 95660 193984 95666 193996
rect 110506 193984 110512 193996
rect 95660 193956 110512 193984
rect 95660 193944 95666 193956
rect 110506 193944 110512 193956
rect 110564 193984 110570 193996
rect 111794 193984 111800 193996
rect 110564 193956 111800 193984
rect 110564 193944 110570 193956
rect 111794 193944 111800 193956
rect 111852 193944 111858 193996
rect 118418 193944 118424 193996
rect 118476 193984 118482 193996
rect 149790 193984 149796 193996
rect 118476 193956 149796 193984
rect 118476 193944 118482 193956
rect 149790 193944 149796 193956
rect 149848 193944 149854 193996
rect 166166 193944 166172 193996
rect 166224 193984 166230 193996
rect 172146 193984 172152 193996
rect 166224 193956 172152 193984
rect 166224 193944 166230 193956
rect 172146 193944 172152 193956
rect 172204 193944 172210 193996
rect 172790 193944 172796 193996
rect 172848 193984 172854 193996
rect 207014 193984 207020 193996
rect 172848 193956 207020 193984
rect 172848 193944 172854 193956
rect 207014 193944 207020 193956
rect 207072 193944 207078 193996
rect 101950 193876 101956 193928
rect 102008 193916 102014 193928
rect 140682 193916 140688 193928
rect 102008 193888 140688 193916
rect 102008 193876 102014 193888
rect 140682 193876 140688 193888
rect 140740 193876 140746 193928
rect 157426 193876 157432 193928
rect 157484 193916 157490 193928
rect 173158 193916 173164 193928
rect 157484 193888 173164 193916
rect 157484 193876 157490 193888
rect 173158 193876 173164 193888
rect 173216 193876 173222 193928
rect 177114 193876 177120 193928
rect 177172 193916 177178 193928
rect 212718 193916 212724 193928
rect 177172 193888 212724 193916
rect 177172 193876 177178 193888
rect 212718 193876 212724 193888
rect 212776 193876 212782 193928
rect 99374 193808 99380 193860
rect 99432 193848 99438 193860
rect 103330 193848 103336 193860
rect 99432 193820 103336 193848
rect 99432 193808 99438 193820
rect 103330 193808 103336 193820
rect 103388 193848 103394 193860
rect 158622 193848 158628 193860
rect 103388 193820 158628 193848
rect 103388 193808 103394 193820
rect 158622 193808 158628 193820
rect 158680 193808 158686 193860
rect 171410 193808 171416 193860
rect 171468 193848 171474 193860
rect 205726 193848 205732 193860
rect 171468 193820 205732 193848
rect 171468 193808 171474 193820
rect 205726 193808 205732 193820
rect 205784 193808 205790 193860
rect 207014 193808 207020 193860
rect 207072 193848 207078 193860
rect 502334 193848 502340 193860
rect 207072 193820 502340 193848
rect 207072 193808 207078 193820
rect 502334 193808 502340 193820
rect 502392 193808 502398 193860
rect 116302 193740 116308 193792
rect 116360 193780 116366 193792
rect 148318 193780 148324 193792
rect 116360 193752 148324 193780
rect 116360 193740 116366 193752
rect 148318 193740 148324 193752
rect 148376 193740 148382 193792
rect 161658 193740 161664 193792
rect 161716 193780 161722 193792
rect 178954 193780 178960 193792
rect 161716 193752 178960 193780
rect 161716 193740 161722 193752
rect 178954 193740 178960 193752
rect 179012 193740 179018 193792
rect 119982 193672 119988 193724
rect 120040 193712 120046 193724
rect 148594 193712 148600 193724
rect 120040 193684 148600 193712
rect 120040 193672 120046 193684
rect 148594 193672 148600 193684
rect 148652 193672 148658 193724
rect 172974 193672 172980 193724
rect 173032 193712 173038 193724
rect 173342 193712 173348 193724
rect 173032 193684 173348 193712
rect 173032 193672 173038 193684
rect 173342 193672 173348 193684
rect 173400 193672 173406 193724
rect 131022 193604 131028 193656
rect 131080 193644 131086 193656
rect 161198 193644 161204 193656
rect 131080 193616 161204 193644
rect 131080 193604 131086 193616
rect 161198 193604 161204 193616
rect 161256 193604 161262 193656
rect 169938 193604 169944 193656
rect 169996 193644 170002 193656
rect 170858 193644 170864 193656
rect 169996 193616 170864 193644
rect 169996 193604 170002 193616
rect 170858 193604 170864 193616
rect 170916 193604 170922 193656
rect 138014 193536 138020 193588
rect 138072 193576 138078 193588
rect 138934 193576 138940 193588
rect 138072 193548 138940 193576
rect 138072 193536 138078 193548
rect 138934 193536 138940 193548
rect 138992 193536 138998 193588
rect 144178 193536 144184 193588
rect 144236 193576 144242 193588
rect 144914 193576 144920 193588
rect 144236 193548 144920 193576
rect 144236 193536 144242 193548
rect 144914 193536 144920 193548
rect 144972 193536 144978 193588
rect 152550 193536 152556 193588
rect 152608 193576 152614 193588
rect 152918 193576 152924 193588
rect 152608 193548 152924 193576
rect 152608 193536 152614 193548
rect 152918 193536 152924 193548
rect 152976 193536 152982 193588
rect 164602 193400 164608 193452
rect 164660 193440 164666 193452
rect 165430 193440 165436 193452
rect 164660 193412 165436 193440
rect 164660 193400 164666 193412
rect 165430 193400 165436 193412
rect 165488 193400 165494 193452
rect 168466 193400 168472 193452
rect 168524 193440 168530 193452
rect 169478 193440 169484 193452
rect 168524 193412 169484 193440
rect 168524 193400 168530 193412
rect 169478 193400 169484 193412
rect 169536 193400 169542 193452
rect 152918 193332 152924 193384
rect 152976 193372 152982 193384
rect 152976 193344 157334 193372
rect 152976 193332 152982 193344
rect 104618 193196 104624 193248
rect 104676 193236 104682 193248
rect 157306 193236 157334 193344
rect 177298 193264 177304 193316
rect 177356 193304 177362 193316
rect 189350 193304 189356 193316
rect 177356 193276 189356 193304
rect 177356 193264 177362 193276
rect 189350 193264 189356 193276
rect 189408 193264 189414 193316
rect 198090 193236 198096 193248
rect 104676 193208 110460 193236
rect 157306 193208 198096 193236
rect 104676 193196 104682 193208
rect 110432 193032 110460 193208
rect 198090 193196 198096 193208
rect 198148 193196 198154 193248
rect 147306 193168 147312 193180
rect 143506 193140 147312 193168
rect 111794 193060 111800 193112
rect 111852 193100 111858 193112
rect 143506 193100 143534 193140
rect 147306 193128 147312 193140
rect 147364 193128 147370 193180
rect 168374 193128 168380 193180
rect 168432 193168 168438 193180
rect 577590 193168 577596 193180
rect 168432 193140 577596 193168
rect 168432 193128 168438 193140
rect 577590 193128 577596 193140
rect 577648 193128 577654 193180
rect 111852 193072 143534 193100
rect 111852 193060 111858 193072
rect 145098 193060 145104 193112
rect 145156 193100 145162 193112
rect 281534 193100 281540 193112
rect 145156 193072 281540 193100
rect 145156 193060 145162 193072
rect 281534 193060 281540 193072
rect 281592 193060 281598 193112
rect 111334 193032 111340 193044
rect 110432 193004 111340 193032
rect 111334 192992 111340 193004
rect 111392 193032 111398 193044
rect 141326 193032 141332 193044
rect 111392 193004 141332 193032
rect 111392 192992 111398 193004
rect 141326 192992 141332 193004
rect 141384 192992 141390 193044
rect 148594 192992 148600 193044
rect 148652 193032 148658 193044
rect 151078 193032 151084 193044
rect 148652 193004 151084 193032
rect 148652 192992 148658 193004
rect 151078 192992 151084 193004
rect 151136 193032 151142 193044
rect 189442 193032 189448 193044
rect 151136 193004 189448 193032
rect 151136 192992 151142 193004
rect 189442 192992 189448 193004
rect 189500 192992 189506 193044
rect 114462 192924 114468 192976
rect 114520 192964 114526 192976
rect 136726 192964 136732 192976
rect 114520 192936 136732 192964
rect 114520 192924 114526 192936
rect 136726 192924 136732 192936
rect 136784 192924 136790 192976
rect 173618 192924 173624 192976
rect 173676 192964 173682 192976
rect 198734 192964 198740 192976
rect 173676 192936 198740 192964
rect 173676 192924 173682 192936
rect 198734 192924 198740 192936
rect 198792 192924 198798 192976
rect 120166 192856 120172 192908
rect 120224 192896 120230 192908
rect 138290 192896 138296 192908
rect 120224 192868 138296 192896
rect 120224 192856 120230 192868
rect 138290 192856 138296 192868
rect 138348 192856 138354 192908
rect 173250 192856 173256 192908
rect 173308 192896 173314 192908
rect 206186 192896 206192 192908
rect 173308 192868 206192 192896
rect 173308 192856 173314 192868
rect 206186 192856 206192 192868
rect 206244 192856 206250 192908
rect 118234 192788 118240 192840
rect 118292 192828 118298 192840
rect 139486 192828 139492 192840
rect 118292 192800 139492 192828
rect 118292 192788 118298 192800
rect 139486 192788 139492 192800
rect 139544 192788 139550 192840
rect 169294 192788 169300 192840
rect 169352 192828 169358 192840
rect 202874 192828 202880 192840
rect 169352 192800 202880 192828
rect 169352 192788 169358 192800
rect 202874 192788 202880 192800
rect 202932 192788 202938 192840
rect 127618 192720 127624 192772
rect 127676 192760 127682 192772
rect 153746 192760 153752 192772
rect 127676 192732 153752 192760
rect 127676 192720 127682 192732
rect 153746 192720 153752 192732
rect 153804 192720 153810 192772
rect 162486 192720 162492 192772
rect 162544 192760 162550 192772
rect 196066 192760 196072 192772
rect 162544 192732 196072 192760
rect 162544 192720 162550 192732
rect 196066 192720 196072 192732
rect 196124 192720 196130 192772
rect 121270 192652 121276 192704
rect 121328 192692 121334 192704
rect 150802 192692 150808 192704
rect 121328 192664 150808 192692
rect 121328 192652 121334 192664
rect 150802 192652 150808 192664
rect 150860 192652 150866 192704
rect 154022 192652 154028 192704
rect 154080 192692 154086 192704
rect 196710 192692 196716 192704
rect 154080 192664 196716 192692
rect 154080 192652 154086 192664
rect 196710 192652 196716 192664
rect 196768 192652 196774 192704
rect 119522 192584 119528 192636
rect 119580 192624 119586 192636
rect 144822 192624 144828 192636
rect 119580 192596 144828 192624
rect 119580 192584 119586 192596
rect 144822 192584 144828 192596
rect 144880 192584 144886 192636
rect 146754 192584 146760 192636
rect 146812 192624 146818 192636
rect 191834 192624 191840 192636
rect 146812 192596 191840 192624
rect 146812 192584 146818 192596
rect 191834 192584 191840 192596
rect 191892 192584 191898 192636
rect 202874 192584 202880 192636
rect 202932 192624 202938 192636
rect 575106 192624 575112 192636
rect 202932 192596 575112 192624
rect 202932 192584 202938 192596
rect 575106 192584 575112 192596
rect 575164 192584 575170 192636
rect 114462 192516 114468 192568
rect 114520 192556 114526 192568
rect 139854 192556 139860 192568
rect 114520 192528 139860 192556
rect 114520 192516 114526 192528
rect 139854 192516 139860 192528
rect 139912 192516 139918 192568
rect 544378 192556 544384 192568
rect 148704 192528 544384 192556
rect 86310 192448 86316 192500
rect 86368 192488 86374 192500
rect 120166 192488 120172 192500
rect 86368 192460 120172 192488
rect 86368 192448 86374 192460
rect 120166 192448 120172 192460
rect 120224 192448 120230 192500
rect 126422 192448 126428 192500
rect 126480 192488 126486 192500
rect 148594 192488 148600 192500
rect 126480 192460 148600 192488
rect 126480 192448 126486 192460
rect 148594 192448 148600 192460
rect 148652 192448 148658 192500
rect 121822 192380 121828 192432
rect 121880 192420 121886 192432
rect 135622 192420 135628 192432
rect 121880 192392 135628 192420
rect 121880 192380 121886 192392
rect 135622 192380 135628 192392
rect 135680 192380 135686 192432
rect 131942 192312 131948 192364
rect 132000 192352 132006 192364
rect 145466 192352 145472 192364
rect 132000 192324 145472 192352
rect 132000 192312 132006 192324
rect 145466 192312 145472 192324
rect 145524 192352 145530 192364
rect 148704 192352 148732 192528
rect 544378 192516 544384 192528
rect 544436 192516 544442 192568
rect 150342 192448 150348 192500
rect 150400 192488 150406 192500
rect 579614 192488 579620 192500
rect 150400 192460 579620 192488
rect 150400 192448 150406 192460
rect 579614 192448 579620 192460
rect 579672 192448 579678 192500
rect 167546 192380 167552 192432
rect 167604 192420 167610 192432
rect 184198 192420 184204 192432
rect 167604 192392 184204 192420
rect 167604 192380 167610 192392
rect 184198 192380 184204 192392
rect 184256 192380 184262 192432
rect 145524 192324 148732 192352
rect 145524 192312 145530 192324
rect 169754 192312 169760 192364
rect 169812 192352 169818 192364
rect 178034 192352 178040 192364
rect 169812 192324 178040 192352
rect 169812 192312 169818 192324
rect 178034 192312 178040 192324
rect 178092 192312 178098 192364
rect 94774 192244 94780 192296
rect 94832 192284 94838 192296
rect 173250 192284 173256 192296
rect 94832 192256 173256 192284
rect 94832 192244 94838 192256
rect 173250 192244 173256 192256
rect 173308 192244 173314 192296
rect 25498 191836 25504 191888
rect 25556 191876 25562 191888
rect 125686 191876 125692 191888
rect 25556 191848 125692 191876
rect 25556 191836 25562 191848
rect 125686 191836 125692 191848
rect 125744 191836 125750 191888
rect 133800 191848 134380 191876
rect 101490 191768 101496 191820
rect 101548 191808 101554 191820
rect 118142 191808 118148 191820
rect 101548 191780 118148 191808
rect 101548 191768 101554 191780
rect 118142 191768 118148 191780
rect 118200 191768 118206 191820
rect 127710 191768 127716 191820
rect 127768 191808 127774 191820
rect 128446 191808 128452 191820
rect 127768 191780 128452 191808
rect 127768 191768 127774 191780
rect 128446 191768 128452 191780
rect 128504 191768 128510 191820
rect 130470 191768 130476 191820
rect 130528 191808 130534 191820
rect 133800 191808 133828 191848
rect 130528 191780 133828 191808
rect 130528 191768 130534 191780
rect 133874 191768 133880 191820
rect 133932 191808 133938 191820
rect 134242 191808 134248 191820
rect 133932 191780 134248 191808
rect 133932 191768 133938 191780
rect 134242 191768 134248 191780
rect 134300 191768 134306 191820
rect 134352 191808 134380 191848
rect 174998 191836 175004 191888
rect 175056 191876 175062 191888
rect 182910 191876 182916 191888
rect 175056 191848 182916 191876
rect 175056 191836 175062 191848
rect 182910 191836 182916 191848
rect 182968 191836 182974 191888
rect 145006 191808 145012 191820
rect 134352 191780 145012 191808
rect 145006 191768 145012 191780
rect 145064 191808 145070 191820
rect 575014 191808 575020 191820
rect 145064 191780 575020 191808
rect 145064 191768 145070 191780
rect 575014 191768 575020 191780
rect 575072 191768 575078 191820
rect 57974 191700 57980 191752
rect 58032 191740 58038 191752
rect 158622 191740 158628 191752
rect 58032 191712 158628 191740
rect 58032 191700 58038 191712
rect 158622 191700 158628 191712
rect 158680 191740 158686 191752
rect 160922 191740 160928 191752
rect 158680 191712 160928 191740
rect 158680 191700 158686 191712
rect 160922 191700 160928 191712
rect 160980 191700 160986 191752
rect 174170 191700 174176 191752
rect 174228 191740 174234 191752
rect 174722 191740 174728 191752
rect 174228 191712 174728 191740
rect 174228 191700 174234 191712
rect 174722 191700 174728 191712
rect 174780 191700 174786 191752
rect 197998 191700 198004 191752
rect 198056 191740 198062 191752
rect 572254 191740 572260 191752
rect 198056 191712 572260 191740
rect 198056 191700 198062 191712
rect 572254 191700 572260 191712
rect 572312 191700 572318 191752
rect 101398 191632 101404 191684
rect 101456 191672 101462 191684
rect 184934 191672 184940 191684
rect 101456 191644 184940 191672
rect 101456 191632 101462 191644
rect 184934 191632 184940 191644
rect 184992 191632 184998 191684
rect 197722 191632 197728 191684
rect 197780 191672 197786 191684
rect 566458 191672 566464 191684
rect 197780 191644 566464 191672
rect 197780 191632 197786 191644
rect 566458 191632 566464 191644
rect 566516 191632 566522 191684
rect 99006 191564 99012 191616
rect 99064 191604 99070 191616
rect 165246 191604 165252 191616
rect 99064 191576 165252 191604
rect 99064 191564 99070 191576
rect 165246 191564 165252 191576
rect 165304 191564 165310 191616
rect 175918 191564 175924 191616
rect 175976 191604 175982 191616
rect 398834 191604 398840 191616
rect 175976 191576 398840 191604
rect 175976 191564 175982 191576
rect 398834 191564 398840 191576
rect 398892 191564 398898 191616
rect 95878 191496 95884 191548
rect 95936 191536 95942 191548
rect 159450 191536 159456 191548
rect 95936 191508 159456 191536
rect 95936 191496 95942 191508
rect 159450 191496 159456 191508
rect 159508 191536 159514 191548
rect 178862 191536 178868 191548
rect 159508 191508 178868 191536
rect 159508 191496 159514 191508
rect 178862 191496 178868 191508
rect 178920 191496 178926 191548
rect 104066 191428 104072 191480
rect 104124 191468 104130 191480
rect 108666 191468 108672 191480
rect 104124 191440 108672 191468
rect 104124 191428 104130 191440
rect 108666 191428 108672 191440
rect 108724 191428 108730 191480
rect 112990 191428 112996 191480
rect 113048 191468 113054 191480
rect 168926 191468 168932 191480
rect 113048 191440 168932 191468
rect 113048 191428 113054 191440
rect 168926 191428 168932 191440
rect 168984 191428 168990 191480
rect 184842 191428 184848 191480
rect 184900 191468 184906 191480
rect 195974 191468 195980 191480
rect 184900 191440 195980 191468
rect 184900 191428 184906 191440
rect 195974 191428 195980 191440
rect 196032 191428 196038 191480
rect 100478 191360 100484 191412
rect 100536 191400 100542 191412
rect 133874 191400 133880 191412
rect 100536 191372 133880 191400
rect 100536 191360 100542 191372
rect 133874 191360 133880 191372
rect 133932 191360 133938 191412
rect 134150 191360 134156 191412
rect 134208 191400 134214 191412
rect 134426 191400 134432 191412
rect 134208 191372 134432 191400
rect 134208 191360 134214 191372
rect 134426 191360 134432 191372
rect 134484 191360 134490 191412
rect 135714 191360 135720 191412
rect 135772 191400 135778 191412
rect 136358 191400 136364 191412
rect 135772 191372 136364 191400
rect 135772 191360 135778 191372
rect 136358 191360 136364 191372
rect 136416 191360 136422 191412
rect 137370 191360 137376 191412
rect 137428 191400 137434 191412
rect 137922 191400 137928 191412
rect 137428 191372 137928 191400
rect 137428 191360 137434 191372
rect 137922 191360 137928 191372
rect 137980 191360 137986 191412
rect 138106 191360 138112 191412
rect 138164 191400 138170 191412
rect 143902 191400 143908 191412
rect 138164 191372 143908 191400
rect 138164 191360 138170 191372
rect 143902 191360 143908 191372
rect 143960 191360 143966 191412
rect 148686 191360 148692 191412
rect 148744 191400 148750 191412
rect 148870 191400 148876 191412
rect 148744 191372 148876 191400
rect 148744 191360 148750 191372
rect 148870 191360 148876 191372
rect 148928 191360 148934 191412
rect 160094 191360 160100 191412
rect 160152 191400 160158 191412
rect 160554 191400 160560 191412
rect 160152 191372 160560 191400
rect 160152 191360 160158 191372
rect 160554 191360 160560 191372
rect 160612 191360 160618 191412
rect 160922 191360 160928 191412
rect 160980 191400 160986 191412
rect 178770 191400 178776 191412
rect 160980 191372 178776 191400
rect 160980 191360 160986 191372
rect 178770 191360 178776 191372
rect 178828 191360 178834 191412
rect 184934 191360 184940 191412
rect 184992 191400 184998 191412
rect 200390 191400 200396 191412
rect 184992 191372 200396 191400
rect 184992 191360 184998 191372
rect 200390 191360 200396 191372
rect 200448 191360 200454 191412
rect 108666 191292 108672 191344
rect 108724 191332 108730 191344
rect 143166 191332 143172 191344
rect 108724 191304 143172 191332
rect 108724 191292 108730 191304
rect 143166 191292 143172 191304
rect 143224 191292 143230 191344
rect 156414 191332 156420 191344
rect 147646 191304 156420 191332
rect 115842 191224 115848 191276
rect 115900 191264 115906 191276
rect 122006 191264 122012 191276
rect 115900 191236 122012 191264
rect 115900 191224 115906 191236
rect 122006 191224 122012 191236
rect 122064 191264 122070 191276
rect 147646 191264 147674 191304
rect 156414 191292 156420 191304
rect 156472 191292 156478 191344
rect 160278 191292 160284 191344
rect 160336 191332 160342 191344
rect 194594 191332 194600 191344
rect 160336 191304 194600 191332
rect 160336 191292 160342 191304
rect 194594 191292 194600 191304
rect 194652 191292 194658 191344
rect 197354 191292 197360 191344
rect 197412 191332 197418 191344
rect 216858 191332 216864 191344
rect 197412 191304 216864 191332
rect 197412 191292 197418 191304
rect 216858 191292 216864 191304
rect 216916 191292 216922 191344
rect 122064 191236 147674 191264
rect 122064 191224 122070 191236
rect 153286 191224 153292 191276
rect 153344 191264 153350 191276
rect 154114 191264 154120 191276
rect 153344 191236 154120 191264
rect 153344 191224 153350 191236
rect 154114 191224 154120 191236
rect 154172 191224 154178 191276
rect 158990 191224 158996 191276
rect 159048 191264 159054 191276
rect 159910 191264 159916 191276
rect 159048 191236 159916 191264
rect 159048 191224 159054 191236
rect 159910 191224 159916 191236
rect 159968 191224 159974 191276
rect 162762 191224 162768 191276
rect 162820 191264 162826 191276
rect 164418 191264 164424 191276
rect 162820 191236 164424 191264
rect 162820 191224 162826 191236
rect 164418 191224 164424 191236
rect 164476 191224 164482 191276
rect 164510 191224 164516 191276
rect 164568 191264 164574 191276
rect 164568 191236 166396 191264
rect 164568 191224 164574 191236
rect 105906 191196 105912 191208
rect 103486 191168 105912 191196
rect 84930 191088 84936 191140
rect 84988 191128 84994 191140
rect 103486 191128 103514 191168
rect 105906 191156 105912 191168
rect 105964 191196 105970 191208
rect 138106 191196 138112 191208
rect 105964 191168 138112 191196
rect 105964 191156 105970 191168
rect 138106 191156 138112 191168
rect 138164 191156 138170 191208
rect 138290 191156 138296 191208
rect 138348 191196 138354 191208
rect 139026 191196 139032 191208
rect 138348 191168 139032 191196
rect 138348 191156 138354 191168
rect 139026 191156 139032 191168
rect 139084 191156 139090 191208
rect 140130 191156 140136 191208
rect 140188 191196 140194 191208
rect 140682 191196 140688 191208
rect 140188 191168 140688 191196
rect 140188 191156 140194 191168
rect 140682 191156 140688 191168
rect 140740 191156 140746 191208
rect 142798 191156 142804 191208
rect 142856 191196 142862 191208
rect 142982 191196 142988 191208
rect 142856 191168 142988 191196
rect 142856 191156 142862 191168
rect 142982 191156 142988 191168
rect 143040 191156 143046 191208
rect 145466 191156 145472 191208
rect 145524 191196 145530 191208
rect 146018 191196 146024 191208
rect 145524 191168 146024 191196
rect 145524 191156 145530 191168
rect 146018 191156 146024 191168
rect 146076 191156 146082 191208
rect 146478 191156 146484 191208
rect 146536 191196 146542 191208
rect 147122 191196 147128 191208
rect 146536 191168 147128 191196
rect 146536 191156 146542 191168
rect 147122 191156 147128 191168
rect 147180 191156 147186 191208
rect 149146 191156 149152 191208
rect 149204 191196 149210 191208
rect 149882 191196 149888 191208
rect 149204 191168 149888 191196
rect 149204 191156 149210 191168
rect 149882 191156 149888 191168
rect 149940 191156 149946 191208
rect 150618 191156 150624 191208
rect 150676 191196 150682 191208
rect 151354 191196 151360 191208
rect 150676 191168 151360 191196
rect 150676 191156 150682 191168
rect 151354 191156 151360 191168
rect 151412 191156 151418 191208
rect 153470 191156 153476 191208
rect 153528 191196 153534 191208
rect 154390 191196 154396 191208
rect 153528 191168 154396 191196
rect 153528 191156 153534 191168
rect 154390 191156 154396 191168
rect 154448 191156 154454 191208
rect 154942 191156 154948 191208
rect 155000 191196 155006 191208
rect 155494 191196 155500 191208
rect 155000 191168 155500 191196
rect 155000 191156 155006 191168
rect 155494 191156 155500 191168
rect 155552 191156 155558 191208
rect 156138 191156 156144 191208
rect 156196 191196 156202 191208
rect 156966 191196 156972 191208
rect 156196 191168 156972 191196
rect 156196 191156 156202 191168
rect 156966 191156 156972 191168
rect 157024 191156 157030 191208
rect 158898 191156 158904 191208
rect 158956 191196 158962 191208
rect 159726 191196 159732 191208
rect 158956 191168 159732 191196
rect 158956 191156 158962 191168
rect 159726 191156 159732 191168
rect 159784 191156 159790 191208
rect 160186 191156 160192 191208
rect 160244 191196 160250 191208
rect 160462 191196 160468 191208
rect 160244 191168 160468 191196
rect 160244 191156 160250 191168
rect 160462 191156 160468 191168
rect 160520 191156 160526 191208
rect 161750 191156 161756 191208
rect 161808 191196 161814 191208
rect 162026 191196 162032 191208
rect 161808 191168 162032 191196
rect 161808 191156 161814 191168
rect 162026 191156 162032 191168
rect 162084 191156 162090 191208
rect 163406 191156 163412 191208
rect 163464 191196 163470 191208
rect 163958 191196 163964 191208
rect 163464 191168 163964 191196
rect 163464 191156 163470 191168
rect 163958 191156 163964 191168
rect 164016 191156 164022 191208
rect 165706 191156 165712 191208
rect 165764 191196 165770 191208
rect 166258 191196 166264 191208
rect 165764 191168 166264 191196
rect 165764 191156 165770 191168
rect 166258 191156 166264 191168
rect 166316 191156 166322 191208
rect 166368 191196 166396 191236
rect 166902 191224 166908 191276
rect 166960 191264 166966 191276
rect 200206 191264 200212 191276
rect 166960 191236 200212 191264
rect 166960 191224 166966 191236
rect 200206 191224 200212 191236
rect 200264 191224 200270 191276
rect 206554 191196 206560 191208
rect 166368 191168 206560 191196
rect 206554 191156 206560 191168
rect 206612 191156 206618 191208
rect 207658 191156 207664 191208
rect 207716 191196 207722 191208
rect 509234 191196 509240 191208
rect 207716 191168 509240 191196
rect 207716 191156 207722 191168
rect 509234 191156 509240 191168
rect 509292 191156 509298 191208
rect 84988 191100 103514 191128
rect 84988 191088 84994 191100
rect 112254 191088 112260 191140
rect 112312 191128 112318 191140
rect 173894 191128 173900 191140
rect 112312 191100 173900 191128
rect 112312 191088 112318 191100
rect 173894 191088 173900 191100
rect 173952 191128 173958 191140
rect 174998 191128 175004 191140
rect 173952 191100 175004 191128
rect 173952 191088 173958 191100
rect 174998 191088 175004 191100
rect 175056 191088 175062 191140
rect 189994 191088 190000 191140
rect 190052 191128 190058 191140
rect 210418 191128 210424 191140
rect 190052 191100 210424 191128
rect 190052 191088 190058 191100
rect 210418 191088 210424 191100
rect 210476 191088 210482 191140
rect 216858 191088 216864 191140
rect 216916 191128 216922 191140
rect 520274 191128 520280 191140
rect 216916 191100 520280 191128
rect 216916 191088 216922 191100
rect 520274 191088 520280 191100
rect 520332 191088 520338 191140
rect 118142 191020 118148 191072
rect 118200 191060 118206 191072
rect 118200 191032 138014 191060
rect 118200 191020 118206 191032
rect 132862 190952 132868 191004
rect 132920 190992 132926 191004
rect 133598 190992 133604 191004
rect 132920 190964 133604 190992
rect 132920 190952 132926 190964
rect 133598 190952 133604 190964
rect 133656 190952 133662 191004
rect 134610 190992 134616 191004
rect 134260 190964 134616 190992
rect 134260 190936 134288 190964
rect 134610 190952 134616 190964
rect 134668 190952 134674 191004
rect 135530 190952 135536 191004
rect 135588 190992 135594 191004
rect 136082 190992 136088 191004
rect 135588 190964 136088 190992
rect 135588 190952 135594 190964
rect 136082 190952 136088 190964
rect 136140 190952 136146 191004
rect 136174 190952 136180 191004
rect 136232 190992 136238 191004
rect 136542 190992 136548 191004
rect 136232 190964 136548 190992
rect 136232 190952 136238 190964
rect 136542 190952 136548 190964
rect 136600 190952 136606 191004
rect 137186 190952 137192 191004
rect 137244 190992 137250 191004
rect 137830 190992 137836 191004
rect 137244 190964 137836 190992
rect 137244 190952 137250 190964
rect 137830 190952 137836 190964
rect 137888 190952 137894 191004
rect 137986 190992 138014 191032
rect 146570 191020 146576 191072
rect 146628 191060 146634 191072
rect 147582 191060 147588 191072
rect 146628 191032 147588 191060
rect 146628 191020 146634 191032
rect 147582 191020 147588 191032
rect 147640 191020 147646 191072
rect 148134 191020 148140 191072
rect 148192 191060 148198 191072
rect 148686 191060 148692 191072
rect 148192 191032 148692 191060
rect 148192 191020 148198 191032
rect 148686 191020 148692 191032
rect 148744 191020 148750 191072
rect 149330 191020 149336 191072
rect 149388 191060 149394 191072
rect 150250 191060 150256 191072
rect 149388 191032 150256 191060
rect 149388 191020 149394 191032
rect 150250 191020 150256 191032
rect 150308 191020 150314 191072
rect 153378 191020 153384 191072
rect 153436 191060 153442 191072
rect 154114 191060 154120 191072
rect 153436 191032 154120 191060
rect 153436 191020 153442 191032
rect 154114 191020 154120 191032
rect 154172 191020 154178 191072
rect 154666 191020 154672 191072
rect 154724 191060 154730 191072
rect 155586 191060 155592 191072
rect 154724 191032 155592 191060
rect 154724 191020 154730 191032
rect 155586 191020 155592 191032
rect 155644 191020 155650 191072
rect 156598 191020 156604 191072
rect 156656 191060 156662 191072
rect 156874 191060 156880 191072
rect 156656 191032 156880 191060
rect 156656 191020 156662 191032
rect 156874 191020 156880 191032
rect 156932 191020 156938 191072
rect 159910 191020 159916 191072
rect 159968 191060 159974 191072
rect 160094 191060 160100 191072
rect 159968 191032 160100 191060
rect 159968 191020 159974 191032
rect 160094 191020 160100 191032
rect 160152 191020 160158 191072
rect 160278 191020 160284 191072
rect 160336 191060 160342 191072
rect 160830 191060 160836 191072
rect 160336 191032 160836 191060
rect 160336 191020 160342 191032
rect 160830 191020 160836 191032
rect 160888 191020 160894 191072
rect 164510 191020 164516 191072
rect 164568 191060 164574 191072
rect 165338 191060 165344 191072
rect 164568 191032 165344 191060
rect 164568 191020 164574 191032
rect 165338 191020 165344 191032
rect 165396 191020 165402 191072
rect 197354 191060 197360 191072
rect 166966 191032 197360 191060
rect 151630 190992 151636 191004
rect 137986 190964 151636 190992
rect 151630 190952 151636 190964
rect 151688 190952 151694 191004
rect 164050 190952 164056 191004
rect 164108 190992 164114 191004
rect 166966 190992 166994 191032
rect 197354 191020 197360 191032
rect 197412 191060 197418 191072
rect 197722 191060 197728 191072
rect 197412 191032 197728 191060
rect 197412 191020 197418 191032
rect 197722 191020 197728 191032
rect 197780 191020 197786 191072
rect 164108 190964 166994 190992
rect 164108 190952 164114 190964
rect 132770 190884 132776 190936
rect 132828 190924 132834 190936
rect 133782 190924 133788 190936
rect 132828 190896 133788 190924
rect 132828 190884 132834 190896
rect 133782 190884 133788 190896
rect 133840 190884 133846 190936
rect 134242 190884 134248 190936
rect 134300 190884 134306 190936
rect 136818 190884 136824 190936
rect 136876 190924 136882 190936
rect 137554 190924 137560 190936
rect 136876 190896 137560 190924
rect 136876 190884 136882 190896
rect 137554 190884 137560 190896
rect 137612 190884 137618 190936
rect 116578 190544 116584 190596
rect 116636 190584 116642 190596
rect 162762 190584 162768 190596
rect 116636 190556 162768 190584
rect 116636 190544 116642 190556
rect 162762 190544 162768 190556
rect 162820 190544 162826 190596
rect 174170 190544 174176 190596
rect 174228 190584 174234 190596
rect 189534 190584 189540 190596
rect 174228 190556 189540 190584
rect 174228 190544 174234 190556
rect 189534 190544 189540 190556
rect 189592 190544 189598 190596
rect 4890 190476 4896 190528
rect 4948 190516 4954 190528
rect 100478 190516 100484 190528
rect 4948 190488 100484 190516
rect 4948 190476 4954 190488
rect 100478 190476 100484 190488
rect 100536 190476 100542 190528
rect 137370 190476 137376 190528
rect 137428 190516 137434 190528
rect 137922 190516 137928 190528
rect 137428 190488 137928 190516
rect 137428 190476 137434 190488
rect 137922 190476 137928 190488
rect 137980 190516 137986 190528
rect 490558 190516 490564 190528
rect 137980 190488 490564 190516
rect 137980 190476 137986 190488
rect 490558 190476 490564 190488
rect 490616 190476 490622 190528
rect 94590 190408 94596 190460
rect 94648 190448 94654 190460
rect 165614 190448 165620 190460
rect 94648 190420 165620 190448
rect 94648 190408 94654 190420
rect 165614 190408 165620 190420
rect 165672 190408 165678 190460
rect 186130 190408 186136 190460
rect 186188 190448 186194 190460
rect 563698 190448 563704 190460
rect 186188 190420 563704 190448
rect 186188 190408 186194 190420
rect 563698 190408 563704 190420
rect 563756 190408 563762 190460
rect 99098 190340 99104 190392
rect 99156 190380 99162 190392
rect 166994 190380 167000 190392
rect 99156 190352 167000 190380
rect 99156 190340 99162 190352
rect 166994 190340 167000 190352
rect 167052 190340 167058 190392
rect 170398 190340 170404 190392
rect 170456 190380 170462 190392
rect 193950 190380 193956 190392
rect 170456 190352 193956 190380
rect 170456 190340 170462 190352
rect 193950 190340 193956 190352
rect 194008 190340 194014 190392
rect 206278 190340 206284 190392
rect 206336 190380 206342 190392
rect 579982 190380 579988 190392
rect 206336 190352 579988 190380
rect 206336 190340 206342 190352
rect 579982 190340 579988 190352
rect 580040 190340 580046 190392
rect 117222 190272 117228 190324
rect 117280 190312 117286 190324
rect 173710 190312 173716 190324
rect 117280 190284 173716 190312
rect 117280 190272 117286 190284
rect 173710 190272 173716 190284
rect 173768 190272 173774 190324
rect 152274 190204 152280 190256
rect 152332 190244 152338 190256
rect 152458 190244 152464 190256
rect 152332 190216 152464 190244
rect 152332 190204 152338 190216
rect 152458 190204 152464 190216
rect 152516 190204 152522 190256
rect 177574 190204 177580 190256
rect 177632 190244 177638 190256
rect 205818 190244 205824 190256
rect 177632 190216 205824 190244
rect 177632 190204 177638 190216
rect 205818 190204 205824 190216
rect 205876 190204 205882 190256
rect 155770 190136 155776 190188
rect 155828 190176 155834 190188
rect 187786 190176 187792 190188
rect 155828 190148 187792 190176
rect 155828 190136 155834 190148
rect 187786 190136 187792 190148
rect 187844 190136 187850 190188
rect 120994 190068 121000 190120
rect 121052 190108 121058 190120
rect 148502 190108 148508 190120
rect 121052 190080 148508 190108
rect 121052 190068 121058 190080
rect 148502 190068 148508 190080
rect 148560 190068 148566 190120
rect 155862 190068 155868 190120
rect 155920 190108 155926 190120
rect 189166 190108 189172 190120
rect 155920 190080 189172 190108
rect 155920 190068 155926 190080
rect 189166 190068 189172 190080
rect 189224 190068 189230 190120
rect 109678 190000 109684 190052
rect 109736 190040 109742 190052
rect 119430 190040 119436 190052
rect 109736 190012 119436 190040
rect 109736 190000 109742 190012
rect 119430 190000 119436 190012
rect 119488 190040 119494 190052
rect 151906 190040 151912 190052
rect 119488 190012 151912 190040
rect 119488 190000 119494 190012
rect 151906 190000 151912 190012
rect 151964 190000 151970 190052
rect 163590 190000 163596 190052
rect 163648 190040 163654 190052
rect 197722 190040 197728 190052
rect 163648 190012 197728 190040
rect 163648 190000 163654 190012
rect 197722 190000 197728 190012
rect 197780 190000 197786 190052
rect 110966 189932 110972 189984
rect 111024 189972 111030 189984
rect 144362 189972 144368 189984
rect 111024 189944 144368 189972
rect 111024 189932 111030 189944
rect 144362 189932 144368 189944
rect 144420 189932 144426 189984
rect 156782 189932 156788 189984
rect 156840 189972 156846 189984
rect 190822 189972 190828 189984
rect 156840 189944 190828 189972
rect 156840 189932 156846 189944
rect 190822 189932 190828 189944
rect 190880 189932 190886 189984
rect 110874 189864 110880 189916
rect 110932 189904 110938 189916
rect 145834 189904 145840 189916
rect 110932 189876 145840 189904
rect 110932 189864 110938 189876
rect 145834 189864 145840 189876
rect 145892 189864 145898 189916
rect 158346 189864 158352 189916
rect 158404 189904 158410 189916
rect 217226 189904 217232 189916
rect 158404 189876 217232 189904
rect 158404 189864 158410 189876
rect 217226 189864 217232 189876
rect 217284 189904 217290 189916
rect 572070 189904 572076 189916
rect 217284 189876 572076 189904
rect 217284 189864 217290 189876
rect 572070 189864 572076 189876
rect 572128 189864 572134 189916
rect 95970 189796 95976 189848
rect 96028 189836 96034 189848
rect 109494 189836 109500 189848
rect 96028 189808 109500 189836
rect 96028 189796 96034 189808
rect 109494 189796 109500 189808
rect 109552 189836 109558 189848
rect 144546 189836 144552 189848
rect 109552 189808 144552 189836
rect 109552 189796 109558 189808
rect 144546 189796 144552 189808
rect 144604 189796 144610 189848
rect 158070 189796 158076 189848
rect 158128 189836 158134 189848
rect 192386 189836 192392 189848
rect 158128 189808 192392 189836
rect 158128 189796 158134 189808
rect 192386 189796 192392 189808
rect 192444 189796 192450 189848
rect 207750 189796 207756 189848
rect 207808 189836 207814 189848
rect 569218 189836 569224 189848
rect 207808 189808 569224 189836
rect 207808 189796 207814 189808
rect 569218 189796 569224 189808
rect 569276 189796 569282 189848
rect 90358 189728 90364 189780
rect 90416 189768 90422 189780
rect 97074 189768 97080 189780
rect 90416 189740 97080 189768
rect 90416 189728 90422 189740
rect 97074 189728 97080 189740
rect 97132 189768 97138 189780
rect 155126 189768 155132 189780
rect 97132 189740 155132 189768
rect 97132 189728 97138 189740
rect 155126 189728 155132 189740
rect 155184 189728 155190 189780
rect 159266 189728 159272 189780
rect 159324 189768 159330 189780
rect 183370 189768 183376 189780
rect 159324 189740 183376 189768
rect 159324 189728 159330 189740
rect 183370 189728 183376 189740
rect 183428 189768 183434 189780
rect 563882 189768 563888 189780
rect 183428 189740 563888 189768
rect 183428 189728 183434 189740
rect 563882 189728 563888 189740
rect 563940 189728 563946 189780
rect 163866 189660 163872 189712
rect 163924 189700 163930 189712
rect 191926 189700 191932 189712
rect 163924 189672 191932 189700
rect 163924 189660 163930 189672
rect 191926 189660 191932 189672
rect 191984 189660 191990 189712
rect 154850 189592 154856 189644
rect 154908 189632 154914 189644
rect 155218 189632 155224 189644
rect 154908 189604 155224 189632
rect 154908 189592 154914 189604
rect 155218 189592 155224 189604
rect 155276 189592 155282 189644
rect 166994 189116 167000 189168
rect 167052 189156 167058 189168
rect 167362 189156 167368 189168
rect 167052 189128 167368 189156
rect 167052 189116 167058 189128
rect 167362 189116 167368 189128
rect 167420 189116 167426 189168
rect 108022 189048 108028 189100
rect 108080 189088 108086 189100
rect 108080 189060 142844 189088
rect 108080 189048 108086 189060
rect 142816 189020 142844 189060
rect 149624 189060 150296 189088
rect 149624 189020 149652 189060
rect 142816 188992 149652 189020
rect 149698 188980 149704 189032
rect 149756 189020 149762 189032
rect 150158 189020 150164 189032
rect 149756 188992 150164 189020
rect 149756 188980 149762 188992
rect 150158 188980 150164 188992
rect 150216 188980 150222 189032
rect 150268 189020 150296 189060
rect 165614 189048 165620 189100
rect 165672 189088 165678 189100
rect 167086 189088 167092 189100
rect 165672 189060 167092 189088
rect 165672 189048 165678 189060
rect 167086 189048 167092 189060
rect 167144 189048 167150 189100
rect 152090 189020 152096 189032
rect 150268 188992 152096 189020
rect 152090 188980 152096 188992
rect 152148 189020 152154 189032
rect 566734 189020 566740 189032
rect 152148 188992 566740 189020
rect 152148 188980 152154 188992
rect 566734 188980 566740 188992
rect 566792 188980 566798 189032
rect 106182 188912 106188 188964
rect 106240 188952 106246 188964
rect 152182 188952 152188 188964
rect 106240 188924 152188 188952
rect 106240 188912 106246 188924
rect 152182 188912 152188 188924
rect 152240 188912 152246 188964
rect 172606 188844 172612 188896
rect 172664 188884 172670 188896
rect 207382 188884 207388 188896
rect 172664 188856 207388 188884
rect 172664 188844 172670 188856
rect 207382 188844 207388 188856
rect 207440 188884 207446 188896
rect 207750 188884 207756 188896
rect 207440 188856 207756 188884
rect 207440 188844 207446 188856
rect 207750 188844 207756 188856
rect 207808 188844 207814 188896
rect 158530 188776 158536 188828
rect 158588 188816 158594 188828
rect 201494 188816 201500 188828
rect 158588 188788 201500 188816
rect 158588 188776 158594 188788
rect 201494 188776 201500 188788
rect 201552 188776 201558 188828
rect 128998 188708 129004 188760
rect 129056 188748 129062 188760
rect 153930 188748 153936 188760
rect 129056 188720 153936 188748
rect 129056 188708 129062 188720
rect 153930 188708 153936 188720
rect 153988 188748 153994 188760
rect 251174 188748 251180 188760
rect 153988 188720 251180 188748
rect 153988 188708 153994 188720
rect 251174 188708 251180 188720
rect 251232 188708 251238 188760
rect 93210 188640 93216 188692
rect 93268 188680 93274 188692
rect 173526 188680 173532 188692
rect 93268 188652 173532 188680
rect 93268 188640 93274 188652
rect 173526 188640 173532 188652
rect 173584 188680 173590 188692
rect 206094 188680 206100 188692
rect 173584 188652 206100 188680
rect 173584 188640 173590 188652
rect 206094 188640 206100 188652
rect 206152 188640 206158 188692
rect 106274 188572 106280 188624
rect 106332 188612 106338 188624
rect 176930 188612 176936 188624
rect 106332 188584 176936 188612
rect 106332 188572 106338 188584
rect 176930 188572 176936 188584
rect 176988 188612 176994 188624
rect 210142 188612 210148 188624
rect 176988 188584 210148 188612
rect 176988 188572 176994 188584
rect 210142 188572 210148 188584
rect 210200 188572 210206 188624
rect 95970 188504 95976 188556
rect 96028 188544 96034 188556
rect 104894 188544 104900 188556
rect 96028 188516 104900 188544
rect 96028 188504 96034 188516
rect 104894 188504 104900 188516
rect 104952 188544 104958 188556
rect 106182 188544 106188 188556
rect 104952 188516 106188 188544
rect 104952 188504 104958 188516
rect 106182 188504 106188 188516
rect 106240 188504 106246 188556
rect 108482 188504 108488 188556
rect 108540 188544 108546 188556
rect 178218 188544 178224 188556
rect 108540 188516 178224 188544
rect 108540 188504 108546 188516
rect 178218 188504 178224 188516
rect 178276 188544 178282 188556
rect 178276 188516 180794 188544
rect 178276 188504 178282 188516
rect 103054 188436 103060 188488
rect 103112 188476 103118 188488
rect 104618 188476 104624 188488
rect 103112 188448 104624 188476
rect 103112 188436 103118 188448
rect 104618 188436 104624 188448
rect 104676 188476 104682 188488
rect 137094 188476 137100 188488
rect 104676 188448 137100 188476
rect 104676 188436 104682 188448
rect 137094 188436 137100 188448
rect 137152 188436 137158 188488
rect 180766 188476 180794 188516
rect 215754 188476 215760 188488
rect 180766 188448 215760 188476
rect 215754 188436 215760 188448
rect 215812 188436 215818 188488
rect 101674 188368 101680 188420
rect 101732 188408 101738 188420
rect 111518 188408 111524 188420
rect 101732 188380 111524 188408
rect 101732 188368 101738 188380
rect 111518 188368 111524 188380
rect 111576 188408 111582 188420
rect 144638 188408 144644 188420
rect 111576 188380 144644 188408
rect 111576 188368 111582 188380
rect 144638 188368 144644 188380
rect 144696 188368 144702 188420
rect 166994 188368 167000 188420
rect 167052 188408 167058 188420
rect 167454 188408 167460 188420
rect 167052 188380 167460 188408
rect 167052 188368 167058 188380
rect 167454 188368 167460 188380
rect 167512 188408 167518 188420
rect 216950 188408 216956 188420
rect 167512 188380 216956 188408
rect 167512 188368 167518 188380
rect 216950 188368 216956 188380
rect 217008 188368 217014 188420
rect 27614 188300 27620 188352
rect 27672 188340 27678 188352
rect 99742 188340 99748 188352
rect 27672 188312 99748 188340
rect 27672 188300 27678 188312
rect 99742 188300 99748 188312
rect 99800 188340 99806 188352
rect 132586 188340 132592 188352
rect 99800 188312 132592 188340
rect 99800 188300 99806 188312
rect 132586 188300 132592 188312
rect 132644 188300 132650 188352
rect 154298 188300 154304 188352
rect 154356 188340 154362 188352
rect 218422 188340 218428 188352
rect 154356 188312 218428 188340
rect 154356 188300 154362 188312
rect 218422 188300 218428 188312
rect 218480 188340 218486 188352
rect 563974 188340 563980 188352
rect 218480 188312 563980 188340
rect 218480 188300 218486 188312
rect 563974 188300 563980 188312
rect 564032 188300 564038 188352
rect 101582 188232 101588 188284
rect 101640 188272 101646 188284
rect 166626 188272 166632 188284
rect 101640 188244 166632 188272
rect 101640 188232 101646 188244
rect 166626 188232 166632 188244
rect 166684 188272 166690 188284
rect 207290 188272 207296 188284
rect 166684 188244 166994 188272
rect 166684 188232 166690 188244
rect 166966 188204 166994 188244
rect 180766 188244 207296 188272
rect 180242 188204 180248 188216
rect 166966 188176 180248 188204
rect 180242 188164 180248 188176
rect 180300 188164 180306 188216
rect 49694 188096 49700 188148
rect 49752 188136 49758 188148
rect 166994 188136 167000 188148
rect 49752 188108 167000 188136
rect 49752 188096 49758 188108
rect 166994 188096 167000 188108
rect 167052 188096 167058 188148
rect 3234 188028 3240 188080
rect 3292 188068 3298 188080
rect 175734 188068 175740 188080
rect 3292 188040 175740 188068
rect 3292 188028 3298 188040
rect 175734 188028 175740 188040
rect 175792 188068 175798 188080
rect 180766 188068 180794 188244
rect 207290 188232 207296 188244
rect 207348 188232 207354 188284
rect 175792 188040 180794 188068
rect 175792 188028 175798 188040
rect 149698 187960 149704 188012
rect 149756 188000 149762 188012
rect 471974 188000 471980 188012
rect 149756 187972 471980 188000
rect 149756 187960 149762 187972
rect 471974 187960 471980 187972
rect 472032 187960 472038 188012
rect 130746 187824 130752 187876
rect 130804 187864 130810 187876
rect 148226 187864 148232 187876
rect 130804 187836 148232 187864
rect 130804 187824 130810 187836
rect 148226 187824 148232 187836
rect 148284 187864 148290 187876
rect 148962 187864 148968 187876
rect 148284 187836 148968 187864
rect 148284 187824 148290 187836
rect 148962 187824 148968 187836
rect 149020 187824 149026 187876
rect 124858 187756 124864 187808
rect 124916 187796 124922 187808
rect 124916 187768 144960 187796
rect 124916 187756 124922 187768
rect 109770 187688 109776 187740
rect 109828 187728 109834 187740
rect 109828 187700 142844 187728
rect 109828 187688 109834 187700
rect 142816 187592 142844 187700
rect 144932 187660 144960 187768
rect 201494 187688 201500 187740
rect 201552 187728 201558 187740
rect 207106 187728 207112 187740
rect 201552 187700 207112 187728
rect 201552 187688 201558 187700
rect 207106 187688 207112 187700
rect 207164 187688 207170 187740
rect 145558 187660 145564 187672
rect 144932 187632 145564 187660
rect 145558 187620 145564 187632
rect 145616 187660 145622 187672
rect 579062 187660 579068 187672
rect 145616 187632 579068 187660
rect 145616 187620 145622 187632
rect 579062 187620 579068 187632
rect 579120 187620 579126 187672
rect 150342 187592 150348 187604
rect 142816 187564 150348 187592
rect 150342 187552 150348 187564
rect 150400 187592 150406 187604
rect 569310 187592 569316 187604
rect 150400 187564 569316 187592
rect 150400 187552 150406 187564
rect 569310 187552 569316 187564
rect 569368 187552 569374 187604
rect 90634 187484 90640 187536
rect 90692 187524 90698 187536
rect 177298 187524 177304 187536
rect 90692 187496 177304 187524
rect 90692 187484 90698 187496
rect 177298 187484 177304 187496
rect 177356 187484 177362 187536
rect 177390 187484 177396 187536
rect 177448 187524 177454 187536
rect 177942 187524 177948 187536
rect 177448 187496 177948 187524
rect 177448 187484 177454 187496
rect 177942 187484 177948 187496
rect 178000 187524 178006 187536
rect 313918 187524 313924 187536
rect 178000 187496 313924 187524
rect 178000 187484 178006 187496
rect 313918 187484 313924 187496
rect 313976 187484 313982 187536
rect 96154 187416 96160 187468
rect 96212 187456 96218 187468
rect 174170 187456 174176 187468
rect 96212 187428 174176 187456
rect 96212 187416 96218 187428
rect 174170 187416 174176 187428
rect 174228 187416 174234 187468
rect 110138 187348 110144 187400
rect 110196 187388 110202 187400
rect 142706 187388 142712 187400
rect 110196 187360 142712 187388
rect 110196 187348 110202 187360
rect 142706 187348 142712 187360
rect 142764 187348 142770 187400
rect 168834 187348 168840 187400
rect 168892 187388 168898 187400
rect 203058 187388 203064 187400
rect 168892 187360 203064 187388
rect 168892 187348 168898 187360
rect 203058 187348 203064 187360
rect 203116 187348 203122 187400
rect 110046 187280 110052 187332
rect 110104 187320 110110 187332
rect 143350 187320 143356 187332
rect 110104 187292 143356 187320
rect 110104 187280 110110 187292
rect 143350 187280 143356 187292
rect 143408 187280 143414 187332
rect 165246 187280 165252 187332
rect 165304 187320 165310 187332
rect 199378 187320 199384 187332
rect 165304 187292 199384 187320
rect 165304 187280 165310 187292
rect 199378 187280 199384 187292
rect 199436 187280 199442 187332
rect 99650 187212 99656 187264
rect 99708 187252 99714 187264
rect 133414 187252 133420 187264
rect 99708 187224 133420 187252
rect 99708 187212 99714 187224
rect 133414 187212 133420 187224
rect 133472 187212 133478 187264
rect 155954 187212 155960 187264
rect 156012 187252 156018 187264
rect 156322 187252 156328 187264
rect 156012 187224 156328 187252
rect 156012 187212 156018 187224
rect 156322 187212 156328 187224
rect 156380 187252 156386 187264
rect 170398 187252 170404 187264
rect 156380 187224 170404 187252
rect 156380 187212 156386 187224
rect 170398 187212 170404 187224
rect 170456 187212 170462 187264
rect 175642 187212 175648 187264
rect 175700 187252 175706 187264
rect 210234 187252 210240 187264
rect 175700 187224 210240 187252
rect 175700 187212 175706 187224
rect 210234 187212 210240 187224
rect 210292 187212 210298 187264
rect 112438 187144 112444 187196
rect 112496 187184 112502 187196
rect 144914 187184 144920 187196
rect 112496 187156 144920 187184
rect 112496 187144 112502 187156
rect 144914 187144 144920 187156
rect 144972 187144 144978 187196
rect 164970 187144 164976 187196
rect 165028 187184 165034 187196
rect 199286 187184 199292 187196
rect 165028 187156 199292 187184
rect 165028 187144 165034 187156
rect 199286 187144 199292 187156
rect 199344 187144 199350 187196
rect 109954 187076 109960 187128
rect 110012 187116 110018 187128
rect 143718 187116 143724 187128
rect 110012 187088 143724 187116
rect 110012 187076 110018 187088
rect 143718 187076 143724 187088
rect 143776 187076 143782 187128
rect 167178 187076 167184 187128
rect 167236 187116 167242 187128
rect 201954 187116 201960 187128
rect 167236 187088 201960 187116
rect 167236 187076 167242 187088
rect 201954 187076 201960 187088
rect 202012 187076 202018 187128
rect 113726 187008 113732 187060
rect 113784 187048 113790 187060
rect 148410 187048 148416 187060
rect 113784 187020 148416 187048
rect 113784 187008 113790 187020
rect 148410 187008 148416 187020
rect 148468 187008 148474 187060
rect 170306 187008 170312 187060
rect 170364 187048 170370 187060
rect 204806 187048 204812 187060
rect 170364 187020 204812 187048
rect 170364 187008 170370 187020
rect 204806 187008 204812 187020
rect 204864 187048 204870 187060
rect 204864 187020 209774 187048
rect 204864 187008 204870 187020
rect 96062 186940 96068 186992
rect 96120 186980 96126 186992
rect 121086 186980 121092 186992
rect 96120 186952 121092 186980
rect 96120 186940 96126 186952
rect 121086 186940 121092 186952
rect 121144 186980 121150 186992
rect 157150 186980 157156 186992
rect 121144 186952 157156 186980
rect 121144 186940 121150 186952
rect 157150 186940 157156 186952
rect 157208 186940 157214 186992
rect 158162 186940 158168 186992
rect 158220 186980 158226 186992
rect 193858 186980 193864 186992
rect 158220 186952 193864 186980
rect 158220 186940 158226 186952
rect 193858 186940 193864 186952
rect 193916 186940 193922 186992
rect 209746 186980 209774 187020
rect 572162 186980 572168 186992
rect 209746 186952 572168 186980
rect 572162 186940 572168 186952
rect 572220 186940 572226 186992
rect 115474 186872 115480 186924
rect 115532 186912 115538 186924
rect 147306 186912 147312 186924
rect 115532 186884 147312 186912
rect 115532 186872 115538 186884
rect 147306 186872 147312 186884
rect 147364 186872 147370 186924
rect 167270 186872 167276 186924
rect 167328 186912 167334 186924
rect 201494 186912 201500 186924
rect 167328 186884 201500 186912
rect 167328 186872 167334 186884
rect 201494 186872 201500 186884
rect 201552 186872 201558 186924
rect 106090 186804 106096 186856
rect 106148 186844 106154 186856
rect 136358 186844 136364 186856
rect 106148 186816 136364 186844
rect 106148 186804 106154 186816
rect 136358 186804 136364 186816
rect 136416 186804 136422 186856
rect 161934 186804 161940 186856
rect 161992 186844 161998 186856
rect 195974 186844 195980 186856
rect 161992 186816 195980 186844
rect 161992 186804 161998 186816
rect 195974 186804 195980 186816
rect 196032 186804 196038 186856
rect 97442 186736 97448 186788
rect 97500 186776 97506 186788
rect 155954 186776 155960 186788
rect 97500 186748 155960 186776
rect 97500 186736 97506 186748
rect 155954 186736 155960 186748
rect 156012 186736 156018 186788
rect 170766 186736 170772 186788
rect 170824 186776 170830 186788
rect 202966 186776 202972 186788
rect 170824 186748 202972 186776
rect 170824 186736 170830 186748
rect 202966 186736 202972 186748
rect 203024 186736 203030 186788
rect 108298 186668 108304 186720
rect 108356 186708 108362 186720
rect 154574 186708 154580 186720
rect 108356 186680 154580 186708
rect 108356 186668 108362 186680
rect 154574 186668 154580 186680
rect 154632 186708 154638 186720
rect 166258 186708 166264 186720
rect 154632 186680 166264 186708
rect 154632 186668 154638 186680
rect 166258 186668 166264 186680
rect 166316 186668 166322 186720
rect 107102 186328 107108 186380
rect 107160 186368 107166 186380
rect 129734 186368 129740 186380
rect 107160 186340 129740 186368
rect 107160 186328 107166 186340
rect 129734 186328 129740 186340
rect 129792 186328 129798 186380
rect 8294 186260 8300 186312
rect 8352 186300 8358 186312
rect 176746 186300 176752 186312
rect 8352 186272 176752 186300
rect 8352 186260 8358 186272
rect 176746 186260 176752 186272
rect 176804 186260 176810 186312
rect 30374 186192 30380 186244
rect 30432 186232 30438 186244
rect 178126 186232 178132 186244
rect 30432 186204 178132 186232
rect 30432 186192 30438 186204
rect 178126 186192 178132 186204
rect 178184 186192 178190 186244
rect 129734 186124 129740 186176
rect 129792 186164 129798 186176
rect 143442 186164 143448 186176
rect 129792 186136 143448 186164
rect 129792 186124 129798 186136
rect 143442 186124 143448 186136
rect 143500 186164 143506 186176
rect 273254 186164 273260 186176
rect 143500 186136 273260 186164
rect 143500 186124 143506 186136
rect 273254 186124 273260 186136
rect 273312 186124 273318 186176
rect 93394 186056 93400 186108
rect 93452 186096 93458 186108
rect 175550 186096 175556 186108
rect 93452 186068 175556 186096
rect 93452 186056 93458 186068
rect 175550 186056 175556 186068
rect 175608 186096 175614 186108
rect 210050 186096 210056 186108
rect 175608 186068 210056 186096
rect 175608 186056 175614 186068
rect 210050 186056 210056 186068
rect 210108 186056 210114 186108
rect 100202 185988 100208 186040
rect 100260 186028 100266 186040
rect 180794 186028 180800 186040
rect 100260 186000 180800 186028
rect 100260 185988 100266 186000
rect 180794 185988 180800 186000
rect 180852 186028 180858 186040
rect 210510 186028 210516 186040
rect 180852 186000 210516 186028
rect 180852 185988 180858 186000
rect 210510 185988 210516 186000
rect 210568 185988 210574 186040
rect 103146 185920 103152 185972
rect 103204 185960 103210 185972
rect 176654 185960 176660 185972
rect 103204 185932 176660 185960
rect 103204 185920 103210 185932
rect 176654 185920 176660 185932
rect 176712 185920 176718 185972
rect 178126 185920 178132 185972
rect 178184 185960 178190 185972
rect 208670 185960 208676 185972
rect 178184 185932 208676 185960
rect 178184 185920 178190 185932
rect 208670 185920 208676 185932
rect 208728 185920 208734 185972
rect 87598 185852 87604 185904
rect 87656 185892 87662 185904
rect 107378 185892 107384 185904
rect 87656 185864 107384 185892
rect 87656 185852 87662 185864
rect 107378 185852 107384 185864
rect 107436 185852 107442 185904
rect 127894 185852 127900 185904
rect 127952 185892 127958 185904
rect 132954 185892 132960 185904
rect 127952 185864 132960 185892
rect 127952 185852 127958 185864
rect 132954 185852 132960 185864
rect 133012 185892 133018 185904
rect 205634 185892 205640 185904
rect 133012 185864 205640 185892
rect 133012 185852 133018 185864
rect 205634 185852 205640 185864
rect 205692 185852 205698 185904
rect 97534 185784 97540 185836
rect 97592 185824 97598 185836
rect 168374 185824 168380 185836
rect 97592 185796 168380 185824
rect 97592 185784 97598 185796
rect 168374 185784 168380 185796
rect 168432 185784 168438 185836
rect 176654 185784 176660 185836
rect 176712 185824 176718 185836
rect 211706 185824 211712 185836
rect 176712 185796 211712 185824
rect 176712 185784 176718 185796
rect 211706 185784 211712 185796
rect 211764 185784 211770 185836
rect 100110 185716 100116 185768
rect 100168 185756 100174 185768
rect 170214 185756 170220 185768
rect 100168 185728 170220 185756
rect 100168 185716 100174 185728
rect 170214 185716 170220 185728
rect 170272 185756 170278 185768
rect 212810 185756 212816 185768
rect 170272 185728 212816 185756
rect 170272 185716 170278 185728
rect 212810 185716 212816 185728
rect 212868 185716 212874 185768
rect 218146 185716 218152 185768
rect 218204 185756 218210 185768
rect 218330 185756 218336 185768
rect 218204 185728 218336 185756
rect 218204 185716 218210 185728
rect 218330 185716 218336 185728
rect 218388 185756 218394 185768
rect 240134 185756 240140 185768
rect 218388 185728 240140 185756
rect 218388 185716 218394 185728
rect 240134 185716 240140 185728
rect 240192 185716 240198 185768
rect 98914 185648 98920 185700
rect 98972 185688 98978 185700
rect 103054 185688 103060 185700
rect 98972 185660 103060 185688
rect 98972 185648 98978 185660
rect 103054 185648 103060 185660
rect 103112 185688 103118 185700
rect 135530 185688 135536 185700
rect 103112 185660 135536 185688
rect 103112 185648 103118 185660
rect 135530 185648 135536 185660
rect 135588 185648 135594 185700
rect 158898 185648 158904 185700
rect 158956 185688 158962 185700
rect 158956 185660 219434 185688
rect 158956 185648 158962 185660
rect 100294 185580 100300 185632
rect 100352 185620 100358 185632
rect 135162 185620 135168 185632
rect 100352 185592 135168 185620
rect 100352 185580 100358 185592
rect 135162 185580 135168 185592
rect 135220 185580 135226 185632
rect 155034 185580 155040 185632
rect 155092 185620 155098 185632
rect 218146 185620 218152 185632
rect 155092 185592 218152 185620
rect 155092 185580 155098 185592
rect 218146 185580 218152 185592
rect 218204 185580 218210 185632
rect 219406 185620 219434 185660
rect 220998 185620 221004 185632
rect 219406 185592 221004 185620
rect 220998 185580 221004 185592
rect 221056 185620 221062 185632
rect 581638 185620 581644 185632
rect 221056 185592 581644 185620
rect 221056 185580 221062 185592
rect 581638 185580 581644 185592
rect 581696 185580 581702 185632
rect 107194 185512 107200 185564
rect 107252 185552 107258 185564
rect 107378 185552 107384 185564
rect 107252 185524 107384 185552
rect 107252 185512 107258 185524
rect 107378 185512 107384 185524
rect 107436 185552 107442 185564
rect 136266 185552 136272 185564
rect 107436 185524 136272 185552
rect 107436 185512 107442 185524
rect 136266 185512 136272 185524
rect 136324 185512 136330 185564
rect 161842 185512 161848 185564
rect 161900 185552 161906 185564
rect 184290 185552 184296 185564
rect 161900 185524 184296 185552
rect 161900 185512 161906 185524
rect 184290 185512 184296 185524
rect 184348 185552 184354 185564
rect 184842 185552 184848 185564
rect 184348 185524 184848 185552
rect 184348 185512 184354 185524
rect 184842 185512 184848 185524
rect 184900 185512 184906 185564
rect 161750 185444 161756 185496
rect 161808 185484 161814 185496
rect 181898 185484 181904 185496
rect 161808 185456 181904 185484
rect 161808 185444 161814 185456
rect 181898 185444 181904 185456
rect 181956 185444 181962 185496
rect 218146 185444 218152 185496
rect 218204 185484 218210 185496
rect 218422 185484 218428 185496
rect 218204 185456 218428 185484
rect 218204 185444 218210 185456
rect 218422 185444 218428 185456
rect 218480 185444 218486 185496
rect 168374 184968 168380 185020
rect 168432 185008 168438 185020
rect 207474 185008 207480 185020
rect 168432 184980 207480 185008
rect 168432 184968 168438 184980
rect 207474 184968 207480 184980
rect 207532 184968 207538 185020
rect 181898 184900 181904 184952
rect 181956 184940 181962 184952
rect 580166 184940 580172 184952
rect 181956 184912 580172 184940
rect 181956 184900 181962 184912
rect 580166 184900 580172 184912
rect 580224 184900 580230 184952
rect 131114 184832 131120 184884
rect 131172 184872 131178 184884
rect 145374 184872 145380 184884
rect 131172 184844 145380 184872
rect 131172 184832 131178 184844
rect 145374 184832 145380 184844
rect 145432 184872 145438 184884
rect 418154 184872 418160 184884
rect 145432 184844 418160 184872
rect 145432 184832 145438 184844
rect 418154 184832 418160 184844
rect 418212 184832 418218 184884
rect 90450 184764 90456 184816
rect 90508 184804 90514 184816
rect 177298 184804 177304 184816
rect 90508 184776 177304 184804
rect 90508 184764 90514 184776
rect 177298 184764 177304 184776
rect 177356 184804 177362 184816
rect 177758 184804 177764 184816
rect 177356 184776 177764 184804
rect 177356 184764 177362 184776
rect 177758 184764 177764 184776
rect 177816 184764 177822 184816
rect 90542 184696 90548 184748
rect 90600 184736 90606 184748
rect 164510 184736 164516 184748
rect 90600 184708 164516 184736
rect 90600 184696 90606 184708
rect 164510 184696 164516 184708
rect 164568 184736 164574 184748
rect 165522 184736 165528 184748
rect 164568 184708 165528 184736
rect 164568 184696 164574 184708
rect 165522 184696 165528 184708
rect 165580 184696 165586 184748
rect 167086 184696 167092 184748
rect 167144 184736 167150 184748
rect 200482 184736 200488 184748
rect 167144 184708 200488 184736
rect 167144 184696 167150 184708
rect 200482 184696 200488 184708
rect 200540 184696 200546 184748
rect 97258 184628 97264 184680
rect 97316 184668 97322 184680
rect 168742 184668 168748 184680
rect 97316 184640 168748 184668
rect 97316 184628 97322 184640
rect 168742 184628 168748 184640
rect 168800 184628 168806 184680
rect 173710 184628 173716 184680
rect 173768 184668 173774 184680
rect 204898 184668 204904 184680
rect 173768 184640 204904 184668
rect 173768 184628 173774 184640
rect 204898 184628 204904 184640
rect 204956 184628 204962 184680
rect 104342 184560 104348 184612
rect 104400 184600 104406 184612
rect 134610 184600 134616 184612
rect 104400 184572 134616 184600
rect 104400 184560 104406 184572
rect 134610 184560 134616 184572
rect 134668 184560 134674 184612
rect 167362 184560 167368 184612
rect 167420 184600 167426 184612
rect 201862 184600 201868 184612
rect 167420 184572 201868 184600
rect 167420 184560 167426 184572
rect 201862 184560 201868 184572
rect 201920 184560 201926 184612
rect 108574 184492 108580 184544
rect 108632 184532 108638 184544
rect 139762 184532 139768 184544
rect 108632 184504 139768 184532
rect 108632 184492 108638 184504
rect 139762 184492 139768 184504
rect 139820 184492 139826 184544
rect 171410 184492 171416 184544
rect 171468 184532 171474 184544
rect 205910 184532 205916 184544
rect 171468 184504 205916 184532
rect 171468 184492 171474 184504
rect 205910 184492 205916 184504
rect 205968 184492 205974 184544
rect 101306 184424 101312 184476
rect 101364 184464 101370 184476
rect 134242 184464 134248 184476
rect 101364 184436 134248 184464
rect 101364 184424 101370 184436
rect 134242 184424 134248 184436
rect 134300 184424 134306 184476
rect 171318 184424 171324 184476
rect 171376 184464 171382 184476
rect 206002 184464 206008 184476
rect 171376 184436 206008 184464
rect 171376 184424 171382 184436
rect 206002 184424 206008 184436
rect 206060 184424 206066 184476
rect 106182 184356 106188 184408
rect 106240 184396 106246 184408
rect 140498 184396 140504 184408
rect 106240 184368 140504 184396
rect 106240 184356 106246 184368
rect 140498 184356 140504 184368
rect 140556 184356 140562 184408
rect 169846 184356 169852 184408
rect 169904 184396 169910 184408
rect 204714 184396 204720 184408
rect 169904 184368 204720 184396
rect 169904 184356 169910 184368
rect 204714 184356 204720 184368
rect 204772 184356 204778 184408
rect 109678 184288 109684 184340
rect 109736 184328 109742 184340
rect 144454 184328 144460 184340
rect 109736 184300 144460 184328
rect 109736 184288 109742 184300
rect 144454 184288 144460 184300
rect 144512 184288 144518 184340
rect 171042 184288 171048 184340
rect 171100 184328 171106 184340
rect 206278 184328 206284 184340
rect 171100 184300 206284 184328
rect 171100 184288 171106 184300
rect 206278 184288 206284 184300
rect 206336 184288 206342 184340
rect 104434 184220 104440 184272
rect 104492 184260 104498 184272
rect 138290 184260 138296 184272
rect 104492 184232 138296 184260
rect 104492 184220 104498 184232
rect 138290 184220 138296 184232
rect 138348 184220 138354 184272
rect 165522 184220 165528 184272
rect 165580 184260 165586 184272
rect 206370 184260 206376 184272
rect 165580 184232 206376 184260
rect 165580 184220 165586 184232
rect 206370 184220 206376 184232
rect 206428 184220 206434 184272
rect 3142 184152 3148 184204
rect 3200 184192 3206 184204
rect 171962 184192 171968 184204
rect 3200 184164 171968 184192
rect 3200 184152 3206 184164
rect 171962 184152 171968 184164
rect 172020 184152 172026 184204
rect 174078 184152 174084 184204
rect 174136 184192 174142 184204
rect 208578 184192 208584 184204
rect 174136 184164 208584 184192
rect 174136 184152 174142 184164
rect 208578 184152 208584 184164
rect 208636 184152 208642 184204
rect 103238 184084 103244 184136
rect 103296 184124 103302 184136
rect 132218 184124 132224 184136
rect 103296 184096 132224 184124
rect 103296 184084 103302 184096
rect 132218 184084 132224 184096
rect 132276 184084 132282 184136
rect 107378 184016 107384 184068
rect 107436 184056 107442 184068
rect 132126 184056 132132 184068
rect 107436 184028 132132 184056
rect 107436 184016 107442 184028
rect 132126 184016 132132 184028
rect 132184 184016 132190 184068
rect 97350 183948 97356 184000
rect 97408 183988 97414 184000
rect 110414 183988 110420 184000
rect 97408 183960 110420 183988
rect 97408 183948 97414 183960
rect 110414 183948 110420 183960
rect 110472 183948 110478 184000
rect 102962 183880 102968 183932
rect 103020 183920 103026 183932
rect 132862 183920 132868 183932
rect 103020 183892 132868 183920
rect 103020 183880 103026 183892
rect 132862 183880 132868 183892
rect 132920 183880 132926 183932
rect 100018 183472 100024 183524
rect 100076 183512 100082 183524
rect 182266 183512 182272 183524
rect 100076 183484 182272 183512
rect 100076 183472 100082 183484
rect 182266 183472 182272 183484
rect 182324 183512 182330 183524
rect 182324 183484 190454 183512
rect 182324 183472 182330 183484
rect 103514 183404 103520 183456
rect 103572 183444 103578 183456
rect 103572 183416 180794 183444
rect 103572 183404 103578 183416
rect 84838 183336 84844 183388
rect 84896 183376 84902 183388
rect 160002 183376 160008 183388
rect 84896 183348 160008 183376
rect 84896 183336 84902 183348
rect 160002 183336 160008 183348
rect 160060 183376 160066 183388
rect 160060 183348 161474 183376
rect 160060 183336 160066 183348
rect 107286 183268 107292 183320
rect 107344 183308 107350 183320
rect 108298 183308 108304 183320
rect 107344 183280 108304 183308
rect 107344 183268 107350 183280
rect 108298 183268 108304 183280
rect 108356 183268 108362 183320
rect 110414 183268 110420 183320
rect 110472 183308 110478 183320
rect 111058 183308 111064 183320
rect 110472 183280 111064 183308
rect 110472 183268 110478 183280
rect 111058 183268 111064 183280
rect 111116 183308 111122 183320
rect 142890 183308 142896 183320
rect 111116 183280 142896 183308
rect 111116 183268 111122 183280
rect 142890 183268 142896 183280
rect 142948 183268 142954 183320
rect 104986 183200 104992 183252
rect 105044 183240 105050 183252
rect 105814 183240 105820 183252
rect 105044 183212 105820 183240
rect 105044 183200 105050 183212
rect 105814 183200 105820 183212
rect 105872 183240 105878 183252
rect 135806 183240 135812 183252
rect 105872 183212 135812 183240
rect 105872 183200 105878 183212
rect 135806 183200 135812 183212
rect 135864 183200 135870 183252
rect 161446 183240 161474 183348
rect 180766 183308 180794 183416
rect 190426 183376 190454 183484
rect 208762 183376 208768 183388
rect 190426 183348 208768 183376
rect 208762 183336 208768 183348
rect 208820 183336 208826 183388
rect 182174 183308 182180 183320
rect 180766 183280 182180 183308
rect 182174 183268 182180 183280
rect 182232 183308 182238 183320
rect 212626 183308 212632 183320
rect 182232 183280 212632 183308
rect 182232 183268 182238 183280
rect 212626 183268 212632 183280
rect 212684 183268 212690 183320
rect 209774 183240 209780 183252
rect 161446 183212 209780 183240
rect 209774 183200 209780 183212
rect 209832 183200 209838 183252
rect 158346 183132 158352 183184
rect 158404 183172 158410 183184
rect 211338 183172 211344 183184
rect 158404 183144 211344 183172
rect 158404 183132 158410 183144
rect 211338 183132 211344 183144
rect 211396 183172 211402 183184
rect 227714 183172 227720 183184
rect 211396 183144 227720 183172
rect 211396 183132 211402 183144
rect 227714 183132 227720 183144
rect 227772 183132 227778 183184
rect 159910 183064 159916 183116
rect 159968 183104 159974 183116
rect 176562 183104 176568 183116
rect 159968 183076 176568 183104
rect 159968 183064 159974 183076
rect 176562 183064 176568 183076
rect 176620 183104 176626 183116
rect 247034 183104 247040 183116
rect 176620 183076 247040 183104
rect 176620 183064 176626 183076
rect 247034 183064 247040 183076
rect 247092 183064 247098 183116
rect 160370 182996 160376 183048
rect 160428 183036 160434 183048
rect 176378 183036 176384 183048
rect 160428 183008 176384 183036
rect 160428 182996 160434 183008
rect 176378 182996 176384 183008
rect 176436 183036 176442 183048
rect 349154 183036 349160 183048
rect 176436 183008 349160 183036
rect 176436 182996 176442 183008
rect 349154 182996 349160 183008
rect 349212 182996 349218 183048
rect 154942 182928 154948 182980
rect 155000 182968 155006 182980
rect 221090 182968 221096 182980
rect 155000 182940 221096 182968
rect 155000 182928 155006 182940
rect 221090 182928 221096 182940
rect 221148 182968 221154 182980
rect 552750 182968 552756 182980
rect 221148 182940 552756 182968
rect 221148 182928 221154 182940
rect 552750 182928 552756 182940
rect 552808 182928 552814 182980
rect 96522 182860 96528 182912
rect 96580 182900 96586 182912
rect 120534 182900 120540 182912
rect 96580 182872 120540 182900
rect 96580 182860 96586 182872
rect 120534 182860 120540 182872
rect 120592 182900 120598 182912
rect 140958 182900 140964 182912
rect 120592 182872 140964 182900
rect 120592 182860 120598 182872
rect 140958 182860 140964 182872
rect 141016 182860 141022 182912
rect 153470 182860 153476 182912
rect 153528 182900 153534 182912
rect 188614 182900 188620 182912
rect 153528 182872 188620 182900
rect 153528 182860 153534 182872
rect 188614 182860 188620 182872
rect 188672 182900 188678 182912
rect 569402 182900 569408 182912
rect 188672 182872 569408 182900
rect 188672 182860 188678 182872
rect 569402 182860 569408 182872
rect 569460 182860 569466 182912
rect 108298 182792 108304 182844
rect 108356 182832 108362 182844
rect 139670 182832 139676 182844
rect 108356 182804 139676 182832
rect 108356 182792 108362 182804
rect 139670 182792 139676 182804
rect 139728 182792 139734 182844
rect 158162 182792 158168 182844
rect 158220 182832 158226 182844
rect 177758 182832 177764 182844
rect 158220 182804 177764 182832
rect 158220 182792 158226 182804
rect 177758 182792 177764 182804
rect 177816 182832 177822 182844
rect 575198 182832 575204 182844
rect 177816 182804 575204 182832
rect 177816 182792 177822 182804
rect 575198 182792 575204 182804
rect 575256 182792 575262 182844
rect 102870 182180 102876 182232
rect 102928 182220 102934 182232
rect 105814 182220 105820 182232
rect 102928 182192 105820 182220
rect 102928 182180 102934 182192
rect 105814 182180 105820 182192
rect 105872 182180 105878 182232
rect 123110 182112 123116 182164
rect 123168 182152 123174 182164
rect 123570 182152 123576 182164
rect 123168 182124 123576 182152
rect 123168 182112 123174 182124
rect 123570 182112 123576 182124
rect 123628 182112 123634 182164
rect 125502 182112 125508 182164
rect 125560 182152 125566 182164
rect 125778 182152 125784 182164
rect 125560 182124 125784 182152
rect 125560 182112 125566 182124
rect 125778 182112 125784 182124
rect 125836 182112 125842 182164
rect 147858 182112 147864 182164
rect 147916 182152 147922 182164
rect 148410 182152 148416 182164
rect 147916 182124 148416 182152
rect 147916 182112 147922 182124
rect 148410 182112 148416 182124
rect 148468 182112 148474 182164
rect 149330 182112 149336 182164
rect 149388 182152 149394 182164
rect 149790 182152 149796 182164
rect 149388 182124 149796 182152
rect 149388 182112 149394 182124
rect 149790 182112 149796 182124
rect 149848 182112 149854 182164
rect 149882 182112 149888 182164
rect 149940 182152 149946 182164
rect 572346 182152 572352 182164
rect 149940 182124 572352 182152
rect 149940 182112 149946 182124
rect 572346 182112 572352 182124
rect 572404 182112 572410 182164
rect 141878 182084 141884 182096
rect 122806 182056 141884 182084
rect 108390 181976 108396 182028
rect 108448 182016 108454 182028
rect 122806 182016 122834 182056
rect 141878 182044 141884 182056
rect 141936 182044 141942 182096
rect 149808 182084 149836 182112
rect 561214 182084 561220 182096
rect 149808 182056 561220 182084
rect 561214 182044 561220 182056
rect 561272 182044 561278 182096
rect 139578 182016 139584 182028
rect 108448 181988 122834 182016
rect 136008 181988 139584 182016
rect 108448 181976 108454 181988
rect 107286 181908 107292 181960
rect 107344 181948 107350 181960
rect 136008 181948 136036 181988
rect 139578 181976 139584 181988
rect 139636 181976 139642 182028
rect 148410 181976 148416 182028
rect 148468 182016 148474 182028
rect 277394 182016 277400 182028
rect 148468 181988 277400 182016
rect 148468 181976 148474 181988
rect 277394 181976 277400 181988
rect 277452 181976 277458 182028
rect 107344 181920 136036 181948
rect 107344 181908 107350 181920
rect 137554 181908 137560 181960
rect 137612 181948 137618 181960
rect 140222 181948 140228 181960
rect 137612 181920 140228 181948
rect 137612 181908 137618 181920
rect 140222 181908 140228 181920
rect 140280 181948 140286 181960
rect 253934 181948 253940 181960
rect 140280 181920 253940 181948
rect 140280 181908 140286 181920
rect 253934 181908 253940 181920
rect 253992 181908 253998 181960
rect 104250 181840 104256 181892
rect 104308 181880 104314 181892
rect 137002 181880 137008 181892
rect 104308 181852 137008 181880
rect 104308 181840 104314 181852
rect 137002 181840 137008 181852
rect 137060 181840 137066 181892
rect 153286 181840 153292 181892
rect 153344 181880 153350 181892
rect 210602 181880 210608 181892
rect 153344 181852 210608 181880
rect 153344 181840 153350 181852
rect 210602 181840 210608 181852
rect 210660 181880 210666 181892
rect 217410 181880 217416 181892
rect 210660 181852 217416 181880
rect 210660 181840 210666 181852
rect 217410 181840 217416 181852
rect 217468 181840 217474 181892
rect 113818 181772 113824 181824
rect 113876 181812 113882 181824
rect 146662 181812 146668 181824
rect 113876 181784 146668 181812
rect 113876 181772 113882 181784
rect 146662 181772 146668 181784
rect 146720 181812 146726 181824
rect 149882 181812 149888 181824
rect 146720 181784 149888 181812
rect 146720 181772 146726 181784
rect 149882 181772 149888 181784
rect 149940 181772 149946 181824
rect 154758 181772 154764 181824
rect 154816 181812 154822 181824
rect 189442 181812 189448 181824
rect 154816 181784 189448 181812
rect 154816 181772 154822 181784
rect 189442 181772 189448 181784
rect 189500 181772 189506 181824
rect 119614 181704 119620 181756
rect 119672 181744 119678 181756
rect 152642 181744 152648 181756
rect 119672 181716 152648 181744
rect 119672 181704 119678 181716
rect 152642 181704 152648 181716
rect 152700 181704 152706 181756
rect 175458 181704 175464 181756
rect 175516 181744 175522 181756
rect 210326 181744 210332 181756
rect 175516 181716 210332 181744
rect 175516 181704 175522 181716
rect 210326 181704 210332 181716
rect 210384 181704 210390 181756
rect 103422 181636 103428 181688
rect 103480 181676 103486 181688
rect 137738 181676 137744 181688
rect 103480 181648 137744 181676
rect 103480 181636 103486 181648
rect 137738 181636 137744 181648
rect 137796 181636 137802 181688
rect 160278 181636 160284 181688
rect 160336 181676 160342 181688
rect 195146 181676 195152 181688
rect 160336 181648 195152 181676
rect 160336 181636 160342 181648
rect 195146 181636 195152 181648
rect 195204 181636 195210 181688
rect 105630 181568 105636 181620
rect 105688 181608 105694 181620
rect 138934 181608 138940 181620
rect 105688 181580 138940 181608
rect 105688 181568 105694 181580
rect 138934 181568 138940 181580
rect 138992 181568 138998 181620
rect 150618 181568 150624 181620
rect 150676 181608 150682 181620
rect 220814 181608 220820 181620
rect 150676 181580 220820 181608
rect 150676 181568 150682 181580
rect 220814 181568 220820 181580
rect 220872 181568 220878 181620
rect 99098 181500 99104 181552
rect 99156 181540 99162 181552
rect 132770 181540 132776 181552
rect 99156 181512 132776 181540
rect 99156 181500 99162 181512
rect 132770 181500 132776 181512
rect 132828 181500 132834 181552
rect 152366 181500 152372 181552
rect 152424 181540 152430 181552
rect 219986 181540 219992 181552
rect 152424 181512 219992 181540
rect 152424 181500 152430 181512
rect 219986 181500 219992 181512
rect 220044 181540 220050 181552
rect 299474 181540 299480 181552
rect 220044 181512 299480 181540
rect 220044 181500 220050 181512
rect 299474 181500 299480 181512
rect 299532 181500 299538 181552
rect 125778 181432 125784 181484
rect 125836 181472 125842 181484
rect 292574 181472 292580 181484
rect 125836 181444 292580 181472
rect 125836 181432 125842 181444
rect 292574 181432 292580 181444
rect 292632 181432 292638 181484
rect 176746 181364 176752 181416
rect 176804 181404 176810 181416
rect 211890 181404 211896 181416
rect 176804 181376 211896 181404
rect 176804 181364 176810 181376
rect 211890 181364 211896 181376
rect 211948 181364 211954 181416
rect 166258 181296 166264 181348
rect 166316 181336 166322 181348
rect 189258 181336 189264 181348
rect 166316 181308 189264 181336
rect 166316 181296 166322 181308
rect 189258 181296 189264 181308
rect 189316 181296 189322 181348
rect 102778 180956 102784 181008
rect 102836 180996 102842 181008
rect 123110 180996 123116 181008
rect 102836 180968 123116 180996
rect 102836 180956 102842 180968
rect 123110 180956 123116 180968
rect 123168 180956 123174 181008
rect 103146 180888 103152 180940
rect 103204 180928 103210 180940
rect 126882 180928 126888 180940
rect 103204 180900 126888 180928
rect 103204 180888 103210 180900
rect 126882 180888 126888 180900
rect 126940 180888 126946 180940
rect 101766 180820 101772 180872
rect 101824 180860 101830 180872
rect 129642 180860 129648 180872
rect 101824 180832 129648 180860
rect 101824 180820 101830 180832
rect 129642 180820 129648 180832
rect 129700 180820 129706 180872
rect 195146 180820 195152 180872
rect 195204 180860 195210 180872
rect 580166 180860 580172 180872
rect 195204 180832 580172 180860
rect 195204 180820 195210 180832
rect 580166 180820 580172 180832
rect 580224 180820 580230 180872
rect 3234 180752 3240 180804
rect 3292 180792 3298 180804
rect 112254 180792 112260 180804
rect 3292 180764 112260 180792
rect 3292 180752 3298 180764
rect 112254 180752 112260 180764
rect 112312 180752 112318 180804
rect 129182 180752 129188 180804
rect 129240 180792 129246 180804
rect 555418 180792 555424 180804
rect 129240 180764 555424 180792
rect 129240 180752 129246 180764
rect 555418 180752 555424 180764
rect 555476 180752 555482 180804
rect 126882 180684 126888 180736
rect 126940 180724 126946 180736
rect 136542 180724 136548 180736
rect 126940 180696 136548 180724
rect 126940 180684 126946 180696
rect 136542 180684 136548 180696
rect 136600 180724 136606 180736
rect 558454 180724 558460 180736
rect 136600 180696 558460 180724
rect 136600 180684 136606 180696
rect 558454 180684 558460 180696
rect 558512 180684 558518 180736
rect 127986 180616 127992 180668
rect 128044 180656 128050 180668
rect 541618 180656 541624 180668
rect 128044 180628 541624 180656
rect 128044 180616 128050 180628
rect 541618 180616 541624 180628
rect 541676 180616 541682 180668
rect 129642 180548 129648 180600
rect 129700 180588 129706 180600
rect 140038 180588 140044 180600
rect 129700 180560 140044 180588
rect 129700 180548 129706 180560
rect 140038 180548 140044 180560
rect 140096 180588 140102 180600
rect 552842 180588 552848 180600
rect 140096 180560 552848 180588
rect 140096 180548 140102 180560
rect 552842 180548 552848 180560
rect 552900 180548 552906 180600
rect 128170 180480 128176 180532
rect 128228 180520 128234 180532
rect 498194 180520 498200 180532
rect 128228 180492 498200 180520
rect 128228 180480 128234 180492
rect 498194 180480 498200 180492
rect 498252 180480 498258 180532
rect 128722 180412 128728 180464
rect 128780 180452 128786 180464
rect 138750 180452 138756 180464
rect 128780 180424 138756 180452
rect 128780 180412 128786 180424
rect 138750 180412 138756 180424
rect 138808 180452 138814 180464
rect 405734 180452 405740 180464
rect 138808 180424 405740 180452
rect 138808 180412 138814 180424
rect 405734 180412 405740 180424
rect 405792 180412 405798 180464
rect 123110 180344 123116 180396
rect 123168 180384 123174 180396
rect 322934 180384 322940 180396
rect 123168 180356 322940 180384
rect 123168 180344 123174 180356
rect 322934 180344 322940 180356
rect 322992 180344 322998 180396
rect 80698 180276 80704 180328
rect 80756 180316 80762 180328
rect 186314 180316 186320 180328
rect 80756 180288 186320 180316
rect 80756 180276 80762 180288
rect 186314 180276 186320 180288
rect 186372 180276 186378 180328
rect 86218 180208 86224 180260
rect 86276 180248 86282 180260
rect 186406 180248 186412 180260
rect 86276 180220 186412 180248
rect 86276 180208 86282 180220
rect 186406 180208 186412 180220
rect 186464 180248 186470 180260
rect 186464 180220 190454 180248
rect 186464 180208 186470 180220
rect 190426 180180 190454 180220
rect 212994 180180 213000 180192
rect 190426 180152 213000 180180
rect 212994 180140 213000 180152
rect 213052 180140 213058 180192
rect 186314 180072 186320 180124
rect 186372 180112 186378 180124
rect 219894 180112 219900 180124
rect 186372 180084 219900 180112
rect 186372 180072 186378 180084
rect 219894 180072 219900 180084
rect 219952 180072 219958 180124
rect 105722 179392 105728 179444
rect 105780 179432 105786 179444
rect 105780 179404 126744 179432
rect 105780 179392 105786 179404
rect 126716 179376 126744 179404
rect 126698 179324 126704 179376
rect 126756 179364 126762 179376
rect 582650 179364 582656 179376
rect 126756 179336 582656 179364
rect 126756 179324 126762 179336
rect 582650 179324 582656 179336
rect 582708 179324 582714 179376
rect 164418 179120 164424 179172
rect 164476 179160 164482 179172
rect 186498 179160 186504 179172
rect 164476 179132 186504 179160
rect 164476 179120 164482 179132
rect 186498 179120 186504 179132
rect 186556 179120 186562 179172
rect 163774 179052 163780 179104
rect 163832 179092 163838 179104
rect 190454 179092 190460 179104
rect 163832 179064 190460 179092
rect 163832 179052 163838 179064
rect 190454 179052 190460 179064
rect 190512 179052 190518 179104
rect 156138 178984 156144 179036
rect 156196 179024 156202 179036
rect 186590 179024 186596 179036
rect 156196 178996 186596 179024
rect 156196 178984 156202 178996
rect 186590 178984 186596 178996
rect 186648 178984 186654 179036
rect 101858 178916 101864 178968
rect 101916 178956 101922 178968
rect 134150 178956 134156 178968
rect 101916 178928 134156 178956
rect 101916 178916 101922 178928
rect 134150 178916 134156 178928
rect 134208 178916 134214 178968
rect 177298 178916 177304 178968
rect 177356 178956 177362 178968
rect 211522 178956 211528 178968
rect 177356 178928 211528 178956
rect 177356 178916 177362 178928
rect 211522 178916 211528 178928
rect 211580 178916 211586 178968
rect 87690 178848 87696 178900
rect 87748 178888 87754 178900
rect 104158 178888 104164 178900
rect 87748 178860 104164 178888
rect 87748 178848 87754 178860
rect 104158 178848 104164 178860
rect 104216 178888 104222 178900
rect 136910 178888 136916 178900
rect 104216 178860 136916 178888
rect 104216 178848 104222 178860
rect 136910 178848 136916 178860
rect 136968 178848 136974 178900
rect 171226 178848 171232 178900
rect 171284 178888 171290 178900
rect 215846 178888 215852 178900
rect 171284 178860 215852 178888
rect 171284 178848 171290 178860
rect 215846 178848 215852 178860
rect 215904 178848 215910 178900
rect 100386 178780 100392 178832
rect 100444 178820 100450 178832
rect 134058 178820 134064 178832
rect 100444 178792 134064 178820
rect 100444 178780 100450 178792
rect 134058 178780 134064 178792
rect 134116 178780 134122 178832
rect 154666 178780 154672 178832
rect 154724 178820 154730 178832
rect 217318 178820 217324 178832
rect 154724 178792 217324 178820
rect 154724 178780 154730 178792
rect 217318 178780 217324 178792
rect 217376 178780 217382 178832
rect 101674 178712 101680 178764
rect 101732 178752 101738 178764
rect 135990 178752 135996 178764
rect 101732 178724 135996 178752
rect 101732 178712 101738 178724
rect 135990 178712 135996 178724
rect 136048 178712 136054 178764
rect 160186 178712 160192 178764
rect 160244 178752 160250 178764
rect 184842 178752 184848 178764
rect 160244 178724 184848 178752
rect 160244 178712 160250 178724
rect 184842 178712 184848 178724
rect 184900 178752 184906 178764
rect 309778 178752 309784 178764
rect 184900 178724 309784 178752
rect 184900 178712 184906 178724
rect 309778 178712 309784 178724
rect 309836 178712 309842 178764
rect 109586 178644 109592 178696
rect 109644 178684 109650 178696
rect 150894 178684 150900 178696
rect 109644 178656 150900 178684
rect 109644 178644 109650 178656
rect 150894 178644 150900 178656
rect 150952 178644 150958 178696
rect 161290 178644 161296 178696
rect 161348 178684 161354 178696
rect 214742 178684 214748 178696
rect 161348 178656 214748 178684
rect 161348 178644 161354 178656
rect 214742 178644 214748 178656
rect 214800 178684 214806 178696
rect 425054 178684 425060 178696
rect 214800 178656 425060 178684
rect 214800 178644 214806 178656
rect 425054 178644 425060 178656
rect 425112 178644 425118 178696
rect 95142 178032 95148 178084
rect 95200 178072 95206 178084
rect 134518 178072 134524 178084
rect 95200 178044 134524 178072
rect 95200 178032 95206 178044
rect 134518 178032 134524 178044
rect 134576 178072 134582 178084
rect 135162 178072 135168 178084
rect 134576 178044 135168 178072
rect 134576 178032 134582 178044
rect 135162 178032 135168 178044
rect 135220 178032 135226 178084
rect 126606 177964 126612 178016
rect 126664 178004 126670 178016
rect 582374 178004 582380 178016
rect 126664 177976 582380 178004
rect 126664 177964 126670 177976
rect 582374 177964 582380 177976
rect 582432 177964 582438 178016
rect 124122 177896 124128 177948
rect 124180 177936 124186 177948
rect 561306 177936 561312 177948
rect 124180 177908 561312 177936
rect 124180 177896 124186 177908
rect 561306 177896 561312 177908
rect 561364 177896 561370 177948
rect 135162 177828 135168 177880
rect 135220 177868 135226 177880
rect 556982 177868 556988 177880
rect 135220 177840 556988 177868
rect 135220 177828 135226 177840
rect 556982 177828 556988 177840
rect 557040 177828 557046 177880
rect 140774 177760 140780 177812
rect 140832 177800 140838 177812
rect 141142 177800 141148 177812
rect 140832 177772 141148 177800
rect 140832 177760 140838 177772
rect 141142 177760 141148 177772
rect 141200 177800 141206 177812
rect 555510 177800 555516 177812
rect 141200 177772 555516 177800
rect 141200 177760 141206 177772
rect 555510 177760 555516 177772
rect 555568 177760 555574 177812
rect 140130 177732 140136 177744
rect 122806 177704 140136 177732
rect 105814 177352 105820 177404
rect 105872 177392 105878 177404
rect 122806 177392 122834 177704
rect 140130 177692 140136 177704
rect 140188 177732 140194 177744
rect 409874 177732 409880 177744
rect 140188 177704 409880 177732
rect 140188 177692 140194 177704
rect 409874 177692 409880 177704
rect 409932 177692 409938 177744
rect 137462 177624 137468 177676
rect 137520 177664 137526 177676
rect 364334 177664 364340 177676
rect 137520 177636 364340 177664
rect 137520 177624 137526 177636
rect 364334 177624 364340 177636
rect 364392 177624 364398 177676
rect 136818 177420 136824 177472
rect 136876 177460 136882 177472
rect 137462 177460 137468 177472
rect 136876 177432 137468 177460
rect 136876 177420 136882 177432
rect 137462 177420 137468 177432
rect 137520 177420 137526 177472
rect 105872 177364 122834 177392
rect 105872 177352 105878 177364
rect 192754 177352 192760 177404
rect 192812 177392 192818 177404
rect 221734 177392 221740 177404
rect 192812 177364 221740 177392
rect 192812 177352 192818 177364
rect 221734 177352 221740 177364
rect 221792 177352 221798 177404
rect 105538 177284 105544 177336
rect 105596 177324 105602 177336
rect 140774 177324 140780 177336
rect 105596 177296 140780 177324
rect 105596 177284 105602 177296
rect 140774 177284 140780 177296
rect 140832 177284 140838 177336
rect 141326 177284 141332 177336
rect 141384 177324 141390 177336
rect 142154 177324 142160 177336
rect 141384 177296 142160 177324
rect 141384 177284 141390 177296
rect 142154 177284 142160 177296
rect 142212 177324 142218 177336
rect 558546 177324 558552 177336
rect 142212 177296 558552 177324
rect 142212 177284 142218 177296
rect 558546 177284 558552 177296
rect 558604 177284 558610 177336
rect 221274 176672 221280 176724
rect 221332 176712 221338 176724
rect 221734 176712 221740 176724
rect 221332 176684 221740 176712
rect 221332 176672 221338 176684
rect 221734 176672 221740 176684
rect 221792 176712 221798 176724
rect 579798 176712 579804 176724
rect 221792 176684 579804 176712
rect 221792 176672 221798 176684
rect 579798 176672 579804 176684
rect 579856 176672 579862 176724
rect 133782 176604 133788 176656
rect 133840 176644 133846 176656
rect 559650 176644 559656 176656
rect 133840 176616 559656 176644
rect 133840 176604 133846 176616
rect 559650 176604 559656 176616
rect 559708 176604 559714 176656
rect 156598 176060 156604 176112
rect 156656 176100 156662 176112
rect 190914 176100 190920 176112
rect 156656 176072 190920 176100
rect 156656 176060 156662 176072
rect 190914 176060 190920 176072
rect 190972 176060 190978 176112
rect 169110 175992 169116 176044
rect 169168 176032 169174 176044
rect 208946 176032 208952 176044
rect 169168 176004 208952 176032
rect 169168 175992 169174 176004
rect 208946 175992 208952 176004
rect 209004 175992 209010 176044
rect 99006 175924 99012 175976
rect 99064 175964 99070 175976
rect 132678 175964 132684 175976
rect 99064 175936 132684 175964
rect 99064 175924 99070 175936
rect 132678 175924 132684 175936
rect 132736 175964 132742 175976
rect 133782 175964 133788 175976
rect 132736 175936 133788 175964
rect 132736 175924 132742 175936
rect 133782 175924 133788 175936
rect 133840 175924 133846 175976
rect 167638 175924 167644 175976
rect 167696 175964 167702 175976
rect 207658 175964 207664 175976
rect 167696 175936 207664 175964
rect 167696 175924 167702 175936
rect 207658 175924 207664 175936
rect 207716 175924 207722 175976
rect 135162 175176 135168 175228
rect 135220 175216 135226 175228
rect 565078 175216 565084 175228
rect 135220 175188 565084 175216
rect 135220 175176 135226 175188
rect 565078 175176 565084 175188
rect 565136 175176 565142 175228
rect 140866 175108 140872 175160
rect 140924 175148 140930 175160
rect 562318 175148 562324 175160
rect 140924 175120 562324 175148
rect 140924 175108 140930 175120
rect 562318 175108 562324 175120
rect 562376 175108 562382 175160
rect 140774 175040 140780 175092
rect 140832 175080 140838 175092
rect 368474 175080 368480 175092
rect 140832 175052 368480 175080
rect 140832 175040 140838 175052
rect 368474 175040 368480 175052
rect 368532 175040 368538 175092
rect 136542 174972 136548 175024
rect 136600 175012 136606 175024
rect 357434 175012 357440 175024
rect 136600 174984 357440 175012
rect 136600 174972 136606 174984
rect 357434 174972 357440 174984
rect 357492 174972 357498 175024
rect 353294 174944 353300 174956
rect 142126 174916 353300 174944
rect 101490 174700 101496 174752
rect 101548 174740 101554 174752
rect 134610 174740 134616 174752
rect 101548 174712 134616 174740
rect 101548 174700 101554 174712
rect 134610 174700 134616 174712
rect 134668 174740 134674 174752
rect 135162 174740 135168 174752
rect 134668 174712 135168 174740
rect 134668 174700 134674 174712
rect 135162 174700 135168 174712
rect 135220 174700 135226 174752
rect 102686 174632 102692 174684
rect 102744 174672 102750 174684
rect 135898 174672 135904 174684
rect 102744 174644 135904 174672
rect 102744 174632 102750 174644
rect 135898 174632 135904 174644
rect 135956 174672 135962 174684
rect 142126 174672 142154 174916
rect 353294 174904 353300 174916
rect 353352 174904 353358 174956
rect 135956 174644 142154 174672
rect 135956 174632 135962 174644
rect 101582 174564 101588 174616
rect 101640 174604 101646 174616
rect 136542 174604 136548 174616
rect 101640 174576 136548 174604
rect 101640 174564 101646 174576
rect 136542 174564 136548 174576
rect 136600 174564 136606 174616
rect 106918 174496 106924 174548
rect 106976 174536 106982 174548
rect 140774 174536 140780 174548
rect 106976 174508 140780 174536
rect 106976 174496 106982 174508
rect 140774 174496 140780 174508
rect 140832 174496 140838 174548
rect 124030 173884 124036 173936
rect 124088 173924 124094 173936
rect 140866 173924 140872 173936
rect 124088 173896 140872 173924
rect 124088 173884 124094 173896
rect 140866 173884 140872 173896
rect 140924 173884 140930 173936
rect 3234 172456 3240 172508
rect 3292 172496 3298 172508
rect 116578 172496 116584 172508
rect 3292 172468 116584 172496
rect 3292 172456 3298 172468
rect 116578 172456 116584 172468
rect 116636 172456 116642 172508
rect 3326 168308 3332 168360
rect 3384 168348 3390 168360
rect 25498 168348 25504 168360
rect 3384 168320 25504 168348
rect 3384 168308 3390 168320
rect 25498 168308 25504 168320
rect 25556 168308 25562 168360
rect 172238 164840 172244 164892
rect 172296 164880 172302 164892
rect 204990 164880 204996 164892
rect 172296 164852 204996 164880
rect 172296 164840 172302 164852
rect 204990 164840 204996 164852
rect 205048 164840 205054 164892
rect 204990 164228 204996 164280
rect 205048 164268 205054 164280
rect 580166 164268 580172 164280
rect 205048 164240 580172 164268
rect 205048 164228 205054 164240
rect 580166 164228 580172 164240
rect 580224 164228 580230 164280
rect 97442 163480 97448 163532
rect 97500 163520 97506 163532
rect 146570 163520 146576 163532
rect 97500 163492 146576 163520
rect 97500 163480 97506 163492
rect 146570 163480 146576 163492
rect 146628 163480 146634 163532
rect 3050 162868 3056 162920
rect 3108 162908 3114 162920
rect 97442 162908 97448 162920
rect 3108 162880 97448 162908
rect 3108 162868 3114 162880
rect 97442 162868 97448 162880
rect 97500 162868 97506 162920
rect 198090 157292 198096 157344
rect 198148 157332 198154 157344
rect 580166 157332 580172 157344
rect 198148 157304 580172 157332
rect 198148 157292 198154 157304
rect 580166 157292 580172 157304
rect 580224 157292 580230 157344
rect 3510 155864 3516 155916
rect 3568 155904 3574 155916
rect 117774 155904 117780 155916
rect 3568 155876 117780 155904
rect 3568 155864 3574 155876
rect 117774 155864 117780 155876
rect 117832 155864 117838 155916
rect 180242 155184 180248 155236
rect 180300 155224 180306 155236
rect 197354 155224 197360 155236
rect 180300 155196 197360 155224
rect 180300 155184 180306 155196
rect 197354 155184 197360 155196
rect 197412 155184 197418 155236
rect 192478 153144 192484 153196
rect 192536 153184 192542 153196
rect 199470 153184 199476 153196
rect 192536 153156 199476 153184
rect 192536 153144 192542 153156
rect 199470 153144 199476 153156
rect 199528 153144 199534 153196
rect 199470 151784 199476 151836
rect 199528 151824 199534 151836
rect 579798 151824 579804 151836
rect 199528 151796 579804 151824
rect 199528 151784 199534 151796
rect 579798 151784 579804 151796
rect 579856 151784 579862 151836
rect 100018 151240 100024 151292
rect 100076 151280 100082 151292
rect 132034 151280 132040 151292
rect 100076 151252 132040 151280
rect 100076 151240 100082 151252
rect 132034 151240 132040 151252
rect 132092 151240 132098 151292
rect 173342 151240 173348 151292
rect 173400 151280 173406 151292
rect 205082 151280 205088 151292
rect 173400 151252 205088 151280
rect 173400 151240 173406 151252
rect 205082 151240 205088 151252
rect 205140 151240 205146 151292
rect 94958 151172 94964 151224
rect 95016 151212 95022 151224
rect 138198 151212 138204 151224
rect 95016 151184 138204 151212
rect 95016 151172 95022 151184
rect 138198 151172 138204 151184
rect 138256 151172 138262 151224
rect 176010 151172 176016 151224
rect 176068 151212 176074 151224
rect 209130 151212 209136 151224
rect 176068 151184 209136 151212
rect 176068 151172 176074 151184
rect 209130 151172 209136 151184
rect 209188 151172 209194 151224
rect 95878 151104 95884 151156
rect 95936 151144 95942 151156
rect 140682 151144 140688 151156
rect 95936 151116 140688 151144
rect 95936 151104 95942 151116
rect 140682 151104 140688 151116
rect 140740 151104 140746 151156
rect 171870 151104 171876 151156
rect 171928 151144 171934 151156
rect 209038 151144 209044 151156
rect 171928 151116 209044 151144
rect 171928 151104 171934 151116
rect 209038 151104 209044 151116
rect 209096 151104 209102 151156
rect 95050 151036 95056 151088
rect 95108 151076 95114 151088
rect 140406 151076 140412 151088
rect 95108 151048 140412 151076
rect 95108 151036 95114 151048
rect 140406 151036 140412 151048
rect 140464 151036 140470 151088
rect 154298 151036 154304 151088
rect 154356 151076 154362 151088
rect 218606 151076 218612 151088
rect 154356 151048 218612 151076
rect 154356 151036 154362 151048
rect 218606 151036 218612 151048
rect 218664 151036 218670 151088
rect 106826 148996 106832 149048
rect 106884 149036 106890 149048
rect 131298 149036 131304 149048
rect 106884 149008 131304 149036
rect 106884 148996 106890 149008
rect 131298 148996 131304 149008
rect 131356 148996 131362 149048
rect 176286 148996 176292 149048
rect 176344 149036 176350 149048
rect 207750 149036 207756 149048
rect 176344 149008 207756 149036
rect 176344 148996 176350 149008
rect 207750 148996 207756 149008
rect 207808 148996 207814 149048
rect 101214 148928 101220 148980
rect 101272 148968 101278 148980
rect 126514 148968 126520 148980
rect 101272 148940 126520 148968
rect 101272 148928 101278 148940
rect 126514 148928 126520 148940
rect 126572 148928 126578 148980
rect 162762 148928 162768 148980
rect 162820 148968 162826 148980
rect 195422 148968 195428 148980
rect 162820 148940 195428 148968
rect 162820 148928 162826 148940
rect 195422 148928 195428 148940
rect 195480 148928 195486 148980
rect 102594 148860 102600 148912
rect 102652 148900 102658 148912
rect 135714 148900 135720 148912
rect 102652 148872 135720 148900
rect 102652 148860 102658 148872
rect 135714 148860 135720 148872
rect 135772 148860 135778 148912
rect 177482 148860 177488 148912
rect 177540 148900 177546 148912
rect 210602 148900 210608 148912
rect 177540 148872 210608 148900
rect 177540 148860 177546 148872
rect 210602 148860 210608 148872
rect 210660 148860 210666 148912
rect 103974 148792 103980 148844
rect 104032 148832 104038 148844
rect 137370 148832 137376 148844
rect 104032 148804 137376 148832
rect 104032 148792 104038 148804
rect 137370 148792 137376 148804
rect 137428 148792 137434 148844
rect 170674 148792 170680 148844
rect 170732 148832 170738 148844
rect 203242 148832 203248 148844
rect 170732 148804 203248 148832
rect 170732 148792 170738 148804
rect 203242 148792 203248 148804
rect 203300 148792 203306 148844
rect 114922 148724 114928 148776
rect 114980 148764 114986 148776
rect 150250 148764 150256 148776
rect 114980 148736 150256 148764
rect 114980 148724 114986 148736
rect 150250 148724 150256 148736
rect 150308 148724 150314 148776
rect 168650 148724 168656 148776
rect 168708 148764 168714 148776
rect 203426 148764 203432 148776
rect 168708 148736 203432 148764
rect 168708 148724 168714 148736
rect 203426 148724 203432 148736
rect 203484 148724 203490 148776
rect 98822 148656 98828 148708
rect 98880 148696 98886 148708
rect 133230 148696 133236 148708
rect 98880 148668 133236 148696
rect 98880 148656 98886 148668
rect 133230 148656 133236 148668
rect 133288 148656 133294 148708
rect 168558 148656 168564 148708
rect 168616 148696 168622 148708
rect 203334 148696 203340 148708
rect 168616 148668 203340 148696
rect 168616 148656 168622 148668
rect 203334 148656 203340 148668
rect 203392 148656 203398 148708
rect 98914 148588 98920 148640
rect 98972 148628 98978 148640
rect 133322 148628 133328 148640
rect 98972 148600 133328 148628
rect 98972 148588 98978 148600
rect 133322 148588 133328 148600
rect 133380 148588 133386 148640
rect 165890 148588 165896 148640
rect 165948 148628 165954 148640
rect 200666 148628 200672 148640
rect 165948 148600 200672 148628
rect 165948 148588 165954 148600
rect 200666 148588 200672 148600
rect 200724 148588 200730 148640
rect 99926 148520 99932 148572
rect 99984 148560 99990 148572
rect 134426 148560 134432 148572
rect 99984 148532 134432 148560
rect 99984 148520 99990 148532
rect 134426 148520 134432 148532
rect 134484 148520 134490 148572
rect 165798 148520 165804 148572
rect 165856 148560 165862 148572
rect 200574 148560 200580 148572
rect 165856 148532 200580 148560
rect 165856 148520 165862 148532
rect 200574 148520 200580 148532
rect 200632 148520 200638 148572
rect 98730 148452 98736 148504
rect 98788 148492 98794 148504
rect 133138 148492 133144 148504
rect 98788 148464 133144 148492
rect 98788 148452 98794 148464
rect 133138 148452 133144 148464
rect 133196 148452 133202 148504
rect 165430 148452 165436 148504
rect 165488 148492 165494 148504
rect 199654 148492 199660 148504
rect 165488 148464 199660 148492
rect 165488 148452 165494 148464
rect 199654 148452 199660 148464
rect 199712 148452 199718 148504
rect 101398 148384 101404 148436
rect 101456 148424 101462 148436
rect 137554 148424 137560 148436
rect 101456 148396 137560 148424
rect 101456 148384 101462 148396
rect 137554 148384 137560 148396
rect 137612 148384 137618 148436
rect 168282 148384 168288 148436
rect 168340 148424 168346 148436
rect 203610 148424 203616 148436
rect 168340 148396 203616 148424
rect 168340 148384 168346 148396
rect 203610 148384 203616 148396
rect 203668 148384 203674 148436
rect 96522 148316 96528 148368
rect 96580 148356 96586 148368
rect 130378 148356 130384 148368
rect 96580 148328 130384 148356
rect 96580 148316 96586 148328
rect 130378 148316 130384 148328
rect 130436 148316 130442 148368
rect 174538 148316 174544 148368
rect 174596 148356 174602 148368
rect 211982 148356 211988 148368
rect 174596 148328 211988 148356
rect 174596 148316 174602 148328
rect 211982 148316 211988 148328
rect 212040 148316 212046 148368
rect 106734 148248 106740 148300
rect 106792 148288 106798 148300
rect 127894 148288 127900 148300
rect 106792 148260 127900 148288
rect 106792 148248 106798 148260
rect 127894 148248 127900 148260
rect 127952 148248 127958 148300
rect 175274 148248 175280 148300
rect 175332 148288 175338 148300
rect 206462 148288 206468 148300
rect 175332 148260 206468 148288
rect 175332 148248 175338 148260
rect 206462 148248 206468 148260
rect 206520 148248 206526 148300
rect 121178 148180 121184 148232
rect 121236 148220 121242 148232
rect 127802 148220 127808 148232
rect 121236 148192 127808 148220
rect 121236 148180 121242 148192
rect 127802 148180 127808 148192
rect 127860 148180 127866 148232
rect 172146 148180 172152 148232
rect 172204 148220 172210 148232
rect 200758 148220 200764 148232
rect 172204 148192 200764 148220
rect 172204 148180 172210 148192
rect 200758 148180 200764 148192
rect 200816 148180 200822 148232
rect 120718 148112 120724 148164
rect 120776 148152 120782 148164
rect 125686 148152 125692 148164
rect 120776 148124 125692 148152
rect 120776 148112 120782 148124
rect 125686 148112 125692 148124
rect 125744 148112 125750 148164
rect 169386 148112 169392 148164
rect 169444 148152 169450 148164
rect 191374 148152 191380 148164
rect 169444 148124 191380 148152
rect 169444 148112 169450 148124
rect 191374 148112 191380 148124
rect 191432 148112 191438 148164
rect 3418 147568 3424 147620
rect 3476 147608 3482 147620
rect 114094 147608 114100 147620
rect 3476 147580 114100 147608
rect 3476 147568 3482 147580
rect 114094 147568 114100 147580
rect 114152 147608 114158 147620
rect 120902 147608 120908 147620
rect 114152 147580 120908 147608
rect 114152 147568 114158 147580
rect 120902 147568 120908 147580
rect 120960 147568 120966 147620
rect 580350 147608 580356 147620
rect 200086 147580 580356 147608
rect 185670 147228 185676 147280
rect 185728 147268 185734 147280
rect 196434 147268 196440 147280
rect 185728 147240 196440 147268
rect 185728 147228 185734 147240
rect 196434 147228 196440 147240
rect 196492 147268 196498 147280
rect 200086 147268 200114 147580
rect 580350 147568 580356 147580
rect 580408 147568 580414 147620
rect 196492 147240 200114 147268
rect 196492 147228 196498 147240
rect 165706 147160 165712 147212
rect 165764 147200 165770 147212
rect 192754 147200 192760 147212
rect 165764 147172 192760 147200
rect 165764 147160 165770 147172
rect 192754 147160 192760 147172
rect 192812 147160 192818 147212
rect 169018 147092 169024 147144
rect 169076 147132 169082 147144
rect 203518 147132 203524 147144
rect 169076 147104 203524 147132
rect 169076 147092 169082 147104
rect 203518 147092 203524 147104
rect 203576 147092 203582 147144
rect 117038 147024 117044 147076
rect 117096 147064 117102 147076
rect 117222 147064 117228 147076
rect 117096 147036 117228 147064
rect 117096 147024 117102 147036
rect 117222 147024 117228 147036
rect 117280 147024 117286 147076
rect 168098 147024 168104 147076
rect 168156 147064 168162 147076
rect 202138 147064 202144 147076
rect 168156 147036 202144 147064
rect 168156 147024 168162 147036
rect 202138 147024 202144 147036
rect 202196 147024 202202 147076
rect 111426 146956 111432 147008
rect 111484 146996 111490 147008
rect 138658 146996 138664 147008
rect 111484 146968 138664 146996
rect 111484 146956 111490 146968
rect 138658 146956 138664 146968
rect 138716 146956 138722 147008
rect 154114 146956 154120 147008
rect 154172 146996 154178 147008
rect 187694 146996 187700 147008
rect 154172 146968 187700 146996
rect 154172 146956 154178 146968
rect 187694 146956 187700 146968
rect 187752 146956 187758 147008
rect 188154 146956 188160 147008
rect 188212 146996 188218 147008
rect 188982 146996 188988 147008
rect 188212 146968 188988 146996
rect 188212 146956 188218 146968
rect 188982 146956 188988 146968
rect 189040 146956 189046 147008
rect 104066 146888 104072 146940
rect 104124 146928 104130 146940
rect 139026 146928 139032 146940
rect 104124 146900 139032 146928
rect 104124 146888 104130 146900
rect 139026 146888 139032 146900
rect 139084 146888 139090 146940
rect 156690 146888 156696 146940
rect 156748 146928 156754 146940
rect 216030 146928 216036 146940
rect 156748 146900 216036 146928
rect 156748 146888 156754 146900
rect 216030 146888 216036 146900
rect 216088 146888 216094 146940
rect 179690 146344 179696 146396
rect 179748 146384 179754 146396
rect 180150 146384 180156 146396
rect 179748 146356 180156 146384
rect 179748 146344 179754 146356
rect 180150 146344 180156 146356
rect 180208 146384 180214 146396
rect 215938 146384 215944 146396
rect 180208 146356 215944 146384
rect 180208 146344 180214 146356
rect 215938 146344 215944 146356
rect 215996 146344 216002 146396
rect 216030 146344 216036 146396
rect 216088 146384 216094 146396
rect 580810 146384 580816 146396
rect 216088 146356 580816 146384
rect 216088 146344 216094 146356
rect 580810 146344 580816 146356
rect 580868 146344 580874 146396
rect 187694 146276 187700 146328
rect 187752 146316 187758 146328
rect 188798 146316 188804 146328
rect 187752 146288 188804 146316
rect 187752 146276 187758 146288
rect 188798 146276 188804 146288
rect 188856 146316 188862 146328
rect 580902 146316 580908 146328
rect 188856 146288 580908 146316
rect 188856 146276 188862 146288
rect 580902 146276 580908 146288
rect 580960 146276 580966 146328
rect 117866 146208 117872 146260
rect 117924 146248 117930 146260
rect 130102 146248 130108 146260
rect 117924 146220 130108 146248
rect 117924 146208 117930 146220
rect 130102 146208 130108 146220
rect 130160 146208 130166 146260
rect 171502 146208 171508 146260
rect 171560 146248 171566 146260
rect 196250 146248 196256 146260
rect 171560 146220 196256 146248
rect 171560 146208 171566 146220
rect 196250 146208 196256 146220
rect 196308 146208 196314 146260
rect 490558 146208 490564 146260
rect 490616 146248 490622 146260
rect 580166 146248 580172 146260
rect 490616 146220 580172 146248
rect 490616 146208 490622 146220
rect 580166 146208 580172 146220
rect 580224 146208 580230 146260
rect 112346 146140 112352 146192
rect 112404 146180 112410 146192
rect 129366 146180 129372 146192
rect 112404 146152 129372 146180
rect 112404 146140 112410 146152
rect 129366 146140 129372 146152
rect 129424 146140 129430 146192
rect 172514 146140 172520 146192
rect 172572 146180 172578 146192
rect 199194 146180 199200 146192
rect 172572 146152 199200 146180
rect 172572 146140 172578 146152
rect 199194 146140 199200 146152
rect 199252 146140 199258 146192
rect 114278 146072 114284 146124
rect 114336 146112 114342 146124
rect 134794 146112 134800 146124
rect 114336 146084 134800 146112
rect 114336 146072 114342 146084
rect 134794 146072 134800 146084
rect 134852 146072 134858 146124
rect 164418 146072 164424 146124
rect 164476 146112 164482 146124
rect 193766 146112 193772 146124
rect 164476 146084 193772 146112
rect 164476 146072 164482 146084
rect 193766 146072 193772 146084
rect 193824 146072 193830 146124
rect 111150 146004 111156 146056
rect 111208 146044 111214 146056
rect 132586 146044 132592 146056
rect 111208 146016 132592 146044
rect 111208 146004 111214 146016
rect 132586 146004 132592 146016
rect 132644 146004 132650 146056
rect 166534 146004 166540 146056
rect 166592 146044 166598 146056
rect 196342 146044 196348 146056
rect 166592 146016 196348 146044
rect 166592 146004 166598 146016
rect 196342 146004 196348 146016
rect 196400 146004 196406 146056
rect 111242 145936 111248 145988
rect 111300 145976 111306 145988
rect 137186 145976 137192 145988
rect 111300 145948 137192 145976
rect 111300 145936 111306 145948
rect 137186 145936 137192 145948
rect 137244 145936 137250 145988
rect 167362 145936 167368 145988
rect 167420 145976 167426 145988
rect 199102 145976 199108 145988
rect 167420 145948 199108 145976
rect 167420 145936 167426 145948
rect 199102 145936 199108 145948
rect 199160 145936 199166 145988
rect 112714 145868 112720 145920
rect 112772 145908 112778 145920
rect 139394 145908 139400 145920
rect 112772 145880 139400 145908
rect 112772 145868 112778 145880
rect 139394 145868 139400 145880
rect 139452 145868 139458 145920
rect 162394 145868 162400 145920
rect 162452 145908 162458 145920
rect 194778 145908 194784 145920
rect 162452 145880 194784 145908
rect 162452 145868 162458 145880
rect 194778 145868 194784 145880
rect 194836 145868 194842 145920
rect 114002 145800 114008 145852
rect 114060 145840 114066 145852
rect 144914 145840 144920 145852
rect 114060 145812 144920 145840
rect 114060 145800 114066 145812
rect 144914 145800 144920 145812
rect 144972 145800 144978 145852
rect 164878 145800 164884 145852
rect 164936 145840 164942 145852
rect 197814 145840 197820 145852
rect 164936 145812 197820 145840
rect 164936 145800 164942 145812
rect 197814 145800 197820 145812
rect 197872 145800 197878 145852
rect 114186 145732 114192 145784
rect 114244 145772 114250 145784
rect 146478 145772 146484 145784
rect 114244 145744 146484 145772
rect 114244 145732 114250 145744
rect 146478 145732 146484 145744
rect 146536 145732 146542 145784
rect 156598 145732 156604 145784
rect 156656 145772 156662 145784
rect 190730 145772 190736 145784
rect 156656 145744 190736 145772
rect 156656 145732 156662 145744
rect 190730 145732 190736 145744
rect 190788 145732 190794 145784
rect 116762 145664 116768 145716
rect 116820 145704 116826 145716
rect 149974 145704 149980 145716
rect 116820 145676 149980 145704
rect 116820 145664 116826 145676
rect 149974 145664 149980 145676
rect 150032 145664 150038 145716
rect 160094 145664 160100 145716
rect 160152 145704 160158 145716
rect 194962 145704 194968 145716
rect 160152 145676 194968 145704
rect 160152 145664 160158 145676
rect 194962 145664 194968 145676
rect 195020 145664 195026 145716
rect 112714 145596 112720 145648
rect 112772 145636 112778 145648
rect 146570 145636 146576 145648
rect 112772 145608 146576 145636
rect 112772 145596 112778 145608
rect 146570 145596 146576 145608
rect 146628 145596 146634 145648
rect 157426 145596 157432 145648
rect 157484 145636 157490 145648
rect 192570 145636 192576 145648
rect 157484 145608 192576 145636
rect 157484 145596 157490 145608
rect 192570 145596 192576 145608
rect 192628 145596 192634 145648
rect 112254 145528 112260 145580
rect 112312 145568 112318 145580
rect 151170 145568 151176 145580
rect 112312 145540 151176 145568
rect 112312 145528 112318 145540
rect 151170 145528 151176 145540
rect 151228 145528 151234 145580
rect 154942 145528 154948 145580
rect 155000 145568 155006 145580
rect 189902 145568 189908 145580
rect 155000 145540 189908 145568
rect 155000 145528 155006 145540
rect 189902 145528 189908 145540
rect 189960 145528 189966 145580
rect 112162 145460 112168 145512
rect 112220 145500 112226 145512
rect 123386 145500 123392 145512
rect 112220 145472 123392 145500
rect 112220 145460 112226 145472
rect 123386 145460 123392 145472
rect 123444 145460 123450 145512
rect 176654 145460 176660 145512
rect 176712 145500 176718 145512
rect 196526 145500 196532 145512
rect 176712 145472 196532 145500
rect 176712 145460 176718 145472
rect 196526 145460 196532 145472
rect 196584 145460 196590 145512
rect 116670 145392 116676 145444
rect 116728 145432 116734 145444
rect 127710 145432 127716 145444
rect 116728 145404 127716 145432
rect 116728 145392 116734 145404
rect 127710 145392 127716 145404
rect 127768 145392 127774 145444
rect 179414 145392 179420 145444
rect 179472 145432 179478 145444
rect 197538 145432 197544 145444
rect 179472 145404 197544 145432
rect 179472 145392 179478 145404
rect 197538 145392 197544 145404
rect 197596 145392 197602 145444
rect 114094 145324 114100 145376
rect 114152 145364 114158 145376
rect 124214 145364 124220 145376
rect 114152 145336 124220 145364
rect 114152 145324 114158 145336
rect 124214 145324 124220 145336
rect 124272 145324 124278 145376
rect 180794 145324 180800 145376
rect 180852 145364 180858 145376
rect 197906 145364 197912 145376
rect 180852 145336 197912 145364
rect 180852 145324 180858 145336
rect 197906 145324 197912 145336
rect 197964 145324 197970 145376
rect 119338 144916 119344 144968
rect 119396 144956 119402 144968
rect 119706 144956 119712 144968
rect 119396 144928 119712 144956
rect 119396 144916 119402 144928
rect 119706 144916 119712 144928
rect 119764 144916 119770 144968
rect 3142 144848 3148 144900
rect 3200 144888 3206 144900
rect 179690 144888 179696 144900
rect 3200 144860 179696 144888
rect 3200 144848 3206 144860
rect 179690 144848 179696 144860
rect 179748 144848 179754 144900
rect 580258 144888 580264 144900
rect 200086 144860 580264 144888
rect 112898 144780 112904 144832
rect 112956 144820 112962 144832
rect 139762 144820 139768 144832
rect 112956 144792 139768 144820
rect 112956 144780 112962 144792
rect 139762 144780 139768 144792
rect 139820 144780 139826 144832
rect 175090 144780 175096 144832
rect 175148 144820 175154 144832
rect 193490 144820 193496 144832
rect 175148 144792 193496 144820
rect 175148 144780 175154 144792
rect 193490 144780 193496 144792
rect 193548 144780 193554 144832
rect 112806 144712 112812 144764
rect 112864 144752 112870 144764
rect 141786 144752 141792 144764
rect 112864 144724 141792 144752
rect 112864 144712 112870 144724
rect 141786 144712 141792 144724
rect 141844 144712 141850 144764
rect 173802 144712 173808 144764
rect 173860 144752 173866 144764
rect 193674 144752 193680 144764
rect 173860 144724 193680 144752
rect 173860 144712 173866 144724
rect 193674 144712 193680 144724
rect 193732 144752 193738 144764
rect 200086 144752 200114 144860
rect 580258 144848 580264 144860
rect 580316 144848 580322 144900
rect 193732 144724 200114 144752
rect 193732 144712 193738 144724
rect 116486 144644 116492 144696
rect 116544 144684 116550 144696
rect 148870 144684 148876 144696
rect 116544 144656 148876 144684
rect 116544 144644 116550 144656
rect 148870 144644 148876 144656
rect 148928 144644 148934 144696
rect 173986 144644 173992 144696
rect 174044 144684 174050 144696
rect 197630 144684 197636 144696
rect 174044 144656 197636 144684
rect 174044 144644 174050 144656
rect 197630 144644 197636 144656
rect 197688 144644 197694 144696
rect 110230 144576 110236 144628
rect 110288 144616 110294 144628
rect 142154 144616 142160 144628
rect 110288 144588 142160 144616
rect 110288 144576 110294 144588
rect 142154 144576 142160 144588
rect 142212 144576 142218 144628
rect 175182 144576 175188 144628
rect 175240 144616 175246 144628
rect 199010 144616 199016 144628
rect 175240 144588 199016 144616
rect 175240 144576 175246 144588
rect 199010 144576 199016 144588
rect 199068 144576 199074 144628
rect 115658 144508 115664 144560
rect 115716 144548 115722 144560
rect 148686 144548 148692 144560
rect 115716 144520 148692 144548
rect 115716 144508 115722 144520
rect 148686 144508 148692 144520
rect 148744 144508 148750 144560
rect 162946 144508 162952 144560
rect 163004 144548 163010 144560
rect 197538 144548 197544 144560
rect 163004 144520 197544 144548
rect 163004 144508 163010 144520
rect 197538 144508 197544 144520
rect 197596 144508 197602 144560
rect 114278 144440 114284 144492
rect 114336 144480 114342 144492
rect 146386 144480 146392 144492
rect 114336 144452 146392 144480
rect 114336 144440 114342 144452
rect 146386 144440 146392 144452
rect 146444 144440 146450 144492
rect 162302 144440 162308 144492
rect 162360 144480 162366 144492
rect 196526 144480 196532 144492
rect 162360 144452 196532 144480
rect 162360 144440 162366 144452
rect 196526 144440 196532 144452
rect 196584 144440 196590 144492
rect 118510 144372 118516 144424
rect 118568 144412 118574 144424
rect 151078 144412 151084 144424
rect 118568 144384 151084 144412
rect 118568 144372 118574 144384
rect 151078 144372 151084 144384
rect 151136 144372 151142 144424
rect 162486 144372 162492 144424
rect 162544 144412 162550 144424
rect 196434 144412 196440 144424
rect 162544 144384 196440 144412
rect 162544 144372 162550 144384
rect 196434 144372 196440 144384
rect 196492 144372 196498 144424
rect 119706 144304 119712 144356
rect 119764 144344 119770 144356
rect 152550 144344 152556 144356
rect 119764 144316 152556 144344
rect 119764 144304 119770 144316
rect 152550 144304 152556 144316
rect 152608 144304 152614 144356
rect 168006 144304 168012 144356
rect 168064 144344 168070 144356
rect 202046 144344 202052 144356
rect 168064 144316 202052 144344
rect 168064 144304 168070 144316
rect 202046 144304 202052 144316
rect 202104 144304 202110 144356
rect 105354 144236 105360 144288
rect 105412 144276 105418 144288
rect 166718 144276 166724 144288
rect 105412 144248 166724 144276
rect 105412 144236 105418 144248
rect 166718 144236 166724 144248
rect 166776 144276 166782 144288
rect 207842 144276 207848 144288
rect 166776 144248 207848 144276
rect 166776 144236 166782 144248
rect 207842 144236 207848 144248
rect 207900 144236 207906 144288
rect 117130 144168 117136 144220
rect 117188 144208 117194 144220
rect 178034 144208 178040 144220
rect 117188 144180 178040 144208
rect 117188 144168 117194 144180
rect 178034 144168 178040 144180
rect 178092 144168 178098 144220
rect 179046 144168 179052 144220
rect 179104 144208 179110 144220
rect 194778 144208 194784 144220
rect 179104 144180 194784 144208
rect 179104 144168 179110 144180
rect 194778 144168 194784 144180
rect 194836 144168 194842 144220
rect 116670 144100 116676 144152
rect 116728 144140 116734 144152
rect 131666 144140 131672 144152
rect 116728 144112 131672 144140
rect 116728 144100 116734 144112
rect 131666 144100 131672 144112
rect 131724 144100 131730 144152
rect 177758 144100 177764 144152
rect 177816 144140 177822 144152
rect 192846 144140 192852 144152
rect 177816 144112 192852 144140
rect 177816 144100 177822 144112
rect 192846 144100 192852 144112
rect 192904 144100 192910 144152
rect 116210 144032 116216 144084
rect 116268 144072 116274 144084
rect 128354 144072 128360 144084
rect 116268 144044 128360 144072
rect 116268 144032 116274 144044
rect 128354 144032 128360 144044
rect 128412 144032 128418 144084
rect 139762 143692 139768 143744
rect 139820 143732 139826 143744
rect 140406 143732 140412 143744
rect 139820 143704 140412 143732
rect 139820 143692 139826 143704
rect 140406 143692 140412 143704
rect 140464 143732 140470 143744
rect 191834 143732 191840 143744
rect 140464 143704 191840 143732
rect 140464 143692 140470 143704
rect 191834 143692 191840 143704
rect 191892 143692 191898 143744
rect 95786 143624 95792 143676
rect 95844 143664 95850 143676
rect 164418 143664 164424 143676
rect 95844 143636 164424 143664
rect 95844 143624 95850 143636
rect 164418 143624 164424 143636
rect 164476 143624 164482 143676
rect 196342 143624 196348 143676
rect 196400 143664 196406 143676
rect 196618 143664 196624 143676
rect 196400 143636 196624 143664
rect 196400 143624 196406 143636
rect 196618 143624 196624 143636
rect 196676 143664 196682 143676
rect 580534 143664 580540 143676
rect 196676 143636 580540 143664
rect 196676 143624 196682 143636
rect 580534 143624 580540 143636
rect 580592 143624 580598 143676
rect 134794 143556 134800 143608
rect 134852 143596 134858 143608
rect 580442 143596 580448 143608
rect 134852 143568 580448 143596
rect 134852 143556 134858 143568
rect 580442 143556 580448 143568
rect 580500 143556 580506 143608
rect 115290 143488 115296 143540
rect 115348 143528 115354 143540
rect 128538 143528 128544 143540
rect 115348 143500 128544 143528
rect 115348 143488 115354 143500
rect 128538 143488 128544 143500
rect 128596 143488 128602 143540
rect 188890 143488 188896 143540
rect 188948 143528 188954 143540
rect 196250 143528 196256 143540
rect 188948 143500 196256 143528
rect 188948 143488 188954 143500
rect 196250 143488 196256 143500
rect 196308 143488 196314 143540
rect 112622 143420 112628 143472
rect 112680 143460 112686 143472
rect 119890 143460 119896 143472
rect 112680 143432 119896 143460
rect 112680 143420 112686 143432
rect 119890 143420 119896 143432
rect 119948 143420 119954 143472
rect 120074 143420 120080 143472
rect 120132 143460 120138 143472
rect 121362 143460 121368 143472
rect 120132 143432 121368 143460
rect 120132 143420 120138 143432
rect 121362 143420 121368 143432
rect 121420 143420 121426 143472
rect 121454 143420 121460 143472
rect 121512 143460 121518 143472
rect 122190 143460 122196 143472
rect 121512 143432 122196 143460
rect 121512 143420 121518 143432
rect 122190 143420 122196 143432
rect 122248 143420 122254 143472
rect 181346 143420 181352 143472
rect 181404 143460 181410 143472
rect 190638 143460 190644 143472
rect 181404 143432 190644 143460
rect 181404 143420 181410 143432
rect 190638 143420 190644 143432
rect 190696 143420 190702 143472
rect 115382 143352 115388 143404
rect 115440 143392 115446 143404
rect 135990 143392 135996 143404
rect 115440 143364 135996 143392
rect 115440 143352 115446 143364
rect 135990 143352 135996 143364
rect 136048 143352 136054 143404
rect 185486 143352 185492 143404
rect 185544 143392 185550 143404
rect 196158 143392 196164 143404
rect 185544 143364 196164 143392
rect 185544 143352 185550 143364
rect 196158 143352 196164 143364
rect 196216 143352 196222 143404
rect 115566 143284 115572 143336
rect 115624 143324 115630 143336
rect 138474 143324 138480 143336
rect 115624 143296 138480 143324
rect 115624 143284 115630 143296
rect 138474 143284 138480 143296
rect 138532 143284 138538 143336
rect 183462 143284 183468 143336
rect 183520 143324 183526 143336
rect 195054 143324 195060 143336
rect 183520 143296 195060 143324
rect 183520 143284 183526 143296
rect 195054 143284 195060 143296
rect 195112 143284 195118 143336
rect 119890 143216 119896 143268
rect 119948 143256 119954 143268
rect 126974 143256 126980 143268
rect 119948 143228 126980 143256
rect 119948 143216 119954 143228
rect 126974 143216 126980 143228
rect 127032 143216 127038 143268
rect 127066 143216 127072 143268
rect 127124 143256 127130 143268
rect 143626 143256 143632 143268
rect 127124 143228 143632 143256
rect 127124 143216 127130 143228
rect 143626 143216 143632 143228
rect 143684 143216 143690 143268
rect 184658 143216 184664 143268
rect 184716 143256 184722 143268
rect 197814 143256 197820 143268
rect 184716 143228 197820 143256
rect 184716 143216 184722 143228
rect 197814 143216 197820 143228
rect 197872 143216 197878 143268
rect 116946 143148 116952 143200
rect 117004 143188 117010 143200
rect 141234 143188 141240 143200
rect 117004 143160 141240 143188
rect 117004 143148 117010 143160
rect 141234 143148 141240 143160
rect 141292 143148 141298 143200
rect 159818 143148 159824 143200
rect 159876 143188 159882 143200
rect 173802 143188 173808 143200
rect 159876 143160 173808 143188
rect 159876 143148 159882 143160
rect 173802 143148 173808 143160
rect 173860 143148 173866 143200
rect 178862 143148 178868 143200
rect 178920 143188 178926 143200
rect 192202 143188 192208 143200
rect 178920 143160 192208 143188
rect 178920 143148 178926 143160
rect 192202 143148 192208 143160
rect 192260 143188 192266 143200
rect 192260 143160 200114 143188
rect 192260 143148 192266 143160
rect 97994 143080 98000 143132
rect 98052 143120 98058 143132
rect 116854 143120 116860 143132
rect 98052 143092 116860 143120
rect 98052 143080 98058 143092
rect 116854 143080 116860 143092
rect 116912 143080 116918 143132
rect 117038 143080 117044 143132
rect 117096 143120 117102 143132
rect 146754 143120 146760 143132
rect 117096 143092 146760 143120
rect 117096 143080 117102 143092
rect 146754 143080 146760 143092
rect 146812 143080 146818 143132
rect 168926 143080 168932 143132
rect 168984 143120 168990 143132
rect 192662 143120 192668 143132
rect 168984 143092 192668 143120
rect 168984 143080 168990 143092
rect 192662 143080 192668 143092
rect 192720 143080 192726 143132
rect 110414 143012 110420 143064
rect 110472 143052 110478 143064
rect 111610 143052 111616 143064
rect 110472 143024 111616 143052
rect 110472 143012 110478 143024
rect 111610 143012 111616 143024
rect 111668 143052 111674 143064
rect 142614 143052 142620 143064
rect 111668 143024 142620 143052
rect 111668 143012 111674 143024
rect 142614 143012 142620 143024
rect 142672 143012 142678 143064
rect 162302 143012 162308 143064
rect 162360 143052 162366 143064
rect 185670 143052 185676 143064
rect 162360 143024 185676 143052
rect 162360 143012 162366 143024
rect 185670 143012 185676 143024
rect 185728 143012 185734 143064
rect 200086 143052 200114 143160
rect 211246 143052 211252 143064
rect 200086 143024 211252 143052
rect 211246 143012 211252 143024
rect 211304 143012 211310 143064
rect 82814 142944 82820 142996
rect 82872 142984 82878 142996
rect 115290 142984 115296 142996
rect 82872 142956 115296 142984
rect 82872 142944 82878 142956
rect 115290 142944 115296 142956
rect 115348 142944 115354 142996
rect 115750 142944 115756 142996
rect 115808 142984 115814 142996
rect 147674 142984 147680 142996
rect 115808 142956 147680 142984
rect 115808 142944 115814 142956
rect 147674 142944 147680 142956
rect 147732 142944 147738 142996
rect 166442 142944 166448 142996
rect 166500 142984 166506 142996
rect 192110 142984 192116 142996
rect 166500 142956 192116 142984
rect 166500 142944 166506 142956
rect 192110 142944 192116 142956
rect 192168 142984 192174 142996
rect 213086 142984 213092 142996
rect 192168 142956 213092 142984
rect 192168 142944 192174 142956
rect 213086 142944 213092 142956
rect 213144 142944 213150 142996
rect 97350 142876 97356 142928
rect 97408 142916 97414 142928
rect 137094 142916 137100 142928
rect 97408 142888 137100 142916
rect 97408 142876 97414 142888
rect 137094 142876 137100 142888
rect 137152 142876 137158 142928
rect 169662 142876 169668 142928
rect 169720 142916 169726 142928
rect 196342 142916 196348 142928
rect 169720 142888 196348 142916
rect 169720 142876 169726 142888
rect 196342 142876 196348 142888
rect 196400 142876 196406 142928
rect 44174 142808 44180 142860
rect 44232 142848 44238 142860
rect 110414 142848 110420 142860
rect 44232 142820 110420 142848
rect 44232 142808 44238 142820
rect 110414 142808 110420 142820
rect 110472 142808 110478 142860
rect 115106 142808 115112 142860
rect 115164 142848 115170 142860
rect 148318 142848 148324 142860
rect 115164 142820 148324 142848
rect 115164 142808 115170 142820
rect 148318 142808 148324 142820
rect 148376 142808 148382 142860
rect 158622 142808 158628 142860
rect 158680 142848 158686 142860
rect 191190 142848 191196 142860
rect 158680 142820 191196 142848
rect 158680 142808 158686 142820
rect 191190 142808 191196 142820
rect 191248 142808 191254 142860
rect 197814 142808 197820 142860
rect 197872 142848 197878 142860
rect 198366 142848 198372 142860
rect 197872 142820 198372 142848
rect 197872 142808 197878 142820
rect 198366 142808 198372 142820
rect 198424 142848 198430 142860
rect 329834 142848 329840 142860
rect 198424 142820 329840 142848
rect 198424 142808 198430 142820
rect 329834 142808 329840 142820
rect 329892 142808 329898 142860
rect 116854 142740 116860 142792
rect 116912 142780 116918 142792
rect 126054 142780 126060 142792
rect 116912 142752 126060 142780
rect 116912 142740 116918 142752
rect 126054 142740 126060 142752
rect 126112 142740 126118 142792
rect 120902 142672 120908 142724
rect 120960 142712 120966 142724
rect 127066 142712 127072 142724
rect 120960 142684 127072 142712
rect 120960 142672 120966 142684
rect 127066 142672 127072 142684
rect 127124 142672 127130 142724
rect 186038 142604 186044 142656
rect 186096 142644 186102 142656
rect 186222 142644 186228 142656
rect 186096 142616 186228 142644
rect 186096 142604 186102 142616
rect 186222 142604 186228 142616
rect 186280 142604 186286 142656
rect 179322 142468 179328 142520
rect 179380 142508 179386 142520
rect 187602 142508 187608 142520
rect 179380 142480 187608 142508
rect 179380 142468 179386 142480
rect 187602 142468 187608 142480
rect 187660 142468 187666 142520
rect 176378 142400 176384 142452
rect 176436 142440 176442 142452
rect 189626 142440 189632 142452
rect 176436 142412 189632 142440
rect 176436 142400 176442 142412
rect 189626 142400 189632 142412
rect 189684 142440 189690 142452
rect 189994 142440 190000 142452
rect 189684 142412 190000 142440
rect 189684 142400 189690 142412
rect 189994 142400 190000 142412
rect 190052 142400 190058 142452
rect 149974 142332 149980 142384
rect 150032 142372 150038 142384
rect 188982 142372 188988 142384
rect 150032 142344 188988 142372
rect 150032 142332 150038 142344
rect 188982 142332 188988 142344
rect 189040 142332 189046 142384
rect 144914 142264 144920 142316
rect 144972 142304 144978 142316
rect 145374 142304 145380 142316
rect 144972 142276 145380 142304
rect 144972 142264 144978 142276
rect 145374 142264 145380 142276
rect 145432 142304 145438 142316
rect 518894 142304 518900 142316
rect 145432 142276 518900 142304
rect 145432 142264 145438 142276
rect 518894 142264 518900 142276
rect 518952 142264 518958 142316
rect 120626 142196 120632 142248
rect 120684 142236 120690 142248
rect 122834 142236 122840 142248
rect 120684 142208 122840 142236
rect 120684 142196 120690 142208
rect 122834 142196 122840 142208
rect 122892 142196 122898 142248
rect 143534 142196 143540 142248
rect 143592 142236 143598 142248
rect 150894 142236 150900 142248
rect 143592 142208 150900 142236
rect 143592 142196 143598 142208
rect 150894 142196 150900 142208
rect 150952 142196 150958 142248
rect 161382 142196 161388 142248
rect 161440 142236 161446 142248
rect 168834 142236 168840 142248
rect 161440 142208 168840 142236
rect 161440 142196 161446 142208
rect 168834 142196 168840 142208
rect 168892 142196 168898 142248
rect 187418 142196 187424 142248
rect 187476 142236 187482 142248
rect 580258 142236 580264 142248
rect 187476 142208 580264 142236
rect 187476 142196 187482 142208
rect 580258 142196 580264 142208
rect 580316 142196 580322 142248
rect 97902 142128 97908 142180
rect 97960 142168 97966 142180
rect 113266 142168 113272 142180
rect 97960 142140 113272 142168
rect 97960 142128 97966 142140
rect 113266 142128 113272 142140
rect 113324 142128 113330 142180
rect 118602 142128 118608 142180
rect 118660 142168 118666 142180
rect 123662 142168 123668 142180
rect 118660 142140 123668 142168
rect 118660 142128 118666 142140
rect 123662 142128 123668 142140
rect 123720 142128 123726 142180
rect 148962 142168 148968 142180
rect 148875 142140 148968 142168
rect 148962 142128 148968 142140
rect 149020 142168 149026 142180
rect 580718 142168 580724 142180
rect 149020 142140 580724 142168
rect 149020 142128 149026 142140
rect 580718 142128 580724 142140
rect 580776 142128 580782 142180
rect 117222 142060 117228 142112
rect 117280 142100 117286 142112
rect 117280 142072 118694 142100
rect 117280 142060 117286 142072
rect 118666 142032 118694 142072
rect 119798 142060 119804 142112
rect 119856 142100 119862 142112
rect 148980 142100 149008 142128
rect 119856 142072 149008 142100
rect 119856 142060 119862 142072
rect 183002 142060 183008 142112
rect 183060 142100 183066 142112
rect 197446 142100 197452 142112
rect 183060 142072 197452 142100
rect 183060 142060 183066 142072
rect 197446 142060 197452 142072
rect 197504 142060 197510 142112
rect 544378 142060 544384 142112
rect 544436 142100 544442 142112
rect 580166 142100 580172 142112
rect 544436 142072 580172 142100
rect 544436 142060 544442 142072
rect 580166 142060 580172 142072
rect 580224 142060 580230 142112
rect 143534 142032 143540 142044
rect 118666 142004 128354 142032
rect 116578 141924 116584 141976
rect 116636 141964 116642 141976
rect 126238 141964 126244 141976
rect 116636 141936 126244 141964
rect 116636 141924 116642 141936
rect 126238 141924 126244 141936
rect 126296 141924 126302 141976
rect 128326 141964 128354 142004
rect 132466 142004 143540 142032
rect 132466 141964 132494 142004
rect 143534 141992 143540 142004
rect 143592 141992 143598 142044
rect 128326 141936 132494 141964
rect 180058 141924 180064 141976
rect 180116 141964 180122 141976
rect 196158 141964 196164 141976
rect 180116 141936 196164 141964
rect 180116 141924 180122 141936
rect 196158 141924 196164 141936
rect 196216 141924 196222 141976
rect 112898 141856 112904 141908
rect 112956 141896 112962 141908
rect 127802 141896 127808 141908
rect 112956 141868 127808 141896
rect 112956 141856 112962 141868
rect 127802 141856 127808 141868
rect 127860 141856 127866 141908
rect 173158 141856 173164 141908
rect 173216 141896 173222 141908
rect 185578 141896 185584 141908
rect 173216 141868 185584 141896
rect 173216 141856 173222 141868
rect 185578 141856 185584 141868
rect 185636 141856 185642 141908
rect 187602 141856 187608 141908
rect 187660 141896 187666 141908
rect 198918 141896 198924 141908
rect 187660 141868 198924 141896
rect 187660 141856 187666 141868
rect 198918 141856 198924 141868
rect 198976 141856 198982 141908
rect 113266 141788 113272 141840
rect 113324 141828 113330 141840
rect 113910 141828 113916 141840
rect 113324 141800 113916 141828
rect 113324 141788 113330 141800
rect 113910 141788 113916 141800
rect 113968 141828 113974 141840
rect 144270 141828 144276 141840
rect 113968 141800 144276 141828
rect 113968 141788 113974 141800
rect 144270 141788 144276 141800
rect 144328 141788 144334 141840
rect 174630 141788 174636 141840
rect 174688 141828 174694 141840
rect 194870 141828 194876 141840
rect 174688 141800 194876 141828
rect 174688 141788 174694 141800
rect 194870 141788 194876 141800
rect 194928 141788 194934 141840
rect 117038 141720 117044 141772
rect 117096 141760 117102 141772
rect 148594 141760 148600 141772
rect 117096 141732 148600 141760
rect 117096 141720 117102 141732
rect 148594 141720 148600 141732
rect 148652 141720 148658 141772
rect 165338 141720 165344 141772
rect 165396 141760 165402 141772
rect 199194 141760 199200 141772
rect 165396 141732 199200 141760
rect 165396 141720 165402 141732
rect 199194 141720 199200 141732
rect 199252 141720 199258 141772
rect 118326 141652 118332 141704
rect 118384 141692 118390 141704
rect 151998 141692 152004 141704
rect 118384 141664 152004 141692
rect 118384 141652 118390 141664
rect 151998 141652 152004 141664
rect 152056 141692 152062 141704
rect 153010 141692 153016 141704
rect 152056 141664 153016 141692
rect 152056 141652 152062 141664
rect 153010 141652 153016 141664
rect 153068 141652 153074 141704
rect 155586 141652 155592 141704
rect 155644 141692 155650 141704
rect 189626 141692 189632 141704
rect 155644 141664 189632 141692
rect 155644 141652 155650 141664
rect 189626 141652 189632 141664
rect 189684 141652 189690 141704
rect 115566 141584 115572 141636
rect 115624 141624 115630 141636
rect 149146 141624 149152 141636
rect 115624 141596 149152 141624
rect 115624 141584 115630 141596
rect 149146 141584 149152 141596
rect 149204 141584 149210 141636
rect 153102 141584 153108 141636
rect 153160 141624 153166 141636
rect 188890 141624 188896 141636
rect 153160 141596 188896 141624
rect 153160 141584 153166 141596
rect 188890 141584 188896 141596
rect 188948 141584 188954 141636
rect 98638 141516 98644 141568
rect 98696 141556 98702 141568
rect 158438 141556 158444 141568
rect 98696 141528 158444 141556
rect 98696 141516 98702 141528
rect 158438 141516 158444 141528
rect 158496 141516 158502 141568
rect 163958 141516 163964 141568
rect 164016 141556 164022 141568
rect 197906 141556 197912 141568
rect 164016 141528 197912 141556
rect 164016 141516 164022 141528
rect 197906 141516 197912 141528
rect 197964 141516 197970 141568
rect 198918 141516 198924 141568
rect 198976 141556 198982 141568
rect 213178 141556 213184 141568
rect 198976 141528 213184 141556
rect 198976 141516 198982 141528
rect 213178 141516 213184 141528
rect 213236 141516 213242 141568
rect 97258 141448 97264 141500
rect 97316 141488 97322 141500
rect 138566 141488 138572 141500
rect 97316 141460 138572 141488
rect 97316 141448 97322 141460
rect 138566 141448 138572 141460
rect 138624 141448 138630 141500
rect 154022 141448 154028 141500
rect 154080 141488 154086 141500
rect 218514 141488 218520 141500
rect 154080 141460 218520 141488
rect 154080 141448 154086 141460
rect 218514 141448 218520 141460
rect 218572 141448 218578 141500
rect 3602 141380 3608 141432
rect 3660 141420 3666 141432
rect 113634 141420 113640 141432
rect 3660 141392 113640 141420
rect 3660 141380 3666 141392
rect 113634 141380 113640 141392
rect 113692 141380 113698 141432
rect 119338 141380 119344 141432
rect 119396 141420 119402 141432
rect 133690 141420 133696 141432
rect 119396 141392 133696 141420
rect 119396 141380 119402 141392
rect 133690 141380 133696 141392
rect 133748 141380 133754 141432
rect 141234 141380 141240 141432
rect 141292 141420 141298 141432
rect 580350 141420 580356 141432
rect 141292 141392 580356 141420
rect 141292 141380 141298 141392
rect 580350 141380 580356 141392
rect 580408 141380 580414 141432
rect 171778 141312 171784 141364
rect 171836 141352 171842 141364
rect 186406 141352 186412 141364
rect 171836 141324 186412 141352
rect 171836 141312 171842 141324
rect 186406 141312 186412 141324
rect 186464 141312 186470 141364
rect 119246 141244 119252 141296
rect 119304 141284 119310 141296
rect 126330 141284 126336 141296
rect 119304 141256 126336 141284
rect 119304 141244 119310 141256
rect 126330 141244 126336 141256
rect 126388 141244 126394 141296
rect 181898 141244 181904 141296
rect 181956 141284 181962 141296
rect 196618 141284 196624 141296
rect 181956 141256 196624 141284
rect 181956 141244 181962 141256
rect 196618 141244 196624 141256
rect 196676 141244 196682 141296
rect 174722 141176 174728 141228
rect 174780 141216 174786 141228
rect 190730 141216 190736 141228
rect 174780 141188 190736 141216
rect 174780 141176 174786 141188
rect 190730 141176 190736 141188
rect 190788 141176 190794 141228
rect 185578 141108 185584 141160
rect 185636 141148 185642 141160
rect 192202 141148 192208 141160
rect 185636 141120 192208 141148
rect 185636 141108 185642 141120
rect 192202 141108 192208 141120
rect 192260 141108 192266 141160
rect 118666 140916 132494 140944
rect 113174 140836 113180 140888
rect 113232 140876 113238 140888
rect 117222 140876 117228 140888
rect 113232 140848 117228 140876
rect 113232 140836 113238 140848
rect 117222 140836 117228 140848
rect 117280 140836 117286 140888
rect 108114 140768 108120 140820
rect 108172 140808 108178 140820
rect 118666 140808 118694 140916
rect 108172 140780 118694 140808
rect 132466 140808 132494 140916
rect 153010 140836 153016 140888
rect 153068 140876 153074 140888
rect 211798 140876 211804 140888
rect 153068 140848 211804 140876
rect 153068 140836 153074 140848
rect 211798 140836 211804 140848
rect 211856 140836 211862 140888
rect 174630 140808 174636 140820
rect 132466 140780 174636 140808
rect 108172 140768 108178 140780
rect 174630 140768 174636 140780
rect 174688 140768 174694 140820
rect 179414 140768 179420 140820
rect 179472 140808 179478 140820
rect 179874 140808 179880 140820
rect 179472 140780 179880 140808
rect 179472 140768 179478 140780
rect 179874 140768 179880 140780
rect 179932 140768 179938 140820
rect 180794 140768 180800 140820
rect 180852 140808 180858 140820
rect 181530 140808 181536 140820
rect 180852 140780 181536 140808
rect 180852 140768 180858 140780
rect 181530 140768 181536 140780
rect 181588 140768 181594 140820
rect 187694 140768 187700 140820
rect 187752 140808 187758 140820
rect 188246 140808 188252 140820
rect 187752 140780 188252 140808
rect 187752 140768 187758 140780
rect 188246 140768 188252 140780
rect 188304 140768 188310 140820
rect 119890 140700 119896 140752
rect 119948 140740 119954 140752
rect 124306 140740 124312 140752
rect 119948 140712 124312 140740
rect 119948 140700 119954 140712
rect 124306 140700 124312 140712
rect 124364 140700 124370 140752
rect 168834 140700 168840 140752
rect 168892 140740 168898 140752
rect 193398 140740 193404 140752
rect 168892 140712 193404 140740
rect 168892 140700 168898 140712
rect 193398 140700 193404 140712
rect 193456 140700 193462 140752
rect 2774 140632 2780 140684
rect 2832 140672 2838 140684
rect 4890 140672 4896 140684
rect 2832 140644 4896 140672
rect 2832 140632 2838 140644
rect 4890 140632 4896 140644
rect 4948 140632 4954 140684
rect 115198 140632 115204 140684
rect 115256 140672 115262 140684
rect 126422 140672 126428 140684
rect 115256 140644 126428 140672
rect 115256 140632 115262 140644
rect 126422 140632 126428 140644
rect 126480 140632 126486 140684
rect 182818 140632 182824 140684
rect 182876 140672 182882 140684
rect 183094 140672 183100 140684
rect 182876 140644 183100 140672
rect 182876 140632 182882 140644
rect 183094 140632 183100 140644
rect 183152 140632 183158 140684
rect 187326 140632 187332 140684
rect 187384 140672 187390 140684
rect 193766 140672 193772 140684
rect 187384 140644 193772 140672
rect 187384 140632 187390 140644
rect 193766 140632 193772 140644
rect 193824 140632 193830 140684
rect 120810 140564 120816 140616
rect 120868 140604 120874 140616
rect 134334 140604 134340 140616
rect 120868 140576 134340 140604
rect 120868 140564 120874 140576
rect 134334 140564 134340 140576
rect 134392 140564 134398 140616
rect 182910 140564 182916 140616
rect 182968 140604 182974 140616
rect 192478 140604 192484 140616
rect 182968 140576 192484 140604
rect 182968 140564 182974 140576
rect 192478 140564 192484 140576
rect 192536 140564 192542 140616
rect 115382 140496 115388 140548
rect 115440 140536 115446 140548
rect 131666 140536 131672 140548
rect 115440 140508 131672 140536
rect 115440 140496 115446 140508
rect 131666 140496 131672 140508
rect 131724 140496 131730 140548
rect 176562 140496 176568 140548
rect 176620 140536 176626 140548
rect 186314 140536 186320 140548
rect 176620 140508 186320 140536
rect 176620 140496 176626 140508
rect 186314 140496 186320 140508
rect 186372 140496 186378 140548
rect 189810 140536 189816 140548
rect 186424 140508 189816 140536
rect 112346 140428 112352 140480
rect 112404 140468 112410 140480
rect 131942 140468 131948 140480
rect 112404 140440 131948 140468
rect 112404 140428 112410 140440
rect 131942 140428 131948 140440
rect 132000 140428 132006 140480
rect 177850 140428 177856 140480
rect 177908 140468 177914 140480
rect 186424 140468 186452 140508
rect 189810 140496 189816 140508
rect 189868 140496 189874 140548
rect 177908 140440 186452 140468
rect 177908 140428 177914 140440
rect 187786 140428 187792 140480
rect 187844 140468 187850 140480
rect 188706 140468 188712 140480
rect 187844 140440 188712 140468
rect 187844 140428 187850 140440
rect 188706 140428 188712 140440
rect 188764 140428 188770 140480
rect 115290 140360 115296 140412
rect 115348 140400 115354 140412
rect 144178 140400 144184 140412
rect 115348 140372 144184 140400
rect 115348 140360 115354 140372
rect 144178 140360 144184 140372
rect 144236 140360 144242 140412
rect 178954 140360 178960 140412
rect 179012 140400 179018 140412
rect 193490 140400 193496 140412
rect 179012 140372 193496 140400
rect 179012 140360 179018 140372
rect 193490 140360 193496 140372
rect 193548 140360 193554 140412
rect 119706 140292 119712 140344
rect 119764 140332 119770 140344
rect 150066 140332 150072 140344
rect 119764 140304 150072 140332
rect 119764 140292 119770 140304
rect 150066 140292 150072 140304
rect 150124 140292 150130 140344
rect 178678 140292 178684 140344
rect 178736 140332 178742 140344
rect 197814 140332 197820 140344
rect 178736 140304 197820 140332
rect 178736 140292 178742 140304
rect 197814 140292 197820 140304
rect 197872 140292 197878 140344
rect 112530 140224 112536 140276
rect 112588 140264 112594 140276
rect 142798 140264 142804 140276
rect 112588 140236 142804 140264
rect 112588 140224 112594 140236
rect 142798 140224 142804 140236
rect 142856 140224 142862 140276
rect 172054 140224 172060 140276
rect 172112 140264 172118 140276
rect 198090 140264 198096 140276
rect 172112 140236 198096 140264
rect 172112 140224 172118 140236
rect 198090 140224 198096 140236
rect 198148 140224 198154 140276
rect 112622 140156 112628 140208
rect 112680 140196 112686 140208
rect 145466 140196 145472 140208
rect 112680 140168 145472 140196
rect 112680 140156 112686 140168
rect 145466 140156 145472 140168
rect 145524 140156 145530 140208
rect 158530 140156 158536 140208
rect 158588 140196 158594 140208
rect 193674 140196 193680 140208
rect 158588 140168 193680 140196
rect 158588 140156 158594 140168
rect 193674 140156 193680 140168
rect 193732 140156 193738 140208
rect 114002 140088 114008 140140
rect 114060 140128 114066 140140
rect 130470 140128 130476 140140
rect 114060 140100 130476 140128
rect 114060 140088 114066 140100
rect 130470 140088 130476 140100
rect 130528 140088 130534 140140
rect 131022 140088 131028 140140
rect 131080 140128 131086 140140
rect 194962 140128 194968 140140
rect 131080 140100 194968 140128
rect 131080 140088 131086 140100
rect 194962 140088 194968 140100
rect 195020 140088 195026 140140
rect 150986 140060 150992 140072
rect 132466 140032 150992 140060
rect 116854 139952 116860 140004
rect 116912 139992 116918 140004
rect 132466 139992 132494 140032
rect 150986 140020 150992 140032
rect 151044 140020 151050 140072
rect 159634 140020 159640 140072
rect 159692 140060 159698 140072
rect 159692 140032 180794 140060
rect 159692 140020 159698 140032
rect 116912 139964 132494 139992
rect 180766 139992 180794 140032
rect 186314 140020 186320 140072
rect 186372 140060 186378 140072
rect 187326 140060 187332 140072
rect 186372 140032 187332 140060
rect 186372 140020 186378 140032
rect 187326 140020 187332 140032
rect 187384 140020 187390 140072
rect 193398 140020 193404 140072
rect 193456 140060 193462 140072
rect 492674 140060 492680 140072
rect 193456 140032 492680 140060
rect 193456 140020 193462 140032
rect 492674 140020 492680 140032
rect 492732 140020 492738 140072
rect 190546 139992 190552 140004
rect 180766 139964 190552 139992
rect 116912 139952 116918 139964
rect 190546 139952 190552 139964
rect 190604 139952 190610 140004
rect 113910 139884 113916 139936
rect 113968 139924 113974 139936
rect 124858 139924 124864 139936
rect 113968 139896 124864 139924
rect 113968 139884 113974 139896
rect 124858 139884 124864 139896
rect 124916 139884 124922 139936
rect 185670 139884 185676 139936
rect 185728 139924 185734 139936
rect 191190 139924 191196 139936
rect 185728 139896 191196 139924
rect 185728 139884 185734 139896
rect 191190 139884 191196 139896
rect 191248 139884 191254 139936
rect 185762 139816 185768 139868
rect 185820 139856 185826 139868
rect 192570 139856 192576 139868
rect 185820 139828 192576 139856
rect 185820 139816 185826 139828
rect 192570 139816 192576 139828
rect 192628 139816 192634 139868
rect 133690 139476 133696 139528
rect 133748 139516 133754 139528
rect 288434 139516 288440 139528
rect 133748 139488 288440 139516
rect 133748 139476 133754 139488
rect 288434 139476 288440 139488
rect 288492 139476 288498 139528
rect 4798 139408 4804 139460
rect 4856 139448 4862 139460
rect 182542 139448 182548 139460
rect 4856 139420 182548 139448
rect 4856 139408 4862 139420
rect 182542 139408 182548 139420
rect 182600 139408 182606 139460
rect 188154 139340 188160 139392
rect 188212 139380 188218 139392
rect 189902 139380 189908 139392
rect 188212 139352 189908 139380
rect 188212 139340 188218 139352
rect 189902 139340 189908 139352
rect 189960 139340 189966 139392
rect 111242 139272 111248 139324
rect 111300 139312 111306 139324
rect 123202 139312 123208 139324
rect 111300 139284 123208 139312
rect 111300 139272 111306 139284
rect 123202 139272 123208 139284
rect 123260 139272 123266 139324
rect 186406 139272 186412 139324
rect 186464 139312 186470 139324
rect 194042 139312 194048 139324
rect 186464 139284 194048 139312
rect 186464 139272 186470 139284
rect 194042 139272 194048 139284
rect 194100 139272 194106 139324
rect 192754 138796 192760 138848
rect 192812 138836 192818 138848
rect 200850 138836 200856 138848
rect 192812 138808 200856 138836
rect 192812 138796 192818 138808
rect 200850 138796 200856 138808
rect 200908 138796 200914 138848
rect 189902 138728 189908 138780
rect 189960 138768 189966 138780
rect 197446 138768 197452 138780
rect 189960 138740 197452 138768
rect 189960 138728 189966 138740
rect 197446 138728 197452 138740
rect 197504 138728 197510 138780
rect 188982 138660 188988 138712
rect 189040 138700 189046 138712
rect 511994 138700 512000 138712
rect 189040 138672 512000 138700
rect 189040 138660 189046 138672
rect 511994 138660 512000 138672
rect 512052 138660 512058 138712
rect 195422 137640 195428 137692
rect 195480 137680 195486 137692
rect 199562 137680 199568 137692
rect 195480 137652 199568 137680
rect 195480 137640 195486 137652
rect 199562 137640 199568 137652
rect 199620 137640 199626 137692
rect 191374 137300 191380 137352
rect 191432 137340 191438 137352
rect 203702 137340 203708 137352
rect 191432 137312 203708 137340
rect 191432 137300 191438 137312
rect 203702 137300 203708 137312
rect 203760 137300 203766 137352
rect 108206 137232 108212 137284
rect 108264 137272 108270 137284
rect 120166 137272 120172 137284
rect 108264 137244 120172 137272
rect 108264 137232 108270 137244
rect 120166 137232 120172 137244
rect 120224 137232 120230 137284
rect 189994 137232 190000 137284
rect 190052 137272 190058 137284
rect 416774 137272 416780 137284
rect 190052 137244 416780 137272
rect 190052 137232 190058 137244
rect 416774 137232 416780 137244
rect 416832 137232 416838 137284
rect 3510 136552 3516 136604
rect 3568 136592 3574 136604
rect 104066 136592 104072 136604
rect 3568 136564 104072 136592
rect 3568 136552 3574 136564
rect 104066 136552 104072 136564
rect 104124 136552 104130 136604
rect 188890 133832 188896 133884
rect 188948 133832 188954 133884
rect 188908 133680 188936 133832
rect 188890 133628 188896 133680
rect 188948 133628 188954 133680
rect 196710 133152 196716 133204
rect 196768 133192 196774 133204
rect 216122 133192 216128 133204
rect 196768 133164 216128 133192
rect 196768 133152 196774 133164
rect 216122 133152 216128 133164
rect 216180 133152 216186 133204
rect 216122 132472 216128 132524
rect 216180 132512 216186 132524
rect 579798 132512 579804 132524
rect 216180 132484 579804 132512
rect 216180 132472 216186 132484
rect 579798 132472 579804 132484
rect 579856 132472 579862 132524
rect 3326 132404 3332 132456
rect 3384 132444 3390 132456
rect 105354 132444 105360 132456
rect 3384 132416 105360 132444
rect 3384 132404 3390 132416
rect 105354 132404 105360 132416
rect 105412 132404 105418 132456
rect 3418 127576 3424 127628
rect 3476 127616 3482 127628
rect 117958 127616 117964 127628
rect 3476 127588 117964 127616
rect 3476 127576 3482 127588
rect 117958 127576 117964 127588
rect 118016 127576 118022 127628
rect 3418 122816 3424 122868
rect 3476 122856 3482 122868
rect 117866 122856 117872 122868
rect 3476 122828 117872 122856
rect 3476 122816 3482 122828
rect 117866 122816 117872 122828
rect 117924 122816 117930 122868
rect 3326 120028 3332 120080
rect 3384 120068 3390 120080
rect 95786 120068 95792 120080
rect 3384 120040 95792 120068
rect 3384 120028 3390 120040
rect 95786 120028 95792 120040
rect 95844 120028 95850 120080
rect 3418 116560 3424 116612
rect 3476 116600 3482 116612
rect 120626 116600 120632 116612
rect 3476 116572 120632 116600
rect 3476 116560 3482 116572
rect 120626 116560 120632 116572
rect 120684 116560 120690 116612
rect 3326 111800 3332 111852
rect 3384 111840 3390 111852
rect 116946 111840 116952 111852
rect 3384 111812 116952 111840
rect 3384 111800 3390 111812
rect 116946 111800 116952 111812
rect 117004 111800 117010 111852
rect 116486 110576 116492 110628
rect 116544 110616 116550 110628
rect 120626 110616 120632 110628
rect 116544 110588 120632 110616
rect 116544 110576 116550 110588
rect 120626 110576 120632 110588
rect 120684 110576 120690 110628
rect 3050 108944 3056 108996
rect 3108 108984 3114 108996
rect 100754 108984 100760 108996
rect 3108 108956 100760 108984
rect 3108 108944 3114 108956
rect 100754 108944 100760 108956
rect 100812 108984 100818 108996
rect 101306 108984 101312 108996
rect 100812 108956 101312 108984
rect 100812 108944 100818 108956
rect 101306 108944 101312 108956
rect 101364 108944 101370 108996
rect 100754 108264 100760 108316
rect 100812 108304 100818 108316
rect 111150 108304 111156 108316
rect 100812 108276 111156 108304
rect 100812 108264 100818 108276
rect 111150 108264 111156 108276
rect 111208 108264 111214 108316
rect 200942 107652 200948 107704
rect 201000 107692 201006 107704
rect 580166 107692 580172 107704
rect 201000 107664 580172 107692
rect 201000 107652 201006 107664
rect 580166 107652 580172 107664
rect 580224 107652 580230 107704
rect 2958 104796 2964 104848
rect 3016 104836 3022 104848
rect 110414 104836 110420 104848
rect 3016 104808 110420 104836
rect 3016 104796 3022 104808
rect 110414 104796 110420 104808
rect 110472 104836 110478 104848
rect 110966 104836 110972 104848
rect 110472 104808 110972 104836
rect 110472 104796 110478 104808
rect 110966 104796 110972 104808
rect 111024 104796 111030 104848
rect 110414 104116 110420 104168
rect 110472 104156 110478 104168
rect 119154 104156 119160 104168
rect 110472 104128 119160 104156
rect 110472 104116 110478 104128
rect 119154 104116 119160 104128
rect 119212 104116 119218 104168
rect 2866 99356 2872 99408
rect 2924 99396 2930 99408
rect 105354 99396 105360 99408
rect 2924 99368 105360 99396
rect 2924 99356 2930 99368
rect 105354 99356 105360 99368
rect 105412 99356 105418 99408
rect 111610 95888 111616 95940
rect 111668 95928 111674 95940
rect 119246 95928 119252 95940
rect 111668 95900 119252 95928
rect 111668 95888 111674 95900
rect 119246 95888 119252 95900
rect 119304 95888 119310 95940
rect 2958 95208 2964 95260
rect 3016 95248 3022 95260
rect 116394 95248 116400 95260
rect 3016 95220 116400 95248
rect 3016 95208 3022 95220
rect 116394 95208 116400 95220
rect 116452 95208 116458 95260
rect 112254 94732 112260 94784
rect 112312 94772 112318 94784
rect 115014 94772 115020 94784
rect 112312 94744 115020 94772
rect 112312 94732 112318 94744
rect 115014 94732 115020 94744
rect 115072 94732 115078 94784
rect 110966 93100 110972 93152
rect 111024 93140 111030 93152
rect 120718 93140 120724 93152
rect 111024 93112 120724 93140
rect 111024 93100 111030 93112
rect 120718 93100 120724 93112
rect 120776 93100 120782 93152
rect 3050 91060 3056 91112
rect 3108 91100 3114 91112
rect 97166 91100 97172 91112
rect 3108 91072 97172 91100
rect 3108 91060 3114 91072
rect 97166 91060 97172 91072
rect 97224 91060 97230 91112
rect 189718 88340 189724 88392
rect 189776 88380 189782 88392
rect 189902 88380 189908 88392
rect 189776 88352 189908 88380
rect 189776 88340 189782 88352
rect 189902 88340 189908 88352
rect 189960 88340 189966 88392
rect 3510 88272 3516 88324
rect 3568 88312 3574 88324
rect 108114 88312 108120 88324
rect 3568 88284 108120 88312
rect 3568 88272 3574 88284
rect 108114 88272 108120 88284
rect 108172 88272 108178 88324
rect 189534 86708 189540 86760
rect 189592 86748 189598 86760
rect 190178 86748 190184 86760
rect 189592 86720 190184 86748
rect 189592 86708 189598 86720
rect 190178 86708 190184 86720
rect 190236 86708 190242 86760
rect 189350 86572 189356 86624
rect 189408 86612 189414 86624
rect 189534 86612 189540 86624
rect 189408 86584 189540 86612
rect 189408 86572 189414 86584
rect 189534 86572 189540 86584
rect 189592 86572 189598 86624
rect 189166 86436 189172 86488
rect 189224 86476 189230 86488
rect 189350 86476 189356 86488
rect 189224 86448 189356 86476
rect 189224 86436 189230 86448
rect 189350 86436 189356 86448
rect 189408 86436 189414 86488
rect 189074 84872 189080 84924
rect 189132 84912 189138 84924
rect 189718 84912 189724 84924
rect 189132 84884 189724 84912
rect 189132 84872 189138 84884
rect 189718 84872 189724 84884
rect 189776 84872 189782 84924
rect 97626 83172 97632 83224
rect 97684 83212 97690 83224
rect 98638 83212 98644 83224
rect 97684 83184 98644 83212
rect 97684 83172 97690 83184
rect 98638 83172 98644 83184
rect 98696 83172 98702 83224
rect 3510 82832 3516 82884
rect 3568 82872 3574 82884
rect 97626 82872 97632 82884
rect 3568 82844 97632 82872
rect 3568 82832 3574 82844
rect 97626 82832 97632 82844
rect 97684 82832 97690 82884
rect 111610 82084 111616 82136
rect 111668 82124 111674 82136
rect 117406 82124 117412 82136
rect 111668 82096 117412 82124
rect 111668 82084 111674 82096
rect 117406 82084 117412 82096
rect 117464 82084 117470 82136
rect 140746 81688 143534 81716
rect 104066 81472 104072 81524
rect 104124 81472 104130 81524
rect 104084 81252 104112 81472
rect 119706 81336 119712 81388
rect 119764 81376 119770 81388
rect 121638 81376 121644 81388
rect 119764 81348 121644 81376
rect 119764 81336 119770 81348
rect 121638 81336 121644 81348
rect 121696 81336 121702 81388
rect 140746 81376 140774 81688
rect 143506 81512 143534 81688
rect 143506 81484 144914 81512
rect 144886 81444 144914 81484
rect 144886 81416 146294 81444
rect 132052 81348 140774 81376
rect 143506 81348 144914 81376
rect 104066 81200 104072 81252
rect 104124 81200 104130 81252
rect 113726 81064 113732 81116
rect 113784 81104 113790 81116
rect 121546 81104 121552 81116
rect 113784 81076 121552 81104
rect 113784 81064 113790 81076
rect 121546 81064 121552 81076
rect 121604 81064 121610 81116
rect 132052 81036 132080 81348
rect 143506 81308 143534 81348
rect 131868 81008 132080 81036
rect 140746 81280 143534 81308
rect 118666 80940 131252 80968
rect 116578 80860 116584 80912
rect 116636 80900 116642 80912
rect 118666 80900 118694 80940
rect 116636 80872 118694 80900
rect 123680 80872 128354 80900
rect 116636 80860 116642 80872
rect 118510 80792 118516 80844
rect 118568 80832 118574 80844
rect 123680 80832 123708 80872
rect 118568 80804 123708 80832
rect 128326 80832 128354 80872
rect 131224 80832 131252 80940
rect 131868 80900 131896 81008
rect 140746 80968 140774 81280
rect 144886 81172 144914 81348
rect 146266 81240 146294 81416
rect 580166 81376 580172 81388
rect 209746 81348 580172 81376
rect 207566 81308 207572 81320
rect 186286 81280 207572 81308
rect 146266 81212 149054 81240
rect 149026 81172 149054 81212
rect 144886 81144 146294 81172
rect 149026 81144 154574 81172
rect 131776 80872 131896 80900
rect 133892 80940 140774 80968
rect 146266 80968 146294 81144
rect 146266 80940 147674 80968
rect 128326 80804 131114 80832
rect 131224 80804 131712 80832
rect 118568 80792 118574 80804
rect 95602 80656 95608 80708
rect 95660 80696 95666 80708
rect 95660 80668 119752 80696
rect 95660 80656 95666 80668
rect 115106 80588 115112 80640
rect 115164 80628 115170 80640
rect 115164 80600 118694 80628
rect 115164 80588 115170 80600
rect 118666 80492 118694 80600
rect 119724 80560 119752 80668
rect 119798 80656 119804 80708
rect 119856 80696 119862 80708
rect 123754 80696 123760 80708
rect 119856 80668 123760 80696
rect 119856 80656 119862 80668
rect 123754 80656 123760 80668
rect 123812 80656 123818 80708
rect 123938 80656 123944 80708
rect 123996 80696 124002 80708
rect 128906 80696 128912 80708
rect 123996 80668 128912 80696
rect 123996 80656 124002 80668
rect 128906 80656 128912 80668
rect 128964 80656 128970 80708
rect 131086 80696 131114 80804
rect 131684 80708 131712 80804
rect 131574 80696 131580 80708
rect 131086 80668 131580 80696
rect 131574 80656 131580 80668
rect 131632 80656 131638 80708
rect 131666 80656 131672 80708
rect 131724 80656 131730 80708
rect 121914 80588 121920 80640
rect 121972 80628 121978 80640
rect 131776 80628 131804 80872
rect 133892 80832 133920 80940
rect 131960 80804 133920 80832
rect 131960 80708 131988 80804
rect 132052 80736 142154 80764
rect 131942 80656 131948 80708
rect 132000 80656 132006 80708
rect 121972 80600 131804 80628
rect 121972 80588 121978 80600
rect 119724 80532 128354 80560
rect 124490 80492 124496 80504
rect 118666 80464 124496 80492
rect 124490 80452 124496 80464
rect 124548 80452 124554 80504
rect 128326 80492 128354 80532
rect 131666 80520 131672 80572
rect 131724 80560 131730 80572
rect 132052 80560 132080 80736
rect 132126 80656 132132 80708
rect 132184 80696 132190 80708
rect 132184 80668 137738 80696
rect 132184 80656 132190 80668
rect 132218 80588 132224 80640
rect 132276 80628 132282 80640
rect 132276 80600 137646 80628
rect 132276 80588 132282 80600
rect 131724 80532 132080 80560
rect 131724 80520 131730 80532
rect 132126 80492 132132 80504
rect 128326 80464 132132 80492
rect 132126 80452 132132 80464
rect 132184 80452 132190 80504
rect 131574 80384 131580 80436
rect 131632 80424 131638 80436
rect 131942 80424 131948 80436
rect 131632 80396 131948 80424
rect 131632 80384 131638 80396
rect 131942 80384 131948 80396
rect 132000 80384 132006 80436
rect 128170 80316 128176 80368
rect 128228 80356 128234 80368
rect 137618 80356 137646 80600
rect 137710 80560 137738 80668
rect 142126 80628 142154 80736
rect 143506 80668 144914 80696
rect 143506 80628 143534 80668
rect 137940 80600 138198 80628
rect 142126 80600 143534 80628
rect 144886 80628 144914 80668
rect 147646 80628 147674 80940
rect 144886 80600 146294 80628
rect 147646 80600 151814 80628
rect 137940 80560 137968 80600
rect 137710 80532 137968 80560
rect 138170 80492 138198 80600
rect 146266 80492 146294 80600
rect 147646 80532 149054 80560
rect 147646 80492 147674 80532
rect 138170 80464 140774 80492
rect 146266 80464 147674 80492
rect 140746 80424 140774 80464
rect 140746 80396 147398 80424
rect 128228 80328 135668 80356
rect 137618 80328 142660 80356
rect 128228 80316 128234 80328
rect 135640 80288 135668 80328
rect 135640 80260 138014 80288
rect 129918 80180 129924 80232
rect 129976 80220 129982 80232
rect 131850 80220 131856 80232
rect 129976 80192 131856 80220
rect 129976 80180 129982 80192
rect 131850 80180 131856 80192
rect 131908 80180 131914 80232
rect 132052 80192 132494 80220
rect 131758 80112 131764 80164
rect 131816 80152 131822 80164
rect 132052 80152 132080 80192
rect 131816 80124 132080 80152
rect 131816 80112 131822 80124
rect 130102 80044 130108 80096
rect 130160 80084 130166 80096
rect 131666 80084 131672 80096
rect 130160 80056 131672 80084
rect 130160 80044 130166 80056
rect 131666 80044 131672 80056
rect 131724 80044 131730 80096
rect 132466 80084 132494 80192
rect 132466 80056 137232 80084
rect 131942 80016 131948 80028
rect 122806 79988 131948 80016
rect 101674 79772 101680 79824
rect 101732 79812 101738 79824
rect 122806 79812 122834 79988
rect 131942 79976 131948 79988
rect 132000 79976 132006 80028
rect 132052 79988 134058 80016
rect 131666 79908 131672 79960
rect 131724 79948 131730 79960
rect 132052 79948 132080 79988
rect 131724 79920 132080 79948
rect 131724 79908 131730 79920
rect 132126 79908 132132 79960
rect 132184 79948 132190 79960
rect 132540 79948 132546 79960
rect 132184 79920 132546 79948
rect 132184 79908 132190 79920
rect 132540 79908 132546 79920
rect 132598 79908 132604 79960
rect 132632 79908 132638 79960
rect 132690 79908 132696 79960
rect 132908 79908 132914 79960
rect 132966 79908 132972 79960
rect 133000 79908 133006 79960
rect 133058 79908 133064 79960
rect 133184 79908 133190 79960
rect 133242 79908 133248 79960
rect 133368 79948 133374 79960
rect 133340 79908 133374 79948
rect 133426 79908 133432 79960
rect 133828 79908 133834 79960
rect 133886 79908 133892 79960
rect 133920 79908 133926 79960
rect 133978 79908 133984 79960
rect 134030 79948 134058 79988
rect 134950 79988 135162 80016
rect 134950 79948 134978 79988
rect 135134 79960 135162 79988
rect 134030 79920 134702 79948
rect 101732 79784 122834 79812
rect 125566 79852 131114 79880
rect 101732 79772 101738 79784
rect 105998 79704 106004 79756
rect 106056 79744 106062 79756
rect 125566 79744 125594 79852
rect 106056 79716 125594 79744
rect 131086 79744 131114 79852
rect 131574 79772 131580 79824
rect 131632 79812 131638 79824
rect 132650 79812 132678 79908
rect 132926 79812 132954 79908
rect 131632 79784 132678 79812
rect 132742 79784 132954 79812
rect 131632 79772 131638 79784
rect 132742 79744 132770 79784
rect 131086 79716 132770 79744
rect 106056 79704 106062 79716
rect 132862 79704 132868 79756
rect 132920 79704 132926 79756
rect 3510 79636 3516 79688
rect 3568 79676 3574 79688
rect 3568 79648 132494 79676
rect 3568 79636 3574 79648
rect 117682 79568 117688 79620
rect 117740 79608 117746 79620
rect 126238 79608 126244 79620
rect 117740 79580 126244 79608
rect 117740 79568 117746 79580
rect 126238 79568 126244 79580
rect 126296 79568 126302 79620
rect 119338 79500 119344 79552
rect 119396 79540 119402 79552
rect 127618 79540 127624 79552
rect 119396 79512 127624 79540
rect 119396 79500 119402 79512
rect 127618 79500 127624 79512
rect 127676 79500 127682 79552
rect 111150 79432 111156 79484
rect 111208 79472 111214 79484
rect 130102 79472 130108 79484
rect 111208 79444 130108 79472
rect 111208 79432 111214 79444
rect 130102 79432 130108 79444
rect 130160 79432 130166 79484
rect 132466 79472 132494 79648
rect 132880 79540 132908 79704
rect 133018 79688 133046 79908
rect 133202 79824 133230 79908
rect 133138 79772 133144 79824
rect 133196 79784 133230 79824
rect 133196 79772 133202 79784
rect 133018 79648 133052 79688
rect 133046 79636 133052 79648
rect 133104 79636 133110 79688
rect 132954 79568 132960 79620
rect 133012 79608 133018 79620
rect 133340 79608 133368 79908
rect 133846 79756 133874 79908
rect 133938 79812 133966 79908
rect 134674 79892 134702 79920
rect 134766 79920 134978 79948
rect 134288 79840 134294 79892
rect 134346 79880 134352 79892
rect 134564 79880 134570 79892
rect 134346 79840 134380 79880
rect 133938 79784 134288 79812
rect 133846 79716 133880 79756
rect 133874 79704 133880 79716
rect 133932 79704 133938 79756
rect 134260 79620 134288 79784
rect 134352 79756 134380 79840
rect 134536 79840 134570 79880
rect 134622 79840 134628 79892
rect 134656 79840 134662 79892
rect 134714 79840 134720 79892
rect 134334 79704 134340 79756
rect 134392 79704 134398 79756
rect 134536 79676 134564 79840
rect 134610 79704 134616 79756
rect 134668 79744 134674 79756
rect 134766 79744 134794 79920
rect 135024 79908 135030 79960
rect 135082 79908 135088 79960
rect 135116 79908 135122 79960
rect 135174 79908 135180 79960
rect 135208 79908 135214 79960
rect 135266 79908 135272 79960
rect 135300 79908 135306 79960
rect 135358 79908 135364 79960
rect 136220 79948 136226 79960
rect 136192 79908 136226 79948
rect 136278 79908 136284 79960
rect 136496 79948 136502 79960
rect 136468 79908 136502 79948
rect 136554 79908 136560 79960
rect 137048 79908 137054 79960
rect 137106 79908 137112 79960
rect 137204 79948 137232 80056
rect 137986 79960 138014 80260
rect 139366 80192 141050 80220
rect 139366 80016 139394 80192
rect 138400 79988 139394 80016
rect 137508 79948 137514 79960
rect 137204 79920 137514 79948
rect 137508 79908 137514 79920
rect 137566 79908 137572 79960
rect 137600 79908 137606 79960
rect 137658 79908 137664 79960
rect 137692 79908 137698 79960
rect 137750 79908 137756 79960
rect 137968 79908 137974 79960
rect 138026 79908 138032 79960
rect 138152 79908 138158 79960
rect 138210 79908 138216 79960
rect 138244 79908 138250 79960
rect 138302 79908 138308 79960
rect 134840 79840 134846 79892
rect 134898 79840 134904 79892
rect 134932 79840 134938 79892
rect 134990 79840 134996 79892
rect 134668 79716 134794 79744
rect 134668 79704 134674 79716
rect 134702 79676 134708 79688
rect 134536 79648 134708 79676
rect 134702 79636 134708 79648
rect 134760 79636 134766 79688
rect 133690 79608 133696 79620
rect 133012 79580 133368 79608
rect 133432 79580 133696 79608
rect 133012 79568 133018 79580
rect 133432 79540 133460 79580
rect 133690 79568 133696 79580
rect 133748 79568 133754 79620
rect 134242 79568 134248 79620
rect 134300 79568 134306 79620
rect 134426 79568 134432 79620
rect 134484 79608 134490 79620
rect 134858 79608 134886 79840
rect 134484 79580 134886 79608
rect 134484 79568 134490 79580
rect 134950 79552 134978 79840
rect 135042 79756 135070 79908
rect 135226 79824 135254 79908
rect 135162 79772 135168 79824
rect 135220 79784 135254 79824
rect 135220 79772 135226 79784
rect 135318 79756 135346 79908
rect 135484 79840 135490 79892
rect 135542 79880 135548 79892
rect 135542 79840 135576 79880
rect 135944 79840 135950 79892
rect 136002 79840 136008 79892
rect 136036 79840 136042 79892
rect 136094 79880 136100 79892
rect 136094 79840 136128 79880
rect 135548 79756 135576 79840
rect 135042 79716 135076 79756
rect 135070 79704 135076 79716
rect 135128 79704 135134 79756
rect 135254 79704 135260 79756
rect 135312 79716 135346 79756
rect 135312 79704 135318 79716
rect 135530 79704 135536 79756
rect 135588 79704 135594 79756
rect 135962 79688 135990 79840
rect 136100 79756 136128 79840
rect 136192 79756 136220 79908
rect 136312 79840 136318 79892
rect 136370 79880 136376 79892
rect 136370 79840 136404 79880
rect 136082 79704 136088 79756
rect 136140 79704 136146 79756
rect 136174 79704 136180 79756
rect 136232 79704 136238 79756
rect 136376 79688 136404 79840
rect 135962 79648 135996 79688
rect 135990 79636 135996 79648
rect 136048 79636 136054 79688
rect 136358 79636 136364 79688
rect 136416 79636 136422 79688
rect 135806 79568 135812 79620
rect 135864 79608 135870 79620
rect 136468 79608 136496 79908
rect 136588 79880 136594 79892
rect 136560 79840 136594 79880
rect 136646 79840 136652 79892
rect 136680 79840 136686 79892
rect 136738 79840 136744 79892
rect 136864 79840 136870 79892
rect 136922 79840 136928 79892
rect 136560 79688 136588 79840
rect 136698 79812 136726 79840
rect 136652 79784 136726 79812
rect 136652 79688 136680 79784
rect 136882 79744 136910 79840
rect 136744 79716 136910 79744
rect 137066 79756 137094 79908
rect 137232 79840 137238 79892
rect 137290 79840 137296 79892
rect 137416 79840 137422 79892
rect 137474 79840 137480 79892
rect 137066 79716 137100 79756
rect 136542 79636 136548 79688
rect 136600 79636 136606 79688
rect 136634 79636 136640 79688
rect 136692 79636 136698 79688
rect 135864 79580 136496 79608
rect 136744 79608 136772 79716
rect 137094 79704 137100 79716
rect 137152 79704 137158 79756
rect 136818 79636 136824 79688
rect 136876 79676 136882 79688
rect 137250 79676 137278 79840
rect 136876 79648 137278 79676
rect 136876 79636 136882 79648
rect 137250 79620 137278 79648
rect 137434 79620 137462 79840
rect 137618 79824 137646 79908
rect 137554 79772 137560 79824
rect 137612 79784 137646 79824
rect 137612 79772 137618 79784
rect 137710 79756 137738 79908
rect 138170 79880 138198 79908
rect 138078 79852 138198 79880
rect 138078 79824 138106 79852
rect 138014 79772 138020 79824
rect 138072 79784 138106 79824
rect 138262 79812 138290 79908
rect 138262 79784 138336 79812
rect 138072 79772 138078 79784
rect 137646 79704 137652 79756
rect 137704 79716 137738 79756
rect 137704 79704 137710 79716
rect 138106 79636 138112 79688
rect 138164 79676 138170 79688
rect 138308 79676 138336 79784
rect 138400 79688 138428 79988
rect 141022 79960 141050 80192
rect 139164 79948 139170 79960
rect 138492 79920 139170 79948
rect 138164 79648 138336 79676
rect 138164 79636 138170 79648
rect 138382 79636 138388 79688
rect 138440 79636 138446 79688
rect 137002 79608 137008 79620
rect 136744 79580 137008 79608
rect 135864 79568 135870 79580
rect 137002 79568 137008 79580
rect 137060 79568 137066 79620
rect 137250 79580 137284 79620
rect 137278 79568 137284 79580
rect 137336 79568 137342 79620
rect 137370 79568 137376 79620
rect 137428 79580 137462 79620
rect 137428 79568 137434 79580
rect 132880 79512 133460 79540
rect 134886 79500 134892 79552
rect 134944 79512 134978 79552
rect 134944 79500 134950 79512
rect 136266 79500 136272 79552
rect 136324 79540 136330 79552
rect 138492 79540 138520 79920
rect 139164 79908 139170 79920
rect 139222 79908 139228 79960
rect 139808 79908 139814 79960
rect 139866 79908 139872 79960
rect 139900 79908 139906 79960
rect 139958 79908 139964 79960
rect 139992 79908 139998 79960
rect 140050 79948 140056 79960
rect 140050 79908 140084 79948
rect 140176 79908 140182 79960
rect 140234 79908 140240 79960
rect 140268 79908 140274 79960
rect 140326 79908 140332 79960
rect 140452 79908 140458 79960
rect 140510 79908 140516 79960
rect 140636 79948 140642 79960
rect 140608 79908 140642 79948
rect 140694 79908 140700 79960
rect 140728 79908 140734 79960
rect 140786 79908 140792 79960
rect 140912 79948 140918 79960
rect 140838 79920 140918 79948
rect 138704 79840 138710 79892
rect 138762 79840 138768 79892
rect 138796 79840 138802 79892
rect 138854 79840 138860 79892
rect 138980 79840 138986 79892
rect 139038 79840 139044 79892
rect 139072 79840 139078 79892
rect 139130 79840 139136 79892
rect 139826 79880 139854 79908
rect 139320 79852 139854 79880
rect 138722 79744 138750 79840
rect 138676 79716 138750 79744
rect 138676 79608 138704 79716
rect 138814 79688 138842 79840
rect 138998 79756 139026 79840
rect 138934 79704 138940 79756
rect 138992 79716 139026 79756
rect 138992 79704 138998 79716
rect 139090 79688 139118 79840
rect 138750 79636 138756 79688
rect 138808 79648 138842 79688
rect 138808 79636 138814 79648
rect 139026 79636 139032 79688
rect 139084 79648 139118 79688
rect 139084 79636 139090 79648
rect 139210 79608 139216 79620
rect 138676 79580 139216 79608
rect 139210 79568 139216 79580
rect 139268 79568 139274 79620
rect 136324 79512 138520 79540
rect 136324 79500 136330 79512
rect 138566 79500 138572 79552
rect 138624 79540 138630 79552
rect 139320 79540 139348 79852
rect 139918 79824 139946 79908
rect 139440 79772 139446 79824
rect 139498 79772 139504 79824
rect 139918 79784 139952 79824
rect 139946 79772 139952 79784
rect 140004 79772 140010 79824
rect 139458 79620 139486 79772
rect 139854 79704 139860 79756
rect 139912 79744 139918 79756
rect 140056 79744 140084 79908
rect 139912 79716 140084 79744
rect 139912 79704 139918 79716
rect 139670 79636 139676 79688
rect 139728 79676 139734 79688
rect 140194 79676 140222 79908
rect 139728 79648 140222 79676
rect 139728 79636 139734 79648
rect 139394 79568 139400 79620
rect 139452 79580 139486 79620
rect 139452 79568 139458 79580
rect 139762 79568 139768 79620
rect 139820 79608 139826 79620
rect 140286 79608 140314 79908
rect 140470 79688 140498 79908
rect 140406 79636 140412 79688
rect 140464 79648 140498 79688
rect 140464 79636 140470 79648
rect 140608 79620 140636 79908
rect 140746 79880 140774 79908
rect 140700 79852 140774 79880
rect 140700 79756 140728 79852
rect 140838 79824 140866 79920
rect 140912 79908 140918 79920
rect 140970 79908 140976 79960
rect 141004 79908 141010 79960
rect 141062 79908 141068 79960
rect 141188 79908 141194 79960
rect 141246 79908 141252 79960
rect 141372 79908 141378 79960
rect 141430 79908 141436 79960
rect 141740 79908 141746 79960
rect 141798 79908 141804 79960
rect 141832 79908 141838 79960
rect 141890 79908 141896 79960
rect 142016 79908 142022 79960
rect 142074 79908 142080 79960
rect 142476 79948 142482 79960
rect 142126 79920 142482 79948
rect 141206 79880 141234 79908
rect 140774 79772 140780 79824
rect 140832 79784 140866 79824
rect 140976 79852 141234 79880
rect 140832 79772 140838 79784
rect 140682 79704 140688 79756
rect 140740 79704 140746 79756
rect 139820 79580 140314 79608
rect 139820 79568 139826 79580
rect 140590 79568 140596 79620
rect 140648 79568 140654 79620
rect 140976 79552 141004 79852
rect 141390 79744 141418 79908
rect 141556 79840 141562 79892
rect 141614 79840 141620 79892
rect 141160 79716 141418 79744
rect 138624 79512 139348 79540
rect 138624 79500 138630 79512
rect 140958 79500 140964 79552
rect 141016 79500 141022 79552
rect 141160 79472 141188 79716
rect 141326 79636 141332 79688
rect 141384 79676 141390 79688
rect 141574 79676 141602 79840
rect 141758 79824 141786 79908
rect 141740 79772 141746 79824
rect 141798 79772 141804 79824
rect 141384 79648 141602 79676
rect 141384 79636 141390 79648
rect 141694 79568 141700 79620
rect 141752 79608 141758 79620
rect 141850 79608 141878 79908
rect 142034 79756 142062 79908
rect 141970 79704 141976 79756
rect 142028 79716 142062 79756
rect 142028 79704 142034 79716
rect 142126 79620 142154 79920
rect 142476 79908 142482 79920
rect 142534 79908 142540 79960
rect 142200 79840 142206 79892
rect 142258 79840 142264 79892
rect 142384 79840 142390 79892
rect 142442 79840 142448 79892
rect 141752 79580 141878 79608
rect 141752 79568 141758 79580
rect 142062 79568 142068 79620
rect 142120 79580 142154 79620
rect 142120 79568 142126 79580
rect 142218 79484 142246 79840
rect 142402 79744 142430 79840
rect 142310 79716 142430 79744
rect 142310 79552 142338 79716
rect 142522 79676 142528 79688
rect 142448 79648 142528 79676
rect 142310 79512 142344 79552
rect 142338 79500 142344 79512
rect 142396 79500 142402 79552
rect 141878 79472 141884 79484
rect 132466 79444 138244 79472
rect 141160 79444 141884 79472
rect 108206 79364 108212 79416
rect 108264 79404 108270 79416
rect 134978 79404 134984 79416
rect 108264 79376 134984 79404
rect 108264 79364 108270 79376
rect 134978 79364 134984 79376
rect 135036 79364 135042 79416
rect 135346 79364 135352 79416
rect 135404 79404 135410 79416
rect 136450 79404 136456 79416
rect 135404 79376 136456 79404
rect 135404 79364 135410 79376
rect 136450 79364 136456 79376
rect 136508 79364 136514 79416
rect 138216 79404 138244 79444
rect 141878 79432 141884 79444
rect 141936 79432 141942 79484
rect 142218 79444 142252 79484
rect 142246 79432 142252 79444
rect 142304 79432 142310 79484
rect 142448 79472 142476 79648
rect 142522 79636 142528 79648
rect 142580 79636 142586 79688
rect 142632 79608 142660 80328
rect 145530 79988 146018 80016
rect 145530 79960 145558 79988
rect 142936 79908 142942 79960
rect 142994 79908 143000 79960
rect 143212 79908 143218 79960
rect 143270 79908 143276 79960
rect 143488 79908 143494 79960
rect 143546 79908 143552 79960
rect 143580 79908 143586 79960
rect 143638 79908 143644 79960
rect 143764 79948 143770 79960
rect 143690 79920 143770 79948
rect 142798 79608 142804 79620
rect 142632 79580 142804 79608
rect 142798 79568 142804 79580
rect 142856 79568 142862 79620
rect 142522 79500 142528 79552
rect 142580 79540 142586 79552
rect 142954 79540 142982 79908
rect 143120 79880 143126 79892
rect 143092 79840 143126 79880
rect 143178 79840 143184 79892
rect 143092 79756 143120 79840
rect 143230 79756 143258 79908
rect 143396 79812 143402 79824
rect 143074 79704 143080 79756
rect 143132 79704 143138 79756
rect 143166 79704 143172 79756
rect 143224 79716 143258 79756
rect 143368 79772 143402 79812
rect 143454 79772 143460 79824
rect 143224 79704 143230 79716
rect 143368 79620 143396 79772
rect 143506 79744 143534 79908
rect 143460 79716 143534 79744
rect 143460 79620 143488 79716
rect 143598 79688 143626 79908
rect 143534 79636 143540 79688
rect 143592 79648 143626 79688
rect 143592 79636 143598 79648
rect 143350 79568 143356 79620
rect 143408 79568 143414 79620
rect 143442 79568 143448 79620
rect 143500 79568 143506 79620
rect 142580 79512 142982 79540
rect 142580 79500 142586 79512
rect 142890 79472 142896 79484
rect 142448 79444 142896 79472
rect 142890 79432 142896 79444
rect 142948 79432 142954 79484
rect 143690 79472 143718 79920
rect 143764 79908 143770 79920
rect 143822 79908 143828 79960
rect 143948 79948 143954 79960
rect 143920 79908 143954 79948
rect 144006 79908 144012 79960
rect 144316 79908 144322 79960
rect 144374 79908 144380 79960
rect 144408 79908 144414 79960
rect 144466 79908 144472 79960
rect 144592 79908 144598 79960
rect 144650 79908 144656 79960
rect 144684 79908 144690 79960
rect 144742 79908 144748 79960
rect 144776 79908 144782 79960
rect 144834 79948 144840 79960
rect 144834 79908 144868 79948
rect 145236 79908 145242 79960
rect 145294 79908 145300 79960
rect 145420 79908 145426 79960
rect 145478 79908 145484 79960
rect 145512 79908 145518 79960
rect 145570 79908 145576 79960
rect 145604 79908 145610 79960
rect 145662 79908 145668 79960
rect 145880 79948 145886 79960
rect 145714 79920 145886 79948
rect 143920 79620 143948 79908
rect 144040 79880 144046 79892
rect 144012 79840 144046 79880
rect 144098 79840 144104 79892
rect 144012 79688 144040 79840
rect 144334 79812 144362 79908
rect 144104 79784 144362 79812
rect 143994 79636 144000 79688
rect 144052 79636 144058 79688
rect 144104 79620 144132 79784
rect 144270 79636 144276 79688
rect 144328 79676 144334 79688
rect 144426 79676 144454 79908
rect 144610 79688 144638 79908
rect 144702 79824 144730 79908
rect 144684 79772 144690 79824
rect 144742 79772 144748 79824
rect 144328 79648 144454 79676
rect 144328 79636 144334 79648
rect 144546 79636 144552 79688
rect 144604 79648 144638 79688
rect 144604 79636 144610 79648
rect 144730 79636 144736 79688
rect 144788 79676 144794 79688
rect 144840 79676 144868 79908
rect 144960 79840 144966 79892
rect 145018 79840 145024 79892
rect 145144 79840 145150 79892
rect 145202 79840 145208 79892
rect 144788 79648 144868 79676
rect 144788 79636 144794 79648
rect 143902 79568 143908 79620
rect 143960 79568 143966 79620
rect 144086 79568 144092 79620
rect 144144 79568 144150 79620
rect 144978 79608 145006 79840
rect 145162 79688 145190 79840
rect 145254 79744 145282 79908
rect 145438 79824 145466 79908
rect 145374 79772 145380 79824
rect 145432 79784 145466 79824
rect 145432 79772 145438 79784
rect 145622 79756 145650 79908
rect 145466 79744 145472 79756
rect 145254 79716 145472 79744
rect 145466 79704 145472 79716
rect 145524 79704 145530 79756
rect 145558 79704 145564 79756
rect 145616 79716 145650 79756
rect 145616 79704 145622 79716
rect 145162 79648 145196 79688
rect 145190 79636 145196 79648
rect 145248 79636 145254 79688
rect 145714 79676 145742 79920
rect 145880 79908 145886 79920
rect 145938 79908 145944 79960
rect 145788 79840 145794 79892
rect 145846 79840 145852 79892
rect 145806 79756 145834 79840
rect 145990 79824 146018 79988
rect 147370 79960 147398 80396
rect 149026 80016 149054 80532
rect 151786 80492 151814 80600
rect 151786 80464 152458 80492
rect 149026 79988 149698 80016
rect 149670 79960 149698 79988
rect 152430 79960 152458 80464
rect 154546 80016 154574 81144
rect 186286 81104 186314 81280
rect 207566 81268 207572 81280
rect 207624 81268 207630 81320
rect 191374 81132 191380 81184
rect 191432 81172 191438 81184
rect 198090 81172 198096 81184
rect 191432 81144 198096 81172
rect 191432 81132 191438 81144
rect 198090 81132 198096 81144
rect 198148 81132 198154 81184
rect 177776 81076 186314 81104
rect 164206 81008 172606 81036
rect 164206 80628 164234 81008
rect 172578 80628 172606 81008
rect 177776 80696 177804 81076
rect 188982 81064 188988 81116
rect 189040 81104 189046 81116
rect 209130 81104 209136 81116
rect 189040 81076 209136 81104
rect 189040 81064 189046 81076
rect 209130 81064 209136 81076
rect 209188 81064 209194 81116
rect 202414 81036 202420 81048
rect 178052 81008 202420 81036
rect 178052 80708 178080 81008
rect 202414 80996 202420 81008
rect 202472 81036 202478 81048
rect 209746 81036 209774 81348
rect 580166 81336 580172 81348
rect 580224 81336 580230 81388
rect 202472 81008 209774 81036
rect 202472 80996 202478 81008
rect 204530 80968 204536 80980
rect 183526 80940 204536 80968
rect 183526 80900 183554 80940
rect 204530 80928 204536 80940
rect 204588 80928 204594 80980
rect 178420 80872 183554 80900
rect 178420 80708 178448 80872
rect 188982 80860 188988 80912
rect 189040 80900 189046 80912
rect 219986 80900 219992 80912
rect 189040 80872 219992 80900
rect 189040 80860 189046 80872
rect 219986 80860 219992 80872
rect 220044 80860 220050 80912
rect 196618 80832 196624 80844
rect 178512 80804 196624 80832
rect 177850 80696 177856 80708
rect 177776 80668 177856 80696
rect 177850 80656 177856 80668
rect 177908 80656 177914 80708
rect 178034 80656 178040 80708
rect 178092 80656 178098 80708
rect 178402 80656 178408 80708
rect 178460 80656 178466 80708
rect 178512 80628 178540 80804
rect 196618 80792 196624 80804
rect 196676 80792 196682 80844
rect 211430 80764 211436 80776
rect 183526 80736 211436 80764
rect 162090 80600 164234 80628
rect 168300 80600 172514 80628
rect 172578 80600 178540 80628
rect 154776 80056 158530 80084
rect 154776 80016 154804 80056
rect 154546 79988 154804 80016
rect 157812 79988 158346 80016
rect 146064 79908 146070 79960
rect 146122 79908 146128 79960
rect 146156 79908 146162 79960
rect 146214 79908 146220 79960
rect 146340 79908 146346 79960
rect 146398 79908 146404 79960
rect 146800 79908 146806 79960
rect 146858 79908 146864 79960
rect 147352 79908 147358 79960
rect 147410 79908 147416 79960
rect 147444 79908 147450 79960
rect 147502 79908 147508 79960
rect 147536 79908 147542 79960
rect 147594 79908 147600 79960
rect 148088 79908 148094 79960
rect 148146 79908 148152 79960
rect 148824 79948 148830 79960
rect 148750 79920 148830 79948
rect 146082 79824 146110 79908
rect 145926 79772 145932 79824
rect 145984 79784 146018 79824
rect 145984 79772 145990 79784
rect 146064 79772 146070 79824
rect 146122 79772 146128 79824
rect 145806 79716 145840 79756
rect 145834 79704 145840 79716
rect 145892 79704 145898 79756
rect 146174 79744 146202 79908
rect 146036 79716 146202 79744
rect 145300 79648 145742 79676
rect 145300 79620 145328 79648
rect 146036 79620 146064 79716
rect 145098 79608 145104 79620
rect 144978 79580 145104 79608
rect 145098 79568 145104 79580
rect 145156 79568 145162 79620
rect 145282 79568 145288 79620
rect 145340 79568 145346 79620
rect 146018 79568 146024 79620
rect 146076 79568 146082 79620
rect 146358 79552 146386 79908
rect 146432 79840 146438 79892
rect 146490 79840 146496 79892
rect 146616 79840 146622 79892
rect 146674 79840 146680 79892
rect 146818 79880 146846 79908
rect 146772 79852 146846 79880
rect 146450 79620 146478 79840
rect 146450 79580 146484 79620
rect 146478 79568 146484 79580
rect 146536 79568 146542 79620
rect 146358 79512 146392 79552
rect 146386 79500 146392 79512
rect 146444 79500 146450 79552
rect 146634 79540 146662 79840
rect 146772 79608 146800 79852
rect 146892 79840 146898 79892
rect 146950 79840 146956 79892
rect 146984 79840 146990 79892
rect 147042 79840 147048 79892
rect 147168 79840 147174 79892
rect 147226 79840 147232 79892
rect 147260 79840 147266 79892
rect 147318 79880 147324 79892
rect 147462 79880 147490 79908
rect 147318 79840 147352 79880
rect 146910 79688 146938 79840
rect 147002 79744 147030 79840
rect 147186 79756 147214 79840
rect 147324 79756 147352 79840
rect 147416 79852 147490 79880
rect 147416 79824 147444 79852
rect 147554 79824 147582 79908
rect 147628 79840 147634 79892
rect 147686 79840 147692 79892
rect 147398 79772 147404 79824
rect 147456 79772 147462 79824
rect 147490 79772 147496 79824
rect 147548 79784 147582 79824
rect 147548 79772 147554 79784
rect 147646 79756 147674 79840
rect 147002 79716 147122 79744
rect 147186 79716 147220 79756
rect 146910 79648 146944 79688
rect 146938 79636 146944 79648
rect 146996 79636 147002 79688
rect 146846 79608 146852 79620
rect 146772 79580 146852 79608
rect 146846 79568 146852 79580
rect 146904 79568 146910 79620
rect 147094 79552 147122 79716
rect 147214 79704 147220 79716
rect 147272 79704 147278 79756
rect 147306 79704 147312 79756
rect 147364 79704 147370 79756
rect 147582 79704 147588 79756
rect 147640 79716 147674 79756
rect 147640 79704 147646 79716
rect 146754 79540 146760 79552
rect 146634 79512 146760 79540
rect 146754 79500 146760 79512
rect 146812 79500 146818 79552
rect 147030 79500 147036 79552
rect 147088 79512 147122 79552
rect 148106 79552 148134 79908
rect 148548 79840 148554 79892
rect 148606 79840 148612 79892
rect 148566 79608 148594 79840
rect 148750 79688 148778 79920
rect 148824 79908 148830 79920
rect 148882 79908 148888 79960
rect 148916 79908 148922 79960
rect 148974 79908 148980 79960
rect 149008 79908 149014 79960
rect 149066 79908 149072 79960
rect 149468 79908 149474 79960
rect 149526 79908 149532 79960
rect 149560 79908 149566 79960
rect 149618 79908 149624 79960
rect 149652 79908 149658 79960
rect 149710 79908 149716 79960
rect 150756 79908 150762 79960
rect 150814 79908 150820 79960
rect 151032 79908 151038 79960
rect 151090 79908 151096 79960
rect 151400 79908 151406 79960
rect 151458 79948 151464 79960
rect 151458 79920 151538 79948
rect 151458 79908 151464 79920
rect 148934 79880 148962 79908
rect 148888 79852 148962 79880
rect 148888 79756 148916 79852
rect 149026 79824 149054 79908
rect 148962 79772 148968 79824
rect 149020 79784 149054 79824
rect 149020 79772 149026 79784
rect 149192 79772 149198 79824
rect 149250 79772 149256 79824
rect 148870 79704 148876 79756
rect 148928 79704 148934 79756
rect 148686 79636 148692 79688
rect 148744 79648 148778 79688
rect 148744 79636 148750 79648
rect 149210 79620 149238 79772
rect 149486 79688 149514 79908
rect 149578 79756 149606 79908
rect 149744 79880 149750 79892
rect 149716 79840 149750 79880
rect 149802 79840 149808 79892
rect 149836 79840 149842 79892
rect 149894 79840 149900 79892
rect 149928 79840 149934 79892
rect 149986 79840 149992 79892
rect 150112 79840 150118 79892
rect 150170 79840 150176 79892
rect 150296 79840 150302 79892
rect 150354 79840 150360 79892
rect 150774 79880 150802 79908
rect 150544 79852 150802 79880
rect 149716 79756 149744 79840
rect 149854 79756 149882 79840
rect 149578 79716 149612 79756
rect 149606 79704 149612 79716
rect 149664 79704 149670 79756
rect 149698 79704 149704 79756
rect 149756 79704 149762 79756
rect 149790 79704 149796 79756
rect 149848 79716 149882 79756
rect 149848 79704 149854 79716
rect 149946 79688 149974 79840
rect 149486 79648 149520 79688
rect 149514 79636 149520 79648
rect 149572 79636 149578 79688
rect 149882 79636 149888 79688
rect 149940 79648 149974 79688
rect 149940 79636 149946 79648
rect 148778 79608 148784 79620
rect 148566 79580 148784 79608
rect 148778 79568 148784 79580
rect 148836 79568 148842 79620
rect 149146 79568 149152 79620
rect 149204 79580 149238 79620
rect 149204 79568 149210 79580
rect 148106 79512 148140 79552
rect 147088 79500 147094 79512
rect 148134 79500 148140 79512
rect 148192 79500 148198 79552
rect 149238 79500 149244 79552
rect 149296 79540 149302 79552
rect 150130 79540 150158 79840
rect 149296 79512 150158 79540
rect 149296 79500 149302 79512
rect 150314 79484 150342 79840
rect 150544 79484 150572 79852
rect 150664 79772 150670 79824
rect 150722 79772 150728 79824
rect 150682 79608 150710 79772
rect 151050 79608 151078 79908
rect 151308 79840 151314 79892
rect 151366 79840 151372 79892
rect 151326 79744 151354 79840
rect 151510 79824 151538 79920
rect 151584 79908 151590 79960
rect 151642 79908 151648 79960
rect 151676 79908 151682 79960
rect 151734 79908 151740 79960
rect 151860 79908 151866 79960
rect 151918 79908 151924 79960
rect 151952 79908 151958 79960
rect 152010 79948 152016 79960
rect 152010 79920 152274 79948
rect 152010 79908 152016 79920
rect 151492 79772 151498 79824
rect 151550 79772 151556 79824
rect 151326 79716 151492 79744
rect 151354 79608 151360 79620
rect 150682 79580 150756 79608
rect 151050 79580 151360 79608
rect 150728 79552 150756 79580
rect 151354 79568 151360 79580
rect 151412 79568 151418 79620
rect 150710 79500 150716 79552
rect 150768 79500 150774 79552
rect 150986 79500 150992 79552
rect 151044 79540 151050 79552
rect 151464 79540 151492 79716
rect 151602 79688 151630 79908
rect 151538 79636 151544 79688
rect 151596 79648 151630 79688
rect 151596 79636 151602 79648
rect 151694 79608 151722 79908
rect 151878 79756 151906 79908
rect 152044 79880 152050 79892
rect 152016 79840 152050 79880
rect 152102 79840 152108 79892
rect 152016 79756 152044 79840
rect 152136 79772 152142 79824
rect 152194 79772 152200 79824
rect 151878 79716 151912 79756
rect 151906 79704 151912 79716
rect 151964 79704 151970 79756
rect 151998 79704 152004 79756
rect 152056 79704 152062 79756
rect 152154 79688 152182 79772
rect 152246 79744 152274 79920
rect 152412 79908 152418 79960
rect 152470 79908 152476 79960
rect 152964 79908 152970 79960
rect 153022 79908 153028 79960
rect 153608 79908 153614 79960
rect 153666 79908 153672 79960
rect 154252 79908 154258 79960
rect 154310 79908 154316 79960
rect 154344 79908 154350 79960
rect 154402 79908 154408 79960
rect 154436 79908 154442 79960
rect 154494 79908 154500 79960
rect 154988 79948 154994 79960
rect 154960 79908 154994 79948
rect 155046 79908 155052 79960
rect 155172 79948 155178 79960
rect 155144 79908 155178 79948
rect 155230 79908 155236 79960
rect 155816 79908 155822 79960
rect 155874 79908 155880 79960
rect 156184 79908 156190 79960
rect 156242 79908 156248 79960
rect 156644 79908 156650 79960
rect 156702 79908 156708 79960
rect 156920 79908 156926 79960
rect 156978 79908 156984 79960
rect 157012 79908 157018 79960
rect 157070 79908 157076 79960
rect 157104 79908 157110 79960
rect 157162 79908 157168 79960
rect 157196 79908 157202 79960
rect 157254 79908 157260 79960
rect 157380 79948 157386 79960
rect 157352 79908 157386 79948
rect 157438 79908 157444 79960
rect 157472 79908 157478 79960
rect 157530 79908 157536 79960
rect 157656 79908 157662 79960
rect 157714 79908 157720 79960
rect 152780 79840 152786 79892
rect 152838 79840 152844 79892
rect 152458 79744 152464 79756
rect 152246 79716 152464 79744
rect 152458 79704 152464 79716
rect 152516 79704 152522 79756
rect 152090 79636 152096 79688
rect 152148 79648 152182 79688
rect 152798 79688 152826 79840
rect 152982 79744 153010 79908
rect 153240 79840 153246 79892
rect 153298 79840 153304 79892
rect 153424 79880 153430 79892
rect 153396 79840 153430 79880
rect 153482 79840 153488 79892
rect 153056 79772 153062 79824
rect 153114 79812 153120 79824
rect 153114 79784 153194 79812
rect 153114 79772 153120 79784
rect 152936 79716 153010 79744
rect 152798 79648 152832 79688
rect 152148 79636 152154 79648
rect 152826 79636 152832 79648
rect 152884 79636 152890 79688
rect 152182 79608 152188 79620
rect 151694 79580 152188 79608
rect 152182 79568 152188 79580
rect 152240 79568 152246 79620
rect 151044 79512 151492 79540
rect 152936 79540 152964 79716
rect 153010 79568 153016 79620
rect 153068 79608 153074 79620
rect 153166 79608 153194 79784
rect 153068 79580 153194 79608
rect 153258 79620 153286 79840
rect 153258 79580 153292 79620
rect 153068 79568 153074 79580
rect 153286 79568 153292 79580
rect 153344 79568 153350 79620
rect 153102 79540 153108 79552
rect 152936 79512 153108 79540
rect 151044 79500 151050 79512
rect 153102 79500 153108 79512
rect 153160 79500 153166 79552
rect 153194 79500 153200 79552
rect 153252 79540 153258 79552
rect 153396 79540 153424 79840
rect 153626 79688 153654 79908
rect 154270 79824 154298 79908
rect 153884 79812 153890 79824
rect 153562 79636 153568 79688
rect 153620 79648 153654 79688
rect 153810 79784 153890 79812
rect 153620 79636 153626 79648
rect 153810 79620 153838 79784
rect 153884 79772 153890 79784
rect 153942 79772 153948 79824
rect 154068 79772 154074 79824
rect 154126 79772 154132 79824
rect 154206 79772 154212 79824
rect 154264 79784 154298 79824
rect 154264 79772 154270 79784
rect 154086 79688 154114 79772
rect 154086 79648 154120 79688
rect 154114 79636 154120 79648
rect 154172 79636 154178 79688
rect 154362 79676 154390 79908
rect 154454 79824 154482 79908
rect 154436 79772 154442 79824
rect 154494 79772 154500 79824
rect 154960 79756 154988 79908
rect 154942 79704 154948 79756
rect 155000 79704 155006 79756
rect 155144 79688 155172 79908
rect 155264 79840 155270 79892
rect 155322 79840 155328 79892
rect 155632 79840 155638 79892
rect 155690 79840 155696 79892
rect 155282 79756 155310 79840
rect 155282 79716 155316 79756
rect 155310 79704 155316 79716
rect 155368 79704 155374 79756
rect 154362 79648 154712 79676
rect 153810 79580 153844 79620
rect 153838 79568 153844 79580
rect 153896 79568 153902 79620
rect 154684 79608 154712 79648
rect 155126 79636 155132 79688
rect 155184 79636 155190 79688
rect 155650 79608 155678 79840
rect 155834 79756 155862 79908
rect 155908 79840 155914 79892
rect 155966 79840 155972 79892
rect 156000 79840 156006 79892
rect 156058 79840 156064 79892
rect 155770 79704 155776 79756
rect 155828 79716 155862 79756
rect 155828 79704 155834 79716
rect 155926 79688 155954 79840
rect 156018 79744 156046 79840
rect 156202 79824 156230 79908
rect 156202 79784 156236 79824
rect 156230 79772 156236 79784
rect 156288 79772 156294 79824
rect 156138 79744 156144 79756
rect 156018 79716 156144 79744
rect 156138 79704 156144 79716
rect 156196 79704 156202 79756
rect 155862 79636 155868 79688
rect 155920 79648 155954 79688
rect 155920 79636 155926 79648
rect 155954 79608 155960 79620
rect 154454 79580 154574 79608
rect 154684 79580 154896 79608
rect 155650 79580 155960 79608
rect 153252 79512 153424 79540
rect 153252 79500 153258 79512
rect 153470 79500 153476 79552
rect 153528 79540 153534 79552
rect 154454 79540 154482 79580
rect 153528 79512 154482 79540
rect 154546 79540 154574 79580
rect 154868 79540 154896 79580
rect 155954 79568 155960 79580
rect 156012 79568 156018 79620
rect 154546 79512 154712 79540
rect 154868 79512 155172 79540
rect 153528 79500 153534 79512
rect 154684 79484 154712 79512
rect 143810 79472 143816 79484
rect 143690 79444 143816 79472
rect 143810 79432 143816 79444
rect 143868 79432 143874 79484
rect 150250 79432 150256 79484
rect 150308 79444 150342 79484
rect 150308 79432 150314 79444
rect 150526 79432 150532 79484
rect 150584 79432 150590 79484
rect 154666 79432 154672 79484
rect 154724 79432 154730 79484
rect 138216 79376 144914 79404
rect 104158 79296 104164 79348
rect 104216 79336 104222 79348
rect 104710 79336 104716 79348
rect 104216 79308 104716 79336
rect 104216 79296 104222 79308
rect 104710 79296 104716 79308
rect 104768 79296 104774 79348
rect 110230 79296 110236 79348
rect 110288 79336 110294 79348
rect 141602 79336 141608 79348
rect 110288 79308 141608 79336
rect 110288 79296 110294 79308
rect 141602 79296 141608 79308
rect 141660 79296 141666 79348
rect 144886 79336 144914 79376
rect 149422 79364 149428 79416
rect 149480 79404 149486 79416
rect 149480 79376 154528 79404
rect 149480 79364 149486 79376
rect 144886 79308 153194 79336
rect 118050 79228 118056 79280
rect 118108 79268 118114 79280
rect 149238 79268 149244 79280
rect 118108 79240 149244 79268
rect 118108 79228 118114 79240
rect 149238 79228 149244 79240
rect 149296 79228 149302 79280
rect 104526 79160 104532 79212
rect 104584 79200 104590 79212
rect 104710 79200 104716 79212
rect 104584 79172 104716 79200
rect 104584 79160 104590 79172
rect 104710 79160 104716 79172
rect 104768 79160 104774 79212
rect 113082 79160 113088 79212
rect 113140 79200 113146 79212
rect 145558 79200 145564 79212
rect 113140 79172 145564 79200
rect 113140 79160 113146 79172
rect 145558 79160 145564 79172
rect 145616 79160 145622 79212
rect 113910 79092 113916 79144
rect 113968 79132 113974 79144
rect 146386 79132 146392 79144
rect 113968 79104 146392 79132
rect 113968 79092 113974 79104
rect 146386 79092 146392 79104
rect 146444 79092 146450 79144
rect 102870 79024 102876 79076
rect 102928 79064 102934 79076
rect 135346 79064 135352 79076
rect 102928 79036 135352 79064
rect 102928 79024 102934 79036
rect 135346 79024 135352 79036
rect 135404 79024 135410 79076
rect 136450 79024 136456 79076
rect 136508 79064 136514 79076
rect 136726 79064 136732 79076
rect 136508 79036 136732 79064
rect 136508 79024 136514 79036
rect 136726 79024 136732 79036
rect 136784 79064 136790 79076
rect 149422 79064 149428 79076
rect 136784 79036 149428 79064
rect 136784 79024 136790 79036
rect 149422 79024 149428 79036
rect 149480 79024 149486 79076
rect 112346 78956 112352 79008
rect 112404 78996 112410 79008
rect 145926 78996 145932 79008
rect 112404 78968 145932 78996
rect 112404 78956 112410 78968
rect 145926 78956 145932 78968
rect 145984 78956 145990 79008
rect 153166 78996 153194 79308
rect 154500 79200 154528 79376
rect 154666 79228 154672 79280
rect 154724 79268 154730 79280
rect 155144 79268 155172 79512
rect 156414 79500 156420 79552
rect 156472 79540 156478 79552
rect 156662 79540 156690 79908
rect 156736 79840 156742 79892
rect 156794 79840 156800 79892
rect 156828 79840 156834 79892
rect 156886 79840 156892 79892
rect 156472 79512 156690 79540
rect 156754 79552 156782 79840
rect 156846 79620 156874 79840
rect 156938 79688 156966 79908
rect 157030 79824 157058 79908
rect 157012 79772 157018 79824
rect 157070 79772 157076 79824
rect 157122 79744 157150 79908
rect 157076 79716 157150 79744
rect 157076 79688 157104 79716
rect 157214 79688 157242 79908
rect 157352 79756 157380 79908
rect 157490 79880 157518 79908
rect 157444 79852 157518 79880
rect 157334 79704 157340 79756
rect 157392 79704 157398 79756
rect 156938 79648 156972 79688
rect 156966 79636 156972 79648
rect 157024 79636 157030 79688
rect 157058 79636 157064 79688
rect 157116 79636 157122 79688
rect 157150 79636 157156 79688
rect 157208 79648 157242 79688
rect 157208 79636 157214 79648
rect 156846 79580 156880 79620
rect 156874 79568 156880 79580
rect 156932 79568 156938 79620
rect 157444 79608 157472 79852
rect 157564 79840 157570 79892
rect 157622 79840 157628 79892
rect 157674 79880 157702 79908
rect 157674 79852 157748 79880
rect 157582 79756 157610 79840
rect 157720 79824 157748 79852
rect 157702 79772 157708 79824
rect 157760 79772 157766 79824
rect 157518 79704 157524 79756
rect 157576 79716 157610 79756
rect 157576 79704 157582 79716
rect 157610 79636 157616 79688
rect 157668 79676 157674 79688
rect 157812 79676 157840 79988
rect 158318 79960 158346 79988
rect 158208 79908 158214 79960
rect 158266 79908 158272 79960
rect 158300 79908 158306 79960
rect 158358 79908 158364 79960
rect 157668 79648 157840 79676
rect 157668 79636 157674 79648
rect 157886 79608 157892 79620
rect 157444 79580 157892 79608
rect 157886 79568 157892 79580
rect 157944 79568 157950 79620
rect 158226 79552 158254 79908
rect 158502 79892 158530 80056
rect 162090 79960 162118 80600
rect 166092 79988 167086 80016
rect 166092 79960 166120 79988
rect 159128 79948 159134 79960
rect 159054 79920 159134 79948
rect 158484 79840 158490 79892
rect 158542 79840 158548 79892
rect 158576 79840 158582 79892
rect 158634 79840 158640 79892
rect 158944 79840 158950 79892
rect 159002 79840 159008 79892
rect 158594 79756 158622 79840
rect 158530 79704 158536 79756
rect 158588 79716 158622 79756
rect 158588 79704 158594 79716
rect 156754 79512 156788 79552
rect 156472 79500 156478 79512
rect 156782 79500 156788 79512
rect 156840 79500 156846 79552
rect 158226 79512 158260 79552
rect 158254 79500 158260 79512
rect 158312 79500 158318 79552
rect 158962 79540 158990 79840
rect 158824 79512 158990 79540
rect 158824 79336 158852 79512
rect 158898 79364 158904 79416
rect 158956 79404 158962 79416
rect 159054 79404 159082 79920
rect 159128 79908 159134 79920
rect 159186 79908 159192 79960
rect 159220 79908 159226 79960
rect 159278 79908 159284 79960
rect 159312 79908 159318 79960
rect 159370 79948 159376 79960
rect 159370 79908 159404 79948
rect 159496 79908 159502 79960
rect 159554 79948 159560 79960
rect 159864 79948 159870 79960
rect 159554 79908 159588 79948
rect 159238 79688 159266 79908
rect 159238 79648 159272 79688
rect 159266 79636 159272 79648
rect 159324 79636 159330 79688
rect 159174 79568 159180 79620
rect 159232 79608 159238 79620
rect 159376 79608 159404 79908
rect 159560 79756 159588 79908
rect 159836 79908 159870 79948
rect 159922 79908 159928 79960
rect 160232 79948 160238 79960
rect 160204 79908 160238 79948
rect 160290 79908 160296 79960
rect 160416 79908 160422 79960
rect 160474 79908 160480 79960
rect 160692 79908 160698 79960
rect 160750 79908 160756 79960
rect 160968 79948 160974 79960
rect 160940 79908 160974 79948
rect 161026 79908 161032 79960
rect 161612 79908 161618 79960
rect 161670 79908 161676 79960
rect 161704 79908 161710 79960
rect 161762 79948 161768 79960
rect 161762 79908 161796 79948
rect 161888 79908 161894 79960
rect 161946 79948 161952 79960
rect 161946 79908 161980 79948
rect 162072 79908 162078 79960
rect 162130 79908 162136 79960
rect 162164 79908 162170 79960
rect 162222 79908 162228 79960
rect 162256 79908 162262 79960
rect 162314 79948 162320 79960
rect 162992 79948 162998 79960
rect 162314 79920 162762 79948
rect 162314 79908 162320 79920
rect 159542 79704 159548 79756
rect 159600 79704 159606 79756
rect 159836 79620 159864 79908
rect 159956 79840 159962 79892
rect 160014 79840 160020 79892
rect 160048 79840 160054 79892
rect 160106 79880 160112 79892
rect 160106 79840 160140 79880
rect 159974 79812 160002 79840
rect 159974 79784 160048 79812
rect 160020 79756 160048 79784
rect 160002 79704 160008 79756
rect 160060 79704 160066 79756
rect 160112 79688 160140 79840
rect 160094 79636 160100 79688
rect 160152 79636 160158 79688
rect 159232 79580 159404 79608
rect 159232 79568 159238 79580
rect 159818 79568 159824 79620
rect 159876 79568 159882 79620
rect 160204 79472 160232 79908
rect 160434 79812 160462 79908
rect 160508 79840 160514 79892
rect 160566 79840 160572 79892
rect 160296 79784 160462 79812
rect 160296 79688 160324 79784
rect 160526 79756 160554 79840
rect 160710 79824 160738 79908
rect 160646 79772 160652 79824
rect 160704 79784 160738 79824
rect 160704 79772 160710 79784
rect 160526 79716 160560 79756
rect 160554 79704 160560 79716
rect 160612 79704 160618 79756
rect 160940 79688 160968 79908
rect 161152 79840 161158 79892
rect 161210 79880 161216 79892
rect 161630 79880 161658 79908
rect 161210 79852 161382 79880
rect 161630 79852 161704 79880
rect 161210 79840 161216 79852
rect 161244 79772 161250 79824
rect 161302 79772 161308 79824
rect 161262 79688 161290 79772
rect 160278 79636 160284 79688
rect 160336 79636 160342 79688
rect 160922 79636 160928 79688
rect 160980 79636 160986 79688
rect 161198 79636 161204 79688
rect 161256 79648 161290 79688
rect 161354 79676 161382 79852
rect 161520 79772 161526 79824
rect 161578 79772 161584 79824
rect 161538 79744 161566 79772
rect 161538 79716 161612 79744
rect 161474 79676 161480 79688
rect 161354 79648 161480 79676
rect 161256 79636 161262 79648
rect 161474 79636 161480 79648
rect 161532 79636 161538 79688
rect 160738 79500 160744 79552
rect 160796 79540 160802 79552
rect 161106 79540 161112 79552
rect 160796 79512 161112 79540
rect 160796 79500 160802 79512
rect 161106 79500 161112 79512
rect 161164 79500 161170 79552
rect 161584 79540 161612 79716
rect 161676 79620 161704 79852
rect 161768 79756 161796 79908
rect 161952 79824 161980 79908
rect 161934 79772 161940 79824
rect 161992 79772 161998 79824
rect 162182 79812 162210 79908
rect 162624 79840 162630 79892
rect 162682 79840 162688 79892
rect 162182 79784 162256 79812
rect 162228 79756 162256 79784
rect 161750 79704 161756 79756
rect 161808 79704 161814 79756
rect 162210 79704 162216 79756
rect 162268 79704 162274 79756
rect 162026 79636 162032 79688
rect 162084 79676 162090 79688
rect 162642 79676 162670 79840
rect 162084 79648 162670 79676
rect 162084 79636 162090 79648
rect 162734 79620 162762 79920
rect 162964 79908 162998 79948
rect 163050 79908 163056 79960
rect 163452 79908 163458 79960
rect 163510 79908 163516 79960
rect 164096 79908 164102 79960
rect 164154 79908 164160 79960
rect 164556 79908 164562 79960
rect 164614 79948 164620 79960
rect 164832 79948 164838 79960
rect 164614 79908 164648 79948
rect 162808 79772 162814 79824
rect 162866 79772 162872 79824
rect 162826 79688 162854 79772
rect 162964 79688 162992 79908
rect 163176 79840 163182 79892
rect 163234 79880 163240 79892
rect 163234 79840 163268 79880
rect 162826 79648 162860 79688
rect 162854 79636 162860 79648
rect 162912 79636 162918 79688
rect 162946 79636 162952 79688
rect 163004 79636 163010 79688
rect 163240 79620 163268 79840
rect 161658 79568 161664 79620
rect 161716 79568 161722 79620
rect 162670 79568 162676 79620
rect 162728 79580 162762 79620
rect 162728 79568 162734 79580
rect 163222 79568 163228 79620
rect 163280 79568 163286 79620
rect 161934 79540 161940 79552
rect 161584 79512 161940 79540
rect 161934 79500 161940 79512
rect 161992 79500 161998 79552
rect 160370 79472 160376 79484
rect 160204 79444 160376 79472
rect 160370 79432 160376 79444
rect 160428 79432 160434 79484
rect 163470 79472 163498 79908
rect 163544 79840 163550 79892
rect 163602 79840 163608 79892
rect 163562 79540 163590 79840
rect 163820 79812 163826 79824
rect 163792 79772 163826 79812
rect 163878 79772 163884 79824
rect 163912 79772 163918 79824
rect 163970 79772 163976 79824
rect 163792 79608 163820 79772
rect 163930 79688 163958 79772
rect 163866 79636 163872 79688
rect 163924 79648 163958 79688
rect 163924 79636 163930 79648
rect 164114 79620 164142 79908
rect 164464 79880 164470 79892
rect 164252 79852 164470 79880
rect 163958 79608 163964 79620
rect 163792 79580 163964 79608
rect 163958 79568 163964 79580
rect 164016 79568 164022 79620
rect 164114 79580 164148 79620
rect 164142 79568 164148 79580
rect 164200 79568 164206 79620
rect 163682 79540 163688 79552
rect 163562 79512 163688 79540
rect 163682 79500 163688 79512
rect 163740 79500 163746 79552
rect 164252 79540 164280 79852
rect 164464 79840 164470 79852
rect 164522 79840 164528 79892
rect 164620 79756 164648 79908
rect 164804 79908 164838 79948
rect 164890 79908 164896 79960
rect 165108 79908 165114 79960
rect 165166 79908 165172 79960
rect 165200 79908 165206 79960
rect 165258 79908 165264 79960
rect 165292 79908 165298 79960
rect 165350 79908 165356 79960
rect 165384 79908 165390 79960
rect 165442 79948 165448 79960
rect 165442 79908 165476 79948
rect 165936 79908 165942 79960
rect 165994 79948 166000 79960
rect 165994 79908 166028 79948
rect 166092 79920 166126 79960
rect 166120 79908 166126 79920
rect 166178 79908 166184 79960
rect 166396 79908 166402 79960
rect 166454 79908 166460 79960
rect 166672 79908 166678 79960
rect 166730 79908 166736 79960
rect 166764 79908 166770 79960
rect 166822 79948 166828 79960
rect 166822 79908 166856 79948
rect 166948 79908 166954 79960
rect 167006 79908 167012 79960
rect 164602 79704 164608 79756
rect 164660 79704 164666 79756
rect 164804 79688 164832 79908
rect 165126 79688 165154 79908
rect 165218 79756 165246 79908
rect 165310 79880 165338 79908
rect 165310 79852 165384 79880
rect 165356 79756 165384 79852
rect 165218 79716 165252 79756
rect 165246 79704 165252 79716
rect 165304 79704 165310 79756
rect 165338 79704 165344 79756
rect 165396 79704 165402 79756
rect 164786 79636 164792 79688
rect 164844 79636 164850 79688
rect 165126 79648 165160 79688
rect 165154 79636 165160 79648
rect 165212 79636 165218 79688
rect 165448 79620 165476 79908
rect 165752 79840 165758 79892
rect 165810 79840 165816 79892
rect 165844 79840 165850 79892
rect 165902 79840 165908 79892
rect 165770 79688 165798 79840
rect 165862 79756 165890 79840
rect 165862 79716 165896 79756
rect 165890 79704 165896 79716
rect 165948 79704 165954 79756
rect 166000 79688 166028 79908
rect 166304 79840 166310 79892
rect 166362 79840 166368 79892
rect 166322 79756 166350 79840
rect 166258 79704 166264 79756
rect 166316 79716 166350 79756
rect 166316 79704 166322 79716
rect 165770 79648 165804 79688
rect 165798 79636 165804 79648
rect 165856 79636 165862 79688
rect 165982 79636 165988 79688
rect 166040 79636 166046 79688
rect 166414 79676 166442 79908
rect 166690 79880 166718 79908
rect 166690 79852 166764 79880
rect 166488 79772 166494 79824
rect 166546 79812 166552 79824
rect 166546 79784 166672 79812
rect 166546 79772 166552 79784
rect 166534 79676 166540 79688
rect 166414 79648 166540 79676
rect 166534 79636 166540 79648
rect 166592 79636 166598 79688
rect 165430 79568 165436 79620
rect 165488 79568 165494 79620
rect 166442 79568 166448 79620
rect 166500 79608 166506 79620
rect 166644 79608 166672 79784
rect 166736 79620 166764 79852
rect 166828 79620 166856 79908
rect 166500 79580 166672 79608
rect 166500 79568 166506 79580
rect 166718 79568 166724 79620
rect 166776 79568 166782 79620
rect 166810 79568 166816 79620
rect 166868 79568 166874 79620
rect 164878 79540 164884 79552
rect 164252 79512 164884 79540
rect 164878 79500 164884 79512
rect 164936 79500 164942 79552
rect 166350 79500 166356 79552
rect 166408 79540 166414 79552
rect 166966 79540 166994 79908
rect 166408 79512 166994 79540
rect 166408 79500 166414 79512
rect 164050 79472 164056 79484
rect 163470 79444 164056 79472
rect 164050 79432 164056 79444
rect 164108 79432 164114 79484
rect 167058 79472 167086 79988
rect 167500 79948 167506 79960
rect 167150 79920 167506 79948
rect 167150 79540 167178 79920
rect 167500 79908 167506 79920
rect 167558 79908 167564 79960
rect 167592 79908 167598 79960
rect 167650 79948 167656 79960
rect 168300 79948 168328 80600
rect 172486 80560 172514 80600
rect 178586 80588 178592 80640
rect 178644 80628 178650 80640
rect 183526 80628 183554 80736
rect 211430 80724 211436 80736
rect 211488 80724 211494 80776
rect 207658 80696 207664 80708
rect 178644 80600 183554 80628
rect 186286 80668 207664 80696
rect 178644 80588 178650 80600
rect 178034 80560 178040 80572
rect 172486 80532 178040 80560
rect 178034 80520 178040 80532
rect 178092 80520 178098 80572
rect 186286 80560 186314 80668
rect 207658 80656 207664 80668
rect 207716 80656 207722 80708
rect 187694 80588 187700 80640
rect 187752 80628 187758 80640
rect 189074 80628 189080 80640
rect 187752 80600 189080 80628
rect 187752 80588 187758 80600
rect 189074 80588 189080 80600
rect 189132 80588 189138 80640
rect 183526 80532 186314 80560
rect 183526 80492 183554 80532
rect 188338 80520 188344 80572
rect 188396 80560 188402 80572
rect 194042 80560 194048 80572
rect 188396 80532 194048 80560
rect 188396 80520 188402 80532
rect 194042 80520 194048 80532
rect 194100 80520 194106 80572
rect 172486 80464 183554 80492
rect 172486 80424 172514 80464
rect 184198 80452 184204 80504
rect 184256 80492 184262 80504
rect 191374 80492 191380 80504
rect 184256 80464 191380 80492
rect 184256 80452 184262 80464
rect 191374 80452 191380 80464
rect 191432 80452 191438 80504
rect 177850 80424 177856 80436
rect 171106 80396 172514 80424
rect 174142 80396 177856 80424
rect 171106 80356 171134 80396
rect 169726 80328 171134 80356
rect 169726 80220 169754 80328
rect 167650 79920 168328 79948
rect 168576 80192 169754 80220
rect 167650 79908 167656 79920
rect 167224 79840 167230 79892
rect 167282 79880 167288 79892
rect 168576 79880 168604 80192
rect 174142 80016 174170 80396
rect 177850 80384 177856 80396
rect 177908 80384 177914 80436
rect 177758 80356 177764 80368
rect 173498 79988 174170 80016
rect 174234 80328 177764 80356
rect 173498 79960 173526 79988
rect 174234 79960 174262 80328
rect 177758 80316 177764 80328
rect 177816 80316 177822 80368
rect 178310 80288 178316 80300
rect 174878 80260 178316 80288
rect 174878 79960 174906 80260
rect 178310 80248 178316 80260
rect 178368 80248 178374 80300
rect 178402 80220 178408 80232
rect 176810 80192 178408 80220
rect 176810 80084 176838 80192
rect 178402 80180 178408 80192
rect 178460 80180 178466 80232
rect 178034 80152 178040 80164
rect 175614 80056 176838 80084
rect 176902 80124 178040 80152
rect 175614 79960 175642 80056
rect 176350 79988 176746 80016
rect 176350 79960 176378 79988
rect 169156 79908 169162 79960
rect 169214 79908 169220 79960
rect 170720 79908 170726 79960
rect 170778 79948 170784 79960
rect 172192 79948 172198 79960
rect 170778 79920 171180 79948
rect 170778 79908 170784 79920
rect 167282 79852 168604 79880
rect 167282 79840 167288 79852
rect 168788 79840 168794 79892
rect 168846 79840 168852 79892
rect 168972 79840 168978 79892
rect 169030 79840 169036 79892
rect 168420 79772 168426 79824
rect 168478 79772 168484 79824
rect 168512 79772 168518 79824
rect 168570 79772 168576 79824
rect 167822 79540 167828 79552
rect 167150 79512 167828 79540
rect 167822 79500 167828 79512
rect 167880 79500 167886 79552
rect 168438 79540 168466 79772
rect 168530 79676 168558 79772
rect 168650 79676 168656 79688
rect 168530 79648 168656 79676
rect 168650 79636 168656 79648
rect 168708 79636 168714 79688
rect 168806 79552 168834 79840
rect 168990 79688 169018 79840
rect 168990 79648 169024 79688
rect 169018 79636 169024 79648
rect 169076 79636 169082 79688
rect 168558 79540 168564 79552
rect 168438 79512 168564 79540
rect 168558 79500 168564 79512
rect 168616 79500 168622 79552
rect 168742 79500 168748 79552
rect 168800 79512 168834 79552
rect 168800 79500 168806 79512
rect 168466 79472 168472 79484
rect 167058 79444 168472 79472
rect 168466 79432 168472 79444
rect 168524 79432 168530 79484
rect 169174 79472 169202 79908
rect 169616 79880 169622 79892
rect 169312 79852 169622 79880
rect 169312 79540 169340 79852
rect 169616 79840 169622 79852
rect 169674 79840 169680 79892
rect 169984 79880 169990 79892
rect 169956 79840 169990 79880
rect 170042 79840 170048 79892
rect 170076 79840 170082 79892
rect 170134 79840 170140 79892
rect 169432 79772 169438 79824
rect 169490 79772 169496 79824
rect 169450 79676 169478 79772
rect 169956 79756 169984 79840
rect 170094 79756 170122 79840
rect 169938 79704 169944 79756
rect 169996 79704 170002 79756
rect 170030 79704 170036 79756
rect 170088 79716 170122 79756
rect 170088 79704 170094 79716
rect 169450 79648 169754 79676
rect 169478 79540 169484 79552
rect 169312 79512 169484 79540
rect 169478 79500 169484 79512
rect 169536 79500 169542 79552
rect 169726 79540 169754 79648
rect 170950 79540 170956 79552
rect 169726 79512 170956 79540
rect 170950 79500 170956 79512
rect 171008 79500 171014 79552
rect 171152 79540 171180 79920
rect 172072 79920 172198 79948
rect 171364 79840 171370 79892
rect 171422 79840 171428 79892
rect 171732 79880 171738 79892
rect 171704 79840 171738 79880
rect 171790 79840 171796 79892
rect 171824 79840 171830 79892
rect 171882 79840 171888 79892
rect 171382 79608 171410 79840
rect 171548 79772 171554 79824
rect 171606 79772 171612 79824
rect 171566 79688 171594 79772
rect 171704 79688 171732 79840
rect 171842 79688 171870 79840
rect 171502 79636 171508 79688
rect 171560 79648 171594 79688
rect 171560 79636 171566 79648
rect 171686 79636 171692 79688
rect 171744 79636 171750 79688
rect 171778 79636 171784 79688
rect 171836 79648 171870 79688
rect 171836 79636 171842 79648
rect 171382 79580 172008 79608
rect 171870 79540 171876 79552
rect 171152 79512 171876 79540
rect 171870 79500 171876 79512
rect 171928 79500 171934 79552
rect 170398 79472 170404 79484
rect 169174 79444 170404 79472
rect 170398 79432 170404 79444
rect 170456 79432 170462 79484
rect 171980 79472 172008 79580
rect 172072 79540 172100 79920
rect 172192 79908 172198 79920
rect 172250 79908 172256 79960
rect 172560 79908 172566 79960
rect 172618 79948 172624 79960
rect 172618 79920 172698 79948
rect 172618 79908 172624 79920
rect 172284 79840 172290 79892
rect 172342 79840 172348 79892
rect 172376 79840 172382 79892
rect 172434 79840 172440 79892
rect 172302 79608 172330 79840
rect 172394 79812 172422 79840
rect 172560 79812 172566 79824
rect 172394 79784 172566 79812
rect 172560 79772 172566 79784
rect 172618 79772 172624 79824
rect 172670 79620 172698 79920
rect 172836 79908 172842 79960
rect 172894 79908 172900 79960
rect 172928 79908 172934 79960
rect 172986 79948 172992 79960
rect 172986 79920 173158 79948
rect 172986 79908 172992 79920
rect 172744 79840 172750 79892
rect 172802 79840 172808 79892
rect 172762 79688 172790 79840
rect 172854 79744 172882 79908
rect 172854 79716 173020 79744
rect 172762 79648 172796 79688
rect 172790 79636 172796 79648
rect 172848 79636 172854 79688
rect 172992 79620 173020 79716
rect 172302 79580 172560 79608
rect 172670 79580 172704 79620
rect 172532 79552 172560 79580
rect 172698 79568 172704 79580
rect 172756 79568 172762 79620
rect 172974 79568 172980 79620
rect 173032 79568 173038 79620
rect 173130 79608 173158 79920
rect 173480 79908 173486 79960
rect 173538 79908 173544 79960
rect 173572 79908 173578 79960
rect 173630 79908 173636 79960
rect 173664 79908 173670 79960
rect 173722 79908 173728 79960
rect 173848 79908 173854 79960
rect 173906 79908 173912 79960
rect 174032 79908 174038 79960
rect 174090 79908 174096 79960
rect 174216 79908 174222 79960
rect 174274 79908 174280 79960
rect 174308 79908 174314 79960
rect 174366 79908 174372 79960
rect 174584 79908 174590 79960
rect 174642 79948 174648 79960
rect 174768 79948 174774 79960
rect 174642 79908 174676 79948
rect 173296 79840 173302 79892
rect 173354 79840 173360 79892
rect 173388 79840 173394 79892
rect 173446 79840 173452 79892
rect 173314 79688 173342 79840
rect 173406 79812 173434 79840
rect 173406 79784 173480 79812
rect 173452 79688 173480 79784
rect 173314 79648 173348 79688
rect 173342 79636 173348 79648
rect 173400 79636 173406 79688
rect 173434 79636 173440 79688
rect 173492 79636 173498 79688
rect 173590 79620 173618 79908
rect 173682 79756 173710 79908
rect 173866 79756 173894 79908
rect 174050 79824 174078 79908
rect 174326 79824 174354 79908
rect 174648 79824 174676 79908
rect 174740 79908 174774 79948
rect 174826 79908 174832 79960
rect 174860 79908 174866 79960
rect 174918 79908 174924 79960
rect 175136 79908 175142 79960
rect 175194 79908 175200 79960
rect 175596 79908 175602 79960
rect 175654 79908 175660 79960
rect 175780 79908 175786 79960
rect 175838 79908 175844 79960
rect 176056 79948 176062 79960
rect 176028 79908 176062 79948
rect 176114 79908 176120 79960
rect 176332 79908 176338 79960
rect 176390 79908 176396 79960
rect 176516 79908 176522 79960
rect 176574 79908 176580 79960
rect 174740 79824 174768 79908
rect 175044 79840 175050 79892
rect 175102 79840 175108 79892
rect 174032 79772 174038 79824
rect 174090 79772 174096 79824
rect 174262 79772 174268 79824
rect 174320 79784 174354 79824
rect 174320 79772 174326 79784
rect 174630 79772 174636 79824
rect 174688 79772 174694 79824
rect 174722 79772 174728 79824
rect 174780 79772 174786 79824
rect 173682 79716 173716 79756
rect 173710 79704 173716 79716
rect 173768 79704 173774 79756
rect 173866 79716 173900 79756
rect 173894 79704 173900 79716
rect 173952 79704 173958 79756
rect 175062 79676 175090 79840
rect 175154 79744 175182 79908
rect 175688 79880 175694 79892
rect 175660 79840 175694 79880
rect 175746 79840 175752 79892
rect 175660 79756 175688 79840
rect 175154 79716 175320 79744
rect 175182 79676 175188 79688
rect 175062 79648 175188 79676
rect 175182 79636 175188 79648
rect 175240 79636 175246 79688
rect 173250 79608 173256 79620
rect 173130 79580 173256 79608
rect 173250 79568 173256 79580
rect 173308 79568 173314 79620
rect 173590 79580 173624 79620
rect 173618 79568 173624 79580
rect 173676 79568 173682 79620
rect 175090 79568 175096 79620
rect 175148 79608 175154 79620
rect 175292 79608 175320 79716
rect 175642 79704 175648 79756
rect 175700 79704 175706 79756
rect 175148 79580 175320 79608
rect 175798 79620 175826 79908
rect 176028 79824 176056 79908
rect 176148 79840 176154 79892
rect 176206 79840 176212 79892
rect 176534 79880 176562 79908
rect 176534 79852 176608 79880
rect 176010 79772 176016 79824
rect 176068 79772 176074 79824
rect 176166 79756 176194 79840
rect 176424 79772 176430 79824
rect 176482 79772 176488 79824
rect 176102 79704 176108 79756
rect 176160 79716 176194 79756
rect 176160 79704 176166 79716
rect 176286 79636 176292 79688
rect 176344 79676 176350 79688
rect 176442 79676 176470 79772
rect 176344 79648 176470 79676
rect 176344 79636 176350 79648
rect 176580 79620 176608 79852
rect 176718 79744 176746 79988
rect 176792 79840 176798 79892
rect 176850 79880 176856 79892
rect 176902 79880 176930 80124
rect 178034 80112 178040 80124
rect 178092 80112 178098 80164
rect 178126 80112 178132 80164
rect 178184 80152 178190 80164
rect 181162 80152 181168 80164
rect 178184 80124 181168 80152
rect 178184 80112 178190 80124
rect 181162 80112 181168 80124
rect 181220 80112 181226 80164
rect 177758 80044 177764 80096
rect 177816 80084 177822 80096
rect 179598 80084 179604 80096
rect 177816 80056 179604 80084
rect 177816 80044 177822 80056
rect 179598 80044 179604 80056
rect 179656 80044 179662 80096
rect 191374 80044 191380 80096
rect 191432 80084 191438 80096
rect 198182 80084 198188 80096
rect 191432 80056 198188 80084
rect 191432 80044 191438 80056
rect 198182 80044 198188 80056
rect 198240 80044 198246 80096
rect 177942 79976 177948 80028
rect 178000 80016 178006 80028
rect 178126 80016 178132 80028
rect 178000 79988 178132 80016
rect 178000 79976 178006 79988
rect 178126 79976 178132 79988
rect 178184 79976 178190 80028
rect 184934 79976 184940 80028
rect 184992 80016 184998 80028
rect 215662 80016 215668 80028
rect 184992 79988 215668 80016
rect 184992 79976 184998 79988
rect 215662 79976 215668 79988
rect 215720 79976 215726 80028
rect 176976 79908 176982 79960
rect 177034 79908 177040 79960
rect 177160 79908 177166 79960
rect 177218 79908 177224 79960
rect 177270 79920 179414 79948
rect 176850 79852 176930 79880
rect 176850 79840 176856 79852
rect 176994 79824 177022 79908
rect 176930 79772 176936 79824
rect 176988 79784 177022 79824
rect 177178 79812 177206 79908
rect 177270 79892 177298 79920
rect 177252 79840 177258 79892
rect 177310 79840 177316 79892
rect 177344 79840 177350 79892
rect 177402 79880 177408 79892
rect 178494 79880 178500 79892
rect 177402 79852 178500 79880
rect 177402 79840 177408 79852
rect 178494 79840 178500 79852
rect 178552 79840 178558 79892
rect 179386 79880 179414 79920
rect 182910 79880 182916 79892
rect 179386 79852 182916 79880
rect 182910 79840 182916 79852
rect 182968 79840 182974 79892
rect 194042 79840 194048 79892
rect 194100 79880 194106 79892
rect 200850 79880 200856 79892
rect 194100 79852 200856 79880
rect 194100 79840 194106 79852
rect 200850 79840 200856 79852
rect 200908 79840 200914 79892
rect 177666 79812 177672 79824
rect 177178 79784 177672 79812
rect 176988 79772 176994 79784
rect 177666 79772 177672 79784
rect 177724 79772 177730 79824
rect 177298 79744 177304 79756
rect 176718 79716 177304 79744
rect 177298 79704 177304 79716
rect 177356 79704 177362 79756
rect 189074 79636 189080 79688
rect 189132 79676 189138 79688
rect 203058 79676 203064 79688
rect 189132 79648 203064 79676
rect 189132 79636 189138 79648
rect 203058 79636 203064 79648
rect 203116 79636 203122 79688
rect 175798 79580 175832 79620
rect 175148 79568 175154 79580
rect 175826 79568 175832 79580
rect 175884 79568 175890 79620
rect 176562 79568 176568 79620
rect 176620 79568 176626 79620
rect 181438 79568 181444 79620
rect 181496 79608 181502 79620
rect 580810 79608 580816 79620
rect 181496 79580 580816 79608
rect 181496 79568 181502 79580
rect 580810 79568 580816 79580
rect 580868 79568 580874 79620
rect 172072 79512 172376 79540
rect 172348 79484 172376 79512
rect 172514 79500 172520 79552
rect 172572 79500 172578 79552
rect 173158 79500 173164 79552
rect 173216 79540 173222 79552
rect 188982 79540 188988 79552
rect 173216 79512 188988 79540
rect 173216 79500 173222 79512
rect 188982 79500 188988 79512
rect 189040 79500 189046 79552
rect 172054 79472 172060 79484
rect 171980 79444 172060 79472
rect 172054 79432 172060 79444
rect 172112 79432 172118 79484
rect 172330 79432 172336 79484
rect 172388 79432 172394 79484
rect 173894 79432 173900 79484
rect 173952 79472 173958 79484
rect 214650 79472 214656 79484
rect 173952 79444 214656 79472
rect 173952 79432 173958 79444
rect 214650 79432 214656 79444
rect 214708 79432 214714 79484
rect 158956 79376 159082 79404
rect 158956 79364 158962 79376
rect 159358 79364 159364 79416
rect 159416 79404 159422 79416
rect 167178 79404 167184 79416
rect 159416 79376 167184 79404
rect 159416 79364 159422 79376
rect 167178 79364 167184 79376
rect 167236 79364 167242 79416
rect 167270 79364 167276 79416
rect 167328 79404 167334 79416
rect 187694 79404 187700 79416
rect 167328 79376 187700 79404
rect 167328 79364 167334 79376
rect 187694 79364 187700 79376
rect 187752 79364 187758 79416
rect 160462 79336 160468 79348
rect 158824 79308 160468 79336
rect 160462 79296 160468 79308
rect 160520 79296 160526 79348
rect 160554 79296 160560 79348
rect 160612 79336 160618 79348
rect 195238 79336 195244 79348
rect 160612 79308 195244 79336
rect 160612 79296 160618 79308
rect 195238 79296 195244 79308
rect 195296 79296 195302 79348
rect 154724 79240 155172 79268
rect 154724 79228 154730 79240
rect 167178 79228 167184 79280
rect 167236 79268 167242 79280
rect 167236 79240 168972 79268
rect 167236 79228 167242 79240
rect 159358 79200 159364 79212
rect 154500 79172 159364 79200
rect 159358 79160 159364 79172
rect 159416 79160 159422 79212
rect 168944 79200 168972 79240
rect 171962 79228 171968 79280
rect 172020 79268 172026 79280
rect 210602 79268 210608 79280
rect 172020 79240 210608 79268
rect 172020 79228 172026 79240
rect 210602 79228 210608 79240
rect 210660 79228 210666 79280
rect 181438 79200 181444 79212
rect 161768 79172 166994 79200
rect 168944 79172 181444 79200
rect 154574 79092 154580 79144
rect 154632 79132 154638 79144
rect 155586 79132 155592 79144
rect 154632 79104 155592 79132
rect 154632 79092 154638 79104
rect 155586 79092 155592 79104
rect 155644 79092 155650 79144
rect 161768 78996 161796 79172
rect 166966 79132 166994 79172
rect 181438 79160 181444 79172
rect 181496 79160 181502 79212
rect 181530 79160 181536 79212
rect 181588 79200 181594 79212
rect 215478 79200 215484 79212
rect 181588 79172 215484 79200
rect 181588 79160 181594 79172
rect 215478 79160 215484 79172
rect 215536 79160 215542 79212
rect 175642 79132 175648 79144
rect 166966 79104 175648 79132
rect 175642 79092 175648 79104
rect 175700 79092 175706 79144
rect 179598 79092 179604 79144
rect 179656 79132 179662 79144
rect 215754 79132 215760 79144
rect 179656 79104 215760 79132
rect 179656 79092 179662 79104
rect 215754 79092 215760 79104
rect 215812 79092 215818 79144
rect 170490 79024 170496 79076
rect 170548 79064 170554 79076
rect 212810 79064 212816 79076
rect 170548 79036 212816 79064
rect 170548 79024 170554 79036
rect 212810 79024 212816 79036
rect 212868 79024 212874 79076
rect 153166 78968 161796 78996
rect 174262 78956 174268 79008
rect 174320 78996 174326 79008
rect 219618 78996 219624 79008
rect 174320 78968 219624 78996
rect 174320 78956 174326 78968
rect 219618 78956 219624 78968
rect 219676 78956 219682 79008
rect 129182 78888 129188 78940
rect 129240 78928 129246 78940
rect 138750 78928 138756 78940
rect 129240 78900 138756 78928
rect 129240 78888 129246 78900
rect 138750 78888 138756 78900
rect 138808 78888 138814 78940
rect 160922 78888 160928 78940
rect 160980 78928 160986 78940
rect 210510 78928 210516 78940
rect 160980 78900 210516 78928
rect 160980 78888 160986 78900
rect 210510 78888 210516 78900
rect 210568 78888 210574 78940
rect 95970 78820 95976 78872
rect 96028 78860 96034 78872
rect 152274 78860 152280 78872
rect 96028 78832 152280 78860
rect 96028 78820 96034 78832
rect 152274 78820 152280 78832
rect 152332 78820 152338 78872
rect 161750 78820 161756 78872
rect 161808 78860 161814 78872
rect 217134 78860 217140 78872
rect 161808 78832 217140 78860
rect 161808 78820 161814 78832
rect 217134 78820 217140 78832
rect 217192 78820 217198 78872
rect 131022 78752 131028 78804
rect 131080 78792 131086 78804
rect 141510 78792 141516 78804
rect 131080 78764 141516 78792
rect 131080 78752 131086 78764
rect 141510 78752 141516 78764
rect 141568 78752 141574 78804
rect 157426 78752 157432 78804
rect 157484 78792 157490 78804
rect 158162 78792 158168 78804
rect 157484 78764 158168 78792
rect 157484 78752 157490 78764
rect 158162 78752 158168 78764
rect 158220 78752 158226 78804
rect 175734 78752 175740 78804
rect 175792 78792 175798 78804
rect 180242 78792 180248 78804
rect 175792 78764 180248 78792
rect 175792 78752 175798 78764
rect 180242 78752 180248 78764
rect 180300 78752 180306 78804
rect 181162 78752 181168 78804
rect 181220 78792 181226 78804
rect 212718 78792 212724 78804
rect 181220 78764 212724 78792
rect 181220 78752 181226 78764
rect 212718 78752 212724 78764
rect 212776 78752 212782 78804
rect 135346 78684 135352 78736
rect 135404 78724 135410 78736
rect 135806 78724 135812 78736
rect 135404 78696 135812 78724
rect 135404 78684 135410 78696
rect 135806 78684 135812 78696
rect 135864 78684 135870 78736
rect 136726 78684 136732 78736
rect 136784 78724 136790 78736
rect 137002 78724 137008 78736
rect 136784 78696 137008 78724
rect 136784 78684 136790 78696
rect 137002 78684 137008 78696
rect 137060 78684 137066 78736
rect 141234 78684 141240 78736
rect 141292 78724 141298 78736
rect 141878 78724 141884 78736
rect 141292 78696 141884 78724
rect 141292 78684 141298 78696
rect 141878 78684 141884 78696
rect 141936 78684 141942 78736
rect 142706 78684 142712 78736
rect 142764 78724 142770 78736
rect 142982 78724 142988 78736
rect 142764 78696 142988 78724
rect 142764 78684 142770 78696
rect 142982 78684 142988 78696
rect 143040 78684 143046 78736
rect 153286 78684 153292 78736
rect 153344 78724 153350 78736
rect 154390 78724 154396 78736
rect 153344 78696 154396 78724
rect 153344 78684 153350 78696
rect 154390 78684 154396 78696
rect 154448 78684 154454 78736
rect 171226 78684 171232 78736
rect 171284 78724 171290 78736
rect 171502 78724 171508 78736
rect 171284 78696 171508 78724
rect 171284 78684 171290 78696
rect 171502 78684 171508 78696
rect 171560 78684 171566 78736
rect 172238 78684 172244 78736
rect 172296 78724 172302 78736
rect 180610 78724 180616 78736
rect 172296 78696 180616 78724
rect 172296 78684 172302 78696
rect 180610 78684 180616 78696
rect 180668 78684 180674 78736
rect 96522 78616 96528 78668
rect 96580 78656 96586 78668
rect 132034 78656 132040 78668
rect 96580 78628 132040 78656
rect 96580 78616 96586 78628
rect 132034 78616 132040 78628
rect 132092 78616 132098 78668
rect 132126 78616 132132 78668
rect 132184 78656 132190 78668
rect 143350 78656 143356 78668
rect 132184 78628 143356 78656
rect 132184 78616 132190 78628
rect 143350 78616 143356 78628
rect 143408 78616 143414 78668
rect 145282 78616 145288 78668
rect 145340 78656 145346 78668
rect 145466 78656 145472 78668
rect 145340 78628 145472 78656
rect 145340 78616 145346 78628
rect 145466 78616 145472 78628
rect 145524 78616 145530 78668
rect 154022 78616 154028 78668
rect 154080 78656 154086 78668
rect 154482 78656 154488 78668
rect 154080 78628 154488 78656
rect 154080 78616 154086 78628
rect 154482 78616 154488 78628
rect 154540 78616 154546 78668
rect 159542 78616 159548 78668
rect 159600 78656 159606 78668
rect 159600 78628 166994 78656
rect 159600 78616 159606 78628
rect 121822 78548 121828 78600
rect 121880 78588 121886 78600
rect 136450 78588 136456 78600
rect 121880 78560 136456 78588
rect 121880 78548 121886 78560
rect 136450 78548 136456 78560
rect 136508 78548 136514 78600
rect 166966 78588 166994 78628
rect 170582 78616 170588 78668
rect 170640 78656 170646 78668
rect 173894 78656 173900 78668
rect 170640 78628 173900 78656
rect 170640 78616 170646 78628
rect 173894 78616 173900 78628
rect 173952 78616 173958 78668
rect 177574 78616 177580 78668
rect 177632 78656 177638 78668
rect 219894 78656 219900 78668
rect 177632 78628 219900 78656
rect 177632 78616 177638 78628
rect 219894 78616 219900 78628
rect 219952 78616 219958 78668
rect 169478 78588 169484 78600
rect 166966 78560 169484 78588
rect 169478 78548 169484 78560
rect 169536 78548 169542 78600
rect 170398 78548 170404 78600
rect 170456 78588 170462 78600
rect 171502 78588 171508 78600
rect 170456 78560 171508 78588
rect 170456 78548 170462 78560
rect 171502 78548 171508 78560
rect 171560 78548 171566 78600
rect 172514 78548 172520 78600
rect 172572 78588 172578 78600
rect 173618 78588 173624 78600
rect 172572 78560 173624 78588
rect 172572 78548 172578 78560
rect 173618 78548 173624 78560
rect 173676 78548 173682 78600
rect 178034 78548 178040 78600
rect 178092 78588 178098 78600
rect 189534 78588 189540 78600
rect 178092 78560 189540 78588
rect 178092 78548 178098 78560
rect 189534 78548 189540 78560
rect 189592 78548 189598 78600
rect 105906 78480 105912 78532
rect 105964 78520 105970 78532
rect 139946 78520 139952 78532
rect 105964 78492 139952 78520
rect 105964 78480 105970 78492
rect 139946 78480 139952 78492
rect 140004 78480 140010 78532
rect 142982 78480 142988 78532
rect 143040 78520 143046 78532
rect 151906 78520 151912 78532
rect 143040 78492 151912 78520
rect 143040 78480 143046 78492
rect 151906 78480 151912 78492
rect 151964 78480 151970 78532
rect 165430 78480 165436 78532
rect 165488 78520 165494 78532
rect 165488 78492 167500 78520
rect 165488 78480 165494 78492
rect 103974 78412 103980 78464
rect 104032 78452 104038 78464
rect 136634 78452 136640 78464
rect 104032 78424 136640 78452
rect 104032 78412 104038 78424
rect 136634 78412 136640 78424
rect 136692 78412 136698 78464
rect 165614 78412 165620 78464
rect 165672 78452 165678 78464
rect 166166 78452 166172 78464
rect 165672 78424 166172 78452
rect 165672 78412 165678 78424
rect 166166 78412 166172 78424
rect 166224 78412 166230 78464
rect 167472 78452 167500 78492
rect 167546 78480 167552 78532
rect 167604 78520 167610 78532
rect 169570 78520 169576 78532
rect 167604 78492 169576 78520
rect 167604 78480 167610 78492
rect 169570 78480 169576 78492
rect 169628 78480 169634 78532
rect 170582 78480 170588 78532
rect 170640 78520 170646 78532
rect 171042 78520 171048 78532
rect 170640 78492 171048 78520
rect 170640 78480 170646 78492
rect 171042 78480 171048 78492
rect 171100 78480 171106 78532
rect 214098 78520 214104 78532
rect 171152 78492 214104 78520
rect 171152 78452 171180 78492
rect 214098 78480 214104 78492
rect 214156 78480 214162 78532
rect 167472 78424 171180 78452
rect 171318 78412 171324 78464
rect 171376 78452 171382 78464
rect 206278 78452 206284 78464
rect 171376 78424 206284 78452
rect 171376 78412 171382 78424
rect 206278 78412 206284 78424
rect 206336 78412 206342 78464
rect 99742 78344 99748 78396
rect 99800 78384 99806 78396
rect 131574 78384 131580 78396
rect 99800 78356 131580 78384
rect 99800 78344 99806 78356
rect 131574 78344 131580 78356
rect 131632 78344 131638 78396
rect 139394 78384 139400 78396
rect 133156 78356 139400 78384
rect 130378 78276 130384 78328
rect 130436 78316 130442 78328
rect 132126 78316 132132 78328
rect 130436 78288 132132 78316
rect 130436 78276 130442 78288
rect 132126 78276 132132 78288
rect 132184 78276 132190 78328
rect 108298 78208 108304 78260
rect 108356 78248 108362 78260
rect 133156 78248 133184 78356
rect 139394 78344 139400 78356
rect 139452 78344 139458 78396
rect 169018 78344 169024 78396
rect 169076 78384 169082 78396
rect 169076 78356 176654 78384
rect 169076 78344 169082 78356
rect 136634 78276 136640 78328
rect 136692 78316 136698 78328
rect 142062 78316 142068 78328
rect 136692 78288 142068 78316
rect 136692 78276 136698 78288
rect 142062 78276 142068 78288
rect 142120 78276 142126 78328
rect 146294 78276 146300 78328
rect 146352 78316 146358 78328
rect 155126 78316 155132 78328
rect 146352 78288 155132 78316
rect 146352 78276 146358 78288
rect 155126 78276 155132 78288
rect 155184 78276 155190 78328
rect 176626 78316 176654 78356
rect 177206 78344 177212 78396
rect 177264 78384 177270 78396
rect 211706 78384 211712 78396
rect 177264 78356 211712 78384
rect 177264 78344 177270 78356
rect 211706 78344 211712 78356
rect 211764 78344 211770 78396
rect 203610 78316 203616 78328
rect 176626 78288 203616 78316
rect 203610 78276 203616 78288
rect 203668 78276 203674 78328
rect 108356 78220 133184 78248
rect 108356 78208 108362 78220
rect 138842 78208 138848 78260
rect 138900 78248 138906 78260
rect 146110 78248 146116 78260
rect 138900 78220 146116 78248
rect 138900 78208 138906 78220
rect 146110 78208 146116 78220
rect 146168 78208 146174 78260
rect 152366 78208 152372 78260
rect 152424 78248 152430 78260
rect 152918 78248 152924 78260
rect 152424 78220 152924 78248
rect 152424 78208 152430 78220
rect 152918 78208 152924 78220
rect 152976 78208 152982 78260
rect 164418 78208 164424 78260
rect 164476 78248 164482 78260
rect 165246 78248 165252 78260
rect 164476 78220 165252 78248
rect 164476 78208 164482 78220
rect 165246 78208 165252 78220
rect 165304 78208 165310 78260
rect 175458 78208 175464 78260
rect 175516 78248 175522 78260
rect 189718 78248 189724 78260
rect 175516 78220 189724 78248
rect 175516 78208 175522 78220
rect 189718 78208 189724 78220
rect 189776 78208 189782 78260
rect 102778 78140 102784 78192
rect 102836 78180 102842 78192
rect 129918 78180 129924 78192
rect 102836 78152 129924 78180
rect 102836 78140 102842 78152
rect 129918 78140 129924 78152
rect 129976 78140 129982 78192
rect 132862 78140 132868 78192
rect 132920 78180 132926 78192
rect 138382 78180 138388 78192
rect 132920 78152 138388 78180
rect 132920 78140 132926 78152
rect 138382 78140 138388 78152
rect 138440 78140 138446 78192
rect 140038 78140 140044 78192
rect 140096 78180 140102 78192
rect 150710 78180 150716 78192
rect 140096 78152 150716 78180
rect 140096 78140 140102 78152
rect 150710 78140 150716 78152
rect 150768 78140 150774 78192
rect 157886 78140 157892 78192
rect 157944 78180 157950 78192
rect 157944 78152 160140 78180
rect 157944 78140 157950 78152
rect 101766 78072 101772 78124
rect 101824 78112 101830 78124
rect 131022 78112 131028 78124
rect 101824 78084 131028 78112
rect 101824 78072 101830 78084
rect 131022 78072 131028 78084
rect 131080 78072 131086 78124
rect 132034 78072 132040 78124
rect 132092 78112 132098 78124
rect 134518 78112 134524 78124
rect 132092 78084 134524 78112
rect 132092 78072 132098 78084
rect 134518 78072 134524 78084
rect 134576 78072 134582 78124
rect 135898 78072 135904 78124
rect 135956 78112 135962 78124
rect 143258 78112 143264 78124
rect 135956 78084 143264 78112
rect 135956 78072 135962 78084
rect 143258 78072 143264 78084
rect 143316 78072 143322 78124
rect 145926 78072 145932 78124
rect 145984 78112 145990 78124
rect 158530 78112 158536 78124
rect 145984 78084 158536 78112
rect 145984 78072 145990 78084
rect 158530 78072 158536 78084
rect 158588 78072 158594 78124
rect 103882 78004 103888 78056
rect 103940 78044 103946 78056
rect 137462 78044 137468 78056
rect 103940 78016 137468 78044
rect 103940 78004 103946 78016
rect 137462 78004 137468 78016
rect 137520 78004 137526 78056
rect 140406 78004 140412 78056
rect 140464 78044 140470 78056
rect 151722 78044 151728 78056
rect 140464 78016 151728 78044
rect 140464 78004 140470 78016
rect 151722 78004 151728 78016
rect 151780 78004 151786 78056
rect 160112 78044 160140 78152
rect 181714 78140 181720 78192
rect 181772 78180 181778 78192
rect 196526 78180 196532 78192
rect 181772 78152 196532 78180
rect 181772 78140 181778 78152
rect 196526 78140 196532 78152
rect 196584 78140 196590 78192
rect 173710 78072 173716 78124
rect 173768 78112 173774 78124
rect 179690 78112 179696 78124
rect 173768 78084 179696 78112
rect 173768 78072 173774 78084
rect 179690 78072 179696 78084
rect 179748 78072 179754 78124
rect 181530 78072 181536 78124
rect 181588 78112 181594 78124
rect 196434 78112 196440 78124
rect 181588 78084 196440 78112
rect 181588 78072 181594 78084
rect 196434 78072 196440 78084
rect 196492 78072 196498 78124
rect 167546 78044 167552 78056
rect 160112 78016 167552 78044
rect 167546 78004 167552 78016
rect 167604 78004 167610 78056
rect 168926 78004 168932 78056
rect 168984 78044 168990 78056
rect 168984 78016 171410 78044
rect 168984 78004 168990 78016
rect 120810 77936 120816 77988
rect 120868 77976 120874 77988
rect 134058 77976 134064 77988
rect 120868 77948 134064 77976
rect 120868 77936 120874 77948
rect 134058 77936 134064 77948
rect 134116 77936 134122 77988
rect 146018 77976 146024 77988
rect 137986 77948 146024 77976
rect 105722 77868 105728 77920
rect 105780 77908 105786 77920
rect 128170 77908 128176 77920
rect 105780 77880 128176 77908
rect 105780 77868 105786 77880
rect 128170 77868 128176 77880
rect 128228 77868 128234 77920
rect 135622 77908 135628 77920
rect 128326 77880 135628 77908
rect 101582 77800 101588 77852
rect 101640 77840 101646 77852
rect 128326 77840 128354 77880
rect 135622 77868 135628 77880
rect 135680 77868 135686 77920
rect 137002 77868 137008 77920
rect 137060 77908 137066 77920
rect 137986 77908 138014 77948
rect 146018 77936 146024 77948
rect 146076 77936 146082 77988
rect 157518 77936 157524 77988
rect 157576 77976 157582 77988
rect 169662 77976 169668 77988
rect 157576 77948 169668 77976
rect 157576 77936 157582 77948
rect 169662 77936 169668 77948
rect 169720 77936 169726 77988
rect 171382 77976 171410 78016
rect 172790 78004 172796 78056
rect 172848 78044 172854 78056
rect 181254 78044 181260 78056
rect 172848 78016 181260 78044
rect 172848 78004 172854 78016
rect 181254 78004 181260 78016
rect 181312 78004 181318 78056
rect 181806 78004 181812 78056
rect 181864 78044 181870 78056
rect 197906 78044 197912 78056
rect 181864 78016 197912 78044
rect 181864 78004 181870 78016
rect 197906 78004 197912 78016
rect 197964 78004 197970 78056
rect 177850 77976 177856 77988
rect 171382 77948 177856 77976
rect 177850 77936 177856 77948
rect 177908 77936 177914 77988
rect 180334 77936 180340 77988
rect 180392 77976 180398 77988
rect 202230 77976 202236 77988
rect 180392 77948 202236 77976
rect 180392 77936 180398 77948
rect 202230 77936 202236 77948
rect 202288 77936 202294 77988
rect 137060 77880 138014 77908
rect 137060 77868 137066 77880
rect 157978 77868 157984 77920
rect 158036 77908 158042 77920
rect 166810 77908 166816 77920
rect 158036 77880 166816 77908
rect 158036 77868 158042 77880
rect 166810 77868 166816 77880
rect 166868 77868 166874 77920
rect 174170 77868 174176 77920
rect 174228 77908 174234 77920
rect 174446 77908 174452 77920
rect 174228 77880 174452 77908
rect 174228 77868 174234 77880
rect 174446 77868 174452 77880
rect 174504 77868 174510 77920
rect 181346 77868 181352 77920
rect 181404 77908 181410 77920
rect 193766 77908 193772 77920
rect 181404 77880 193772 77908
rect 181404 77868 181410 77880
rect 193766 77868 193772 77880
rect 193824 77868 193830 77920
rect 101640 77812 128354 77840
rect 101640 77800 101646 77812
rect 135714 77800 135720 77852
rect 135772 77840 135778 77852
rect 148870 77840 148876 77852
rect 135772 77812 148876 77840
rect 135772 77800 135778 77812
rect 148870 77800 148876 77812
rect 148928 77800 148934 77852
rect 171594 77800 171600 77852
rect 171652 77840 171658 77852
rect 181438 77840 181444 77852
rect 171652 77812 181444 77840
rect 171652 77800 171658 77812
rect 181438 77800 181444 77812
rect 181496 77800 181502 77852
rect 103054 77732 103060 77784
rect 103112 77772 103118 77784
rect 134978 77772 134984 77784
rect 103112 77744 134984 77772
rect 103112 77732 103118 77744
rect 134978 77732 134984 77744
rect 135036 77732 135042 77784
rect 166626 77732 166632 77784
rect 166684 77772 166690 77784
rect 171870 77772 171876 77784
rect 166684 77744 171876 77772
rect 166684 77732 166690 77744
rect 171870 77732 171876 77744
rect 171928 77732 171934 77784
rect 174630 77732 174636 77784
rect 174688 77772 174694 77784
rect 189994 77772 190000 77784
rect 174688 77744 190000 77772
rect 174688 77732 174694 77744
rect 189994 77732 190000 77744
rect 190052 77732 190058 77784
rect 136818 77664 136824 77716
rect 136876 77704 136882 77716
rect 144546 77704 144552 77716
rect 136876 77676 144552 77704
rect 136876 77664 136882 77676
rect 144546 77664 144552 77676
rect 144604 77664 144610 77716
rect 166718 77664 166724 77716
rect 166776 77704 166782 77716
rect 173894 77704 173900 77716
rect 166776 77676 173900 77704
rect 166776 77664 166782 77676
rect 173894 77664 173900 77676
rect 173952 77664 173958 77716
rect 142890 77596 142896 77648
rect 142948 77636 142954 77648
rect 154114 77636 154120 77648
rect 142948 77608 154120 77636
rect 142948 77596 142954 77608
rect 154114 77596 154120 77608
rect 154172 77596 154178 77648
rect 155494 77596 155500 77648
rect 155552 77636 155558 77648
rect 173158 77636 173164 77648
rect 155552 77608 173164 77636
rect 155552 77596 155558 77608
rect 173158 77596 173164 77608
rect 173216 77596 173222 77648
rect 173802 77596 173808 77648
rect 173860 77636 173866 77648
rect 210418 77636 210424 77648
rect 173860 77608 210424 77636
rect 173860 77596 173866 77608
rect 210418 77596 210424 77608
rect 210476 77596 210482 77648
rect 159082 77460 159088 77512
rect 159140 77500 159146 77512
rect 162578 77500 162584 77512
rect 159140 77472 162584 77500
rect 159140 77460 159146 77472
rect 162578 77460 162584 77472
rect 162636 77460 162642 77512
rect 169110 77460 169116 77512
rect 169168 77500 169174 77512
rect 170674 77500 170680 77512
rect 169168 77472 170680 77500
rect 169168 77460 169174 77472
rect 170674 77460 170680 77472
rect 170732 77460 170738 77512
rect 164602 77392 164608 77444
rect 164660 77432 164666 77444
rect 165522 77432 165528 77444
rect 164660 77404 165528 77432
rect 164660 77392 164666 77404
rect 165522 77392 165528 77404
rect 165580 77392 165586 77444
rect 168834 77324 168840 77376
rect 168892 77364 168898 77376
rect 174630 77364 174636 77376
rect 168892 77336 174636 77364
rect 168892 77324 168898 77336
rect 174630 77324 174636 77336
rect 174688 77324 174694 77376
rect 136082 77256 136088 77308
rect 136140 77296 136146 77308
rect 138934 77296 138940 77308
rect 136140 77268 138940 77296
rect 136140 77256 136146 77268
rect 138934 77256 138940 77268
rect 138992 77256 138998 77308
rect 97166 77188 97172 77240
rect 97224 77228 97230 77240
rect 97224 77200 103514 77228
rect 97224 77188 97230 77200
rect 103486 77160 103514 77200
rect 116394 77188 116400 77240
rect 116452 77228 116458 77240
rect 156690 77228 156696 77240
rect 116452 77200 156696 77228
rect 116452 77188 116458 77200
rect 156690 77188 156696 77200
rect 156748 77188 156754 77240
rect 163498 77188 163504 77240
rect 163556 77228 163562 77240
rect 164142 77228 164148 77240
rect 163556 77200 164148 77228
rect 163556 77188 163562 77200
rect 164142 77188 164148 77200
rect 164200 77188 164206 77240
rect 165890 77188 165896 77240
rect 165948 77228 165954 77240
rect 166166 77228 166172 77240
rect 165948 77200 166172 77228
rect 165948 77188 165954 77200
rect 166166 77188 166172 77200
rect 166224 77188 166230 77240
rect 177666 77188 177672 77240
rect 177724 77228 177730 77240
rect 201678 77228 201684 77240
rect 177724 77200 201684 77228
rect 177724 77188 177730 77200
rect 201678 77188 201684 77200
rect 201736 77188 201742 77240
rect 168466 77160 168472 77172
rect 103486 77132 168472 77160
rect 168466 77120 168472 77132
rect 168524 77120 168530 77172
rect 177298 77120 177304 77172
rect 177356 77160 177362 77172
rect 191190 77160 191196 77172
rect 177356 77132 191196 77160
rect 177356 77120 177362 77132
rect 191190 77120 191196 77132
rect 191248 77120 191254 77172
rect 107010 77052 107016 77104
rect 107068 77092 107074 77104
rect 139486 77092 139492 77104
rect 107068 77064 139492 77092
rect 107068 77052 107074 77064
rect 139486 77052 139492 77064
rect 139544 77052 139550 77104
rect 147950 77052 147956 77104
rect 148008 77092 148014 77104
rect 149974 77092 149980 77104
rect 148008 77064 149980 77092
rect 148008 77052 148014 77064
rect 149974 77052 149980 77064
rect 150032 77092 150038 77104
rect 200942 77092 200948 77104
rect 150032 77064 200948 77092
rect 150032 77052 150038 77064
rect 200942 77052 200948 77064
rect 201000 77052 201006 77104
rect 116946 76984 116952 77036
rect 117004 77024 117010 77036
rect 167270 77024 167276 77036
rect 117004 76996 167276 77024
rect 117004 76984 117010 76996
rect 167270 76984 167276 76996
rect 167328 76984 167334 77036
rect 173342 76984 173348 77036
rect 173400 77024 173406 77036
rect 209038 77024 209044 77036
rect 173400 76996 209044 77024
rect 173400 76984 173406 76996
rect 209038 76984 209044 76996
rect 209096 76984 209102 77036
rect 117866 76916 117872 76968
rect 117924 76956 117930 76968
rect 117924 76928 155770 76956
rect 117924 76916 117930 76928
rect 2866 76848 2872 76900
rect 2924 76888 2930 76900
rect 120074 76888 120080 76900
rect 2924 76860 120080 76888
rect 2924 76848 2930 76860
rect 120074 76848 120080 76860
rect 120132 76848 120138 76900
rect 121270 76848 121276 76900
rect 121328 76888 121334 76900
rect 153194 76888 153200 76900
rect 121328 76860 153200 76888
rect 121328 76848 121334 76860
rect 153166 76848 153200 76860
rect 153252 76848 153258 76900
rect 102962 76780 102968 76832
rect 103020 76820 103026 76832
rect 133230 76820 133236 76832
rect 103020 76792 133236 76820
rect 103020 76780 103026 76792
rect 133230 76780 133236 76792
rect 133288 76780 133294 76832
rect 134334 76780 134340 76832
rect 134392 76820 134398 76832
rect 134978 76820 134984 76832
rect 134392 76792 134984 76820
rect 134392 76780 134398 76792
rect 134978 76780 134984 76792
rect 135036 76780 135042 76832
rect 146662 76780 146668 76832
rect 146720 76820 146726 76832
rect 147030 76820 147036 76832
rect 146720 76792 147036 76820
rect 146720 76780 146726 76792
rect 147030 76780 147036 76792
rect 147088 76780 147094 76832
rect 117406 76712 117412 76764
rect 117464 76752 117470 76764
rect 148962 76752 148968 76764
rect 117464 76724 148968 76752
rect 117464 76712 117470 76724
rect 148962 76712 148968 76724
rect 149020 76712 149026 76764
rect 109494 76644 109500 76696
rect 109552 76684 109558 76696
rect 136818 76684 136824 76696
rect 109552 76656 136824 76684
rect 109552 76644 109558 76656
rect 136818 76644 136824 76656
rect 136876 76644 136882 76696
rect 148226 76644 148232 76696
rect 148284 76684 148290 76696
rect 148594 76684 148600 76696
rect 148284 76656 148600 76684
rect 148284 76644 148290 76656
rect 148594 76644 148600 76656
rect 148652 76644 148658 76696
rect 150710 76644 150716 76696
rect 150768 76684 150774 76696
rect 150894 76684 150900 76696
rect 150768 76656 150900 76684
rect 150768 76644 150774 76656
rect 150894 76644 150900 76656
rect 150952 76644 150958 76696
rect 119154 76576 119160 76628
rect 119212 76616 119218 76628
rect 144086 76616 144092 76628
rect 119212 76588 144092 76616
rect 119212 76576 119218 76588
rect 144086 76576 144092 76588
rect 144144 76576 144150 76628
rect 146754 76576 146760 76628
rect 146812 76616 146818 76628
rect 147030 76616 147036 76628
rect 146812 76588 147036 76616
rect 146812 76576 146818 76588
rect 147030 76576 147036 76588
rect 147088 76576 147094 76628
rect 153166 76616 153194 76848
rect 155742 76820 155770 76928
rect 156690 76916 156696 76968
rect 156748 76956 156754 76968
rect 159266 76956 159272 76968
rect 156748 76928 159272 76956
rect 156748 76916 156754 76928
rect 159266 76916 159272 76928
rect 159324 76956 159330 76968
rect 193950 76956 193956 76968
rect 159324 76928 193956 76956
rect 159324 76916 159330 76928
rect 193950 76916 193956 76928
rect 194008 76916 194014 76968
rect 160094 76848 160100 76900
rect 160152 76888 160158 76900
rect 164142 76888 164148 76900
rect 160152 76860 164148 76888
rect 160152 76848 160158 76860
rect 164142 76848 164148 76860
rect 164200 76848 164206 76900
rect 178494 76848 178500 76900
rect 178552 76888 178558 76900
rect 211890 76888 211896 76900
rect 178552 76860 211896 76888
rect 178552 76848 178558 76860
rect 211890 76848 211896 76860
rect 211948 76848 211954 76900
rect 156782 76820 156788 76832
rect 155742 76792 156788 76820
rect 156782 76780 156788 76792
rect 156840 76820 156846 76832
rect 190822 76820 190828 76832
rect 156840 76792 190828 76820
rect 156840 76780 156846 76792
rect 190822 76780 190828 76792
rect 190880 76780 190886 76832
rect 168466 76712 168472 76764
rect 168524 76752 168530 76764
rect 200298 76752 200304 76764
rect 168524 76724 200304 76752
rect 168524 76712 168530 76724
rect 200298 76712 200304 76724
rect 200356 76712 200362 76764
rect 154942 76644 154948 76696
rect 155000 76684 155006 76696
rect 155770 76684 155776 76696
rect 155000 76656 155776 76684
rect 155000 76644 155006 76656
rect 155770 76644 155776 76656
rect 155828 76644 155834 76696
rect 156782 76644 156788 76696
rect 156840 76684 156846 76696
rect 157150 76684 157156 76696
rect 156840 76656 157156 76684
rect 156840 76644 156846 76656
rect 157150 76644 157156 76656
rect 157208 76644 157214 76696
rect 157794 76644 157800 76696
rect 157852 76684 157858 76696
rect 158438 76684 158444 76696
rect 157852 76656 158444 76684
rect 157852 76644 157858 76656
rect 158438 76644 158444 76656
rect 158496 76644 158502 76696
rect 160094 76644 160100 76696
rect 160152 76684 160158 76696
rect 160370 76684 160376 76696
rect 160152 76656 160376 76684
rect 160152 76644 160158 76656
rect 160370 76644 160376 76656
rect 160428 76644 160434 76696
rect 165706 76644 165712 76696
rect 165764 76684 165770 76696
rect 199378 76684 199384 76696
rect 165764 76656 199384 76684
rect 165764 76644 165770 76656
rect 199378 76644 199384 76656
rect 199436 76644 199442 76696
rect 182910 76616 182916 76628
rect 153166 76588 182916 76616
rect 182910 76576 182916 76588
rect 182968 76576 182974 76628
rect 104526 76508 104532 76560
rect 104584 76548 104590 76560
rect 136266 76548 136272 76560
rect 104584 76520 136272 76548
rect 104584 76508 104590 76520
rect 136266 76508 136272 76520
rect 136324 76508 136330 76560
rect 136818 76508 136824 76560
rect 136876 76548 136882 76560
rect 137646 76548 137652 76560
rect 136876 76520 137652 76548
rect 136876 76508 136882 76520
rect 137646 76508 137652 76520
rect 137704 76508 137710 76560
rect 138290 76508 138296 76560
rect 138348 76548 138354 76560
rect 138474 76548 138480 76560
rect 138348 76520 138480 76548
rect 138348 76508 138354 76520
rect 138474 76508 138480 76520
rect 138532 76508 138538 76560
rect 140774 76508 140780 76560
rect 140832 76548 140838 76560
rect 141326 76548 141332 76560
rect 140832 76520 141332 76548
rect 140832 76508 140838 76520
rect 141326 76508 141332 76520
rect 141384 76508 141390 76560
rect 141510 76508 141516 76560
rect 141568 76548 141574 76560
rect 143074 76548 143080 76560
rect 141568 76520 143080 76548
rect 141568 76508 141574 76520
rect 143074 76508 143080 76520
rect 143132 76508 143138 76560
rect 148134 76508 148140 76560
rect 148192 76548 148198 76560
rect 148594 76548 148600 76560
rect 148192 76520 148600 76548
rect 148192 76508 148198 76520
rect 148594 76508 148600 76520
rect 148652 76508 148658 76560
rect 150894 76508 150900 76560
rect 150952 76548 150958 76560
rect 151630 76548 151636 76560
rect 150952 76520 151636 76548
rect 150952 76508 150958 76520
rect 151630 76508 151636 76520
rect 151688 76508 151694 76560
rect 155954 76508 155960 76560
rect 156012 76548 156018 76560
rect 196434 76548 196440 76560
rect 156012 76520 196440 76548
rect 156012 76508 156018 76520
rect 196434 76508 196440 76520
rect 196492 76508 196498 76560
rect 131850 76440 131856 76492
rect 131908 76480 131914 76492
rect 150802 76480 150808 76492
rect 131908 76452 150808 76480
rect 131908 76440 131914 76452
rect 150802 76440 150808 76452
rect 150860 76440 150866 76492
rect 155126 76440 155132 76492
rect 155184 76480 155190 76492
rect 155862 76480 155868 76492
rect 155184 76452 155868 76480
rect 155184 76440 155190 76452
rect 155862 76440 155868 76452
rect 155920 76440 155926 76492
rect 158530 76440 158536 76492
rect 158588 76480 158594 76492
rect 217226 76480 217232 76492
rect 158588 76452 217232 76480
rect 158588 76440 158594 76452
rect 217226 76440 217232 76452
rect 217284 76440 217290 76492
rect 120074 76372 120080 76424
rect 120132 76412 120138 76424
rect 120994 76412 121000 76424
rect 120132 76384 121000 76412
rect 120132 76372 120138 76384
rect 120994 76372 121000 76384
rect 121052 76412 121058 76424
rect 153930 76412 153936 76424
rect 121052 76384 153936 76412
rect 121052 76372 121058 76384
rect 153930 76372 153936 76384
rect 153988 76372 153994 76424
rect 171318 76372 171324 76424
rect 171376 76412 171382 76424
rect 171778 76412 171784 76424
rect 171376 76384 171784 76412
rect 171376 76372 171382 76384
rect 171778 76372 171784 76384
rect 171836 76372 171842 76424
rect 214558 76412 214564 76424
rect 179386 76384 214564 76412
rect 138014 76304 138020 76356
rect 138072 76344 138078 76356
rect 138474 76344 138480 76356
rect 138072 76316 138480 76344
rect 138072 76304 138078 76316
rect 138474 76304 138480 76316
rect 138532 76304 138538 76356
rect 146754 76304 146760 76356
rect 146812 76344 146818 76356
rect 147306 76344 147312 76356
rect 146812 76316 147312 76344
rect 146812 76304 146818 76316
rect 147306 76304 147312 76316
rect 147364 76304 147370 76356
rect 174998 76304 175004 76356
rect 175056 76344 175062 76356
rect 179386 76344 179414 76384
rect 214558 76372 214564 76384
rect 214616 76372 214622 76424
rect 175056 76316 179414 76344
rect 175056 76304 175062 76316
rect 140866 76168 140872 76220
rect 140924 76208 140930 76220
rect 141142 76208 141148 76220
rect 140924 76180 141148 76208
rect 140924 76168 140930 76180
rect 141142 76168 141148 76180
rect 141200 76168 141206 76220
rect 134058 76100 134064 76152
rect 134116 76140 134122 76152
rect 134518 76140 134524 76152
rect 134116 76112 134524 76140
rect 134116 76100 134122 76112
rect 134518 76100 134524 76112
rect 134576 76100 134582 76152
rect 156230 76100 156236 76152
rect 156288 76140 156294 76152
rect 156966 76140 156972 76152
rect 156288 76112 156972 76140
rect 156288 76100 156294 76112
rect 156966 76100 156972 76112
rect 157024 76100 157030 76152
rect 163682 76100 163688 76152
rect 163740 76140 163746 76152
rect 165062 76140 165068 76152
rect 163740 76112 165068 76140
rect 163740 76100 163746 76112
rect 165062 76100 165068 76112
rect 165120 76100 165126 76152
rect 137186 76032 137192 76084
rect 137244 76072 137250 76084
rect 138566 76072 138572 76084
rect 137244 76044 138572 76072
rect 137244 76032 137250 76044
rect 138566 76032 138572 76044
rect 138624 76032 138630 76084
rect 146846 75964 146852 76016
rect 146904 76004 146910 76016
rect 147214 76004 147220 76016
rect 146904 75976 147220 76004
rect 146904 75964 146910 75976
rect 147214 75964 147220 75976
rect 147272 75964 147278 76016
rect 126330 75896 126336 75948
rect 126388 75936 126394 75948
rect 132034 75936 132040 75948
rect 126388 75908 132040 75936
rect 126388 75896 126394 75908
rect 132034 75896 132040 75908
rect 132092 75896 132098 75948
rect 143534 75896 143540 75948
rect 143592 75936 143598 75948
rect 152366 75936 152372 75948
rect 143592 75908 152372 75936
rect 143592 75896 143598 75908
rect 152366 75896 152372 75908
rect 152424 75896 152430 75948
rect 155218 75896 155224 75948
rect 155276 75936 155282 75948
rect 158254 75936 158260 75948
rect 155276 75908 158260 75936
rect 155276 75896 155282 75908
rect 158254 75896 158260 75908
rect 158312 75896 158318 75948
rect 162670 75896 162676 75948
rect 162728 75936 162734 75948
rect 170858 75936 170864 75948
rect 162728 75908 170864 75936
rect 162728 75896 162734 75908
rect 170858 75896 170864 75908
rect 170916 75896 170922 75948
rect 172514 75896 172520 75948
rect 172572 75936 172578 75948
rect 172974 75936 172980 75948
rect 172572 75908 172980 75936
rect 172572 75896 172578 75908
rect 172974 75896 172980 75908
rect 173032 75896 173038 75948
rect 173986 75896 173992 75948
rect 174044 75936 174050 75948
rect 174814 75936 174820 75948
rect 174044 75908 174820 75936
rect 174044 75896 174050 75908
rect 174814 75896 174820 75908
rect 174872 75896 174878 75948
rect 99650 75828 99656 75880
rect 99708 75868 99714 75880
rect 102778 75868 102784 75880
rect 99708 75840 102784 75868
rect 99708 75828 99714 75840
rect 102778 75828 102784 75840
rect 102836 75828 102842 75880
rect 124490 75828 124496 75880
rect 124548 75868 124554 75880
rect 135714 75868 135720 75880
rect 124548 75840 135720 75868
rect 124548 75828 124554 75840
rect 135714 75828 135720 75840
rect 135772 75828 135778 75880
rect 138198 75828 138204 75880
rect 138256 75868 138262 75880
rect 145650 75868 145656 75880
rect 138256 75840 145656 75868
rect 138256 75828 138262 75840
rect 145650 75828 145656 75840
rect 145708 75828 145714 75880
rect 157334 75828 157340 75880
rect 157392 75868 157398 75880
rect 157610 75868 157616 75880
rect 157392 75840 157616 75868
rect 157392 75828 157398 75840
rect 157610 75828 157616 75840
rect 157668 75828 157674 75880
rect 174262 75828 174268 75880
rect 174320 75868 174326 75880
rect 175090 75868 175096 75880
rect 174320 75840 175096 75868
rect 174320 75828 174326 75840
rect 175090 75828 175096 75840
rect 175148 75828 175154 75880
rect 196434 75828 196440 75880
rect 196492 75868 196498 75880
rect 217318 75868 217324 75880
rect 196492 75840 217324 75868
rect 196492 75828 196498 75840
rect 217318 75828 217324 75840
rect 217376 75828 217382 75880
rect 97442 75760 97448 75812
rect 97500 75800 97506 75812
rect 97500 75772 103514 75800
rect 97500 75760 97506 75772
rect 103486 75732 103514 75772
rect 130838 75760 130844 75812
rect 130896 75800 130902 75812
rect 133322 75800 133328 75812
rect 130896 75772 133328 75800
rect 130896 75760 130902 75772
rect 133322 75760 133328 75772
rect 133380 75760 133386 75812
rect 137922 75760 137928 75812
rect 137980 75800 137986 75812
rect 153102 75800 153108 75812
rect 137980 75772 153108 75800
rect 137980 75760 137986 75772
rect 153102 75760 153108 75772
rect 153160 75760 153166 75812
rect 167086 75760 167092 75812
rect 167144 75800 167150 75812
rect 174354 75800 174360 75812
rect 167144 75772 174360 75800
rect 167144 75760 167150 75772
rect 174354 75760 174360 75772
rect 174412 75800 174418 75812
rect 192294 75800 192300 75812
rect 174412 75772 192300 75800
rect 174412 75760 174418 75772
rect 192294 75760 192300 75772
rect 192352 75760 192358 75812
rect 147582 75732 147588 75744
rect 103486 75704 147588 75732
rect 147582 75692 147588 75704
rect 147640 75692 147646 75744
rect 162118 75692 162124 75744
rect 162176 75732 162182 75744
rect 171042 75732 171048 75744
rect 162176 75704 171048 75732
rect 162176 75692 162182 75704
rect 171042 75692 171048 75704
rect 171100 75692 171106 75744
rect 175826 75692 175832 75744
rect 175884 75732 175890 75744
rect 214282 75732 214288 75744
rect 175884 75704 214288 75732
rect 175884 75692 175890 75704
rect 214282 75692 214288 75704
rect 214340 75692 214346 75744
rect 114370 75624 114376 75676
rect 114428 75664 114434 75676
rect 142062 75664 142068 75676
rect 114428 75636 142068 75664
rect 114428 75624 114434 75636
rect 142062 75624 142068 75636
rect 142120 75624 142126 75676
rect 156046 75624 156052 75676
rect 156104 75664 156110 75676
rect 156874 75664 156880 75676
rect 156104 75636 156880 75664
rect 156104 75624 156110 75636
rect 156874 75624 156880 75636
rect 156932 75624 156938 75676
rect 157334 75624 157340 75676
rect 157392 75664 157398 75676
rect 158070 75664 158076 75676
rect 157392 75636 158076 75664
rect 157392 75624 157398 75636
rect 158070 75624 158076 75636
rect 158128 75624 158134 75676
rect 160370 75624 160376 75676
rect 160428 75664 160434 75676
rect 161198 75664 161204 75676
rect 160428 75636 161204 75664
rect 160428 75624 160434 75636
rect 161198 75624 161204 75636
rect 161256 75624 161262 75676
rect 162670 75624 162676 75676
rect 162728 75664 162734 75676
rect 164970 75664 164976 75676
rect 162728 75636 164976 75664
rect 162728 75624 162734 75636
rect 164970 75624 164976 75636
rect 165028 75664 165034 75676
rect 199286 75664 199292 75676
rect 165028 75636 199292 75664
rect 165028 75624 165034 75636
rect 199286 75624 199292 75636
rect 199344 75624 199350 75676
rect 116762 75556 116768 75608
rect 116820 75596 116826 75608
rect 117130 75596 117136 75608
rect 116820 75568 117136 75596
rect 116820 75556 116826 75568
rect 117130 75556 117136 75568
rect 117188 75596 117194 75608
rect 149146 75596 149152 75608
rect 117188 75568 149152 75596
rect 117188 75556 117194 75568
rect 149146 75556 149152 75568
rect 149204 75556 149210 75608
rect 181254 75556 181260 75608
rect 181312 75596 181318 75608
rect 182082 75596 182088 75608
rect 181312 75568 182088 75596
rect 181312 75556 181318 75568
rect 182082 75556 182088 75568
rect 182140 75596 182146 75608
rect 214190 75596 214196 75608
rect 182140 75568 214196 75596
rect 182140 75556 182146 75568
rect 214190 75556 214196 75568
rect 214248 75556 214254 75608
rect 116302 75488 116308 75540
rect 116360 75528 116366 75540
rect 148502 75528 148508 75540
rect 116360 75500 148508 75528
rect 116360 75488 116366 75500
rect 148502 75488 148508 75500
rect 148560 75488 148566 75540
rect 175366 75488 175372 75540
rect 175424 75528 175430 75540
rect 175918 75528 175924 75540
rect 175424 75500 175924 75528
rect 175424 75488 175430 75500
rect 175918 75488 175924 75500
rect 175976 75488 175982 75540
rect 179690 75488 179696 75540
rect 179748 75528 179754 75540
rect 205082 75528 205088 75540
rect 179748 75500 205088 75528
rect 179748 75488 179754 75500
rect 205082 75488 205088 75500
rect 205140 75488 205146 75540
rect 118234 75420 118240 75472
rect 118292 75460 118298 75472
rect 140498 75460 140504 75472
rect 118292 75432 140504 75460
rect 118292 75420 118298 75432
rect 140498 75420 140504 75432
rect 140556 75420 140562 75472
rect 142338 75460 142344 75472
rect 140746 75432 142344 75460
rect 114462 75352 114468 75404
rect 114520 75392 114526 75404
rect 140746 75392 140774 75432
rect 142338 75420 142344 75432
rect 142396 75460 142402 75472
rect 143074 75460 143080 75472
rect 142396 75432 143080 75460
rect 142396 75420 142402 75432
rect 143074 75420 143080 75432
rect 143132 75420 143138 75472
rect 146570 75420 146576 75472
rect 146628 75460 146634 75472
rect 147398 75460 147404 75472
rect 146628 75432 147404 75460
rect 146628 75420 146634 75432
rect 147398 75420 147404 75432
rect 147456 75420 147462 75472
rect 148134 75420 148140 75472
rect 148192 75460 148198 75472
rect 148410 75460 148416 75472
rect 148192 75432 148416 75460
rect 148192 75420 148198 75432
rect 148410 75420 148416 75432
rect 148468 75420 148474 75472
rect 158806 75420 158812 75472
rect 158864 75460 158870 75472
rect 159082 75460 159088 75472
rect 158864 75432 159088 75460
rect 158864 75420 158870 75432
rect 159082 75420 159088 75432
rect 159140 75420 159146 75472
rect 175826 75420 175832 75472
rect 175884 75460 175890 75472
rect 176470 75460 176476 75472
rect 175884 75432 176476 75460
rect 175884 75420 175890 75432
rect 176470 75420 176476 75432
rect 176528 75460 176534 75472
rect 198826 75460 198832 75472
rect 176528 75432 198832 75460
rect 176528 75420 176534 75432
rect 198826 75420 198832 75432
rect 198884 75420 198890 75472
rect 114520 75364 140774 75392
rect 114520 75352 114526 75364
rect 141050 75352 141056 75404
rect 141108 75392 141114 75404
rect 142062 75392 142068 75404
rect 141108 75364 142068 75392
rect 141108 75352 141114 75364
rect 142062 75352 142068 75364
rect 142120 75352 142126 75404
rect 158714 75352 158720 75404
rect 158772 75392 158778 75404
rect 159266 75392 159272 75404
rect 158772 75364 159272 75392
rect 158772 75352 158778 75364
rect 159266 75352 159272 75364
rect 159324 75352 159330 75404
rect 165798 75352 165804 75404
rect 165856 75392 165862 75404
rect 166258 75392 166264 75404
rect 165856 75364 166264 75392
rect 165856 75352 165862 75364
rect 166258 75352 166264 75364
rect 166316 75352 166322 75404
rect 170214 75352 170220 75404
rect 170272 75392 170278 75404
rect 192570 75392 192576 75404
rect 170272 75364 192576 75392
rect 170272 75352 170278 75364
rect 192570 75352 192576 75364
rect 192628 75352 192634 75404
rect 119522 75284 119528 75336
rect 119580 75324 119586 75336
rect 138198 75324 138204 75336
rect 119580 75296 138204 75324
rect 119580 75284 119586 75296
rect 138198 75284 138204 75296
rect 138256 75284 138262 75336
rect 138658 75284 138664 75336
rect 138716 75324 138722 75336
rect 143902 75324 143908 75336
rect 138716 75296 143908 75324
rect 138716 75284 138722 75296
rect 143902 75284 143908 75296
rect 143960 75284 143966 75336
rect 158806 75284 158812 75336
rect 158864 75324 158870 75336
rect 159726 75324 159732 75336
rect 158864 75296 159732 75324
rect 158864 75284 158870 75296
rect 159726 75284 159732 75296
rect 159784 75284 159790 75336
rect 165706 75284 165712 75336
rect 165764 75324 165770 75336
rect 166534 75324 166540 75336
rect 165764 75296 166540 75324
rect 165764 75284 165770 75296
rect 166534 75284 166540 75296
rect 166592 75284 166598 75336
rect 166994 75284 167000 75336
rect 167052 75324 167058 75336
rect 168282 75324 168288 75336
rect 167052 75296 168288 75324
rect 167052 75284 167058 75296
rect 168282 75284 168288 75296
rect 168340 75284 168346 75336
rect 171686 75284 171692 75336
rect 171744 75324 171750 75336
rect 171962 75324 171968 75336
rect 171744 75296 171968 75324
rect 171744 75284 171750 75296
rect 171962 75284 171968 75296
rect 172020 75284 172026 75336
rect 174446 75284 174452 75336
rect 174504 75324 174510 75336
rect 192478 75324 192484 75336
rect 174504 75296 192484 75324
rect 174504 75284 174510 75296
rect 192478 75284 192484 75296
rect 192536 75284 192542 75336
rect 107654 75216 107660 75268
rect 107712 75256 107718 75268
rect 126330 75256 126336 75268
rect 107712 75228 126336 75256
rect 107712 75216 107718 75228
rect 126330 75216 126336 75228
rect 126388 75216 126394 75268
rect 133046 75216 133052 75268
rect 133104 75256 133110 75268
rect 133782 75256 133788 75268
rect 133104 75228 133788 75256
rect 133104 75216 133110 75228
rect 133782 75216 133788 75228
rect 133840 75216 133846 75268
rect 135530 75216 135536 75268
rect 135588 75256 135594 75268
rect 135990 75256 135996 75268
rect 135588 75228 135996 75256
rect 135588 75216 135594 75228
rect 135990 75216 135996 75228
rect 136048 75216 136054 75268
rect 138566 75216 138572 75268
rect 138624 75256 138630 75268
rect 139302 75256 139308 75268
rect 138624 75228 139308 75256
rect 138624 75216 138630 75228
rect 139302 75216 139308 75228
rect 139360 75216 139366 75268
rect 146846 75216 146852 75268
rect 146904 75256 146910 75268
rect 147490 75256 147496 75268
rect 146904 75228 147496 75256
rect 146904 75216 146910 75228
rect 147490 75216 147496 75228
rect 147548 75216 147554 75268
rect 150434 75216 150440 75268
rect 150492 75256 150498 75268
rect 151170 75256 151176 75268
rect 150492 75228 151176 75256
rect 150492 75216 150498 75228
rect 151170 75216 151176 75228
rect 151228 75216 151234 75268
rect 158714 75216 158720 75268
rect 158772 75256 158778 75268
rect 158990 75256 158996 75268
rect 158772 75228 158996 75256
rect 158772 75216 158778 75228
rect 158990 75216 158996 75228
rect 159048 75216 159054 75268
rect 161566 75216 161572 75268
rect 161624 75256 161630 75268
rect 162210 75256 162216 75268
rect 161624 75228 162216 75256
rect 161624 75216 161630 75228
rect 162210 75216 162216 75228
rect 162268 75216 162274 75268
rect 165890 75216 165896 75268
rect 165948 75256 165954 75268
rect 166442 75256 166448 75268
rect 165948 75228 166448 75256
rect 165948 75216 165954 75228
rect 166442 75216 166448 75228
rect 166500 75216 166506 75268
rect 167178 75216 167184 75268
rect 167236 75256 167242 75268
rect 167730 75256 167736 75268
rect 167236 75228 167736 75256
rect 167236 75216 167242 75228
rect 167730 75216 167736 75228
rect 167788 75216 167794 75268
rect 168466 75216 168472 75268
rect 168524 75256 168530 75268
rect 169202 75256 169208 75268
rect 168524 75228 169208 75256
rect 168524 75216 168530 75228
rect 169202 75216 169208 75228
rect 169260 75216 169266 75268
rect 175274 75216 175280 75268
rect 175332 75256 175338 75268
rect 176194 75256 176200 75268
rect 175332 75228 176200 75256
rect 175332 75216 175338 75228
rect 176194 75216 176200 75228
rect 176252 75216 176258 75268
rect 40034 75148 40040 75200
rect 40092 75188 40098 75200
rect 117130 75188 117136 75200
rect 40092 75160 117136 75188
rect 40092 75148 40098 75160
rect 117130 75148 117136 75160
rect 117188 75148 117194 75200
rect 120074 75148 120080 75200
rect 120132 75188 120138 75200
rect 167086 75188 167092 75200
rect 120132 75160 167092 75188
rect 120132 75148 120138 75160
rect 167086 75148 167092 75160
rect 167144 75148 167150 75200
rect 167270 75148 167276 75200
rect 167328 75188 167334 75200
rect 168098 75188 168104 75200
rect 167328 75160 168104 75188
rect 167328 75148 167334 75160
rect 168098 75148 168104 75160
rect 168156 75148 168162 75200
rect 168190 75148 168196 75200
rect 168248 75188 168254 75200
rect 177942 75188 177948 75200
rect 168248 75160 177948 75188
rect 168248 75148 168254 75160
rect 177942 75148 177948 75160
rect 178000 75148 178006 75200
rect 194502 75148 194508 75200
rect 194560 75188 194566 75200
rect 269114 75188 269120 75200
rect 194560 75160 269120 75188
rect 194560 75148 194566 75160
rect 269114 75148 269120 75160
rect 269172 75148 269178 75200
rect 135622 75080 135628 75132
rect 135680 75120 135686 75132
rect 136542 75120 136548 75132
rect 135680 75092 136548 75120
rect 135680 75080 135686 75092
rect 136542 75080 136548 75092
rect 136600 75080 136606 75132
rect 139578 75080 139584 75132
rect 139636 75120 139642 75132
rect 140314 75120 140320 75132
rect 139636 75092 140320 75120
rect 139636 75080 139642 75092
rect 140314 75080 140320 75092
rect 140372 75080 140378 75132
rect 141050 75080 141056 75132
rect 141108 75120 141114 75132
rect 141878 75120 141884 75132
rect 141108 75092 141884 75120
rect 141108 75080 141114 75092
rect 141878 75080 141884 75092
rect 141936 75080 141942 75132
rect 153746 75080 153752 75132
rect 153804 75120 153810 75132
rect 216122 75120 216128 75132
rect 153804 75092 216128 75120
rect 153804 75080 153810 75092
rect 216122 75080 216128 75092
rect 216180 75080 216186 75132
rect 141786 75052 141792 75064
rect 137986 75024 141792 75052
rect 93670 74944 93676 74996
rect 93728 74984 93734 74996
rect 137986 74984 138014 75024
rect 141786 75012 141792 75024
rect 141844 75012 141850 75064
rect 158990 75012 158996 75064
rect 159048 75052 159054 75064
rect 160002 75052 160008 75064
rect 159048 75024 160008 75052
rect 159048 75012 159054 75024
rect 160002 75012 160008 75024
rect 160060 75012 160066 75064
rect 162854 75012 162860 75064
rect 162912 75052 162918 75064
rect 163498 75052 163504 75064
rect 162912 75024 163504 75052
rect 162912 75012 162918 75024
rect 163498 75012 163504 75024
rect 163556 75012 163562 75064
rect 170582 75012 170588 75064
rect 170640 75052 170646 75064
rect 214374 75052 214380 75064
rect 170640 75024 214380 75052
rect 170640 75012 170646 75024
rect 214374 75012 214380 75024
rect 214432 75012 214438 75064
rect 93728 74956 138014 74984
rect 93728 74944 93734 74956
rect 139578 74944 139584 74996
rect 139636 74984 139642 74996
rect 140682 74984 140688 74996
rect 139636 74956 140688 74984
rect 139636 74944 139642 74956
rect 140682 74944 140688 74956
rect 140740 74944 140746 74996
rect 145558 74944 145564 74996
rect 145616 74984 145622 74996
rect 146110 74984 146116 74996
rect 145616 74956 146116 74984
rect 145616 74944 145622 74956
rect 146110 74944 146116 74956
rect 146168 74944 146174 74996
rect 173066 74944 173072 74996
rect 173124 74984 173130 74996
rect 193214 74984 193220 74996
rect 173124 74956 193220 74984
rect 173124 74944 173130 74956
rect 193214 74944 193220 74956
rect 193272 74944 193278 74996
rect 95694 74876 95700 74928
rect 95752 74916 95758 74928
rect 145374 74916 145380 74928
rect 95752 74888 145380 74916
rect 95752 74876 95758 74888
rect 145374 74876 145380 74888
rect 145432 74876 145438 74928
rect 162578 74876 162584 74928
rect 162636 74916 162642 74928
rect 181346 74916 181352 74928
rect 162636 74888 181352 74916
rect 162636 74876 162642 74888
rect 181346 74876 181352 74888
rect 181404 74876 181410 74928
rect 140498 74808 140504 74860
rect 140556 74848 140562 74860
rect 147214 74848 147220 74860
rect 140556 74820 147220 74848
rect 140556 74808 140562 74820
rect 147214 74808 147220 74820
rect 147272 74808 147278 74860
rect 170030 74808 170036 74860
rect 170088 74848 170094 74860
rect 172146 74848 172152 74860
rect 170088 74820 172152 74848
rect 170088 74808 170094 74820
rect 172146 74808 172152 74820
rect 172204 74808 172210 74860
rect 107010 74740 107016 74792
rect 107068 74780 107074 74792
rect 107470 74780 107476 74792
rect 107068 74752 107476 74780
rect 107068 74740 107074 74752
rect 107470 74740 107476 74752
rect 107528 74740 107534 74792
rect 128906 74740 128912 74792
rect 128964 74780 128970 74792
rect 137922 74780 137928 74792
rect 128964 74752 137928 74780
rect 128964 74740 128970 74752
rect 137922 74740 137928 74752
rect 137980 74740 137986 74792
rect 151814 74740 151820 74792
rect 151872 74780 151878 74792
rect 154206 74780 154212 74792
rect 151872 74752 154212 74780
rect 151872 74740 151878 74752
rect 154206 74740 154212 74752
rect 154264 74740 154270 74792
rect 107470 74604 107476 74656
rect 107528 74644 107534 74656
rect 107654 74644 107660 74656
rect 107528 74616 107660 74644
rect 107528 74604 107534 74616
rect 107654 74604 107660 74616
rect 107712 74604 107718 74656
rect 137278 74604 137284 74656
rect 137336 74644 137342 74656
rect 142798 74644 142804 74656
rect 137336 74616 142804 74644
rect 137336 74604 137342 74616
rect 142798 74604 142804 74616
rect 142856 74604 142862 74656
rect 101858 74468 101864 74520
rect 101916 74508 101922 74520
rect 106274 74508 106280 74520
rect 101916 74480 106280 74508
rect 101916 74468 101922 74480
rect 106274 74468 106280 74480
rect 106332 74468 106338 74520
rect 118142 74468 118148 74520
rect 118200 74508 118206 74520
rect 140406 74508 140412 74520
rect 118200 74480 140412 74508
rect 118200 74468 118206 74480
rect 140406 74468 140412 74480
rect 140464 74468 140470 74520
rect 169478 74468 169484 74520
rect 169536 74508 169542 74520
rect 193858 74508 193864 74520
rect 169536 74480 193864 74508
rect 169536 74468 169542 74480
rect 193858 74468 193864 74480
rect 193916 74468 193922 74520
rect 97626 74400 97632 74452
rect 97684 74440 97690 74452
rect 157702 74440 157708 74452
rect 97684 74412 157708 74440
rect 97684 74400 97690 74412
rect 157702 74400 157708 74412
rect 157760 74400 157766 74452
rect 163314 74400 163320 74452
rect 163372 74440 163378 74452
rect 216858 74440 216864 74452
rect 163372 74412 216864 74440
rect 163372 74400 163378 74412
rect 216858 74400 216864 74412
rect 216916 74400 216922 74452
rect 114002 74332 114008 74384
rect 114060 74372 114066 74384
rect 143810 74372 143816 74384
rect 114060 74344 143816 74372
rect 114060 74332 114066 74344
rect 143810 74332 143816 74344
rect 143868 74332 143874 74384
rect 172054 74332 172060 74384
rect 172112 74372 172118 74384
rect 215386 74372 215392 74384
rect 172112 74344 215392 74372
rect 172112 74332 172118 74344
rect 215386 74332 215392 74344
rect 215444 74332 215450 74384
rect 118418 74264 118424 74316
rect 118476 74304 118482 74316
rect 152642 74304 152648 74316
rect 118476 74276 152648 74304
rect 118476 74264 118482 74276
rect 152642 74264 152648 74276
rect 152700 74264 152706 74316
rect 164602 74264 164608 74316
rect 164660 74304 164666 74316
rect 200390 74304 200396 74316
rect 164660 74276 200396 74304
rect 164660 74264 164666 74276
rect 200390 74264 200396 74276
rect 200448 74264 200454 74316
rect 117222 74196 117228 74248
rect 117280 74236 117286 74248
rect 150710 74236 150716 74248
rect 117280 74208 150716 74236
rect 117280 74196 117286 74208
rect 150710 74196 150716 74208
rect 150768 74196 150774 74248
rect 154666 74196 154672 74248
rect 154724 74236 154730 74248
rect 155402 74236 155408 74248
rect 154724 74208 155408 74236
rect 154724 74196 154730 74208
rect 155402 74196 155408 74208
rect 155460 74196 155466 74248
rect 161474 74196 161480 74248
rect 161532 74236 161538 74248
rect 162486 74236 162492 74248
rect 161532 74208 162492 74236
rect 161532 74196 161538 74208
rect 162486 74196 162492 74208
rect 162544 74196 162550 74248
rect 177850 74196 177856 74248
rect 177908 74236 177914 74248
rect 208946 74236 208952 74248
rect 177908 74208 208952 74236
rect 177908 74196 177914 74208
rect 208946 74196 208952 74208
rect 209004 74196 209010 74248
rect 108758 74128 108764 74180
rect 108816 74168 108822 74180
rect 142246 74168 142252 74180
rect 108816 74140 142252 74168
rect 108816 74128 108822 74140
rect 142246 74128 142252 74140
rect 142304 74128 142310 74180
rect 169018 74128 169024 74180
rect 169076 74168 169082 74180
rect 195054 74168 195060 74180
rect 169076 74140 195060 74168
rect 169076 74128 169082 74140
rect 195054 74128 195060 74140
rect 195112 74128 195118 74180
rect 112530 74060 112536 74112
rect 112588 74100 112594 74112
rect 146110 74100 146116 74112
rect 112588 74072 146116 74100
rect 112588 74060 112594 74072
rect 146110 74060 146116 74072
rect 146168 74060 146174 74112
rect 163774 74060 163780 74112
rect 163832 74100 163838 74112
rect 197998 74100 198004 74112
rect 163832 74072 198004 74100
rect 163832 74060 163838 74072
rect 197998 74060 198004 74072
rect 198056 74060 198062 74112
rect 102686 73992 102692 74044
rect 102744 74032 102750 74044
rect 135806 74032 135812 74044
rect 102744 74004 135812 74032
rect 102744 73992 102750 74004
rect 135806 73992 135812 74004
rect 135864 73992 135870 74044
rect 145098 73992 145104 74044
rect 145156 74032 145162 74044
rect 145558 74032 145564 74044
rect 145156 74004 145564 74032
rect 145156 73992 145162 74004
rect 145558 73992 145564 74004
rect 145616 73992 145622 74044
rect 145650 73992 145656 74044
rect 145708 74032 145714 74044
rect 145926 74032 145932 74044
rect 145708 74004 145932 74032
rect 145708 73992 145714 74004
rect 145926 73992 145932 74004
rect 145984 73992 145990 74044
rect 149330 73992 149336 74044
rect 149388 74032 149394 74044
rect 149882 74032 149888 74044
rect 149388 74004 149888 74032
rect 149388 73992 149394 74004
rect 149882 73992 149888 74004
rect 149940 73992 149946 74044
rect 173434 73992 173440 74044
rect 173492 74032 173498 74044
rect 206186 74032 206192 74044
rect 173492 74004 206192 74032
rect 173492 73992 173498 74004
rect 206186 73992 206192 74004
rect 206244 73992 206250 74044
rect 111334 73924 111340 73976
rect 111392 73964 111398 73976
rect 142614 73964 142620 73976
rect 111392 73936 142620 73964
rect 111392 73924 111398 73936
rect 142614 73924 142620 73936
rect 142672 73924 142678 73976
rect 174722 73924 174728 73976
rect 174780 73964 174786 73976
rect 207014 73964 207020 73976
rect 174780 73936 207020 73964
rect 174780 73924 174786 73936
rect 207014 73924 207020 73936
rect 207072 73924 207078 73976
rect 74534 73856 74540 73908
rect 74592 73896 74598 73908
rect 117222 73896 117228 73908
rect 74592 73868 117228 73896
rect 74592 73856 74598 73868
rect 117222 73856 117228 73868
rect 117280 73856 117286 73908
rect 152458 73856 152464 73908
rect 152516 73896 152522 73908
rect 162670 73896 162676 73908
rect 152516 73868 162676 73896
rect 152516 73856 152522 73868
rect 162670 73856 162676 73868
rect 162728 73856 162734 73908
rect 189166 73856 189172 73908
rect 189224 73896 189230 73908
rect 189810 73896 189816 73908
rect 189224 73868 189816 73896
rect 189224 73856 189230 73868
rect 189810 73856 189816 73868
rect 189868 73896 189874 73908
rect 321554 73896 321560 73908
rect 189868 73868 321560 73896
rect 189868 73856 189874 73868
rect 321554 73856 321560 73868
rect 321612 73856 321618 73908
rect 35158 73788 35164 73840
rect 35216 73828 35222 73840
rect 100294 73828 100300 73840
rect 35216 73800 100300 73828
rect 35216 73788 35222 73800
rect 100294 73788 100300 73800
rect 100352 73788 100358 73840
rect 115290 73788 115296 73840
rect 115348 73828 115354 73840
rect 145098 73828 145104 73840
rect 115348 73800 145104 73828
rect 115348 73788 115354 73800
rect 145098 73788 145104 73800
rect 145156 73788 145162 73840
rect 161290 73788 161296 73840
rect 161348 73828 161354 73840
rect 184934 73828 184940 73840
rect 161348 73800 184940 73828
rect 161348 73788 161354 73800
rect 184934 73788 184940 73800
rect 184992 73788 184998 73840
rect 215386 73788 215392 73840
rect 215444 73828 215450 73840
rect 560938 73828 560944 73840
rect 215444 73800 560944 73828
rect 215444 73788 215450 73800
rect 560938 73788 560944 73800
rect 560996 73788 561002 73840
rect 112622 73720 112628 73772
rect 112680 73760 112686 73772
rect 138198 73760 138204 73772
rect 112680 73732 138204 73760
rect 112680 73720 112686 73732
rect 138198 73720 138204 73732
rect 138256 73760 138262 73772
rect 138842 73760 138848 73772
rect 138256 73732 138848 73760
rect 138256 73720 138262 73732
rect 138842 73720 138848 73732
rect 138900 73720 138906 73772
rect 149698 73720 149704 73772
rect 149756 73760 149762 73772
rect 221274 73760 221280 73772
rect 149756 73732 221280 73760
rect 149756 73720 149762 73732
rect 221274 73720 221280 73732
rect 221332 73720 221338 73772
rect 115198 73652 115204 73704
rect 115256 73692 115262 73704
rect 151262 73692 151268 73704
rect 115256 73664 151268 73692
rect 115256 73652 115262 73664
rect 151262 73652 151268 73664
rect 151320 73652 151326 73704
rect 154574 73652 154580 73704
rect 154632 73692 154638 73704
rect 189166 73692 189172 73704
rect 154632 73664 189172 73692
rect 154632 73652 154638 73664
rect 189166 73652 189172 73664
rect 189224 73652 189230 73704
rect 100294 73584 100300 73636
rect 100352 73624 100358 73636
rect 135162 73624 135168 73636
rect 100352 73596 135168 73624
rect 100352 73584 100358 73596
rect 135162 73584 135168 73596
rect 135220 73584 135226 73636
rect 106274 73516 106280 73568
rect 106332 73556 106338 73568
rect 107470 73556 107476 73568
rect 106332 73528 107476 73556
rect 106332 73516 106338 73528
rect 107470 73516 107476 73528
rect 107528 73516 107534 73568
rect 131758 73448 131764 73500
rect 131816 73488 131822 73500
rect 137738 73488 137744 73500
rect 131816 73460 137744 73488
rect 131816 73448 131822 73460
rect 137738 73448 137744 73460
rect 137796 73448 137802 73500
rect 153378 73312 153384 73364
rect 153436 73352 153442 73364
rect 154022 73352 154028 73364
rect 153436 73324 154028 73352
rect 153436 73312 153442 73324
rect 154022 73312 154028 73324
rect 154080 73312 154086 73364
rect 149330 73176 149336 73228
rect 149388 73216 149394 73228
rect 182818 73216 182824 73228
rect 149388 73188 182824 73216
rect 149388 73176 149394 73188
rect 182818 73176 182824 73188
rect 182876 73176 182882 73228
rect 3142 73108 3148 73160
rect 3200 73148 3206 73160
rect 152458 73148 152464 73160
rect 3200 73120 152464 73148
rect 3200 73108 3206 73120
rect 152458 73108 152464 73120
rect 152516 73108 152522 73160
rect 171870 73108 171876 73160
rect 171928 73148 171934 73160
rect 197354 73148 197360 73160
rect 171928 73120 197360 73148
rect 171928 73108 171934 73120
rect 197354 73108 197360 73120
rect 197412 73108 197418 73160
rect 218054 73108 218060 73160
rect 218112 73148 218118 73160
rect 218606 73148 218612 73160
rect 218112 73120 218612 73148
rect 218112 73108 218118 73120
rect 218606 73108 218612 73120
rect 218664 73148 218670 73160
rect 580166 73148 580172 73160
rect 218664 73120 580172 73148
rect 218664 73108 218670 73120
rect 580166 73108 580172 73120
rect 580224 73108 580230 73160
rect 121086 73040 121092 73092
rect 121144 73080 121150 73092
rect 121144 73052 149744 73080
rect 121144 73040 121150 73052
rect 114830 72972 114836 73024
rect 114888 73012 114894 73024
rect 149238 73012 149244 73024
rect 114888 72984 149244 73012
rect 114888 72972 114894 72984
rect 149238 72972 149244 72984
rect 149296 72972 149302 73024
rect 149716 73012 149744 73052
rect 149790 73040 149796 73092
rect 149848 73080 149854 73092
rect 150342 73080 150348 73092
rect 149848 73052 150348 73080
rect 149848 73040 149854 73052
rect 150342 73040 150348 73052
rect 150400 73040 150406 73092
rect 171042 73040 171048 73092
rect 171100 73080 171106 73092
rect 195974 73080 195980 73092
rect 171100 73052 195980 73080
rect 171100 73040 171106 73052
rect 195974 73040 195980 73052
rect 196032 73040 196038 73092
rect 157150 73012 157156 73024
rect 149716 72984 157156 73012
rect 157150 72972 157156 72984
rect 157208 72972 157214 73024
rect 173894 72972 173900 73024
rect 173952 73012 173958 73024
rect 200482 73012 200488 73024
rect 173952 72984 200488 73012
rect 173952 72972 173958 72984
rect 200482 72972 200488 72984
rect 200540 72972 200546 73024
rect 119890 72904 119896 72956
rect 119948 72944 119954 72956
rect 152274 72944 152280 72956
rect 119948 72916 152280 72944
rect 119948 72904 119954 72916
rect 152274 72904 152280 72916
rect 152332 72904 152338 72956
rect 156506 72904 156512 72956
rect 156564 72944 156570 72956
rect 190914 72944 190920 72956
rect 156564 72916 190920 72944
rect 156564 72904 156570 72916
rect 190914 72904 190920 72916
rect 190972 72904 190978 72956
rect 126238 72836 126244 72888
rect 126296 72876 126302 72888
rect 153010 72876 153016 72888
rect 126296 72848 153016 72876
rect 126296 72836 126302 72848
rect 153010 72836 153016 72848
rect 153068 72836 153074 72888
rect 161382 72836 161388 72888
rect 161440 72876 161446 72888
rect 194962 72876 194968 72888
rect 161440 72848 194968 72876
rect 161440 72836 161446 72848
rect 194962 72836 194968 72848
rect 195020 72836 195026 72888
rect 114094 72768 114100 72820
rect 114152 72808 114158 72820
rect 148778 72808 148784 72820
rect 114152 72780 148784 72808
rect 114152 72768 114158 72780
rect 148778 72768 148784 72780
rect 148836 72768 148842 72820
rect 162762 72768 162768 72820
rect 162820 72808 162826 72820
rect 163958 72808 163964 72820
rect 162820 72780 163964 72808
rect 162820 72768 162826 72780
rect 163958 72768 163964 72780
rect 164016 72768 164022 72820
rect 167914 72768 167920 72820
rect 167972 72808 167978 72820
rect 201954 72808 201960 72820
rect 167972 72780 201960 72808
rect 167972 72768 167978 72780
rect 201954 72768 201960 72780
rect 202012 72808 202018 72820
rect 202012 72780 209774 72808
rect 202012 72768 202018 72780
rect 114922 72700 114928 72752
rect 114980 72740 114986 72752
rect 149054 72740 149060 72752
rect 114980 72712 149060 72740
rect 114980 72700 114986 72712
rect 149054 72700 149060 72712
rect 149112 72700 149118 72752
rect 163406 72700 163412 72752
rect 163464 72740 163470 72752
rect 197722 72740 197728 72752
rect 163464 72712 197728 72740
rect 163464 72700 163470 72712
rect 197722 72700 197728 72712
rect 197780 72700 197786 72752
rect 111702 72632 111708 72684
rect 111760 72672 111766 72684
rect 143534 72672 143540 72684
rect 111760 72644 143540 72672
rect 111760 72632 111766 72644
rect 143534 72632 143540 72644
rect 143592 72632 143598 72684
rect 153562 72632 153568 72684
rect 153620 72672 153626 72684
rect 158346 72672 158352 72684
rect 153620 72644 158352 72672
rect 153620 72632 153626 72644
rect 158346 72632 158352 72644
rect 158404 72632 158410 72684
rect 177942 72632 177948 72684
rect 178000 72672 178006 72684
rect 208394 72672 208400 72684
rect 178000 72644 208400 72672
rect 178000 72632 178006 72644
rect 208394 72632 208400 72644
rect 208452 72632 208458 72684
rect 120902 72564 120908 72616
rect 120960 72604 120966 72616
rect 151814 72604 151820 72616
rect 120960 72576 151820 72604
rect 120960 72564 120966 72576
rect 151814 72564 151820 72576
rect 151872 72564 151878 72616
rect 173710 72564 173716 72616
rect 173768 72604 173774 72616
rect 204898 72604 204904 72616
rect 173768 72576 204904 72604
rect 173768 72564 173774 72576
rect 204898 72564 204904 72576
rect 204956 72564 204962 72616
rect 115382 72496 115388 72548
rect 115440 72536 115446 72548
rect 146938 72536 146944 72548
rect 115440 72508 146944 72536
rect 115440 72496 115446 72508
rect 146938 72496 146944 72508
rect 146996 72496 147002 72548
rect 159910 72496 159916 72548
rect 159968 72536 159974 72548
rect 193490 72536 193496 72548
rect 159968 72508 193496 72536
rect 159968 72496 159974 72508
rect 193490 72496 193496 72508
rect 193548 72496 193554 72548
rect 52454 72428 52460 72480
rect 52512 72468 52518 72480
rect 98822 72468 98828 72480
rect 52512 72440 98828 72468
rect 52512 72428 52518 72440
rect 98822 72428 98828 72440
rect 98880 72428 98886 72480
rect 124214 72428 124220 72480
rect 124272 72468 124278 72480
rect 175458 72468 175464 72480
rect 124272 72440 175464 72468
rect 124272 72428 124278 72440
rect 175458 72428 175464 72440
rect 175516 72428 175522 72480
rect 184934 72428 184940 72480
rect 184992 72468 184998 72480
rect 186222 72468 186228 72480
rect 184992 72440 186228 72468
rect 184992 72428 184998 72440
rect 186222 72428 186228 72440
rect 186280 72468 186286 72480
rect 194594 72468 194600 72480
rect 186280 72440 194600 72468
rect 186280 72428 186286 72440
rect 194594 72428 194600 72440
rect 194652 72428 194658 72480
rect 209746 72468 209774 72780
rect 253934 72468 253940 72480
rect 209746 72440 253940 72468
rect 253934 72428 253940 72440
rect 253992 72428 253998 72480
rect 119982 72360 119988 72412
rect 120040 72400 120046 72412
rect 149790 72400 149796 72412
rect 120040 72372 149796 72400
rect 120040 72360 120046 72372
rect 149790 72360 149796 72372
rect 149848 72360 149854 72412
rect 155586 72360 155592 72412
rect 155644 72400 155650 72412
rect 218054 72400 218060 72412
rect 155644 72372 218060 72400
rect 155644 72360 155650 72372
rect 218054 72360 218060 72372
rect 218112 72360 218118 72412
rect 98822 72292 98828 72344
rect 98880 72332 98886 72344
rect 133138 72332 133144 72344
rect 98880 72304 133144 72332
rect 98880 72292 98886 72304
rect 133138 72292 133144 72304
rect 133196 72292 133202 72344
rect 161106 72292 161112 72344
rect 161164 72332 161170 72344
rect 195146 72332 195152 72344
rect 161164 72304 195152 72332
rect 161164 72292 161170 72304
rect 195146 72292 195152 72304
rect 195204 72292 195210 72344
rect 98730 72224 98736 72276
rect 98788 72264 98794 72276
rect 133874 72264 133880 72276
rect 98788 72236 133880 72264
rect 98788 72224 98794 72236
rect 133874 72224 133880 72236
rect 133932 72224 133938 72276
rect 157426 72224 157432 72276
rect 157484 72264 157490 72276
rect 192386 72264 192392 72276
rect 157484 72236 192392 72264
rect 157484 72224 157490 72236
rect 192386 72224 192392 72236
rect 192444 72224 192450 72276
rect 133138 72156 133144 72208
rect 133196 72196 133202 72208
rect 133598 72196 133604 72208
rect 133196 72168 133604 72196
rect 133196 72156 133202 72168
rect 133598 72156 133604 72168
rect 133656 72156 133662 72208
rect 165522 72156 165528 72208
rect 165580 72196 165586 72208
rect 184198 72196 184204 72208
rect 165580 72168 184204 72196
rect 165580 72156 165586 72168
rect 184198 72156 184204 72168
rect 184256 72156 184262 72208
rect 121730 71680 121736 71732
rect 121788 71720 121794 71732
rect 142982 71720 142988 71732
rect 121788 71692 142988 71720
rect 121788 71680 121794 71692
rect 142982 71680 142988 71692
rect 143040 71680 143046 71732
rect 148410 71680 148416 71732
rect 148468 71720 148474 71732
rect 148686 71720 148692 71732
rect 148468 71692 148692 71720
rect 148468 71680 148474 71692
rect 148686 71680 148692 71692
rect 148744 71680 148750 71732
rect 158622 71680 158628 71732
rect 158680 71720 158686 71732
rect 219710 71720 219716 71732
rect 158680 71692 219716 71720
rect 158680 71680 158686 71692
rect 219710 71680 219716 71692
rect 219768 71680 219774 71732
rect 116854 71612 116860 71664
rect 116912 71652 116918 71664
rect 151354 71652 151360 71664
rect 116912 71624 151360 71652
rect 116912 71612 116918 71624
rect 151354 71612 151360 71624
rect 151412 71652 151418 71664
rect 151722 71652 151728 71664
rect 151412 71624 151728 71652
rect 151412 71612 151418 71624
rect 151722 71612 151728 71624
rect 151780 71612 151786 71664
rect 172238 71612 172244 71664
rect 172296 71652 172302 71664
rect 215846 71652 215852 71664
rect 172296 71624 215852 71652
rect 172296 71612 172302 71624
rect 215846 71612 215852 71624
rect 215904 71612 215910 71664
rect 123478 71544 123484 71596
rect 123536 71584 123542 71596
rect 142890 71584 142896 71596
rect 123536 71556 142896 71584
rect 123536 71544 123542 71556
rect 142890 71544 142896 71556
rect 142948 71544 142954 71596
rect 175182 71584 175188 71596
rect 157306 71556 175188 71584
rect 111058 71476 111064 71528
rect 111116 71516 111122 71528
rect 141694 71516 141700 71528
rect 111116 71488 141700 71516
rect 111116 71476 111122 71488
rect 141694 71476 141700 71488
rect 141752 71476 141758 71528
rect 115658 71408 115664 71460
rect 115716 71448 115722 71460
rect 147674 71448 147680 71460
rect 115716 71420 147680 71448
rect 115716 71408 115722 71420
rect 147674 71408 147680 71420
rect 147732 71448 147738 71460
rect 148318 71448 148324 71460
rect 147732 71420 148324 71448
rect 147732 71408 147738 71420
rect 148318 71408 148324 71420
rect 148376 71408 148382 71460
rect 117038 71340 117044 71392
rect 117096 71380 117102 71392
rect 148410 71380 148416 71392
rect 117096 71352 148416 71380
rect 117096 71340 117102 71352
rect 148410 71340 148416 71352
rect 148468 71340 148474 71392
rect 108850 71272 108856 71324
rect 108908 71312 108914 71324
rect 139118 71312 139124 71324
rect 108908 71284 139124 71312
rect 108908 71272 108914 71284
rect 139118 71272 139124 71284
rect 139176 71272 139182 71324
rect 106734 71204 106740 71256
rect 106792 71244 106798 71256
rect 130838 71244 130844 71256
rect 106792 71216 130844 71244
rect 106792 71204 106798 71216
rect 130838 71204 130844 71216
rect 130896 71204 130902 71256
rect 153102 71204 153108 71256
rect 153160 71244 153166 71256
rect 157306 71244 157334 71556
rect 175182 71544 175188 71556
rect 175240 71584 175246 71596
rect 197630 71584 197636 71596
rect 175240 71556 197636 71584
rect 175240 71544 175246 71556
rect 197630 71544 197636 71556
rect 197688 71544 197694 71596
rect 172698 71476 172704 71528
rect 172756 71516 172762 71528
rect 207382 71516 207388 71528
rect 172756 71488 207388 71516
rect 172756 71476 172762 71488
rect 207382 71476 207388 71488
rect 207440 71476 207446 71528
rect 176930 71408 176936 71460
rect 176988 71448 176994 71460
rect 210142 71448 210148 71460
rect 176988 71420 210148 71448
rect 176988 71408 176994 71420
rect 210142 71408 210148 71420
rect 210200 71408 210206 71460
rect 176746 71340 176752 71392
rect 176804 71380 176810 71392
rect 209866 71380 209872 71392
rect 176804 71352 209872 71380
rect 176804 71340 176810 71352
rect 209866 71340 209872 71352
rect 209924 71340 209930 71392
rect 172146 71272 172152 71324
rect 172204 71312 172210 71324
rect 204438 71312 204444 71324
rect 172204 71284 204444 71312
rect 172204 71272 172210 71284
rect 204438 71272 204444 71284
rect 204496 71272 204502 71324
rect 153160 71216 157334 71244
rect 153160 71204 153166 71216
rect 176102 71204 176108 71256
rect 176160 71244 176166 71256
rect 207290 71244 207296 71256
rect 176160 71216 207296 71244
rect 176160 71204 176166 71216
rect 207290 71204 207296 71216
rect 207348 71204 207354 71256
rect 110966 71136 110972 71188
rect 111024 71176 111030 71188
rect 137186 71176 137192 71188
rect 111024 71148 137192 71176
rect 111024 71136 111030 71148
rect 137186 71136 137192 71148
rect 137244 71136 137250 71188
rect 171502 71136 171508 71188
rect 171560 71176 171566 71188
rect 202874 71176 202880 71188
rect 171560 71148 202880 71176
rect 171560 71136 171566 71148
rect 202874 71136 202880 71148
rect 202932 71136 202938 71188
rect 151722 71068 151728 71120
rect 151780 71108 151786 71120
rect 306374 71108 306380 71120
rect 151780 71080 306380 71108
rect 151780 71068 151786 71080
rect 306374 71068 306380 71080
rect 306432 71068 306438 71120
rect 2774 71000 2780 71052
rect 2832 71040 2838 71052
rect 157426 71040 157432 71052
rect 2832 71012 157432 71040
rect 2832 71000 2838 71012
rect 157426 71000 157432 71012
rect 157484 71000 157490 71052
rect 176010 71000 176016 71052
rect 176068 71040 176074 71052
rect 176286 71040 176292 71052
rect 176068 71012 176292 71040
rect 176068 71000 176074 71012
rect 176286 71000 176292 71012
rect 176344 71040 176350 71052
rect 206462 71040 206468 71052
rect 176344 71012 206468 71040
rect 176344 71000 176350 71012
rect 206462 71000 206468 71012
rect 206520 71000 206526 71052
rect 215846 71000 215852 71052
rect 215904 71040 215910 71052
rect 484394 71040 484400 71052
rect 215904 71012 484400 71040
rect 215904 71000 215910 71012
rect 484394 71000 484400 71012
rect 484452 71000 484458 71052
rect 93762 70932 93768 70984
rect 93820 70972 93826 70984
rect 156966 70972 156972 70984
rect 93820 70944 156972 70972
rect 93820 70932 93826 70944
rect 156966 70932 156972 70944
rect 157024 70932 157030 70984
rect 180242 70932 180248 70984
rect 180300 70972 180306 70984
rect 188982 70972 188988 70984
rect 180300 70944 188988 70972
rect 180300 70932 180306 70944
rect 188982 70932 188988 70944
rect 189040 70972 189046 70984
rect 207750 70972 207756 70984
rect 189040 70944 207756 70972
rect 189040 70932 189046 70944
rect 207750 70932 207756 70944
rect 207808 70932 207814 70984
rect 114186 70864 114192 70916
rect 114244 70904 114250 70916
rect 147122 70904 147128 70916
rect 114244 70876 147128 70904
rect 114244 70864 114250 70876
rect 147122 70864 147128 70876
rect 147180 70864 147186 70916
rect 156322 70864 156328 70916
rect 156380 70904 156386 70916
rect 192018 70904 192024 70916
rect 156380 70876 192024 70904
rect 156380 70864 156386 70876
rect 192018 70864 192024 70876
rect 192076 70864 192082 70916
rect 106826 70796 106832 70848
rect 106884 70836 106890 70848
rect 132402 70836 132408 70848
rect 106884 70808 132408 70836
rect 106884 70796 106890 70808
rect 132402 70796 132408 70808
rect 132460 70796 132466 70848
rect 127618 70728 127624 70780
rect 127676 70768 127682 70780
rect 150526 70768 150532 70780
rect 127676 70740 150532 70768
rect 127676 70728 127682 70740
rect 150526 70728 150532 70740
rect 150584 70728 150590 70780
rect 160462 70728 160468 70780
rect 160520 70768 160526 70780
rect 161382 70768 161388 70780
rect 160520 70740 161388 70768
rect 160520 70728 160526 70740
rect 161382 70728 161388 70740
rect 161440 70728 161446 70780
rect 108942 70320 108948 70372
rect 109000 70360 109006 70372
rect 135898 70360 135904 70372
rect 109000 70332 135904 70360
rect 109000 70320 109006 70332
rect 135898 70320 135904 70332
rect 135956 70320 135962 70372
rect 166166 70320 166172 70372
rect 166224 70360 166230 70372
rect 207842 70360 207848 70372
rect 166224 70332 207848 70360
rect 166224 70320 166230 70332
rect 207842 70320 207848 70332
rect 207900 70320 207906 70372
rect 118602 70252 118608 70304
rect 118660 70292 118666 70304
rect 150986 70292 150992 70304
rect 118660 70264 150992 70292
rect 118660 70252 118666 70264
rect 150986 70252 150992 70264
rect 151044 70252 151050 70304
rect 164694 70252 164700 70304
rect 164752 70292 164758 70304
rect 199470 70292 199476 70304
rect 164752 70264 199476 70292
rect 164752 70252 164758 70264
rect 199470 70252 199476 70264
rect 199528 70252 199534 70304
rect 109770 70184 109776 70236
rect 109828 70224 109834 70236
rect 151170 70224 151176 70236
rect 109828 70196 151176 70224
rect 109828 70184 109834 70196
rect 151170 70184 151176 70196
rect 151228 70184 151234 70236
rect 175550 70184 175556 70236
rect 175608 70224 175614 70236
rect 210234 70224 210240 70236
rect 175608 70196 210240 70224
rect 175608 70184 175614 70196
rect 210234 70184 210240 70196
rect 210292 70184 210298 70236
rect 115566 70116 115572 70168
rect 115624 70156 115630 70168
rect 149330 70156 149336 70168
rect 115624 70128 149336 70156
rect 115624 70116 115630 70128
rect 149330 70116 149336 70128
rect 149388 70116 149394 70168
rect 167086 70116 167092 70168
rect 167144 70156 167150 70168
rect 167454 70156 167460 70168
rect 167144 70128 167460 70156
rect 167144 70116 167150 70128
rect 167454 70116 167460 70128
rect 167512 70156 167518 70168
rect 202138 70156 202144 70168
rect 167512 70128 202144 70156
rect 167512 70116 167518 70128
rect 202138 70116 202144 70128
rect 202196 70116 202202 70168
rect 117958 70048 117964 70100
rect 118016 70088 118022 70100
rect 152918 70088 152924 70100
rect 118016 70060 152924 70088
rect 118016 70048 118022 70060
rect 152918 70048 152924 70060
rect 152976 70048 152982 70100
rect 157610 70048 157616 70100
rect 157668 70088 157674 70100
rect 158530 70088 158536 70100
rect 157668 70060 158536 70088
rect 157668 70048 157674 70060
rect 158530 70048 158536 70060
rect 158588 70088 158594 70100
rect 192202 70088 192208 70100
rect 158588 70060 192208 70088
rect 158588 70048 158594 70060
rect 192202 70048 192208 70060
rect 192260 70048 192266 70100
rect 122006 69980 122012 70032
rect 122064 70020 122070 70032
rect 156690 70020 156696 70032
rect 122064 69992 156696 70020
rect 122064 69980 122070 69992
rect 156690 69980 156696 69992
rect 156748 69980 156754 70032
rect 160278 69980 160284 70032
rect 160336 70020 160342 70032
rect 161198 70020 161204 70032
rect 160336 69992 161204 70020
rect 160336 69980 160342 69992
rect 161198 69980 161204 69992
rect 161256 70020 161262 70032
rect 194778 70020 194784 70032
rect 161256 69992 194784 70020
rect 161256 69980 161262 69992
rect 194778 69980 194784 69992
rect 194836 69980 194842 70032
rect 99006 69912 99012 69964
rect 99064 69952 99070 69964
rect 133782 69952 133788 69964
rect 99064 69924 133788 69952
rect 99064 69912 99070 69924
rect 133782 69912 133788 69924
rect 133840 69912 133846 69964
rect 172514 69912 172520 69964
rect 172572 69952 172578 69964
rect 206094 69952 206100 69964
rect 172572 69924 206100 69952
rect 172572 69912 172578 69924
rect 206094 69912 206100 69924
rect 206152 69912 206158 69964
rect 108666 69844 108672 69896
rect 108724 69884 108730 69896
rect 141510 69884 141516 69896
rect 108724 69856 141516 69884
rect 108724 69844 108730 69856
rect 141510 69844 141516 69856
rect 141568 69844 141574 69896
rect 172606 69844 172612 69896
rect 172664 69884 172670 69896
rect 173158 69884 173164 69896
rect 172664 69856 173164 69884
rect 172664 69844 172670 69856
rect 173158 69844 173164 69856
rect 173216 69884 173222 69896
rect 205818 69884 205824 69896
rect 173216 69856 205824 69884
rect 173216 69844 173222 69856
rect 205818 69844 205824 69856
rect 205876 69844 205882 69896
rect 113818 69776 113824 69828
rect 113876 69816 113882 69828
rect 147398 69816 147404 69828
rect 113876 69788 147404 69816
rect 113876 69776 113882 69788
rect 147398 69776 147404 69788
rect 147456 69776 147462 69828
rect 157702 69776 157708 69828
rect 157760 69816 157766 69828
rect 158622 69816 158628 69828
rect 157760 69788 158628 69816
rect 157760 69776 157766 69788
rect 158622 69776 158628 69788
rect 158680 69816 158686 69828
rect 190730 69816 190736 69828
rect 158680 69788 190736 69816
rect 158680 69776 158686 69788
rect 190730 69776 190736 69788
rect 190788 69776 190794 69828
rect 13078 69708 13084 69760
rect 13136 69748 13142 69760
rect 94958 69748 94964 69760
rect 13136 69720 94964 69748
rect 13136 69708 13142 69720
rect 94958 69708 94964 69720
rect 95016 69748 95022 69760
rect 95142 69748 95148 69760
rect 95016 69720 95148 69748
rect 95016 69708 95022 69720
rect 95142 69708 95148 69720
rect 95200 69708 95206 69760
rect 126238 69708 126244 69760
rect 126296 69748 126302 69760
rect 167086 69748 167092 69760
rect 126296 69720 167092 69748
rect 126296 69708 126302 69720
rect 167086 69708 167092 69720
rect 167144 69708 167150 69760
rect 172698 69708 172704 69760
rect 172756 69748 172762 69760
rect 198734 69748 198740 69760
rect 172756 69720 198740 69748
rect 172756 69708 172762 69720
rect 198734 69708 198740 69720
rect 198792 69748 198798 69760
rect 198792 69720 200114 69748
rect 198792 69708 198798 69720
rect 78674 69640 78680 69692
rect 78732 69680 78738 69692
rect 160462 69680 160468 69692
rect 78732 69652 160468 69680
rect 78732 69640 78738 69652
rect 160462 69640 160468 69652
rect 160520 69640 160526 69692
rect 166166 69640 166172 69692
rect 166224 69680 166230 69692
rect 197814 69680 197820 69692
rect 166224 69652 197820 69680
rect 166224 69640 166230 69652
rect 197814 69640 197820 69652
rect 197872 69640 197878 69692
rect 200086 69680 200114 69720
rect 314654 69680 314660 69692
rect 200086 69652 314660 69680
rect 314654 69640 314660 69652
rect 314712 69640 314718 69692
rect 108022 69572 108028 69624
rect 108080 69612 108086 69624
rect 152182 69612 152188 69624
rect 108080 69584 152188 69612
rect 108080 69572 108086 69584
rect 152182 69572 152188 69584
rect 152240 69572 152246 69624
rect 160370 69572 160376 69624
rect 160428 69612 160434 69624
rect 161382 69612 161388 69624
rect 160428 69584 161388 69612
rect 160428 69572 160434 69584
rect 161382 69572 161388 69584
rect 161440 69612 161446 69624
rect 192662 69612 192668 69624
rect 161440 69584 192668 69612
rect 161440 69572 161446 69584
rect 192662 69572 192668 69584
rect 192720 69572 192726 69624
rect 95142 69504 95148 69556
rect 95200 69544 95206 69556
rect 139210 69544 139216 69556
rect 95200 69516 139216 69544
rect 95200 69504 95206 69516
rect 139210 69504 139216 69516
rect 139268 69504 139274 69556
rect 162118 69504 162124 69556
rect 162176 69544 162182 69556
rect 162578 69544 162584 69556
rect 162176 69516 162584 69544
rect 162176 69504 162182 69516
rect 162578 69504 162584 69516
rect 162636 69504 162642 69556
rect 165154 69504 165160 69556
rect 165212 69544 165218 69556
rect 174538 69544 174544 69556
rect 165212 69516 174544 69544
rect 165212 69504 165218 69516
rect 174538 69504 174544 69516
rect 174596 69504 174602 69556
rect 164142 69436 164148 69488
rect 164200 69476 164206 69488
rect 181622 69476 181628 69488
rect 164200 69448 181628 69476
rect 164200 69436 164206 69448
rect 181622 69436 181628 69448
rect 181680 69436 181686 69488
rect 162578 69368 162584 69420
rect 162636 69408 162642 69420
rect 181530 69408 181536 69420
rect 162636 69380 181536 69408
rect 162636 69368 162642 69380
rect 181530 69368 181536 69380
rect 181588 69368 181594 69420
rect 107194 68960 107200 69012
rect 107252 69000 107258 69012
rect 136450 69000 136456 69012
rect 107252 68972 136456 69000
rect 107252 68960 107258 68972
rect 136450 68960 136456 68972
rect 136508 68960 136514 69012
rect 162026 68960 162032 69012
rect 162084 69000 162090 69012
rect 162670 69000 162676 69012
rect 162084 68972 162676 69000
rect 162084 68960 162090 68972
rect 162670 68960 162676 68972
rect 162728 68960 162734 69012
rect 163130 68960 163136 69012
rect 163188 69000 163194 69012
rect 164050 69000 164056 69012
rect 163188 68972 164056 69000
rect 163188 68960 163194 68972
rect 164050 68960 164056 68972
rect 164108 68960 164114 69012
rect 166626 68960 166632 69012
rect 166684 69000 166690 69012
rect 191098 69000 191104 69012
rect 166684 68972 191104 69000
rect 166684 68960 166690 68972
rect 191098 68960 191104 68972
rect 191156 68960 191162 69012
rect 111242 68892 111248 68944
rect 111300 68932 111306 68944
rect 138658 68932 138664 68944
rect 111300 68904 138664 68932
rect 111300 68892 111306 68904
rect 138658 68892 138664 68904
rect 138716 68892 138722 68944
rect 160186 68892 160192 68944
rect 160244 68932 160250 68944
rect 194870 68932 194876 68944
rect 160244 68904 194876 68932
rect 160244 68892 160250 68904
rect 194870 68892 194876 68904
rect 194928 68892 194934 68944
rect 110322 68824 110328 68876
rect 110380 68864 110386 68876
rect 156230 68864 156236 68876
rect 110380 68836 156236 68864
rect 110380 68824 110386 68836
rect 156230 68824 156236 68836
rect 156288 68824 156294 68876
rect 167362 68824 167368 68876
rect 167420 68864 167426 68876
rect 201862 68864 201868 68876
rect 167420 68836 201868 68864
rect 167420 68824 167426 68836
rect 201862 68824 201868 68836
rect 201920 68824 201926 68876
rect 104158 68756 104164 68808
rect 104216 68796 104222 68808
rect 138566 68796 138572 68808
rect 104216 68768 138572 68796
rect 104216 68756 104222 68768
rect 138566 68756 138572 68768
rect 138624 68756 138630 68808
rect 155862 68756 155868 68808
rect 155920 68796 155926 68808
rect 189442 68796 189448 68808
rect 155920 68768 189448 68796
rect 155920 68756 155926 68768
rect 189442 68756 189448 68768
rect 189500 68756 189506 68808
rect 112162 68688 112168 68740
rect 112220 68728 112226 68740
rect 146478 68728 146484 68740
rect 112220 68700 146484 68728
rect 112220 68688 112226 68700
rect 146478 68688 146484 68700
rect 146536 68688 146542 68740
rect 164050 68688 164056 68740
rect 164108 68728 164114 68740
rect 197538 68728 197544 68740
rect 164108 68700 197544 68728
rect 164108 68688 164114 68700
rect 197538 68688 197544 68700
rect 197596 68688 197602 68740
rect 99190 68620 99196 68672
rect 99248 68660 99254 68672
rect 133138 68660 133144 68672
rect 99248 68632 133144 68660
rect 99248 68620 99254 68632
rect 133138 68620 133144 68632
rect 133196 68620 133202 68672
rect 161842 68620 161848 68672
rect 161900 68660 161906 68672
rect 196250 68660 196256 68672
rect 161900 68632 196256 68660
rect 161900 68620 161906 68632
rect 196250 68620 196256 68632
rect 196308 68620 196314 68672
rect 114278 68552 114284 68604
rect 114336 68592 114342 68604
rect 146846 68592 146852 68604
rect 114336 68564 146852 68592
rect 114336 68552 114342 68564
rect 146846 68552 146852 68564
rect 146904 68552 146910 68604
rect 159174 68552 159180 68604
rect 159232 68592 159238 68604
rect 193306 68592 193312 68604
rect 159232 68564 193312 68592
rect 159232 68552 159238 68564
rect 193306 68552 193312 68564
rect 193364 68552 193370 68604
rect 116210 68484 116216 68536
rect 116268 68524 116274 68536
rect 148594 68524 148600 68536
rect 116268 68496 148600 68524
rect 116268 68484 116274 68496
rect 148594 68484 148600 68496
rect 148652 68484 148658 68536
rect 159266 68484 159272 68536
rect 159324 68524 159330 68536
rect 194226 68524 194232 68536
rect 159324 68496 194232 68524
rect 159324 68484 159330 68496
rect 194226 68484 194232 68496
rect 194284 68484 194290 68536
rect 111518 68416 111524 68468
rect 111576 68456 111582 68468
rect 141418 68456 141424 68468
rect 111576 68428 141424 68456
rect 111576 68416 111582 68428
rect 141418 68416 141424 68428
rect 141476 68416 141482 68468
rect 174630 68416 174636 68468
rect 174688 68456 174694 68468
rect 207474 68456 207480 68468
rect 174688 68428 207480 68456
rect 174688 68416 174694 68428
rect 207474 68416 207480 68428
rect 207532 68416 207538 68468
rect 120718 68348 120724 68400
rect 120776 68388 120782 68400
rect 150066 68388 150072 68400
rect 120776 68360 150072 68388
rect 120776 68348 120782 68360
rect 150066 68348 150072 68360
rect 150124 68348 150130 68400
rect 150434 68348 150440 68400
rect 150492 68388 150498 68400
rect 310514 68388 310520 68400
rect 150492 68360 310520 68388
rect 150492 68348 150498 68360
rect 310514 68348 310520 68360
rect 310572 68348 310578 68400
rect 95878 68280 95884 68332
rect 95936 68320 95942 68332
rect 132494 68320 132500 68332
rect 95936 68292 132500 68320
rect 95936 68280 95942 68292
rect 132494 68280 132500 68292
rect 132552 68320 132558 68332
rect 139854 68320 139860 68332
rect 132552 68292 139860 68320
rect 132552 68280 132558 68292
rect 139854 68280 139860 68292
rect 139912 68280 139918 68332
rect 149238 68280 149244 68332
rect 149296 68320 149302 68332
rect 462314 68320 462320 68332
rect 149296 68292 462320 68320
rect 149296 68280 149302 68292
rect 462314 68280 462320 68292
rect 462372 68280 462378 68332
rect 107010 68212 107016 68264
rect 107068 68252 107074 68264
rect 135530 68252 135536 68264
rect 107068 68224 135536 68252
rect 107068 68212 107074 68224
rect 135530 68212 135536 68224
rect 135588 68212 135594 68264
rect 162670 68212 162676 68264
rect 162728 68252 162734 68264
rect 181438 68252 181444 68264
rect 162728 68224 181444 68252
rect 162728 68212 162734 68224
rect 181438 68212 181444 68224
rect 181496 68212 181502 68264
rect 182174 68212 182180 68264
rect 182232 68252 182238 68264
rect 211154 68252 211160 68264
rect 182232 68224 211160 68252
rect 182232 68212 182238 68224
rect 211154 68212 211160 68224
rect 211212 68212 211218 68264
rect 3510 68144 3516 68196
rect 3568 68184 3574 68196
rect 153102 68184 153108 68196
rect 3568 68156 153108 68184
rect 3568 68144 3574 68156
rect 153102 68144 153108 68156
rect 153160 68144 153166 68196
rect 163314 68144 163320 68196
rect 163372 68184 163378 68196
rect 208762 68184 208768 68196
rect 163372 68156 208768 68184
rect 163372 68144 163378 68156
rect 208762 68144 208768 68156
rect 208820 68144 208826 68196
rect 105354 68076 105360 68128
rect 105412 68116 105418 68128
rect 155034 68116 155040 68128
rect 105412 68088 155040 68116
rect 105412 68076 105418 68088
rect 155034 68076 155040 68088
rect 155092 68116 155098 68128
rect 155862 68116 155868 68128
rect 155092 68088 155868 68116
rect 155092 68076 155098 68088
rect 155862 68076 155868 68088
rect 155920 68076 155926 68128
rect 156230 68008 156236 68060
rect 156288 68048 156294 68060
rect 156690 68048 156696 68060
rect 156288 68020 156696 68048
rect 156288 68008 156294 68020
rect 156690 68008 156696 68020
rect 156748 68008 156754 68060
rect 109678 67532 109684 67584
rect 109736 67572 109742 67584
rect 144362 67572 144368 67584
rect 109736 67544 144368 67572
rect 109736 67532 109742 67544
rect 144362 67532 144368 67544
rect 144420 67532 144426 67584
rect 145466 67532 145472 67584
rect 145524 67572 145530 67584
rect 145650 67572 145656 67584
rect 145524 67544 145656 67572
rect 145524 67532 145530 67544
rect 145650 67532 145656 67544
rect 145708 67532 145714 67584
rect 164510 67532 164516 67584
rect 164568 67572 164574 67584
rect 165430 67572 165436 67584
rect 164568 67544 165436 67572
rect 164568 67532 164574 67544
rect 165430 67532 165436 67544
rect 165488 67532 165494 67584
rect 165982 67532 165988 67584
rect 166040 67572 166046 67584
rect 166810 67572 166816 67584
rect 166040 67544 166816 67572
rect 166040 67532 166046 67544
rect 166810 67532 166816 67544
rect 166868 67532 166874 67584
rect 167730 67532 167736 67584
rect 167788 67572 167794 67584
rect 192846 67572 192852 67584
rect 167788 67544 192852 67572
rect 167788 67532 167794 67544
rect 192846 67532 192852 67544
rect 192904 67532 192910 67584
rect 104434 67464 104440 67516
rect 104492 67504 104498 67516
rect 136634 67504 136640 67516
rect 104492 67476 136640 67504
rect 104492 67464 104498 67476
rect 136634 67464 136640 67476
rect 136692 67464 136698 67516
rect 136818 67464 136824 67516
rect 136876 67504 136882 67516
rect 137278 67504 137284 67516
rect 136876 67476 137284 67504
rect 136876 67464 136882 67476
rect 137278 67464 137284 67476
rect 137336 67464 137342 67516
rect 138750 67464 138756 67516
rect 138808 67504 138814 67516
rect 138934 67504 138940 67516
rect 138808 67476 138940 67504
rect 138808 67464 138814 67476
rect 138934 67464 138940 67476
rect 138992 67464 138998 67516
rect 157518 67464 157524 67516
rect 157576 67504 157582 67516
rect 207198 67504 207204 67516
rect 157576 67476 207204 67504
rect 157576 67464 157582 67476
rect 207198 67464 207204 67476
rect 207256 67464 207262 67516
rect 109954 67396 109960 67448
rect 110012 67436 110018 67448
rect 143626 67436 143632 67448
rect 110012 67408 143632 67436
rect 110012 67396 110018 67408
rect 143626 67396 143632 67408
rect 143684 67436 143690 67448
rect 144270 67436 144276 67448
rect 143684 67408 144276 67436
rect 143684 67396 143690 67408
rect 144270 67396 144276 67408
rect 144328 67396 144334 67448
rect 165890 67396 165896 67448
rect 165948 67436 165954 67448
rect 166902 67436 166908 67448
rect 165948 67408 166908 67436
rect 165948 67396 165954 67408
rect 166902 67396 166908 67408
rect 166960 67396 166966 67448
rect 169938 67396 169944 67448
rect 169996 67436 170002 67448
rect 211982 67436 211988 67448
rect 169996 67408 211988 67436
rect 169996 67396 170002 67408
rect 211982 67396 211988 67408
rect 212040 67396 212046 67448
rect 110874 67328 110880 67380
rect 110932 67368 110938 67380
rect 145650 67368 145656 67380
rect 110932 67340 145656 67368
rect 110932 67328 110938 67340
rect 145650 67328 145656 67340
rect 145708 67328 145714 67380
rect 153470 67328 153476 67380
rect 153528 67368 153534 67380
rect 188798 67368 188804 67380
rect 153528 67340 188804 67368
rect 153528 67328 153534 67340
rect 188798 67328 188804 67340
rect 188856 67328 188862 67380
rect 104342 67260 104348 67312
rect 104400 67300 104406 67312
rect 136818 67300 136824 67312
rect 104400 67272 136824 67300
rect 104400 67260 104406 67272
rect 136818 67260 136824 67272
rect 136876 67260 136882 67312
rect 161842 67260 161848 67312
rect 161900 67300 161906 67312
rect 165614 67300 165620 67312
rect 161900 67272 165620 67300
rect 161900 67260 161906 67272
rect 165614 67260 165620 67272
rect 165672 67300 165678 67312
rect 200758 67300 200764 67312
rect 165672 67272 200764 67300
rect 165672 67260 165678 67272
rect 200758 67260 200764 67272
rect 200816 67260 200822 67312
rect 104710 67192 104716 67244
rect 104768 67232 104774 67244
rect 136910 67232 136916 67244
rect 104768 67204 136916 67232
rect 104768 67192 104774 67204
rect 136910 67192 136916 67204
rect 136968 67192 136974 67244
rect 168834 67192 168840 67244
rect 168892 67232 168898 67244
rect 169202 67232 169208 67244
rect 168892 67204 169208 67232
rect 168892 67192 168898 67204
rect 169202 67192 169208 67204
rect 169260 67232 169266 67244
rect 203702 67232 203708 67244
rect 169260 67204 203708 67232
rect 169260 67192 169266 67204
rect 203702 67192 203708 67204
rect 203760 67192 203766 67244
rect 104618 67124 104624 67176
rect 104676 67164 104682 67176
rect 136726 67164 136732 67176
rect 104676 67136 136732 67164
rect 104676 67124 104682 67136
rect 136726 67124 136732 67136
rect 136784 67124 136790 67176
rect 166902 67124 166908 67176
rect 166960 67164 166966 67176
rect 200666 67164 200672 67176
rect 166960 67136 200672 67164
rect 166960 67124 166966 67136
rect 200666 67124 200672 67136
rect 200724 67124 200730 67176
rect 103238 67056 103244 67108
rect 103296 67096 103302 67108
rect 134886 67096 134892 67108
rect 103296 67068 134892 67096
rect 103296 67056 103302 67068
rect 134886 67056 134892 67068
rect 134944 67056 134950 67108
rect 136634 67056 136640 67108
rect 136692 67096 136698 67108
rect 138750 67096 138756 67108
rect 136692 67068 138756 67096
rect 136692 67056 136698 67068
rect 138750 67056 138756 67068
rect 138808 67056 138814 67108
rect 165430 67056 165436 67108
rect 165488 67096 165494 67108
rect 199654 67096 199660 67108
rect 165488 67068 199660 67096
rect 165488 67056 165494 67068
rect 199654 67056 199660 67068
rect 199712 67056 199718 67108
rect 93854 66988 93860 67040
rect 93912 67028 93918 67040
rect 166166 67028 166172 67040
rect 93912 67000 166172 67028
rect 93912 66988 93918 67000
rect 166166 66988 166172 67000
rect 166224 66988 166230 67040
rect 175366 66988 175372 67040
rect 175424 67028 175430 67040
rect 210050 67028 210056 67040
rect 175424 67000 210056 67028
rect 175424 66988 175430 67000
rect 210050 66988 210056 67000
rect 210108 66988 210114 67040
rect 121546 66920 121552 66972
rect 121604 66960 121610 66972
rect 148134 66960 148140 66972
rect 121604 66932 148140 66960
rect 121604 66920 121610 66932
rect 148134 66920 148140 66932
rect 148192 66920 148198 66972
rect 161750 66920 161756 66972
rect 161808 66960 161814 66972
rect 196342 66960 196348 66972
rect 161808 66932 196348 66960
rect 161808 66920 161814 66932
rect 196342 66920 196348 66932
rect 196400 66960 196406 66972
rect 386414 66960 386420 66972
rect 196400 66932 386420 66960
rect 196400 66920 196406 66932
rect 386414 66920 386420 66932
rect 386472 66920 386478 66972
rect 26234 66852 26240 66904
rect 26292 66892 26298 66904
rect 104250 66892 104256 66904
rect 26292 66864 104256 66892
rect 26292 66852 26298 66864
rect 104250 66852 104256 66864
rect 104308 66892 104314 66904
rect 104710 66892 104716 66904
rect 104308 66864 104716 66892
rect 104308 66852 104314 66864
rect 104710 66852 104716 66864
rect 104768 66852 104774 66904
rect 129734 66852 129740 66904
rect 129792 66892 129798 66904
rect 130378 66892 130384 66904
rect 129792 66864 130384 66892
rect 129792 66852 129798 66864
rect 130378 66852 130384 66864
rect 130436 66852 130442 66904
rect 145926 66852 145932 66904
rect 145984 66892 145990 66904
rect 488534 66892 488540 66904
rect 145984 66864 488540 66892
rect 145984 66852 145990 66864
rect 488534 66852 488540 66864
rect 488592 66852 488598 66904
rect 120626 66784 120632 66836
rect 120684 66824 120690 66836
rect 148226 66824 148232 66836
rect 120684 66796 148232 66824
rect 120684 66784 120690 66796
rect 148226 66784 148232 66796
rect 148284 66784 148290 66836
rect 166810 66784 166816 66836
rect 166868 66824 166874 66836
rect 200574 66824 200580 66836
rect 166868 66796 200580 66824
rect 166868 66784 166874 66796
rect 200574 66784 200580 66796
rect 200632 66784 200638 66836
rect 121638 66716 121644 66768
rect 121696 66756 121702 66768
rect 149606 66756 149612 66768
rect 121696 66728 149612 66756
rect 121696 66716 121702 66728
rect 149606 66716 149612 66728
rect 149664 66716 149670 66768
rect 156138 66716 156144 66768
rect 156196 66756 156202 66768
rect 216030 66756 216036 66768
rect 156196 66728 216036 66756
rect 156196 66716 156202 66728
rect 216030 66716 216036 66728
rect 216088 66716 216094 66768
rect 110046 66648 110052 66700
rect 110104 66688 110110 66700
rect 129734 66688 129740 66700
rect 110104 66660 129740 66688
rect 110104 66648 110110 66660
rect 129734 66648 129740 66660
rect 129792 66648 129798 66700
rect 89714 66580 89720 66632
rect 89772 66620 89778 66632
rect 168834 66620 168840 66632
rect 89772 66592 168840 66620
rect 89772 66580 89778 66592
rect 168834 66580 168840 66592
rect 168892 66580 168898 66632
rect 121178 66172 121184 66224
rect 121236 66212 121242 66224
rect 135990 66212 135996 66224
rect 121236 66184 135996 66212
rect 121236 66172 121242 66184
rect 135990 66172 135996 66184
rect 136048 66172 136054 66224
rect 158990 66172 158996 66224
rect 159048 66212 159054 66224
rect 220998 66212 221004 66224
rect 159048 66184 221004 66212
rect 159048 66172 159054 66184
rect 220998 66172 221004 66184
rect 221056 66172 221062 66224
rect 120534 66104 120540 66156
rect 120592 66144 120598 66156
rect 141050 66144 141056 66156
rect 120592 66116 141056 66144
rect 120592 66104 120598 66116
rect 141050 66104 141056 66116
rect 141108 66104 141114 66156
rect 157334 66104 157340 66156
rect 157392 66144 157398 66156
rect 211338 66144 211344 66156
rect 157392 66116 211344 66144
rect 157392 66104 157398 66116
rect 211338 66104 211344 66116
rect 211396 66104 211402 66156
rect 100386 66036 100392 66088
rect 100444 66076 100450 66088
rect 134334 66076 134340 66088
rect 100444 66048 134340 66076
rect 100444 66036 100450 66048
rect 134334 66036 134340 66048
rect 134392 66036 134398 66088
rect 154850 66036 154856 66088
rect 154908 66076 154914 66088
rect 189258 66076 189264 66088
rect 154908 66048 189264 66076
rect 154908 66036 154914 66048
rect 189258 66036 189264 66048
rect 189316 66036 189322 66088
rect 98914 65968 98920 66020
rect 98972 66008 98978 66020
rect 133138 66008 133144 66020
rect 98972 65980 133144 66008
rect 98972 65968 98978 65980
rect 133138 65968 133144 65980
rect 133196 66008 133202 66020
rect 133414 66008 133420 66020
rect 133196 65980 133420 66008
rect 133196 65968 133202 65980
rect 133414 65968 133420 65980
rect 133472 65968 133478 66020
rect 156874 65968 156880 66020
rect 156932 66008 156938 66020
rect 191006 66008 191012 66020
rect 156932 65980 191012 66008
rect 156932 65968 156938 65980
rect 191006 65968 191012 65980
rect 191064 65968 191070 66020
rect 104066 65900 104072 65952
rect 104124 65940 104130 65952
rect 138474 65940 138480 65952
rect 104124 65912 138480 65940
rect 104124 65900 104130 65912
rect 138474 65900 138480 65912
rect 138532 65900 138538 65952
rect 169754 65900 169760 65952
rect 169812 65940 169818 65952
rect 171042 65940 171048 65952
rect 169812 65912 171048 65940
rect 169812 65900 169818 65912
rect 171042 65900 171048 65912
rect 171100 65940 171106 65952
rect 204714 65940 204720 65952
rect 171100 65912 204720 65940
rect 171100 65900 171106 65912
rect 204714 65900 204720 65912
rect 204772 65900 204778 65952
rect 105446 65832 105452 65884
rect 105504 65872 105510 65884
rect 140314 65872 140320 65884
rect 105504 65844 140320 65872
rect 105504 65832 105510 65844
rect 140314 65832 140320 65844
rect 140372 65832 140378 65884
rect 171318 65832 171324 65884
rect 171376 65872 171382 65884
rect 172330 65872 172336 65884
rect 171376 65844 172336 65872
rect 171376 65832 171382 65844
rect 172330 65832 172336 65844
rect 172388 65832 172394 65884
rect 174078 65832 174084 65884
rect 174136 65872 174142 65884
rect 175090 65872 175096 65884
rect 174136 65844 175096 65872
rect 174136 65832 174142 65844
rect 175090 65832 175096 65844
rect 175148 65832 175154 65884
rect 175274 65832 175280 65884
rect 175332 65872 175338 65884
rect 176562 65872 176568 65884
rect 175332 65844 176568 65872
rect 175332 65832 175338 65844
rect 176562 65832 176568 65844
rect 176620 65832 176626 65884
rect 176654 65832 176660 65884
rect 176712 65872 176718 65884
rect 205910 65872 205916 65884
rect 176712 65844 205916 65872
rect 176712 65832 176718 65844
rect 205910 65832 205916 65844
rect 205968 65832 205974 65884
rect 100570 65764 100576 65816
rect 100628 65804 100634 65816
rect 134150 65804 134156 65816
rect 100628 65776 134156 65804
rect 100628 65764 100634 65776
rect 134150 65764 134156 65776
rect 134208 65804 134214 65816
rect 135898 65804 135904 65816
rect 134208 65776 135904 65804
rect 134208 65764 134214 65776
rect 135898 65764 135904 65776
rect 135956 65764 135962 65816
rect 172348 65804 172376 65832
rect 206002 65804 206008 65816
rect 172348 65776 206008 65804
rect 206002 65764 206008 65776
rect 206060 65764 206066 65816
rect 107562 65696 107568 65748
rect 107620 65736 107626 65748
rect 141142 65736 141148 65748
rect 107620 65708 141148 65736
rect 107620 65696 107626 65708
rect 141142 65696 141148 65708
rect 141200 65696 141206 65748
rect 160094 65696 160100 65748
rect 160152 65736 160158 65748
rect 195514 65736 195520 65748
rect 160152 65708 195520 65736
rect 160152 65696 160158 65708
rect 195514 65696 195520 65708
rect 195572 65696 195578 65748
rect 167270 65628 167276 65680
rect 167328 65668 167334 65680
rect 201770 65668 201776 65680
rect 167328 65640 201776 65668
rect 167328 65628 167334 65640
rect 201770 65628 201776 65640
rect 201828 65628 201834 65680
rect 102594 65560 102600 65612
rect 102652 65600 102658 65612
rect 135438 65600 135444 65612
rect 102652 65572 135444 65600
rect 102652 65560 102658 65572
rect 135438 65560 135444 65572
rect 135496 65560 135502 65612
rect 147214 65560 147220 65612
rect 147272 65600 147278 65612
rect 260834 65600 260840 65612
rect 147272 65572 260840 65600
rect 147272 65560 147278 65572
rect 260834 65560 260840 65572
rect 260892 65560 260898 65612
rect 67634 65492 67640 65544
rect 67692 65532 67698 65544
rect 110138 65532 110144 65544
rect 67692 65504 110144 65532
rect 67692 65492 67698 65504
rect 110138 65492 110144 65504
rect 110196 65532 110202 65544
rect 142706 65532 142712 65544
rect 110196 65504 142712 65532
rect 110196 65492 110202 65504
rect 142706 65492 142712 65504
rect 142764 65492 142770 65544
rect 146018 65492 146024 65544
rect 146076 65532 146082 65544
rect 408494 65532 408500 65544
rect 146076 65504 408500 65532
rect 146076 65492 146082 65504
rect 408494 65492 408500 65504
rect 408552 65492 408558 65544
rect 111426 65424 111432 65476
rect 111484 65464 111490 65476
rect 140866 65464 140872 65476
rect 111484 65436 140872 65464
rect 111484 65424 111490 65436
rect 140866 65424 140872 65436
rect 140924 65464 140930 65476
rect 141510 65464 141516 65476
rect 140924 65436 141516 65464
rect 140924 65424 140930 65436
rect 141510 65424 141516 65436
rect 141568 65424 141574 65476
rect 171226 65424 171232 65476
rect 171284 65464 171290 65476
rect 172422 65464 172428 65476
rect 171284 65436 172428 65464
rect 171284 65424 171290 65436
rect 172422 65424 172428 65436
rect 172480 65424 172486 65476
rect 175090 65424 175096 65476
rect 175148 65464 175154 65476
rect 208578 65464 208584 65476
rect 175148 65436 208584 65464
rect 175148 65424 175154 65436
rect 208578 65424 208584 65436
rect 208636 65424 208642 65476
rect 101398 65356 101404 65408
rect 101456 65396 101462 65408
rect 140590 65396 140596 65408
rect 101456 65368 140596 65396
rect 101456 65356 101462 65368
rect 140590 65356 140596 65368
rect 140648 65356 140654 65408
rect 158346 65356 158352 65408
rect 158404 65396 158410 65408
rect 188614 65396 188620 65408
rect 158404 65368 188620 65396
rect 158404 65356 158410 65368
rect 188614 65356 188620 65368
rect 188672 65356 188678 65408
rect 100018 65288 100024 65340
rect 100076 65328 100082 65340
rect 134702 65328 134708 65340
rect 100076 65300 134708 65328
rect 100076 65288 100082 65300
rect 134702 65288 134708 65300
rect 134760 65288 134766 65340
rect 176562 65288 176568 65340
rect 176620 65328 176626 65340
rect 210326 65328 210332 65340
rect 176620 65300 210332 65328
rect 176620 65288 176626 65300
rect 210326 65288 210332 65300
rect 210384 65288 210390 65340
rect 100478 65220 100484 65272
rect 100536 65260 100542 65272
rect 134978 65260 134984 65272
rect 100536 65232 134984 65260
rect 100536 65220 100542 65232
rect 134978 65220 134984 65232
rect 135036 65220 135042 65272
rect 172422 65220 172428 65272
rect 172480 65260 172486 65272
rect 176654 65260 176660 65272
rect 172480 65232 176660 65260
rect 172480 65220 172486 65232
rect 176654 65220 176660 65232
rect 176712 65220 176718 65272
rect 106090 64812 106096 64864
rect 106148 64852 106154 64864
rect 135622 64852 135628 64864
rect 106148 64824 135628 64852
rect 106148 64812 106154 64824
rect 135622 64812 135628 64824
rect 135680 64812 135686 64864
rect 138290 64812 138296 64864
rect 138348 64852 138354 64864
rect 580718 64852 580724 64864
rect 138348 64824 580724 64852
rect 138348 64812 138354 64824
rect 580718 64812 580724 64824
rect 580776 64812 580782 64864
rect 112898 64744 112904 64796
rect 112956 64784 112962 64796
rect 141326 64784 141332 64796
rect 112956 64756 141332 64784
rect 112956 64744 112962 64756
rect 141326 64744 141332 64756
rect 141384 64744 141390 64796
rect 154758 64744 154764 64796
rect 154816 64784 154822 64796
rect 215938 64784 215944 64796
rect 154816 64756 215944 64784
rect 154816 64744 154822 64756
rect 215938 64744 215944 64756
rect 215996 64744 216002 64796
rect 96338 64676 96344 64728
rect 96396 64716 96402 64728
rect 136082 64716 136088 64728
rect 96396 64688 136088 64716
rect 96396 64676 96402 64688
rect 136082 64676 136088 64688
rect 136140 64676 136146 64728
rect 168742 64676 168748 64728
rect 168800 64716 168806 64728
rect 212534 64716 212540 64728
rect 168800 64688 212540 64716
rect 168800 64676 168806 64688
rect 212534 64676 212540 64688
rect 212592 64676 212598 64728
rect 99098 64608 99104 64660
rect 99156 64648 99162 64660
rect 133230 64648 133236 64660
rect 99156 64620 133236 64648
rect 99156 64608 99162 64620
rect 133230 64608 133236 64620
rect 133288 64608 133294 64660
rect 175182 64608 175188 64660
rect 175240 64648 175246 64660
rect 213914 64648 213920 64660
rect 175240 64620 213920 64648
rect 175240 64608 175246 64620
rect 213914 64608 213920 64620
rect 213972 64608 213978 64660
rect 100662 64540 100668 64592
rect 100720 64580 100726 64592
rect 134610 64580 134616 64592
rect 100720 64552 134616 64580
rect 100720 64540 100726 64552
rect 134610 64540 134616 64552
rect 134668 64540 134674 64592
rect 158898 64540 158904 64592
rect 158956 64580 158962 64592
rect 188338 64580 188344 64592
rect 158956 64552 188344 64580
rect 158956 64540 158962 64552
rect 188338 64540 188344 64552
rect 188396 64540 188402 64592
rect 99926 64472 99932 64524
rect 99984 64512 99990 64524
rect 134426 64512 134432 64524
rect 99984 64484 134432 64512
rect 99984 64472 99990 64484
rect 134426 64472 134432 64484
rect 134484 64472 134490 64524
rect 165062 64472 165068 64524
rect 165120 64512 165126 64524
rect 191374 64512 191380 64524
rect 165120 64484 191380 64512
rect 165120 64472 165126 64484
rect 191374 64472 191380 64484
rect 191432 64472 191438 64524
rect 108390 64404 108396 64456
rect 108448 64444 108454 64456
rect 141418 64444 141424 64456
rect 108448 64416 141424 64444
rect 108448 64404 108454 64416
rect 141418 64404 141424 64416
rect 141476 64444 141482 64456
rect 142062 64444 142068 64456
rect 141476 64416 142068 64444
rect 141476 64404 141482 64416
rect 142062 64404 142068 64416
rect 142120 64404 142126 64456
rect 163038 64404 163044 64456
rect 163096 64444 163102 64456
rect 188890 64444 188896 64456
rect 163096 64416 188896 64444
rect 163096 64404 163102 64416
rect 188890 64404 188896 64416
rect 188948 64404 188954 64456
rect 107286 64336 107292 64388
rect 107344 64376 107350 64388
rect 139762 64376 139768 64388
rect 107344 64348 139768 64376
rect 107344 64336 107350 64348
rect 139762 64336 139768 64348
rect 139820 64336 139826 64388
rect 107378 64268 107384 64320
rect 107436 64308 107442 64320
rect 139670 64308 139676 64320
rect 107436 64280 139676 64308
rect 107436 64268 107442 64280
rect 139670 64268 139676 64280
rect 139728 64268 139734 64320
rect 148226 64268 148232 64320
rect 148284 64308 148290 64320
rect 184934 64308 184940 64320
rect 148284 64280 184940 64308
rect 148284 64268 148290 64280
rect 184934 64268 184940 64280
rect 184992 64268 184998 64320
rect 102778 64200 102784 64252
rect 102836 64240 102842 64252
rect 132954 64240 132960 64252
rect 102836 64212 132960 64240
rect 102836 64200 102842 64212
rect 132954 64200 132960 64212
rect 133012 64200 133018 64252
rect 133322 64200 133328 64252
rect 133380 64240 133386 64252
rect 264974 64240 264980 64252
rect 133380 64212 264980 64240
rect 133380 64200 133386 64212
rect 264974 64200 264980 64212
rect 265032 64200 265038 64252
rect 63494 64132 63500 64184
rect 63552 64172 63558 64184
rect 106090 64172 106096 64184
rect 63552 64144 106096 64172
rect 63552 64132 63558 64144
rect 106090 64132 106096 64144
rect 106148 64132 106154 64184
rect 108574 64132 108580 64184
rect 108632 64172 108638 64184
rect 139578 64172 139584 64184
rect 108632 64144 139584 64172
rect 108632 64132 108638 64144
rect 139578 64132 139584 64144
rect 139636 64132 139642 64184
rect 142890 64132 142896 64184
rect 142948 64172 142954 64184
rect 477494 64172 477500 64184
rect 142948 64144 477500 64172
rect 142948 64132 142954 64144
rect 477494 64132 477500 64144
rect 477552 64132 477558 64184
rect 97258 64064 97264 64116
rect 97316 64104 97322 64116
rect 138658 64104 138664 64116
rect 97316 64076 138664 64104
rect 97316 64064 97322 64076
rect 138658 64064 138664 64076
rect 138716 64064 138722 64116
rect 97350 63996 97356 64048
rect 97408 64036 97414 64048
rect 137094 64036 137100 64048
rect 97408 64008 137100 64036
rect 97408 63996 97414 64008
rect 137094 63996 137100 64008
rect 137152 63996 137158 64048
rect 133874 63860 133880 63912
rect 133932 63900 133938 63912
rect 134426 63900 134432 63912
rect 133932 63872 134432 63900
rect 133932 63860 133938 63872
rect 134426 63860 134432 63872
rect 134484 63860 134490 63912
rect 139670 63588 139676 63640
rect 139728 63628 139734 63640
rect 140130 63628 140136 63640
rect 139728 63600 140136 63628
rect 139728 63588 139734 63600
rect 140130 63588 140136 63600
rect 140188 63588 140194 63640
rect 173986 63588 173992 63640
rect 174044 63628 174050 63640
rect 175182 63628 175188 63640
rect 174044 63600 175188 63628
rect 174044 63588 174050 63600
rect 175182 63588 175188 63600
rect 175240 63588 175246 63640
rect 102134 63520 102140 63572
rect 102192 63560 102198 63572
rect 102778 63560 102784 63572
rect 102192 63532 102784 63560
rect 102192 63520 102198 63532
rect 102778 63520 102784 63532
rect 102836 63520 102842 63572
rect 137094 63520 137100 63572
rect 137152 63560 137158 63572
rect 137370 63560 137376 63572
rect 137152 63532 137376 63560
rect 137152 63520 137158 63532
rect 137370 63520 137376 63532
rect 137428 63520 137434 63572
rect 139762 63520 139768 63572
rect 139820 63560 139826 63572
rect 140038 63560 140044 63572
rect 139820 63532 140044 63560
rect 139820 63520 139826 63532
rect 140038 63520 140044 63532
rect 140096 63520 140102 63572
rect 97810 63452 97816 63504
rect 97868 63492 97874 63504
rect 158806 63492 158812 63504
rect 97868 63464 158812 63492
rect 97868 63452 97874 63464
rect 158806 63452 158812 63464
rect 158864 63452 158870 63504
rect 162762 63452 162768 63504
rect 162820 63492 162826 63504
rect 211522 63492 211528 63504
rect 162820 63464 211528 63492
rect 162820 63452 162826 63464
rect 211522 63452 211528 63464
rect 211580 63452 211586 63504
rect 96430 63384 96436 63436
rect 96488 63424 96494 63436
rect 150802 63424 150808 63436
rect 96488 63396 150808 63424
rect 96488 63384 96494 63396
rect 150802 63384 150808 63396
rect 150860 63384 150866 63436
rect 168650 63384 168656 63436
rect 168708 63424 168714 63436
rect 212626 63424 212632 63436
rect 168708 63396 212632 63424
rect 168708 63384 168714 63396
rect 212626 63384 212632 63396
rect 212684 63384 212690 63436
rect 101950 63316 101956 63368
rect 102008 63356 102014 63368
rect 142522 63356 142528 63368
rect 102008 63328 142528 63356
rect 102008 63316 102014 63328
rect 142522 63316 142528 63328
rect 142580 63356 142586 63368
rect 143442 63356 143448 63368
rect 142580 63328 143448 63356
rect 142580 63316 142586 63328
rect 143442 63316 143448 63328
rect 143500 63316 143506 63368
rect 162854 63316 162860 63368
rect 162912 63356 162918 63368
rect 204254 63356 204260 63368
rect 162912 63328 204260 63356
rect 162912 63316 162918 63328
rect 204254 63316 204260 63328
rect 204312 63316 204318 63368
rect 115014 63248 115020 63300
rect 115072 63288 115078 63300
rect 153378 63288 153384 63300
rect 115072 63260 153384 63288
rect 115072 63248 115078 63260
rect 153378 63248 153384 63260
rect 153436 63248 153442 63300
rect 165522 63248 165528 63300
rect 165580 63288 165586 63300
rect 206554 63288 206560 63300
rect 165580 63260 206560 63288
rect 165580 63248 165586 63260
rect 206554 63248 206560 63260
rect 206612 63248 206618 63300
rect 119614 63180 119620 63232
rect 119672 63220 119678 63232
rect 151906 63220 151912 63232
rect 119672 63192 151912 63220
rect 119672 63180 119678 63192
rect 151906 63180 151912 63192
rect 151964 63220 151970 63232
rect 152550 63220 152556 63232
rect 151964 63192 152556 63220
rect 151964 63180 151970 63192
rect 152550 63180 152556 63192
rect 152608 63180 152614 63232
rect 169570 63180 169576 63232
rect 169628 63220 169634 63232
rect 209774 63220 209780 63232
rect 169628 63192 209780 63220
rect 169628 63180 169634 63192
rect 209774 63180 209780 63192
rect 209832 63180 209838 63232
rect 109586 63112 109592 63164
rect 109644 63152 109650 63164
rect 131114 63152 131120 63164
rect 109644 63124 131120 63152
rect 109644 63112 109650 63124
rect 131114 63112 131120 63124
rect 131172 63112 131178 63164
rect 164326 63112 164332 63164
rect 164384 63152 164390 63164
rect 199562 63152 199568 63164
rect 164384 63124 199568 63152
rect 164384 63112 164390 63124
rect 199562 63112 199568 63124
rect 199620 63112 199626 63164
rect 168282 63044 168288 63096
rect 168340 63084 168346 63096
rect 202046 63084 202052 63096
rect 168340 63056 202052 63084
rect 168340 63044 168346 63056
rect 202046 63044 202052 63056
rect 202104 63044 202110 63096
rect 165614 62976 165620 63028
rect 165672 63016 165678 63028
rect 213178 63016 213184 63028
rect 165672 62988 213184 63016
rect 165672 62976 165678 62988
rect 213178 62976 213184 62988
rect 213236 62976 213242 63028
rect 146294 62908 146300 62960
rect 146352 62948 146358 62960
rect 213086 62948 213092 62960
rect 146352 62920 213092 62948
rect 146352 62908 146358 62920
rect 213086 62908 213092 62920
rect 213144 62908 213150 62960
rect 148502 62840 148508 62892
rect 148560 62880 148566 62892
rect 302234 62880 302240 62892
rect 148560 62852 302240 62880
rect 148560 62840 148566 62852
rect 302234 62840 302240 62852
rect 302292 62840 302298 62892
rect 8938 62772 8944 62824
rect 8996 62812 9002 62824
rect 97810 62812 97816 62824
rect 8996 62784 97816 62812
rect 8996 62772 9002 62784
rect 97810 62772 97816 62784
rect 97868 62772 97874 62824
rect 168558 62772 168564 62824
rect 168616 62812 168622 62824
rect 203426 62812 203432 62824
rect 168616 62784 203432 62812
rect 168616 62772 168622 62784
rect 203426 62772 203432 62784
rect 203484 62812 203490 62824
rect 425054 62812 425060 62824
rect 203484 62784 425060 62812
rect 203484 62772 203490 62784
rect 425054 62772 425060 62784
rect 425112 62772 425118 62824
rect 162946 62704 162952 62756
rect 163004 62744 163010 62756
rect 197446 62744 197452 62756
rect 163004 62716 197452 62744
rect 163004 62704 163010 62716
rect 197446 62704 197452 62716
rect 197504 62704 197510 62756
rect 170674 62636 170680 62688
rect 170732 62676 170738 62688
rect 203518 62676 203524 62688
rect 170732 62648 203524 62676
rect 170732 62636 170738 62648
rect 203518 62636 203524 62648
rect 203576 62636 203582 62688
rect 166718 62568 166724 62620
rect 166776 62608 166782 62620
rect 194042 62608 194048 62620
rect 166776 62580 194048 62608
rect 166776 62568 166782 62580
rect 194042 62568 194048 62580
rect 194100 62568 194106 62620
rect 164418 62500 164424 62552
rect 164476 62540 164482 62552
rect 165522 62540 165528 62552
rect 164476 62512 165528 62540
rect 164476 62500 164482 62512
rect 165522 62500 165528 62512
rect 165580 62500 165586 62552
rect 131114 62432 131120 62484
rect 131172 62472 131178 62484
rect 131850 62472 131856 62484
rect 131172 62444 131856 62472
rect 131172 62432 131178 62444
rect 131850 62432 131856 62444
rect 131908 62432 131914 62484
rect 165798 62364 165804 62416
rect 165856 62404 165862 62416
rect 166718 62404 166724 62416
rect 165856 62376 166724 62404
rect 165856 62364 165862 62376
rect 166718 62364 166724 62376
rect 166776 62364 166782 62416
rect 153378 62092 153384 62144
rect 153436 62132 153442 62144
rect 153838 62132 153844 62144
rect 153436 62104 153844 62132
rect 153436 62092 153442 62104
rect 153838 62092 153844 62104
rect 153896 62092 153902 62144
rect 96062 62024 96068 62076
rect 96120 62064 96126 62076
rect 96246 62064 96252 62076
rect 96120 62036 96252 62064
rect 96120 62024 96126 62036
rect 96246 62024 96252 62036
rect 96304 62064 96310 62076
rect 161566 62064 161572 62076
rect 96304 62036 161572 62064
rect 96304 62024 96310 62036
rect 161566 62024 161572 62036
rect 161624 62024 161630 62076
rect 168466 62024 168472 62076
rect 168524 62064 168530 62076
rect 203334 62064 203340 62076
rect 168524 62036 203340 62064
rect 168524 62024 168530 62036
rect 203334 62024 203340 62036
rect 203392 62024 203398 62076
rect 149790 61412 149796 61464
rect 149848 61452 149854 61464
rect 295334 61452 295340 61464
rect 149848 61424 295340 61452
rect 149848 61412 149854 61424
rect 295334 61412 295340 61424
rect 295392 61412 295398 61464
rect 6914 61344 6920 61396
rect 6972 61384 6978 61396
rect 96062 61384 96068 61396
rect 6972 61356 96068 61384
rect 6972 61344 6978 61356
rect 96062 61344 96068 61356
rect 96120 61344 96126 61396
rect 203334 61344 203340 61396
rect 203392 61384 203398 61396
rect 496078 61384 496084 61396
rect 203392 61356 496084 61384
rect 203392 61344 203398 61356
rect 496078 61344 496084 61356
rect 496136 61344 496142 61396
rect 3510 60664 3516 60716
rect 3568 60704 3574 60716
rect 161842 60704 161848 60716
rect 3568 60676 161848 60704
rect 3568 60664 3574 60676
rect 161842 60664 161848 60676
rect 161900 60664 161906 60716
rect 174446 60664 174452 60716
rect 174504 60704 174510 60716
rect 198734 60704 198740 60716
rect 174504 60676 198740 60704
rect 174504 60664 174510 60676
rect 198734 60664 198740 60676
rect 198792 60704 198798 60716
rect 199010 60704 199016 60716
rect 198792 60676 199016 60704
rect 198792 60664 198798 60676
rect 199010 60664 199016 60676
rect 199068 60664 199074 60716
rect 156782 60596 156788 60648
rect 156840 60636 156846 60648
rect 190638 60636 190644 60648
rect 156840 60608 190644 60636
rect 156840 60596 156846 60608
rect 190638 60596 190644 60608
rect 190696 60636 190702 60648
rect 192478 60636 192484 60648
rect 190696 60608 192484 60636
rect 190696 60596 190702 60608
rect 192478 60596 192484 60608
rect 192536 60596 192542 60648
rect 134242 59984 134248 60036
rect 134300 60024 134306 60036
rect 454034 60024 454040 60036
rect 134300 59996 454040 60024
rect 134300 59984 134306 59996
rect 454034 59984 454040 59996
rect 454092 59984 454098 60036
rect 198734 59848 198740 59900
rect 198792 59888 198798 59900
rect 200114 59888 200120 59900
rect 198792 59860 200120 59888
rect 198792 59848 198798 59860
rect 200114 59848 200120 59860
rect 200172 59848 200178 59900
rect 134886 58760 134892 58812
rect 134944 58800 134950 58812
rect 215294 58800 215300 58812
rect 134944 58772 215300 58800
rect 134944 58760 134950 58772
rect 215294 58760 215300 58772
rect 215352 58760 215358 58812
rect 31018 58692 31024 58744
rect 31076 58732 31082 58744
rect 162854 58732 162860 58744
rect 31076 58704 162860 58732
rect 31076 58692 31082 58704
rect 162854 58692 162860 58704
rect 162912 58692 162918 58744
rect 143442 58624 143448 58676
rect 143500 58664 143506 58676
rect 545758 58664 545764 58676
rect 143500 58636 545764 58664
rect 143500 58624 143506 58636
rect 545758 58624 545764 58636
rect 545816 58624 545822 58676
rect 105630 57876 105636 57928
rect 105688 57916 105694 57928
rect 106182 57916 106188 57928
rect 105688 57888 106188 57916
rect 105688 57876 105694 57888
rect 106182 57876 106188 57888
rect 106240 57916 106246 57928
rect 140222 57916 140228 57928
rect 106240 57888 140228 57916
rect 106240 57876 106246 57888
rect 140222 57876 140228 57888
rect 140280 57876 140286 57928
rect 154666 57876 154672 57928
rect 154724 57916 154730 57928
rect 218054 57916 218060 57928
rect 154724 57888 218060 57916
rect 154724 57876 154730 57888
rect 218054 57876 218060 57888
rect 218112 57916 218118 57928
rect 218514 57916 218520 57928
rect 218112 57888 218520 57916
rect 218112 57876 218118 57888
rect 218514 57876 218520 57888
rect 218572 57876 218578 57928
rect 158438 57808 158444 57860
rect 158496 57848 158502 57860
rect 191926 57848 191932 57860
rect 158496 57820 191932 57848
rect 158496 57808 158502 57820
rect 191926 57808 191932 57820
rect 191984 57848 191990 57860
rect 193122 57848 193128 57860
rect 191984 57820 193128 57848
rect 191984 57808 191990 57820
rect 193122 57808 193128 57820
rect 193180 57808 193186 57860
rect 193122 57264 193128 57316
rect 193180 57304 193186 57316
rect 256694 57304 256700 57316
rect 193180 57276 256700 57304
rect 193180 57264 193186 57276
rect 256694 57264 256700 57276
rect 256752 57264 256758 57316
rect 71774 57196 71780 57248
rect 71832 57236 71838 57248
rect 105630 57236 105636 57248
rect 71832 57208 105636 57236
rect 71832 57196 71838 57208
rect 105630 57196 105636 57208
rect 105688 57196 105694 57248
rect 218054 57196 218060 57248
rect 218112 57236 218118 57248
rect 470594 57236 470600 57248
rect 218112 57208 470600 57236
rect 218112 57196 218118 57208
rect 470594 57196 470600 57208
rect 470652 57196 470658 57248
rect 150434 56584 150440 56636
rect 150492 56624 150498 56636
rect 151906 56624 151912 56636
rect 150492 56596 151912 56624
rect 150492 56584 150498 56596
rect 151906 56584 151912 56596
rect 151964 56584 151970 56636
rect 186222 56516 186228 56568
rect 186280 56556 186286 56568
rect 579890 56556 579896 56568
rect 186280 56528 579896 56556
rect 186280 56516 186286 56528
rect 579890 56516 579896 56528
rect 579948 56516 579954 56568
rect 164234 55972 164240 56024
rect 164292 56012 164298 56024
rect 184842 56012 184848 56024
rect 164292 55984 184848 56012
rect 164292 55972 164298 55984
rect 184842 55972 184848 55984
rect 184900 55972 184906 56024
rect 17954 55904 17960 55956
rect 18012 55944 18018 55956
rect 176010 55944 176016 55956
rect 18012 55916 176016 55944
rect 18012 55904 18018 55916
rect 176010 55904 176016 55916
rect 176068 55904 176074 55956
rect 141510 55836 141516 55888
rect 141568 55876 141574 55888
rect 345014 55876 345020 55888
rect 141568 55848 345020 55876
rect 141568 55836 141574 55848
rect 345014 55836 345020 55848
rect 345072 55836 345078 55888
rect 95050 55156 95056 55208
rect 95108 55196 95114 55208
rect 139946 55196 139952 55208
rect 95108 55168 139952 55196
rect 95108 55156 95114 55168
rect 139946 55156 139952 55168
rect 140004 55156 140010 55208
rect 165706 55156 165712 55208
rect 165764 55196 165770 55208
rect 200206 55196 200212 55208
rect 165764 55168 200212 55196
rect 165764 55156 165770 55168
rect 200206 55156 200212 55168
rect 200264 55196 200270 55208
rect 201402 55196 201408 55208
rect 200264 55168 201408 55196
rect 200264 55156 200270 55168
rect 201402 55156 201408 55168
rect 201460 55156 201466 55208
rect 184842 55088 184848 55140
rect 184900 55128 184906 55140
rect 199102 55128 199108 55140
rect 184900 55100 199108 55128
rect 184900 55088 184906 55100
rect 199102 55088 199108 55100
rect 199160 55088 199166 55140
rect 145650 54544 145656 54596
rect 145708 54584 145714 54596
rect 234614 54584 234620 54596
rect 145708 54556 234620 54584
rect 145708 54544 145714 54556
rect 234614 54544 234620 54556
rect 234672 54544 234678 54596
rect 48314 54476 48320 54528
rect 48372 54516 48378 54528
rect 95050 54516 95056 54528
rect 48372 54488 95056 54516
rect 48372 54476 48378 54488
rect 95050 54476 95056 54488
rect 95108 54476 95114 54528
rect 201402 54476 201408 54528
rect 201460 54516 201466 54528
rect 578878 54516 578884 54528
rect 201460 54488 578884 54516
rect 201460 54476 201466 54488
rect 578878 54476 578884 54488
rect 578936 54476 578942 54528
rect 167086 53728 167092 53780
rect 167144 53768 167150 53780
rect 201494 53768 201500 53780
rect 167144 53740 201500 53768
rect 167144 53728 167150 53740
rect 201494 53728 201500 53740
rect 201552 53768 201558 53780
rect 202782 53768 202788 53780
rect 201552 53740 202788 53768
rect 201552 53728 201558 53740
rect 202782 53728 202788 53740
rect 202840 53728 202846 53780
rect 202782 53116 202788 53168
rect 202840 53156 202846 53168
rect 276014 53156 276020 53168
rect 202840 53128 276020 53156
rect 202840 53116 202846 53128
rect 276014 53116 276020 53128
rect 276072 53116 276078 53168
rect 147122 53048 147128 53100
rect 147180 53088 147186 53100
rect 542354 53088 542360 53100
rect 147180 53060 542360 53088
rect 147180 53048 147186 53060
rect 542354 53048 542360 53060
rect 542412 53048 542418 53100
rect 3510 52368 3516 52420
rect 3568 52408 3574 52420
rect 8938 52408 8944 52420
rect 3568 52380 8944 52408
rect 3568 52368 3574 52380
rect 8938 52368 8944 52380
rect 8996 52368 9002 52420
rect 182910 52368 182916 52420
rect 182968 52408 182974 52420
rect 579890 52408 579896 52420
rect 182968 52380 579896 52408
rect 182968 52368 182974 52380
rect 579890 52368 579896 52380
rect 579948 52368 579954 52420
rect 154390 51756 154396 51808
rect 154448 51796 154454 51808
rect 186222 51796 186228 51808
rect 154448 51768 186228 51796
rect 154448 51756 154454 51768
rect 186222 51756 186228 51768
rect 186280 51796 186286 51808
rect 188706 51796 188712 51808
rect 186280 51768 188712 51796
rect 186280 51756 186286 51768
rect 188706 51756 188712 51768
rect 188764 51756 188770 51808
rect 133230 51688 133236 51740
rect 133288 51728 133294 51740
rect 502978 51728 502984 51740
rect 133288 51700 502984 51728
rect 133288 51688 133294 51700
rect 502978 51688 502984 51700
rect 503036 51688 503042 51740
rect 135990 51008 135996 51060
rect 136048 51048 136054 51060
rect 144178 51048 144184 51060
rect 136048 51020 144184 51048
rect 136048 51008 136054 51020
rect 144178 51008 144184 51020
rect 144236 51008 144242 51060
rect 166994 51008 167000 51060
rect 167052 51048 167058 51060
rect 196158 51048 196164 51060
rect 167052 51020 196164 51048
rect 167052 51008 167058 51020
rect 196158 51008 196164 51020
rect 196216 51008 196222 51060
rect 144362 50396 144368 50448
rect 144420 50436 144426 50448
rect 400858 50436 400864 50448
rect 144420 50408 400864 50436
rect 144420 50396 144426 50408
rect 400858 50396 400864 50408
rect 400916 50396 400922 50448
rect 196158 50328 196164 50380
rect 196216 50368 196222 50380
rect 553394 50368 553400 50380
rect 196216 50340 553400 50368
rect 196216 50328 196222 50340
rect 553394 50328 553400 50340
rect 553452 50328 553458 50380
rect 169754 49648 169760 49700
rect 169812 49688 169818 49700
rect 173158 49688 173164 49700
rect 169812 49660 173164 49688
rect 169812 49648 169818 49660
rect 173158 49648 173164 49660
rect 173216 49648 173222 49700
rect 174538 49648 174544 49700
rect 174596 49688 174602 49700
rect 199194 49688 199200 49700
rect 174596 49660 199200 49688
rect 174596 49648 174602 49660
rect 199194 49648 199200 49660
rect 199252 49688 199258 49700
rect 580166 49688 580172 49700
rect 199252 49660 580172 49688
rect 199252 49648 199258 49660
rect 580166 49648 580172 49660
rect 580224 49648 580230 49700
rect 140130 48968 140136 49020
rect 140188 49008 140194 49020
rect 374638 49008 374644 49020
rect 140188 48980 374644 49008
rect 140188 48968 140194 48980
rect 374638 48968 374644 48980
rect 374696 48968 374702 49020
rect 3510 48220 3516 48272
rect 3568 48260 3574 48272
rect 122098 48260 122104 48272
rect 3568 48232 122104 48260
rect 3568 48220 3574 48232
rect 122098 48220 122104 48232
rect 122156 48260 122162 48272
rect 144454 48260 144460 48272
rect 122156 48232 144460 48260
rect 122156 48220 122162 48232
rect 144454 48220 144460 48232
rect 144512 48220 144518 48272
rect 150894 48220 150900 48272
rect 150952 48260 150958 48272
rect 220814 48260 220820 48272
rect 150952 48232 220820 48260
rect 150952 48220 150958 48232
rect 220814 48220 220820 48232
rect 220872 48260 220878 48272
rect 222102 48260 222108 48272
rect 220872 48232 222108 48260
rect 220872 48220 220878 48232
rect 222102 48220 222108 48232
rect 222160 48220 222166 48272
rect 169846 48152 169852 48204
rect 169904 48192 169910 48204
rect 203242 48192 203248 48204
rect 169904 48164 203248 48192
rect 169904 48152 169910 48164
rect 203242 48152 203248 48164
rect 203300 48192 203306 48204
rect 204162 48192 204168 48204
rect 203300 48164 204168 48192
rect 203300 48152 203306 48164
rect 204162 48152 204168 48164
rect 204220 48152 204226 48204
rect 204162 47608 204168 47660
rect 204220 47648 204226 47660
rect 284294 47648 284300 47660
rect 204220 47620 284300 47648
rect 204220 47608 204226 47620
rect 284294 47608 284300 47620
rect 284352 47608 284358 47660
rect 222102 47540 222108 47592
rect 222160 47580 222166 47592
rect 420914 47580 420920 47592
rect 222160 47552 420920 47580
rect 222160 47540 222166 47552
rect 420914 47540 420920 47552
rect 420972 47540 420978 47592
rect 168374 46860 168380 46912
rect 168432 46900 168438 46912
rect 203150 46900 203156 46912
rect 168432 46872 203156 46900
rect 168432 46860 168438 46872
rect 203150 46860 203156 46872
rect 203208 46900 203214 46912
rect 204162 46900 204168 46912
rect 203208 46872 204168 46900
rect 203208 46860 203214 46872
rect 204162 46860 204168 46872
rect 204220 46860 204226 46912
rect 171134 46792 171140 46844
rect 171192 46832 171198 46844
rect 205634 46832 205640 46844
rect 171192 46804 205640 46832
rect 171192 46792 171198 46804
rect 205634 46792 205640 46804
rect 205692 46792 205698 46844
rect 205634 46248 205640 46300
rect 205692 46288 205698 46300
rect 230474 46288 230480 46300
rect 205692 46260 230480 46288
rect 205692 46248 205698 46260
rect 230474 46248 230480 46260
rect 230532 46248 230538 46300
rect 204162 46180 204168 46232
rect 204220 46220 204226 46232
rect 556798 46220 556804 46232
rect 204220 46192 556804 46220
rect 204220 46180 204226 46192
rect 556798 46180 556804 46192
rect 556856 46180 556862 46232
rect 153930 45500 153936 45552
rect 153988 45540 153994 45552
rect 579982 45540 579988 45552
rect 153988 45512 579988 45540
rect 153988 45500 153994 45512
rect 579982 45500 579988 45512
rect 580040 45500 580046 45552
rect 137370 44820 137376 44872
rect 137428 44860 137434 44872
rect 436094 44860 436100 44872
rect 137428 44832 436100 44860
rect 137428 44820 137434 44832
rect 436094 44820 436100 44832
rect 436152 44820 436158 44872
rect 3510 44072 3516 44124
rect 3568 44112 3574 44124
rect 103422 44112 103428 44124
rect 3568 44084 103428 44112
rect 3568 44072 3574 44084
rect 103422 44072 103428 44084
rect 103480 44112 103486 44124
rect 131758 44112 131764 44124
rect 103480 44084 131764 44112
rect 103480 44072 103486 44084
rect 131758 44072 131764 44084
rect 131816 44072 131822 44124
rect 147030 43460 147036 43512
rect 147088 43500 147094 43512
rect 394694 43500 394700 43512
rect 147088 43472 394700 43500
rect 147088 43460 147094 43472
rect 394694 43460 394700 43472
rect 394752 43460 394758 43512
rect 138842 43392 138848 43444
rect 138900 43432 138906 43444
rect 557534 43432 557540 43444
rect 138900 43404 557540 43432
rect 138900 43392 138906 43404
rect 557534 43392 557540 43404
rect 557592 43392 557598 43444
rect 133138 42100 133144 42152
rect 133196 42140 133202 42152
rect 377398 42140 377404 42152
rect 133196 42112 377404 42140
rect 133196 42100 133202 42112
rect 377398 42100 377404 42112
rect 377456 42100 377462 42152
rect 148410 42032 148416 42084
rect 148468 42072 148474 42084
rect 503714 42072 503720 42084
rect 148468 42044 503720 42072
rect 148468 42032 148474 42044
rect 503714 42032 503720 42044
rect 503772 42032 503778 42084
rect 158254 41352 158260 41404
rect 158312 41392 158318 41404
rect 190454 41392 190460 41404
rect 158312 41364 190460 41392
rect 158312 41352 158318 41364
rect 190454 41352 190460 41364
rect 190512 41392 190518 41404
rect 580166 41392 580172 41404
rect 190512 41364 580172 41392
rect 190512 41352 190518 41364
rect 580166 41352 580172 41364
rect 580224 41352 580230 41404
rect 138750 40672 138756 40724
rect 138808 40712 138814 40724
rect 390554 40712 390560 40724
rect 138808 40684 390560 40712
rect 138808 40672 138814 40684
rect 390554 40672 390560 40684
rect 390612 40672 390618 40724
rect 3510 39992 3516 40044
rect 3568 40032 3574 40044
rect 126238 40032 126244 40044
rect 3568 40004 126244 40032
rect 3568 39992 3574 40004
rect 126238 39992 126244 40004
rect 126296 39992 126302 40044
rect 164050 39380 164056 39432
rect 164108 39420 164114 39432
rect 245654 39420 245660 39432
rect 164108 39392 245660 39420
rect 164108 39380 164114 39392
rect 245654 39380 245660 39392
rect 245712 39380 245718 39432
rect 176562 39312 176568 39364
rect 176620 39352 176626 39364
rect 340874 39352 340880 39364
rect 176620 39324 340880 39352
rect 176620 39312 176626 39324
rect 340874 39312 340880 39324
rect 340932 39312 340938 39364
rect 155586 38564 155592 38616
rect 155644 38604 155650 38616
rect 189166 38604 189172 38616
rect 155644 38576 189172 38604
rect 155644 38564 155650 38576
rect 189166 38564 189172 38576
rect 189224 38604 189230 38616
rect 189626 38604 189632 38616
rect 189224 38576 189632 38604
rect 189224 38564 189230 38576
rect 189626 38564 189632 38576
rect 189684 38564 189690 38616
rect 189166 37952 189172 38004
rect 189224 37992 189230 38004
rect 378134 37992 378140 38004
rect 189224 37964 378140 37992
rect 189224 37952 189230 37964
rect 378134 37952 378140 37964
rect 378192 37952 378198 38004
rect 137278 37884 137284 37936
rect 137336 37924 137342 37936
rect 442258 37924 442264 37936
rect 137336 37896 442264 37924
rect 137336 37884 137342 37896
rect 442258 37884 442264 37896
rect 442316 37884 442322 37936
rect 3142 37204 3148 37256
rect 3200 37244 3206 37256
rect 133874 37244 133880 37256
rect 3200 37216 133880 37244
rect 3200 37204 3206 37216
rect 133874 37204 133880 37216
rect 133932 37204 133938 37256
rect 192478 37204 192484 37256
rect 192536 37244 192542 37256
rect 580166 37244 580172 37256
rect 192536 37216 580172 37244
rect 192536 37204 192542 37216
rect 580166 37204 580172 37216
rect 580224 37204 580230 37256
rect 144270 36524 144276 36576
rect 144328 36564 144334 36576
rect 219434 36564 219440 36576
rect 144328 36536 219440 36564
rect 144328 36524 144334 36536
rect 219434 36524 219440 36536
rect 219492 36524 219498 36576
rect 158530 35232 158536 35284
rect 158588 35272 158594 35284
rect 371234 35272 371240 35284
rect 158588 35244 371240 35272
rect 158588 35232 158594 35244
rect 371234 35232 371240 35244
rect 371292 35232 371298 35284
rect 168282 35164 168288 35216
rect 168340 35204 168346 35216
rect 548518 35204 548524 35216
rect 168340 35176 548524 35204
rect 168340 35164 168346 35176
rect 548518 35164 548524 35176
rect 548576 35164 548582 35216
rect 158714 34416 158720 34468
rect 158772 34456 158778 34468
rect 190546 34456 190552 34468
rect 158772 34428 190552 34456
rect 158772 34416 158778 34428
rect 190546 34416 190552 34428
rect 190604 34456 190610 34468
rect 191742 34456 191748 34468
rect 190604 34428 191748 34456
rect 190604 34416 190610 34428
rect 191742 34416 191748 34428
rect 191800 34416 191806 34468
rect 161474 34348 161480 34400
rect 161532 34388 161538 34400
rect 191926 34388 191932 34400
rect 161532 34360 191932 34388
rect 161532 34348 161538 34360
rect 191926 34348 191932 34360
rect 191984 34388 191990 34400
rect 193122 34388 193128 34400
rect 191984 34360 193128 34388
rect 191984 34348 191990 34360
rect 193122 34348 193128 34360
rect 193180 34348 193186 34400
rect 191742 33736 191748 33788
rect 191800 33776 191806 33788
rect 356054 33776 356060 33788
rect 191800 33748 356060 33776
rect 191800 33736 191806 33748
rect 356054 33736 356060 33748
rect 356112 33736 356118 33788
rect 193122 33124 193128 33176
rect 193180 33164 193186 33176
rect 571978 33164 571984 33176
rect 193180 33136 571984 33164
rect 193180 33124 193186 33136
rect 571978 33124 571984 33136
rect 572036 33124 572042 33176
rect 152458 33056 152464 33108
rect 152516 33096 152522 33108
rect 580166 33096 580172 33108
rect 152516 33068 580172 33096
rect 152516 33056 152522 33068
rect 580166 33056 580172 33068
rect 580224 33056 580230 33108
rect 161198 31084 161204 31136
rect 161256 31124 161262 31136
rect 364334 31124 364340 31136
rect 161256 31096 364340 31124
rect 161256 31084 161262 31096
rect 364334 31084 364340 31096
rect 364392 31084 364398 31136
rect 166718 31016 166724 31068
rect 166776 31056 166782 31068
rect 563698 31056 563704 31068
rect 166776 31028 563704 31056
rect 166776 31016 166782 31028
rect 563698 31016 563704 31028
rect 563756 31016 563762 31068
rect 154022 30268 154028 30320
rect 154080 30308 154086 30320
rect 189166 30308 189172 30320
rect 154080 30280 189172 30308
rect 154080 30268 154086 30280
rect 189166 30268 189172 30280
rect 189224 30268 189230 30320
rect 165430 29656 165436 29708
rect 165488 29696 165494 29708
rect 332594 29696 332600 29708
rect 165488 29668 332600 29696
rect 165488 29656 165494 29668
rect 332594 29656 332600 29668
rect 332652 29656 332658 29708
rect 189166 29588 189172 29640
rect 189224 29628 189230 29640
rect 189902 29628 189908 29640
rect 189224 29600 189908 29628
rect 189224 29588 189230 29600
rect 189902 29588 189908 29600
rect 189960 29628 189966 29640
rect 500218 29628 500224 29640
rect 189960 29600 500224 29628
rect 189960 29588 189966 29600
rect 500218 29588 500224 29600
rect 500276 29588 500282 29640
rect 3142 28908 3148 28960
rect 3200 28948 3206 28960
rect 138198 28948 138204 28960
rect 3200 28920 138204 28948
rect 3200 28908 3206 28920
rect 138198 28908 138204 28920
rect 138256 28908 138262 28960
rect 188982 28908 188988 28960
rect 189040 28948 189046 28960
rect 580166 28948 580172 28960
rect 189040 28920 580172 28948
rect 189040 28908 189046 28920
rect 580166 28908 580172 28920
rect 580224 28908 580230 28960
rect 141418 28228 141424 28280
rect 141476 28268 141482 28280
rect 207658 28268 207664 28280
rect 141476 28240 207664 28268
rect 141476 28228 141482 28240
rect 207658 28228 207664 28240
rect 207716 28228 207722 28280
rect 166810 26936 166816 26988
rect 166868 26976 166874 26988
rect 249794 26976 249800 26988
rect 166868 26948 249800 26976
rect 166868 26936 166874 26948
rect 249794 26936 249800 26948
rect 249852 26936 249858 26988
rect 148318 26868 148324 26920
rect 148376 26908 148382 26920
rect 347774 26908 347780 26920
rect 148376 26880 347780 26908
rect 148376 26868 148382 26880
rect 347774 26868 347780 26880
rect 347832 26868 347838 26920
rect 162670 25508 162676 25560
rect 162728 25548 162734 25560
rect 473354 25548 473360 25560
rect 162728 25520 473360 25548
rect 162728 25508 162734 25520
rect 473354 25508 473360 25520
rect 473412 25508 473418 25560
rect 182082 24760 182088 24812
rect 182140 24800 182146 24812
rect 580166 24800 580172 24812
rect 182140 24772 580172 24800
rect 182140 24760 182146 24772
rect 580166 24760 580172 24772
rect 580224 24760 580230 24812
rect 134702 24080 134708 24132
rect 134760 24120 134766 24132
rect 210418 24120 210424 24132
rect 134760 24092 210424 24120
rect 134760 24080 134766 24092
rect 210418 24080 210424 24092
rect 210476 24080 210482 24132
rect 171042 22720 171048 22772
rect 171100 22760 171106 22772
rect 514018 22760 514024 22772
rect 171100 22732 514024 22760
rect 171100 22720 171106 22732
rect 514018 22720 514024 22732
rect 514076 22720 514082 22772
rect 166902 21360 166908 21412
rect 166960 21400 166966 21412
rect 466454 21400 466460 21412
rect 166960 21372 466460 21400
rect 166960 21360 166966 21372
rect 466454 21360 466460 21372
rect 466512 21360 466518 21412
rect 3142 20612 3148 20664
rect 3200 20652 3206 20664
rect 139578 20652 139584 20664
rect 3200 20624 139584 20652
rect 3200 20612 3206 20624
rect 139578 20612 139584 20624
rect 139636 20612 139642 20664
rect 161290 20612 161296 20664
rect 161348 20652 161354 20664
rect 580166 20652 580172 20664
rect 161348 20624 580172 20652
rect 161348 20612 161354 20624
rect 580166 20612 580172 20624
rect 580224 20612 580230 20664
rect 146938 18640 146944 18692
rect 146996 18680 147002 18692
rect 226334 18680 226340 18692
rect 146996 18652 226340 18680
rect 146996 18640 147002 18652
rect 226334 18640 226340 18652
rect 226392 18640 226398 18692
rect 175090 18572 175096 18624
rect 175148 18612 175154 18624
rect 481634 18612 481640 18624
rect 175148 18584 481640 18612
rect 175148 18572 175154 18584
rect 481634 18572 481640 18584
rect 481692 18572 481698 18624
rect 161382 17212 161388 17264
rect 161440 17252 161446 17264
rect 527174 17252 527180 17264
rect 161440 17224 527180 17252
rect 161440 17212 161446 17224
rect 527174 17212 527180 17224
rect 527232 17212 527238 17264
rect 3326 16532 3332 16584
rect 3384 16572 3390 16584
rect 131114 16572 131120 16584
rect 3384 16544 131120 16572
rect 3384 16532 3390 16544
rect 131114 16532 131120 16544
rect 131172 16532 131178 16584
rect 182818 16532 182824 16584
rect 182876 16572 182882 16584
rect 580166 16572 580172 16584
rect 182876 16544 580172 16572
rect 182876 16532 182882 16544
rect 580166 16532 580172 16544
rect 580224 16532 580230 16584
rect 156690 15852 156696 15904
rect 156748 15892 156754 15904
rect 178402 15892 178408 15904
rect 156748 15864 178408 15892
rect 156748 15852 156754 15864
rect 178402 15852 178408 15864
rect 178460 15852 178466 15904
rect 153838 14560 153844 14612
rect 153896 14600 153902 14612
rect 204346 14600 204352 14612
rect 153896 14572 204352 14600
rect 153896 14560 153902 14572
rect 204346 14560 204352 14572
rect 204404 14560 204410 14612
rect 172330 14492 172336 14544
rect 172388 14532 172394 14544
rect 352466 14532 352472 14544
rect 172388 14504 352472 14532
rect 172388 14492 172394 14504
rect 352466 14492 352472 14504
rect 352524 14492 352530 14544
rect 140038 14424 140044 14476
rect 140096 14464 140102 14476
rect 459186 14464 459192 14476
rect 140096 14436 459192 14464
rect 140096 14424 140102 14436
rect 459186 14424 459192 14436
rect 459244 14424 459250 14476
rect 162946 13200 162952 13252
rect 163004 13240 163010 13252
rect 175918 13240 175924 13252
rect 163004 13212 175924 13240
rect 163004 13200 163010 13212
rect 175918 13200 175924 13212
rect 175976 13200 175982 13252
rect 175182 13132 175188 13184
rect 175240 13172 175246 13184
rect 447594 13172 447600 13184
rect 175240 13144 447600 13172
rect 175240 13132 175246 13144
rect 447594 13132 447600 13144
rect 447652 13132 447658 13184
rect 134518 13064 134524 13116
rect 134576 13104 134582 13116
rect 531314 13104 531320 13116
rect 134576 13076 531320 13104
rect 134576 13064 134582 13076
rect 531314 13064 531320 13076
rect 531372 13064 531378 13116
rect 3050 12384 3056 12436
rect 3108 12424 3114 12436
rect 129734 12424 129740 12436
rect 3108 12396 129740 12424
rect 3108 12384 3114 12396
rect 129734 12384 129740 12396
rect 129792 12384 129798 12436
rect 186222 12384 186228 12436
rect 186280 12424 186286 12436
rect 580166 12424 580172 12436
rect 186280 12396 580172 12424
rect 186280 12384 186286 12396
rect 580166 12384 580172 12396
rect 580224 12384 580230 12436
rect 149698 11704 149704 11756
rect 149756 11744 149762 11756
rect 193214 11744 193220 11756
rect 149756 11716 193220 11744
rect 149756 11704 149762 11716
rect 193214 11704 193220 11716
rect 193272 11704 193278 11756
rect 172422 10344 172428 10396
rect 172480 10384 172486 10396
rect 299474 10384 299480 10396
rect 172480 10356 299480 10384
rect 172480 10344 172486 10356
rect 299474 10344 299480 10356
rect 299532 10344 299538 10396
rect 157242 10276 157248 10328
rect 157300 10316 157306 10328
rect 562318 10316 562324 10328
rect 157300 10288 562324 10316
rect 157300 10276 157306 10288
rect 562318 10276 562324 10288
rect 562376 10276 562382 10328
rect 134610 8916 134616 8968
rect 134668 8956 134674 8968
rect 241698 8956 241704 8968
rect 134668 8928 241704 8956
rect 134668 8916 134674 8928
rect 241698 8916 241704 8928
rect 241756 8916 241762 8968
rect 2958 8236 2964 8288
rect 3016 8276 3022 8288
rect 151814 8276 151820 8288
rect 3016 8248 151820 8276
rect 3016 8236 3022 8248
rect 151814 8236 151820 8248
rect 151872 8236 151878 8288
rect 560938 8236 560944 8288
rect 560996 8276 561002 8288
rect 580166 8276 580172 8288
rect 560996 8248 580172 8276
rect 560996 8236 561002 8248
rect 580166 8236 580172 8248
rect 580224 8236 580230 8288
rect 162578 7624 162584 7676
rect 162636 7664 162642 7676
rect 318794 7664 318800 7676
rect 162636 7636 318800 7664
rect 162636 7624 162642 7636
rect 318794 7624 318800 7636
rect 318852 7624 318858 7676
rect 164142 7556 164148 7608
rect 164200 7596 164206 7608
rect 360654 7596 360660 7608
rect 164200 7568 360660 7596
rect 164200 7556 164206 7568
rect 360654 7556 360660 7568
rect 360712 7556 360718 7608
rect 110138 6196 110144 6248
rect 110196 6236 110202 6248
rect 147674 6236 147680 6248
rect 110196 6208 147680 6236
rect 110196 6196 110202 6208
rect 147674 6196 147680 6208
rect 147732 6196 147738 6248
rect 158622 6196 158628 6248
rect 158680 6236 158686 6248
rect 398650 6236 398656 6248
rect 158680 6208 398656 6236
rect 158680 6196 158686 6208
rect 398650 6196 398656 6208
rect 398708 6196 398714 6248
rect 138658 6128 138664 6180
rect 138716 6168 138722 6180
rect 432782 6168 432788 6180
rect 138716 6140 432788 6168
rect 138716 6128 138722 6140
rect 432782 6128 432788 6140
rect 432840 6128 432846 6180
rect 184842 5448 184848 5500
rect 184900 5488 184906 5500
rect 580166 5488 580172 5500
rect 184900 5460 580172 5488
rect 184900 5448 184906 5460
rect 580166 5448 580172 5460
rect 580224 5448 580230 5500
rect 145558 4768 145564 4820
rect 145616 4808 145622 4820
rect 155218 4808 155224 4820
rect 145616 4780 155224 4808
rect 145616 4768 145622 4780
rect 155218 4768 155224 4780
rect 155276 4768 155282 4820
rect 165522 4768 165528 4820
rect 165580 4808 165586 4820
rect 280798 4808 280804 4820
rect 165580 4780 280804 4808
rect 165580 4768 165586 4780
rect 280798 4768 280804 4780
rect 280856 4768 280862 4820
rect 2774 4020 2780 4072
rect 2832 4060 2838 4072
rect 4798 4060 4804 4072
rect 2832 4032 4804 4060
rect 2832 4020 2838 4032
rect 4798 4020 4804 4032
rect 4856 4020 4862 4072
rect 117222 3544 117228 3596
rect 117280 3584 117286 3596
rect 156598 3584 156604 3596
rect 117280 3556 156604 3584
rect 117280 3544 117286 3556
rect 156598 3544 156604 3556
rect 156656 3544 156662 3596
rect 165614 3544 165620 3596
rect 165672 3584 165678 3596
rect 166810 3584 166816 3596
rect 165672 3556 166816 3584
rect 165672 3544 165678 3556
rect 166810 3544 166816 3556
rect 166868 3544 166874 3596
rect 174538 3544 174544 3596
rect 174596 3584 174602 3596
rect 191834 3584 191840 3596
rect 174596 3556 191840 3584
rect 174596 3544 174602 3556
rect 191834 3544 191840 3556
rect 191892 3544 191898 3596
rect 207658 3544 207664 3596
rect 207716 3584 207722 3596
rect 208670 3584 208676 3596
rect 207716 3556 208676 3584
rect 207716 3544 207722 3556
rect 208670 3544 208676 3556
rect 208728 3544 208734 3596
rect 210418 3544 210424 3596
rect 210476 3584 210482 3596
rect 242802 3584 242808 3596
rect 210476 3556 242808 3584
rect 210476 3544 210482 3556
rect 242802 3544 242808 3556
rect 242860 3544 242866 3596
rect 377398 3544 377404 3596
rect 377456 3584 377462 3596
rect 377456 3556 383654 3584
rect 377456 3544 377462 3556
rect 30282 3476 30288 3528
rect 30340 3516 30346 3528
rect 31018 3516 31024 3528
rect 30340 3488 31024 3516
rect 30340 3476 30346 3488
rect 31018 3476 31024 3488
rect 31076 3476 31082 3528
rect 34146 3476 34152 3528
rect 34204 3516 34210 3528
rect 35158 3516 35164 3528
rect 34204 3488 35164 3516
rect 34204 3476 34210 3488
rect 35158 3476 35164 3488
rect 35216 3476 35222 3528
rect 97902 3476 97908 3528
rect 97960 3516 97966 3528
rect 128814 3516 128820 3528
rect 97960 3488 128820 3516
rect 97960 3476 97966 3488
rect 128814 3476 128820 3488
rect 128872 3476 128878 3528
rect 136542 3476 136548 3528
rect 136600 3516 136606 3528
rect 211246 3516 211252 3528
rect 136600 3488 211252 3516
rect 136600 3476 136606 3488
rect 211246 3476 211252 3488
rect 211304 3476 211310 3528
rect 211798 3476 211804 3528
rect 211856 3516 211862 3528
rect 212534 3516 212540 3528
rect 211856 3488 212540 3516
rect 211856 3476 211862 3488
rect 212534 3476 212540 3488
rect 212592 3476 212598 3528
rect 241698 3476 241704 3528
rect 241756 3516 241762 3528
rect 326522 3516 326528 3528
rect 241756 3488 326528 3516
rect 241756 3476 241762 3488
rect 326522 3476 326528 3488
rect 326580 3476 326586 3528
rect 374638 3476 374644 3528
rect 374696 3516 374702 3528
rect 375466 3516 375472 3528
rect 374696 3488 375472 3516
rect 374696 3476 374702 3488
rect 375466 3476 375472 3488
rect 375524 3476 375530 3528
rect 378134 3476 378140 3528
rect 378192 3516 378198 3528
rect 379330 3516 379336 3528
rect 378192 3488 379336 3516
rect 378192 3476 378198 3488
rect 379330 3476 379336 3488
rect 379388 3476 379394 3528
rect 383626 3516 383654 3556
rect 508774 3516 508780 3528
rect 383626 3488 508780 3516
rect 508774 3476 508780 3488
rect 508832 3476 508838 3528
rect 545758 3476 545764 3528
rect 545816 3516 545822 3528
rect 546770 3516 546776 3528
rect 545816 3488 546776 3516
rect 545816 3476 545822 3488
rect 546770 3476 546776 3488
rect 546828 3476 546834 3528
rect 571978 3476 571984 3528
rect 572036 3516 572042 3528
rect 573174 3516 573180 3528
rect 572036 3488 573180 3516
rect 572036 3476 572042 3488
rect 573174 3476 573180 3488
rect 573232 3476 573238 3528
rect 14 3408 20 3460
rect 72 3448 78 3460
rect 13078 3448 13084 3460
rect 72 3420 13084 3448
rect 72 3408 78 3420
rect 13078 3408 13084 3420
rect 13136 3408 13142 3460
rect 14826 3408 14832 3460
rect 14884 3448 14890 3460
rect 135438 3448 135444 3460
rect 14884 3420 135444 3448
rect 14884 3408 14890 3420
rect 135438 3408 135444 3420
rect 135496 3408 135502 3460
rect 142798 3408 142804 3460
rect 142856 3448 142862 3460
rect 144270 3448 144276 3460
rect 142856 3420 144276 3448
rect 142856 3408 142862 3420
rect 144270 3408 144276 3420
rect 144328 3408 144334 3460
rect 146294 3408 146300 3460
rect 146352 3448 146358 3460
rect 147490 3448 147496 3460
rect 146352 3420 147496 3448
rect 146352 3408 146358 3420
rect 147490 3408 147496 3420
rect 147548 3408 147554 3460
rect 383194 3448 383200 3460
rect 151786 3420 383200 3448
rect 144178 3340 144184 3392
rect 144236 3380 144242 3392
rect 151786 3380 151814 3420
rect 383194 3408 383200 3420
rect 383252 3408 383258 3460
rect 400858 3408 400864 3460
rect 400916 3448 400922 3460
rect 402514 3448 402520 3460
rect 400916 3420 402520 3448
rect 400916 3408 400922 3420
rect 402514 3408 402520 3420
rect 402572 3408 402578 3460
rect 442258 3408 442264 3460
rect 442316 3448 442322 3460
rect 443730 3448 443736 3460
rect 442316 3420 443736 3448
rect 442316 3408 442322 3420
rect 443730 3408 443736 3420
rect 443788 3408 443794 3460
rect 454034 3408 454040 3460
rect 454092 3448 454098 3460
rect 455322 3448 455328 3460
rect 454092 3420 455328 3448
rect 454092 3408 454098 3420
rect 455322 3408 455328 3420
rect 455380 3408 455386 3460
rect 473354 3408 473360 3460
rect 473412 3448 473418 3460
rect 474642 3448 474648 3460
rect 473412 3420 474648 3448
rect 473412 3408 473418 3420
rect 474642 3408 474648 3420
rect 474700 3408 474706 3460
rect 496078 3408 496084 3460
rect 496136 3448 496142 3460
rect 497182 3448 497188 3460
rect 496136 3420 497188 3448
rect 496136 3408 496142 3420
rect 497182 3408 497188 3420
rect 497240 3408 497246 3460
rect 502978 3408 502984 3460
rect 503036 3448 503042 3460
rect 539042 3448 539048 3460
rect 503036 3420 539048 3448
rect 503036 3408 503042 3420
rect 539042 3408 539048 3420
rect 539100 3408 539106 3460
rect 556798 3408 556804 3460
rect 556856 3448 556862 3460
rect 561582 3448 561588 3460
rect 556856 3420 561588 3448
rect 556856 3408 556862 3420
rect 561582 3408 561588 3420
rect 561640 3408 561646 3460
rect 562318 3408 562324 3460
rect 562376 3448 562382 3460
rect 562376 3420 567194 3448
rect 562376 3408 562382 3420
rect 144236 3352 151814 3380
rect 567166 3380 567194 3420
rect 577038 3380 577044 3392
rect 567166 3352 577044 3380
rect 144236 3340 144242 3352
rect 577038 3340 577044 3352
rect 577096 3340 577102 3392
rect 135898 3272 135904 3324
rect 135956 3312 135962 3324
rect 140406 3312 140412 3324
rect 135956 3284 140412 3312
rect 135956 3272 135962 3284
rect 140406 3272 140412 3284
rect 140464 3272 140470 3324
rect 548518 3068 548524 3120
rect 548576 3108 548582 3120
rect 550634 3108 550640 3120
rect 548576 3080 550640 3108
rect 548576 3068 548582 3080
rect 550634 3068 550640 3080
rect 550692 3068 550698 3120
rect 514018 3000 514024 3052
rect 514076 3040 514082 3052
rect 515858 3040 515864 3052
rect 514076 3012 515864 3040
rect 514076 3000 514082 3012
rect 515858 3000 515864 3012
rect 515916 3000 515922 3052
rect 563698 3000 563704 3052
rect 563756 3040 563762 3052
rect 565446 3040 565452 3052
rect 563756 3012 565452 3040
rect 563756 3000 563762 3012
rect 565446 3000 565452 3012
rect 565504 3000 565510 3052
rect 500218 2864 500224 2916
rect 500276 2904 500282 2916
rect 501046 2904 501052 2916
rect 500276 2876 501052 2904
rect 500276 2864 500282 2876
rect 501046 2864 501052 2876
rect 501104 2864 501110 2916
<< via1 >>
rect 30380 702992 30432 703044
rect 31576 702992 31628 703044
rect 405740 702992 405792 703044
rect 407028 702992 407080 703044
rect 425060 702992 425112 703044
rect 426348 702992 426400 703044
rect 436100 702992 436152 703044
rect 437296 702992 437348 703044
rect 455420 702992 455472 703044
rect 456616 702992 456668 703044
rect 544384 702448 544436 702500
rect 580172 702448 580224 702500
rect 3424 701020 3476 701072
rect 131120 701020 131172 701072
rect 88248 700680 88300 700732
rect 102784 700680 102836 700732
rect 65708 700612 65760 700664
rect 79324 700612 79376 700664
rect 80520 700612 80572 700664
rect 88984 700612 89036 700664
rect 95976 700612 96028 700664
rect 122840 700612 122892 700664
rect 4528 700544 4580 700596
rect 26884 700544 26936 700596
rect 46388 700544 46440 700596
rect 98736 700544 98788 700596
rect 179052 700544 179104 700596
rect 189540 700544 189592 700596
rect 19984 700476 20036 700528
rect 48964 700476 49016 700528
rect 54116 700476 54168 700528
rect 117964 700476 118016 700528
rect 133972 700476 134024 700528
rect 149704 700476 149756 700528
rect 168104 700476 168156 700528
rect 191840 700476 191892 700528
rect 23848 700408 23900 700460
rect 109040 700408 109092 700460
rect 117228 700408 117280 700460
rect 137836 700408 137888 700460
rect 164240 700408 164292 700460
rect 193220 700408 193272 700460
rect 543004 700408 543056 700460
rect 574468 700408 574520 700460
rect 12256 700340 12308 700392
rect 100116 700340 100168 700392
rect 115848 700340 115900 700392
rect 141700 700340 141752 700392
rect 175832 700340 175884 700392
rect 189448 700340 189500 700392
rect 189724 700340 189776 700392
rect 244096 700340 244148 700392
rect 514024 700340 514076 700392
rect 566740 700340 566792 700392
rect 664 700272 716 700324
rect 100024 700272 100076 700324
rect 120724 700272 120776 700324
rect 198372 700272 198424 700324
rect 239404 700272 239456 700324
rect 555148 700272 555200 700324
rect 190644 699728 190696 699780
rect 195980 699728 196032 699780
rect 42524 699660 42576 699712
rect 43444 699660 43496 699712
rect 144184 699660 144236 699712
rect 144920 699660 144972 699712
rect 192484 699660 192536 699712
rect 194508 699660 194560 699712
rect 260104 699660 260156 699712
rect 262772 699660 262824 699712
rect 305644 699660 305696 699712
rect 308496 699660 308548 699712
rect 309784 699660 309836 699712
rect 312360 699660 312412 699712
rect 313924 699660 313976 699712
rect 316224 699660 316276 699712
rect 327724 699660 327776 699712
rect 331036 699660 331088 699712
rect 359464 699660 359516 699712
rect 361948 699660 362000 699712
rect 377404 699660 377456 699712
rect 380624 699660 380676 699712
rect 381544 699660 381596 699712
rect 384488 699660 384540 699712
rect 428464 699660 428516 699712
rect 430212 699660 430264 699712
rect 431224 699660 431276 699712
rect 434076 699660 434128 699712
rect 476764 699660 476816 699712
rect 479156 699660 479208 699712
rect 548524 699660 548576 699712
rect 551284 699660 551336 699712
rect 558184 699660 558236 699712
rect 559012 699660 559064 699712
rect 16120 698912 16172 698964
rect 62764 698912 62816 698964
rect 199384 698300 199436 698352
rect 580172 698300 580224 698352
rect 67640 697552 67692 697604
rect 68928 697552 68980 697604
rect 531320 697552 531372 697604
rect 532608 697552 532660 697604
rect 3056 696940 3108 696992
rect 98644 696940 98696 696992
rect 299480 696600 299532 696652
rect 300768 696600 300820 696652
rect 512000 696600 512052 696652
rect 513288 696600 513340 696652
rect 559564 694152 559616 694204
rect 580172 694152 580224 694204
rect 552664 690004 552716 690056
rect 580172 690004 580224 690056
rect 3424 688644 3476 688696
rect 14464 688644 14516 688696
rect 556804 685856 556856 685908
rect 579804 685856 579856 685908
rect 3148 684496 3200 684548
rect 93124 684496 93176 684548
rect 552756 681708 552808 681760
rect 580172 681708 580224 681760
rect 3424 680348 3476 680400
rect 104164 680348 104216 680400
rect 566464 677560 566516 677612
rect 580172 677560 580224 677612
rect 3424 676200 3476 676252
rect 93308 676200 93360 676252
rect 200764 673480 200816 673532
rect 580172 673480 580224 673532
rect 548616 669332 548668 669384
rect 580172 669332 580224 669384
rect 3240 663756 3292 663808
rect 112444 663756 112496 663808
rect 3424 661036 3476 661088
rect 86224 661036 86276 661088
rect 541624 661036 541676 661088
rect 580172 661036 580224 661088
rect 124312 658248 124364 658300
rect 580172 658248 580224 658300
rect 566556 654100 566608 654152
rect 580172 654100 580224 654152
rect 3056 652740 3108 652792
rect 108304 652740 108356 652792
rect 179328 645872 179380 645924
rect 580172 645872 580224 645924
rect 3424 644444 3476 644496
rect 89076 644444 89128 644496
rect 558276 641724 558328 641776
rect 580172 641724 580224 641776
rect 3148 640296 3200 640348
rect 94504 640296 94556 640348
rect 3148 636216 3200 636268
rect 13084 636216 13136 636268
rect 3424 632068 3476 632120
rect 90364 632068 90416 632120
rect 570604 625132 570656 625184
rect 580172 625132 580224 625184
rect 3240 623772 3292 623824
rect 102876 623772 102928 623824
rect 3424 620984 3476 621036
rect 104256 620984 104308 621036
rect 576124 620984 576176 621036
rect 579804 620984 579856 621036
rect 3148 616836 3200 616888
rect 21364 616836 21416 616888
rect 3148 612756 3200 612808
rect 64144 612756 64196 612808
rect 120080 605820 120132 605872
rect 580172 605820 580224 605872
rect 3056 604460 3108 604512
rect 104348 604460 104400 604512
rect 560944 601672 560996 601724
rect 580172 601672 580224 601724
rect 3516 600312 3568 600364
rect 115940 600312 115992 600364
rect 3056 596164 3108 596216
rect 104900 596164 104952 596216
rect 3148 592016 3200 592068
rect 80704 592016 80756 592068
rect 574744 589296 574796 589348
rect 580172 589296 580224 589348
rect 3240 587868 3292 587920
rect 180800 587868 180852 587920
rect 3148 583720 3200 583772
rect 84844 583720 84896 583772
rect 3332 581000 3384 581052
rect 90456 581000 90508 581052
rect 3516 576852 3568 576904
rect 80796 576852 80848 576904
rect 2872 568556 2924 568608
rect 94596 568556 94648 568608
rect 562324 568556 562376 568608
rect 580172 568556 580224 568608
rect 130384 565836 130436 565888
rect 580172 565836 580224 565888
rect 3056 560260 3108 560312
rect 106924 560260 106976 560312
rect 3056 556180 3108 556232
rect 97264 556180 97316 556232
rect 576216 553392 576268 553444
rect 580172 553392 580224 553444
rect 3516 552032 3568 552084
rect 84936 552032 84988 552084
rect 571984 549244 572036 549296
rect 580172 549244 580224 549296
rect 3056 547884 3108 547936
rect 98828 547884 98880 547936
rect 558368 545096 558420 545148
rect 579896 545096 579948 545148
rect 3148 543736 3200 543788
rect 110512 543736 110564 543788
rect 3516 540948 3568 541000
rect 94688 540948 94740 541000
rect 565084 540948 565136 541000
rect 580172 540948 580224 541000
rect 3332 536800 3384 536852
rect 97356 536800 97408 536852
rect 120172 536800 120224 536852
rect 580172 536800 580224 536852
rect 3332 532720 3384 532772
rect 167092 532720 167144 532772
rect 577504 529048 577556 529100
rect 579804 529048 579856 529100
rect 3516 528572 3568 528624
rect 95884 528572 95936 528624
rect 3516 524424 3568 524476
rect 86316 524424 86368 524476
rect 555424 524424 555476 524476
rect 580172 524424 580224 524476
rect 2872 520276 2924 520328
rect 115204 520276 115256 520328
rect 189816 520276 189868 520328
rect 580172 520276 580224 520328
rect 2964 516128 3016 516180
rect 97448 516128 97500 516180
rect 3056 511980 3108 512032
rect 108396 511980 108448 512032
rect 574836 509260 574888 509312
rect 580172 509260 580224 509312
rect 3516 507832 3568 507884
rect 95976 507832 96028 507884
rect 138664 507832 138716 507884
rect 144184 507832 144236 507884
rect 554044 505112 554096 505164
rect 580080 505112 580132 505164
rect 3056 503684 3108 503736
rect 127164 503684 127216 503736
rect 576308 500964 576360 501016
rect 580080 500964 580132 501016
rect 3332 496816 3384 496868
rect 108488 496816 108540 496868
rect 554136 496816 554188 496868
rect 579896 496816 579948 496868
rect 3516 492668 3568 492720
rect 90548 492668 90600 492720
rect 574928 492668 574980 492720
rect 580172 492668 580224 492720
rect 3332 488520 3384 488572
rect 111064 488520 111116 488572
rect 566648 488520 566700 488572
rect 580172 488520 580224 488572
rect 3516 484372 3568 484424
rect 104440 484372 104492 484424
rect 215944 484372 215996 484424
rect 580172 484372 580224 484424
rect 3516 480224 3568 480276
rect 101404 480224 101456 480276
rect 561036 480224 561088 480276
rect 580172 480224 580224 480276
rect 2872 476076 2924 476128
rect 102968 476076 103020 476128
rect 567844 476076 567896 476128
rect 580172 476076 580224 476128
rect 561128 473356 561180 473408
rect 580172 473356 580224 473408
rect 2872 471996 2924 472048
rect 87604 471996 87656 472048
rect 128360 469820 128412 469872
rect 147680 469820 147732 469872
rect 2964 467848 3016 467900
rect 100208 467848 100260 467900
rect 3516 465060 3568 465112
rect 93216 465060 93268 465112
rect 573364 465060 573416 465112
rect 580172 465060 580224 465112
rect 3516 460912 3568 460964
rect 113824 460912 113876 460964
rect 556896 460912 556948 460964
rect 580080 460912 580132 460964
rect 3240 456764 3292 456816
rect 105544 456764 105596 456816
rect 119988 456764 120040 456816
rect 580080 456764 580132 456816
rect 3332 452616 3384 452668
rect 126244 452616 126296 452668
rect 3332 448536 3384 448588
rect 120816 448536 120868 448588
rect 563704 448536 563756 448588
rect 579712 448536 579764 448588
rect 3516 444388 3568 444440
rect 109132 444388 109184 444440
rect 570696 444388 570748 444440
rect 580172 444388 580224 444440
rect 3332 440240 3384 440292
rect 119344 440240 119396 440292
rect 572076 440240 572128 440292
rect 580172 440240 580224 440292
rect 3516 436092 3568 436144
rect 183652 436092 183704 436144
rect 567936 436092 567988 436144
rect 579620 436092 579672 436144
rect 3516 431944 3568 431996
rect 93400 431944 93452 431996
rect 563796 431944 563848 431996
rect 580172 431944 580224 431996
rect 563888 429156 563940 429208
rect 579988 429156 580040 429208
rect 2872 427796 2924 427848
rect 108580 427796 108632 427848
rect 577596 425076 577648 425128
rect 579620 425076 579672 425128
rect 3516 416780 3568 416832
rect 112536 416780 112588 416832
rect 3516 412632 3568 412684
rect 118056 412632 118108 412684
rect 572168 412632 572220 412684
rect 580172 412632 580224 412684
rect 3516 408484 3568 408536
rect 104992 408484 105044 408536
rect 149704 407736 149756 407788
rect 182272 407736 182324 407788
rect 552848 404336 552900 404388
rect 580172 404336 580224 404388
rect 3240 400188 3292 400240
rect 184940 400188 184992 400240
rect 191748 400188 191800 400240
rect 580172 400188 580224 400240
rect 3608 396040 3660 396092
rect 79416 396040 79468 396092
rect 569224 391960 569276 392012
rect 580172 391960 580224 392012
rect 2964 387812 3016 387864
rect 87696 387812 87748 387864
rect 121276 385024 121328 385076
rect 579804 385024 579856 385076
rect 3148 383664 3200 383716
rect 94780 383664 94832 383716
rect 196624 380876 196676 380928
rect 579988 380876 580040 380928
rect 3332 379516 3384 379568
rect 107016 379516 107068 379568
rect 3332 376728 3384 376780
rect 90640 376728 90692 376780
rect 569316 376728 569368 376780
rect 580172 376728 580224 376780
rect 3332 372580 3384 372632
rect 194600 372580 194652 372632
rect 556988 372580 557040 372632
rect 580172 372580 580224 372632
rect 3332 368500 3384 368552
rect 97540 368500 97592 368552
rect 559656 368500 559708 368552
rect 580172 368500 580224 368552
rect 3332 364488 3384 364540
rect 7564 364488 7616 364540
rect 191104 364352 191156 364404
rect 579620 364352 579672 364404
rect 3332 360204 3384 360256
rect 103060 360204 103112 360256
rect 561220 360204 561272 360256
rect 579620 360204 579672 360256
rect 3332 356056 3384 356108
rect 98920 356056 98972 356108
rect 192576 356056 192628 356108
rect 580172 356056 580224 356108
rect 563980 353268 564032 353320
rect 579620 353268 579672 353320
rect 3240 351908 3292 351960
rect 96068 351908 96120 351960
rect 194508 349120 194560 349172
rect 580172 349120 580224 349172
rect 3148 347760 3200 347812
rect 120908 347760 120960 347812
rect 558460 345040 558512 345092
rect 580172 345040 580224 345092
rect 3332 343612 3384 343664
rect 107108 343612 107160 343664
rect 575020 340892 575072 340944
rect 580172 340892 580224 340944
rect 3148 339464 3200 339516
rect 113916 339464 113968 339516
rect 128452 336744 128504 336796
rect 579988 336744 580040 336796
rect 171048 335996 171100 336048
rect 359464 335996 359516 336048
rect 3332 335316 3384 335368
rect 103152 335316 103204 335368
rect 3332 332596 3384 332648
rect 101496 332596 101548 332648
rect 572260 332596 572312 332648
rect 579988 332596 580040 332648
rect 3332 328448 3384 328500
rect 99012 328448 99064 328500
rect 3332 324300 3384 324352
rect 96160 324300 96212 324352
rect 3148 320152 3200 320204
rect 125692 320152 125744 320204
rect 575112 320152 575164 320204
rect 579620 320152 579672 320204
rect 3332 316004 3384 316056
rect 119436 316004 119488 316056
rect 566740 316004 566792 316056
rect 579620 316004 579672 316056
rect 577688 313284 577740 313336
rect 580632 313284 580684 313336
rect 555516 309136 555568 309188
rect 580172 309136 580224 309188
rect 3332 307776 3384 307828
rect 107200 307776 107252 307828
rect 572352 304988 572404 305040
rect 579620 304988 579672 305040
rect 3056 303628 3108 303680
rect 104624 303628 104676 303680
rect 577780 300840 577832 300892
rect 580632 300840 580684 300892
rect 3148 299480 3200 299532
rect 104072 299480 104124 299532
rect 180064 296692 180116 296744
rect 580172 296692 580224 296744
rect 3332 295332 3384 295384
rect 10324 295332 10376 295384
rect 569408 292544 569460 292596
rect 579988 292544 580040 292596
rect 3148 291184 3200 291236
rect 122104 291184 122156 291236
rect 561312 288396 561364 288448
rect 579988 288396 580040 288448
rect 3332 287036 3384 287088
rect 108672 287036 108724 287088
rect 3332 284316 3384 284368
rect 101588 284316 101640 284368
rect 3332 280168 3384 280220
rect 99104 280168 99156 280220
rect 558552 280168 558604 280220
rect 580172 280168 580224 280220
rect 13084 277992 13136 278044
rect 174544 277992 174596 278044
rect 564072 276020 564124 276072
rect 580172 276020 580224 276072
rect 124864 275272 124916 275324
rect 396080 275272 396132 275324
rect 14464 273912 14516 273964
rect 109224 273912 109276 273964
rect 109224 273232 109276 273284
rect 110236 273232 110288 273284
rect 133880 273232 133932 273284
rect 575204 273232 575256 273284
rect 580172 273232 580224 273284
rect 3148 271872 3200 271924
rect 145564 271872 145616 271924
rect 7564 271124 7616 271176
rect 165620 271124 165672 271176
rect 148968 269832 149020 269884
rect 288440 269832 288492 269884
rect 10324 269764 10376 269816
rect 161480 269764 161532 269816
rect 79416 268336 79468 268388
rect 156052 268336 156104 268388
rect 153108 267044 153160 267096
rect 199384 267044 199436 267096
rect 21364 266976 21416 267028
rect 115388 266976 115440 267028
rect 191656 266976 191708 267028
rect 440240 266976 440292 267028
rect 155684 266364 155736 266416
rect 190552 266364 190604 266416
rect 191656 266364 191708 266416
rect 145564 265820 145616 265872
rect 169760 265820 169812 265872
rect 155960 265752 156012 265804
rect 190460 265752 190512 265804
rect 151820 265684 151872 265736
rect 196072 265684 196124 265736
rect 67640 265616 67692 265668
rect 173072 265616 173124 265668
rect 179328 265140 179380 265192
rect 197544 265140 197596 265192
rect 174544 265072 174596 265124
rect 193496 265072 193548 265124
rect 162768 265004 162820 265056
rect 193312 265004 193364 265056
rect 196624 265004 196676 265056
rect 112536 264936 112588 264988
rect 115756 264936 115808 264988
rect 146760 264936 146812 264988
rect 161480 264936 161532 264988
rect 194784 264936 194836 264988
rect 566832 264936 566884 264988
rect 580172 264936 580224 264988
rect 146208 264256 146260 264308
rect 180064 264256 180116 264308
rect 34520 264188 34572 264240
rect 118700 264188 118752 264240
rect 115020 264052 115072 264104
rect 148968 264052 149020 264104
rect 115572 263984 115624 264036
rect 135444 263984 135496 264036
rect 112720 263916 112772 263968
rect 138664 263916 138716 263968
rect 117688 263848 117740 263900
rect 145380 263848 145432 263900
rect 192576 264188 192628 264240
rect 195060 264188 195112 264240
rect 215944 264188 215996 264240
rect 117136 263780 117188 263832
rect 146208 263780 146260 263832
rect 121000 263712 121052 263764
rect 152004 263712 152056 263764
rect 153108 263712 153160 263764
rect 118700 263644 118752 263696
rect 119068 263644 119120 263696
rect 152556 263644 152608 263696
rect 185492 263644 185544 263696
rect 194692 263644 194744 263696
rect 195060 263644 195112 263696
rect 3332 263576 3384 263628
rect 107292 263576 107344 263628
rect 113916 263576 113968 263628
rect 115572 263576 115624 263628
rect 159824 263576 159876 263628
rect 194968 263576 195020 263628
rect 200764 263576 200816 263628
rect 113916 263168 113968 263220
rect 143540 263168 143592 263220
rect 160652 263168 160704 263220
rect 193404 263168 193456 263220
rect 111616 263100 111668 263152
rect 141792 263100 141844 263152
rect 169668 263100 169720 263152
rect 198924 263100 198976 263152
rect 112536 263032 112588 263084
rect 131304 263032 131356 263084
rect 126244 262964 126296 263016
rect 127900 262964 127952 263016
rect 157248 263032 157300 263084
rect 182180 263032 182232 263084
rect 183468 263032 183520 263084
rect 198740 263032 198792 263084
rect 285680 263032 285732 263084
rect 327080 262964 327132 263016
rect 122104 262896 122156 262948
rect 188160 262896 188212 262948
rect 38660 262828 38712 262880
rect 117044 262760 117096 262812
rect 150072 262760 150124 262812
rect 183468 262828 183520 262880
rect 192576 262828 192628 262880
rect 164424 262760 164476 262812
rect 197820 262760 197872 262812
rect 114284 262692 114336 262744
rect 133512 262692 133564 262744
rect 183468 262692 183520 262744
rect 198372 262692 198424 262744
rect 444380 262896 444432 262948
rect 198924 262828 198976 262880
rect 199568 262828 199620 262880
rect 467840 262828 467892 262880
rect 116952 262624 117004 262676
rect 140136 262624 140188 262676
rect 177212 262624 177264 262676
rect 198464 262624 198516 262676
rect 112904 262556 112956 262608
rect 139400 262556 139452 262608
rect 165528 262556 165580 262608
rect 192116 262556 192168 262608
rect 119896 262488 119948 262540
rect 147680 262488 147732 262540
rect 172244 262488 172296 262540
rect 198740 262488 198792 262540
rect 199200 262488 199252 262540
rect 114100 262420 114152 262472
rect 142620 262420 142672 262472
rect 168932 262420 168984 262472
rect 196624 262420 196676 262472
rect 115296 262352 115348 262404
rect 126980 262352 127032 262404
rect 135260 262352 135312 262404
rect 179880 262352 179932 262404
rect 190644 262352 190696 262404
rect 127716 262284 127768 262336
rect 116860 262216 116912 262268
rect 125232 262216 125284 262268
rect 132776 262284 132828 262336
rect 135444 262284 135496 262336
rect 137652 262284 137704 262336
rect 187608 262284 187660 262336
rect 211160 262284 211212 262336
rect 119712 262148 119764 262200
rect 127900 262216 127952 262268
rect 136824 262216 136876 262268
rect 177948 262216 178000 262268
rect 192208 262216 192260 262268
rect 53104 260992 53156 261044
rect 179880 260992 179932 261044
rect 182088 260992 182140 261044
rect 197452 260992 197504 261044
rect 114376 260924 114428 260976
rect 189080 260924 189132 260976
rect 176384 260856 176436 260908
rect 192760 260856 192812 260908
rect 577872 260856 577924 260908
rect 580724 260856 580776 260908
rect 118608 260788 118660 260840
rect 122840 260788 122892 260840
rect 114008 260176 114060 260228
rect 111248 260108 111300 260160
rect 126244 260176 126296 260228
rect 128452 260176 128504 260228
rect 129694 260176 129746 260228
rect 158168 260312 158220 260364
rect 191196 260312 191248 260364
rect 156052 260244 156104 260296
rect 190736 260244 190788 260296
rect 144598 260176 144650 260228
rect 161158 260176 161210 260228
rect 196440 260176 196492 260228
rect 116676 260040 116728 260092
rect 127210 260108 127262 260160
rect 117872 259972 117924 260024
rect 158674 260108 158726 260160
rect 193680 260108 193732 260160
rect 124036 259904 124088 259956
rect 149566 260040 149618 260092
rect 182686 260040 182738 260092
rect 195060 260040 195112 260092
rect 181352 259972 181404 260024
rect 197912 259972 197964 260024
rect 168104 259904 168156 259956
rect 192668 259904 192720 259956
rect 112628 259836 112680 259888
rect 126060 259836 126112 259888
rect 169760 259836 169812 259888
rect 170956 259836 171008 259888
rect 196256 259836 196308 259888
rect 112352 259768 112404 259820
rect 128360 259768 128412 259820
rect 166448 259768 166500 259820
rect 196348 259768 196400 259820
rect 111156 259700 111208 259752
rect 131120 259700 131172 259752
rect 131856 259700 131908 259752
rect 163964 259700 164016 259752
rect 193772 259700 193824 259752
rect 113640 259632 113692 259684
rect 135996 259632 136048 259684
rect 184664 259632 184716 259684
rect 196164 259632 196216 259684
rect 115112 259564 115164 259616
rect 123576 259564 123628 259616
rect 124864 259564 124916 259616
rect 178868 259564 178920 259616
rect 198924 259564 198976 259616
rect 118332 259496 118384 259548
rect 150900 259496 150952 259548
rect 175372 259496 175424 259548
rect 189632 259496 189684 259548
rect 3056 259428 3108 259480
rect 101680 259428 101732 259480
rect 119252 259428 119304 259480
rect 124404 259428 124456 259480
rect 173808 259428 173860 259480
rect 194876 259428 194928 259480
rect 116768 259292 116820 259344
rect 124036 259292 124088 259344
rect 120080 259224 120132 259276
rect 121276 259224 121328 259276
rect 120448 258748 120500 258800
rect 121000 258748 121052 258800
rect 3148 255280 3200 255332
rect 117412 255280 117464 255332
rect 120172 253376 120224 253428
rect 120080 253172 120132 253224
rect 192760 252560 192812 252612
rect 196532 252560 196584 252612
rect 579804 252560 579856 252612
rect 3148 251200 3200 251252
rect 119528 251200 119580 251252
rect 191288 248412 191340 248464
rect 579804 248412 579856 248464
rect 3332 247052 3384 247104
rect 96528 247052 96580 247104
rect 190092 244264 190144 244316
rect 580172 244264 580224 244316
rect 3148 242904 3200 242956
rect 119620 242904 119672 242956
rect 3332 240048 3384 240100
rect 53104 240048 53156 240100
rect 191656 237396 191708 237448
rect 580172 237396 580224 237448
rect 3332 235968 3384 236020
rect 109684 235968 109736 236020
rect 3332 231820 3384 231872
rect 112996 231820 113048 231872
rect 3332 227740 3384 227792
rect 92480 227740 92532 227792
rect 3332 223592 3384 223644
rect 120632 223592 120684 223644
rect 208400 220804 208452 220856
rect 580172 220804 580224 220856
rect 3240 220736 3292 220788
rect 114376 220736 114428 220788
rect 191196 217268 191248 217320
rect 580172 217268 580224 217320
rect 3332 215296 3384 215348
rect 96436 215296 96488 215348
rect 119160 215296 119212 215348
rect 190460 208904 190512 208956
rect 190828 208904 190880 208956
rect 202788 206252 202840 206304
rect 580632 206252 580684 206304
rect 191380 205640 191432 205692
rect 201684 205640 201736 205692
rect 202788 205640 202840 205692
rect 576400 205572 576452 205624
rect 579988 205572 580040 205624
rect 115940 202784 115992 202836
rect 116584 202784 116636 202836
rect 96988 201560 97040 201612
rect 116584 201560 116636 201612
rect 96344 201492 96396 201544
rect 117412 201492 117464 201544
rect 117780 201492 117832 201544
rect 211068 200880 211120 200932
rect 474740 200880 474792 200932
rect 191748 200812 191800 200864
rect 204536 200812 204588 200864
rect 221004 200812 221056 200864
rect 531320 200812 531372 200864
rect 3516 200744 3568 200796
rect 92480 200744 92532 200796
rect 113824 200744 113876 200796
rect 115204 200676 115256 200728
rect 119620 200608 119672 200660
rect 131856 200608 131908 200660
rect 119436 200200 119488 200252
rect 122840 200200 122892 200252
rect 92480 200132 92532 200184
rect 93676 200132 93728 200184
rect 132040 200336 132092 200388
rect 124864 200200 124916 200252
rect 131948 199928 132000 199980
rect 128544 199860 128596 199912
rect 131764 199860 131816 199912
rect 132224 199860 132276 199912
rect 132822 199860 132874 199912
rect 133926 199860 133978 199912
rect 117964 199792 118016 199844
rect 124864 199792 124916 199844
rect 124956 199792 125008 199844
rect 133282 199792 133334 199844
rect 133650 199792 133702 199844
rect 133742 199792 133794 199844
rect 110328 199724 110380 199776
rect 88984 199588 89036 199640
rect 108120 199588 108172 199640
rect 132132 199724 132184 199776
rect 132500 199724 132552 199776
rect 133006 199724 133058 199776
rect 133098 199724 133150 199776
rect 125508 199656 125560 199708
rect 131672 199656 131724 199708
rect 75920 199520 75972 199572
rect 108212 199520 108264 199572
rect 118056 199520 118108 199572
rect 124312 199520 124364 199572
rect 125508 199520 125560 199572
rect 71780 199452 71832 199504
rect 132224 199588 132276 199640
rect 132776 199588 132828 199640
rect 131764 199520 131816 199572
rect 133374 199724 133426 199776
rect 133236 199588 133288 199640
rect 133604 199588 133656 199640
rect 133696 199588 133748 199640
rect 134294 199860 134346 199912
rect 134478 199860 134530 199912
rect 134570 199860 134622 199912
rect 134340 199656 134392 199708
rect 134432 199656 134484 199708
rect 134524 199656 134576 199708
rect 134064 199588 134116 199640
rect 134248 199588 134300 199640
rect 134846 199860 134898 199912
rect 135122 199860 135174 199912
rect 135306 199860 135358 199912
rect 135398 199860 135450 199912
rect 135490 199860 135542 199912
rect 135674 199860 135726 199912
rect 135766 199860 135818 199912
rect 136042 199860 136094 199912
rect 136410 199860 136462 199912
rect 136594 199860 136646 199912
rect 136686 199860 136738 199912
rect 136778 199860 136830 199912
rect 136870 199860 136922 199912
rect 137146 199860 137198 199912
rect 134800 199724 134852 199776
rect 134938 199724 134990 199776
rect 134892 199588 134944 199640
rect 134340 199520 134392 199572
rect 134984 199520 135036 199572
rect 135352 199724 135404 199776
rect 135444 199656 135496 199708
rect 135950 199792 136002 199844
rect 135720 199656 135772 199708
rect 135996 199656 136048 199708
rect 135904 199588 135956 199640
rect 136640 199724 136692 199776
rect 136456 199588 136508 199640
rect 135260 199520 135312 199572
rect 135628 199520 135680 199572
rect 135812 199520 135864 199572
rect 136824 199520 136876 199572
rect 136916 199520 136968 199572
rect 137008 199520 137060 199572
rect 137606 199860 137658 199912
rect 137790 199860 137842 199912
rect 137974 199860 138026 199912
rect 138618 199860 138670 199912
rect 138710 199860 138762 199912
rect 139078 199860 139130 199912
rect 137514 199792 137566 199844
rect 137560 199656 137612 199708
rect 137376 199588 137428 199640
rect 137928 199724 137980 199776
rect 138158 199724 138210 199776
rect 138342 199724 138394 199776
rect 137836 199656 137888 199708
rect 138894 199792 138946 199844
rect 138664 199724 138716 199776
rect 138756 199656 138808 199708
rect 138940 199656 138992 199708
rect 139170 199792 139222 199844
rect 139354 199792 139406 199844
rect 139124 199656 139176 199708
rect 139216 199656 139268 199708
rect 138848 199588 138900 199640
rect 139032 199588 139084 199640
rect 139308 199588 139360 199640
rect 139998 199860 140050 199912
rect 139630 199792 139682 199844
rect 140182 199792 140234 199844
rect 139584 199656 139636 199708
rect 139952 199656 140004 199708
rect 140136 199588 140188 199640
rect 140826 199860 140878 199912
rect 141102 199860 141154 199912
rect 141378 199860 141430 199912
rect 140458 199792 140510 199844
rect 140504 199656 140556 199708
rect 137744 199520 137796 199572
rect 138388 199520 138440 199572
rect 140320 199520 140372 199572
rect 3424 199384 3476 199436
rect 108764 199384 108816 199436
rect 119344 199384 119396 199436
rect 126796 199384 126848 199436
rect 131212 199384 131264 199436
rect 132224 199384 132276 199436
rect 140228 199452 140280 199504
rect 142022 199860 142074 199912
rect 141470 199792 141522 199844
rect 141746 199792 141798 199844
rect 141930 199792 141982 199844
rect 140688 199520 140740 199572
rect 140596 199452 140648 199504
rect 142574 199860 142626 199912
rect 142666 199860 142718 199912
rect 142758 199860 142810 199912
rect 142528 199656 142580 199708
rect 143310 199860 143362 199912
rect 143586 199860 143638 199912
rect 142942 199792 142994 199844
rect 142160 199588 142212 199640
rect 142344 199588 142396 199640
rect 142804 199588 142856 199640
rect 142620 199520 142672 199572
rect 142712 199520 142764 199572
rect 143126 199724 143178 199776
rect 142988 199656 143040 199708
rect 143080 199588 143132 199640
rect 143172 199588 143224 199640
rect 143494 199724 143546 199776
rect 143402 199656 143454 199708
rect 141424 199452 141476 199504
rect 141700 199452 141752 199504
rect 141884 199452 141936 199504
rect 143264 199452 143316 199504
rect 143356 199452 143408 199504
rect 143540 199588 143592 199640
rect 144138 199860 144190 199912
rect 144414 199860 144466 199912
rect 144874 199860 144926 199912
rect 144966 199860 145018 199912
rect 145150 199860 145202 199912
rect 145242 199860 145294 199912
rect 145334 199860 145386 199912
rect 145426 199860 145478 199912
rect 145518 199860 145570 199912
rect 145702 199860 145754 199912
rect 145886 199860 145938 199912
rect 145978 199860 146030 199912
rect 146070 199860 146122 199912
rect 146254 199860 146306 199912
rect 146346 199860 146398 199912
rect 146438 199860 146490 199912
rect 146530 199860 146582 199912
rect 143770 199792 143822 199844
rect 143862 199724 143914 199776
rect 143908 199520 143960 199572
rect 144368 199724 144420 199776
rect 144276 199588 144328 199640
rect 144368 199520 144420 199572
rect 144460 199520 144512 199572
rect 144782 199792 144834 199844
rect 144828 199656 144880 199708
rect 144920 199656 144972 199708
rect 145012 199520 145064 199572
rect 143816 199452 143868 199504
rect 145196 199724 145248 199776
rect 145380 199588 145432 199640
rect 145288 199520 145340 199572
rect 145564 199656 145616 199708
rect 145656 199656 145708 199708
rect 146208 199724 146260 199776
rect 146300 199724 146352 199776
rect 146392 199724 146444 199776
rect 146024 199656 146076 199708
rect 145840 199588 145892 199640
rect 145932 199588 145984 199640
rect 146484 199520 146536 199572
rect 147082 199860 147134 199912
rect 147542 199860 147594 199912
rect 147726 199860 147778 199912
rect 147910 199860 147962 199912
rect 148002 199860 148054 199912
rect 148370 199860 148422 199912
rect 146760 199520 146812 199572
rect 146852 199452 146904 199504
rect 147772 199724 147824 199776
rect 147680 199588 147732 199640
rect 148738 199860 148790 199912
rect 149014 199860 149066 199912
rect 149750 199860 149802 199912
rect 148140 199588 148192 199640
rect 148416 199588 148468 199640
rect 148600 199588 148652 199640
rect 148876 199588 148928 199640
rect 149290 199792 149342 199844
rect 149382 199792 149434 199844
rect 149428 199656 149480 199708
rect 149336 199588 149388 199640
rect 149612 199520 149664 199572
rect 150026 199724 150078 199776
rect 147404 199452 147456 199504
rect 149336 199452 149388 199504
rect 149888 199452 149940 199504
rect 149980 199452 150032 199504
rect 150486 199792 150538 199844
rect 150348 199520 150400 199572
rect 150440 199520 150492 199572
rect 151038 199792 151090 199844
rect 150992 199588 151044 199640
rect 151682 199860 151734 199912
rect 151406 199792 151458 199844
rect 151498 199792 151550 199844
rect 147956 199384 148008 199436
rect 148508 199384 148560 199436
rect 150532 199384 150584 199436
rect 150716 199384 150768 199436
rect 119436 199316 119488 199368
rect 121920 199316 121972 199368
rect 148968 199316 149020 199368
rect 140504 199248 140556 199300
rect 144092 199248 144144 199300
rect 150348 199316 150400 199368
rect 151958 199860 152010 199912
rect 152234 199860 152286 199912
rect 152326 199860 152378 199912
rect 152510 199860 152562 199912
rect 152602 199860 152654 199912
rect 152694 199860 152746 199912
rect 152878 199860 152930 199912
rect 151452 199656 151504 199708
rect 151728 199588 151780 199640
rect 152464 199724 152516 199776
rect 152280 199656 152332 199708
rect 152372 199588 152424 199640
rect 152556 199588 152608 199640
rect 151912 199520 151964 199572
rect 152832 199588 152884 199640
rect 178224 200676 178276 200728
rect 580724 200744 580776 200796
rect 153430 199860 153482 199912
rect 153338 199792 153390 199844
rect 153614 199860 153666 199912
rect 153706 199860 153758 199912
rect 153798 199860 153850 199912
rect 153890 199860 153942 199912
rect 153752 199724 153804 199776
rect 153568 199656 153620 199708
rect 153292 199588 153344 199640
rect 153476 199588 153528 199640
rect 153384 199520 153436 199572
rect 153844 199588 153896 199640
rect 154074 199860 154126 199912
rect 153936 199520 153988 199572
rect 154350 199860 154402 199912
rect 154442 199860 154494 199912
rect 154534 199860 154586 199912
rect 154626 199860 154678 199912
rect 154994 199860 155046 199912
rect 154304 199656 154356 199708
rect 154488 199656 154540 199708
rect 154580 199656 154632 199708
rect 154856 199588 154908 199640
rect 154764 199520 154816 199572
rect 151360 199452 151412 199504
rect 152004 199452 152056 199504
rect 152372 199452 152424 199504
rect 153660 199452 153712 199504
rect 152648 199384 152700 199436
rect 155270 199860 155322 199912
rect 155362 199860 155414 199912
rect 155454 199860 155506 199912
rect 155546 199860 155598 199912
rect 155638 199860 155690 199912
rect 155316 199724 155368 199776
rect 155408 199724 155460 199776
rect 155592 199656 155644 199708
rect 155500 199588 155552 199640
rect 155914 199860 155966 199912
rect 155868 199520 155920 199572
rect 156466 199860 156518 199912
rect 156558 199860 156610 199912
rect 156742 199860 156794 199912
rect 156512 199724 156564 199776
rect 157110 199860 157162 199912
rect 157202 199860 157254 199912
rect 157386 199860 157438 199912
rect 157570 199860 157622 199912
rect 157754 199860 157806 199912
rect 157156 199656 157208 199708
rect 156788 199588 156840 199640
rect 156972 199588 157024 199640
rect 157248 199588 157300 199640
rect 157938 199860 157990 199912
rect 158030 199860 158082 199912
rect 158122 199860 158174 199912
rect 158214 199860 158266 199912
rect 158306 199860 158358 199912
rect 158490 199860 158542 199912
rect 158674 199860 158726 199912
rect 157800 199724 157852 199776
rect 157892 199724 157944 199776
rect 158076 199724 158128 199776
rect 157984 199656 158036 199708
rect 157616 199588 157668 199640
rect 158168 199588 158220 199640
rect 157432 199520 157484 199572
rect 158260 199520 158312 199572
rect 156420 199384 156472 199436
rect 158950 199860 159002 199912
rect 159134 199860 159186 199912
rect 159226 199860 159278 199912
rect 159686 199860 159738 199912
rect 159870 199860 159922 199912
rect 160054 199860 160106 199912
rect 160698 199860 160750 199912
rect 160790 199860 160842 199912
rect 160882 199860 160934 199912
rect 161066 199860 161118 199912
rect 161158 199860 161210 199912
rect 161434 199860 161486 199912
rect 158996 199724 159048 199776
rect 159088 199724 159140 199776
rect 159364 199588 159416 199640
rect 158812 199384 158864 199436
rect 152372 199316 152424 199368
rect 153752 199316 153804 199368
rect 132224 199180 132276 199232
rect 153108 199180 153160 199232
rect 119528 199112 119580 199164
rect 122932 199112 122984 199164
rect 144000 199112 144052 199164
rect 145656 199112 145708 199164
rect 147864 199112 147916 199164
rect 147956 199112 148008 199164
rect 119160 199044 119212 199096
rect 148508 199044 148560 199096
rect 108120 198976 108172 199028
rect 108948 198976 109000 199028
rect 142160 198976 142212 199028
rect 108212 198908 108264 198960
rect 108856 198908 108908 198960
rect 142252 198908 142304 198960
rect 149520 199112 149572 199164
rect 149888 199112 149940 199164
rect 154396 199180 154448 199232
rect 159548 199384 159600 199436
rect 160330 199792 160382 199844
rect 160422 199792 160474 199844
rect 159824 199588 159876 199640
rect 160284 199588 160336 199640
rect 160744 199724 160796 199776
rect 161342 199792 161394 199844
rect 161204 199724 161256 199776
rect 161112 199656 161164 199708
rect 161296 199656 161348 199708
rect 161618 199792 161670 199844
rect 161388 199588 161440 199640
rect 160836 199520 160888 199572
rect 160376 199384 160428 199436
rect 160192 199316 160244 199368
rect 161802 199860 161854 199912
rect 161664 199384 161716 199436
rect 160928 199316 160980 199368
rect 162170 199860 162222 199912
rect 162354 199860 162406 199912
rect 162446 199860 162498 199912
rect 162538 199860 162590 199912
rect 162400 199724 162452 199776
rect 162630 199792 162682 199844
rect 162492 199656 162544 199708
rect 162584 199656 162636 199708
rect 162216 199588 162268 199640
rect 162124 199520 162176 199572
rect 177856 200608 177908 200660
rect 178040 200608 178092 200660
rect 181904 200676 181956 200728
rect 182824 200676 182876 200728
rect 428464 200676 428516 200728
rect 191288 200608 191340 200660
rect 177764 200540 177816 200592
rect 179144 200540 179196 200592
rect 177948 200472 178000 200524
rect 162998 199860 163050 199912
rect 163090 199860 163142 199912
rect 163182 199860 163234 199912
rect 163366 199860 163418 199912
rect 163458 199860 163510 199912
rect 163044 199656 163096 199708
rect 163412 199656 163464 199708
rect 163320 199588 163372 199640
rect 163136 199520 163188 199572
rect 163734 199860 163786 199912
rect 164010 199860 164062 199912
rect 164286 199860 164338 199912
rect 163964 199724 164016 199776
rect 163688 199520 163740 199572
rect 164240 199656 164292 199708
rect 164240 199452 164292 199504
rect 164470 199860 164522 199912
rect 164654 199860 164706 199912
rect 164930 199860 164982 199912
rect 165206 199860 165258 199912
rect 164516 199724 164568 199776
rect 165482 199860 165534 199912
rect 165758 199860 165810 199912
rect 165942 199860 165994 199912
rect 166034 199860 166086 199912
rect 166218 199860 166270 199912
rect 166310 199860 166362 199912
rect 166402 199860 166454 199912
rect 166586 199860 166638 199912
rect 166862 199860 166914 199912
rect 166954 199860 167006 199912
rect 167138 199860 167190 199912
rect 167690 199860 167742 199912
rect 168058 199860 168110 199912
rect 168150 199860 168202 199912
rect 168334 199860 168386 199912
rect 168426 199860 168478 199912
rect 168518 199860 168570 199912
rect 168610 199860 168662 199912
rect 168886 199860 168938 199912
rect 168978 199860 169030 199912
rect 169070 199860 169122 199912
rect 169622 199860 169674 199912
rect 169806 199860 169858 199912
rect 169898 199860 169950 199912
rect 169990 199860 170042 199912
rect 170082 199860 170134 199912
rect 170174 199860 170226 199912
rect 165068 199588 165120 199640
rect 165160 199588 165212 199640
rect 165252 199588 165304 199640
rect 165804 199588 165856 199640
rect 166264 199724 166316 199776
rect 166356 199724 166408 199776
rect 166172 199588 166224 199640
rect 166540 199588 166592 199640
rect 166908 199724 166960 199776
rect 167598 199792 167650 199844
rect 167552 199588 167604 199640
rect 168196 199724 168248 199776
rect 168288 199724 168340 199776
rect 168012 199588 168064 199640
rect 166724 199520 166776 199572
rect 166816 199520 166868 199572
rect 167368 199520 167420 199572
rect 167736 199520 167788 199572
rect 168472 199656 168524 199708
rect 168656 199588 168708 199640
rect 168748 199588 168800 199640
rect 168564 199520 168616 199572
rect 168840 199520 168892 199572
rect 169760 199724 169812 199776
rect 169668 199656 169720 199708
rect 169852 199656 169904 199708
rect 169576 199588 169628 199640
rect 170128 199724 170180 199776
rect 170634 199860 170686 199912
rect 170818 199860 170870 199912
rect 171002 199860 171054 199912
rect 171094 199860 171146 199912
rect 171186 199860 171238 199912
rect 170772 199724 170824 199776
rect 171048 199724 171100 199776
rect 171140 199724 171192 199776
rect 164792 199452 164844 199504
rect 165988 199452 166040 199504
rect 169116 199452 169168 199504
rect 170404 199452 170456 199504
rect 171324 199452 171376 199504
rect 171738 199860 171790 199912
rect 171922 199860 171974 199912
rect 172106 199860 172158 199912
rect 172290 199860 172342 199912
rect 171784 199588 171836 199640
rect 172060 199588 172112 199640
rect 172520 199452 172572 199504
rect 162032 199384 162084 199436
rect 162308 199384 162360 199436
rect 162860 199384 162912 199436
rect 165896 199384 165948 199436
rect 167920 199384 167972 199436
rect 168380 199384 168432 199436
rect 161204 199248 161256 199300
rect 161480 199248 161532 199300
rect 167092 199316 167144 199368
rect 167368 199316 167420 199368
rect 167736 199316 167788 199368
rect 170220 199316 170272 199368
rect 170588 199316 170640 199368
rect 171600 199384 171652 199436
rect 172842 199860 172894 199912
rect 172934 199860 172986 199912
rect 173026 199860 173078 199912
rect 173302 199860 173354 199912
rect 173394 199860 173446 199912
rect 173486 199860 173538 199912
rect 173578 199860 173630 199912
rect 173670 199860 173722 199912
rect 173762 199860 173814 199912
rect 173854 199860 173906 199912
rect 172796 199724 172848 199776
rect 173256 199724 173308 199776
rect 173348 199724 173400 199776
rect 173532 199724 173584 199776
rect 173624 199724 173676 199776
rect 173716 199520 173768 199572
rect 174590 199860 174642 199912
rect 174636 199588 174688 199640
rect 178592 200404 178644 200456
rect 191748 200540 191800 200592
rect 194508 200404 194560 200456
rect 200120 200404 200172 200456
rect 190460 200336 190512 200388
rect 191656 200336 191708 200388
rect 214104 200336 214156 200388
rect 177856 200268 177908 200320
rect 179052 200268 179104 200320
rect 209964 200268 210016 200320
rect 211068 200268 211120 200320
rect 221004 200200 221056 200252
rect 177948 200132 178000 200184
rect 188988 200132 189040 200184
rect 580172 200132 580224 200184
rect 179052 200064 179104 200116
rect 179236 200064 179288 200116
rect 182916 200064 182968 200116
rect 174958 199860 175010 199912
rect 175510 199860 175562 199912
rect 175602 199860 175654 199912
rect 175694 199860 175746 199912
rect 175786 199860 175838 199912
rect 175648 199656 175700 199708
rect 175556 199588 175608 199640
rect 177948 199996 178000 200048
rect 177764 199928 177816 199980
rect 181904 199928 181956 199980
rect 176062 199860 176114 199912
rect 176430 199860 176482 199912
rect 176522 199860 176574 199912
rect 176982 199860 177034 199912
rect 177258 199860 177310 199912
rect 177442 199860 177494 199912
rect 181812 199860 181864 199912
rect 176154 199792 176206 199844
rect 176108 199656 176160 199708
rect 172980 199452 173032 199504
rect 173900 199452 173952 199504
rect 176108 199452 176160 199504
rect 174452 199384 174504 199436
rect 172980 199316 173032 199368
rect 174912 199248 174964 199300
rect 177028 199724 177080 199776
rect 177948 199724 178000 199776
rect 176844 199588 176896 199640
rect 177304 199588 177356 199640
rect 179512 199588 179564 199640
rect 180340 199588 180392 199640
rect 176660 199520 176712 199572
rect 180984 199724 181036 199776
rect 303620 199724 303672 199776
rect 180708 199656 180760 199708
rect 191104 199656 191156 199708
rect 218428 199656 218480 199708
rect 402980 199656 403032 199708
rect 180524 199588 180576 199640
rect 184940 199588 184992 199640
rect 186228 199588 186280 199640
rect 448520 199588 448572 199640
rect 528560 199520 528612 199572
rect 176844 199452 176896 199504
rect 539600 199452 539652 199504
rect 176384 199384 176436 199436
rect 176476 199384 176528 199436
rect 177304 199384 177356 199436
rect 177672 199384 177724 199436
rect 582472 199384 582524 199436
rect 179236 199316 179288 199368
rect 176384 199248 176436 199300
rect 160652 199180 160704 199232
rect 161020 199112 161072 199164
rect 161480 199112 161532 199164
rect 161572 199112 161624 199164
rect 162124 199112 162176 199164
rect 170956 199180 171008 199232
rect 192484 199248 192536 199300
rect 177212 199180 177264 199232
rect 185400 199180 185452 199232
rect 184940 199112 184992 199164
rect 179696 199044 179748 199096
rect 180708 199044 180760 199096
rect 165436 198976 165488 199028
rect 156880 198908 156932 198960
rect 156972 198908 157024 198960
rect 163688 198908 163740 198960
rect 165344 198908 165396 198960
rect 190460 198976 190512 199028
rect 167092 198908 167144 198960
rect 188896 198908 188948 198960
rect 190092 198908 190144 198960
rect 106004 198840 106056 198892
rect 120724 198840 120776 198892
rect 121000 198840 121052 198892
rect 3516 198772 3568 198824
rect 119436 198772 119488 198824
rect 120816 198772 120868 198824
rect 124220 198772 124272 198824
rect 142068 198772 142120 198824
rect 117964 198704 118016 198756
rect 118700 198704 118752 198756
rect 120908 198704 120960 198756
rect 131304 198704 131356 198756
rect 132408 198704 132460 198756
rect 132500 198704 132552 198756
rect 137008 198704 137060 198756
rect 120724 198636 120776 198688
rect 133052 198636 133104 198688
rect 126888 198568 126940 198620
rect 130936 198568 130988 198620
rect 151268 198840 151320 198892
rect 154580 198840 154632 198892
rect 160928 198840 160980 198892
rect 166540 198840 166592 198892
rect 167920 198840 167972 198892
rect 194508 198840 194560 198892
rect 146392 198772 146444 198824
rect 146852 198772 146904 198824
rect 149428 198772 149480 198824
rect 161848 198772 161900 198824
rect 165344 198772 165396 198824
rect 165436 198772 165488 198824
rect 170956 198772 171008 198824
rect 171048 198772 171100 198824
rect 218060 198772 218112 198824
rect 218428 198772 218480 198824
rect 147680 198704 147732 198756
rect 153108 198704 153160 198756
rect 153844 198704 153896 198756
rect 154028 198704 154080 198756
rect 157800 198704 157852 198756
rect 158444 198704 158496 198756
rect 148968 198636 149020 198688
rect 154396 198636 154448 198688
rect 160744 198636 160796 198688
rect 165620 198636 165672 198688
rect 149428 198568 149480 198620
rect 149888 198568 149940 198620
rect 176476 198704 176528 198756
rect 176936 198704 176988 198756
rect 177120 198704 177172 198756
rect 182916 198704 182968 198756
rect 185584 198704 185636 198756
rect 189724 198704 189776 198756
rect 168472 198636 168524 198688
rect 168748 198636 168800 198688
rect 169300 198636 169352 198688
rect 194600 198636 194652 198688
rect 172520 198568 172572 198620
rect 177488 198568 177540 198620
rect 129188 198500 129240 198552
rect 140964 198500 141016 198552
rect 142252 198500 142304 198552
rect 147036 198500 147088 198552
rect 151452 198500 151504 198552
rect 125508 198432 125560 198484
rect 138020 198432 138072 198484
rect 153016 198432 153068 198484
rect 161020 198432 161072 198484
rect 163228 198432 163280 198484
rect 128176 198364 128228 198416
rect 141240 198364 141292 198416
rect 151084 198364 151136 198416
rect 154856 198364 154908 198416
rect 159824 198364 159876 198416
rect 166540 198364 166592 198416
rect 166908 198364 166960 198416
rect 167736 198364 167788 198416
rect 169760 198432 169812 198484
rect 170036 198432 170088 198484
rect 170680 198500 170732 198552
rect 171692 198500 171744 198552
rect 171968 198500 172020 198552
rect 190828 198568 190880 198620
rect 191748 198568 191800 198620
rect 185400 198500 185452 198552
rect 191380 198500 191432 198552
rect 172428 198432 172480 198484
rect 172796 198432 172848 198484
rect 173072 198432 173124 198484
rect 175556 198432 175608 198484
rect 175924 198432 175976 198484
rect 176016 198432 176068 198484
rect 176660 198432 176712 198484
rect 176752 198432 176804 198484
rect 189540 198432 189592 198484
rect 129648 198296 129700 198348
rect 140872 198296 140924 198348
rect 142896 198296 142948 198348
rect 143908 198296 143960 198348
rect 163872 198296 163924 198348
rect 165620 198296 165672 198348
rect 166724 198296 166776 198348
rect 172520 198296 172572 198348
rect 126520 198228 126572 198280
rect 134156 198228 134208 198280
rect 137100 198228 137152 198280
rect 137652 198228 137704 198280
rect 140964 198228 141016 198280
rect 141884 198228 141936 198280
rect 158168 198228 158220 198280
rect 159456 198228 159508 198280
rect 168564 198228 168616 198280
rect 171784 198228 171836 198280
rect 172428 198228 172480 198280
rect 176016 198296 176068 198348
rect 177396 198296 177448 198348
rect 173072 198228 173124 198280
rect 177764 198228 177816 198280
rect 193220 198228 193272 198280
rect 204352 198228 204404 198280
rect 100668 198160 100720 198212
rect 129740 198160 129792 198212
rect 137284 198160 137336 198212
rect 139676 198160 139728 198212
rect 140044 198160 140096 198212
rect 140320 198160 140372 198212
rect 142344 198160 142396 198212
rect 143448 198160 143500 198212
rect 159824 198160 159876 198212
rect 160928 198160 160980 198212
rect 161296 198160 161348 198212
rect 163688 198160 163740 198212
rect 166908 198160 166960 198212
rect 180800 198160 180852 198212
rect 181076 198160 181128 198212
rect 196072 198160 196124 198212
rect 201592 198160 201644 198212
rect 114468 198092 114520 198144
rect 128452 198092 128504 198144
rect 129648 198092 129700 198144
rect 141884 198092 141936 198144
rect 150808 198092 150860 198144
rect 159456 198092 159508 198144
rect 159732 198092 159784 198144
rect 164700 198092 164752 198144
rect 184940 198092 184992 198144
rect 194600 198092 194652 198144
rect 212540 198092 212592 198144
rect 100576 198024 100628 198076
rect 131948 198024 132000 198076
rect 132960 198024 133012 198076
rect 133236 198024 133288 198076
rect 62764 197956 62816 198008
rect 99196 197956 99248 198008
rect 133512 197956 133564 198008
rect 139860 198024 139912 198076
rect 140688 198024 140740 198076
rect 141700 198024 141752 198076
rect 144736 198024 144788 198076
rect 145012 198024 145064 198076
rect 156880 198024 156932 198076
rect 180156 198024 180208 198076
rect 191748 198024 191800 198076
rect 211436 198024 211488 198076
rect 127992 197888 128044 197940
rect 131764 197888 131816 197940
rect 127808 197820 127860 197872
rect 135352 197888 135404 197940
rect 138388 197956 138440 198008
rect 139308 197956 139360 198008
rect 139952 197956 140004 198008
rect 141056 197956 141108 198008
rect 142068 197956 142120 198008
rect 139768 197888 139820 197940
rect 140780 197888 140832 197940
rect 125692 197616 125744 197668
rect 139584 197820 139636 197872
rect 139952 197820 140004 197872
rect 140320 197820 140372 197872
rect 154856 197956 154908 198008
rect 165068 197956 165120 198008
rect 144276 197888 144328 197940
rect 145288 197888 145340 197940
rect 150716 197888 150768 197940
rect 151636 197888 151688 197940
rect 132132 197548 132184 197600
rect 140780 197752 140832 197804
rect 141148 197752 141200 197804
rect 141516 197752 141568 197804
rect 142068 197752 142120 197804
rect 146116 197820 146168 197872
rect 161480 197820 161532 197872
rect 166908 197956 166960 198008
rect 168656 197956 168708 198008
rect 167092 197888 167144 197940
rect 169760 197888 169812 197940
rect 173164 197888 173216 197940
rect 173348 197888 173400 197940
rect 174544 197956 174596 198008
rect 174820 197956 174872 198008
rect 177948 197956 178000 198008
rect 178224 197956 178276 198008
rect 180708 197956 180760 198008
rect 582564 197956 582616 198008
rect 182180 197888 182232 197940
rect 166540 197820 166592 197872
rect 168196 197820 168248 197872
rect 172704 197820 172756 197872
rect 177580 197820 177632 197872
rect 177856 197820 177908 197872
rect 186412 197820 186464 197872
rect 145288 197752 145340 197804
rect 158260 197752 158312 197804
rect 166724 197752 166776 197804
rect 172520 197752 172572 197804
rect 174544 197752 174596 197804
rect 177672 197752 177724 197804
rect 186320 197752 186372 197804
rect 136732 197684 136784 197736
rect 148232 197684 148284 197736
rect 159364 197684 159416 197736
rect 165896 197684 165948 197736
rect 171784 197684 171836 197736
rect 182088 197684 182140 197736
rect 140044 197616 140096 197668
rect 140688 197616 140740 197668
rect 142252 197616 142304 197668
rect 145012 197616 145064 197668
rect 146392 197616 146444 197668
rect 165620 197616 165672 197668
rect 177764 197616 177816 197668
rect 137100 197548 137152 197600
rect 173072 197548 173124 197600
rect 174728 197548 174780 197600
rect 174912 197548 174964 197600
rect 175280 197548 175332 197600
rect 182640 197548 182692 197600
rect 126612 197480 126664 197532
rect 137284 197480 137336 197532
rect 95700 197412 95752 197464
rect 109132 197412 109184 197464
rect 119988 197412 120040 197464
rect 125600 197412 125652 197464
rect 126888 197412 126940 197464
rect 94688 197344 94740 197396
rect 99288 197344 99340 197396
rect 128360 197344 128412 197396
rect 133144 197344 133196 197396
rect 133880 197344 133932 197396
rect 137100 197344 137152 197396
rect 139492 197344 139544 197396
rect 140320 197344 140372 197396
rect 146576 197480 146628 197532
rect 155040 197480 155092 197532
rect 144184 197412 144236 197464
rect 144644 197412 144696 197464
rect 146392 197412 146444 197464
rect 147680 197412 147732 197464
rect 133972 197276 134024 197328
rect 134340 197276 134392 197328
rect 139308 197276 139360 197328
rect 142988 197344 143040 197396
rect 145196 197344 145248 197396
rect 141516 197276 141568 197328
rect 144828 197276 144880 197328
rect 108580 197208 108632 197260
rect 156604 197208 156656 197260
rect 156880 197208 156932 197260
rect 168196 197480 168248 197532
rect 168840 197480 168892 197532
rect 164240 197412 164292 197464
rect 172060 197412 172112 197464
rect 165344 197344 165396 197396
rect 173440 197344 173492 197396
rect 165068 197276 165120 197328
rect 167092 197276 167144 197328
rect 169944 197276 169996 197328
rect 170680 197276 170732 197328
rect 175188 197276 175240 197328
rect 175464 197276 175516 197328
rect 189080 197276 189132 197328
rect 167276 197208 167328 197260
rect 175924 197208 175976 197260
rect 176568 197208 176620 197260
rect 185676 197208 185728 197260
rect 111064 197140 111116 197192
rect 158168 197140 158220 197192
rect 163780 197140 163832 197192
rect 109132 197072 109184 197124
rect 144276 197072 144328 197124
rect 146208 197072 146260 197124
rect 149060 197072 149112 197124
rect 130660 197004 130712 197056
rect 141884 197004 141936 197056
rect 133972 196936 134024 196988
rect 145656 197004 145708 197056
rect 159088 197004 159140 197056
rect 186504 197140 186556 197192
rect 164884 197072 164936 197124
rect 192484 197072 192536 197124
rect 171140 197004 171192 197056
rect 200764 197004 200816 197056
rect 125416 196868 125468 196920
rect 152832 196936 152884 196988
rect 166080 196936 166132 196988
rect 200304 196936 200356 196988
rect 162768 196868 162820 196920
rect 168564 196868 168616 196920
rect 168748 196868 168800 196920
rect 169116 196868 169168 196920
rect 170404 196868 170456 196920
rect 204720 196868 204772 196920
rect 104808 196800 104860 196852
rect 138572 196800 138624 196852
rect 117964 196732 118016 196784
rect 151912 196800 151964 196852
rect 152280 196800 152332 196852
rect 153016 196800 153068 196852
rect 169024 196800 169076 196852
rect 169300 196800 169352 196852
rect 169576 196800 169628 196852
rect 141332 196732 141384 196784
rect 142804 196732 142856 196784
rect 97724 196664 97776 196716
rect 109040 196664 109092 196716
rect 117780 196664 117832 196716
rect 159180 196732 159232 196784
rect 171784 196732 171836 196784
rect 171968 196732 172020 196784
rect 173256 196732 173308 196784
rect 149796 196664 149848 196716
rect 150072 196664 150124 196716
rect 150808 196664 150860 196716
rect 153476 196664 153528 196716
rect 164240 196664 164292 196716
rect 164516 196664 164568 196716
rect 166356 196664 166408 196716
rect 166908 196664 166960 196716
rect 169852 196664 169904 196716
rect 170680 196664 170732 196716
rect 178408 196800 178460 196852
rect 214196 196800 214248 196852
rect 178592 196732 178644 196784
rect 213920 196732 213972 196784
rect 174544 196664 174596 196716
rect 175188 196664 175240 196716
rect 214012 196664 214064 196716
rect 102048 196596 102100 196648
rect 135444 196596 135496 196648
rect 137468 196596 137520 196648
rect 138572 196596 138624 196648
rect 146944 196596 146996 196648
rect 149152 196596 149204 196648
rect 151636 196596 151688 196648
rect 192760 196596 192812 196648
rect 145380 196528 145432 196580
rect 145748 196528 145800 196580
rect 164516 196528 164568 196580
rect 165160 196528 165212 196580
rect 165252 196528 165304 196580
rect 165528 196528 165580 196580
rect 165896 196528 165948 196580
rect 170404 196528 170456 196580
rect 171324 196528 171376 196580
rect 171876 196528 171928 196580
rect 132224 196460 132276 196512
rect 134984 196460 135036 196512
rect 137468 196460 137520 196512
rect 144092 196460 144144 196512
rect 148508 196460 148560 196512
rect 154120 196460 154172 196512
rect 168564 196460 168616 196512
rect 169208 196460 169260 196512
rect 174176 196460 174228 196512
rect 178224 196460 178276 196512
rect 107016 196392 107068 196444
rect 131764 196324 131816 196376
rect 139308 196324 139360 196376
rect 140044 196324 140096 196376
rect 141792 196324 141844 196376
rect 142528 196324 142580 196376
rect 143080 196324 143132 196376
rect 170588 196324 170640 196376
rect 176568 196324 176620 196376
rect 168104 196256 168156 196308
rect 169208 196256 169260 196308
rect 134984 196188 135036 196240
rect 135812 196188 135864 196240
rect 135996 196188 136048 196240
rect 136180 196188 136232 196240
rect 144828 196188 144880 196240
rect 145564 196188 145616 196240
rect 152556 196188 152608 196240
rect 152740 196188 152792 196240
rect 167184 196188 167236 196240
rect 167644 196188 167696 196240
rect 171232 196188 171284 196240
rect 172244 196188 172296 196240
rect 134892 196120 134944 196172
rect 135628 196120 135680 196172
rect 156604 196120 156656 196172
rect 159548 196120 159600 196172
rect 175280 196120 175332 196172
rect 176384 196120 176436 196172
rect 3608 196052 3660 196104
rect 124404 196052 124456 196104
rect 125416 196052 125468 196104
rect 136180 196052 136232 196104
rect 138204 196052 138256 196104
rect 3516 195984 3568 196036
rect 128360 195984 128412 196036
rect 133972 195984 134024 196036
rect 135812 195984 135864 196036
rect 136548 195984 136600 196036
rect 136916 195984 136968 196036
rect 137100 195984 137152 196036
rect 138112 195984 138164 196036
rect 143816 196052 143868 196104
rect 157800 196052 157852 196104
rect 158352 196052 158404 196104
rect 175464 196052 175516 196104
rect 176292 196052 176344 196104
rect 204444 196052 204496 196104
rect 204720 196052 204772 196104
rect 580172 196052 580224 196104
rect 145564 195984 145616 196036
rect 146300 195984 146352 196036
rect 147772 195984 147824 196036
rect 148048 195984 148100 196036
rect 156972 195984 157024 196036
rect 157248 195984 157300 196036
rect 161848 195984 161900 196036
rect 162124 195984 162176 196036
rect 173992 195984 174044 196036
rect 175004 195984 175056 196036
rect 175740 195984 175792 196036
rect 176016 195984 176068 196036
rect 176752 195984 176804 196036
rect 177304 195984 177356 196036
rect 186504 195984 186556 196036
rect 187516 195984 187568 196036
rect 580632 195984 580684 196036
rect 130384 195916 130436 195968
rect 132316 195916 132368 195968
rect 580264 195916 580316 195968
rect 109868 195848 109920 195900
rect 142344 195848 142396 195900
rect 577688 195848 577740 195900
rect 104532 195780 104584 195832
rect 138112 195780 138164 195832
rect 141976 195780 142028 195832
rect 327724 195780 327776 195832
rect 104440 195712 104492 195764
rect 176936 195712 176988 195764
rect 102968 195644 103020 195696
rect 133052 195576 133104 195628
rect 142804 195576 142856 195628
rect 154212 195576 154264 195628
rect 155408 195576 155460 195628
rect 98828 195508 98880 195560
rect 152556 195508 152608 195560
rect 97816 195440 97868 195492
rect 152464 195440 152516 195492
rect 160008 195644 160060 195696
rect 160192 195644 160244 195696
rect 163596 195644 163648 195696
rect 167276 195576 167328 195628
rect 167828 195576 167880 195628
rect 160376 195508 160428 195560
rect 161664 195508 161716 195560
rect 164148 195508 164200 195560
rect 170772 195644 170824 195696
rect 193588 195644 193640 195696
rect 170496 195576 170548 195628
rect 172888 195576 172940 195628
rect 193220 195576 193272 195628
rect 198004 195508 198056 195560
rect 96252 195372 96304 195424
rect 155960 195372 156012 195424
rect 170956 195372 171008 195424
rect 175832 195440 175884 195492
rect 176292 195440 176344 195492
rect 176936 195440 176988 195492
rect 178040 195440 178092 195492
rect 214288 195440 214340 195492
rect 204260 195372 204312 195424
rect 3424 195304 3476 195356
rect 120172 195236 120224 195288
rect 121460 195236 121512 195288
rect 126336 195236 126388 195288
rect 133052 195236 133104 195288
rect 138664 195236 138716 195288
rect 140780 195236 140832 195288
rect 160376 195304 160428 195356
rect 160560 195304 160612 195356
rect 177304 195304 177356 195356
rect 214564 195304 214616 195356
rect 167644 195236 167696 195288
rect 200764 195236 200816 195288
rect 214380 195236 214432 195288
rect 580816 195236 580868 195288
rect 111708 195168 111760 195220
rect 143264 195168 143316 195220
rect 124128 195100 124180 195152
rect 134984 195100 135036 195152
rect 152464 195100 152516 195152
rect 156604 195100 156656 195152
rect 156696 195032 156748 195084
rect 192024 195168 192076 195220
rect 168288 195100 168340 195152
rect 175188 195100 175240 195152
rect 167736 195032 167788 195084
rect 178684 195032 178736 195084
rect 142804 194964 142856 195016
rect 149336 194964 149388 195016
rect 206284 194964 206336 195016
rect 108396 194896 108448 194948
rect 175188 194896 175240 194948
rect 180064 194896 180116 194948
rect 174912 194828 174964 194880
rect 177304 194828 177356 194880
rect 132040 194760 132092 194812
rect 134524 194760 134576 194812
rect 152556 194760 152608 194812
rect 157616 194760 157668 194812
rect 160744 194760 160796 194812
rect 139860 194556 139912 194608
rect 142436 194556 142488 194608
rect 114836 194488 114888 194540
rect 149244 194488 149296 194540
rect 149796 194488 149848 194540
rect 152740 194488 152792 194540
rect 578976 194488 579028 194540
rect 107108 194420 107160 194472
rect 114468 194420 114520 194472
rect 122104 194420 122156 194472
rect 141516 194420 141568 194472
rect 142620 194420 142672 194472
rect 567844 194420 567896 194472
rect 107476 194352 107528 194404
rect 118700 194352 118752 194404
rect 139952 194352 140004 194404
rect 564072 194352 564124 194404
rect 104256 194284 104308 194336
rect 177120 194284 177172 194336
rect 107200 194216 107252 194268
rect 161940 194216 161992 194268
rect 174360 194216 174412 194268
rect 192300 194216 192352 194268
rect 108672 194148 108724 194200
rect 163320 194148 163372 194200
rect 163596 194148 163648 194200
rect 174084 194148 174136 194200
rect 175096 194148 175148 194200
rect 176476 194148 176528 194200
rect 198832 194148 198884 194200
rect 107016 194080 107068 194132
rect 139952 194080 140004 194132
rect 157708 194080 157760 194132
rect 158444 194080 158496 194132
rect 158720 194080 158772 194132
rect 185768 194080 185820 194132
rect 189540 194080 189592 194132
rect 104716 194012 104768 194064
rect 135076 194012 135128 194064
rect 162400 194012 162452 194064
rect 189724 194012 189776 194064
rect 209872 194012 209924 194064
rect 95608 193944 95660 193996
rect 110512 193944 110564 193996
rect 111800 193944 111852 193996
rect 118424 193944 118476 193996
rect 149796 193944 149848 193996
rect 166172 193944 166224 193996
rect 172152 193944 172204 193996
rect 172796 193944 172848 193996
rect 207020 193944 207072 193996
rect 101956 193876 102008 193928
rect 140688 193876 140740 193928
rect 157432 193876 157484 193928
rect 173164 193876 173216 193928
rect 177120 193876 177172 193928
rect 212724 193876 212776 193928
rect 99380 193808 99432 193860
rect 103336 193808 103388 193860
rect 158628 193808 158680 193860
rect 171416 193808 171468 193860
rect 205732 193808 205784 193860
rect 207020 193808 207072 193860
rect 502340 193808 502392 193860
rect 116308 193740 116360 193792
rect 148324 193740 148376 193792
rect 161664 193740 161716 193792
rect 178960 193740 179012 193792
rect 119988 193672 120040 193724
rect 148600 193672 148652 193724
rect 172980 193672 173032 193724
rect 173348 193672 173400 193724
rect 131028 193604 131080 193656
rect 161204 193604 161256 193656
rect 169944 193604 169996 193656
rect 170864 193604 170916 193656
rect 138020 193536 138072 193588
rect 138940 193536 138992 193588
rect 144184 193536 144236 193588
rect 144920 193536 144972 193588
rect 152556 193536 152608 193588
rect 152924 193536 152976 193588
rect 164608 193400 164660 193452
rect 165436 193400 165488 193452
rect 168472 193400 168524 193452
rect 169484 193400 169536 193452
rect 152924 193332 152976 193384
rect 104624 193196 104676 193248
rect 177304 193264 177356 193316
rect 189356 193264 189408 193316
rect 198096 193196 198148 193248
rect 111800 193060 111852 193112
rect 147312 193128 147364 193180
rect 168380 193128 168432 193180
rect 577596 193128 577648 193180
rect 145104 193060 145156 193112
rect 281540 193060 281592 193112
rect 111340 192992 111392 193044
rect 141332 192992 141384 193044
rect 148600 192992 148652 193044
rect 151084 192992 151136 193044
rect 189448 192992 189500 193044
rect 114468 192924 114520 192976
rect 136732 192924 136784 192976
rect 173624 192924 173676 192976
rect 198740 192924 198792 192976
rect 120172 192856 120224 192908
rect 138296 192856 138348 192908
rect 173256 192856 173308 192908
rect 206192 192856 206244 192908
rect 118240 192788 118292 192840
rect 139492 192788 139544 192840
rect 169300 192788 169352 192840
rect 202880 192788 202932 192840
rect 127624 192720 127676 192772
rect 153752 192720 153804 192772
rect 162492 192720 162544 192772
rect 196072 192720 196124 192772
rect 121276 192652 121328 192704
rect 150808 192652 150860 192704
rect 154028 192652 154080 192704
rect 196716 192652 196768 192704
rect 119528 192584 119580 192636
rect 144828 192584 144880 192636
rect 146760 192584 146812 192636
rect 191840 192584 191892 192636
rect 202880 192584 202932 192636
rect 575112 192584 575164 192636
rect 114468 192516 114520 192568
rect 139860 192516 139912 192568
rect 86316 192448 86368 192500
rect 120172 192448 120224 192500
rect 126428 192448 126480 192500
rect 148600 192448 148652 192500
rect 121828 192380 121880 192432
rect 135628 192380 135680 192432
rect 131948 192312 132000 192364
rect 145472 192312 145524 192364
rect 544384 192516 544436 192568
rect 150348 192448 150400 192500
rect 579620 192448 579672 192500
rect 167552 192380 167604 192432
rect 184204 192380 184256 192432
rect 169760 192312 169812 192364
rect 178040 192312 178092 192364
rect 94780 192244 94832 192296
rect 173256 192244 173308 192296
rect 25504 191836 25556 191888
rect 125692 191836 125744 191888
rect 101496 191768 101548 191820
rect 118148 191768 118200 191820
rect 127716 191768 127768 191820
rect 128452 191768 128504 191820
rect 130476 191768 130528 191820
rect 133880 191768 133932 191820
rect 134248 191768 134300 191820
rect 175004 191836 175056 191888
rect 182916 191836 182968 191888
rect 145012 191768 145064 191820
rect 575020 191768 575072 191820
rect 57980 191700 58032 191752
rect 158628 191700 158680 191752
rect 160928 191700 160980 191752
rect 174176 191700 174228 191752
rect 174728 191700 174780 191752
rect 198004 191700 198056 191752
rect 572260 191700 572312 191752
rect 101404 191632 101456 191684
rect 184940 191632 184992 191684
rect 197728 191632 197780 191684
rect 566464 191632 566516 191684
rect 99012 191564 99064 191616
rect 165252 191564 165304 191616
rect 175924 191564 175976 191616
rect 398840 191564 398892 191616
rect 95884 191496 95936 191548
rect 159456 191496 159508 191548
rect 178868 191496 178920 191548
rect 104072 191428 104124 191480
rect 108672 191428 108724 191480
rect 112996 191428 113048 191480
rect 168932 191428 168984 191480
rect 184848 191428 184900 191480
rect 195980 191428 196032 191480
rect 100484 191360 100536 191412
rect 133880 191360 133932 191412
rect 134156 191360 134208 191412
rect 134432 191360 134484 191412
rect 135720 191360 135772 191412
rect 136364 191360 136416 191412
rect 137376 191360 137428 191412
rect 137928 191360 137980 191412
rect 138112 191360 138164 191412
rect 143908 191360 143960 191412
rect 148692 191360 148744 191412
rect 148876 191360 148928 191412
rect 160100 191360 160152 191412
rect 160560 191360 160612 191412
rect 160928 191360 160980 191412
rect 178776 191360 178828 191412
rect 184940 191360 184992 191412
rect 200396 191360 200448 191412
rect 108672 191292 108724 191344
rect 143172 191292 143224 191344
rect 115848 191224 115900 191276
rect 122012 191224 122064 191276
rect 156420 191292 156472 191344
rect 160284 191292 160336 191344
rect 194600 191292 194652 191344
rect 197360 191292 197412 191344
rect 216864 191292 216916 191344
rect 153292 191224 153344 191276
rect 154120 191224 154172 191276
rect 158996 191224 159048 191276
rect 159916 191224 159968 191276
rect 162768 191224 162820 191276
rect 164424 191224 164476 191276
rect 164516 191224 164568 191276
rect 84936 191088 84988 191140
rect 105912 191156 105964 191208
rect 138112 191156 138164 191208
rect 138296 191156 138348 191208
rect 139032 191156 139084 191208
rect 140136 191156 140188 191208
rect 140688 191156 140740 191208
rect 142804 191156 142856 191208
rect 142988 191156 143040 191208
rect 145472 191156 145524 191208
rect 146024 191156 146076 191208
rect 146484 191156 146536 191208
rect 147128 191156 147180 191208
rect 149152 191156 149204 191208
rect 149888 191156 149940 191208
rect 150624 191156 150676 191208
rect 151360 191156 151412 191208
rect 153476 191156 153528 191208
rect 154396 191156 154448 191208
rect 154948 191156 155000 191208
rect 155500 191156 155552 191208
rect 156144 191156 156196 191208
rect 156972 191156 157024 191208
rect 158904 191156 158956 191208
rect 159732 191156 159784 191208
rect 160192 191156 160244 191208
rect 160468 191156 160520 191208
rect 161756 191156 161808 191208
rect 162032 191156 162084 191208
rect 163412 191156 163464 191208
rect 163964 191156 164016 191208
rect 165712 191156 165764 191208
rect 166264 191156 166316 191208
rect 166908 191224 166960 191276
rect 200212 191224 200264 191276
rect 206560 191156 206612 191208
rect 207664 191156 207716 191208
rect 509240 191156 509292 191208
rect 112260 191088 112312 191140
rect 173900 191088 173952 191140
rect 175004 191088 175056 191140
rect 190000 191088 190052 191140
rect 210424 191088 210476 191140
rect 216864 191088 216916 191140
rect 520280 191088 520332 191140
rect 118148 191020 118200 191072
rect 132868 190952 132920 191004
rect 133604 190952 133656 191004
rect 134616 190952 134668 191004
rect 135536 190952 135588 191004
rect 136088 190952 136140 191004
rect 136180 190952 136232 191004
rect 136548 190952 136600 191004
rect 137192 190952 137244 191004
rect 137836 190952 137888 191004
rect 146576 191020 146628 191072
rect 147588 191020 147640 191072
rect 148140 191020 148192 191072
rect 148692 191020 148744 191072
rect 149336 191020 149388 191072
rect 150256 191020 150308 191072
rect 153384 191020 153436 191072
rect 154120 191020 154172 191072
rect 154672 191020 154724 191072
rect 155592 191020 155644 191072
rect 156604 191020 156656 191072
rect 156880 191020 156932 191072
rect 159916 191020 159968 191072
rect 160100 191020 160152 191072
rect 160284 191020 160336 191072
rect 160836 191020 160888 191072
rect 164516 191020 164568 191072
rect 165344 191020 165396 191072
rect 151636 190952 151688 191004
rect 164056 190952 164108 191004
rect 197360 191020 197412 191072
rect 197728 191020 197780 191072
rect 132776 190884 132828 190936
rect 133788 190884 133840 190936
rect 134248 190884 134300 190936
rect 136824 190884 136876 190936
rect 137560 190884 137612 190936
rect 116584 190544 116636 190596
rect 162768 190544 162820 190596
rect 174176 190544 174228 190596
rect 189540 190544 189592 190596
rect 4896 190476 4948 190528
rect 100484 190476 100536 190528
rect 137376 190476 137428 190528
rect 137928 190476 137980 190528
rect 490564 190476 490616 190528
rect 94596 190408 94648 190460
rect 165620 190408 165672 190460
rect 186136 190408 186188 190460
rect 563704 190408 563756 190460
rect 99104 190340 99156 190392
rect 167000 190340 167052 190392
rect 170404 190340 170456 190392
rect 193956 190340 194008 190392
rect 206284 190340 206336 190392
rect 579988 190340 580040 190392
rect 117228 190272 117280 190324
rect 173716 190272 173768 190324
rect 152280 190204 152332 190256
rect 152464 190204 152516 190256
rect 177580 190204 177632 190256
rect 205824 190204 205876 190256
rect 155776 190136 155828 190188
rect 187792 190136 187844 190188
rect 121000 190068 121052 190120
rect 148508 190068 148560 190120
rect 155868 190068 155920 190120
rect 189172 190068 189224 190120
rect 109684 190000 109736 190052
rect 119436 190000 119488 190052
rect 151912 190000 151964 190052
rect 163596 190000 163648 190052
rect 197728 190000 197780 190052
rect 110972 189932 111024 189984
rect 144368 189932 144420 189984
rect 156788 189932 156840 189984
rect 190828 189932 190880 189984
rect 110880 189864 110932 189916
rect 145840 189864 145892 189916
rect 158352 189864 158404 189916
rect 217232 189864 217284 189916
rect 572076 189864 572128 189916
rect 95976 189796 96028 189848
rect 109500 189796 109552 189848
rect 144552 189796 144604 189848
rect 158076 189796 158128 189848
rect 192392 189796 192444 189848
rect 207756 189796 207808 189848
rect 569224 189796 569276 189848
rect 90364 189728 90416 189780
rect 97080 189728 97132 189780
rect 155132 189728 155184 189780
rect 159272 189728 159324 189780
rect 183376 189728 183428 189780
rect 563888 189728 563940 189780
rect 163872 189660 163924 189712
rect 191932 189660 191984 189712
rect 154856 189592 154908 189644
rect 155224 189592 155276 189644
rect 167000 189116 167052 189168
rect 167368 189116 167420 189168
rect 108028 189048 108080 189100
rect 149704 188980 149756 189032
rect 150164 188980 150216 189032
rect 165620 189048 165672 189100
rect 167092 189048 167144 189100
rect 152096 188980 152148 189032
rect 566740 188980 566792 189032
rect 106188 188912 106240 188964
rect 152188 188912 152240 188964
rect 172612 188844 172664 188896
rect 207388 188844 207440 188896
rect 207756 188844 207808 188896
rect 158536 188776 158588 188828
rect 201500 188776 201552 188828
rect 129004 188708 129056 188760
rect 153936 188708 153988 188760
rect 251180 188708 251232 188760
rect 93216 188640 93268 188692
rect 173532 188640 173584 188692
rect 206100 188640 206152 188692
rect 106280 188572 106332 188624
rect 176936 188572 176988 188624
rect 210148 188572 210200 188624
rect 95976 188504 96028 188556
rect 104900 188504 104952 188556
rect 106188 188504 106240 188556
rect 108488 188504 108540 188556
rect 178224 188504 178276 188556
rect 103060 188436 103112 188488
rect 104624 188436 104676 188488
rect 137100 188436 137152 188488
rect 215760 188436 215812 188488
rect 101680 188368 101732 188420
rect 111524 188368 111576 188420
rect 144644 188368 144696 188420
rect 167000 188368 167052 188420
rect 167460 188368 167512 188420
rect 216956 188368 217008 188420
rect 27620 188300 27672 188352
rect 99748 188300 99800 188352
rect 132592 188300 132644 188352
rect 154304 188300 154356 188352
rect 218428 188300 218480 188352
rect 563980 188300 564032 188352
rect 101588 188232 101640 188284
rect 166632 188232 166684 188284
rect 180248 188164 180300 188216
rect 49700 188096 49752 188148
rect 167000 188096 167052 188148
rect 3240 188028 3292 188080
rect 175740 188028 175792 188080
rect 207296 188232 207348 188284
rect 149704 187960 149756 188012
rect 471980 187960 472032 188012
rect 130752 187824 130804 187876
rect 148232 187824 148284 187876
rect 148968 187824 149020 187876
rect 124864 187756 124916 187808
rect 109776 187688 109828 187740
rect 201500 187688 201552 187740
rect 207112 187688 207164 187740
rect 145564 187620 145616 187672
rect 579068 187620 579120 187672
rect 150348 187552 150400 187604
rect 569316 187552 569368 187604
rect 90640 187484 90692 187536
rect 177304 187484 177356 187536
rect 177396 187484 177448 187536
rect 177948 187484 178000 187536
rect 313924 187484 313976 187536
rect 96160 187416 96212 187468
rect 174176 187416 174228 187468
rect 110144 187348 110196 187400
rect 142712 187348 142764 187400
rect 168840 187348 168892 187400
rect 203064 187348 203116 187400
rect 110052 187280 110104 187332
rect 143356 187280 143408 187332
rect 165252 187280 165304 187332
rect 199384 187280 199436 187332
rect 99656 187212 99708 187264
rect 133420 187212 133472 187264
rect 155960 187212 156012 187264
rect 156328 187212 156380 187264
rect 170404 187212 170456 187264
rect 175648 187212 175700 187264
rect 210240 187212 210292 187264
rect 112444 187144 112496 187196
rect 144920 187144 144972 187196
rect 164976 187144 165028 187196
rect 199292 187144 199344 187196
rect 109960 187076 110012 187128
rect 143724 187076 143776 187128
rect 167184 187076 167236 187128
rect 201960 187076 202012 187128
rect 113732 187008 113784 187060
rect 148416 187008 148468 187060
rect 170312 187008 170364 187060
rect 204812 187008 204864 187060
rect 96068 186940 96120 186992
rect 121092 186940 121144 186992
rect 157156 186940 157208 186992
rect 158168 186940 158220 186992
rect 193864 186940 193916 186992
rect 572168 186940 572220 186992
rect 115480 186872 115532 186924
rect 147312 186872 147364 186924
rect 167276 186872 167328 186924
rect 201500 186872 201552 186924
rect 106096 186804 106148 186856
rect 136364 186804 136416 186856
rect 161940 186804 161992 186856
rect 195980 186804 196032 186856
rect 97448 186736 97500 186788
rect 155960 186736 156012 186788
rect 170772 186736 170824 186788
rect 202972 186736 203024 186788
rect 108304 186668 108356 186720
rect 154580 186668 154632 186720
rect 166264 186668 166316 186720
rect 107108 186328 107160 186380
rect 129740 186328 129792 186380
rect 8300 186260 8352 186312
rect 176752 186260 176804 186312
rect 30380 186192 30432 186244
rect 178132 186192 178184 186244
rect 129740 186124 129792 186176
rect 143448 186124 143500 186176
rect 273260 186124 273312 186176
rect 93400 186056 93452 186108
rect 175556 186056 175608 186108
rect 210056 186056 210108 186108
rect 100208 185988 100260 186040
rect 180800 185988 180852 186040
rect 210516 185988 210568 186040
rect 103152 185920 103204 185972
rect 176660 185920 176712 185972
rect 178132 185920 178184 185972
rect 208676 185920 208728 185972
rect 87604 185852 87656 185904
rect 107384 185852 107436 185904
rect 127900 185852 127952 185904
rect 132960 185852 133012 185904
rect 205640 185852 205692 185904
rect 97540 185784 97592 185836
rect 168380 185784 168432 185836
rect 176660 185784 176712 185836
rect 211712 185784 211764 185836
rect 100116 185716 100168 185768
rect 170220 185716 170272 185768
rect 212816 185716 212868 185768
rect 218152 185716 218204 185768
rect 218336 185716 218388 185768
rect 240140 185716 240192 185768
rect 98920 185648 98972 185700
rect 103060 185648 103112 185700
rect 135536 185648 135588 185700
rect 158904 185648 158956 185700
rect 100300 185580 100352 185632
rect 135168 185580 135220 185632
rect 155040 185580 155092 185632
rect 218152 185580 218204 185632
rect 221004 185580 221056 185632
rect 581644 185580 581696 185632
rect 107200 185512 107252 185564
rect 107384 185512 107436 185564
rect 136272 185512 136324 185564
rect 161848 185512 161900 185564
rect 184296 185512 184348 185564
rect 184848 185512 184900 185564
rect 161756 185444 161808 185496
rect 181904 185444 181956 185496
rect 218152 185444 218204 185496
rect 218428 185444 218480 185496
rect 168380 184968 168432 185020
rect 207480 184968 207532 185020
rect 181904 184900 181956 184952
rect 580172 184900 580224 184952
rect 131120 184832 131172 184884
rect 145380 184832 145432 184884
rect 418160 184832 418212 184884
rect 90456 184764 90508 184816
rect 177304 184764 177356 184816
rect 177764 184764 177816 184816
rect 90548 184696 90600 184748
rect 164516 184696 164568 184748
rect 165528 184696 165580 184748
rect 167092 184696 167144 184748
rect 200488 184696 200540 184748
rect 97264 184628 97316 184680
rect 168748 184628 168800 184680
rect 173716 184628 173768 184680
rect 204904 184628 204956 184680
rect 104348 184560 104400 184612
rect 134616 184560 134668 184612
rect 167368 184560 167420 184612
rect 201868 184560 201920 184612
rect 108580 184492 108632 184544
rect 139768 184492 139820 184544
rect 171416 184492 171468 184544
rect 205916 184492 205968 184544
rect 101312 184424 101364 184476
rect 134248 184424 134300 184476
rect 171324 184424 171376 184476
rect 206008 184424 206060 184476
rect 106188 184356 106240 184408
rect 140504 184356 140556 184408
rect 169852 184356 169904 184408
rect 204720 184356 204772 184408
rect 109684 184288 109736 184340
rect 144460 184288 144512 184340
rect 171048 184288 171100 184340
rect 206284 184288 206336 184340
rect 104440 184220 104492 184272
rect 138296 184220 138348 184272
rect 165528 184220 165580 184272
rect 206376 184220 206428 184272
rect 3148 184152 3200 184204
rect 171968 184152 172020 184204
rect 174084 184152 174136 184204
rect 208584 184152 208636 184204
rect 103244 184084 103296 184136
rect 132224 184084 132276 184136
rect 107384 184016 107436 184068
rect 132132 184016 132184 184068
rect 97356 183948 97408 184000
rect 110420 183948 110472 184000
rect 102968 183880 103020 183932
rect 132868 183880 132920 183932
rect 100024 183472 100076 183524
rect 182272 183472 182324 183524
rect 103520 183404 103572 183456
rect 84844 183336 84896 183388
rect 160008 183336 160060 183388
rect 107292 183268 107344 183320
rect 108304 183268 108356 183320
rect 110420 183268 110472 183320
rect 111064 183268 111116 183320
rect 142896 183268 142948 183320
rect 104992 183200 105044 183252
rect 105820 183200 105872 183252
rect 135812 183200 135864 183252
rect 208768 183336 208820 183388
rect 182180 183268 182232 183320
rect 212632 183268 212684 183320
rect 209780 183200 209832 183252
rect 158352 183132 158404 183184
rect 211344 183132 211396 183184
rect 227720 183132 227772 183184
rect 159916 183064 159968 183116
rect 176568 183064 176620 183116
rect 247040 183064 247092 183116
rect 160376 182996 160428 183048
rect 176384 182996 176436 183048
rect 349160 182996 349212 183048
rect 154948 182928 155000 182980
rect 221096 182928 221148 182980
rect 552756 182928 552808 182980
rect 96528 182860 96580 182912
rect 120540 182860 120592 182912
rect 140964 182860 141016 182912
rect 153476 182860 153528 182912
rect 188620 182860 188672 182912
rect 569408 182860 569460 182912
rect 108304 182792 108356 182844
rect 139676 182792 139728 182844
rect 158168 182792 158220 182844
rect 177764 182792 177816 182844
rect 575204 182792 575256 182844
rect 102876 182180 102928 182232
rect 105820 182180 105872 182232
rect 123116 182112 123168 182164
rect 123576 182112 123628 182164
rect 125508 182112 125560 182164
rect 125784 182112 125836 182164
rect 147864 182112 147916 182164
rect 148416 182112 148468 182164
rect 149336 182112 149388 182164
rect 149796 182112 149848 182164
rect 149888 182112 149940 182164
rect 572352 182112 572404 182164
rect 108396 181976 108448 182028
rect 141884 182044 141936 182096
rect 561220 182044 561272 182096
rect 107292 181908 107344 181960
rect 139584 181976 139636 182028
rect 148416 181976 148468 182028
rect 277400 181976 277452 182028
rect 137560 181908 137612 181960
rect 140228 181908 140280 181960
rect 253940 181908 253992 181960
rect 104256 181840 104308 181892
rect 137008 181840 137060 181892
rect 153292 181840 153344 181892
rect 210608 181840 210660 181892
rect 217416 181840 217468 181892
rect 113824 181772 113876 181824
rect 146668 181772 146720 181824
rect 149888 181772 149940 181824
rect 154764 181772 154816 181824
rect 189448 181772 189500 181824
rect 119620 181704 119672 181756
rect 152648 181704 152700 181756
rect 175464 181704 175516 181756
rect 210332 181704 210384 181756
rect 103428 181636 103480 181688
rect 137744 181636 137796 181688
rect 160284 181636 160336 181688
rect 195152 181636 195204 181688
rect 105636 181568 105688 181620
rect 138940 181568 138992 181620
rect 150624 181568 150676 181620
rect 220820 181568 220872 181620
rect 99104 181500 99156 181552
rect 132776 181500 132828 181552
rect 152372 181500 152424 181552
rect 219992 181500 220044 181552
rect 299480 181500 299532 181552
rect 125784 181432 125836 181484
rect 292580 181432 292632 181484
rect 176752 181364 176804 181416
rect 211896 181364 211948 181416
rect 166264 181296 166316 181348
rect 189264 181296 189316 181348
rect 102784 180956 102836 181008
rect 123116 180956 123168 181008
rect 103152 180888 103204 180940
rect 126888 180888 126940 180940
rect 101772 180820 101824 180872
rect 129648 180820 129700 180872
rect 195152 180820 195204 180872
rect 580172 180820 580224 180872
rect 3240 180752 3292 180804
rect 112260 180752 112312 180804
rect 129188 180752 129240 180804
rect 555424 180752 555476 180804
rect 126888 180684 126940 180736
rect 136548 180684 136600 180736
rect 558460 180684 558512 180736
rect 127992 180616 128044 180668
rect 541624 180616 541676 180668
rect 129648 180548 129700 180600
rect 140044 180548 140096 180600
rect 552848 180548 552900 180600
rect 128176 180480 128228 180532
rect 498200 180480 498252 180532
rect 128728 180412 128780 180464
rect 138756 180412 138808 180464
rect 405740 180412 405792 180464
rect 123116 180344 123168 180396
rect 322940 180344 322992 180396
rect 80704 180276 80756 180328
rect 186320 180276 186372 180328
rect 86224 180208 86276 180260
rect 186412 180208 186464 180260
rect 213000 180140 213052 180192
rect 186320 180072 186372 180124
rect 219900 180072 219952 180124
rect 105728 179392 105780 179444
rect 126704 179324 126756 179376
rect 582656 179324 582708 179376
rect 164424 179120 164476 179172
rect 186504 179120 186556 179172
rect 163780 179052 163832 179104
rect 190460 179052 190512 179104
rect 156144 178984 156196 179036
rect 186596 178984 186648 179036
rect 101864 178916 101916 178968
rect 134156 178916 134208 178968
rect 177304 178916 177356 178968
rect 211528 178916 211580 178968
rect 87696 178848 87748 178900
rect 104164 178848 104216 178900
rect 136916 178848 136968 178900
rect 171232 178848 171284 178900
rect 215852 178848 215904 178900
rect 100392 178780 100444 178832
rect 134064 178780 134116 178832
rect 154672 178780 154724 178832
rect 217324 178780 217376 178832
rect 101680 178712 101732 178764
rect 135996 178712 136048 178764
rect 160192 178712 160244 178764
rect 184848 178712 184900 178764
rect 309784 178712 309836 178764
rect 109592 178644 109644 178696
rect 150900 178644 150952 178696
rect 161296 178644 161348 178696
rect 214748 178644 214800 178696
rect 425060 178644 425112 178696
rect 95148 178032 95200 178084
rect 134524 178032 134576 178084
rect 135168 178032 135220 178084
rect 126612 177964 126664 178016
rect 582380 177964 582432 178016
rect 124128 177896 124180 177948
rect 561312 177896 561364 177948
rect 135168 177828 135220 177880
rect 556988 177828 557040 177880
rect 140780 177760 140832 177812
rect 141148 177760 141200 177812
rect 555516 177760 555568 177812
rect 105820 177352 105872 177404
rect 140136 177692 140188 177744
rect 409880 177692 409932 177744
rect 137468 177624 137520 177676
rect 364340 177624 364392 177676
rect 136824 177420 136876 177472
rect 137468 177420 137520 177472
rect 192760 177352 192812 177404
rect 221740 177352 221792 177404
rect 105544 177284 105596 177336
rect 140780 177284 140832 177336
rect 141332 177284 141384 177336
rect 142160 177284 142212 177336
rect 558552 177284 558604 177336
rect 221280 176672 221332 176724
rect 221740 176672 221792 176724
rect 579804 176672 579856 176724
rect 133788 176604 133840 176656
rect 559656 176604 559708 176656
rect 156604 176060 156656 176112
rect 190920 176060 190972 176112
rect 169116 175992 169168 176044
rect 208952 175992 209004 176044
rect 99012 175924 99064 175976
rect 132684 175924 132736 175976
rect 133788 175924 133840 175976
rect 167644 175924 167696 175976
rect 207664 175924 207716 175976
rect 135168 175176 135220 175228
rect 565084 175176 565136 175228
rect 140872 175108 140924 175160
rect 562324 175108 562376 175160
rect 140780 175040 140832 175092
rect 368480 175040 368532 175092
rect 136548 174972 136600 175024
rect 357440 174972 357492 175024
rect 101496 174700 101548 174752
rect 134616 174700 134668 174752
rect 135168 174700 135220 174752
rect 102692 174632 102744 174684
rect 135904 174632 135956 174684
rect 353300 174904 353352 174956
rect 101588 174564 101640 174616
rect 136548 174564 136600 174616
rect 106924 174496 106976 174548
rect 140780 174496 140832 174548
rect 124036 173884 124088 173936
rect 140872 173884 140924 173936
rect 3240 172456 3292 172508
rect 116584 172456 116636 172508
rect 3332 168308 3384 168360
rect 25504 168308 25556 168360
rect 172244 164840 172296 164892
rect 204996 164840 205048 164892
rect 204996 164228 205048 164280
rect 580172 164228 580224 164280
rect 97448 163480 97500 163532
rect 146576 163480 146628 163532
rect 3056 162868 3108 162920
rect 97448 162868 97500 162920
rect 198096 157292 198148 157344
rect 580172 157292 580224 157344
rect 3516 155864 3568 155916
rect 117780 155864 117832 155916
rect 180248 155184 180300 155236
rect 197360 155184 197412 155236
rect 192484 153144 192536 153196
rect 199476 153144 199528 153196
rect 199476 151784 199528 151836
rect 579804 151784 579856 151836
rect 100024 151240 100076 151292
rect 132040 151240 132092 151292
rect 173348 151240 173400 151292
rect 205088 151240 205140 151292
rect 94964 151172 95016 151224
rect 138204 151172 138256 151224
rect 176016 151172 176068 151224
rect 209136 151172 209188 151224
rect 95884 151104 95936 151156
rect 140688 151104 140740 151156
rect 171876 151104 171928 151156
rect 209044 151104 209096 151156
rect 95056 151036 95108 151088
rect 140412 151036 140464 151088
rect 154304 151036 154356 151088
rect 218612 151036 218664 151088
rect 106832 148996 106884 149048
rect 131304 148996 131356 149048
rect 176292 148996 176344 149048
rect 207756 148996 207808 149048
rect 101220 148928 101272 148980
rect 126520 148928 126572 148980
rect 162768 148928 162820 148980
rect 195428 148928 195480 148980
rect 102600 148860 102652 148912
rect 135720 148860 135772 148912
rect 177488 148860 177540 148912
rect 210608 148860 210660 148912
rect 103980 148792 104032 148844
rect 137376 148792 137428 148844
rect 170680 148792 170732 148844
rect 203248 148792 203300 148844
rect 114928 148724 114980 148776
rect 150256 148724 150308 148776
rect 168656 148724 168708 148776
rect 203432 148724 203484 148776
rect 98828 148656 98880 148708
rect 133236 148656 133288 148708
rect 168564 148656 168616 148708
rect 203340 148656 203392 148708
rect 98920 148588 98972 148640
rect 133328 148588 133380 148640
rect 165896 148588 165948 148640
rect 200672 148588 200724 148640
rect 99932 148520 99984 148572
rect 134432 148520 134484 148572
rect 165804 148520 165856 148572
rect 200580 148520 200632 148572
rect 98736 148452 98788 148504
rect 133144 148452 133196 148504
rect 165436 148452 165488 148504
rect 199660 148452 199712 148504
rect 101404 148384 101456 148436
rect 137560 148384 137612 148436
rect 168288 148384 168340 148436
rect 203616 148384 203668 148436
rect 96528 148316 96580 148368
rect 130384 148316 130436 148368
rect 174544 148316 174596 148368
rect 211988 148316 212040 148368
rect 106740 148248 106792 148300
rect 127900 148248 127952 148300
rect 175280 148248 175332 148300
rect 206468 148248 206520 148300
rect 121184 148180 121236 148232
rect 127808 148180 127860 148232
rect 172152 148180 172204 148232
rect 200764 148180 200816 148232
rect 120724 148112 120776 148164
rect 125692 148112 125744 148164
rect 169392 148112 169444 148164
rect 191380 148112 191432 148164
rect 3424 147568 3476 147620
rect 114100 147568 114152 147620
rect 120908 147568 120960 147620
rect 185676 147228 185728 147280
rect 196440 147228 196492 147280
rect 580356 147568 580408 147620
rect 165712 147160 165764 147212
rect 192760 147160 192812 147212
rect 169024 147092 169076 147144
rect 203524 147092 203576 147144
rect 117044 147024 117096 147076
rect 117228 147024 117280 147076
rect 168104 147024 168156 147076
rect 202144 147024 202196 147076
rect 111432 146956 111484 147008
rect 138664 146956 138716 147008
rect 154120 146956 154172 147008
rect 187700 146956 187752 147008
rect 188160 146956 188212 147008
rect 188988 146956 189040 147008
rect 104072 146888 104124 146940
rect 139032 146888 139084 146940
rect 156696 146888 156748 146940
rect 216036 146888 216088 146940
rect 179696 146344 179748 146396
rect 180156 146344 180208 146396
rect 215944 146344 215996 146396
rect 216036 146344 216088 146396
rect 580816 146344 580868 146396
rect 187700 146276 187752 146328
rect 188804 146276 188856 146328
rect 580908 146276 580960 146328
rect 117872 146208 117924 146260
rect 130108 146208 130160 146260
rect 171508 146208 171560 146260
rect 196256 146208 196308 146260
rect 490564 146208 490616 146260
rect 580172 146208 580224 146260
rect 112352 146140 112404 146192
rect 129372 146140 129424 146192
rect 172520 146140 172572 146192
rect 199200 146140 199252 146192
rect 114284 146072 114336 146124
rect 134800 146072 134852 146124
rect 164424 146072 164476 146124
rect 193772 146072 193824 146124
rect 111156 146004 111208 146056
rect 132592 146004 132644 146056
rect 166540 146004 166592 146056
rect 196348 146004 196400 146056
rect 111248 145936 111300 145988
rect 137192 145936 137244 145988
rect 167368 145936 167420 145988
rect 199108 145936 199160 145988
rect 112720 145868 112772 145920
rect 139400 145868 139452 145920
rect 162400 145868 162452 145920
rect 194784 145868 194836 145920
rect 114008 145800 114060 145852
rect 144920 145800 144972 145852
rect 164884 145800 164936 145852
rect 197820 145800 197872 145852
rect 114192 145732 114244 145784
rect 146484 145732 146536 145784
rect 156604 145732 156656 145784
rect 190736 145732 190788 145784
rect 116768 145664 116820 145716
rect 149980 145664 150032 145716
rect 160100 145664 160152 145716
rect 194968 145664 195020 145716
rect 112720 145596 112772 145648
rect 146576 145596 146628 145648
rect 157432 145596 157484 145648
rect 192576 145596 192628 145648
rect 112260 145528 112312 145580
rect 151176 145528 151228 145580
rect 154948 145528 155000 145580
rect 189908 145528 189960 145580
rect 112168 145460 112220 145512
rect 123392 145460 123444 145512
rect 176660 145460 176712 145512
rect 196532 145460 196584 145512
rect 116676 145392 116728 145444
rect 127716 145392 127768 145444
rect 179420 145392 179472 145444
rect 197544 145392 197596 145444
rect 114100 145324 114152 145376
rect 124220 145324 124272 145376
rect 180800 145324 180852 145376
rect 197912 145324 197964 145376
rect 119344 144916 119396 144968
rect 119712 144916 119764 144968
rect 3148 144848 3200 144900
rect 179696 144848 179748 144900
rect 112904 144780 112956 144832
rect 139768 144780 139820 144832
rect 175096 144780 175148 144832
rect 193496 144780 193548 144832
rect 112812 144712 112864 144764
rect 141792 144712 141844 144764
rect 173808 144712 173860 144764
rect 193680 144712 193732 144764
rect 580264 144848 580316 144900
rect 116492 144644 116544 144696
rect 148876 144644 148928 144696
rect 173992 144644 174044 144696
rect 197636 144644 197688 144696
rect 110236 144576 110288 144628
rect 142160 144576 142212 144628
rect 175188 144576 175240 144628
rect 199016 144576 199068 144628
rect 115664 144508 115716 144560
rect 148692 144508 148744 144560
rect 162952 144508 163004 144560
rect 197544 144508 197596 144560
rect 114284 144440 114336 144492
rect 146392 144440 146444 144492
rect 162308 144440 162360 144492
rect 196532 144440 196584 144492
rect 118516 144372 118568 144424
rect 151084 144372 151136 144424
rect 162492 144372 162544 144424
rect 196440 144372 196492 144424
rect 119712 144304 119764 144356
rect 152556 144304 152608 144356
rect 168012 144304 168064 144356
rect 202052 144304 202104 144356
rect 105360 144236 105412 144288
rect 166724 144236 166776 144288
rect 207848 144236 207900 144288
rect 117136 144168 117188 144220
rect 178040 144168 178092 144220
rect 179052 144168 179104 144220
rect 194784 144168 194836 144220
rect 116676 144100 116728 144152
rect 131672 144100 131724 144152
rect 177764 144100 177816 144152
rect 192852 144100 192904 144152
rect 116216 144032 116268 144084
rect 128360 144032 128412 144084
rect 139768 143692 139820 143744
rect 140412 143692 140464 143744
rect 191840 143692 191892 143744
rect 95792 143624 95844 143676
rect 164424 143624 164476 143676
rect 196348 143624 196400 143676
rect 196624 143624 196676 143676
rect 580540 143624 580592 143676
rect 134800 143556 134852 143608
rect 580448 143556 580500 143608
rect 115296 143488 115348 143540
rect 128544 143488 128596 143540
rect 188896 143488 188948 143540
rect 196256 143488 196308 143540
rect 112628 143420 112680 143472
rect 119896 143420 119948 143472
rect 120080 143420 120132 143472
rect 121368 143420 121420 143472
rect 121460 143420 121512 143472
rect 122196 143420 122248 143472
rect 181352 143420 181404 143472
rect 190644 143420 190696 143472
rect 115388 143352 115440 143404
rect 135996 143352 136048 143404
rect 185492 143352 185544 143404
rect 196164 143352 196216 143404
rect 115572 143284 115624 143336
rect 138480 143284 138532 143336
rect 183468 143284 183520 143336
rect 195060 143284 195112 143336
rect 119896 143216 119948 143268
rect 126980 143216 127032 143268
rect 127072 143216 127124 143268
rect 143632 143216 143684 143268
rect 184664 143216 184716 143268
rect 197820 143216 197872 143268
rect 116952 143148 117004 143200
rect 141240 143148 141292 143200
rect 159824 143148 159876 143200
rect 173808 143148 173860 143200
rect 178868 143148 178920 143200
rect 192208 143148 192260 143200
rect 98000 143080 98052 143132
rect 116860 143080 116912 143132
rect 117044 143080 117096 143132
rect 146760 143080 146812 143132
rect 168932 143080 168984 143132
rect 192668 143080 192720 143132
rect 110420 143012 110472 143064
rect 111616 143012 111668 143064
rect 142620 143012 142672 143064
rect 162308 143012 162360 143064
rect 185676 143012 185728 143064
rect 211252 143012 211304 143064
rect 82820 142944 82872 142996
rect 115296 142944 115348 142996
rect 115756 142944 115808 142996
rect 147680 142944 147732 142996
rect 166448 142944 166500 142996
rect 192116 142944 192168 142996
rect 213092 142944 213144 142996
rect 97356 142876 97408 142928
rect 137100 142876 137152 142928
rect 169668 142876 169720 142928
rect 196348 142876 196400 142928
rect 44180 142808 44232 142860
rect 110420 142808 110472 142860
rect 115112 142808 115164 142860
rect 148324 142808 148376 142860
rect 158628 142808 158680 142860
rect 191196 142808 191248 142860
rect 197820 142808 197872 142860
rect 198372 142808 198424 142860
rect 329840 142808 329892 142860
rect 116860 142740 116912 142792
rect 126060 142740 126112 142792
rect 120908 142672 120960 142724
rect 127072 142672 127124 142724
rect 186044 142604 186096 142656
rect 186228 142604 186280 142656
rect 179328 142468 179380 142520
rect 187608 142468 187660 142520
rect 176384 142400 176436 142452
rect 189632 142400 189684 142452
rect 190000 142400 190052 142452
rect 149980 142332 150032 142384
rect 188988 142332 189040 142384
rect 144920 142264 144972 142316
rect 145380 142264 145432 142316
rect 518900 142264 518952 142316
rect 120632 142196 120684 142248
rect 122840 142196 122892 142248
rect 143540 142196 143592 142248
rect 150900 142196 150952 142248
rect 161388 142196 161440 142248
rect 168840 142196 168892 142248
rect 187424 142196 187476 142248
rect 580264 142196 580316 142248
rect 97908 142128 97960 142180
rect 113272 142128 113324 142180
rect 118608 142128 118660 142180
rect 123668 142128 123720 142180
rect 148968 142128 149020 142180
rect 580724 142128 580776 142180
rect 117228 142060 117280 142112
rect 119804 142060 119856 142112
rect 183008 142060 183060 142112
rect 197452 142060 197504 142112
rect 544384 142060 544436 142112
rect 580172 142060 580224 142112
rect 116584 141924 116636 141976
rect 126244 141924 126296 141976
rect 143540 141992 143592 142044
rect 180064 141924 180116 141976
rect 196164 141924 196216 141976
rect 112904 141856 112956 141908
rect 127808 141856 127860 141908
rect 173164 141856 173216 141908
rect 185584 141856 185636 141908
rect 187608 141856 187660 141908
rect 198924 141856 198976 141908
rect 113272 141788 113324 141840
rect 113916 141788 113968 141840
rect 144276 141788 144328 141840
rect 174636 141788 174688 141840
rect 194876 141788 194928 141840
rect 117044 141720 117096 141772
rect 148600 141720 148652 141772
rect 165344 141720 165396 141772
rect 199200 141720 199252 141772
rect 118332 141652 118384 141704
rect 152004 141652 152056 141704
rect 153016 141652 153068 141704
rect 155592 141652 155644 141704
rect 189632 141652 189684 141704
rect 115572 141584 115624 141636
rect 149152 141584 149204 141636
rect 153108 141584 153160 141636
rect 188896 141584 188948 141636
rect 98644 141516 98696 141568
rect 158444 141516 158496 141568
rect 163964 141516 164016 141568
rect 197912 141516 197964 141568
rect 198924 141516 198976 141568
rect 213184 141516 213236 141568
rect 97264 141448 97316 141500
rect 138572 141448 138624 141500
rect 154028 141448 154080 141500
rect 218520 141448 218572 141500
rect 3608 141380 3660 141432
rect 113640 141380 113692 141432
rect 119344 141380 119396 141432
rect 133696 141380 133748 141432
rect 141240 141380 141292 141432
rect 580356 141380 580408 141432
rect 171784 141312 171836 141364
rect 186412 141312 186464 141364
rect 119252 141244 119304 141296
rect 126336 141244 126388 141296
rect 181904 141244 181956 141296
rect 196624 141244 196676 141296
rect 174728 141176 174780 141228
rect 190736 141176 190788 141228
rect 185584 141108 185636 141160
rect 192208 141108 192260 141160
rect 113180 140836 113232 140888
rect 117228 140836 117280 140888
rect 108120 140768 108172 140820
rect 153016 140836 153068 140888
rect 211804 140836 211856 140888
rect 174636 140768 174688 140820
rect 179420 140768 179472 140820
rect 179880 140768 179932 140820
rect 180800 140768 180852 140820
rect 181536 140768 181588 140820
rect 187700 140768 187752 140820
rect 188252 140768 188304 140820
rect 119896 140700 119948 140752
rect 124312 140700 124364 140752
rect 168840 140700 168892 140752
rect 193404 140700 193456 140752
rect 2780 140632 2832 140684
rect 4896 140632 4948 140684
rect 115204 140632 115256 140684
rect 126428 140632 126480 140684
rect 182824 140632 182876 140684
rect 183100 140632 183152 140684
rect 187332 140632 187384 140684
rect 193772 140632 193824 140684
rect 120816 140564 120868 140616
rect 134340 140564 134392 140616
rect 182916 140564 182968 140616
rect 192484 140564 192536 140616
rect 115388 140496 115440 140548
rect 131672 140496 131724 140548
rect 176568 140496 176620 140548
rect 186320 140496 186372 140548
rect 112352 140428 112404 140480
rect 131948 140428 132000 140480
rect 177856 140428 177908 140480
rect 189816 140496 189868 140548
rect 187792 140428 187844 140480
rect 188712 140428 188764 140480
rect 115296 140360 115348 140412
rect 144184 140360 144236 140412
rect 178960 140360 179012 140412
rect 193496 140360 193548 140412
rect 119712 140292 119764 140344
rect 150072 140292 150124 140344
rect 178684 140292 178736 140344
rect 197820 140292 197872 140344
rect 112536 140224 112588 140276
rect 142804 140224 142856 140276
rect 172060 140224 172112 140276
rect 198096 140224 198148 140276
rect 112628 140156 112680 140208
rect 145472 140156 145524 140208
rect 158536 140156 158588 140208
rect 193680 140156 193732 140208
rect 114008 140088 114060 140140
rect 130476 140088 130528 140140
rect 131028 140088 131080 140140
rect 194968 140088 195020 140140
rect 116860 139952 116912 140004
rect 150992 140020 151044 140072
rect 159640 140020 159692 140072
rect 186320 140020 186372 140072
rect 187332 140020 187384 140072
rect 193404 140020 193456 140072
rect 492680 140020 492732 140072
rect 190552 139952 190604 140004
rect 113916 139884 113968 139936
rect 124864 139884 124916 139936
rect 185676 139884 185728 139936
rect 191196 139884 191248 139936
rect 185768 139816 185820 139868
rect 192576 139816 192628 139868
rect 133696 139476 133748 139528
rect 288440 139476 288492 139528
rect 4804 139408 4856 139460
rect 182548 139408 182600 139460
rect 188160 139340 188212 139392
rect 189908 139340 189960 139392
rect 111248 139272 111300 139324
rect 123208 139272 123260 139324
rect 186412 139272 186464 139324
rect 194048 139272 194100 139324
rect 192760 138796 192812 138848
rect 200856 138796 200908 138848
rect 189908 138728 189960 138780
rect 197452 138728 197504 138780
rect 188988 138660 189040 138712
rect 512000 138660 512052 138712
rect 195428 137640 195480 137692
rect 199568 137640 199620 137692
rect 191380 137300 191432 137352
rect 203708 137300 203760 137352
rect 108212 137232 108264 137284
rect 120172 137232 120224 137284
rect 190000 137232 190052 137284
rect 416780 137232 416832 137284
rect 3516 136552 3568 136604
rect 104072 136552 104124 136604
rect 188896 133832 188948 133884
rect 188896 133628 188948 133680
rect 196716 133152 196768 133204
rect 216128 133152 216180 133204
rect 216128 132472 216180 132524
rect 579804 132472 579856 132524
rect 3332 132404 3384 132456
rect 105360 132404 105412 132456
rect 3424 127576 3476 127628
rect 117964 127576 118016 127628
rect 3424 122816 3476 122868
rect 117872 122816 117924 122868
rect 3332 120028 3384 120080
rect 95792 120028 95844 120080
rect 3424 116560 3476 116612
rect 120632 116560 120684 116612
rect 3332 111800 3384 111852
rect 116952 111800 117004 111852
rect 116492 110576 116544 110628
rect 120632 110576 120684 110628
rect 3056 108944 3108 108996
rect 100760 108944 100812 108996
rect 101312 108944 101364 108996
rect 100760 108264 100812 108316
rect 111156 108264 111208 108316
rect 200948 107652 201000 107704
rect 580172 107652 580224 107704
rect 2964 104796 3016 104848
rect 110420 104796 110472 104848
rect 110972 104796 111024 104848
rect 110420 104116 110472 104168
rect 119160 104116 119212 104168
rect 2872 99356 2924 99408
rect 105360 99356 105412 99408
rect 111616 95888 111668 95940
rect 119252 95888 119304 95940
rect 2964 95208 3016 95260
rect 116400 95208 116452 95260
rect 112260 94732 112312 94784
rect 115020 94732 115072 94784
rect 110972 93100 111024 93152
rect 120724 93100 120776 93152
rect 3056 91060 3108 91112
rect 97172 91060 97224 91112
rect 189724 88340 189776 88392
rect 189908 88340 189960 88392
rect 3516 88272 3568 88324
rect 108120 88272 108172 88324
rect 189540 86708 189592 86760
rect 190184 86708 190236 86760
rect 189356 86572 189408 86624
rect 189540 86572 189592 86624
rect 189172 86436 189224 86488
rect 189356 86436 189408 86488
rect 189080 84872 189132 84924
rect 189724 84872 189776 84924
rect 97632 83172 97684 83224
rect 98644 83172 98696 83224
rect 3516 82832 3568 82884
rect 97632 82832 97684 82884
rect 111616 82084 111668 82136
rect 117412 82084 117464 82136
rect 104072 81472 104124 81524
rect 119712 81336 119764 81388
rect 121644 81336 121696 81388
rect 104072 81200 104124 81252
rect 113732 81064 113784 81116
rect 121552 81064 121604 81116
rect 116584 80860 116636 80912
rect 118516 80792 118568 80844
rect 95608 80656 95660 80708
rect 115112 80588 115164 80640
rect 119804 80656 119856 80708
rect 123760 80656 123812 80708
rect 123944 80656 123996 80708
rect 128912 80656 128964 80708
rect 131580 80656 131632 80708
rect 131672 80656 131724 80708
rect 121920 80588 121972 80640
rect 131948 80656 132000 80708
rect 124496 80452 124548 80504
rect 131672 80520 131724 80572
rect 132132 80656 132184 80708
rect 132224 80588 132276 80640
rect 132132 80452 132184 80504
rect 131580 80384 131632 80436
rect 131948 80384 132000 80436
rect 128176 80316 128228 80368
rect 129924 80180 129976 80232
rect 131856 80180 131908 80232
rect 131764 80112 131816 80164
rect 130108 80044 130160 80096
rect 131672 80044 131724 80096
rect 101680 79772 101732 79824
rect 131948 79976 132000 80028
rect 131672 79908 131724 79960
rect 132132 79908 132184 79960
rect 132546 79908 132598 79960
rect 132638 79908 132690 79960
rect 132914 79908 132966 79960
rect 133006 79908 133058 79960
rect 133190 79908 133242 79960
rect 133374 79908 133426 79960
rect 133834 79908 133886 79960
rect 133926 79908 133978 79960
rect 106004 79704 106056 79756
rect 131580 79772 131632 79824
rect 132868 79704 132920 79756
rect 3516 79636 3568 79688
rect 117688 79568 117740 79620
rect 126244 79568 126296 79620
rect 119344 79500 119396 79552
rect 127624 79500 127676 79552
rect 111156 79432 111208 79484
rect 130108 79432 130160 79484
rect 133144 79772 133196 79824
rect 133052 79636 133104 79688
rect 132960 79568 133012 79620
rect 134294 79840 134346 79892
rect 133880 79704 133932 79756
rect 134570 79840 134622 79892
rect 134662 79840 134714 79892
rect 134340 79704 134392 79756
rect 134616 79704 134668 79756
rect 135030 79908 135082 79960
rect 135122 79908 135174 79960
rect 135214 79908 135266 79960
rect 135306 79908 135358 79960
rect 136226 79908 136278 79960
rect 136502 79908 136554 79960
rect 137054 79908 137106 79960
rect 137514 79908 137566 79960
rect 137606 79908 137658 79960
rect 137698 79908 137750 79960
rect 137974 79908 138026 79960
rect 138158 79908 138210 79960
rect 138250 79908 138302 79960
rect 134846 79840 134898 79892
rect 134938 79840 134990 79892
rect 134708 79636 134760 79688
rect 133696 79568 133748 79620
rect 134248 79568 134300 79620
rect 134432 79568 134484 79620
rect 135168 79772 135220 79824
rect 135490 79840 135542 79892
rect 135950 79840 136002 79892
rect 136042 79840 136094 79892
rect 135076 79704 135128 79756
rect 135260 79704 135312 79756
rect 135536 79704 135588 79756
rect 136318 79840 136370 79892
rect 136088 79704 136140 79756
rect 136180 79704 136232 79756
rect 135996 79636 136048 79688
rect 136364 79636 136416 79688
rect 135812 79568 135864 79620
rect 136594 79840 136646 79892
rect 136686 79840 136738 79892
rect 136870 79840 136922 79892
rect 137238 79840 137290 79892
rect 137422 79840 137474 79892
rect 136548 79636 136600 79688
rect 136640 79636 136692 79688
rect 137100 79704 137152 79756
rect 136824 79636 136876 79688
rect 137560 79772 137612 79824
rect 138020 79772 138072 79824
rect 137652 79704 137704 79756
rect 138112 79636 138164 79688
rect 138388 79636 138440 79688
rect 137008 79568 137060 79620
rect 137284 79568 137336 79620
rect 137376 79568 137428 79620
rect 134892 79500 134944 79552
rect 136272 79500 136324 79552
rect 139170 79908 139222 79960
rect 139814 79908 139866 79960
rect 139906 79908 139958 79960
rect 139998 79908 140050 79960
rect 140182 79908 140234 79960
rect 140274 79908 140326 79960
rect 140458 79908 140510 79960
rect 140642 79908 140694 79960
rect 140734 79908 140786 79960
rect 138710 79840 138762 79892
rect 138802 79840 138854 79892
rect 138986 79840 139038 79892
rect 139078 79840 139130 79892
rect 138940 79704 138992 79756
rect 138756 79636 138808 79688
rect 139032 79636 139084 79688
rect 139216 79568 139268 79620
rect 138572 79500 138624 79552
rect 139446 79772 139498 79824
rect 139952 79772 140004 79824
rect 139860 79704 139912 79756
rect 139676 79636 139728 79688
rect 139400 79568 139452 79620
rect 139768 79568 139820 79620
rect 140412 79636 140464 79688
rect 140918 79908 140970 79960
rect 141010 79908 141062 79960
rect 141194 79908 141246 79960
rect 141378 79908 141430 79960
rect 141746 79908 141798 79960
rect 141838 79908 141890 79960
rect 142022 79908 142074 79960
rect 140780 79772 140832 79824
rect 140688 79704 140740 79756
rect 140596 79568 140648 79620
rect 141562 79840 141614 79892
rect 140964 79500 141016 79552
rect 141332 79636 141384 79688
rect 141746 79772 141798 79824
rect 141700 79568 141752 79620
rect 141976 79704 142028 79756
rect 142482 79908 142534 79960
rect 142206 79840 142258 79892
rect 142390 79840 142442 79892
rect 142068 79568 142120 79620
rect 142344 79500 142396 79552
rect 108212 79364 108264 79416
rect 134984 79364 135036 79416
rect 135352 79364 135404 79416
rect 136456 79364 136508 79416
rect 141884 79432 141936 79484
rect 142252 79432 142304 79484
rect 142528 79636 142580 79688
rect 142942 79908 142994 79960
rect 143218 79908 143270 79960
rect 143494 79908 143546 79960
rect 143586 79908 143638 79960
rect 142804 79568 142856 79620
rect 142528 79500 142580 79552
rect 143126 79840 143178 79892
rect 143080 79704 143132 79756
rect 143172 79704 143224 79756
rect 143402 79772 143454 79824
rect 143540 79636 143592 79688
rect 143356 79568 143408 79620
rect 143448 79568 143500 79620
rect 142896 79432 142948 79484
rect 143770 79908 143822 79960
rect 143954 79908 144006 79960
rect 144322 79908 144374 79960
rect 144414 79908 144466 79960
rect 144598 79908 144650 79960
rect 144690 79908 144742 79960
rect 144782 79908 144834 79960
rect 145242 79908 145294 79960
rect 145426 79908 145478 79960
rect 145518 79908 145570 79960
rect 145610 79908 145662 79960
rect 144046 79840 144098 79892
rect 144000 79636 144052 79688
rect 144276 79636 144328 79688
rect 144690 79772 144742 79824
rect 144552 79636 144604 79688
rect 144736 79636 144788 79688
rect 144966 79840 145018 79892
rect 145150 79840 145202 79892
rect 143908 79568 143960 79620
rect 144092 79568 144144 79620
rect 145380 79772 145432 79824
rect 145472 79704 145524 79756
rect 145564 79704 145616 79756
rect 145196 79636 145248 79688
rect 145886 79908 145938 79960
rect 145794 79840 145846 79892
rect 207572 81268 207624 81320
rect 191380 81132 191432 81184
rect 198096 81132 198148 81184
rect 188988 81064 189040 81116
rect 209136 81064 209188 81116
rect 202420 80996 202472 81048
rect 580172 81336 580224 81388
rect 204536 80928 204588 80980
rect 188988 80860 189040 80912
rect 219992 80860 220044 80912
rect 177856 80656 177908 80708
rect 178040 80656 178092 80708
rect 178408 80656 178460 80708
rect 196624 80792 196676 80844
rect 146070 79908 146122 79960
rect 146162 79908 146214 79960
rect 146346 79908 146398 79960
rect 146806 79908 146858 79960
rect 147358 79908 147410 79960
rect 147450 79908 147502 79960
rect 147542 79908 147594 79960
rect 148094 79908 148146 79960
rect 145932 79772 145984 79824
rect 146070 79772 146122 79824
rect 145840 79704 145892 79756
rect 145104 79568 145156 79620
rect 145288 79568 145340 79620
rect 146024 79568 146076 79620
rect 146438 79840 146490 79892
rect 146622 79840 146674 79892
rect 146484 79568 146536 79620
rect 146392 79500 146444 79552
rect 146898 79840 146950 79892
rect 146990 79840 147042 79892
rect 147174 79840 147226 79892
rect 147266 79840 147318 79892
rect 147634 79840 147686 79892
rect 147404 79772 147456 79824
rect 147496 79772 147548 79824
rect 146944 79636 146996 79688
rect 146852 79568 146904 79620
rect 147220 79704 147272 79756
rect 147312 79704 147364 79756
rect 147588 79704 147640 79756
rect 146760 79500 146812 79552
rect 147036 79500 147088 79552
rect 148554 79840 148606 79892
rect 148830 79908 148882 79960
rect 148922 79908 148974 79960
rect 149014 79908 149066 79960
rect 149474 79908 149526 79960
rect 149566 79908 149618 79960
rect 149658 79908 149710 79960
rect 150762 79908 150814 79960
rect 151038 79908 151090 79960
rect 151406 79908 151458 79960
rect 148968 79772 149020 79824
rect 149198 79772 149250 79824
rect 148876 79704 148928 79756
rect 148692 79636 148744 79688
rect 149750 79840 149802 79892
rect 149842 79840 149894 79892
rect 149934 79840 149986 79892
rect 150118 79840 150170 79892
rect 150302 79840 150354 79892
rect 149612 79704 149664 79756
rect 149704 79704 149756 79756
rect 149796 79704 149848 79756
rect 149520 79636 149572 79688
rect 149888 79636 149940 79688
rect 148784 79568 148836 79620
rect 149152 79568 149204 79620
rect 148140 79500 148192 79552
rect 149244 79500 149296 79552
rect 150670 79772 150722 79824
rect 151314 79840 151366 79892
rect 151590 79908 151642 79960
rect 151682 79908 151734 79960
rect 151866 79908 151918 79960
rect 151958 79908 152010 79960
rect 151498 79772 151550 79824
rect 151360 79568 151412 79620
rect 150716 79500 150768 79552
rect 150992 79500 151044 79552
rect 151544 79636 151596 79688
rect 152050 79840 152102 79892
rect 152142 79772 152194 79824
rect 151912 79704 151964 79756
rect 152004 79704 152056 79756
rect 152418 79908 152470 79960
rect 152970 79908 153022 79960
rect 153614 79908 153666 79960
rect 154258 79908 154310 79960
rect 154350 79908 154402 79960
rect 154442 79908 154494 79960
rect 154994 79908 155046 79960
rect 155178 79908 155230 79960
rect 155822 79908 155874 79960
rect 156190 79908 156242 79960
rect 156650 79908 156702 79960
rect 156926 79908 156978 79960
rect 157018 79908 157070 79960
rect 157110 79908 157162 79960
rect 157202 79908 157254 79960
rect 157386 79908 157438 79960
rect 157478 79908 157530 79960
rect 157662 79908 157714 79960
rect 152786 79840 152838 79892
rect 152464 79704 152516 79756
rect 152096 79636 152148 79688
rect 153246 79840 153298 79892
rect 153430 79840 153482 79892
rect 153062 79772 153114 79824
rect 152832 79636 152884 79688
rect 152188 79568 152240 79620
rect 153016 79568 153068 79620
rect 153292 79568 153344 79620
rect 153108 79500 153160 79552
rect 153200 79500 153252 79552
rect 153568 79636 153620 79688
rect 153890 79772 153942 79824
rect 154074 79772 154126 79824
rect 154212 79772 154264 79824
rect 154120 79636 154172 79688
rect 154442 79772 154494 79824
rect 154948 79704 155000 79756
rect 155270 79840 155322 79892
rect 155638 79840 155690 79892
rect 155316 79704 155368 79756
rect 153844 79568 153896 79620
rect 155132 79636 155184 79688
rect 155914 79840 155966 79892
rect 156006 79840 156058 79892
rect 155776 79704 155828 79756
rect 156236 79772 156288 79824
rect 156144 79704 156196 79756
rect 155868 79636 155920 79688
rect 153476 79500 153528 79552
rect 155960 79568 156012 79620
rect 143816 79432 143868 79484
rect 150256 79432 150308 79484
rect 150532 79432 150584 79484
rect 154672 79432 154724 79484
rect 104164 79296 104216 79348
rect 104716 79296 104768 79348
rect 110236 79296 110288 79348
rect 141608 79296 141660 79348
rect 149428 79364 149480 79416
rect 118056 79228 118108 79280
rect 149244 79228 149296 79280
rect 104532 79160 104584 79212
rect 104716 79160 104768 79212
rect 113088 79160 113140 79212
rect 145564 79160 145616 79212
rect 113916 79092 113968 79144
rect 146392 79092 146444 79144
rect 102876 79024 102928 79076
rect 135352 79024 135404 79076
rect 136456 79024 136508 79076
rect 136732 79024 136784 79076
rect 149428 79024 149480 79076
rect 112352 78956 112404 79008
rect 145932 78956 145984 79008
rect 154672 79228 154724 79280
rect 156420 79500 156472 79552
rect 156742 79840 156794 79892
rect 156834 79840 156886 79892
rect 157018 79772 157070 79824
rect 157340 79704 157392 79756
rect 156972 79636 157024 79688
rect 157064 79636 157116 79688
rect 157156 79636 157208 79688
rect 156880 79568 156932 79620
rect 157570 79840 157622 79892
rect 157708 79772 157760 79824
rect 157524 79704 157576 79756
rect 157616 79636 157668 79688
rect 158214 79908 158266 79960
rect 158306 79908 158358 79960
rect 157892 79568 157944 79620
rect 158490 79840 158542 79892
rect 158582 79840 158634 79892
rect 158950 79840 159002 79892
rect 158536 79704 158588 79756
rect 156788 79500 156840 79552
rect 158260 79500 158312 79552
rect 158904 79364 158956 79416
rect 159134 79908 159186 79960
rect 159226 79908 159278 79960
rect 159318 79908 159370 79960
rect 159502 79908 159554 79960
rect 159272 79636 159324 79688
rect 159180 79568 159232 79620
rect 159870 79908 159922 79960
rect 160238 79908 160290 79960
rect 160422 79908 160474 79960
rect 160698 79908 160750 79960
rect 160974 79908 161026 79960
rect 161618 79908 161670 79960
rect 161710 79908 161762 79960
rect 161894 79908 161946 79960
rect 162078 79908 162130 79960
rect 162170 79908 162222 79960
rect 162262 79908 162314 79960
rect 159548 79704 159600 79756
rect 159962 79840 160014 79892
rect 160054 79840 160106 79892
rect 160008 79704 160060 79756
rect 160100 79636 160152 79688
rect 159824 79568 159876 79620
rect 160514 79840 160566 79892
rect 160652 79772 160704 79824
rect 160560 79704 160612 79756
rect 161158 79840 161210 79892
rect 161250 79772 161302 79824
rect 160284 79636 160336 79688
rect 160928 79636 160980 79688
rect 161204 79636 161256 79688
rect 161526 79772 161578 79824
rect 161480 79636 161532 79688
rect 160744 79500 160796 79552
rect 161112 79500 161164 79552
rect 161940 79772 161992 79824
rect 162630 79840 162682 79892
rect 161756 79704 161808 79756
rect 162216 79704 162268 79756
rect 162032 79636 162084 79688
rect 162998 79908 163050 79960
rect 163458 79908 163510 79960
rect 164102 79908 164154 79960
rect 164562 79908 164614 79960
rect 162814 79772 162866 79824
rect 163182 79840 163234 79892
rect 162860 79636 162912 79688
rect 162952 79636 163004 79688
rect 161664 79568 161716 79620
rect 162676 79568 162728 79620
rect 163228 79568 163280 79620
rect 161940 79500 161992 79552
rect 160376 79432 160428 79484
rect 163550 79840 163602 79892
rect 163826 79772 163878 79824
rect 163918 79772 163970 79824
rect 163872 79636 163924 79688
rect 163964 79568 164016 79620
rect 164148 79568 164200 79620
rect 163688 79500 163740 79552
rect 164470 79840 164522 79892
rect 164838 79908 164890 79960
rect 165114 79908 165166 79960
rect 165206 79908 165258 79960
rect 165298 79908 165350 79960
rect 165390 79908 165442 79960
rect 165942 79908 165994 79960
rect 166126 79908 166178 79960
rect 166402 79908 166454 79960
rect 166678 79908 166730 79960
rect 166770 79908 166822 79960
rect 166954 79908 167006 79960
rect 164608 79704 164660 79756
rect 165252 79704 165304 79756
rect 165344 79704 165396 79756
rect 164792 79636 164844 79688
rect 165160 79636 165212 79688
rect 165758 79840 165810 79892
rect 165850 79840 165902 79892
rect 165896 79704 165948 79756
rect 166310 79840 166362 79892
rect 166264 79704 166316 79756
rect 165804 79636 165856 79688
rect 165988 79636 166040 79688
rect 166494 79772 166546 79824
rect 166540 79636 166592 79688
rect 165436 79568 165488 79620
rect 166448 79568 166500 79620
rect 166724 79568 166776 79620
rect 166816 79568 166868 79620
rect 164884 79500 164936 79552
rect 166356 79500 166408 79552
rect 164056 79432 164108 79484
rect 167506 79908 167558 79960
rect 167598 79908 167650 79960
rect 178592 80588 178644 80640
rect 211436 80724 211488 80776
rect 178040 80520 178092 80572
rect 207664 80656 207716 80708
rect 187700 80588 187752 80640
rect 189080 80588 189132 80640
rect 188344 80520 188396 80572
rect 194048 80520 194100 80572
rect 184204 80452 184256 80504
rect 191380 80452 191432 80504
rect 167230 79840 167282 79892
rect 177856 80384 177908 80436
rect 177764 80316 177816 80368
rect 178316 80248 178368 80300
rect 178408 80180 178460 80232
rect 169162 79908 169214 79960
rect 170726 79908 170778 79960
rect 168794 79840 168846 79892
rect 168978 79840 169030 79892
rect 168426 79772 168478 79824
rect 168518 79772 168570 79824
rect 167828 79500 167880 79552
rect 168656 79636 168708 79688
rect 169024 79636 169076 79688
rect 168564 79500 168616 79552
rect 168748 79500 168800 79552
rect 168472 79432 168524 79484
rect 169622 79840 169674 79892
rect 169990 79840 170042 79892
rect 170082 79840 170134 79892
rect 169438 79772 169490 79824
rect 169944 79704 169996 79756
rect 170036 79704 170088 79756
rect 169484 79500 169536 79552
rect 170956 79500 171008 79552
rect 171370 79840 171422 79892
rect 171738 79840 171790 79892
rect 171830 79840 171882 79892
rect 171554 79772 171606 79824
rect 171508 79636 171560 79688
rect 171692 79636 171744 79688
rect 171784 79636 171836 79688
rect 171876 79500 171928 79552
rect 170404 79432 170456 79484
rect 172198 79908 172250 79960
rect 172566 79908 172618 79960
rect 172290 79840 172342 79892
rect 172382 79840 172434 79892
rect 172566 79772 172618 79824
rect 172842 79908 172894 79960
rect 172934 79908 172986 79960
rect 172750 79840 172802 79892
rect 172796 79636 172848 79688
rect 172704 79568 172756 79620
rect 172980 79568 173032 79620
rect 173486 79908 173538 79960
rect 173578 79908 173630 79960
rect 173670 79908 173722 79960
rect 173854 79908 173906 79960
rect 174038 79908 174090 79960
rect 174222 79908 174274 79960
rect 174314 79908 174366 79960
rect 174590 79908 174642 79960
rect 173302 79840 173354 79892
rect 173394 79840 173446 79892
rect 173348 79636 173400 79688
rect 173440 79636 173492 79688
rect 174774 79908 174826 79960
rect 174866 79908 174918 79960
rect 175142 79908 175194 79960
rect 175602 79908 175654 79960
rect 175786 79908 175838 79960
rect 176062 79908 176114 79960
rect 176338 79908 176390 79960
rect 176522 79908 176574 79960
rect 175050 79840 175102 79892
rect 174038 79772 174090 79824
rect 174268 79772 174320 79824
rect 174636 79772 174688 79824
rect 174728 79772 174780 79824
rect 173716 79704 173768 79756
rect 173900 79704 173952 79756
rect 175694 79840 175746 79892
rect 175188 79636 175240 79688
rect 173256 79568 173308 79620
rect 173624 79568 173676 79620
rect 175096 79568 175148 79620
rect 175648 79704 175700 79756
rect 176154 79840 176206 79892
rect 176016 79772 176068 79824
rect 176430 79772 176482 79824
rect 176108 79704 176160 79756
rect 176292 79636 176344 79688
rect 176798 79840 176850 79892
rect 178040 80112 178092 80164
rect 178132 80112 178184 80164
rect 181168 80112 181220 80164
rect 177764 80044 177816 80096
rect 179604 80044 179656 80096
rect 191380 80044 191432 80096
rect 198188 80044 198240 80096
rect 177948 79976 178000 80028
rect 178132 79976 178184 80028
rect 184940 79976 184992 80028
rect 215668 79976 215720 80028
rect 176982 79908 177034 79960
rect 177166 79908 177218 79960
rect 176936 79772 176988 79824
rect 177258 79840 177310 79892
rect 177350 79840 177402 79892
rect 178500 79840 178552 79892
rect 182916 79840 182968 79892
rect 194048 79840 194100 79892
rect 200856 79840 200908 79892
rect 177672 79772 177724 79824
rect 177304 79704 177356 79756
rect 189080 79636 189132 79688
rect 203064 79636 203116 79688
rect 175832 79568 175884 79620
rect 176568 79568 176620 79620
rect 181444 79568 181496 79620
rect 580816 79568 580868 79620
rect 172520 79500 172572 79552
rect 173164 79500 173216 79552
rect 188988 79500 189040 79552
rect 172060 79432 172112 79484
rect 172336 79432 172388 79484
rect 173900 79432 173952 79484
rect 214656 79432 214708 79484
rect 159364 79364 159416 79416
rect 167184 79364 167236 79416
rect 167276 79364 167328 79416
rect 187700 79364 187752 79416
rect 160468 79296 160520 79348
rect 160560 79296 160612 79348
rect 195244 79296 195296 79348
rect 167184 79228 167236 79280
rect 159364 79160 159416 79212
rect 171968 79228 172020 79280
rect 210608 79228 210660 79280
rect 154580 79092 154632 79144
rect 155592 79092 155644 79144
rect 181444 79160 181496 79212
rect 181536 79160 181588 79212
rect 215484 79160 215536 79212
rect 175648 79092 175700 79144
rect 179604 79092 179656 79144
rect 215760 79092 215812 79144
rect 170496 79024 170548 79076
rect 212816 79024 212868 79076
rect 174268 78956 174320 79008
rect 219624 78956 219676 79008
rect 129188 78888 129240 78940
rect 138756 78888 138808 78940
rect 160928 78888 160980 78940
rect 210516 78888 210568 78940
rect 95976 78820 96028 78872
rect 152280 78820 152332 78872
rect 161756 78820 161808 78872
rect 217140 78820 217192 78872
rect 131028 78752 131080 78804
rect 141516 78752 141568 78804
rect 157432 78752 157484 78804
rect 158168 78752 158220 78804
rect 175740 78752 175792 78804
rect 180248 78752 180300 78804
rect 181168 78752 181220 78804
rect 212724 78752 212776 78804
rect 135352 78684 135404 78736
rect 135812 78684 135864 78736
rect 136732 78684 136784 78736
rect 137008 78684 137060 78736
rect 141240 78684 141292 78736
rect 141884 78684 141936 78736
rect 142712 78684 142764 78736
rect 142988 78684 143040 78736
rect 153292 78684 153344 78736
rect 154396 78684 154448 78736
rect 171232 78684 171284 78736
rect 171508 78684 171560 78736
rect 172244 78684 172296 78736
rect 180616 78684 180668 78736
rect 96528 78616 96580 78668
rect 132040 78616 132092 78668
rect 132132 78616 132184 78668
rect 143356 78616 143408 78668
rect 145288 78616 145340 78668
rect 145472 78616 145524 78668
rect 154028 78616 154080 78668
rect 154488 78616 154540 78668
rect 159548 78616 159600 78668
rect 121828 78548 121880 78600
rect 136456 78548 136508 78600
rect 170588 78616 170640 78668
rect 173900 78616 173952 78668
rect 177580 78616 177632 78668
rect 219900 78616 219952 78668
rect 169484 78548 169536 78600
rect 170404 78548 170456 78600
rect 171508 78548 171560 78600
rect 172520 78548 172572 78600
rect 173624 78548 173676 78600
rect 178040 78548 178092 78600
rect 189540 78548 189592 78600
rect 105912 78480 105964 78532
rect 139952 78480 140004 78532
rect 142988 78480 143040 78532
rect 151912 78480 151964 78532
rect 165436 78480 165488 78532
rect 103980 78412 104032 78464
rect 136640 78412 136692 78464
rect 165620 78412 165672 78464
rect 166172 78412 166224 78464
rect 167552 78480 167604 78532
rect 169576 78480 169628 78532
rect 170588 78480 170640 78532
rect 171048 78480 171100 78532
rect 214104 78480 214156 78532
rect 171324 78412 171376 78464
rect 206284 78412 206336 78464
rect 99748 78344 99800 78396
rect 131580 78344 131632 78396
rect 130384 78276 130436 78328
rect 132132 78276 132184 78328
rect 108304 78208 108356 78260
rect 139400 78344 139452 78396
rect 169024 78344 169076 78396
rect 136640 78276 136692 78328
rect 142068 78276 142120 78328
rect 146300 78276 146352 78328
rect 155132 78276 155184 78328
rect 177212 78344 177264 78396
rect 211712 78344 211764 78396
rect 203616 78276 203668 78328
rect 138848 78208 138900 78260
rect 146116 78208 146168 78260
rect 152372 78208 152424 78260
rect 152924 78208 152976 78260
rect 164424 78208 164476 78260
rect 165252 78208 165304 78260
rect 175464 78208 175516 78260
rect 189724 78208 189776 78260
rect 102784 78140 102836 78192
rect 129924 78140 129976 78192
rect 132868 78140 132920 78192
rect 138388 78140 138440 78192
rect 140044 78140 140096 78192
rect 150716 78140 150768 78192
rect 157892 78140 157944 78192
rect 101772 78072 101824 78124
rect 131028 78072 131080 78124
rect 132040 78072 132092 78124
rect 134524 78072 134576 78124
rect 135904 78072 135956 78124
rect 143264 78072 143316 78124
rect 145932 78072 145984 78124
rect 158536 78072 158588 78124
rect 103888 78004 103940 78056
rect 137468 78004 137520 78056
rect 140412 78004 140464 78056
rect 151728 78004 151780 78056
rect 181720 78140 181772 78192
rect 196532 78140 196584 78192
rect 173716 78072 173768 78124
rect 179696 78072 179748 78124
rect 181536 78072 181588 78124
rect 196440 78072 196492 78124
rect 167552 78004 167604 78056
rect 168932 78004 168984 78056
rect 120816 77936 120868 77988
rect 134064 77936 134116 77988
rect 105728 77868 105780 77920
rect 128176 77868 128228 77920
rect 101588 77800 101640 77852
rect 135628 77868 135680 77920
rect 137008 77868 137060 77920
rect 146024 77936 146076 77988
rect 157524 77936 157576 77988
rect 169668 77936 169720 77988
rect 172796 78004 172848 78056
rect 181260 78004 181312 78056
rect 181812 78004 181864 78056
rect 197912 78004 197964 78056
rect 177856 77936 177908 77988
rect 180340 77936 180392 77988
rect 202236 77936 202288 77988
rect 157984 77868 158036 77920
rect 166816 77868 166868 77920
rect 174176 77868 174228 77920
rect 174452 77868 174504 77920
rect 181352 77868 181404 77920
rect 193772 77868 193824 77920
rect 135720 77800 135772 77852
rect 148876 77800 148928 77852
rect 171600 77800 171652 77852
rect 181444 77800 181496 77852
rect 103060 77732 103112 77784
rect 134984 77732 135036 77784
rect 166632 77732 166684 77784
rect 171876 77732 171928 77784
rect 174636 77732 174688 77784
rect 190000 77732 190052 77784
rect 136824 77664 136876 77716
rect 144552 77664 144604 77716
rect 166724 77664 166776 77716
rect 173900 77664 173952 77716
rect 142896 77596 142948 77648
rect 154120 77596 154172 77648
rect 155500 77596 155552 77648
rect 173164 77596 173216 77648
rect 173808 77596 173860 77648
rect 210424 77596 210476 77648
rect 159088 77460 159140 77512
rect 162584 77460 162636 77512
rect 169116 77460 169168 77512
rect 170680 77460 170732 77512
rect 164608 77392 164660 77444
rect 165528 77392 165580 77444
rect 168840 77324 168892 77376
rect 174636 77324 174688 77376
rect 136088 77256 136140 77308
rect 138940 77256 138992 77308
rect 97172 77188 97224 77240
rect 116400 77188 116452 77240
rect 156696 77188 156748 77240
rect 163504 77188 163556 77240
rect 164148 77188 164200 77240
rect 165896 77188 165948 77240
rect 166172 77188 166224 77240
rect 177672 77188 177724 77240
rect 201684 77188 201736 77240
rect 168472 77120 168524 77172
rect 177304 77120 177356 77172
rect 191196 77120 191248 77172
rect 107016 77052 107068 77104
rect 139492 77052 139544 77104
rect 147956 77052 148008 77104
rect 149980 77052 150032 77104
rect 200948 77052 201000 77104
rect 116952 76984 117004 77036
rect 167276 76984 167328 77036
rect 173348 76984 173400 77036
rect 209044 76984 209096 77036
rect 117872 76916 117924 76968
rect 2872 76848 2924 76900
rect 120080 76848 120132 76900
rect 121276 76848 121328 76900
rect 153200 76848 153252 76900
rect 102968 76780 103020 76832
rect 133236 76780 133288 76832
rect 134340 76780 134392 76832
rect 134984 76780 135036 76832
rect 146668 76780 146720 76832
rect 147036 76780 147088 76832
rect 117412 76712 117464 76764
rect 148968 76712 149020 76764
rect 109500 76644 109552 76696
rect 136824 76644 136876 76696
rect 148232 76644 148284 76696
rect 148600 76644 148652 76696
rect 150716 76644 150768 76696
rect 150900 76644 150952 76696
rect 119160 76576 119212 76628
rect 144092 76576 144144 76628
rect 146760 76576 146812 76628
rect 147036 76576 147088 76628
rect 156696 76916 156748 76968
rect 159272 76916 159324 76968
rect 193956 76916 194008 76968
rect 160100 76848 160152 76900
rect 164148 76848 164200 76900
rect 178500 76848 178552 76900
rect 211896 76848 211948 76900
rect 156788 76780 156840 76832
rect 190828 76780 190880 76832
rect 168472 76712 168524 76764
rect 200304 76712 200356 76764
rect 154948 76644 155000 76696
rect 155776 76644 155828 76696
rect 156788 76644 156840 76696
rect 157156 76644 157208 76696
rect 157800 76644 157852 76696
rect 158444 76644 158496 76696
rect 160100 76644 160152 76696
rect 160376 76644 160428 76696
rect 165712 76644 165764 76696
rect 199384 76644 199436 76696
rect 182916 76576 182968 76628
rect 104532 76508 104584 76560
rect 136272 76508 136324 76560
rect 136824 76508 136876 76560
rect 137652 76508 137704 76560
rect 138296 76508 138348 76560
rect 138480 76508 138532 76560
rect 140780 76508 140832 76560
rect 141332 76508 141384 76560
rect 141516 76508 141568 76560
rect 143080 76508 143132 76560
rect 148140 76508 148192 76560
rect 148600 76508 148652 76560
rect 150900 76508 150952 76560
rect 151636 76508 151688 76560
rect 155960 76508 156012 76560
rect 196440 76508 196492 76560
rect 131856 76440 131908 76492
rect 150808 76440 150860 76492
rect 155132 76440 155184 76492
rect 155868 76440 155920 76492
rect 158536 76440 158588 76492
rect 217232 76440 217284 76492
rect 120080 76372 120132 76424
rect 121000 76372 121052 76424
rect 153936 76372 153988 76424
rect 171324 76372 171376 76424
rect 171784 76372 171836 76424
rect 138020 76304 138072 76356
rect 138480 76304 138532 76356
rect 146760 76304 146812 76356
rect 147312 76304 147364 76356
rect 175004 76304 175056 76356
rect 214564 76372 214616 76424
rect 140872 76168 140924 76220
rect 141148 76168 141200 76220
rect 134064 76100 134116 76152
rect 134524 76100 134576 76152
rect 156236 76100 156288 76152
rect 156972 76100 157024 76152
rect 163688 76100 163740 76152
rect 165068 76100 165120 76152
rect 137192 76032 137244 76084
rect 138572 76032 138624 76084
rect 146852 75964 146904 76016
rect 147220 75964 147272 76016
rect 126336 75896 126388 75948
rect 132040 75896 132092 75948
rect 143540 75896 143592 75948
rect 152372 75896 152424 75948
rect 155224 75896 155276 75948
rect 158260 75896 158312 75948
rect 162676 75896 162728 75948
rect 170864 75896 170916 75948
rect 172520 75896 172572 75948
rect 172980 75896 173032 75948
rect 173992 75896 174044 75948
rect 174820 75896 174872 75948
rect 99656 75828 99708 75880
rect 102784 75828 102836 75880
rect 124496 75828 124548 75880
rect 135720 75828 135772 75880
rect 138204 75828 138256 75880
rect 145656 75828 145708 75880
rect 157340 75828 157392 75880
rect 157616 75828 157668 75880
rect 174268 75828 174320 75880
rect 175096 75828 175148 75880
rect 196440 75828 196492 75880
rect 217324 75828 217376 75880
rect 97448 75760 97500 75812
rect 130844 75760 130896 75812
rect 133328 75760 133380 75812
rect 137928 75760 137980 75812
rect 153108 75760 153160 75812
rect 167092 75760 167144 75812
rect 174360 75760 174412 75812
rect 192300 75760 192352 75812
rect 147588 75692 147640 75744
rect 162124 75692 162176 75744
rect 171048 75692 171100 75744
rect 175832 75692 175884 75744
rect 214288 75692 214340 75744
rect 114376 75624 114428 75676
rect 142068 75624 142120 75676
rect 156052 75624 156104 75676
rect 156880 75624 156932 75676
rect 157340 75624 157392 75676
rect 158076 75624 158128 75676
rect 160376 75624 160428 75676
rect 161204 75624 161256 75676
rect 162676 75624 162728 75676
rect 164976 75624 165028 75676
rect 199292 75624 199344 75676
rect 116768 75556 116820 75608
rect 117136 75556 117188 75608
rect 149152 75556 149204 75608
rect 181260 75556 181312 75608
rect 182088 75556 182140 75608
rect 214196 75556 214248 75608
rect 116308 75488 116360 75540
rect 148508 75488 148560 75540
rect 175372 75488 175424 75540
rect 175924 75488 175976 75540
rect 179696 75488 179748 75540
rect 205088 75488 205140 75540
rect 118240 75420 118292 75472
rect 140504 75420 140556 75472
rect 114468 75352 114520 75404
rect 142344 75420 142396 75472
rect 143080 75420 143132 75472
rect 146576 75420 146628 75472
rect 147404 75420 147456 75472
rect 148140 75420 148192 75472
rect 148416 75420 148468 75472
rect 158812 75420 158864 75472
rect 159088 75420 159140 75472
rect 175832 75420 175884 75472
rect 176476 75420 176528 75472
rect 198832 75420 198884 75472
rect 141056 75352 141108 75404
rect 142068 75352 142120 75404
rect 158720 75352 158772 75404
rect 159272 75352 159324 75404
rect 165804 75352 165856 75404
rect 166264 75352 166316 75404
rect 170220 75352 170272 75404
rect 192576 75352 192628 75404
rect 119528 75284 119580 75336
rect 138204 75284 138256 75336
rect 138664 75284 138716 75336
rect 143908 75284 143960 75336
rect 158812 75284 158864 75336
rect 159732 75284 159784 75336
rect 165712 75284 165764 75336
rect 166540 75284 166592 75336
rect 167000 75284 167052 75336
rect 168288 75284 168340 75336
rect 171692 75284 171744 75336
rect 171968 75284 172020 75336
rect 174452 75284 174504 75336
rect 192484 75284 192536 75336
rect 107660 75216 107712 75268
rect 126336 75216 126388 75268
rect 133052 75216 133104 75268
rect 133788 75216 133840 75268
rect 135536 75216 135588 75268
rect 135996 75216 136048 75268
rect 138572 75216 138624 75268
rect 139308 75216 139360 75268
rect 146852 75216 146904 75268
rect 147496 75216 147548 75268
rect 150440 75216 150492 75268
rect 151176 75216 151228 75268
rect 158720 75216 158772 75268
rect 158996 75216 159048 75268
rect 161572 75216 161624 75268
rect 162216 75216 162268 75268
rect 165896 75216 165948 75268
rect 166448 75216 166500 75268
rect 167184 75216 167236 75268
rect 167736 75216 167788 75268
rect 168472 75216 168524 75268
rect 169208 75216 169260 75268
rect 175280 75216 175332 75268
rect 176200 75216 176252 75268
rect 40040 75148 40092 75200
rect 117136 75148 117188 75200
rect 120080 75148 120132 75200
rect 167092 75148 167144 75200
rect 167276 75148 167328 75200
rect 168104 75148 168156 75200
rect 168196 75148 168248 75200
rect 177948 75148 178000 75200
rect 194508 75148 194560 75200
rect 269120 75148 269172 75200
rect 135628 75080 135680 75132
rect 136548 75080 136600 75132
rect 139584 75080 139636 75132
rect 140320 75080 140372 75132
rect 141056 75080 141108 75132
rect 141884 75080 141936 75132
rect 153752 75080 153804 75132
rect 216128 75080 216180 75132
rect 93676 74944 93728 74996
rect 141792 75012 141844 75064
rect 158996 75012 159048 75064
rect 160008 75012 160060 75064
rect 162860 75012 162912 75064
rect 163504 75012 163556 75064
rect 170588 75012 170640 75064
rect 214380 75012 214432 75064
rect 139584 74944 139636 74996
rect 140688 74944 140740 74996
rect 145564 74944 145616 74996
rect 146116 74944 146168 74996
rect 173072 74944 173124 74996
rect 193220 74944 193272 74996
rect 95700 74876 95752 74928
rect 145380 74876 145432 74928
rect 162584 74876 162636 74928
rect 181352 74876 181404 74928
rect 140504 74808 140556 74860
rect 147220 74808 147272 74860
rect 170036 74808 170088 74860
rect 172152 74808 172204 74860
rect 107016 74740 107068 74792
rect 107476 74740 107528 74792
rect 128912 74740 128964 74792
rect 137928 74740 137980 74792
rect 151820 74740 151872 74792
rect 154212 74740 154264 74792
rect 107476 74604 107528 74656
rect 107660 74604 107712 74656
rect 137284 74604 137336 74656
rect 142804 74604 142856 74656
rect 101864 74468 101916 74520
rect 106280 74468 106332 74520
rect 118148 74468 118200 74520
rect 140412 74468 140464 74520
rect 169484 74468 169536 74520
rect 193864 74468 193916 74520
rect 97632 74400 97684 74452
rect 157708 74400 157760 74452
rect 163320 74400 163372 74452
rect 216864 74400 216916 74452
rect 114008 74332 114060 74384
rect 143816 74332 143868 74384
rect 172060 74332 172112 74384
rect 215392 74332 215444 74384
rect 118424 74264 118476 74316
rect 152648 74264 152700 74316
rect 164608 74264 164660 74316
rect 200396 74264 200448 74316
rect 117228 74196 117280 74248
rect 150716 74196 150768 74248
rect 154672 74196 154724 74248
rect 155408 74196 155460 74248
rect 161480 74196 161532 74248
rect 162492 74196 162544 74248
rect 177856 74196 177908 74248
rect 208952 74196 209004 74248
rect 108764 74128 108816 74180
rect 142252 74128 142304 74180
rect 169024 74128 169076 74180
rect 195060 74128 195112 74180
rect 112536 74060 112588 74112
rect 146116 74060 146168 74112
rect 163780 74060 163832 74112
rect 198004 74060 198056 74112
rect 102692 73992 102744 74044
rect 135812 73992 135864 74044
rect 145104 73992 145156 74044
rect 145564 73992 145616 74044
rect 145656 73992 145708 74044
rect 145932 73992 145984 74044
rect 149336 73992 149388 74044
rect 149888 73992 149940 74044
rect 173440 73992 173492 74044
rect 206192 73992 206244 74044
rect 111340 73924 111392 73976
rect 142620 73924 142672 73976
rect 174728 73924 174780 73976
rect 207020 73924 207072 73976
rect 74540 73856 74592 73908
rect 117228 73856 117280 73908
rect 152464 73856 152516 73908
rect 162676 73856 162728 73908
rect 189172 73856 189224 73908
rect 189816 73856 189868 73908
rect 321560 73856 321612 73908
rect 35164 73788 35216 73840
rect 100300 73788 100352 73840
rect 115296 73788 115348 73840
rect 145104 73788 145156 73840
rect 161296 73788 161348 73840
rect 184940 73788 184992 73840
rect 215392 73788 215444 73840
rect 560944 73788 560996 73840
rect 112628 73720 112680 73772
rect 138204 73720 138256 73772
rect 138848 73720 138900 73772
rect 149704 73720 149756 73772
rect 221280 73720 221332 73772
rect 115204 73652 115256 73704
rect 151268 73652 151320 73704
rect 154580 73652 154632 73704
rect 189172 73652 189224 73704
rect 100300 73584 100352 73636
rect 135168 73584 135220 73636
rect 106280 73516 106332 73568
rect 107476 73516 107528 73568
rect 131764 73448 131816 73500
rect 137744 73448 137796 73500
rect 153384 73312 153436 73364
rect 154028 73312 154080 73364
rect 149336 73176 149388 73228
rect 182824 73176 182876 73228
rect 3148 73108 3200 73160
rect 152464 73108 152516 73160
rect 171876 73108 171928 73160
rect 197360 73108 197412 73160
rect 218060 73108 218112 73160
rect 218612 73108 218664 73160
rect 580172 73108 580224 73160
rect 121092 73040 121144 73092
rect 114836 72972 114888 73024
rect 149244 72972 149296 73024
rect 149796 73040 149848 73092
rect 150348 73040 150400 73092
rect 171048 73040 171100 73092
rect 195980 73040 196032 73092
rect 157156 72972 157208 73024
rect 173900 72972 173952 73024
rect 200488 72972 200540 73024
rect 119896 72904 119948 72956
rect 152280 72904 152332 72956
rect 156512 72904 156564 72956
rect 190920 72904 190972 72956
rect 126244 72836 126296 72888
rect 153016 72836 153068 72888
rect 161388 72836 161440 72888
rect 194968 72836 195020 72888
rect 114100 72768 114152 72820
rect 148784 72768 148836 72820
rect 162768 72768 162820 72820
rect 163964 72768 164016 72820
rect 167920 72768 167972 72820
rect 201960 72768 202012 72820
rect 114928 72700 114980 72752
rect 149060 72700 149112 72752
rect 163412 72700 163464 72752
rect 197728 72700 197780 72752
rect 111708 72632 111760 72684
rect 143540 72632 143592 72684
rect 153568 72632 153620 72684
rect 158352 72632 158404 72684
rect 177948 72632 178000 72684
rect 208400 72632 208452 72684
rect 120908 72564 120960 72616
rect 151820 72564 151872 72616
rect 173716 72564 173768 72616
rect 204904 72564 204956 72616
rect 115388 72496 115440 72548
rect 146944 72496 146996 72548
rect 159916 72496 159968 72548
rect 193496 72496 193548 72548
rect 52460 72428 52512 72480
rect 98828 72428 98880 72480
rect 124220 72428 124272 72480
rect 175464 72428 175516 72480
rect 184940 72428 184992 72480
rect 186228 72428 186280 72480
rect 194600 72428 194652 72480
rect 253940 72428 253992 72480
rect 119988 72360 120040 72412
rect 149796 72360 149848 72412
rect 155592 72360 155644 72412
rect 218060 72360 218112 72412
rect 98828 72292 98880 72344
rect 133144 72292 133196 72344
rect 161112 72292 161164 72344
rect 195152 72292 195204 72344
rect 98736 72224 98788 72276
rect 133880 72224 133932 72276
rect 157432 72224 157484 72276
rect 192392 72224 192444 72276
rect 133144 72156 133196 72208
rect 133604 72156 133656 72208
rect 165528 72156 165580 72208
rect 184204 72156 184256 72208
rect 121736 71680 121788 71732
rect 142988 71680 143040 71732
rect 148416 71680 148468 71732
rect 148692 71680 148744 71732
rect 158628 71680 158680 71732
rect 219716 71680 219768 71732
rect 116860 71612 116912 71664
rect 151360 71612 151412 71664
rect 151728 71612 151780 71664
rect 172244 71612 172296 71664
rect 215852 71612 215904 71664
rect 123484 71544 123536 71596
rect 142896 71544 142948 71596
rect 111064 71476 111116 71528
rect 141700 71476 141752 71528
rect 115664 71408 115716 71460
rect 147680 71408 147732 71460
rect 148324 71408 148376 71460
rect 117044 71340 117096 71392
rect 148416 71340 148468 71392
rect 108856 71272 108908 71324
rect 139124 71272 139176 71324
rect 106740 71204 106792 71256
rect 130844 71204 130896 71256
rect 153108 71204 153160 71256
rect 175188 71544 175240 71596
rect 197636 71544 197688 71596
rect 172704 71476 172756 71528
rect 207388 71476 207440 71528
rect 176936 71408 176988 71460
rect 210148 71408 210200 71460
rect 176752 71340 176804 71392
rect 209872 71340 209924 71392
rect 172152 71272 172204 71324
rect 204444 71272 204496 71324
rect 176108 71204 176160 71256
rect 207296 71204 207348 71256
rect 110972 71136 111024 71188
rect 137192 71136 137244 71188
rect 171508 71136 171560 71188
rect 202880 71136 202932 71188
rect 151728 71068 151780 71120
rect 306380 71068 306432 71120
rect 2780 71000 2832 71052
rect 157432 71000 157484 71052
rect 176016 71000 176068 71052
rect 176292 71000 176344 71052
rect 206468 71000 206520 71052
rect 215852 71000 215904 71052
rect 484400 71000 484452 71052
rect 93768 70932 93820 70984
rect 156972 70932 157024 70984
rect 180248 70932 180300 70984
rect 188988 70932 189040 70984
rect 207756 70932 207808 70984
rect 114192 70864 114244 70916
rect 147128 70864 147180 70916
rect 156328 70864 156380 70916
rect 192024 70864 192076 70916
rect 106832 70796 106884 70848
rect 132408 70796 132460 70848
rect 127624 70728 127676 70780
rect 150532 70728 150584 70780
rect 160468 70728 160520 70780
rect 161388 70728 161440 70780
rect 108948 70320 109000 70372
rect 135904 70320 135956 70372
rect 166172 70320 166224 70372
rect 207848 70320 207900 70372
rect 118608 70252 118660 70304
rect 150992 70252 151044 70304
rect 164700 70252 164752 70304
rect 199476 70252 199528 70304
rect 109776 70184 109828 70236
rect 151176 70184 151228 70236
rect 175556 70184 175608 70236
rect 210240 70184 210292 70236
rect 115572 70116 115624 70168
rect 149336 70116 149388 70168
rect 167092 70116 167144 70168
rect 167460 70116 167512 70168
rect 202144 70116 202196 70168
rect 117964 70048 118016 70100
rect 152924 70048 152976 70100
rect 157616 70048 157668 70100
rect 158536 70048 158588 70100
rect 192208 70048 192260 70100
rect 122012 69980 122064 70032
rect 156696 69980 156748 70032
rect 160284 69980 160336 70032
rect 161204 69980 161256 70032
rect 194784 69980 194836 70032
rect 99012 69912 99064 69964
rect 133788 69912 133840 69964
rect 172520 69912 172572 69964
rect 206100 69912 206152 69964
rect 108672 69844 108724 69896
rect 141516 69844 141568 69896
rect 172612 69844 172664 69896
rect 173164 69844 173216 69896
rect 205824 69844 205876 69896
rect 113824 69776 113876 69828
rect 147404 69776 147456 69828
rect 157708 69776 157760 69828
rect 158628 69776 158680 69828
rect 190736 69776 190788 69828
rect 13084 69708 13136 69760
rect 94964 69708 95016 69760
rect 95148 69708 95200 69760
rect 126244 69708 126296 69760
rect 167092 69708 167144 69760
rect 172704 69708 172756 69760
rect 198740 69708 198792 69760
rect 78680 69640 78732 69692
rect 160468 69640 160520 69692
rect 166172 69640 166224 69692
rect 197820 69640 197872 69692
rect 314660 69640 314712 69692
rect 108028 69572 108080 69624
rect 152188 69572 152240 69624
rect 160376 69572 160428 69624
rect 161388 69572 161440 69624
rect 192668 69572 192720 69624
rect 95148 69504 95200 69556
rect 139216 69504 139268 69556
rect 162124 69504 162176 69556
rect 162584 69504 162636 69556
rect 165160 69504 165212 69556
rect 174544 69504 174596 69556
rect 164148 69436 164200 69488
rect 181628 69436 181680 69488
rect 162584 69368 162636 69420
rect 181536 69368 181588 69420
rect 107200 68960 107252 69012
rect 136456 68960 136508 69012
rect 162032 68960 162084 69012
rect 162676 68960 162728 69012
rect 163136 68960 163188 69012
rect 164056 68960 164108 69012
rect 166632 68960 166684 69012
rect 191104 68960 191156 69012
rect 111248 68892 111300 68944
rect 138664 68892 138716 68944
rect 160192 68892 160244 68944
rect 194876 68892 194928 68944
rect 110328 68824 110380 68876
rect 156236 68824 156288 68876
rect 167368 68824 167420 68876
rect 201868 68824 201920 68876
rect 104164 68756 104216 68808
rect 138572 68756 138624 68808
rect 155868 68756 155920 68808
rect 189448 68756 189500 68808
rect 112168 68688 112220 68740
rect 146484 68688 146536 68740
rect 164056 68688 164108 68740
rect 197544 68688 197596 68740
rect 99196 68620 99248 68672
rect 133144 68620 133196 68672
rect 161848 68620 161900 68672
rect 196256 68620 196308 68672
rect 114284 68552 114336 68604
rect 146852 68552 146904 68604
rect 159180 68552 159232 68604
rect 193312 68552 193364 68604
rect 116216 68484 116268 68536
rect 148600 68484 148652 68536
rect 159272 68484 159324 68536
rect 194232 68484 194284 68536
rect 111524 68416 111576 68468
rect 141424 68416 141476 68468
rect 174636 68416 174688 68468
rect 207480 68416 207532 68468
rect 120724 68348 120776 68400
rect 150072 68348 150124 68400
rect 150440 68348 150492 68400
rect 310520 68348 310572 68400
rect 95884 68280 95936 68332
rect 132500 68280 132552 68332
rect 139860 68280 139912 68332
rect 149244 68280 149296 68332
rect 462320 68280 462372 68332
rect 107016 68212 107068 68264
rect 135536 68212 135588 68264
rect 162676 68212 162728 68264
rect 181444 68212 181496 68264
rect 182180 68212 182232 68264
rect 211160 68212 211212 68264
rect 3516 68144 3568 68196
rect 153108 68144 153160 68196
rect 163320 68144 163372 68196
rect 208768 68144 208820 68196
rect 105360 68076 105412 68128
rect 155040 68076 155092 68128
rect 155868 68076 155920 68128
rect 156236 68008 156288 68060
rect 156696 68008 156748 68060
rect 109684 67532 109736 67584
rect 144368 67532 144420 67584
rect 145472 67532 145524 67584
rect 145656 67532 145708 67584
rect 164516 67532 164568 67584
rect 165436 67532 165488 67584
rect 165988 67532 166040 67584
rect 166816 67532 166868 67584
rect 167736 67532 167788 67584
rect 192852 67532 192904 67584
rect 104440 67464 104492 67516
rect 136640 67464 136692 67516
rect 136824 67464 136876 67516
rect 137284 67464 137336 67516
rect 138756 67464 138808 67516
rect 138940 67464 138992 67516
rect 157524 67464 157576 67516
rect 207204 67464 207256 67516
rect 109960 67396 110012 67448
rect 143632 67396 143684 67448
rect 144276 67396 144328 67448
rect 165896 67396 165948 67448
rect 166908 67396 166960 67448
rect 169944 67396 169996 67448
rect 211988 67396 212040 67448
rect 110880 67328 110932 67380
rect 145656 67328 145708 67380
rect 153476 67328 153528 67380
rect 188804 67328 188856 67380
rect 104348 67260 104400 67312
rect 136824 67260 136876 67312
rect 161848 67260 161900 67312
rect 165620 67260 165672 67312
rect 200764 67260 200816 67312
rect 104716 67192 104768 67244
rect 136916 67192 136968 67244
rect 168840 67192 168892 67244
rect 169208 67192 169260 67244
rect 203708 67192 203760 67244
rect 104624 67124 104676 67176
rect 136732 67124 136784 67176
rect 166908 67124 166960 67176
rect 200672 67124 200724 67176
rect 103244 67056 103296 67108
rect 134892 67056 134944 67108
rect 136640 67056 136692 67108
rect 138756 67056 138808 67108
rect 165436 67056 165488 67108
rect 199660 67056 199712 67108
rect 93860 66988 93912 67040
rect 166172 66988 166224 67040
rect 175372 66988 175424 67040
rect 210056 66988 210108 67040
rect 121552 66920 121604 66972
rect 148140 66920 148192 66972
rect 161756 66920 161808 66972
rect 196348 66920 196400 66972
rect 386420 66920 386472 66972
rect 26240 66852 26292 66904
rect 104256 66852 104308 66904
rect 104716 66852 104768 66904
rect 129740 66852 129792 66904
rect 130384 66852 130436 66904
rect 145932 66852 145984 66904
rect 488540 66852 488592 66904
rect 120632 66784 120684 66836
rect 148232 66784 148284 66836
rect 166816 66784 166868 66836
rect 200580 66784 200632 66836
rect 121644 66716 121696 66768
rect 149612 66716 149664 66768
rect 156144 66716 156196 66768
rect 216036 66716 216088 66768
rect 110052 66648 110104 66700
rect 129740 66648 129792 66700
rect 89720 66580 89772 66632
rect 168840 66580 168892 66632
rect 121184 66172 121236 66224
rect 135996 66172 136048 66224
rect 158996 66172 159048 66224
rect 221004 66172 221056 66224
rect 120540 66104 120592 66156
rect 141056 66104 141108 66156
rect 157340 66104 157392 66156
rect 211344 66104 211396 66156
rect 100392 66036 100444 66088
rect 134340 66036 134392 66088
rect 154856 66036 154908 66088
rect 189264 66036 189316 66088
rect 98920 65968 98972 66020
rect 133144 65968 133196 66020
rect 133420 65968 133472 66020
rect 156880 65968 156932 66020
rect 191012 65968 191064 66020
rect 104072 65900 104124 65952
rect 138480 65900 138532 65952
rect 169760 65900 169812 65952
rect 171048 65900 171100 65952
rect 204720 65900 204772 65952
rect 105452 65832 105504 65884
rect 140320 65832 140372 65884
rect 171324 65832 171376 65884
rect 172336 65832 172388 65884
rect 174084 65832 174136 65884
rect 175096 65832 175148 65884
rect 175280 65832 175332 65884
rect 176568 65832 176620 65884
rect 176660 65832 176712 65884
rect 205916 65832 205968 65884
rect 100576 65764 100628 65816
rect 134156 65764 134208 65816
rect 135904 65764 135956 65816
rect 206008 65764 206060 65816
rect 107568 65696 107620 65748
rect 141148 65696 141200 65748
rect 160100 65696 160152 65748
rect 195520 65696 195572 65748
rect 167276 65628 167328 65680
rect 201776 65628 201828 65680
rect 102600 65560 102652 65612
rect 135444 65560 135496 65612
rect 147220 65560 147272 65612
rect 260840 65560 260892 65612
rect 67640 65492 67692 65544
rect 110144 65492 110196 65544
rect 142712 65492 142764 65544
rect 146024 65492 146076 65544
rect 408500 65492 408552 65544
rect 111432 65424 111484 65476
rect 140872 65424 140924 65476
rect 141516 65424 141568 65476
rect 171232 65424 171284 65476
rect 172428 65424 172480 65476
rect 175096 65424 175148 65476
rect 208584 65424 208636 65476
rect 101404 65356 101456 65408
rect 140596 65356 140648 65408
rect 158352 65356 158404 65408
rect 188620 65356 188672 65408
rect 100024 65288 100076 65340
rect 134708 65288 134760 65340
rect 176568 65288 176620 65340
rect 210332 65288 210384 65340
rect 100484 65220 100536 65272
rect 134984 65220 135036 65272
rect 172428 65220 172480 65272
rect 176660 65220 176712 65272
rect 106096 64812 106148 64864
rect 135628 64812 135680 64864
rect 138296 64812 138348 64864
rect 580724 64812 580776 64864
rect 112904 64744 112956 64796
rect 141332 64744 141384 64796
rect 154764 64744 154816 64796
rect 215944 64744 215996 64796
rect 96344 64676 96396 64728
rect 136088 64676 136140 64728
rect 168748 64676 168800 64728
rect 212540 64676 212592 64728
rect 99104 64608 99156 64660
rect 133236 64608 133288 64660
rect 175188 64608 175240 64660
rect 213920 64608 213972 64660
rect 100668 64540 100720 64592
rect 134616 64540 134668 64592
rect 158904 64540 158956 64592
rect 188344 64540 188396 64592
rect 99932 64472 99984 64524
rect 134432 64472 134484 64524
rect 165068 64472 165120 64524
rect 191380 64472 191432 64524
rect 108396 64404 108448 64456
rect 141424 64404 141476 64456
rect 142068 64404 142120 64456
rect 163044 64404 163096 64456
rect 188896 64404 188948 64456
rect 107292 64336 107344 64388
rect 139768 64336 139820 64388
rect 107384 64268 107436 64320
rect 139676 64268 139728 64320
rect 148232 64268 148284 64320
rect 184940 64268 184992 64320
rect 102784 64200 102836 64252
rect 132960 64200 133012 64252
rect 133328 64200 133380 64252
rect 264980 64200 265032 64252
rect 63500 64132 63552 64184
rect 106096 64132 106148 64184
rect 108580 64132 108632 64184
rect 139584 64132 139636 64184
rect 142896 64132 142948 64184
rect 477500 64132 477552 64184
rect 97264 64064 97316 64116
rect 138664 64064 138716 64116
rect 97356 63996 97408 64048
rect 137100 63996 137152 64048
rect 133880 63860 133932 63912
rect 134432 63860 134484 63912
rect 139676 63588 139728 63640
rect 140136 63588 140188 63640
rect 173992 63588 174044 63640
rect 175188 63588 175240 63640
rect 102140 63520 102192 63572
rect 102784 63520 102836 63572
rect 137100 63520 137152 63572
rect 137376 63520 137428 63572
rect 139768 63520 139820 63572
rect 140044 63520 140096 63572
rect 97816 63452 97868 63504
rect 158812 63452 158864 63504
rect 162768 63452 162820 63504
rect 211528 63452 211580 63504
rect 96436 63384 96488 63436
rect 150808 63384 150860 63436
rect 168656 63384 168708 63436
rect 212632 63384 212684 63436
rect 101956 63316 102008 63368
rect 142528 63316 142580 63368
rect 143448 63316 143500 63368
rect 162860 63316 162912 63368
rect 204260 63316 204312 63368
rect 115020 63248 115072 63300
rect 153384 63248 153436 63300
rect 165528 63248 165580 63300
rect 206560 63248 206612 63300
rect 119620 63180 119672 63232
rect 151912 63180 151964 63232
rect 152556 63180 152608 63232
rect 169576 63180 169628 63232
rect 209780 63180 209832 63232
rect 109592 63112 109644 63164
rect 131120 63112 131172 63164
rect 164332 63112 164384 63164
rect 199568 63112 199620 63164
rect 168288 63044 168340 63096
rect 202052 63044 202104 63096
rect 165620 62976 165672 63028
rect 213184 62976 213236 63028
rect 146300 62908 146352 62960
rect 213092 62908 213144 62960
rect 148508 62840 148560 62892
rect 302240 62840 302292 62892
rect 8944 62772 8996 62824
rect 97816 62772 97868 62824
rect 168564 62772 168616 62824
rect 203432 62772 203484 62824
rect 425060 62772 425112 62824
rect 162952 62704 163004 62756
rect 197452 62704 197504 62756
rect 170680 62636 170732 62688
rect 203524 62636 203576 62688
rect 166724 62568 166776 62620
rect 194048 62568 194100 62620
rect 164424 62500 164476 62552
rect 165528 62500 165580 62552
rect 131120 62432 131172 62484
rect 131856 62432 131908 62484
rect 165804 62364 165856 62416
rect 166724 62364 166776 62416
rect 153384 62092 153436 62144
rect 153844 62092 153896 62144
rect 96068 62024 96120 62076
rect 96252 62024 96304 62076
rect 161572 62024 161624 62076
rect 168472 62024 168524 62076
rect 203340 62024 203392 62076
rect 149796 61412 149848 61464
rect 295340 61412 295392 61464
rect 6920 61344 6972 61396
rect 96068 61344 96120 61396
rect 203340 61344 203392 61396
rect 496084 61344 496136 61396
rect 3516 60664 3568 60716
rect 161848 60664 161900 60716
rect 174452 60664 174504 60716
rect 198740 60664 198792 60716
rect 199016 60664 199068 60716
rect 156788 60596 156840 60648
rect 190644 60596 190696 60648
rect 192484 60596 192536 60648
rect 134248 59984 134300 60036
rect 454040 59984 454092 60036
rect 198740 59848 198792 59900
rect 200120 59848 200172 59900
rect 134892 58760 134944 58812
rect 215300 58760 215352 58812
rect 31024 58692 31076 58744
rect 162860 58692 162912 58744
rect 143448 58624 143500 58676
rect 545764 58624 545816 58676
rect 105636 57876 105688 57928
rect 106188 57876 106240 57928
rect 140228 57876 140280 57928
rect 154672 57876 154724 57928
rect 218060 57876 218112 57928
rect 218520 57876 218572 57928
rect 158444 57808 158496 57860
rect 191932 57808 191984 57860
rect 193128 57808 193180 57860
rect 193128 57264 193180 57316
rect 256700 57264 256752 57316
rect 71780 57196 71832 57248
rect 105636 57196 105688 57248
rect 218060 57196 218112 57248
rect 470600 57196 470652 57248
rect 150440 56584 150492 56636
rect 151912 56584 151964 56636
rect 186228 56516 186280 56568
rect 579896 56516 579948 56568
rect 164240 55972 164292 56024
rect 184848 55972 184900 56024
rect 17960 55904 18012 55956
rect 176016 55904 176068 55956
rect 141516 55836 141568 55888
rect 345020 55836 345072 55888
rect 95056 55156 95108 55208
rect 139952 55156 140004 55208
rect 165712 55156 165764 55208
rect 200212 55156 200264 55208
rect 201408 55156 201460 55208
rect 184848 55088 184900 55140
rect 199108 55088 199160 55140
rect 145656 54544 145708 54596
rect 234620 54544 234672 54596
rect 48320 54476 48372 54528
rect 95056 54476 95108 54528
rect 201408 54476 201460 54528
rect 578884 54476 578936 54528
rect 167092 53728 167144 53780
rect 201500 53728 201552 53780
rect 202788 53728 202840 53780
rect 202788 53116 202840 53168
rect 276020 53116 276072 53168
rect 147128 53048 147180 53100
rect 542360 53048 542412 53100
rect 3516 52368 3568 52420
rect 8944 52368 8996 52420
rect 182916 52368 182968 52420
rect 579896 52368 579948 52420
rect 154396 51756 154448 51808
rect 186228 51756 186280 51808
rect 188712 51756 188764 51808
rect 133236 51688 133288 51740
rect 502984 51688 503036 51740
rect 135996 51008 136048 51060
rect 144184 51008 144236 51060
rect 167000 51008 167052 51060
rect 196164 51008 196216 51060
rect 144368 50396 144420 50448
rect 400864 50396 400916 50448
rect 196164 50328 196216 50380
rect 553400 50328 553452 50380
rect 169760 49648 169812 49700
rect 173164 49648 173216 49700
rect 174544 49648 174596 49700
rect 199200 49648 199252 49700
rect 580172 49648 580224 49700
rect 140136 48968 140188 49020
rect 374644 48968 374696 49020
rect 3516 48220 3568 48272
rect 122104 48220 122156 48272
rect 144460 48220 144512 48272
rect 150900 48220 150952 48272
rect 220820 48220 220872 48272
rect 222108 48220 222160 48272
rect 169852 48152 169904 48204
rect 203248 48152 203300 48204
rect 204168 48152 204220 48204
rect 204168 47608 204220 47660
rect 284300 47608 284352 47660
rect 222108 47540 222160 47592
rect 420920 47540 420972 47592
rect 168380 46860 168432 46912
rect 203156 46860 203208 46912
rect 204168 46860 204220 46912
rect 171140 46792 171192 46844
rect 205640 46792 205692 46844
rect 205640 46248 205692 46300
rect 230480 46248 230532 46300
rect 204168 46180 204220 46232
rect 556804 46180 556856 46232
rect 153936 45500 153988 45552
rect 579988 45500 580040 45552
rect 137376 44820 137428 44872
rect 436100 44820 436152 44872
rect 3516 44072 3568 44124
rect 103428 44072 103480 44124
rect 131764 44072 131816 44124
rect 147036 43460 147088 43512
rect 394700 43460 394752 43512
rect 138848 43392 138900 43444
rect 557540 43392 557592 43444
rect 133144 42100 133196 42152
rect 377404 42100 377456 42152
rect 148416 42032 148468 42084
rect 503720 42032 503772 42084
rect 158260 41352 158312 41404
rect 190460 41352 190512 41404
rect 580172 41352 580224 41404
rect 138756 40672 138808 40724
rect 390560 40672 390612 40724
rect 3516 39992 3568 40044
rect 126244 39992 126296 40044
rect 164056 39380 164108 39432
rect 245660 39380 245712 39432
rect 176568 39312 176620 39364
rect 340880 39312 340932 39364
rect 155592 38564 155644 38616
rect 189172 38564 189224 38616
rect 189632 38564 189684 38616
rect 189172 37952 189224 38004
rect 378140 37952 378192 38004
rect 137284 37884 137336 37936
rect 442264 37884 442316 37936
rect 3148 37204 3200 37256
rect 133880 37204 133932 37256
rect 192484 37204 192536 37256
rect 580172 37204 580224 37256
rect 144276 36524 144328 36576
rect 219440 36524 219492 36576
rect 158536 35232 158588 35284
rect 371240 35232 371292 35284
rect 168288 35164 168340 35216
rect 548524 35164 548576 35216
rect 158720 34416 158772 34468
rect 190552 34416 190604 34468
rect 191748 34416 191800 34468
rect 161480 34348 161532 34400
rect 191932 34348 191984 34400
rect 193128 34348 193180 34400
rect 191748 33736 191800 33788
rect 356060 33736 356112 33788
rect 193128 33124 193180 33176
rect 571984 33124 572036 33176
rect 152464 33056 152516 33108
rect 580172 33056 580224 33108
rect 161204 31084 161256 31136
rect 364340 31084 364392 31136
rect 166724 31016 166776 31068
rect 563704 31016 563756 31068
rect 154028 30268 154080 30320
rect 189172 30268 189224 30320
rect 165436 29656 165488 29708
rect 332600 29656 332652 29708
rect 189172 29588 189224 29640
rect 189908 29588 189960 29640
rect 500224 29588 500276 29640
rect 3148 28908 3200 28960
rect 138204 28908 138256 28960
rect 188988 28908 189040 28960
rect 580172 28908 580224 28960
rect 141424 28228 141476 28280
rect 207664 28228 207716 28280
rect 166816 26936 166868 26988
rect 249800 26936 249852 26988
rect 148324 26868 148376 26920
rect 347780 26868 347832 26920
rect 162676 25508 162728 25560
rect 473360 25508 473412 25560
rect 182088 24760 182140 24812
rect 580172 24760 580224 24812
rect 134708 24080 134760 24132
rect 210424 24080 210476 24132
rect 171048 22720 171100 22772
rect 514024 22720 514076 22772
rect 166908 21360 166960 21412
rect 466460 21360 466512 21412
rect 3148 20612 3200 20664
rect 139584 20612 139636 20664
rect 161296 20612 161348 20664
rect 580172 20612 580224 20664
rect 146944 18640 146996 18692
rect 226340 18640 226392 18692
rect 175096 18572 175148 18624
rect 481640 18572 481692 18624
rect 161388 17212 161440 17264
rect 527180 17212 527232 17264
rect 3332 16532 3384 16584
rect 131120 16532 131172 16584
rect 182824 16532 182876 16584
rect 580172 16532 580224 16584
rect 156696 15852 156748 15904
rect 178408 15852 178460 15904
rect 153844 14560 153896 14612
rect 204352 14560 204404 14612
rect 172336 14492 172388 14544
rect 352472 14492 352524 14544
rect 140044 14424 140096 14476
rect 459192 14424 459244 14476
rect 162952 13200 163004 13252
rect 175924 13200 175976 13252
rect 175188 13132 175240 13184
rect 447600 13132 447652 13184
rect 134524 13064 134576 13116
rect 531320 13064 531372 13116
rect 3056 12384 3108 12436
rect 129740 12384 129792 12436
rect 186228 12384 186280 12436
rect 580172 12384 580224 12436
rect 149704 11704 149756 11756
rect 193220 11704 193272 11756
rect 172428 10344 172480 10396
rect 299480 10344 299532 10396
rect 157248 10276 157300 10328
rect 562324 10276 562376 10328
rect 134616 8916 134668 8968
rect 241704 8916 241756 8968
rect 2964 8236 3016 8288
rect 151820 8236 151872 8288
rect 560944 8236 560996 8288
rect 580172 8236 580224 8288
rect 162584 7624 162636 7676
rect 318800 7624 318852 7676
rect 164148 7556 164200 7608
rect 360660 7556 360712 7608
rect 110144 6196 110196 6248
rect 147680 6196 147732 6248
rect 158628 6196 158680 6248
rect 398656 6196 398708 6248
rect 138664 6128 138716 6180
rect 432788 6128 432840 6180
rect 184848 5448 184900 5500
rect 580172 5448 580224 5500
rect 145564 4768 145616 4820
rect 155224 4768 155276 4820
rect 165528 4768 165580 4820
rect 280804 4768 280856 4820
rect 2780 4020 2832 4072
rect 4804 4020 4856 4072
rect 117228 3544 117280 3596
rect 156604 3544 156656 3596
rect 165620 3544 165672 3596
rect 166816 3544 166868 3596
rect 174544 3544 174596 3596
rect 191840 3544 191892 3596
rect 207664 3544 207716 3596
rect 208676 3544 208728 3596
rect 210424 3544 210476 3596
rect 242808 3544 242860 3596
rect 377404 3544 377456 3596
rect 30288 3476 30340 3528
rect 31024 3476 31076 3528
rect 34152 3476 34204 3528
rect 35164 3476 35216 3528
rect 97908 3476 97960 3528
rect 128820 3476 128872 3528
rect 136548 3476 136600 3528
rect 211252 3476 211304 3528
rect 211804 3476 211856 3528
rect 212540 3476 212592 3528
rect 241704 3476 241756 3528
rect 326528 3476 326580 3528
rect 374644 3476 374696 3528
rect 375472 3476 375524 3528
rect 378140 3476 378192 3528
rect 379336 3476 379388 3528
rect 508780 3476 508832 3528
rect 545764 3476 545816 3528
rect 546776 3476 546828 3528
rect 571984 3476 572036 3528
rect 573180 3476 573232 3528
rect 20 3408 72 3460
rect 13084 3408 13136 3460
rect 14832 3408 14884 3460
rect 135444 3408 135496 3460
rect 142804 3408 142856 3460
rect 144276 3408 144328 3460
rect 146300 3408 146352 3460
rect 147496 3408 147548 3460
rect 144184 3340 144236 3392
rect 383200 3408 383252 3460
rect 400864 3408 400916 3460
rect 402520 3408 402572 3460
rect 442264 3408 442316 3460
rect 443736 3408 443788 3460
rect 454040 3408 454092 3460
rect 455328 3408 455380 3460
rect 473360 3408 473412 3460
rect 474648 3408 474700 3460
rect 496084 3408 496136 3460
rect 497188 3408 497240 3460
rect 502984 3408 503036 3460
rect 539048 3408 539100 3460
rect 556804 3408 556856 3460
rect 561588 3408 561640 3460
rect 562324 3408 562376 3460
rect 577044 3340 577096 3392
rect 135904 3272 135956 3324
rect 140412 3272 140464 3324
rect 548524 3068 548576 3120
rect 550640 3068 550692 3120
rect 514024 3000 514076 3052
rect 515864 3000 515916 3052
rect 563704 3000 563756 3052
rect 565452 3000 565504 3052
rect 500224 2864 500276 2916
rect 501052 2864 501104 2916
<< metal2 >>
rect 634 703520 746 704960
rect 4498 703520 4610 704960
rect 8362 703520 8474 704960
rect 12226 703520 12338 704960
rect 16090 703520 16202 704960
rect 19954 703520 20066 704960
rect 23818 703520 23930 704960
rect 27682 703520 27794 704960
rect 31546 703520 31658 704960
rect 34766 703520 34878 704960
rect 38630 703520 38742 704960
rect 42494 703520 42606 704960
rect 46358 703520 46470 704960
rect 49712 703582 50108 703610
rect 676 700330 704 703520
rect 3422 701176 3478 701185
rect 3422 701111 3478 701120
rect 3436 701078 3464 701111
rect 3424 701072 3476 701078
rect 3424 701014 3476 701020
rect 4540 700602 4568 703520
rect 4528 700596 4580 700602
rect 4528 700538 4580 700544
rect 664 700324 716 700330
rect 664 700266 716 700272
rect 3054 697776 3110 697785
rect 3054 697711 3110 697720
rect 3068 696998 3096 697711
rect 3056 696992 3108 696998
rect 3056 696934 3108 696940
rect 3422 689616 3478 689625
rect 3422 689551 3478 689560
rect 3436 688702 3464 689551
rect 3424 688696 3476 688702
rect 3424 688638 3476 688644
rect 3146 685536 3202 685545
rect 3146 685471 3202 685480
rect 3160 684554 3188 685471
rect 3148 684548 3200 684554
rect 3148 684490 3200 684496
rect 8404 683114 8432 703520
rect 12268 700398 12296 703520
rect 12256 700392 12308 700398
rect 12256 700334 12308 700340
rect 16132 698970 16160 703520
rect 19996 700534 20024 703520
rect 19984 700528 20036 700534
rect 19984 700470 20036 700476
rect 23860 700466 23888 703520
rect 26884 700596 26936 700602
rect 26884 700538 26936 700544
rect 23848 700460 23900 700466
rect 23848 700402 23900 700408
rect 16120 698964 16172 698970
rect 16120 698906 16172 698912
rect 14464 688696 14516 688702
rect 14464 688638 14516 688644
rect 8312 683086 8432 683114
rect 3422 681456 3478 681465
rect 3422 681391 3478 681400
rect 3436 680406 3464 681391
rect 3424 680400 3476 680406
rect 3424 680342 3476 680348
rect 3422 677376 3478 677385
rect 3422 677311 3478 677320
rect 3436 676258 3464 677311
rect 3424 676252 3476 676258
rect 3424 676194 3476 676200
rect 3238 665136 3294 665145
rect 3238 665071 3294 665080
rect 3252 663814 3280 665071
rect 3240 663808 3292 663814
rect 3240 663750 3292 663756
rect 3424 661088 3476 661094
rect 3422 661056 3424 661065
rect 3476 661056 3478 661065
rect 3422 660991 3478 661000
rect 3054 653576 3110 653585
rect 3054 653511 3110 653520
rect 3068 652798 3096 653511
rect 3056 652792 3108 652798
rect 3056 652734 3108 652740
rect 3422 645416 3478 645425
rect 3422 645351 3478 645360
rect 3436 644502 3464 645351
rect 3424 644496 3476 644502
rect 3424 644438 3476 644444
rect 3146 641336 3202 641345
rect 3146 641271 3202 641280
rect 3160 640354 3188 641271
rect 3148 640348 3200 640354
rect 3148 640290 3200 640296
rect 3146 637256 3202 637265
rect 3146 637191 3202 637200
rect 3160 636274 3188 637191
rect 3148 636268 3200 636274
rect 3148 636210 3200 636216
rect 3422 633176 3478 633185
rect 3422 633111 3478 633120
rect 3436 632126 3464 633111
rect 3424 632120 3476 632126
rect 3424 632062 3476 632068
rect 3238 625016 3294 625025
rect 3238 624951 3294 624960
rect 3252 623830 3280 624951
rect 3240 623824 3292 623830
rect 3240 623766 3292 623772
rect 3422 621616 3478 621625
rect 3422 621551 3478 621560
rect 3436 621042 3464 621551
rect 3424 621036 3476 621042
rect 3424 620978 3476 620984
rect 3146 617536 3202 617545
rect 3146 617471 3202 617480
rect 3160 616894 3188 617471
rect 3148 616888 3200 616894
rect 3148 616830 3200 616836
rect 3146 613456 3202 613465
rect 3146 613391 3202 613400
rect 3160 612814 3188 613391
rect 3148 612808 3200 612814
rect 3148 612750 3200 612756
rect 3422 609376 3478 609385
rect 3422 609311 3478 609320
rect 3054 605296 3110 605305
rect 3054 605231 3110 605240
rect 3068 604518 3096 605231
rect 3056 604512 3108 604518
rect 3056 604454 3108 604460
rect 3054 597136 3110 597145
rect 3054 597071 3110 597080
rect 3068 596222 3096 597071
rect 3056 596216 3108 596222
rect 3056 596158 3108 596164
rect 3146 593056 3202 593065
rect 3146 592991 3202 593000
rect 3160 592074 3188 592991
rect 3148 592068 3200 592074
rect 3148 592010 3200 592016
rect 3238 588976 3294 588985
rect 3238 588911 3294 588920
rect 3252 587926 3280 588911
rect 3240 587920 3292 587926
rect 3240 587862 3292 587868
rect 3146 584896 3202 584905
rect 3146 584831 3202 584840
rect 3160 583778 3188 584831
rect 3148 583772 3200 583778
rect 3148 583714 3200 583720
rect 3330 581496 3386 581505
rect 3330 581431 3386 581440
rect 3344 581058 3372 581431
rect 3332 581052 3384 581058
rect 3332 580994 3384 581000
rect 2870 569256 2926 569265
rect 2870 569191 2926 569200
rect 2884 568614 2912 569191
rect 2872 568608 2924 568614
rect 2872 568550 2924 568556
rect 3054 561096 3110 561105
rect 3054 561031 3110 561040
rect 3068 560318 3096 561031
rect 3056 560312 3108 560318
rect 3056 560254 3108 560260
rect 3054 557016 3110 557025
rect 3054 556951 3110 556960
rect 3068 556238 3096 556951
rect 3056 556232 3108 556238
rect 3056 556174 3108 556180
rect 3054 548856 3110 548865
rect 3054 548791 3110 548800
rect 3068 547942 3096 548791
rect 3056 547936 3108 547942
rect 3056 547878 3108 547884
rect 3146 544776 3202 544785
rect 3146 544711 3202 544720
rect 3160 543794 3188 544711
rect 3148 543788 3200 543794
rect 3148 543730 3200 543736
rect 3330 537296 3386 537305
rect 3330 537231 3386 537240
rect 3344 536858 3372 537231
rect 3332 536852 3384 536858
rect 3332 536794 3384 536800
rect 3330 533216 3386 533225
rect 3330 533151 3386 533160
rect 3344 532778 3372 533151
rect 3332 532772 3384 532778
rect 3332 532714 3384 532720
rect 2870 520976 2926 520985
rect 2870 520911 2926 520920
rect 2884 520334 2912 520911
rect 2872 520328 2924 520334
rect 2872 520270 2924 520276
rect 2962 516896 3018 516905
rect 2962 516831 3018 516840
rect 2976 516186 3004 516831
rect 2964 516180 3016 516186
rect 2964 516122 3016 516128
rect 3054 512816 3110 512825
rect 3054 512751 3110 512760
rect 3068 512038 3096 512751
rect 3056 512032 3108 512038
rect 3056 511974 3108 511980
rect 3054 504656 3110 504665
rect 3054 504591 3110 504600
rect 3068 503742 3096 504591
rect 3056 503736 3108 503742
rect 3056 503678 3108 503684
rect 3330 497176 3386 497185
rect 3330 497111 3386 497120
rect 3344 496874 3372 497111
rect 3332 496868 3384 496874
rect 3332 496810 3384 496816
rect 3330 489016 3386 489025
rect 3330 488951 3386 488960
rect 3344 488578 3372 488951
rect 3332 488572 3384 488578
rect 3332 488514 3384 488520
rect 2870 476776 2926 476785
rect 2870 476711 2926 476720
rect 2884 476134 2912 476711
rect 2872 476128 2924 476134
rect 2872 476070 2924 476076
rect 2870 472696 2926 472705
rect 2870 472631 2926 472640
rect 2884 472054 2912 472631
rect 2872 472048 2924 472054
rect 2872 471990 2924 471996
rect 2962 468616 3018 468625
rect 2962 468551 3018 468560
rect 2976 467906 3004 468551
rect 2964 467900 3016 467906
rect 2964 467842 3016 467848
rect 3238 457056 3294 457065
rect 3238 456991 3294 457000
rect 3252 456822 3280 456991
rect 3240 456816 3292 456822
rect 3240 456758 3292 456764
rect 3330 452976 3386 452985
rect 3330 452911 3386 452920
rect 3344 452674 3372 452911
rect 3332 452668 3384 452674
rect 3332 452610 3384 452616
rect 3330 448896 3386 448905
rect 3330 448831 3386 448840
rect 3344 448594 3372 448831
rect 3332 448588 3384 448594
rect 3332 448530 3384 448536
rect 3330 440736 3386 440745
rect 3330 440671 3386 440680
rect 3344 440298 3372 440671
rect 3332 440292 3384 440298
rect 3332 440234 3384 440240
rect 2870 428496 2926 428505
rect 2870 428431 2926 428440
rect 2884 427854 2912 428431
rect 2872 427848 2924 427854
rect 2872 427790 2924 427796
rect 3238 400616 3294 400625
rect 3238 400551 3294 400560
rect 3252 400246 3280 400551
rect 3240 400240 3292 400246
rect 3240 400182 3292 400188
rect 2962 388376 3018 388385
rect 2962 388311 3018 388320
rect 2976 387870 3004 388311
rect 2964 387864 3016 387870
rect 2964 387806 3016 387812
rect 3146 384976 3202 384985
rect 3146 384911 3202 384920
rect 3160 383722 3188 384911
rect 3148 383716 3200 383722
rect 3148 383658 3200 383664
rect 3330 380896 3386 380905
rect 3330 380831 3386 380840
rect 3344 379574 3372 380831
rect 3332 379568 3384 379574
rect 3332 379510 3384 379516
rect 3330 376816 3386 376825
rect 3330 376751 3332 376760
rect 3384 376751 3386 376760
rect 3332 376722 3384 376728
rect 3330 372736 3386 372745
rect 3330 372671 3386 372680
rect 3344 372638 3372 372671
rect 3332 372632 3384 372638
rect 3332 372574 3384 372580
rect 3330 368656 3386 368665
rect 3330 368591 3386 368600
rect 3344 368558 3372 368591
rect 3332 368552 3384 368558
rect 3332 368494 3384 368500
rect 3330 364576 3386 364585
rect 3330 364511 3332 364520
rect 3384 364511 3386 364520
rect 3332 364482 3384 364488
rect 3330 360496 3386 360505
rect 3330 360431 3386 360440
rect 3344 360262 3372 360431
rect 3332 360256 3384 360262
rect 3332 360198 3384 360204
rect 3330 356416 3386 356425
rect 3330 356351 3386 356360
rect 3344 356114 3372 356351
rect 3332 356108 3384 356114
rect 3332 356050 3384 356056
rect 3238 352336 3294 352345
rect 3238 352271 3294 352280
rect 3252 351966 3280 352271
rect 3240 351960 3292 351966
rect 3240 351902 3292 351908
rect 3146 348936 3202 348945
rect 3146 348871 3202 348880
rect 3160 347818 3188 348871
rect 3148 347812 3200 347818
rect 3148 347754 3200 347760
rect 3330 344856 3386 344865
rect 3330 344791 3386 344800
rect 3344 343670 3372 344791
rect 3332 343664 3384 343670
rect 3332 343606 3384 343612
rect 3146 340776 3202 340785
rect 3146 340711 3202 340720
rect 3160 339522 3188 340711
rect 3148 339516 3200 339522
rect 3148 339458 3200 339464
rect 3330 336696 3386 336705
rect 3330 336631 3386 336640
rect 3344 335374 3372 336631
rect 3332 335368 3384 335374
rect 3332 335310 3384 335316
rect 3332 332648 3384 332654
rect 3330 332616 3332 332625
rect 3384 332616 3386 332625
rect 3330 332551 3386 332560
rect 3330 328536 3386 328545
rect 3330 328471 3332 328480
rect 3384 328471 3386 328480
rect 3332 328442 3384 328448
rect 3330 324456 3386 324465
rect 3330 324391 3386 324400
rect 3344 324358 3372 324391
rect 3332 324352 3384 324358
rect 3332 324294 3384 324300
rect 3146 320376 3202 320385
rect 3146 320311 3202 320320
rect 3160 320210 3188 320311
rect 3148 320204 3200 320210
rect 3148 320146 3200 320152
rect 3330 316296 3386 316305
rect 3330 316231 3386 316240
rect 3344 316062 3372 316231
rect 3332 316056 3384 316062
rect 3332 315998 3384 316004
rect 3330 308816 3386 308825
rect 3330 308751 3386 308760
rect 3344 307834 3372 308751
rect 3332 307828 3384 307834
rect 3332 307770 3384 307776
rect 3054 304736 3110 304745
rect 3054 304671 3110 304680
rect 3068 303686 3096 304671
rect 3056 303680 3108 303686
rect 3056 303622 3108 303628
rect 3146 300656 3202 300665
rect 3146 300591 3202 300600
rect 3160 299538 3188 300591
rect 3148 299532 3200 299538
rect 3148 299474 3200 299480
rect 3330 296576 3386 296585
rect 3330 296511 3386 296520
rect 3344 295390 3372 296511
rect 3332 295384 3384 295390
rect 3332 295326 3384 295332
rect 3146 292496 3202 292505
rect 3146 292431 3202 292440
rect 3160 291242 3188 292431
rect 3148 291236 3200 291242
rect 3148 291178 3200 291184
rect 3330 288416 3386 288425
rect 3330 288351 3386 288360
rect 3344 287094 3372 288351
rect 3332 287088 3384 287094
rect 3332 287030 3384 287036
rect 3332 284368 3384 284374
rect 3330 284336 3332 284345
rect 3384 284336 3386 284345
rect 3330 284271 3386 284280
rect 3330 280256 3386 280265
rect 3330 280191 3332 280200
rect 3384 280191 3386 280200
rect 3332 280162 3384 280168
rect 3146 272096 3202 272105
rect 3146 272031 3202 272040
rect 3160 271930 3188 272031
rect 3148 271924 3200 271930
rect 3148 271866 3200 271872
rect 3330 264616 3386 264625
rect 3330 264551 3386 264560
rect 3344 263634 3372 264551
rect 3332 263628 3384 263634
rect 3332 263570 3384 263576
rect 3054 260536 3110 260545
rect 3054 260471 3110 260480
rect 3068 259486 3096 260471
rect 3056 259480 3108 259486
rect 3056 259422 3108 259428
rect 3146 256456 3202 256465
rect 3146 256391 3202 256400
rect 3160 255338 3188 256391
rect 3148 255332 3200 255338
rect 3148 255274 3200 255280
rect 3146 252376 3202 252385
rect 3146 252311 3202 252320
rect 3160 251258 3188 252311
rect 3148 251252 3200 251258
rect 3148 251194 3200 251200
rect 3330 248296 3386 248305
rect 3330 248231 3386 248240
rect 3344 247110 3372 248231
rect 3332 247104 3384 247110
rect 3332 247046 3384 247052
rect 3146 244216 3202 244225
rect 3146 244151 3202 244160
rect 3160 242962 3188 244151
rect 3148 242956 3200 242962
rect 3148 242898 3200 242904
rect 3330 240136 3386 240145
rect 3330 240071 3332 240080
rect 3384 240071 3386 240080
rect 3332 240042 3384 240048
rect 3330 236056 3386 236065
rect 3330 235991 3332 236000
rect 3384 235991 3386 236000
rect 3332 235962 3384 235968
rect 3330 232656 3386 232665
rect 3330 232591 3386 232600
rect 3344 231878 3372 232591
rect 3332 231872 3384 231878
rect 3332 231814 3384 231820
rect 3330 228576 3386 228585
rect 3330 228511 3386 228520
rect 3344 227798 3372 228511
rect 3332 227792 3384 227798
rect 3332 227734 3384 227740
rect 3330 224496 3386 224505
rect 3330 224431 3386 224440
rect 3344 223650 3372 224431
rect 3332 223644 3384 223650
rect 3332 223586 3384 223592
rect 3240 220788 3292 220794
rect 3240 220730 3292 220736
rect 3252 220425 3280 220730
rect 3238 220416 3294 220425
rect 3238 220351 3294 220360
rect 3330 216336 3386 216345
rect 3330 216271 3386 216280
rect 3344 215354 3372 216271
rect 3332 215348 3384 215354
rect 3332 215290 3384 215296
rect 3436 199442 3464 609311
rect 3514 601216 3570 601225
rect 3514 601151 3570 601160
rect 3528 600370 3556 601151
rect 3516 600364 3568 600370
rect 3516 600306 3568 600312
rect 3514 577416 3570 577425
rect 3514 577351 3570 577360
rect 3528 576910 3556 577351
rect 3516 576904 3568 576910
rect 3516 576846 3568 576852
rect 3514 552936 3570 552945
rect 3514 552871 3570 552880
rect 3528 552090 3556 552871
rect 3516 552084 3568 552090
rect 3516 552026 3568 552032
rect 3514 541376 3570 541385
rect 3514 541311 3570 541320
rect 3528 541006 3556 541311
rect 3516 541000 3568 541006
rect 3516 540942 3568 540948
rect 3514 529136 3570 529145
rect 3514 529071 3570 529080
rect 3528 528630 3556 529071
rect 3516 528624 3568 528630
rect 3516 528566 3568 528572
rect 3514 525056 3570 525065
rect 3514 524991 3570 525000
rect 3528 524482 3556 524991
rect 3516 524476 3568 524482
rect 3516 524418 3568 524424
rect 3514 508736 3570 508745
rect 3514 508671 3570 508680
rect 3528 507890 3556 508671
rect 3516 507884 3568 507890
rect 3516 507826 3568 507832
rect 3514 493096 3570 493105
rect 3514 493031 3570 493040
rect 3528 492726 3556 493031
rect 3516 492720 3568 492726
rect 3516 492662 3568 492668
rect 3514 484936 3570 484945
rect 3514 484871 3570 484880
rect 3528 484430 3556 484871
rect 3516 484424 3568 484430
rect 3516 484366 3568 484372
rect 3514 480856 3570 480865
rect 3514 480791 3570 480800
rect 3528 480282 3556 480791
rect 3516 480276 3568 480282
rect 3516 480218 3568 480224
rect 3514 465216 3570 465225
rect 3514 465151 3570 465160
rect 3528 465118 3556 465151
rect 3516 465112 3568 465118
rect 3516 465054 3568 465060
rect 3514 461136 3570 461145
rect 3514 461071 3570 461080
rect 3528 460970 3556 461071
rect 3516 460964 3568 460970
rect 3516 460906 3568 460912
rect 3514 444816 3570 444825
rect 3514 444751 3570 444760
rect 3528 444446 3556 444751
rect 3516 444440 3568 444446
rect 3516 444382 3568 444388
rect 3514 436656 3570 436665
rect 3514 436591 3570 436600
rect 3528 436150 3556 436591
rect 3516 436144 3568 436150
rect 3516 436086 3568 436092
rect 3514 432576 3570 432585
rect 3514 432511 3570 432520
rect 3528 432002 3556 432511
rect 3516 431996 3568 432002
rect 3516 431938 3568 431944
rect 3514 416936 3570 416945
rect 3514 416871 3570 416880
rect 3528 416838 3556 416871
rect 3516 416832 3568 416838
rect 3516 416774 3568 416780
rect 3514 412856 3570 412865
rect 3514 412791 3570 412800
rect 3528 412690 3556 412791
rect 3516 412684 3568 412690
rect 3516 412626 3568 412632
rect 3514 408776 3570 408785
rect 3514 408711 3570 408720
rect 3528 408542 3556 408711
rect 3516 408536 3568 408542
rect 3516 408478 3568 408484
rect 3514 404696 3570 404705
rect 3514 404631 3570 404640
rect 3528 200802 3556 404631
rect 3606 396536 3662 396545
rect 3606 396471 3662 396480
rect 3620 396098 3648 396471
rect 3608 396092 3660 396098
rect 3608 396034 3660 396040
rect 7564 364540 7616 364546
rect 7564 364482 7616 364488
rect 7576 271182 7604 364482
rect 7564 271176 7616 271182
rect 7564 271118 7616 271124
rect 3516 200796 3568 200802
rect 3516 200738 3568 200744
rect 3514 200016 3570 200025
rect 3514 199951 3570 199960
rect 3424 199436 3476 199442
rect 3424 199378 3476 199384
rect 3528 198830 3556 199951
rect 3516 198824 3568 198830
rect 3516 198766 3568 198772
rect 3608 196104 3660 196110
rect 3608 196046 3660 196052
rect 3516 196036 3568 196042
rect 3516 195978 3568 195984
rect 3422 195936 3478 195945
rect 3422 195871 3478 195880
rect 3436 195362 3464 195871
rect 3424 195356 3476 195362
rect 3424 195298 3476 195304
rect 3422 192536 3478 192545
rect 3422 192471 3478 192480
rect 3238 188456 3294 188465
rect 3238 188391 3294 188400
rect 3252 188086 3280 188391
rect 3240 188080 3292 188086
rect 3240 188022 3292 188028
rect 3146 184376 3202 184385
rect 3146 184311 3202 184320
rect 3160 184210 3188 184311
rect 3148 184204 3200 184210
rect 3148 184146 3200 184152
rect 3240 180804 3292 180810
rect 3240 180746 3292 180752
rect 3252 180305 3280 180746
rect 3238 180296 3294 180305
rect 3238 180231 3294 180240
rect 3240 172508 3292 172514
rect 3240 172450 3292 172456
rect 3252 172145 3280 172450
rect 3238 172136 3294 172145
rect 3238 172071 3294 172080
rect 3332 168360 3384 168366
rect 3332 168302 3384 168308
rect 3344 168065 3372 168302
rect 3330 168056 3386 168065
rect 3330 167991 3386 168000
rect 3054 163976 3110 163985
rect 3054 163911 3110 163920
rect 3068 162926 3096 163911
rect 3056 162920 3108 162926
rect 3056 162862 3108 162868
rect 3436 147626 3464 192471
rect 3528 156074 3556 195978
rect 3620 159905 3648 196046
rect 4896 190528 4948 190534
rect 4896 190470 4948 190476
rect 3606 159896 3662 159905
rect 3606 159831 3662 159840
rect 3528 156046 3648 156074
rect 3516 155916 3568 155922
rect 3516 155858 3568 155864
rect 3528 155825 3556 155858
rect 3514 155816 3570 155825
rect 3514 155751 3570 155760
rect 3620 152425 3648 156046
rect 3606 152416 3662 152425
rect 3606 152351 3662 152360
rect 3424 147620 3476 147626
rect 3424 147562 3476 147568
rect 3148 144900 3200 144906
rect 3148 144842 3200 144848
rect 3160 144265 3188 144842
rect 3146 144256 3202 144265
rect 3146 144191 3202 144200
rect 3608 141432 3660 141438
rect 3608 141374 3660 141380
rect 2780 140684 2832 140690
rect 2780 140626 2832 140632
rect 2792 140185 2820 140626
rect 2778 140176 2834 140185
rect 2778 140111 2834 140120
rect 3516 136604 3568 136610
rect 3516 136546 3568 136552
rect 3528 136105 3556 136546
rect 3514 136096 3570 136105
rect 3514 136031 3570 136040
rect 3332 132456 3384 132462
rect 3332 132398 3384 132404
rect 3344 132025 3372 132398
rect 3330 132016 3386 132025
rect 3330 131951 3386 131960
rect 3422 127936 3478 127945
rect 3422 127871 3478 127880
rect 3436 127634 3464 127871
rect 3424 127628 3476 127634
rect 3424 127570 3476 127576
rect 3422 123856 3478 123865
rect 3422 123791 3478 123800
rect 3436 122874 3464 123791
rect 3424 122868 3476 122874
rect 3620 122834 3648 141374
rect 4908 140690 4936 190470
rect 8312 186318 8340 683086
rect 13084 636268 13136 636274
rect 13084 636210 13136 636216
rect 10324 295384 10376 295390
rect 10324 295326 10376 295332
rect 10336 269822 10364 295326
rect 13096 278050 13124 636210
rect 13084 278044 13136 278050
rect 13084 277986 13136 277992
rect 14476 273970 14504 688638
rect 21364 616888 21416 616894
rect 21364 616830 21416 616836
rect 14464 273964 14516 273970
rect 14464 273906 14516 273912
rect 10324 269816 10376 269822
rect 10324 269758 10376 269764
rect 21376 267034 21404 616830
rect 21364 267028 21416 267034
rect 21364 266970 21416 266976
rect 26896 199481 26924 700538
rect 27724 683114 27752 703520
rect 31588 703050 31616 703520
rect 30380 703044 30432 703050
rect 30380 702986 30432 702992
rect 31576 703044 31628 703050
rect 31576 702986 31628 702992
rect 27632 683086 27752 683114
rect 26882 199472 26938 199481
rect 26882 199407 26938 199416
rect 25504 191888 25556 191894
rect 25504 191830 25556 191836
rect 8300 186312 8352 186318
rect 8300 186254 8352 186260
rect 25516 168366 25544 191830
rect 27632 188358 27660 683086
rect 27620 188352 27672 188358
rect 27620 188294 27672 188300
rect 30392 186250 30420 702986
rect 34808 702434 34836 703520
rect 34532 702406 34836 702434
rect 34532 264246 34560 702406
rect 34520 264240 34572 264246
rect 34520 264182 34572 264188
rect 38672 262886 38700 703520
rect 42536 699718 42564 703520
rect 46400 700602 46428 703520
rect 46388 700596 46440 700602
rect 46388 700538 46440 700544
rect 48964 700528 49016 700534
rect 48964 700470 49016 700476
rect 42524 699712 42576 699718
rect 42524 699654 42576 699660
rect 43444 699712 43496 699718
rect 43444 699654 43496 699660
rect 38660 262880 38712 262886
rect 38660 262822 38712 262828
rect 43456 199753 43484 699654
rect 48976 200705 49004 700470
rect 48962 200696 49018 200705
rect 48962 200631 49018 200640
rect 43442 199744 43498 199753
rect 43442 199679 43498 199688
rect 49712 188154 49740 703582
rect 50080 703474 50108 703582
rect 50222 703520 50334 704960
rect 54086 703520 54198 704960
rect 57950 703520 58062 704960
rect 60752 703582 61700 703610
rect 50264 703474 50292 703520
rect 50080 703446 50292 703474
rect 54128 700534 54156 703520
rect 54116 700528 54168 700534
rect 54116 700470 54168 700476
rect 53104 261044 53156 261050
rect 53104 260986 53156 260992
rect 53116 240106 53144 260986
rect 53104 240100 53156 240106
rect 53104 240042 53156 240048
rect 57992 191758 58020 703520
rect 57980 191752 58032 191758
rect 57980 191694 58032 191700
rect 60752 190369 60780 703582
rect 61672 703474 61700 703582
rect 61814 703520 61926 704960
rect 65678 703520 65790 704960
rect 68898 703520 69010 704960
rect 72762 703520 72874 704960
rect 76626 703520 76738 704960
rect 80490 703520 80602 704960
rect 84354 703520 84466 704960
rect 88218 703520 88330 704960
rect 92082 703520 92194 704960
rect 95946 703520 96058 704960
rect 99810 703520 99922 704960
rect 103674 703520 103786 704960
rect 106292 703582 106780 703610
rect 61856 703474 61884 703520
rect 61672 703446 61884 703474
rect 65720 700670 65748 703520
rect 65708 700664 65760 700670
rect 65708 700606 65760 700612
rect 62764 698964 62816 698970
rect 62764 698906 62816 698912
rect 62776 198014 62804 698906
rect 68940 697610 68968 703520
rect 72804 702434 72832 703520
rect 76668 702434 76696 703520
rect 71792 702406 72832 702434
rect 75932 702406 76696 702434
rect 67640 697604 67692 697610
rect 67640 697546 67692 697552
rect 68928 697604 68980 697610
rect 68928 697546 68980 697552
rect 64144 612808 64196 612814
rect 64144 612750 64196 612756
rect 62764 198008 62816 198014
rect 62764 197950 62816 197956
rect 60738 190360 60794 190369
rect 60738 190295 60794 190304
rect 49700 188148 49752 188154
rect 49700 188090 49752 188096
rect 30380 186244 30432 186250
rect 30380 186186 30432 186192
rect 25504 168360 25556 168366
rect 25504 168302 25556 168308
rect 64156 145625 64184 612750
rect 67652 265674 67680 697546
rect 67640 265668 67692 265674
rect 67640 265610 67692 265616
rect 71792 199510 71820 702406
rect 75932 199578 75960 702406
rect 80532 700670 80560 703520
rect 79324 700664 79376 700670
rect 79324 700606 79376 700612
rect 80520 700664 80572 700670
rect 80520 700606 80572 700612
rect 79336 200841 79364 700606
rect 84396 683114 84424 703520
rect 88260 700738 88288 703520
rect 92124 702434 92152 703520
rect 91112 702406 92152 702434
rect 88248 700732 88300 700738
rect 88248 700674 88300 700680
rect 88984 700664 89036 700670
rect 88984 700606 89036 700612
rect 84212 683086 84424 683114
rect 80704 592068 80756 592074
rect 80704 592010 80756 592016
rect 79416 396092 79468 396098
rect 79416 396034 79468 396040
rect 79428 268394 79456 396034
rect 79416 268388 79468 268394
rect 79416 268330 79468 268336
rect 79322 200832 79378 200841
rect 79322 200767 79378 200776
rect 75920 199572 75972 199578
rect 75920 199514 75972 199520
rect 71780 199504 71832 199510
rect 71780 199446 71832 199452
rect 80716 180334 80744 592010
rect 80796 576904 80848 576910
rect 80796 576846 80848 576852
rect 80808 191185 80836 576846
rect 84212 194585 84240 683086
rect 86224 661088 86276 661094
rect 86224 661030 86276 661036
rect 84844 583772 84896 583778
rect 84844 583714 84896 583720
rect 84198 194576 84254 194585
rect 84198 194511 84254 194520
rect 80794 191176 80850 191185
rect 80794 191111 80850 191120
rect 84856 183394 84884 583714
rect 84936 552084 84988 552090
rect 84936 552026 84988 552032
rect 84948 191146 84976 552026
rect 84936 191140 84988 191146
rect 84936 191082 84988 191088
rect 84844 183388 84896 183394
rect 84844 183330 84896 183336
rect 80704 180328 80756 180334
rect 80704 180270 80756 180276
rect 86236 180266 86264 661030
rect 86316 524476 86368 524482
rect 86316 524418 86368 524424
rect 86328 192506 86356 524418
rect 87604 472048 87656 472054
rect 87604 471990 87656 471996
rect 86316 192500 86368 192506
rect 86316 192442 86368 192448
rect 87616 185910 87644 471990
rect 87696 387864 87748 387870
rect 87696 387806 87748 387812
rect 87604 185904 87656 185910
rect 87604 185846 87656 185852
rect 86224 180260 86276 180266
rect 86224 180202 86276 180208
rect 87708 178906 87736 387806
rect 88996 199646 89024 700606
rect 89076 644496 89128 644502
rect 89076 644438 89128 644444
rect 88984 199640 89036 199646
rect 88984 199582 89036 199588
rect 89088 192953 89116 644438
rect 90364 632120 90416 632126
rect 90364 632062 90416 632068
rect 89074 192944 89130 192953
rect 89074 192879 89130 192888
rect 90376 189786 90404 632062
rect 90456 581052 90508 581058
rect 90456 580994 90508 581000
rect 90364 189780 90416 189786
rect 90364 189722 90416 189728
rect 90468 184822 90496 580994
rect 90548 492720 90600 492726
rect 90548 492662 90600 492668
rect 90456 184816 90508 184822
rect 90456 184758 90508 184764
rect 90560 184754 90588 492662
rect 90640 376780 90692 376786
rect 90640 376722 90692 376728
rect 90652 187542 90680 376722
rect 91112 195945 91140 702406
rect 95988 700670 96016 703520
rect 99852 702434 99880 703520
rect 99392 702406 99880 702434
rect 95976 700664 96028 700670
rect 95976 700606 96028 700612
rect 98736 700596 98788 700602
rect 98736 700538 98788 700544
rect 98644 696992 98696 696998
rect 98644 696934 98696 696940
rect 93124 684548 93176 684554
rect 93124 684490 93176 684496
rect 92480 227792 92532 227798
rect 92478 227760 92480 227769
rect 92532 227760 92534 227769
rect 92478 227695 92534 227704
rect 92480 200796 92532 200802
rect 92480 200738 92532 200744
rect 92492 200190 92520 200738
rect 92480 200184 92532 200190
rect 92480 200126 92532 200132
rect 91098 195936 91154 195945
rect 91098 195871 91154 195880
rect 93136 191729 93164 684490
rect 93308 676252 93360 676258
rect 93308 676194 93360 676200
rect 93216 465112 93268 465118
rect 93216 465054 93268 465060
rect 93122 191720 93178 191729
rect 93122 191655 93178 191664
rect 93228 188698 93256 465054
rect 93320 191049 93348 676194
rect 94504 640348 94556 640354
rect 94504 640290 94556 640296
rect 93400 431996 93452 432002
rect 93400 431938 93452 431944
rect 93306 191040 93362 191049
rect 93306 190975 93362 190984
rect 93216 188692 93268 188698
rect 93216 188634 93268 188640
rect 90640 187536 90692 187542
rect 90640 187478 90692 187484
rect 93412 186114 93440 431938
rect 93766 227760 93822 227769
rect 93766 227695 93822 227704
rect 93676 200184 93728 200190
rect 93676 200126 93728 200132
rect 93400 186108 93452 186114
rect 93400 186050 93452 186056
rect 90548 184748 90600 184754
rect 90548 184690 90600 184696
rect 87696 178900 87748 178906
rect 87696 178842 87748 178848
rect 64142 145616 64198 145625
rect 64142 145551 64198 145560
rect 82820 142996 82872 143002
rect 82820 142938 82872 142944
rect 44180 142860 44232 142866
rect 44180 142802 44232 142808
rect 4896 140684 4948 140690
rect 4896 140626 4948 140632
rect 4804 139460 4856 139466
rect 4804 139402 4856 139408
rect 3424 122810 3476 122816
rect 3528 122806 3648 122834
rect 3332 120080 3384 120086
rect 3332 120022 3384 120028
rect 3344 119785 3372 120022
rect 3330 119776 3386 119785
rect 3330 119711 3386 119720
rect 3424 116612 3476 116618
rect 3424 116554 3476 116560
rect 3330 112296 3386 112305
rect 3330 112231 3386 112240
rect 3344 111858 3372 112231
rect 3332 111852 3384 111858
rect 3332 111794 3384 111800
rect 3056 108996 3108 109002
rect 3056 108938 3108 108944
rect 3068 108225 3096 108938
rect 3054 108216 3110 108225
rect 3054 108151 3110 108160
rect 2964 104848 3016 104854
rect 2964 104790 3016 104796
rect 2976 104145 3004 104790
rect 2962 104136 3018 104145
rect 2962 104071 3018 104080
rect 2870 100056 2926 100065
rect 2870 99991 2926 100000
rect 2884 99414 2912 99991
rect 2872 99408 2924 99414
rect 2872 99350 2924 99356
rect 2962 95976 3018 95985
rect 2962 95911 3018 95920
rect 2976 95266 3004 95911
rect 2964 95260 3016 95266
rect 2964 95202 3016 95208
rect 3054 91896 3110 91905
rect 3054 91831 3110 91840
rect 3068 91118 3096 91831
rect 3056 91112 3108 91118
rect 3056 91054 3108 91060
rect 2872 76900 2924 76906
rect 2872 76842 2924 76848
rect 2884 76265 2912 76842
rect 2870 76256 2926 76265
rect 2870 76191 2926 76200
rect 3148 73160 3200 73166
rect 3148 73102 3200 73108
rect 3160 72185 3188 73102
rect 3146 72176 3202 72185
rect 3146 72111 3202 72120
rect 2780 71052 2832 71058
rect 2780 70994 2832 71000
rect 2792 16574 2820 70994
rect 3148 37256 3200 37262
rect 3148 37198 3200 37204
rect 3160 36145 3188 37198
rect 3146 36136 3202 36145
rect 3146 36071 3202 36080
rect 3148 28960 3200 28966
rect 3148 28902 3200 28908
rect 3160 27985 3188 28902
rect 3146 27976 3202 27985
rect 3146 27911 3202 27920
rect 3436 23905 3464 116554
rect 3528 116385 3556 122806
rect 3514 116376 3570 116385
rect 3514 116311 3570 116320
rect 3516 88324 3568 88330
rect 3516 88266 3568 88272
rect 3528 87825 3556 88266
rect 3514 87816 3570 87825
rect 3514 87751 3570 87760
rect 3514 83736 3570 83745
rect 3514 83671 3570 83680
rect 3528 82890 3556 83671
rect 3516 82884 3568 82890
rect 3516 82826 3568 82832
rect 3516 79688 3568 79694
rect 3514 79656 3516 79665
rect 3568 79656 3570 79665
rect 3514 79591 3570 79600
rect 3516 68196 3568 68202
rect 3516 68138 3568 68144
rect 3528 68105 3556 68138
rect 3514 68096 3570 68105
rect 3514 68031 3570 68040
rect 3516 60716 3568 60722
rect 3516 60658 3568 60664
rect 3528 59945 3556 60658
rect 3514 59936 3570 59945
rect 3514 59871 3570 59880
rect 3516 52420 3568 52426
rect 3516 52362 3568 52368
rect 3528 51785 3556 52362
rect 3514 51776 3570 51785
rect 3514 51711 3570 51720
rect 3516 48272 3568 48278
rect 3516 48214 3568 48220
rect 3528 47705 3556 48214
rect 3514 47696 3570 47705
rect 3514 47631 3570 47640
rect 3516 44124 3568 44130
rect 3516 44066 3568 44072
rect 3528 43625 3556 44066
rect 3514 43616 3570 43625
rect 3514 43551 3570 43560
rect 3516 40044 3568 40050
rect 3516 39986 3568 39992
rect 3528 39545 3556 39986
rect 3514 39536 3570 39545
rect 3514 39471 3570 39480
rect 3422 23896 3478 23905
rect 3422 23831 3478 23840
rect 3148 20664 3200 20670
rect 3148 20606 3200 20612
rect 3160 19825 3188 20606
rect 3146 19816 3202 19825
rect 3146 19751 3202 19760
rect 3332 16584 3384 16590
rect 2792 16546 3280 16574
rect 3056 12436 3108 12442
rect 3056 12378 3108 12384
rect 3068 11665 3096 12378
rect 3054 11656 3110 11665
rect 3054 11591 3110 11600
rect 2964 8288 3016 8294
rect 2964 8230 3016 8236
rect 2976 7585 3004 8230
rect 2962 7576 3018 7585
rect 2962 7511 3018 7520
rect 2780 4072 2832 4078
rect 2780 4014 2832 4020
rect 2792 3505 2820 4014
rect 2778 3496 2834 3505
rect 20 3460 72 3466
rect 2778 3431 2834 3440
rect 20 3402 72 3408
rect 32 480 60 3402
rect 3252 480 3280 16546
rect 3332 16526 3384 16532
rect 3344 15745 3372 16526
rect 3330 15736 3386 15745
rect 3330 15671 3386 15680
rect 4816 4078 4844 139402
rect 40040 75200 40092 75206
rect 40040 75142 40092 75148
rect 35164 73840 35216 73846
rect 35164 73782 35216 73788
rect 13084 69760 13136 69766
rect 13084 69702 13136 69708
rect 8944 62824 8996 62830
rect 8944 62766 8996 62772
rect 6920 61396 6972 61402
rect 6920 61338 6972 61344
rect 6932 16574 6960 61338
rect 8956 52426 8984 62766
rect 8944 52420 8996 52426
rect 8944 52362 8996 52368
rect 6932 16546 7144 16574
rect 4804 4072 4856 4078
rect 4804 4014 4856 4020
rect 7116 480 7144 16546
rect 13096 3466 13124 69702
rect 26240 66904 26292 66910
rect 26240 66846 26292 66852
rect 17960 55956 18012 55962
rect 17960 55898 18012 55904
rect 17972 16574 18000 55898
rect 26252 16574 26280 66846
rect 31024 58744 31076 58750
rect 31024 58686 31076 58692
rect 17972 16546 18736 16574
rect 26252 16546 26464 16574
rect 13084 3460 13136 3466
rect 13084 3402 13136 3408
rect 14832 3460 14884 3466
rect 14832 3402 14884 3408
rect 14844 480 14872 3402
rect 18708 480 18736 16546
rect 26436 480 26464 16546
rect 31036 3534 31064 58686
rect 35176 3534 35204 73782
rect 40052 16574 40080 75142
rect 44192 16574 44220 142802
rect 74540 73908 74592 73914
rect 74540 73850 74592 73856
rect 52460 72480 52512 72486
rect 52460 72422 52512 72428
rect 48320 54528 48372 54534
rect 48320 54470 48372 54476
rect 48332 16574 48360 54470
rect 40052 16546 40816 16574
rect 44192 16546 44680 16574
rect 48332 16546 48544 16574
rect 30288 3528 30340 3534
rect 30288 3470 30340 3476
rect 31024 3528 31076 3534
rect 31024 3470 31076 3476
rect 34152 3528 34204 3534
rect 34152 3470 34204 3476
rect 35164 3528 35216 3534
rect 35164 3470 35216 3476
rect 30300 480 30328 3470
rect 34164 480 34192 3470
rect -10 -960 102 480
rect 3210 -960 3322 480
rect 7074 -960 7186 480
rect 10938 -960 11050 480
rect 14802 -960 14914 480
rect 18666 -960 18778 480
rect 22530 -960 22642 480
rect 26394 -960 26506 480
rect 30258 -960 30370 480
rect 34122 -960 34234 480
rect 37342 -960 37454 480
rect 40788 354 40816 16546
rect 41206 354 41318 480
rect 40788 326 41318 354
rect 44652 354 44680 16546
rect 45070 354 45182 480
rect 44652 326 45182 354
rect 48516 354 48544 16546
rect 48934 354 49046 480
rect 48516 326 49046 354
rect 52472 354 52500 72422
rect 67640 65544 67692 65550
rect 67640 65486 67692 65492
rect 63500 64184 63552 64190
rect 63500 64126 63552 64132
rect 63512 16574 63540 64126
rect 67652 16574 67680 65486
rect 71780 57248 71832 57254
rect 71780 57190 71832 57196
rect 63512 16546 64000 16574
rect 67652 16546 67864 16574
rect 52798 354 52910 480
rect 52472 326 52910 354
rect 41206 -960 41318 326
rect 45070 -960 45182 326
rect 48934 -960 49046 326
rect 52798 -960 52910 326
rect 56662 -960 56774 480
rect 60526 -960 60638 480
rect 63972 354 64000 16546
rect 64390 354 64502 480
rect 63972 326 64502 354
rect 67836 354 67864 16546
rect 68254 354 68366 480
rect 67836 326 68366 354
rect 71792 354 71820 57190
rect 74552 16574 74580 73850
rect 78680 69692 78732 69698
rect 78680 69634 78732 69640
rect 78692 16574 78720 69634
rect 82832 16574 82860 142938
rect 93688 75002 93716 200126
rect 93676 74996 93728 75002
rect 93676 74938 93728 74944
rect 93780 70990 93808 227695
rect 94516 186153 94544 640290
rect 94596 568608 94648 568614
rect 94596 568550 94648 568556
rect 94608 190466 94636 568550
rect 97264 556232 97316 556238
rect 97264 556174 97316 556180
rect 94688 541000 94740 541006
rect 94688 540942 94740 540948
rect 94700 197402 94728 540942
rect 95884 528624 95936 528630
rect 95884 528566 95936 528572
rect 94780 383716 94832 383722
rect 94780 383658 94832 383664
rect 94688 197396 94740 197402
rect 94688 197338 94740 197344
rect 94792 192302 94820 383658
rect 95700 197464 95752 197470
rect 95700 197406 95752 197412
rect 95608 193996 95660 194002
rect 95608 193938 95660 193944
rect 94780 192296 94832 192302
rect 94780 192238 94832 192244
rect 94596 190460 94648 190466
rect 94596 190402 94648 190408
rect 94502 186144 94558 186153
rect 94502 186079 94558 186088
rect 95148 178084 95200 178090
rect 95148 178026 95200 178032
rect 94964 151224 95016 151230
rect 94964 151166 95016 151172
rect 93768 70984 93820 70990
rect 93768 70926 93820 70932
rect 94976 69766 95004 151166
rect 95056 151088 95108 151094
rect 95056 151030 95108 151036
rect 94964 69760 95016 69766
rect 94964 69702 95016 69708
rect 93860 67040 93912 67046
rect 93860 66982 93912 66988
rect 89720 66632 89772 66638
rect 89720 66574 89772 66580
rect 89732 16574 89760 66574
rect 93872 16574 93900 66982
rect 95068 55214 95096 151030
rect 95160 76537 95188 178026
rect 95620 80714 95648 193938
rect 95608 80708 95660 80714
rect 95608 80650 95660 80656
rect 95146 76528 95202 76537
rect 95146 76463 95202 76472
rect 95712 74934 95740 197406
rect 95896 191554 95924 528566
rect 95976 507884 96028 507890
rect 95976 507826 96028 507832
rect 95884 191548 95936 191554
rect 95884 191490 95936 191496
rect 95988 189854 96016 507826
rect 96068 351960 96120 351966
rect 96068 351902 96120 351908
rect 95976 189848 96028 189854
rect 95976 189790 96028 189796
rect 95976 188556 96028 188562
rect 95976 188498 96028 188504
rect 95884 151156 95936 151162
rect 95884 151098 95936 151104
rect 95792 143676 95844 143682
rect 95792 143618 95844 143624
rect 95804 120086 95832 143618
rect 95792 120080 95844 120086
rect 95792 120022 95844 120028
rect 95700 74928 95752 74934
rect 95700 74870 95752 74876
rect 95148 69760 95200 69766
rect 95148 69702 95200 69708
rect 95160 69562 95188 69702
rect 95148 69556 95200 69562
rect 95148 69498 95200 69504
rect 95896 68338 95924 151098
rect 95988 78878 96016 188498
rect 96080 186998 96108 351902
rect 96160 324352 96212 324358
rect 96160 324294 96212 324300
rect 96172 187474 96200 324294
rect 96528 247104 96580 247110
rect 96528 247046 96580 247052
rect 96436 215348 96488 215354
rect 96436 215290 96488 215296
rect 96344 201544 96396 201550
rect 96344 201486 96396 201492
rect 96252 195424 96304 195430
rect 96252 195366 96304 195372
rect 96160 187468 96212 187474
rect 96160 187410 96212 187416
rect 96068 186992 96120 186998
rect 96068 186934 96120 186940
rect 95976 78872 96028 78878
rect 95976 78814 96028 78820
rect 95884 68332 95936 68338
rect 95884 68274 95936 68280
rect 96264 62082 96292 195366
rect 96356 64734 96384 201486
rect 96344 64728 96396 64734
rect 96344 64670 96396 64676
rect 96448 63442 96476 215290
rect 96540 182918 96568 247046
rect 96988 201612 97040 201618
rect 96988 201554 97040 201560
rect 96528 182912 96580 182918
rect 96528 182854 96580 182860
rect 96528 148368 96580 148374
rect 96528 148310 96580 148316
rect 96540 78674 96568 148310
rect 97000 81977 97028 201554
rect 97080 189780 97132 189786
rect 97080 189722 97132 189728
rect 96986 81968 97042 81977
rect 96986 81903 97042 81912
rect 96528 78668 96580 78674
rect 96528 78610 96580 78616
rect 97092 71777 97120 189722
rect 97276 184686 97304 556174
rect 97356 536852 97408 536858
rect 97356 536794 97408 536800
rect 97264 184680 97316 184686
rect 97264 184622 97316 184628
rect 97368 184006 97396 536794
rect 97448 516180 97500 516186
rect 97448 516122 97500 516128
rect 97460 186794 97488 516122
rect 97540 368552 97592 368558
rect 97540 368494 97592 368500
rect 97448 186788 97500 186794
rect 97448 186730 97500 186736
rect 97552 185842 97580 368494
rect 97724 196716 97776 196722
rect 97724 196658 97776 196664
rect 97540 185836 97592 185842
rect 97540 185778 97592 185784
rect 97356 184000 97408 184006
rect 97356 183942 97408 183948
rect 97448 163532 97500 163538
rect 97448 163474 97500 163480
rect 97460 162926 97488 163474
rect 97448 162920 97500 162926
rect 97448 162862 97500 162868
rect 97356 142928 97408 142934
rect 97356 142870 97408 142876
rect 97264 141500 97316 141506
rect 97264 141442 97316 141448
rect 97172 91112 97224 91118
rect 97172 91054 97224 91060
rect 97184 77246 97212 91054
rect 97172 77240 97224 77246
rect 97172 77182 97224 77188
rect 97078 71768 97134 71777
rect 97078 71703 97134 71712
rect 97276 64122 97304 141442
rect 97264 64116 97316 64122
rect 97264 64058 97316 64064
rect 97368 64054 97396 142870
rect 97460 75818 97488 162862
rect 97632 83224 97684 83230
rect 97632 83166 97684 83172
rect 97644 82890 97672 83166
rect 97632 82884 97684 82890
rect 97632 82826 97684 82832
rect 97448 75812 97500 75818
rect 97448 75754 97500 75760
rect 97644 74458 97672 82826
rect 97632 74452 97684 74458
rect 97632 74394 97684 74400
rect 97736 67425 97764 196658
rect 97816 195492 97868 195498
rect 97816 195434 97868 195440
rect 97722 67416 97778 67425
rect 97722 67351 97778 67360
rect 97356 64048 97408 64054
rect 97356 63990 97408 63996
rect 97828 63510 97856 195434
rect 98656 191321 98684 696934
rect 98748 200977 98776 700538
rect 98828 547936 98880 547942
rect 98828 547878 98880 547884
rect 98734 200968 98790 200977
rect 98734 200903 98790 200912
rect 98840 195566 98868 547878
rect 98920 356108 98972 356114
rect 98920 356050 98972 356056
rect 98828 195560 98880 195566
rect 98828 195502 98880 195508
rect 98642 191312 98698 191321
rect 98642 191247 98698 191256
rect 98932 185706 98960 356050
rect 99012 328500 99064 328506
rect 99012 328442 99064 328448
rect 99024 191622 99052 328442
rect 99104 280220 99156 280226
rect 99104 280162 99156 280168
rect 99012 191616 99064 191622
rect 99012 191558 99064 191564
rect 99116 190398 99144 280162
rect 99196 198008 99248 198014
rect 99196 197950 99248 197956
rect 99104 190392 99156 190398
rect 99104 190334 99156 190340
rect 98920 185700 98972 185706
rect 98920 185642 98972 185648
rect 99104 181552 99156 181558
rect 99104 181494 99156 181500
rect 99012 175976 99064 175982
rect 99012 175918 99064 175924
rect 98828 148708 98880 148714
rect 98828 148650 98880 148656
rect 98736 148504 98788 148510
rect 98736 148446 98788 148452
rect 98000 143132 98052 143138
rect 98000 143074 98052 143080
rect 97908 142180 97960 142186
rect 97908 142122 97960 142128
rect 97816 63504 97868 63510
rect 97816 63446 97868 63452
rect 96436 63436 96488 63442
rect 96436 63378 96488 63384
rect 97828 62830 97856 63446
rect 97816 62824 97868 62830
rect 97816 62766 97868 62772
rect 96068 62076 96120 62082
rect 96068 62018 96120 62024
rect 96252 62076 96304 62082
rect 96252 62018 96304 62024
rect 96080 61402 96108 62018
rect 96068 61396 96120 61402
rect 96068 61338 96120 61344
rect 95056 55208 95108 55214
rect 95056 55150 95108 55156
rect 95068 54534 95096 55150
rect 95056 54528 95108 54534
rect 95056 54470 95108 54476
rect 74552 16546 75408 16574
rect 78692 16546 79272 16574
rect 82832 16546 83136 16574
rect 89732 16546 90864 16574
rect 93872 16546 94728 16574
rect 75380 480 75408 16546
rect 79244 480 79272 16546
rect 83108 480 83136 16546
rect 90836 480 90864 16546
rect 94700 480 94728 16546
rect 97920 3534 97948 142122
rect 98012 16574 98040 143074
rect 98644 141568 98696 141574
rect 98644 141510 98696 141516
rect 98656 83230 98684 141510
rect 98644 83224 98696 83230
rect 98644 83166 98696 83172
rect 98748 72282 98776 148446
rect 98840 72486 98868 148650
rect 98920 148640 98972 148646
rect 98920 148582 98972 148588
rect 98828 72480 98880 72486
rect 98828 72422 98880 72428
rect 98840 72350 98868 72422
rect 98828 72344 98880 72350
rect 98828 72286 98880 72292
rect 98736 72276 98788 72282
rect 98736 72218 98788 72224
rect 98932 66026 98960 148582
rect 99024 69970 99052 175918
rect 99012 69964 99064 69970
rect 99012 69906 99064 69912
rect 98920 66020 98972 66026
rect 98920 65962 98972 65968
rect 99116 64666 99144 181494
rect 99208 68678 99236 197950
rect 99288 197396 99340 197402
rect 99288 197338 99340 197344
rect 99196 68672 99248 68678
rect 99196 68614 99248 68620
rect 99300 67153 99328 197338
rect 99392 193866 99420 702406
rect 102784 700732 102836 700738
rect 102784 700674 102836 700680
rect 100116 700392 100168 700398
rect 100116 700334 100168 700340
rect 100024 700324 100076 700330
rect 100024 700266 100076 700272
rect 99380 193860 99432 193866
rect 99380 193802 99432 193808
rect 99748 188352 99800 188358
rect 99748 188294 99800 188300
rect 99656 187264 99708 187270
rect 99656 187206 99708 187212
rect 99668 75886 99696 187206
rect 99760 78402 99788 188294
rect 100036 183530 100064 700266
rect 100128 185774 100156 700334
rect 101404 480276 101456 480282
rect 101404 480218 101456 480224
rect 100208 467900 100260 467906
rect 100208 467842 100260 467848
rect 100220 186046 100248 467842
rect 100668 198212 100720 198218
rect 100668 198154 100720 198160
rect 100576 198076 100628 198082
rect 100576 198018 100628 198024
rect 100484 191412 100536 191418
rect 100484 191354 100536 191360
rect 100496 190534 100524 191354
rect 100484 190528 100536 190534
rect 100484 190470 100536 190476
rect 100208 186040 100260 186046
rect 100208 185982 100260 185988
rect 100116 185768 100168 185774
rect 100116 185710 100168 185716
rect 100300 185632 100352 185638
rect 100300 185574 100352 185580
rect 100024 183524 100076 183530
rect 100024 183466 100076 183472
rect 100024 151292 100076 151298
rect 100024 151234 100076 151240
rect 99932 148572 99984 148578
rect 99932 148514 99984 148520
rect 99838 148472 99894 148481
rect 99838 148407 99894 148416
rect 99748 78396 99800 78402
rect 99748 78338 99800 78344
rect 99656 75880 99708 75886
rect 99656 75822 99708 75828
rect 99852 69601 99880 148407
rect 99838 69592 99894 69601
rect 99838 69527 99894 69536
rect 99286 67144 99342 67153
rect 99286 67079 99342 67088
rect 99104 64660 99156 64666
rect 99104 64602 99156 64608
rect 99944 64530 99972 148514
rect 100036 65346 100064 151234
rect 100312 73846 100340 185574
rect 100392 178832 100444 178838
rect 100392 178774 100444 178780
rect 100300 73840 100352 73846
rect 100300 73782 100352 73788
rect 100312 73642 100340 73782
rect 100300 73636 100352 73642
rect 100300 73578 100352 73584
rect 100404 66094 100432 178774
rect 100392 66088 100444 66094
rect 100392 66030 100444 66036
rect 100024 65340 100076 65346
rect 100024 65282 100076 65288
rect 100496 65278 100524 190470
rect 100588 65822 100616 198018
rect 100576 65816 100628 65822
rect 100576 65758 100628 65764
rect 100484 65272 100536 65278
rect 100484 65214 100536 65220
rect 100680 64598 100708 198154
rect 101416 191690 101444 480218
rect 101496 332648 101548 332654
rect 101496 332590 101548 332596
rect 101508 191826 101536 332590
rect 101588 284368 101640 284374
rect 101588 284310 101640 284316
rect 101496 191820 101548 191826
rect 101496 191762 101548 191768
rect 101404 191684 101456 191690
rect 101404 191626 101456 191632
rect 101600 188290 101628 284310
rect 101680 259480 101732 259486
rect 101680 259422 101732 259428
rect 101692 188426 101720 259422
rect 102796 199617 102824 700674
rect 103716 683114 103744 703520
rect 103532 683086 103744 683114
rect 102876 623824 102928 623830
rect 102876 623766 102928 623772
rect 102782 199608 102838 199617
rect 102782 199543 102838 199552
rect 102888 197033 102916 623766
rect 102968 476128 103020 476134
rect 102968 476070 103020 476076
rect 102874 197024 102930 197033
rect 102874 196959 102930 196968
rect 102048 196648 102100 196654
rect 102048 196590 102100 196596
rect 101956 193928 102008 193934
rect 101956 193870 102008 193876
rect 101680 188420 101732 188426
rect 101680 188362 101732 188368
rect 101588 188284 101640 188290
rect 101588 188226 101640 188232
rect 101312 184476 101364 184482
rect 101312 184418 101364 184424
rect 101220 148980 101272 148986
rect 101220 148922 101272 148928
rect 100760 108996 100812 109002
rect 100760 108938 100812 108944
rect 100772 108322 100800 108938
rect 100760 108316 100812 108322
rect 100760 108258 100812 108264
rect 101232 81841 101260 148922
rect 101324 109002 101352 184418
rect 101772 180872 101824 180878
rect 101772 180814 101824 180820
rect 101680 178764 101732 178770
rect 101680 178706 101732 178712
rect 101496 174752 101548 174758
rect 101496 174694 101548 174700
rect 101404 148436 101456 148442
rect 101404 148378 101456 148384
rect 101312 108996 101364 109002
rect 101312 108938 101364 108944
rect 101218 81832 101274 81841
rect 101218 81767 101274 81776
rect 101416 65414 101444 148378
rect 101508 81025 101536 174694
rect 101588 174616 101640 174622
rect 101588 174558 101640 174564
rect 101494 81016 101550 81025
rect 101494 80951 101550 80960
rect 101600 77858 101628 174558
rect 101692 79830 101720 178706
rect 101680 79824 101732 79830
rect 101680 79766 101732 79772
rect 101784 78130 101812 180814
rect 101864 178968 101916 178974
rect 101864 178910 101916 178916
rect 101772 78124 101824 78130
rect 101772 78066 101824 78072
rect 101588 77852 101640 77858
rect 101588 77794 101640 77800
rect 101876 74526 101904 178910
rect 101864 74520 101916 74526
rect 101864 74462 101916 74468
rect 101404 65408 101456 65414
rect 101404 65350 101456 65356
rect 100668 64592 100720 64598
rect 100668 64534 100720 64540
rect 99932 64524 99984 64530
rect 99932 64466 99984 64472
rect 101968 63374 101996 193870
rect 102060 64841 102088 196590
rect 102980 195702 103008 476070
rect 103060 360256 103112 360262
rect 103060 360198 103112 360204
rect 102968 195696 103020 195702
rect 102968 195638 103020 195644
rect 103072 188494 103100 360198
rect 103152 335368 103204 335374
rect 103152 335310 103204 335316
rect 103060 188488 103112 188494
rect 103060 188430 103112 188436
rect 103164 185978 103192 335310
rect 103336 193860 103388 193866
rect 103336 193802 103388 193808
rect 103152 185972 103204 185978
rect 103152 185914 103204 185920
rect 103060 185700 103112 185706
rect 103060 185642 103112 185648
rect 102968 183932 103020 183938
rect 102968 183874 103020 183880
rect 102876 182232 102928 182238
rect 102876 182174 102928 182180
rect 102784 181008 102836 181014
rect 102784 180950 102836 180956
rect 102692 174684 102744 174690
rect 102692 174626 102744 174632
rect 102600 148912 102652 148918
rect 102600 148854 102652 148860
rect 102612 65618 102640 148854
rect 102704 74050 102732 174626
rect 102796 78198 102824 180950
rect 102888 79082 102916 182174
rect 102876 79076 102928 79082
rect 102876 79018 102928 79024
rect 102784 78192 102836 78198
rect 102784 78134 102836 78140
rect 102980 76838 103008 183874
rect 103072 77790 103100 185642
rect 103244 184136 103296 184142
rect 103244 184078 103296 184084
rect 103152 180940 103204 180946
rect 103152 180882 103204 180888
rect 103060 77784 103112 77790
rect 103060 77726 103112 77732
rect 102968 76832 103020 76838
rect 102968 76774 103020 76780
rect 102784 75880 102836 75886
rect 102784 75822 102836 75828
rect 102692 74044 102744 74050
rect 102692 73986 102744 73992
rect 102600 65612 102652 65618
rect 102600 65554 102652 65560
rect 102046 64832 102102 64841
rect 102046 64767 102102 64776
rect 102796 64258 102824 75822
rect 103164 68649 103192 180882
rect 103150 68640 103206 68649
rect 103150 68575 103206 68584
rect 103256 67114 103284 184078
rect 103348 67561 103376 193802
rect 103532 183462 103560 683086
rect 104164 680400 104216 680406
rect 104164 680342 104216 680348
rect 104072 299532 104124 299538
rect 104072 299474 104124 299480
rect 104084 191486 104112 299474
rect 104176 195809 104204 680342
rect 104256 621036 104308 621042
rect 104256 620978 104308 620984
rect 104162 195800 104218 195809
rect 104162 195735 104218 195744
rect 104268 194342 104296 620978
rect 104348 604512 104400 604518
rect 104348 604454 104400 604460
rect 104256 194336 104308 194342
rect 104256 194278 104308 194284
rect 104360 192545 104388 604454
rect 104900 596216 104952 596222
rect 104900 596158 104952 596164
rect 104440 484424 104492 484430
rect 104440 484366 104492 484372
rect 104452 195770 104480 484366
rect 104624 303680 104676 303686
rect 104624 303622 104676 303628
rect 104532 195832 104584 195838
rect 104532 195774 104584 195780
rect 104440 195764 104492 195770
rect 104440 195706 104492 195712
rect 104346 192536 104402 192545
rect 104346 192471 104402 192480
rect 104072 191480 104124 191486
rect 104072 191422 104124 191428
rect 104348 184612 104400 184618
rect 104348 184554 104400 184560
rect 103520 183456 103572 183462
rect 103520 183398 103572 183404
rect 104256 181892 104308 181898
rect 104256 181834 104308 181840
rect 103428 181688 103480 181694
rect 103428 181630 103480 181636
rect 103334 67552 103390 67561
rect 103334 67487 103390 67496
rect 103244 67108 103296 67114
rect 103244 67050 103296 67056
rect 102784 64252 102836 64258
rect 102784 64194 102836 64200
rect 102796 63578 102824 64194
rect 102140 63572 102192 63578
rect 102140 63514 102192 63520
rect 102784 63572 102836 63578
rect 102784 63514 102836 63520
rect 101956 63368 102008 63374
rect 101956 63310 102008 63316
rect 102152 16574 102180 63514
rect 103440 44130 103468 181630
rect 104164 178900 104216 178906
rect 104164 178842 104216 178848
rect 103980 148844 104032 148850
rect 103980 148786 104032 148792
rect 103992 84194 104020 148786
rect 104072 146940 104124 146946
rect 104072 146882 104124 146888
rect 104084 136610 104112 146882
rect 104072 136604 104124 136610
rect 104072 136546 104124 136552
rect 103900 84166 104020 84194
rect 103900 78062 103928 84166
rect 104084 81530 104112 136546
rect 104072 81524 104124 81530
rect 104072 81466 104124 81472
rect 104176 81410 104204 178842
rect 103992 81382 104204 81410
rect 103992 78470 104020 81382
rect 104072 81252 104124 81258
rect 104072 81194 104124 81200
rect 103980 78464 104032 78470
rect 103980 78406 104032 78412
rect 103888 78056 103940 78062
rect 103888 77998 103940 78004
rect 104084 65958 104112 81194
rect 104164 79348 104216 79354
rect 104164 79290 104216 79296
rect 104176 68814 104204 79290
rect 104164 68808 104216 68814
rect 104164 68750 104216 68756
rect 104268 66910 104296 181834
rect 104360 67318 104388 184554
rect 104440 184272 104492 184278
rect 104440 184214 104492 184220
rect 104452 67522 104480 184214
rect 104544 79218 104572 195774
rect 104636 193254 104664 303622
rect 104808 196852 104860 196858
rect 104808 196794 104860 196800
rect 104716 194064 104768 194070
rect 104716 194006 104768 194012
rect 104624 193248 104676 193254
rect 104624 193190 104676 193196
rect 104624 188488 104676 188494
rect 104624 188430 104676 188436
rect 104532 79212 104584 79218
rect 104532 79154 104584 79160
rect 104530 77208 104586 77217
rect 104530 77143 104586 77152
rect 104544 76566 104572 77143
rect 104532 76560 104584 76566
rect 104532 76502 104584 76508
rect 104440 67516 104492 67522
rect 104440 67458 104492 67464
rect 104348 67312 104400 67318
rect 104348 67254 104400 67260
rect 104636 67182 104664 188430
rect 104728 79354 104756 194006
rect 104716 79348 104768 79354
rect 104716 79290 104768 79296
rect 104716 79212 104768 79218
rect 104716 79154 104768 79160
rect 104728 75857 104756 79154
rect 104714 75848 104770 75857
rect 104714 75783 104770 75792
rect 104820 67289 104848 196794
rect 104912 188562 104940 596158
rect 105544 456816 105596 456822
rect 105544 456758 105596 456764
rect 104992 408536 105044 408542
rect 104992 408478 105044 408484
rect 104900 188556 104952 188562
rect 104900 188498 104952 188504
rect 105004 183258 105032 408478
rect 105556 195265 105584 456758
rect 106004 198892 106056 198898
rect 106004 198834 106056 198840
rect 105542 195256 105598 195265
rect 105542 195191 105598 195200
rect 105912 191208 105964 191214
rect 105912 191150 105964 191156
rect 104992 183252 105044 183258
rect 104992 183194 105044 183200
rect 105820 183252 105872 183258
rect 105820 183194 105872 183200
rect 105832 182238 105860 183194
rect 105820 182232 105872 182238
rect 105820 182174 105872 182180
rect 105636 181620 105688 181626
rect 105636 181562 105688 181568
rect 105544 177336 105596 177342
rect 105544 177278 105596 177284
rect 105360 144288 105412 144294
rect 105360 144230 105412 144236
rect 105372 132462 105400 144230
rect 105450 135960 105506 135969
rect 105450 135895 105506 135904
rect 105360 132456 105412 132462
rect 105360 132398 105412 132404
rect 105360 99408 105412 99414
rect 105360 99350 105412 99356
rect 105372 68134 105400 99350
rect 105360 68128 105412 68134
rect 105360 68070 105412 68076
rect 104806 67280 104862 67289
rect 104716 67244 104768 67250
rect 104806 67215 104862 67224
rect 104716 67186 104768 67192
rect 104624 67176 104676 67182
rect 104624 67118 104676 67124
rect 104728 66910 104756 67186
rect 104256 66904 104308 66910
rect 104256 66846 104308 66852
rect 104716 66904 104768 66910
rect 104716 66846 104768 66852
rect 104072 65952 104124 65958
rect 104072 65894 104124 65900
rect 105464 65890 105492 135895
rect 105556 80889 105584 177278
rect 105542 80880 105598 80889
rect 105542 80815 105598 80824
rect 105648 79529 105676 181562
rect 105728 179444 105780 179450
rect 105728 179386 105780 179392
rect 105634 79520 105690 79529
rect 105634 79455 105690 79464
rect 105740 77926 105768 179386
rect 105820 177404 105872 177410
rect 105820 177346 105872 177352
rect 105728 77920 105780 77926
rect 105728 77862 105780 77868
rect 105832 71097 105860 177346
rect 105924 78538 105952 191150
rect 106016 79762 106044 198834
rect 106188 188964 106240 188970
rect 106188 188906 106240 188912
rect 106200 188562 106228 188906
rect 106292 188630 106320 703582
rect 106752 703474 106780 703582
rect 106894 703520 107006 704960
rect 110432 703582 110644 703610
rect 106936 703474 106964 703520
rect 106752 703446 106964 703474
rect 109040 700460 109092 700466
rect 109040 700402 109092 700408
rect 108304 652792 108356 652798
rect 108304 652734 108356 652740
rect 106924 560312 106976 560318
rect 106924 560254 106976 560260
rect 106936 196897 106964 560254
rect 107016 379568 107068 379574
rect 107016 379510 107068 379516
rect 106922 196888 106978 196897
rect 106922 196823 106978 196832
rect 107028 196450 107056 379510
rect 107108 343664 107160 343670
rect 107108 343606 107160 343612
rect 107016 196444 107068 196450
rect 107016 196386 107068 196392
rect 107120 194478 107148 343606
rect 107200 307828 107252 307834
rect 107200 307770 107252 307776
rect 107108 194472 107160 194478
rect 107108 194414 107160 194420
rect 107212 194274 107240 307770
rect 107292 263628 107344 263634
rect 107292 263570 107344 263576
rect 107200 194268 107252 194274
rect 107200 194210 107252 194216
rect 107016 194132 107068 194138
rect 107016 194074 107068 194080
rect 106280 188624 106332 188630
rect 106280 188566 106332 188572
rect 106188 188556 106240 188562
rect 106188 188498 106240 188504
rect 106096 186856 106148 186862
rect 106096 186798 106148 186804
rect 106004 79756 106056 79762
rect 106004 79698 106056 79704
rect 105912 78532 105964 78538
rect 105912 78474 105964 78480
rect 105818 71088 105874 71097
rect 105818 71023 105874 71032
rect 105452 65884 105504 65890
rect 105452 65826 105504 65832
rect 106108 64870 106136 186798
rect 106188 184408 106240 184414
rect 106188 184350 106240 184356
rect 106096 64864 106148 64870
rect 106096 64806 106148 64812
rect 106108 64190 106136 64806
rect 106096 64184 106148 64190
rect 106096 64126 106148 64132
rect 106200 57934 106228 184350
rect 106924 174548 106976 174554
rect 106924 174490 106976 174496
rect 106832 149048 106884 149054
rect 106832 148990 106884 148996
rect 106740 148300 106792 148306
rect 106740 148242 106792 148248
rect 106280 74520 106332 74526
rect 106280 74462 106332 74468
rect 106292 73574 106320 74462
rect 106280 73568 106332 73574
rect 106280 73510 106332 73516
rect 105636 57928 105688 57934
rect 105636 57870 105688 57876
rect 106188 57928 106240 57934
rect 106188 57870 106240 57876
rect 105648 57254 105676 57870
rect 105636 57248 105688 57254
rect 105636 57190 105688 57196
rect 103428 44124 103480 44130
rect 103428 44066 103480 44072
rect 98012 16546 98592 16574
rect 102152 16546 102456 16574
rect 97908 3528 97960 3534
rect 97908 3470 97960 3476
rect 98564 480 98592 16546
rect 102428 480 102456 16546
rect 106292 480 106320 73510
rect 106752 71262 106780 148242
rect 106740 71256 106792 71262
rect 106740 71198 106792 71204
rect 106844 70854 106872 148990
rect 106832 70848 106884 70854
rect 106832 70790 106884 70796
rect 106936 70281 106964 174490
rect 107028 77110 107056 194074
rect 107108 186380 107160 186386
rect 107108 186322 107160 186328
rect 107016 77104 107068 77110
rect 107016 77046 107068 77052
rect 107016 74792 107068 74798
rect 107016 74734 107068 74740
rect 106922 70272 106978 70281
rect 106922 70207 106978 70216
rect 107028 68270 107056 74734
rect 107120 69465 107148 186322
rect 107200 185564 107252 185570
rect 107200 185506 107252 185512
rect 107106 69456 107162 69465
rect 107106 69391 107162 69400
rect 107212 69018 107240 185506
rect 107304 183326 107332 263570
rect 107566 200696 107622 200705
rect 107566 200631 107622 200640
rect 107580 200297 107608 200631
rect 107566 200288 107622 200297
rect 107566 200223 107622 200232
rect 107476 194404 107528 194410
rect 107476 194346 107528 194352
rect 107384 185904 107436 185910
rect 107384 185846 107436 185852
rect 107396 185570 107424 185846
rect 107384 185564 107436 185570
rect 107384 185506 107436 185512
rect 107384 184068 107436 184074
rect 107384 184010 107436 184016
rect 107292 183320 107344 183326
rect 107292 183262 107344 183268
rect 107292 181960 107344 181966
rect 107292 181902 107344 181908
rect 107200 69012 107252 69018
rect 107200 68954 107252 68960
rect 107016 68264 107068 68270
rect 107016 68206 107068 68212
rect 107304 64394 107332 181902
rect 107292 64388 107344 64394
rect 107292 64330 107344 64336
rect 107396 64326 107424 184010
rect 107488 74798 107516 194346
rect 107476 74792 107528 74798
rect 107476 74734 107528 74740
rect 107476 74656 107528 74662
rect 107476 74598 107528 74604
rect 107488 73574 107516 74598
rect 107476 73568 107528 73574
rect 107476 73510 107528 73516
rect 107580 65754 107608 200223
rect 108120 199640 108172 199646
rect 108120 199582 108172 199588
rect 108132 199034 108160 199582
rect 108212 199572 108264 199578
rect 108212 199514 108264 199520
rect 108120 199028 108172 199034
rect 108120 198970 108172 198976
rect 108224 198966 108252 199514
rect 108212 198960 108264 198966
rect 108212 198902 108264 198908
rect 108028 189100 108080 189106
rect 108028 189042 108080 189048
rect 107660 75268 107712 75274
rect 107660 75210 107712 75216
rect 107672 74662 107700 75210
rect 107660 74656 107712 74662
rect 107660 74598 107712 74604
rect 108040 69630 108068 189042
rect 108316 186726 108344 652734
rect 108396 512032 108448 512038
rect 108396 511974 108448 511980
rect 108408 194954 108436 511974
rect 108488 496868 108540 496874
rect 108488 496810 108540 496816
rect 108396 194948 108448 194954
rect 108396 194890 108448 194896
rect 108500 188562 108528 496810
rect 108580 427848 108632 427854
rect 108580 427790 108632 427796
rect 108592 197266 108620 427790
rect 108672 287088 108724 287094
rect 108672 287030 108724 287036
rect 108580 197260 108632 197266
rect 108580 197202 108632 197208
rect 108684 194206 108712 287030
rect 108764 199436 108816 199442
rect 108764 199378 108816 199384
rect 108672 194200 108724 194206
rect 108672 194142 108724 194148
rect 108672 191480 108724 191486
rect 108672 191422 108724 191428
rect 108684 191350 108712 191422
rect 108672 191344 108724 191350
rect 108672 191286 108724 191292
rect 108488 188556 108540 188562
rect 108488 188498 108540 188504
rect 108304 186720 108356 186726
rect 108304 186662 108356 186668
rect 108580 184544 108632 184550
rect 108580 184486 108632 184492
rect 108304 183320 108356 183326
rect 108304 183262 108356 183268
rect 108316 182850 108344 183262
rect 108304 182844 108356 182850
rect 108304 182786 108356 182792
rect 108120 140820 108172 140826
rect 108120 140762 108172 140768
rect 108132 88330 108160 140762
rect 108212 137284 108264 137290
rect 108212 137226 108264 137232
rect 108120 88324 108172 88330
rect 108120 88266 108172 88272
rect 108224 79422 108252 137226
rect 108212 79416 108264 79422
rect 108212 79358 108264 79364
rect 108316 78266 108344 182786
rect 108396 182028 108448 182034
rect 108396 181970 108448 181976
rect 108304 78260 108356 78266
rect 108304 78202 108356 78208
rect 108028 69624 108080 69630
rect 108028 69566 108080 69572
rect 107568 65748 107620 65754
rect 107568 65690 107620 65696
rect 108408 64462 108436 181970
rect 108396 64456 108448 64462
rect 108396 64398 108448 64404
rect 107384 64320 107436 64326
rect 107384 64262 107436 64268
rect 108592 64190 108620 184486
rect 108684 69902 108712 191286
rect 108776 74186 108804 199378
rect 108948 199028 109000 199034
rect 108948 198970 109000 198976
rect 108856 198960 108908 198966
rect 108856 198902 108908 198908
rect 108764 74180 108816 74186
rect 108764 74122 108816 74128
rect 108868 71330 108896 198902
rect 108856 71324 108908 71330
rect 108856 71266 108908 71272
rect 108960 70378 108988 198970
rect 109052 197305 109080 700402
rect 109132 444440 109184 444446
rect 109132 444382 109184 444388
rect 109144 197470 109172 444382
rect 109224 273964 109276 273970
rect 109224 273906 109276 273912
rect 109236 273290 109264 273906
rect 109224 273284 109276 273290
rect 109224 273226 109276 273232
rect 110236 273284 110288 273290
rect 110236 273226 110288 273232
rect 109684 236020 109736 236026
rect 109684 235962 109736 235968
rect 109132 197464 109184 197470
rect 109132 197406 109184 197412
rect 109038 197296 109094 197305
rect 109038 197231 109094 197240
rect 109052 196722 109080 197231
rect 109144 197130 109172 197406
rect 109132 197124 109184 197130
rect 109132 197066 109184 197072
rect 109040 196716 109092 196722
rect 109040 196658 109092 196664
rect 109696 190058 109724 235962
rect 109868 195900 109920 195906
rect 109868 195842 109920 195848
rect 109684 190052 109736 190058
rect 109684 189994 109736 190000
rect 109500 189848 109552 189854
rect 109500 189790 109552 189796
rect 109512 76702 109540 189790
rect 109776 187740 109828 187746
rect 109776 187682 109828 187688
rect 109684 184340 109736 184346
rect 109684 184282 109736 184288
rect 109592 178696 109644 178702
rect 109592 178638 109644 178644
rect 109500 76696 109552 76702
rect 109500 76638 109552 76644
rect 108948 70372 109000 70378
rect 108948 70314 109000 70320
rect 108672 69896 108724 69902
rect 108672 69838 108724 69844
rect 108580 64184 108632 64190
rect 108580 64126 108632 64132
rect 109604 63170 109632 178638
rect 109696 67590 109724 184282
rect 109788 70242 109816 187682
rect 109880 75449 109908 195842
rect 110144 187400 110196 187406
rect 110144 187342 110196 187348
rect 110052 187332 110104 187338
rect 110052 187274 110104 187280
rect 109960 187128 110012 187134
rect 109960 187070 110012 187076
rect 109866 75440 109922 75449
rect 109866 75375 109922 75384
rect 109776 70236 109828 70242
rect 109776 70178 109828 70184
rect 109684 67584 109736 67590
rect 109684 67526 109736 67532
rect 109972 67454 110000 187070
rect 109960 67448 110012 67454
rect 109960 67390 110012 67396
rect 110064 66706 110092 187274
rect 110052 66700 110104 66706
rect 110052 66642 110104 66648
rect 110156 65550 110184 187342
rect 110248 145897 110276 273226
rect 110328 199776 110380 199782
rect 110328 199718 110380 199724
rect 110234 145888 110290 145897
rect 110234 145823 110290 145832
rect 110236 144628 110288 144634
rect 110236 144570 110288 144576
rect 110248 79354 110276 144570
rect 110236 79348 110288 79354
rect 110236 79290 110288 79296
rect 110340 68882 110368 199718
rect 110432 190233 110460 703582
rect 110616 703474 110644 703582
rect 110758 703520 110870 704960
rect 114622 703520 114734 704960
rect 117332 703582 118372 703610
rect 110800 703474 110828 703520
rect 110616 703446 110828 703474
rect 114664 702434 114692 703520
rect 114572 702406 114692 702434
rect 114572 699802 114600 702406
rect 117228 700460 117280 700466
rect 117228 700402 117280 700408
rect 115848 700392 115900 700398
rect 115848 700334 115900 700340
rect 114480 699774 114600 699802
rect 112444 663808 112496 663814
rect 112444 663750 112496 663756
rect 110512 543788 110564 543794
rect 110512 543730 110564 543736
rect 110524 194002 110552 543730
rect 111064 488572 111116 488578
rect 111064 488514 111116 488520
rect 111076 197198 111104 488514
rect 111616 263152 111668 263158
rect 111616 263094 111668 263100
rect 111248 260160 111300 260166
rect 111248 260102 111300 260108
rect 111156 259752 111208 259758
rect 111156 259694 111208 259700
rect 111064 197192 111116 197198
rect 111064 197134 111116 197140
rect 110512 193996 110564 194002
rect 110512 193938 110564 193944
rect 110418 190224 110474 190233
rect 110418 190159 110474 190168
rect 110972 189984 111024 189990
rect 110972 189926 111024 189932
rect 110880 189916 110932 189922
rect 110880 189858 110932 189864
rect 110420 184000 110472 184006
rect 110420 183942 110472 183948
rect 110432 183326 110460 183942
rect 110420 183320 110472 183326
rect 110420 183262 110472 183268
rect 110420 143064 110472 143070
rect 110420 143006 110472 143012
rect 110432 142866 110460 143006
rect 110420 142860 110472 142866
rect 110420 142802 110472 142808
rect 110420 104848 110472 104854
rect 110420 104790 110472 104796
rect 110432 104174 110460 104790
rect 110420 104168 110472 104174
rect 110420 104110 110472 104116
rect 110328 68876 110380 68882
rect 110328 68818 110380 68824
rect 110892 67386 110920 189858
rect 110984 104854 111012 189926
rect 111064 183320 111116 183326
rect 111064 183262 111116 183268
rect 110972 104848 111024 104854
rect 110972 104790 111024 104796
rect 110972 93152 111024 93158
rect 110972 93094 111024 93100
rect 110984 71194 111012 93094
rect 111076 71534 111104 183262
rect 111168 146062 111196 259694
rect 111156 146056 111208 146062
rect 111156 145998 111208 146004
rect 111260 145994 111288 260102
rect 111340 193044 111392 193050
rect 111340 192986 111392 192992
rect 111248 145988 111300 145994
rect 111248 145930 111300 145936
rect 111248 139324 111300 139330
rect 111248 139266 111300 139272
rect 111156 108316 111208 108322
rect 111156 108258 111208 108264
rect 111168 79490 111196 108258
rect 111156 79484 111208 79490
rect 111156 79426 111208 79432
rect 111064 71528 111116 71534
rect 111064 71470 111116 71476
rect 110972 71188 111024 71194
rect 110972 71130 111024 71136
rect 111260 68950 111288 139266
rect 111352 73982 111380 192986
rect 111524 188420 111576 188426
rect 111524 188362 111576 188368
rect 111432 147008 111484 147014
rect 111432 146950 111484 146956
rect 111340 73976 111392 73982
rect 111340 73918 111392 73924
rect 111248 68944 111300 68950
rect 111248 68886 111300 68892
rect 110880 67380 110932 67386
rect 110880 67322 110932 67328
rect 110144 65544 110196 65550
rect 110144 65486 110196 65492
rect 111444 65482 111472 146950
rect 111536 68474 111564 188362
rect 111628 143070 111656 263094
rect 112352 259820 112404 259826
rect 112352 259762 112404 259768
rect 111798 200968 111854 200977
rect 111798 200903 111854 200912
rect 111812 200433 111840 200903
rect 111798 200424 111854 200433
rect 111798 200359 111854 200368
rect 111708 195220 111760 195226
rect 111708 195162 111760 195168
rect 111616 143064 111668 143070
rect 111616 143006 111668 143012
rect 111616 95940 111668 95946
rect 111616 95882 111668 95888
rect 111628 82142 111656 95882
rect 111616 82136 111668 82142
rect 111616 82078 111668 82084
rect 111720 72690 111748 195162
rect 111800 193996 111852 194002
rect 111800 193938 111852 193944
rect 111812 193118 111840 193938
rect 111800 193112 111852 193118
rect 111800 193054 111852 193060
rect 112260 191140 112312 191146
rect 112260 191082 112312 191088
rect 112272 180810 112300 191082
rect 112260 180804 112312 180810
rect 112260 180746 112312 180752
rect 112364 146198 112392 259762
rect 112456 189961 112484 663750
rect 113824 460964 113876 460970
rect 113824 460906 113876 460912
rect 112536 416832 112588 416838
rect 112536 416774 112588 416780
rect 112548 264994 112576 416774
rect 112536 264988 112588 264994
rect 112536 264930 112588 264936
rect 112720 263968 112772 263974
rect 112720 263910 112772 263916
rect 112536 263084 112588 263090
rect 112536 263026 112588 263032
rect 112442 189952 112498 189961
rect 112442 189887 112498 189896
rect 112444 187196 112496 187202
rect 112444 187138 112496 187144
rect 112352 146192 112404 146198
rect 112352 146134 112404 146140
rect 112260 145580 112312 145586
rect 112260 145522 112312 145528
rect 112168 145512 112220 145518
rect 112168 145454 112220 145460
rect 111708 72684 111760 72690
rect 111708 72626 111760 72632
rect 112180 68746 112208 145454
rect 112272 94790 112300 145522
rect 112352 140480 112404 140486
rect 112352 140422 112404 140428
rect 112260 94784 112312 94790
rect 112260 94726 112312 94732
rect 112364 79014 112392 140422
rect 112352 79008 112404 79014
rect 112352 78950 112404 78956
rect 112456 72593 112484 187138
rect 112548 146033 112576 263026
rect 112628 259888 112680 259894
rect 112628 259830 112680 259836
rect 112534 146024 112590 146033
rect 112534 145959 112590 145968
rect 112640 143478 112668 259830
rect 112732 145926 112760 263910
rect 112904 262608 112956 262614
rect 112904 262550 112956 262556
rect 112810 262440 112866 262449
rect 112810 262375 112866 262384
rect 112720 145920 112772 145926
rect 112720 145862 112772 145868
rect 112720 145648 112772 145654
rect 112720 145590 112772 145596
rect 112628 143472 112680 143478
rect 112628 143414 112680 143420
rect 112536 140276 112588 140282
rect 112536 140218 112588 140224
rect 112548 74118 112576 140218
rect 112628 140208 112680 140214
rect 112628 140150 112680 140156
rect 112536 74112 112588 74118
rect 112536 74054 112588 74060
rect 112640 73778 112668 140150
rect 112628 73772 112680 73778
rect 112628 73714 112680 73720
rect 112442 72584 112498 72593
rect 112442 72519 112498 72528
rect 112732 72457 112760 145590
rect 112824 144770 112852 262375
rect 112916 144838 112944 262550
rect 113640 259684 113692 259690
rect 113640 259626 113692 259632
rect 112996 231872 113048 231878
rect 112996 231814 113048 231820
rect 113008 191486 113036 231814
rect 113086 200424 113142 200433
rect 113086 200359 113142 200368
rect 112996 191480 113048 191486
rect 112996 191422 113048 191428
rect 112994 189952 113050 189961
rect 112994 189887 113050 189896
rect 112904 144832 112956 144838
rect 112904 144774 112956 144780
rect 112812 144764 112864 144770
rect 112812 144706 112864 144712
rect 112904 141908 112956 141914
rect 112904 141850 112956 141856
rect 112718 72448 112774 72457
rect 112718 72383 112774 72392
rect 112168 68740 112220 68746
rect 112168 68682 112220 68688
rect 111524 68468 111576 68474
rect 111524 68410 111576 68416
rect 111432 65476 111484 65482
rect 111432 65418 111484 65424
rect 112916 64802 112944 141850
rect 113008 71233 113036 189887
rect 113100 79218 113128 200359
rect 113652 142225 113680 259626
rect 113836 200802 113864 460906
rect 113916 339516 113968 339522
rect 113916 339458 113968 339464
rect 113928 263634 113956 339458
rect 113916 263628 113968 263634
rect 113916 263570 113968 263576
rect 113916 263220 113968 263226
rect 113916 263162 113968 263168
rect 113824 200796 113876 200802
rect 113824 200738 113876 200744
rect 113732 187060 113784 187066
rect 113732 187002 113784 187008
rect 113638 142216 113694 142225
rect 113272 142180 113324 142186
rect 113638 142151 113694 142160
rect 113272 142122 113324 142128
rect 113284 141846 113312 142122
rect 113272 141840 113324 141846
rect 113272 141782 113324 141788
rect 113652 141438 113680 142151
rect 113640 141432 113692 141438
rect 113640 141374 113692 141380
rect 113180 140888 113232 140894
rect 113180 140830 113232 140836
rect 113088 79212 113140 79218
rect 113088 79154 113140 79160
rect 112994 71224 113050 71233
rect 112994 71159 113050 71168
rect 112904 64796 112956 64802
rect 112904 64738 112956 64744
rect 109592 63164 109644 63170
rect 109592 63106 109644 63112
rect 110144 6248 110196 6254
rect 110144 6190 110196 6196
rect 110156 480 110184 6190
rect 72118 354 72230 480
rect 71792 326 72230 354
rect 64390 -960 64502 326
rect 68254 -960 68366 326
rect 72118 -960 72230 326
rect 75338 -960 75450 480
rect 79202 -960 79314 480
rect 83066 -960 83178 480
rect 86930 -960 87042 480
rect 90794 -960 90906 480
rect 94658 -960 94770 480
rect 98522 -960 98634 480
rect 102386 -960 102498 480
rect 106250 -960 106362 480
rect 110114 -960 110226 480
rect 113192 354 113220 140830
rect 113744 81122 113772 187002
rect 113824 181824 113876 181830
rect 113824 181766 113876 181772
rect 113732 81116 113784 81122
rect 113732 81058 113784 81064
rect 113836 69834 113864 181766
rect 113928 141846 113956 263162
rect 114284 262744 114336 262750
rect 114284 262686 114336 262692
rect 114100 262472 114152 262478
rect 114100 262414 114152 262420
rect 114008 260228 114060 260234
rect 114008 260170 114060 260176
rect 114020 145858 114048 260170
rect 114112 147626 114140 262414
rect 114100 147620 114152 147626
rect 114100 147562 114152 147568
rect 114296 146130 114324 262686
rect 114376 260976 114428 260982
rect 114376 260918 114428 260924
rect 114388 220794 114416 260918
rect 114376 220788 114428 220794
rect 114376 220730 114428 220736
rect 114480 198150 114508 699774
rect 115204 520328 115256 520334
rect 115204 520270 115256 520276
rect 115020 264104 115072 264110
rect 115020 264046 115072 264052
rect 114468 198144 114520 198150
rect 114468 198086 114520 198092
rect 114836 194540 114888 194546
rect 114836 194482 114888 194488
rect 114468 194472 114520 194478
rect 114468 194414 114520 194420
rect 114480 192982 114508 194414
rect 114468 192976 114520 192982
rect 114468 192918 114520 192924
rect 114480 192658 114508 192918
rect 114388 192630 114508 192658
rect 114284 146124 114336 146130
rect 114284 146066 114336 146072
rect 114008 145852 114060 145858
rect 114008 145794 114060 145800
rect 114192 145784 114244 145790
rect 114192 145726 114244 145732
rect 114100 145376 114152 145382
rect 114100 145318 114152 145324
rect 113916 141840 113968 141846
rect 113916 141782 113968 141788
rect 114008 140140 114060 140146
rect 114008 140082 114060 140088
rect 113916 139936 113968 139942
rect 113916 139878 113968 139884
rect 113928 79150 113956 139878
rect 113916 79144 113968 79150
rect 113916 79086 113968 79092
rect 114020 74390 114048 140082
rect 114008 74384 114060 74390
rect 114008 74326 114060 74332
rect 114112 72826 114140 145318
rect 114100 72820 114152 72826
rect 114100 72762 114152 72768
rect 114204 70922 114232 145726
rect 114284 144492 114336 144498
rect 114284 144434 114336 144440
rect 114192 70916 114244 70922
rect 114192 70858 114244 70864
rect 113824 69828 113876 69834
rect 113824 69770 113876 69776
rect 114296 68610 114324 144434
rect 114388 75682 114416 192630
rect 114468 192568 114520 192574
rect 114468 192510 114520 192516
rect 114376 75676 114428 75682
rect 114376 75618 114428 75624
rect 114480 75410 114508 192510
rect 114468 75404 114520 75410
rect 114468 75346 114520 75352
rect 114848 73030 114876 194482
rect 114928 148776 114980 148782
rect 114928 148718 114980 148724
rect 114836 73024 114888 73030
rect 114836 72966 114888 72972
rect 114940 72758 114968 148718
rect 115032 142769 115060 264046
rect 115112 259616 115164 259622
rect 115112 259558 115164 259564
rect 115124 143313 115152 259558
rect 115216 200734 115244 520270
rect 115388 267028 115440 267034
rect 115388 266970 115440 266976
rect 115400 262857 115428 266970
rect 115756 264988 115808 264994
rect 115756 264930 115808 264936
rect 115572 264036 115624 264042
rect 115572 263978 115624 263984
rect 115584 263634 115612 263978
rect 115572 263628 115624 263634
rect 115572 263570 115624 263576
rect 115386 262848 115442 262857
rect 115386 262783 115442 262792
rect 115296 262404 115348 262410
rect 115296 262346 115348 262352
rect 115204 200728 115256 200734
rect 115204 200670 115256 200676
rect 115308 143546 115336 262346
rect 115296 143540 115348 143546
rect 115296 143482 115348 143488
rect 115110 143304 115166 143313
rect 115110 143239 115166 143248
rect 115308 143002 115336 143482
rect 115400 143410 115428 262783
rect 115480 186924 115532 186930
rect 115480 186866 115532 186872
rect 115388 143404 115440 143410
rect 115388 143346 115440 143352
rect 115296 142996 115348 143002
rect 115296 142938 115348 142944
rect 115112 142860 115164 142866
rect 115112 142802 115164 142808
rect 115018 142760 115074 142769
rect 115018 142695 115074 142704
rect 115020 94784 115072 94790
rect 115020 94726 115072 94732
rect 114928 72752 114980 72758
rect 114928 72694 114980 72700
rect 114284 68604 114336 68610
rect 114284 68546 114336 68552
rect 115032 63306 115060 94726
rect 115124 80646 115152 142802
rect 115204 140684 115256 140690
rect 115204 140626 115256 140632
rect 115112 80640 115164 80646
rect 115112 80582 115164 80588
rect 115216 73710 115244 140626
rect 115388 140548 115440 140554
rect 115388 140490 115440 140496
rect 115296 140412 115348 140418
rect 115296 140354 115348 140360
rect 115308 73846 115336 140354
rect 115296 73840 115348 73846
rect 115296 73782 115348 73788
rect 115204 73704 115256 73710
rect 115204 73646 115256 73652
rect 115400 72554 115428 140490
rect 115388 72548 115440 72554
rect 115388 72490 115440 72496
rect 115492 67017 115520 186866
rect 115584 143342 115612 263570
rect 115664 144560 115716 144566
rect 115664 144502 115716 144508
rect 115572 143336 115624 143342
rect 115572 143278 115624 143284
rect 115572 141636 115624 141642
rect 115572 141578 115624 141584
rect 115584 70174 115612 141578
rect 115676 71466 115704 144502
rect 115768 143002 115796 264930
rect 115860 191282 115888 700334
rect 115940 600364 115992 600370
rect 115940 600306 115992 600312
rect 115952 202842 115980 600306
rect 117136 263832 117188 263838
rect 117136 263774 117188 263780
rect 117044 262812 117096 262818
rect 117044 262754 117096 262760
rect 116952 262676 117004 262682
rect 116952 262618 117004 262624
rect 116860 262268 116912 262274
rect 116860 262210 116912 262216
rect 116676 260092 116728 260098
rect 116676 260034 116728 260040
rect 115940 202836 115992 202842
rect 115940 202778 115992 202784
rect 116584 202836 116636 202842
rect 116584 202778 116636 202784
rect 116596 201618 116624 202778
rect 116584 201612 116636 201618
rect 116584 201554 116636 201560
rect 116596 199209 116624 201554
rect 116582 199200 116638 199209
rect 116582 199135 116638 199144
rect 116308 193792 116360 193798
rect 116308 193734 116360 193740
rect 115848 191276 115900 191282
rect 115848 191218 115900 191224
rect 116216 144084 116268 144090
rect 116216 144026 116268 144032
rect 115756 142996 115808 143002
rect 115756 142938 115808 142944
rect 115664 71460 115716 71466
rect 115664 71402 115716 71408
rect 115572 70168 115624 70174
rect 115572 70110 115624 70116
rect 116228 68542 116256 144026
rect 116320 75546 116348 193734
rect 116584 190596 116636 190602
rect 116584 190538 116636 190544
rect 116596 172514 116624 190538
rect 116584 172508 116636 172514
rect 116584 172450 116636 172456
rect 116688 145450 116716 260034
rect 116768 259344 116820 259350
rect 116768 259286 116820 259292
rect 116780 145722 116808 259286
rect 116768 145716 116820 145722
rect 116768 145658 116820 145664
rect 116676 145444 116728 145450
rect 116676 145386 116728 145392
rect 116492 144696 116544 144702
rect 116492 144638 116544 144644
rect 116504 110634 116532 144638
rect 116676 144152 116728 144158
rect 116676 144094 116728 144100
rect 116584 141976 116636 141982
rect 116584 141918 116636 141924
rect 116492 110628 116544 110634
rect 116492 110570 116544 110576
rect 116400 95260 116452 95266
rect 116400 95202 116452 95208
rect 116412 77246 116440 95202
rect 116596 80918 116624 141918
rect 116688 81705 116716 144094
rect 116872 143138 116900 262210
rect 116964 143206 116992 262618
rect 117056 147082 117084 262754
rect 117044 147076 117096 147082
rect 117044 147018 117096 147024
rect 117148 146826 117176 263774
rect 117240 190330 117268 700402
rect 117332 193225 117360 703582
rect 118344 703474 118372 703582
rect 118486 703520 118598 704960
rect 122350 703520 122462 704960
rect 126214 703520 126326 704960
rect 130078 703520 130190 704960
rect 133942 703520 134054 704960
rect 137806 703520 137918 704960
rect 141670 703520 141782 704960
rect 144890 703520 145002 704960
rect 148754 703520 148866 704960
rect 152618 703520 152730 704960
rect 156482 703520 156594 704960
rect 160346 703520 160458 704960
rect 164210 703520 164322 704960
rect 168074 703520 168186 704960
rect 171938 703520 172050 704960
rect 175802 703520 175914 704960
rect 179022 703520 179134 704960
rect 182192 703582 182772 703610
rect 118528 703474 118556 703520
rect 118344 703446 118556 703474
rect 131120 701072 131172 701078
rect 131120 701014 131172 701020
rect 122840 700664 122892 700670
rect 122840 700606 122892 700612
rect 117964 700528 118016 700534
rect 117964 700470 118016 700476
rect 117688 263900 117740 263906
rect 117688 263842 117740 263848
rect 117412 255332 117464 255338
rect 117412 255274 117464 255280
rect 117424 201550 117452 255274
rect 117412 201544 117464 201550
rect 117412 201486 117464 201492
rect 117318 193216 117374 193225
rect 117318 193151 117374 193160
rect 117228 190324 117280 190330
rect 117228 190266 117280 190272
rect 117228 147076 117280 147082
rect 117228 147018 117280 147024
rect 117056 146798 117176 146826
rect 116952 143200 117004 143206
rect 116952 143142 117004 143148
rect 117056 143138 117084 146798
rect 117136 144220 117188 144226
rect 117136 144162 117188 144168
rect 116860 143132 116912 143138
rect 116860 143074 116912 143080
rect 117044 143132 117096 143138
rect 117044 143074 117096 143080
rect 116872 142798 116900 143074
rect 116860 142792 116912 142798
rect 116860 142734 116912 142740
rect 117044 141772 117096 141778
rect 117044 141714 117096 141720
rect 116860 140004 116912 140010
rect 116860 139946 116912 139952
rect 116766 138680 116822 138689
rect 116766 138615 116822 138624
rect 116674 81696 116730 81705
rect 116674 81631 116730 81640
rect 116584 80912 116636 80918
rect 116584 80854 116636 80860
rect 116400 77240 116452 77246
rect 116400 77182 116452 77188
rect 116780 75614 116808 138615
rect 116768 75608 116820 75614
rect 116768 75550 116820 75556
rect 116308 75540 116360 75546
rect 116308 75482 116360 75488
rect 116872 71670 116900 139946
rect 116952 111852 117004 111858
rect 116952 111794 117004 111800
rect 116964 77042 116992 111794
rect 116952 77036 117004 77042
rect 116952 76978 117004 76984
rect 116860 71664 116912 71670
rect 116860 71606 116912 71612
rect 117056 71398 117084 141714
rect 117148 132494 117176 144162
rect 117240 142118 117268 147018
rect 117700 143041 117728 263842
rect 117872 260024 117924 260030
rect 117872 259966 117924 259972
rect 117780 201544 117832 201550
rect 117780 201486 117832 201492
rect 117792 200705 117820 201486
rect 117778 200696 117834 200705
rect 117778 200631 117834 200640
rect 117780 196716 117832 196722
rect 117780 196658 117832 196664
rect 117792 155922 117820 196658
rect 117780 155916 117832 155922
rect 117780 155858 117832 155864
rect 117884 146266 117912 259966
rect 117976 199850 118004 700470
rect 120724 700324 120776 700330
rect 120724 700266 120776 700272
rect 120080 605872 120132 605878
rect 120080 605814 120132 605820
rect 119988 456816 120040 456822
rect 119988 456758 120040 456764
rect 119344 440292 119396 440298
rect 119344 440234 119396 440240
rect 118056 412684 118108 412690
rect 118056 412626 118108 412632
rect 117964 199844 118016 199850
rect 117964 199786 118016 199792
rect 117976 198762 118004 199786
rect 118068 199578 118096 412626
rect 118700 264240 118752 264246
rect 118700 264182 118752 264188
rect 118712 263702 118740 264182
rect 118700 263696 118752 263702
rect 118700 263638 118752 263644
rect 119068 263696 119120 263702
rect 119068 263638 119120 263644
rect 118608 260840 118660 260846
rect 118608 260782 118660 260788
rect 118332 259548 118384 259554
rect 118332 259490 118384 259496
rect 118056 199572 118108 199578
rect 118056 199514 118108 199520
rect 117964 198756 118016 198762
rect 117964 198698 118016 198704
rect 117964 196784 118016 196790
rect 117964 196726 118016 196732
rect 117872 146260 117924 146266
rect 117872 146202 117924 146208
rect 117686 143032 117742 143041
rect 117686 142967 117742 142976
rect 117228 142112 117280 142118
rect 117228 142054 117280 142060
rect 117240 140894 117268 142054
rect 117686 141944 117742 141953
rect 117686 141879 117742 141888
rect 117228 140888 117280 140894
rect 117228 140830 117280 140836
rect 117148 132466 117268 132494
rect 117136 75608 117188 75614
rect 117136 75550 117188 75556
rect 117148 75206 117176 75550
rect 117136 75200 117188 75206
rect 117136 75142 117188 75148
rect 117240 74254 117268 132466
rect 117412 82136 117464 82142
rect 117412 82078 117464 82084
rect 117424 76770 117452 82078
rect 117700 79626 117728 141879
rect 117976 127634 118004 196726
rect 118240 192840 118292 192846
rect 118240 192782 118292 192788
rect 118054 192536 118110 192545
rect 118054 192471 118110 192480
rect 117964 127628 118016 127634
rect 117964 127570 118016 127576
rect 117872 122868 117924 122874
rect 117872 122810 117924 122816
rect 117688 79620 117740 79626
rect 117688 79562 117740 79568
rect 117884 76974 117912 122810
rect 117872 76968 117924 76974
rect 117872 76910 117924 76916
rect 117412 76764 117464 76770
rect 117412 76706 117464 76712
rect 117228 74248 117280 74254
rect 117228 74190 117280 74196
rect 117240 73914 117268 74190
rect 117228 73908 117280 73914
rect 117228 73850 117280 73856
rect 117044 71392 117096 71398
rect 117044 71334 117096 71340
rect 117976 70106 118004 127570
rect 118068 79286 118096 192471
rect 118148 191820 118200 191826
rect 118148 191762 118200 191768
rect 118160 191078 118188 191762
rect 118148 191072 118200 191078
rect 118148 191014 118200 191020
rect 118056 79280 118108 79286
rect 118056 79222 118108 79228
rect 118160 74526 118188 191014
rect 118252 75478 118280 192782
rect 118344 141710 118372 259490
rect 118424 193996 118476 194002
rect 118424 193938 118476 193944
rect 118332 141704 118384 141710
rect 118332 141646 118384 141652
rect 118240 75472 118292 75478
rect 118240 75414 118292 75420
rect 118148 74520 118200 74526
rect 118148 74462 118200 74468
rect 118436 74322 118464 193938
rect 118516 144424 118568 144430
rect 118516 144366 118568 144372
rect 118528 80850 118556 144366
rect 118620 142186 118648 260782
rect 118700 198756 118752 198762
rect 118700 198698 118752 198704
rect 118712 194410 118740 198698
rect 118700 194404 118752 194410
rect 118700 194346 118752 194352
rect 119080 142905 119108 263638
rect 119252 259480 119304 259486
rect 119252 259422 119304 259428
rect 119160 215348 119212 215354
rect 119160 215290 119212 215296
rect 119172 199102 119200 215290
rect 119160 199096 119212 199102
rect 119160 199038 119212 199044
rect 119264 144945 119292 259422
rect 119356 199442 119384 440234
rect 119436 316056 119488 316062
rect 119436 315998 119488 316004
rect 119448 200258 119476 315998
rect 119896 262540 119948 262546
rect 119896 262482 119948 262488
rect 119712 262200 119764 262206
rect 119712 262142 119764 262148
rect 119528 251252 119580 251258
rect 119528 251194 119580 251200
rect 119436 200252 119488 200258
rect 119436 200194 119488 200200
rect 119344 199436 119396 199442
rect 119344 199378 119396 199384
rect 119436 199368 119488 199374
rect 119436 199310 119488 199316
rect 119448 198830 119476 199310
rect 119540 199170 119568 251194
rect 119620 242956 119672 242962
rect 119620 242898 119672 242904
rect 119632 200666 119660 242898
rect 119620 200660 119672 200666
rect 119620 200602 119672 200608
rect 119528 199164 119580 199170
rect 119528 199106 119580 199112
rect 119436 198824 119488 198830
rect 119436 198766 119488 198772
rect 119528 192636 119580 192642
rect 119528 192578 119580 192584
rect 119436 190052 119488 190058
rect 119436 189994 119488 190000
rect 119344 144968 119396 144974
rect 119250 144936 119306 144945
rect 119344 144910 119396 144916
rect 119250 144871 119306 144880
rect 119066 142896 119122 142905
rect 119066 142831 119122 142840
rect 118608 142180 118660 142186
rect 118608 142122 118660 142128
rect 119356 141438 119384 144910
rect 119344 141432 119396 141438
rect 119344 141374 119396 141380
rect 119252 141296 119304 141302
rect 119252 141238 119304 141244
rect 118606 139360 118662 139369
rect 118606 139295 118662 139304
rect 118516 80844 118568 80850
rect 118516 80786 118568 80792
rect 118424 74316 118476 74322
rect 118424 74258 118476 74264
rect 118620 70310 118648 139295
rect 119160 104168 119212 104174
rect 119160 104110 119212 104116
rect 119172 76634 119200 104110
rect 119264 95946 119292 141238
rect 119342 138952 119398 138961
rect 119342 138887 119398 138896
rect 119252 95940 119304 95946
rect 119252 95882 119304 95888
rect 119250 95160 119306 95169
rect 119250 95095 119306 95104
rect 119160 76628 119212 76634
rect 119160 76570 119212 76576
rect 119264 74905 119292 95095
rect 119356 79558 119384 138887
rect 119448 89865 119476 189994
rect 119434 89856 119490 89865
rect 119434 89791 119490 89800
rect 119344 79552 119396 79558
rect 119344 79494 119396 79500
rect 119540 75342 119568 192578
rect 119620 181756 119672 181762
rect 119620 181698 119672 181704
rect 119528 75336 119580 75342
rect 119528 75278 119580 75284
rect 119250 74896 119306 74905
rect 119250 74831 119306 74840
rect 118608 70304 118660 70310
rect 118608 70246 118660 70252
rect 117964 70100 118016 70106
rect 117964 70042 118016 70048
rect 116216 68536 116268 68542
rect 116216 68478 116268 68484
rect 115478 67008 115534 67017
rect 115478 66943 115534 66952
rect 115020 63300 115072 63306
rect 115020 63242 115072 63248
rect 119632 63238 119660 181698
rect 119724 144974 119752 262142
rect 119908 147674 119936 262482
rect 120000 197470 120028 456758
rect 120092 259282 120120 605814
rect 120172 536852 120224 536858
rect 120172 536794 120224 536800
rect 120184 267734 120212 536794
rect 120184 267706 120488 267734
rect 120460 259298 120488 267706
rect 120080 259276 120132 259282
rect 120080 259218 120132 259224
rect 120184 259270 120612 259298
rect 120092 253314 120120 259218
rect 120184 253434 120212 259270
rect 120448 258800 120500 258806
rect 120448 258742 120500 258748
rect 120172 253428 120224 253434
rect 120172 253370 120224 253376
rect 120092 253286 120212 253314
rect 120080 253224 120132 253230
rect 120080 253166 120132 253172
rect 119988 197464 120040 197470
rect 119988 197406 120040 197412
rect 119988 193724 120040 193730
rect 119988 193666 120040 193672
rect 119816 147646 119936 147674
rect 119712 144968 119764 144974
rect 119712 144910 119764 144916
rect 119712 144356 119764 144362
rect 119712 144298 119764 144304
rect 119724 141114 119752 144298
rect 119816 142118 119844 147646
rect 119896 143472 119948 143478
rect 119896 143414 119948 143420
rect 119908 143274 119936 143414
rect 119896 143268 119948 143274
rect 119896 143210 119948 143216
rect 119804 142112 119856 142118
rect 119804 142054 119856 142060
rect 119724 141086 119844 141114
rect 119712 140344 119764 140350
rect 119712 140286 119764 140292
rect 119724 81394 119752 140286
rect 119712 81388 119764 81394
rect 119712 81330 119764 81336
rect 119816 80714 119844 141086
rect 119896 140752 119948 140758
rect 119896 140694 119948 140700
rect 119804 80708 119856 80714
rect 119804 80650 119856 80656
rect 119802 78568 119858 78577
rect 119802 78503 119858 78512
rect 119816 72865 119844 78503
rect 119908 72962 119936 140694
rect 119896 72956 119948 72962
rect 119896 72898 119948 72904
rect 119802 72856 119858 72865
rect 119802 72791 119858 72800
rect 120000 72418 120028 193666
rect 120092 143478 120120 253166
rect 120184 195294 120212 253286
rect 120262 198656 120318 198665
rect 120262 198591 120318 198600
rect 120276 197985 120304 198591
rect 120262 197976 120318 197985
rect 120262 197911 120318 197920
rect 120172 195288 120224 195294
rect 120172 195230 120224 195236
rect 120172 192908 120224 192914
rect 120172 192850 120224 192856
rect 120184 192506 120212 192850
rect 120172 192500 120224 192506
rect 120172 192442 120224 192448
rect 120080 143472 120132 143478
rect 120080 143414 120132 143420
rect 120184 137290 120212 192442
rect 120460 145761 120488 258742
rect 120632 223644 120684 223650
rect 120632 223586 120684 223592
rect 120644 223553 120672 223586
rect 120630 223544 120686 223553
rect 120630 223479 120686 223488
rect 120736 198898 120764 700266
rect 120816 448588 120868 448594
rect 120816 448530 120868 448536
rect 120724 198892 120776 198898
rect 120724 198834 120776 198840
rect 120736 198694 120764 198834
rect 120828 198830 120856 448530
rect 121276 385076 121328 385082
rect 121276 385018 121328 385024
rect 120908 347812 120960 347818
rect 120908 347754 120960 347760
rect 120816 198824 120868 198830
rect 120816 198766 120868 198772
rect 120920 198762 120948 347754
rect 121000 263764 121052 263770
rect 121000 263706 121052 263712
rect 121012 258806 121040 263706
rect 121288 259536 121316 385018
rect 122104 291236 122156 291242
rect 122104 291178 122156 291184
rect 122116 262954 122144 291178
rect 122104 262948 122156 262954
rect 122104 262890 122156 262896
rect 122852 260846 122880 700606
rect 124312 658300 124364 658306
rect 124312 658242 124364 658248
rect 122840 260840 122892 260846
rect 122840 260782 122892 260788
rect 122852 259978 122880 260782
rect 122852 259950 123096 259978
rect 124036 259956 124088 259962
rect 124036 259898 124088 259904
rect 123576 259616 123628 259622
rect 122562 259584 122618 259593
rect 122268 259542 122562 259570
rect 121196 259508 121316 259536
rect 123628 259564 123924 259570
rect 123576 259558 123924 259564
rect 123588 259542 123924 259558
rect 122562 259519 122618 259528
rect 121000 258800 121052 258806
rect 121000 258742 121052 258748
rect 121196 253934 121224 259508
rect 124048 259350 124076 259898
rect 124324 259570 124352 658242
rect 130384 565888 130436 565894
rect 130384 565830 130436 565836
rect 127164 503736 127216 503742
rect 127164 503678 127216 503684
rect 126244 452668 126296 452674
rect 126244 452610 126296 452616
rect 125692 320204 125744 320210
rect 125692 320146 125744 320152
rect 124864 275324 124916 275330
rect 124864 275266 124916 275272
rect 124876 259622 124904 275266
rect 125704 267734 125732 320146
rect 125704 267706 126008 267734
rect 125980 263594 126008 267706
rect 125980 263566 126100 263594
rect 125232 262268 125284 262274
rect 125232 262210 125284 262216
rect 125244 259978 125272 262210
rect 125244 259950 125580 259978
rect 126072 259894 126100 263566
rect 126256 263022 126284 452610
rect 126244 263016 126296 263022
rect 126244 262958 126296 262964
rect 126256 260234 126284 262958
rect 126978 262848 127034 262857
rect 126978 262783 127034 262792
rect 126992 262410 127020 262783
rect 126980 262404 127032 262410
rect 126980 262346 127032 262352
rect 127176 260250 127204 503678
rect 128360 469872 128412 469878
rect 128360 469814 128412 469820
rect 127900 263016 127952 263022
rect 127900 262958 127952 262964
rect 127716 262336 127768 262342
rect 127716 262278 127768 262284
rect 126244 260228 126296 260234
rect 127176 260222 127250 260250
rect 126244 260170 126296 260176
rect 127222 260166 127250 260222
rect 127210 260160 127262 260166
rect 127210 260102 127262 260108
rect 127222 259964 127250 260102
rect 127728 259978 127756 262278
rect 127912 262274 127940 262958
rect 127900 262268 127952 262274
rect 127900 262210 127952 262216
rect 128372 259978 128400 469814
rect 128452 336796 128504 336802
rect 128452 336738 128504 336744
rect 128464 260234 128492 336738
rect 130396 263673 130424 565830
rect 130382 263664 130438 263673
rect 130382 263599 130438 263608
rect 128452 260228 128504 260234
rect 128452 260170 128504 260176
rect 129694 260228 129746 260234
rect 129694 260170 129746 260176
rect 127728 259950 128064 259978
rect 128372 259950 128892 259978
rect 129706 259964 129734 260170
rect 130396 259978 130424 263599
rect 130396 259950 130548 259978
rect 126060 259888 126112 259894
rect 126112 259836 126408 259842
rect 126060 259830 126408 259836
rect 126072 259814 126408 259830
rect 128372 259826 128400 259950
rect 128360 259820 128412 259826
rect 128360 259762 128412 259768
rect 131132 259758 131160 701014
rect 133984 700534 134012 703520
rect 133972 700528 134024 700534
rect 133972 700470 134024 700476
rect 137848 700466 137876 703520
rect 137836 700460 137888 700466
rect 137836 700402 137888 700408
rect 141712 700398 141740 703520
rect 141700 700392 141752 700398
rect 141700 700334 141752 700340
rect 144932 699718 144960 703520
rect 148796 702434 148824 703520
rect 152660 702434 152688 703520
rect 156524 702434 156552 703520
rect 147692 702406 148824 702434
rect 151832 702406 152688 702434
rect 155972 702406 156552 702434
rect 144184 699712 144236 699718
rect 144184 699654 144236 699660
rect 144920 699712 144972 699718
rect 144920 699654 144972 699660
rect 144196 507890 144224 699654
rect 138664 507884 138716 507890
rect 138664 507826 138716 507832
rect 144184 507884 144236 507890
rect 144184 507826 144236 507832
rect 133880 273284 133932 273290
rect 133880 273226 133932 273232
rect 133892 267734 133920 273226
rect 133892 267706 134288 267734
rect 131304 263084 131356 263090
rect 131304 263026 131356 263032
rect 131316 259978 131344 263026
rect 133512 262744 133564 262750
rect 133512 262686 133564 262692
rect 132776 262336 132828 262342
rect 132776 262278 132828 262284
rect 132788 259978 132816 262278
rect 133524 259978 133552 262686
rect 134260 259978 134288 267706
rect 135444 264036 135496 264042
rect 135444 263978 135496 263984
rect 135260 262404 135312 262410
rect 135260 262346 135312 262352
rect 135272 259978 135300 262346
rect 135456 262342 135484 263978
rect 138676 263974 138704 507826
rect 147692 469878 147720 702406
rect 149704 700528 149756 700534
rect 149704 700470 149756 700476
rect 147680 469872 147732 469878
rect 147680 469814 147732 469820
rect 149716 407794 149744 700470
rect 149704 407788 149756 407794
rect 149704 407730 149756 407736
rect 145564 271924 145616 271930
rect 145564 271866 145616 271872
rect 145576 265878 145604 271866
rect 148968 269884 149020 269890
rect 148968 269826 149020 269832
rect 145564 265872 145616 265878
rect 145564 265814 145616 265820
rect 146760 264988 146812 264994
rect 146760 264930 146812 264936
rect 146208 264308 146260 264314
rect 146208 264250 146260 264256
rect 138664 263968 138716 263974
rect 138664 263910 138716 263916
rect 135444 262336 135496 262342
rect 135444 262278 135496 262284
rect 137652 262336 137704 262342
rect 137652 262278 137704 262284
rect 136824 262268 136876 262274
rect 136824 262210 136876 262216
rect 136836 259978 136864 262210
rect 137664 259978 137692 262278
rect 138676 259978 138704 263910
rect 145380 263900 145432 263906
rect 145380 263842 145432 263848
rect 143540 263220 143592 263226
rect 143540 263162 143592 263168
rect 141792 263152 141844 263158
rect 141792 263094 141844 263100
rect 140136 262676 140188 262682
rect 140136 262618 140188 262624
rect 139400 262608 139452 262614
rect 139400 262550 139452 262556
rect 139412 259978 139440 262550
rect 140148 259978 140176 262618
rect 141238 262440 141294 262449
rect 141238 262375 141294 262384
rect 141252 259978 141280 262375
rect 141804 259978 141832 263094
rect 142620 262472 142672 262478
rect 142620 262414 142672 262420
rect 142632 259978 142660 262414
rect 143552 259978 143580 263162
rect 144598 260228 144650 260234
rect 144598 260170 144650 260176
rect 131316 259950 131376 259978
rect 132788 259950 133032 259978
rect 133524 259950 133860 259978
rect 134260 259950 134688 259978
rect 135272 259950 135516 259978
rect 136836 259950 137172 259978
rect 137664 259950 138000 259978
rect 138676 259950 138828 259978
rect 139412 259950 139656 259978
rect 140148 259950 140484 259978
rect 141252 259950 141312 259978
rect 141804 259950 142140 259978
rect 142632 259950 142968 259978
rect 143552 259950 143796 259978
rect 144610 259964 144638 260170
rect 145392 259842 145420 263842
rect 146220 263838 146248 264250
rect 146208 263832 146260 263838
rect 146208 263774 146260 263780
rect 146220 259978 146248 263774
rect 146772 259978 146800 264930
rect 148980 264110 149008 269826
rect 151832 265742 151860 702406
rect 153108 267096 153160 267102
rect 153108 267038 153160 267044
rect 151820 265736 151872 265742
rect 151820 265678 151872 265684
rect 148968 264104 149020 264110
rect 148968 264046 149020 264052
rect 147680 262540 147732 262546
rect 147680 262482 147732 262488
rect 147692 259978 147720 262482
rect 148980 259978 149008 264046
rect 153120 263770 153148 267038
rect 155684 266416 155736 266422
rect 155684 266358 155736 266364
rect 152004 263764 152056 263770
rect 152004 263706 152056 263712
rect 153108 263764 153160 263770
rect 153108 263706 153160 263712
rect 150072 262812 150124 262818
rect 150072 262754 150124 262760
rect 149566 260092 149618 260098
rect 149566 260034 149618 260040
rect 146220 259950 146280 259978
rect 146772 259950 147108 259978
rect 147692 259950 147936 259978
rect 148764 259950 149008 259978
rect 149578 259964 149606 260034
rect 150084 259978 150112 262754
rect 150084 259950 150420 259978
rect 152016 259842 152044 263706
rect 152556 263696 152608 263702
rect 152556 263638 152608 263644
rect 152568 259978 152596 263638
rect 154486 262576 154542 262585
rect 154486 262511 154542 262520
rect 154500 259978 154528 262511
rect 155696 259978 155724 266358
rect 155972 265810 156000 702406
rect 164252 700466 164280 703520
rect 168116 700534 168144 703520
rect 171980 702434 172008 703520
rect 171152 702406 172008 702434
rect 168104 700528 168156 700534
rect 168104 700470 168156 700476
rect 164240 700460 164292 700466
rect 164240 700402 164292 700408
rect 167092 532772 167144 532778
rect 167092 532714 167144 532720
rect 165620 271176 165672 271182
rect 165620 271118 165672 271124
rect 161480 269816 161532 269822
rect 161480 269758 161532 269764
rect 156052 268388 156104 268394
rect 156052 268330 156104 268336
rect 155960 265804 156012 265810
rect 155960 265746 156012 265752
rect 156064 260302 156092 268330
rect 161492 264994 161520 269758
rect 165632 267734 165660 271118
rect 167104 267734 167132 532714
rect 171048 336048 171100 336054
rect 171048 335990 171100 335996
rect 165632 267706 165752 267734
rect 167104 267706 167408 267734
rect 162768 265056 162820 265062
rect 162768 264998 162820 265004
rect 161480 264988 161532 264994
rect 161480 264930 161532 264936
rect 159824 263628 159876 263634
rect 159824 263570 159876 263576
rect 157248 263084 157300 263090
rect 157248 263026 157300 263032
rect 156052 260296 156104 260302
rect 156052 260238 156104 260244
rect 152568 259950 152904 259978
rect 154500 259950 154560 259978
rect 155388 259950 155724 259978
rect 156064 259978 156092 260238
rect 157260 259978 157288 263026
rect 158168 260364 158220 260370
rect 158168 260306 158220 260312
rect 158180 259978 158208 260306
rect 158674 260160 158726 260166
rect 158674 260102 158726 260108
rect 156064 259950 156216 259978
rect 157044 259950 157288 259978
rect 157872 259950 158208 259978
rect 158686 259964 158714 260102
rect 159836 259978 159864 263570
rect 160652 263220 160704 263226
rect 160652 263162 160704 263168
rect 160664 259978 160692 263162
rect 161158 260228 161210 260234
rect 161158 260170 161210 260176
rect 159528 259950 159864 259978
rect 160356 259950 160692 259978
rect 161170 259964 161198 260170
rect 161492 259978 161520 264930
rect 162780 259978 162808 264998
rect 164424 262812 164476 262818
rect 164424 262754 164476 262760
rect 161492 259950 162012 259978
rect 162780 259950 162840 259978
rect 164436 259842 164464 262754
rect 165528 262608 165580 262614
rect 165528 262550 165580 262556
rect 165540 259978 165568 262550
rect 165324 259950 165568 259978
rect 165724 259978 165752 267706
rect 166906 262440 166962 262449
rect 166906 262375 166962 262384
rect 166920 259978 166948 262375
rect 167380 259978 167408 267706
rect 169760 265872 169812 265878
rect 169760 265814 169812 265820
rect 169668 263152 169720 263158
rect 169668 263094 169720 263100
rect 168932 262472 168984 262478
rect 168932 262414 168984 262420
rect 168944 259978 168972 262414
rect 169680 259978 169708 263094
rect 165724 259950 166488 259978
rect 166920 259950 166980 259978
rect 167380 259962 168144 259978
rect 167380 259956 168156 259962
rect 167380 259950 168104 259956
rect 145392 259814 145452 259842
rect 152016 259814 152076 259842
rect 164436 259814 164496 259842
rect 166460 259826 166488 259950
rect 168636 259950 168972 259978
rect 169464 259950 169708 259978
rect 168104 259898 168156 259904
rect 169772 259894 169800 265814
rect 171060 263673 171088 335990
rect 170586 263664 170642 263673
rect 170586 263599 170642 263608
rect 171046 263664 171102 263673
rect 171046 263599 171102 263608
rect 170600 259978 170628 263599
rect 171152 260137 171180 702406
rect 175844 700398 175872 703520
rect 179064 700602 179092 703520
rect 179052 700596 179104 700602
rect 179052 700538 179104 700544
rect 175832 700392 175884 700398
rect 175832 700334 175884 700340
rect 179328 645924 179380 645930
rect 179328 645866 179380 645872
rect 174544 278044 174596 278050
rect 174544 277986 174596 277992
rect 173072 265668 173124 265674
rect 173072 265610 173124 265616
rect 173084 263809 173112 265610
rect 174556 265130 174584 277986
rect 179340 265198 179368 645866
rect 180800 587920 180852 587926
rect 180800 587862 180852 587868
rect 180064 296744 180116 296750
rect 180064 296686 180116 296692
rect 179328 265192 179380 265198
rect 179328 265134 179380 265140
rect 174544 265124 174596 265130
rect 174544 265066 174596 265072
rect 173070 263800 173126 263809
rect 173070 263735 173126 263744
rect 172244 262540 172296 262546
rect 172244 262482 172296 262488
rect 171138 260128 171194 260137
rect 171138 260063 171194 260072
rect 172256 259978 172284 262482
rect 173084 259978 173112 263735
rect 174556 259978 174584 265066
rect 177212 262676 177264 262682
rect 177212 262618 177264 262624
rect 176384 260908 176436 260914
rect 176384 260850 176436 260856
rect 176396 259978 176424 260850
rect 177224 259978 177252 262618
rect 177948 262268 178000 262274
rect 177948 262210 178000 262216
rect 177960 259978 177988 262210
rect 170292 259950 170628 259978
rect 171948 259950 172284 259978
rect 172776 259950 173112 259978
rect 174432 259950 174584 259978
rect 176088 259950 176424 259978
rect 176916 259950 177252 259978
rect 177744 259950 177988 259978
rect 179340 259978 179368 265134
rect 180076 264314 180104 296686
rect 180064 264308 180116 264314
rect 180064 264250 180116 264256
rect 179880 262404 179932 262410
rect 179880 262346 179932 262352
rect 179892 261050 179920 262346
rect 179880 261044 179932 261050
rect 179880 260986 179932 260992
rect 179892 259978 179920 260986
rect 180812 259978 180840 587862
rect 182192 263090 182220 703582
rect 182744 703474 182772 703582
rect 182886 703520 182998 704960
rect 186750 703520 186862 704960
rect 190614 703520 190726 704960
rect 194478 703520 194590 704960
rect 198342 703520 198454 704960
rect 201512 703582 202092 703610
rect 182928 703474 182956 703520
rect 182744 703446 182956 703474
rect 189540 700596 189592 700602
rect 189540 700538 189592 700544
rect 189448 700392 189500 700398
rect 189448 700334 189500 700340
rect 183652 436144 183704 436150
rect 183652 436086 183704 436092
rect 182272 407788 182324 407794
rect 182272 407730 182324 407736
rect 182180 263084 182232 263090
rect 182180 263026 182232 263032
rect 182088 261044 182140 261050
rect 182088 260986 182140 260992
rect 181352 260024 181404 260030
rect 179340 259950 179400 259978
rect 179892 259950 180228 259978
rect 180812 259972 181352 259978
rect 182100 259978 182128 260986
rect 180812 259966 181404 259972
rect 180812 259950 181392 259966
rect 181884 259950 182128 259978
rect 182284 259978 182312 407730
rect 183664 267734 183692 436086
rect 184940 400240 184992 400246
rect 184940 400182 184992 400188
rect 183664 267706 183968 267734
rect 183468 263084 183520 263090
rect 183468 263026 183520 263032
rect 183480 262886 183508 263026
rect 183468 262880 183520 262886
rect 183468 262822 183520 262828
rect 183468 262744 183520 262750
rect 183468 262686 183520 262692
rect 182686 260092 182738 260098
rect 182686 260034 182738 260040
rect 182698 259978 182726 260034
rect 182284 259964 182726 259978
rect 183480 259978 183508 262686
rect 183940 259978 183968 267706
rect 184952 260001 184980 400182
rect 185492 263696 185544 263702
rect 185492 263638 185544 263644
rect 184938 259992 184994 260001
rect 182284 259950 182712 259964
rect 183480 259950 183540 259978
rect 183940 259950 184704 259978
rect 169760 259888 169812 259894
rect 169760 259830 169812 259836
rect 170956 259888 171008 259894
rect 171008 259836 171120 259842
rect 170956 259830 171120 259836
rect 166448 259820 166500 259826
rect 170968 259814 171120 259830
rect 166448 259762 166500 259768
rect 131120 259752 131172 259758
rect 131120 259694 131172 259700
rect 131856 259752 131908 259758
rect 163964 259752 164016 259758
rect 154026 259720 154082 259729
rect 131908 259700 132204 259706
rect 131856 259694 132204 259700
rect 131868 259678 132204 259694
rect 136008 259690 136344 259706
rect 135996 259684 136344 259690
rect 136048 259678 136344 259684
rect 153732 259678 154026 259706
rect 163668 259700 163964 259706
rect 163668 259694 164016 259700
rect 163668 259678 164004 259694
rect 184676 259690 184704 259950
rect 185504 259978 185532 263638
rect 188160 262948 188212 262954
rect 188160 262890 188212 262896
rect 187608 262336 187660 262342
rect 187608 262278 187660 262284
rect 185196 259950 185532 259978
rect 185858 259992 185914 260001
rect 184938 259927 184994 259936
rect 187620 259978 187648 262278
rect 188172 259978 188200 262890
rect 189080 260976 189132 260982
rect 189080 260918 189132 260924
rect 189092 259978 189120 260918
rect 185914 259950 186024 259978
rect 187620 259950 187680 259978
rect 188172 259950 188508 259978
rect 189092 259950 189336 259978
rect 185858 259927 185914 259936
rect 184664 259684 184716 259690
rect 154026 259655 154082 259664
rect 135996 259626 136048 259632
rect 184664 259626 184716 259632
rect 124864 259616 124916 259622
rect 124324 259542 124752 259570
rect 178868 259616 178920 259622
rect 124864 259558 124916 259564
rect 150912 259554 151248 259570
rect 150900 259548 151248 259554
rect 124416 259486 124444 259542
rect 150952 259542 151248 259548
rect 173604 259542 173848 259570
rect 175260 259554 175412 259570
rect 178572 259564 178868 259570
rect 187146 259584 187202 259593
rect 178572 259558 178920 259564
rect 175260 259548 175424 259554
rect 175260 259542 175372 259548
rect 150900 259490 150952 259496
rect 173820 259486 173848 259542
rect 178572 259542 178908 259558
rect 186852 259542 187146 259570
rect 187146 259519 187202 259528
rect 175372 259490 175424 259496
rect 124404 259480 124456 259486
rect 124404 259422 124456 259428
rect 173808 259480 173860 259486
rect 173808 259422 173860 259428
rect 124036 259344 124088 259350
rect 121288 259282 121440 259298
rect 124036 259286 124088 259292
rect 121276 259276 121440 259282
rect 121328 259270 121440 259276
rect 121276 259218 121328 259224
rect 121196 253906 121316 253934
rect 120998 223544 121054 223553
rect 120998 223479 121054 223488
rect 121012 198898 121040 223479
rect 121000 198892 121052 198898
rect 121000 198834 121052 198840
rect 120908 198756 120960 198762
rect 120908 198698 120960 198704
rect 120724 198688 120776 198694
rect 121288 198665 121316 253906
rect 178224 200728 178276 200734
rect 178224 200670 178276 200676
rect 181904 200728 181956 200734
rect 181904 200670 181956 200676
rect 182824 200728 182876 200734
rect 182824 200670 182876 200676
rect 187606 200696 187662 200705
rect 131856 200660 131908 200666
rect 131856 200602 131908 200608
rect 177856 200660 177908 200666
rect 177856 200602 177908 200608
rect 178040 200660 178092 200666
rect 178040 200602 178092 200608
rect 131670 200560 131726 200569
rect 131670 200495 131726 200504
rect 122840 200252 122892 200258
rect 122840 200194 122892 200200
rect 124864 200252 124916 200258
rect 124864 200194 124916 200200
rect 121920 199368 121972 199374
rect 121920 199310 121972 199316
rect 120724 198630 120776 198636
rect 121274 198656 121330 198665
rect 121274 198591 121330 198600
rect 121460 195288 121512 195294
rect 121460 195230 121512 195236
rect 121276 192704 121328 192710
rect 121276 192646 121328 192652
rect 121000 190120 121052 190126
rect 121000 190062 121052 190068
rect 120540 182912 120592 182918
rect 120540 182854 120592 182860
rect 120446 145752 120502 145761
rect 120446 145687 120502 145696
rect 120172 137284 120224 137290
rect 120172 137226 120224 137232
rect 120080 76900 120132 76906
rect 120080 76842 120132 76848
rect 120092 76430 120120 76842
rect 120080 76424 120132 76430
rect 120080 76366 120132 76372
rect 120080 75200 120132 75206
rect 120080 75142 120132 75148
rect 119988 72412 120040 72418
rect 119988 72354 120040 72360
rect 119620 63232 119672 63238
rect 119620 63174 119672 63180
rect 120092 16574 120120 75142
rect 120552 66162 120580 182854
rect 120724 148164 120776 148170
rect 120724 148106 120776 148112
rect 120632 142248 120684 142254
rect 120632 142190 120684 142196
rect 120644 116618 120672 142190
rect 120632 116612 120684 116618
rect 120632 116554 120684 116560
rect 120632 110628 120684 110634
rect 120632 110570 120684 110576
rect 120644 66842 120672 110570
rect 120736 93158 120764 148106
rect 120908 147620 120960 147626
rect 120908 147562 120960 147568
rect 120920 142730 120948 147562
rect 120908 142724 120960 142730
rect 120908 142666 120960 142672
rect 120816 140616 120868 140622
rect 120816 140558 120868 140564
rect 120724 93152 120776 93158
rect 120724 93094 120776 93100
rect 120722 80200 120778 80209
rect 120722 80135 120778 80144
rect 120736 68406 120764 80135
rect 120828 77994 120856 140558
rect 120906 139360 120962 139369
rect 120906 139295 120962 139304
rect 120816 77988 120868 77994
rect 120816 77930 120868 77936
rect 120920 72622 120948 139295
rect 121012 76430 121040 190062
rect 121092 186992 121144 186998
rect 121092 186934 121144 186940
rect 121000 76424 121052 76430
rect 121000 76366 121052 76372
rect 121104 73098 121132 186934
rect 121184 148232 121236 148238
rect 121184 148174 121236 148180
rect 121092 73092 121144 73098
rect 121092 73034 121144 73040
rect 120908 72616 120960 72622
rect 120908 72558 120960 72564
rect 120724 68400 120776 68406
rect 120724 68342 120776 68348
rect 120632 66836 120684 66842
rect 120632 66778 120684 66784
rect 121196 66230 121224 148174
rect 121288 76906 121316 192646
rect 121472 143478 121500 195230
rect 121828 192432 121880 192438
rect 121828 192374 121880 192380
rect 121368 143472 121420 143478
rect 121368 143414 121420 143420
rect 121460 143472 121512 143478
rect 121460 143414 121512 143420
rect 121380 139890 121408 143414
rect 121380 139862 121440 139890
rect 121734 138816 121790 138825
rect 121734 138751 121790 138760
rect 121748 138553 121776 138751
rect 121734 138544 121790 138553
rect 121734 138479 121790 138488
rect 121734 138136 121790 138145
rect 121734 138071 121790 138080
rect 121748 135969 121776 138071
rect 121734 135960 121790 135969
rect 121734 135895 121790 135904
rect 121734 89856 121790 89865
rect 121734 89791 121790 89800
rect 121644 81388 121696 81394
rect 121644 81330 121696 81336
rect 121552 81116 121604 81122
rect 121552 81058 121604 81064
rect 121276 76900 121328 76906
rect 121276 76842 121328 76848
rect 121564 66978 121592 81058
rect 121552 66972 121604 66978
rect 121552 66914 121604 66920
rect 121656 66774 121684 81330
rect 121748 71738 121776 89791
rect 121840 78606 121868 192374
rect 121932 80646 121960 199310
rect 122852 197849 122880 200194
rect 124876 199850 124904 200194
rect 129738 200016 129794 200025
rect 129738 199951 129794 199960
rect 128544 199912 128596 199918
rect 128358 199880 128414 199889
rect 124864 199844 124916 199850
rect 124864 199786 124916 199792
rect 124956 199844 125008 199850
rect 128544 199854 128596 199860
rect 128358 199815 128414 199824
rect 124956 199786 125008 199792
rect 124312 199572 124364 199578
rect 124312 199514 124364 199520
rect 122932 199164 122984 199170
rect 122932 199106 122984 199112
rect 122838 197840 122894 197849
rect 122838 197775 122894 197784
rect 122470 197432 122526 197441
rect 122470 197367 122526 197376
rect 122484 195945 122512 197367
rect 122470 195936 122526 195945
rect 122470 195871 122526 195880
rect 122838 195936 122894 195945
rect 122838 195871 122894 195880
rect 122104 194472 122156 194478
rect 122104 194414 122156 194420
rect 122012 191276 122064 191282
rect 122012 191218 122064 191224
rect 121920 80640 121972 80646
rect 121920 80582 121972 80588
rect 121828 78600 121880 78606
rect 121828 78542 121880 78548
rect 121736 71732 121788 71738
rect 121736 71674 121788 71680
rect 122024 70038 122052 191218
rect 122012 70032 122064 70038
rect 122012 69974 122064 69980
rect 121644 66768 121696 66774
rect 121644 66710 121696 66716
rect 121184 66224 121236 66230
rect 121184 66166 121236 66172
rect 120540 66156 120592 66162
rect 120540 66098 120592 66104
rect 122116 48278 122144 194414
rect 122484 190505 122512 195871
rect 122470 190496 122526 190505
rect 122470 190431 122526 190440
rect 122746 189544 122802 189553
rect 122746 189479 122802 189488
rect 122760 181529 122788 189479
rect 122746 181520 122802 181529
rect 122746 181455 122802 181464
rect 122746 180704 122802 180713
rect 122746 180639 122802 180648
rect 122760 171193 122788 180639
rect 122746 171184 122802 171193
rect 122746 171119 122802 171128
rect 122746 171048 122802 171057
rect 122746 170983 122802 170992
rect 122760 161537 122788 170983
rect 122746 161528 122802 161537
rect 122746 161463 122802 161472
rect 122746 161392 122802 161401
rect 122746 161327 122802 161336
rect 122760 151881 122788 161327
rect 122746 151872 122802 151881
rect 122746 151807 122802 151816
rect 122746 151736 122802 151745
rect 122746 151671 122802 151680
rect 122760 147665 122788 151671
rect 122746 147656 122802 147665
rect 122746 147591 122802 147600
rect 122196 143472 122248 143478
rect 122196 143414 122248 143420
rect 122208 139890 122236 143414
rect 122852 142254 122880 195871
rect 122944 151814 122972 199106
rect 124220 198824 124272 198830
rect 124220 198766 124272 198772
rect 123482 197840 123538 197849
rect 123482 197775 123538 197784
rect 123116 182164 123168 182170
rect 123116 182106 123168 182112
rect 123128 181014 123156 182106
rect 123116 181008 123168 181014
rect 123116 180950 123168 180956
rect 123128 180402 123156 180950
rect 123116 180396 123168 180402
rect 123116 180338 123168 180344
rect 123496 151814 123524 197775
rect 124128 195152 124180 195158
rect 124128 195094 124180 195100
rect 123574 194304 123630 194313
rect 123574 194239 123630 194248
rect 123588 182170 123616 194239
rect 123576 182164 123628 182170
rect 123576 182106 123628 182112
rect 124140 177954 124168 195094
rect 124128 177948 124180 177954
rect 124128 177890 124180 177896
rect 124036 173936 124088 173942
rect 124036 173878 124088 173884
rect 124048 151814 124076 173878
rect 122944 151786 123248 151814
rect 122840 142248 122892 142254
rect 122840 142190 122892 142196
rect 122852 139890 122880 142190
rect 122208 139862 122268 139890
rect 122852 139862 123096 139890
rect 123220 139330 123248 151786
rect 123404 151786 123524 151814
rect 123588 151786 124076 151814
rect 123404 145518 123432 151786
rect 123392 145512 123444 145518
rect 123392 145454 123444 145460
rect 123588 139369 123616 151786
rect 123668 142180 123720 142186
rect 123668 142122 123720 142128
rect 123680 139890 123708 142122
rect 123680 139862 123924 139890
rect 124140 139369 124168 177890
rect 124232 145382 124260 198766
rect 124220 145376 124272 145382
rect 124220 145318 124272 145324
rect 124324 143528 124352 199514
rect 124968 199209 124996 199786
rect 125508 199708 125560 199714
rect 125508 199650 125560 199656
rect 125520 199578 125548 199650
rect 125508 199572 125560 199578
rect 125508 199514 125560 199520
rect 126796 199436 126848 199442
rect 126796 199378 126848 199384
rect 124954 199200 125010 199209
rect 124954 199135 125010 199144
rect 125508 198484 125560 198490
rect 125508 198426 125560 198432
rect 125416 196920 125468 196926
rect 125416 196862 125468 196868
rect 125428 196110 125456 196862
rect 124404 196104 124456 196110
rect 124404 196046 124456 196052
rect 125416 196104 125468 196110
rect 125416 196046 125468 196052
rect 124232 143500 124352 143528
rect 124232 139641 124260 143500
rect 124416 143426 124444 196046
rect 124864 187808 124916 187814
rect 124864 187750 124916 187756
rect 124324 143398 124444 143426
rect 124324 140758 124352 143398
rect 124402 143304 124458 143313
rect 124402 143239 124458 143248
rect 124312 140752 124364 140758
rect 124312 140694 124364 140700
rect 124416 139890 124444 143239
rect 124876 139942 124904 187750
rect 125520 182170 125548 198426
rect 126520 198280 126572 198286
rect 126520 198222 126572 198228
rect 126426 197976 126482 197985
rect 126256 197934 126426 197962
rect 125692 197668 125744 197674
rect 125692 197610 125744 197616
rect 125600 197464 125652 197470
rect 125600 197406 125652 197412
rect 125508 182164 125560 182170
rect 125508 182106 125560 182112
rect 125612 148617 125640 197406
rect 125704 191894 125732 197610
rect 125692 191888 125744 191894
rect 125692 191830 125744 191836
rect 125598 148608 125654 148617
rect 125598 148543 125654 148552
rect 125704 148170 125732 191830
rect 125784 182164 125836 182170
rect 125784 182106 125836 182112
rect 125796 181490 125824 182106
rect 125784 181484 125836 181490
rect 125784 181426 125836 181432
rect 125796 148481 125824 181426
rect 125782 148472 125838 148481
rect 125782 148407 125838 148416
rect 125692 148164 125744 148170
rect 125692 148106 125744 148112
rect 125230 144936 125286 144945
rect 125230 144871 125286 144880
rect 124864 139936 124916 139942
rect 124416 139862 124752 139890
rect 124864 139878 124916 139884
rect 125244 139890 125272 144871
rect 126060 142792 126112 142798
rect 126060 142734 126112 142740
rect 126072 139890 126100 142734
rect 126256 141982 126284 197934
rect 126426 197911 126482 197920
rect 126336 195288 126388 195294
rect 126336 195230 126388 195236
rect 126244 141976 126296 141982
rect 126244 141918 126296 141924
rect 126348 141302 126376 195230
rect 126428 192500 126480 192506
rect 126428 192442 126480 192448
rect 126336 141296 126388 141302
rect 126336 141238 126388 141244
rect 126440 140690 126468 192442
rect 126532 148986 126560 198222
rect 126808 197985 126836 199378
rect 126888 198620 126940 198626
rect 126888 198562 126940 198568
rect 126794 197976 126850 197985
rect 126794 197911 126850 197920
rect 126612 197532 126664 197538
rect 126612 197474 126664 197480
rect 126624 178129 126652 197474
rect 126900 197470 126928 198562
rect 128176 198416 128228 198422
rect 128176 198358 128228 198364
rect 127992 197940 128044 197946
rect 127992 197882 128044 197888
rect 127808 197872 127860 197878
rect 127808 197814 127860 197820
rect 126888 197464 126940 197470
rect 126888 197406 126940 197412
rect 126702 194440 126758 194449
rect 126702 194375 126758 194384
rect 126716 179382 126744 194375
rect 127624 192772 127676 192778
rect 127624 192714 127676 192720
rect 126888 180940 126940 180946
rect 126888 180882 126940 180888
rect 126900 180742 126928 180882
rect 126888 180736 126940 180742
rect 126888 180678 126940 180684
rect 126704 179376 126756 179382
rect 126704 179318 126756 179324
rect 126610 178120 126666 178129
rect 126610 178055 126666 178064
rect 126624 178022 126652 178055
rect 126612 178016 126664 178022
rect 126612 177958 126664 177964
rect 126520 148980 126572 148986
rect 126520 148922 126572 148928
rect 126980 143268 127032 143274
rect 126980 143210 127032 143216
rect 127072 143268 127124 143274
rect 127072 143210 127124 143216
rect 126428 140684 126480 140690
rect 126428 140626 126480 140632
rect 126992 139890 127020 143210
rect 127084 142730 127112 143210
rect 127072 142724 127124 142730
rect 127072 142666 127124 142672
rect 125244 139862 125580 139890
rect 126072 139862 126408 139890
rect 126992 139862 127236 139890
rect 124218 139632 124274 139641
rect 124218 139567 124274 139576
rect 127636 139369 127664 192714
rect 127716 191820 127768 191826
rect 127716 191762 127768 191768
rect 127728 147674 127756 191762
rect 127820 148238 127848 197814
rect 127900 185904 127952 185910
rect 127900 185846 127952 185852
rect 127912 148306 127940 185846
rect 128004 181257 128032 197882
rect 127990 181248 128046 181257
rect 127990 181183 128046 181192
rect 128004 180674 128032 181183
rect 128188 180849 128216 198358
rect 128372 197402 128400 199815
rect 128452 198144 128504 198150
rect 128452 198086 128504 198092
rect 128360 197396 128412 197402
rect 128360 197338 128412 197344
rect 128360 196036 128412 196042
rect 128360 195978 128412 195984
rect 128174 180840 128230 180849
rect 128174 180775 128230 180784
rect 127992 180668 128044 180674
rect 127992 180610 128044 180616
rect 128188 180538 128216 180775
rect 128176 180532 128228 180538
rect 128176 180474 128228 180480
rect 127900 148300 127952 148306
rect 127900 148242 127952 148248
rect 127808 148232 127860 148238
rect 127808 148174 127860 148180
rect 127728 147646 127848 147674
rect 127716 145444 127768 145450
rect 127716 145386 127768 145392
rect 127728 139890 127756 145386
rect 127820 141914 127848 147646
rect 128372 144090 128400 195978
rect 128464 191826 128492 198086
rect 128556 194041 128584 199854
rect 129188 198552 129240 198558
rect 129188 198494 129240 198500
rect 128542 194032 128598 194041
rect 128542 193967 128598 193976
rect 128452 191820 128504 191826
rect 128452 191762 128504 191768
rect 129094 189000 129150 189009
rect 129094 188935 129150 188944
rect 129004 188760 129056 188766
rect 129004 188702 129056 188708
rect 128726 181112 128782 181121
rect 128726 181047 128782 181056
rect 128740 180470 128768 181047
rect 128728 180464 128780 180470
rect 128728 180406 128780 180412
rect 128360 144084 128412 144090
rect 128360 144026 128412 144032
rect 128544 143540 128596 143546
rect 128544 143482 128596 143488
rect 127808 141908 127860 141914
rect 127808 141850 127860 141856
rect 128556 139890 128584 143482
rect 129016 142154 129044 188702
rect 129108 148753 129136 188935
rect 129200 180985 129228 198494
rect 129648 198348 129700 198354
rect 129648 198290 129700 198296
rect 129660 198150 129688 198290
rect 129752 198218 129780 199951
rect 131684 199714 131712 200495
rect 131764 199912 131816 199918
rect 131764 199854 131816 199860
rect 131672 199708 131724 199714
rect 131672 199650 131724 199656
rect 131776 199578 131804 199854
rect 131764 199572 131816 199578
rect 131764 199514 131816 199520
rect 131212 199436 131264 199442
rect 131212 199378 131264 199384
rect 130934 199200 130990 199209
rect 130934 199135 130990 199144
rect 130948 198626 130976 199135
rect 130936 198620 130988 198626
rect 130936 198562 130988 198568
rect 129740 198212 129792 198218
rect 129740 198154 129792 198160
rect 129648 198144 129700 198150
rect 129648 198086 129700 198092
rect 130660 197056 130712 197062
rect 130660 196998 130712 197004
rect 129646 196480 129702 196489
rect 129646 196415 129702 196424
rect 129660 189009 129688 196415
rect 130384 195968 130436 195974
rect 130384 195910 130436 195916
rect 129646 189000 129702 189009
rect 129646 188935 129702 188944
rect 129740 186380 129792 186386
rect 129740 186322 129792 186328
rect 129752 186182 129780 186322
rect 129740 186176 129792 186182
rect 129740 186118 129792 186124
rect 129186 180976 129242 180985
rect 129186 180911 129242 180920
rect 129200 180810 129228 180911
rect 129648 180872 129700 180878
rect 129648 180814 129700 180820
rect 129188 180804 129240 180810
rect 129188 180746 129240 180752
rect 129660 180606 129688 180814
rect 129648 180600 129700 180606
rect 129648 180542 129700 180548
rect 129094 148744 129150 148753
rect 129094 148679 129150 148688
rect 130396 148374 130424 195910
rect 130476 191820 130528 191826
rect 130476 191762 130528 191768
rect 130384 148368 130436 148374
rect 130384 148310 130436 148316
rect 130108 146260 130160 146266
rect 130108 146202 130160 146208
rect 129372 146192 129424 146198
rect 129372 146134 129424 146140
rect 129016 142126 129228 142154
rect 127728 139862 128064 139890
rect 128556 139862 128892 139890
rect 129200 139369 129228 142126
rect 129384 139890 129412 146134
rect 130120 139890 130148 146202
rect 130488 140146 130516 191762
rect 130476 140140 130528 140146
rect 130476 140082 130528 140088
rect 129384 139862 129720 139890
rect 130120 139862 130548 139890
rect 123574 139360 123630 139369
rect 123208 139324 123260 139330
rect 123574 139295 123630 139304
rect 124126 139360 124182 139369
rect 124126 139295 124182 139304
rect 127622 139360 127678 139369
rect 127622 139295 127678 139304
rect 129186 139360 129242 139369
rect 130672 139346 130700 196998
rect 131028 193656 131080 193662
rect 131028 193598 131080 193604
rect 130752 187876 130804 187882
rect 130752 187818 130804 187824
rect 130764 151814 130792 187818
rect 130764 151786 130884 151814
rect 130856 139505 130884 151786
rect 131040 140146 131068 193598
rect 131118 185056 131174 185065
rect 131118 184991 131174 185000
rect 131132 184890 131160 184991
rect 131120 184884 131172 184890
rect 131120 184826 131172 184832
rect 131118 143168 131174 143177
rect 131118 143103 131174 143112
rect 131028 140140 131080 140146
rect 131028 140082 131080 140088
rect 131132 139890 131160 143103
rect 131224 141953 131252 199378
rect 131762 199336 131818 199345
rect 131762 199271 131818 199280
rect 131304 198756 131356 198762
rect 131304 198698 131356 198704
rect 131316 149054 131344 198698
rect 131776 197946 131804 199271
rect 131868 198801 131896 200602
rect 177764 200592 177816 200598
rect 177764 200534 177816 200540
rect 177776 200433 177804 200534
rect 177762 200424 177818 200433
rect 132040 200388 132092 200394
rect 177762 200359 177818 200368
rect 132040 200330 132092 200336
rect 131948 199980 132000 199986
rect 131948 199922 132000 199928
rect 131854 198792 131910 198801
rect 131854 198727 131910 198736
rect 131764 197940 131816 197946
rect 131764 197882 131816 197888
rect 131764 196376 131816 196382
rect 131764 196318 131816 196324
rect 131776 151814 131804 196318
rect 131592 151786 131804 151814
rect 131304 149048 131356 149054
rect 131304 148990 131356 148996
rect 131592 142154 131620 151786
rect 131868 146282 131896 198727
rect 131960 198082 131988 199922
rect 132052 199209 132080 200330
rect 177868 200326 177896 200602
rect 177948 200524 178000 200530
rect 177948 200466 178000 200472
rect 177856 200320 177908 200326
rect 177856 200262 177908 200268
rect 177960 200190 177988 200466
rect 177948 200184 178000 200190
rect 132374 200114 132402 200124
rect 132328 200086 132402 200114
rect 132224 199912 132276 199918
rect 132224 199854 132276 199860
rect 132132 199776 132184 199782
rect 132132 199718 132184 199724
rect 132038 199200 132094 199209
rect 132038 199135 132094 199144
rect 132144 198665 132172 199718
rect 132236 199646 132264 199854
rect 132224 199640 132276 199646
rect 132224 199582 132276 199588
rect 132224 199436 132276 199442
rect 132224 199378 132276 199384
rect 132236 199238 132264 199378
rect 132224 199232 132276 199238
rect 132224 199174 132276 199180
rect 132130 198656 132186 198665
rect 132130 198591 132186 198600
rect 131948 198076 132000 198082
rect 131948 198018 132000 198024
rect 132132 197600 132184 197606
rect 132132 197542 132184 197548
rect 132040 194812 132092 194818
rect 132040 194754 132092 194760
rect 131948 192364 132000 192370
rect 131948 192306 132000 192312
rect 131684 146254 131896 146282
rect 131684 144158 131712 146254
rect 131854 146024 131910 146033
rect 131854 145959 131910 145968
rect 131672 144152 131724 144158
rect 131672 144094 131724 144100
rect 131592 142126 131712 142154
rect 131210 141944 131266 141953
rect 131210 141879 131266 141888
rect 131684 140554 131712 142126
rect 131672 140548 131724 140554
rect 131672 140490 131724 140496
rect 131868 139890 131896 145959
rect 131960 140486 131988 192306
rect 132052 151298 132080 194754
rect 132144 184074 132172 197542
rect 132224 196512 132276 196518
rect 132224 196454 132276 196460
rect 132236 184142 132264 196454
rect 132328 195974 132356 200086
rect 132466 199968 132494 200124
rect 132420 199940 132494 199968
rect 132420 198762 132448 199940
rect 132558 199866 132586 200124
rect 132512 199838 132586 199866
rect 132512 199782 132540 199838
rect 132500 199776 132552 199782
rect 132650 199764 132678 200124
rect 132742 199889 132770 200124
rect 132834 199918 132862 200124
rect 132822 199912 132874 199918
rect 132728 199880 132784 199889
rect 132822 199854 132874 199860
rect 132728 199815 132784 199824
rect 132500 199718 132552 199724
rect 132604 199736 132678 199764
rect 132498 199336 132554 199345
rect 132498 199271 132554 199280
rect 132512 198762 132540 199271
rect 132408 198756 132460 198762
rect 132408 198698 132460 198704
rect 132500 198756 132552 198762
rect 132500 198698 132552 198704
rect 132316 195968 132368 195974
rect 132316 195910 132368 195916
rect 132604 188358 132632 199736
rect 132776 199640 132828 199646
rect 132926 199628 132954 200124
rect 133018 199782 133046 200124
rect 133110 199889 133138 200124
rect 133096 199880 133152 199889
rect 133096 199815 133152 199824
rect 133006 199776 133058 199782
rect 133006 199718 133058 199724
rect 133098 199776 133150 199782
rect 133202 199764 133230 200124
rect 133294 199850 133322 200124
rect 133282 199844 133334 199850
rect 133282 199786 133334 199792
rect 133386 199782 133414 200124
rect 133150 199736 133230 199764
rect 133374 199776 133426 199782
rect 133098 199718 133150 199724
rect 133374 199718 133426 199724
rect 133236 199640 133288 199646
rect 132926 199600 133092 199628
rect 132776 199582 132828 199588
rect 132788 191834 132816 199582
rect 133064 198694 133092 199600
rect 133236 199582 133288 199588
rect 133142 199336 133198 199345
rect 133142 199271 133198 199280
rect 133052 198688 133104 198694
rect 133052 198630 133104 198636
rect 132960 198076 133012 198082
rect 132960 198018 133012 198024
rect 132696 191806 132816 191834
rect 132592 188352 132644 188358
rect 132592 188294 132644 188300
rect 132224 184136 132276 184142
rect 132224 184078 132276 184084
rect 132132 184068 132184 184074
rect 132132 184010 132184 184016
rect 132696 175982 132724 191806
rect 132868 191004 132920 191010
rect 132868 190946 132920 190952
rect 132776 190936 132828 190942
rect 132776 190878 132828 190884
rect 132788 181558 132816 190878
rect 132880 183938 132908 190946
rect 132972 185910 133000 198018
rect 133156 197520 133184 199271
rect 133248 198082 133276 199582
rect 133478 199560 133506 200124
rect 133570 199889 133598 200124
rect 133556 199880 133612 199889
rect 133662 199850 133690 200124
rect 133754 199850 133782 200124
rect 133556 199815 133612 199824
rect 133650 199844 133702 199850
rect 133650 199786 133702 199792
rect 133742 199844 133794 199850
rect 133742 199786 133794 199792
rect 133846 199730 133874 200124
rect 133938 199918 133966 200124
rect 133926 199912 133978 199918
rect 133926 199854 133978 199860
rect 134030 199764 134058 200124
rect 134122 199889 134150 200124
rect 134108 199880 134164 199889
rect 134108 199815 134164 199824
rect 133984 199736 134058 199764
rect 134214 199764 134242 200124
rect 134306 199918 134334 200124
rect 134294 199912 134346 199918
rect 134398 199889 134426 200124
rect 134490 199918 134518 200124
rect 134582 199918 134610 200124
rect 134478 199912 134530 199918
rect 134294 199854 134346 199860
rect 134384 199880 134440 199889
rect 134478 199854 134530 199860
rect 134570 199912 134622 199918
rect 134570 199854 134622 199860
rect 134384 199815 134440 199824
rect 134674 199764 134702 200124
rect 134766 199923 134794 200124
rect 134752 199914 134808 199923
rect 134858 199918 134886 200124
rect 134752 199849 134808 199858
rect 134846 199912 134898 199918
rect 134846 199854 134898 199860
rect 134950 199782 134978 200124
rect 134214 199736 134288 199764
rect 133846 199702 133920 199730
rect 133604 199640 133656 199646
rect 133604 199582 133656 199588
rect 133696 199640 133748 199646
rect 133696 199582 133748 199588
rect 133478 199532 133552 199560
rect 133524 199345 133552 199532
rect 133510 199336 133566 199345
rect 133510 199271 133566 199280
rect 133510 199200 133566 199209
rect 133510 199135 133566 199144
rect 133418 198792 133474 198801
rect 133418 198727 133474 198736
rect 133236 198076 133288 198082
rect 133236 198018 133288 198024
rect 133156 197492 133276 197520
rect 133144 197396 133196 197402
rect 133144 197338 133196 197344
rect 133052 195628 133104 195634
rect 133052 195570 133104 195576
rect 133064 195294 133092 195570
rect 133052 195288 133104 195294
rect 133052 195230 133104 195236
rect 132960 185904 133012 185910
rect 132960 185846 133012 185852
rect 132868 183932 132920 183938
rect 132868 183874 132920 183880
rect 132776 181552 132828 181558
rect 132776 181494 132828 181500
rect 132684 175976 132736 175982
rect 132684 175918 132736 175924
rect 132040 151292 132092 151298
rect 132040 151234 132092 151240
rect 133156 148510 133184 197338
rect 133248 148714 133276 197492
rect 133432 187270 133460 198727
rect 133524 198014 133552 199135
rect 133512 198008 133564 198014
rect 133512 197950 133564 197956
rect 133510 195936 133566 195945
rect 133510 195871 133566 195880
rect 133420 187264 133472 187270
rect 133420 187206 133472 187212
rect 133524 186314 133552 195871
rect 133616 191010 133644 199582
rect 133708 191834 133736 199582
rect 133786 199200 133842 199209
rect 133786 199135 133842 199144
rect 133800 194313 133828 199135
rect 133892 197402 133920 199702
rect 133880 197396 133932 197402
rect 133880 197338 133932 197344
rect 133984 197334 134012 199736
rect 134260 199730 134288 199736
rect 134628 199736 134702 199764
rect 134800 199776 134852 199782
rect 134260 199714 134380 199730
rect 134260 199708 134392 199714
rect 134260 199702 134340 199708
rect 134340 199650 134392 199656
rect 134432 199708 134484 199714
rect 134432 199650 134484 199656
rect 134524 199708 134576 199714
rect 134524 199650 134576 199656
rect 134064 199640 134116 199646
rect 134064 199582 134116 199588
rect 134248 199640 134300 199646
rect 134248 199582 134300 199588
rect 133972 197328 134024 197334
rect 133972 197270 134024 197276
rect 133972 196988 134024 196994
rect 133972 196930 134024 196936
rect 133984 196042 134012 196930
rect 133972 196036 134024 196042
rect 133972 195978 134024 195984
rect 133786 194304 133842 194313
rect 133786 194239 133842 194248
rect 133708 191806 133828 191834
rect 133604 191004 133656 191010
rect 133604 190946 133656 190952
rect 133800 190942 133828 191806
rect 133880 191820 133932 191826
rect 133880 191762 133932 191768
rect 133892 191418 133920 191762
rect 133880 191412 133932 191418
rect 133880 191354 133932 191360
rect 133788 190936 133840 190942
rect 133788 190878 133840 190884
rect 133340 186286 133552 186314
rect 133236 148708 133288 148714
rect 133236 148650 133288 148656
rect 133340 148646 133368 186286
rect 134076 178838 134104 199582
rect 134154 199336 134210 199345
rect 134154 199271 134210 199280
rect 134168 198286 134196 199271
rect 134156 198280 134208 198286
rect 134156 198222 134208 198228
rect 134260 191826 134288 199582
rect 134340 199572 134392 199578
rect 134340 199514 134392 199520
rect 134352 198801 134380 199514
rect 134338 198792 134394 198801
rect 134338 198727 134394 198736
rect 134340 197328 134392 197334
rect 134340 197270 134392 197276
rect 134248 191820 134300 191826
rect 134248 191762 134300 191768
rect 134352 191706 134380 197270
rect 134260 191678 134380 191706
rect 134156 191412 134208 191418
rect 134156 191354 134208 191360
rect 134168 178974 134196 191354
rect 134260 191026 134288 191678
rect 134444 191418 134472 199650
rect 134536 194818 134564 199650
rect 134524 194812 134576 194818
rect 134524 194754 134576 194760
rect 134432 191412 134484 191418
rect 134432 191354 134484 191360
rect 134260 190998 134380 191026
rect 134628 191010 134656 199736
rect 134800 199718 134852 199724
rect 134938 199776 134990 199782
rect 134938 199718 134990 199724
rect 134812 199424 134840 199718
rect 135042 199696 135070 200124
rect 135134 199918 135162 200124
rect 135122 199912 135174 199918
rect 135122 199854 135174 199860
rect 135226 199696 135254 200124
rect 135318 199918 135346 200124
rect 135410 199918 135438 200124
rect 135502 199918 135530 200124
rect 135306 199912 135358 199918
rect 135306 199854 135358 199860
rect 135398 199912 135450 199918
rect 135398 199854 135450 199860
rect 135490 199912 135542 199918
rect 135490 199854 135542 199860
rect 135352 199776 135404 199782
rect 135352 199718 135404 199724
rect 135042 199668 135116 199696
rect 134892 199640 134944 199646
rect 134892 199582 134944 199588
rect 134720 199396 134840 199424
rect 134720 191834 134748 199396
rect 134798 198792 134854 198801
rect 134798 198727 134854 198736
rect 134904 198734 134932 199582
rect 134984 199572 135036 199578
rect 134984 199514 135036 199520
rect 134996 199345 135024 199514
rect 134982 199336 135038 199345
rect 134982 199271 135038 199280
rect 135088 198801 135116 199668
rect 135180 199668 135254 199696
rect 135074 198792 135130 198801
rect 134812 193905 134840 198727
rect 134904 198706 135024 198734
rect 135074 198727 135130 198736
rect 134996 196518 135024 198706
rect 135074 197160 135130 197169
rect 135074 197095 135130 197104
rect 134984 196512 135036 196518
rect 134984 196454 135036 196460
rect 134984 196240 135036 196246
rect 134984 196182 135036 196188
rect 134892 196172 134944 196178
rect 134892 196114 134944 196120
rect 134798 193896 134854 193905
rect 134798 193831 134854 193840
rect 134720 191806 134840 191834
rect 134248 190936 134300 190942
rect 134248 190878 134300 190884
rect 134260 184482 134288 190878
rect 134248 184476 134300 184482
rect 134248 184418 134300 184424
rect 134156 178968 134208 178974
rect 134156 178910 134208 178916
rect 134064 178832 134116 178838
rect 134064 178774 134116 178780
rect 133788 176656 133840 176662
rect 133788 176598 133840 176604
rect 133800 175982 133828 176598
rect 133788 175976 133840 175982
rect 133788 175918 133840 175924
rect 133328 148640 133380 148646
rect 133328 148582 133380 148588
rect 133144 148504 133196 148510
rect 133144 148446 133196 148452
rect 132592 146056 132644 146062
rect 132592 145998 132644 146004
rect 131948 140480 132000 140486
rect 131948 140422 132000 140428
rect 132604 139890 132632 145998
rect 133696 141432 133748 141438
rect 133696 141374 133748 141380
rect 131132 139862 131376 139890
rect 131868 139862 132204 139890
rect 132604 139862 133032 139890
rect 133708 139534 133736 141374
rect 134352 140622 134380 190998
rect 134616 191004 134668 191010
rect 134616 190946 134668 190952
rect 134812 190890 134840 191806
rect 134444 190862 134840 190890
rect 134444 148578 134472 190862
rect 134522 190768 134578 190777
rect 134522 190703 134578 190712
rect 134536 180794 134564 190703
rect 134904 186314 134932 196114
rect 134996 195158 135024 196182
rect 134984 195152 135036 195158
rect 134984 195094 135036 195100
rect 135088 194070 135116 197095
rect 135076 194064 135128 194070
rect 135076 194006 135128 194012
rect 134628 186286 134932 186314
rect 134628 184618 134656 186286
rect 135180 185638 135208 199668
rect 135260 199572 135312 199578
rect 135260 199514 135312 199520
rect 135272 194041 135300 199514
rect 135364 197946 135392 199718
rect 135444 199708 135496 199714
rect 135594 199696 135622 200124
rect 135686 199918 135714 200124
rect 135778 199918 135806 200124
rect 135674 199912 135726 199918
rect 135674 199854 135726 199860
rect 135766 199912 135818 199918
rect 135766 199854 135818 199860
rect 135870 199764 135898 200124
rect 135962 199850 135990 200124
rect 136054 199918 136082 200124
rect 136042 199912 136094 199918
rect 136042 199854 136094 199860
rect 135950 199844 136002 199850
rect 135950 199786 136002 199792
rect 135824 199736 135898 199764
rect 135444 199650 135496 199656
rect 135548 199668 135622 199696
rect 135720 199708 135772 199714
rect 135352 197940 135404 197946
rect 135352 197882 135404 197888
rect 135456 196654 135484 199650
rect 135548 198393 135576 199668
rect 135720 199650 135772 199656
rect 135628 199572 135680 199578
rect 135628 199514 135680 199520
rect 135640 199322 135668 199514
rect 135732 199424 135760 199650
rect 135824 199578 135852 199736
rect 135996 199708 136048 199714
rect 136146 199696 136174 200124
rect 136238 199923 136266 200124
rect 136224 199914 136280 199923
rect 136224 199849 136280 199858
rect 136146 199668 136220 199696
rect 135996 199650 136048 199656
rect 135904 199640 135956 199646
rect 135904 199582 135956 199588
rect 135812 199572 135864 199578
rect 135812 199514 135864 199520
rect 135732 199396 135852 199424
rect 135640 199294 135760 199322
rect 135626 198792 135682 198801
rect 135626 198727 135682 198736
rect 135534 198384 135590 198393
rect 135534 198319 135590 198328
rect 135444 196648 135496 196654
rect 135444 196590 135496 196596
rect 135640 196178 135668 198727
rect 135628 196172 135680 196178
rect 135628 196114 135680 196120
rect 135258 194032 135314 194041
rect 135258 193967 135314 193976
rect 135732 193214 135760 199294
rect 135824 196246 135852 199396
rect 135812 196240 135864 196246
rect 135812 196182 135864 196188
rect 135812 196036 135864 196042
rect 135812 195978 135864 195984
rect 135640 193186 135760 193214
rect 135640 192438 135668 193186
rect 135628 192432 135680 192438
rect 135628 192374 135680 192380
rect 135720 191412 135772 191418
rect 135720 191354 135772 191360
rect 135536 191004 135588 191010
rect 135536 190946 135588 190952
rect 135548 185706 135576 190946
rect 135536 185700 135588 185706
rect 135536 185642 135588 185648
rect 135168 185632 135220 185638
rect 135168 185574 135220 185580
rect 134616 184612 134668 184618
rect 134616 184554 134668 184560
rect 134536 180766 134656 180794
rect 134522 178936 134578 178945
rect 134522 178871 134578 178880
rect 134536 178090 134564 178871
rect 134524 178084 134576 178090
rect 134524 178026 134576 178032
rect 134628 174758 134656 180766
rect 135168 178084 135220 178090
rect 135168 178026 135220 178032
rect 135180 177886 135208 178026
rect 135168 177880 135220 177886
rect 135168 177822 135220 177828
rect 135168 175228 135220 175234
rect 135168 175170 135220 175176
rect 135180 174758 135208 175170
rect 134616 174752 134668 174758
rect 134616 174694 134668 174700
rect 135168 174752 135220 174758
rect 135168 174694 135220 174700
rect 135732 148918 135760 191354
rect 135824 183258 135852 195978
rect 135812 183252 135864 183258
rect 135812 183194 135864 183200
rect 135916 174690 135944 199582
rect 136008 199345 136036 199650
rect 135994 199336 136050 199345
rect 135994 199271 136050 199280
rect 136192 198734 136220 199668
rect 136330 199628 136358 200124
rect 136422 199918 136450 200124
rect 136410 199912 136462 199918
rect 136410 199854 136462 199860
rect 136514 199764 136542 200124
rect 136606 199918 136634 200124
rect 136698 199918 136726 200124
rect 136790 199918 136818 200124
rect 136882 199918 136910 200124
rect 136594 199912 136646 199918
rect 136594 199854 136646 199860
rect 136686 199912 136738 199918
rect 136686 199854 136738 199860
rect 136778 199912 136830 199918
rect 136778 199854 136830 199860
rect 136870 199912 136922 199918
rect 136870 199854 136922 199860
rect 136640 199776 136692 199782
rect 136514 199736 136588 199764
rect 136456 199640 136508 199646
rect 136330 199600 136404 199628
rect 136376 198734 136404 199600
rect 136456 199582 136508 199588
rect 136100 198706 136220 198734
rect 136284 198706 136404 198734
rect 135996 196240 136048 196246
rect 135996 196182 136048 196188
rect 136008 193089 136036 196182
rect 135994 193080 136050 193089
rect 135994 193015 136050 193024
rect 136008 178770 136036 193015
rect 136100 191010 136128 198706
rect 136178 198520 136234 198529
rect 136178 198455 136234 198464
rect 136192 196246 136220 198455
rect 136180 196240 136232 196246
rect 136180 196182 136232 196188
rect 136180 196104 136232 196110
rect 136180 196046 136232 196052
rect 136192 191010 136220 196046
rect 136088 191004 136140 191010
rect 136088 190946 136140 190952
rect 136180 191004 136232 191010
rect 136180 190946 136232 190952
rect 136284 185570 136312 198706
rect 136468 197354 136496 199582
rect 136560 199345 136588 199736
rect 136974 199764 137002 200124
rect 136836 199736 137002 199764
rect 136836 199730 136864 199736
rect 136640 199718 136692 199724
rect 136546 199336 136602 199345
rect 136546 199271 136602 199280
rect 136468 197326 136588 197354
rect 136560 196042 136588 197326
rect 136548 196036 136600 196042
rect 136548 195978 136600 195984
rect 136362 195936 136418 195945
rect 136362 195871 136418 195880
rect 136376 191418 136404 195871
rect 136652 191834 136680 199718
rect 136744 199702 136864 199730
rect 136744 199345 136772 199702
rect 137066 199696 137094 200124
rect 137158 199918 137186 200124
rect 137146 199912 137198 199918
rect 137146 199854 137198 199860
rect 137066 199668 137140 199696
rect 136824 199572 136876 199578
rect 136824 199514 136876 199520
rect 136916 199572 136968 199578
rect 136916 199514 136968 199520
rect 137008 199572 137060 199578
rect 137008 199514 137060 199520
rect 136730 199336 136786 199345
rect 136730 199271 136786 199280
rect 136732 197736 136784 197742
rect 136732 197678 136784 197684
rect 136744 192982 136772 197678
rect 136836 196081 136864 199514
rect 136822 196072 136878 196081
rect 136928 196042 136956 199514
rect 137020 198762 137048 199514
rect 137008 198756 137060 198762
rect 137008 198698 137060 198704
rect 137006 198520 137062 198529
rect 137006 198455 137062 198464
rect 136822 196007 136878 196016
rect 136916 196036 136968 196042
rect 136916 195978 136968 195984
rect 136732 192976 136784 192982
rect 136732 192918 136784 192924
rect 136914 192808 136970 192817
rect 136914 192743 136970 192752
rect 136560 191806 136680 191834
rect 136364 191412 136416 191418
rect 136364 191354 136416 191360
rect 136560 191162 136588 191806
rect 136376 191134 136588 191162
rect 136376 186862 136404 191134
rect 136548 191004 136600 191010
rect 136548 190946 136600 190952
rect 136364 186856 136416 186862
rect 136364 186798 136416 186804
rect 136272 185564 136324 185570
rect 136272 185506 136324 185512
rect 136560 180742 136588 190946
rect 136824 190936 136876 190942
rect 136824 190878 136876 190884
rect 136548 180736 136600 180742
rect 136548 180678 136600 180684
rect 135996 178764 136048 178770
rect 135996 178706 136048 178712
rect 136836 177478 136864 190878
rect 136928 178906 136956 192743
rect 137020 181898 137048 198455
rect 137112 198286 137140 199668
rect 137250 199560 137278 200124
rect 137342 199923 137370 200124
rect 137328 199914 137384 199923
rect 137328 199849 137384 199858
rect 137434 199730 137462 200124
rect 137526 199850 137554 200124
rect 137618 199918 137646 200124
rect 137606 199912 137658 199918
rect 137606 199854 137658 199860
rect 137514 199844 137566 199850
rect 137514 199786 137566 199792
rect 137434 199702 137508 199730
rect 137376 199640 137428 199646
rect 137376 199582 137428 199588
rect 137204 199532 137278 199560
rect 137204 198393 137232 199532
rect 137388 199424 137416 199582
rect 137296 199396 137416 199424
rect 137296 199209 137324 199396
rect 137374 199336 137430 199345
rect 137374 199271 137430 199280
rect 137282 199200 137338 199209
rect 137282 199135 137338 199144
rect 137190 198384 137246 198393
rect 137190 198319 137246 198328
rect 137100 198280 137152 198286
rect 137100 198222 137152 198228
rect 137284 198212 137336 198218
rect 137284 198154 137336 198160
rect 137100 197600 137152 197606
rect 137100 197542 137152 197548
rect 137112 197402 137140 197542
rect 137296 197538 137324 198154
rect 137284 197532 137336 197538
rect 137284 197474 137336 197480
rect 137100 197396 137152 197402
rect 137100 197338 137152 197344
rect 137100 196036 137152 196042
rect 137100 195978 137152 195984
rect 137112 188494 137140 195978
rect 137388 191418 137416 199271
rect 137480 196654 137508 199702
rect 137560 199708 137612 199714
rect 137710 199696 137738 200124
rect 137802 199918 137830 200124
rect 137894 199923 137922 200124
rect 137790 199912 137842 199918
rect 137790 199854 137842 199860
rect 137880 199914 137936 199923
rect 137986 199918 138014 200124
rect 137880 199849 137936 199858
rect 137974 199912 138026 199918
rect 137974 199854 138026 199860
rect 137928 199776 137980 199782
rect 138078 199730 138106 200124
rect 138170 199782 138198 200124
rect 137928 199718 137980 199724
rect 137560 199650 137612 199656
rect 137664 199668 137738 199696
rect 137836 199708 137888 199714
rect 137468 196648 137520 196654
rect 137468 196590 137520 196596
rect 137468 196512 137520 196518
rect 137468 196454 137520 196460
rect 137376 191412 137428 191418
rect 137376 191354 137428 191360
rect 137480 191162 137508 196454
rect 137296 191134 137508 191162
rect 137192 191004 137244 191010
rect 137192 190946 137244 190952
rect 137100 188488 137152 188494
rect 137100 188430 137152 188436
rect 137008 181892 137060 181898
rect 137008 181834 137060 181840
rect 136916 178900 136968 178906
rect 136916 178842 136968 178848
rect 136824 177472 136876 177478
rect 136824 177414 136876 177420
rect 136546 176624 136602 176633
rect 136546 176559 136602 176568
rect 136560 175030 136588 176559
rect 136548 175024 136600 175030
rect 136548 174966 136600 174972
rect 135904 174684 135956 174690
rect 135904 174626 135956 174632
rect 136560 174622 136588 174966
rect 136548 174616 136600 174622
rect 136548 174558 136600 174564
rect 137204 151814 137232 190946
rect 137112 151786 137232 151814
rect 135720 148912 135772 148918
rect 135720 148854 135772 148860
rect 134432 148572 134484 148578
rect 134432 148514 134484 148520
rect 134800 146124 134852 146130
rect 134800 146066 134852 146072
rect 134812 143614 134840 146066
rect 135350 145888 135406 145897
rect 135350 145823 135406 145832
rect 134800 143608 134852 143614
rect 134800 143550 134852 143556
rect 134340 140616 134392 140622
rect 134340 140558 134392 140564
rect 134812 139890 134840 143550
rect 134688 139862 134840 139890
rect 135364 139890 135392 145823
rect 135996 143404 136048 143410
rect 135996 143346 136048 143352
rect 136008 139890 136036 143346
rect 137112 142934 137140 151786
rect 137192 145988 137244 145994
rect 137192 145930 137244 145936
rect 137100 142928 137152 142934
rect 137100 142870 137152 142876
rect 136822 142216 136878 142225
rect 136822 142151 136878 142160
rect 136836 139890 136864 142151
rect 137204 140162 137232 145930
rect 137296 140593 137324 191134
rect 137572 190942 137600 199650
rect 137664 198801 137692 199668
rect 137836 199650 137888 199656
rect 137744 199572 137796 199578
rect 137744 199514 137796 199520
rect 137650 198792 137706 198801
rect 137650 198727 137706 198736
rect 137652 198280 137704 198286
rect 137652 198222 137704 198228
rect 137560 190936 137612 190942
rect 137560 190878 137612 190884
rect 137376 190528 137428 190534
rect 137376 190470 137428 190476
rect 137388 148850 137416 190470
rect 137560 181960 137612 181966
rect 137560 181902 137612 181908
rect 137468 177676 137520 177682
rect 137468 177618 137520 177624
rect 137480 177478 137508 177618
rect 137468 177472 137520 177478
rect 137468 177414 137520 177420
rect 137376 148844 137428 148850
rect 137376 148786 137428 148792
rect 137480 144265 137508 177414
rect 137572 148442 137600 181902
rect 137664 175001 137692 198222
rect 137756 181694 137784 199514
rect 137848 199345 137876 199650
rect 137834 199336 137890 199345
rect 137834 199271 137890 199280
rect 137834 199200 137890 199209
rect 137834 199135 137890 199144
rect 137848 191010 137876 199135
rect 137940 194449 137968 199718
rect 138032 199702 138106 199730
rect 138158 199776 138210 199782
rect 138158 199718 138210 199724
rect 138032 198490 138060 199702
rect 138262 199628 138290 200124
rect 138354 199782 138382 200124
rect 138446 199923 138474 200124
rect 138432 199914 138488 199923
rect 138432 199849 138488 199858
rect 138342 199776 138394 199782
rect 138342 199718 138394 199724
rect 138538 199730 138566 200124
rect 138630 199918 138658 200124
rect 138722 199918 138750 200124
rect 138814 199923 138842 200124
rect 138618 199912 138670 199918
rect 138618 199854 138670 199860
rect 138710 199912 138762 199918
rect 138710 199854 138762 199860
rect 138800 199914 138856 199923
rect 138800 199849 138856 199858
rect 138906 199850 138934 200124
rect 138894 199844 138946 199850
rect 138894 199786 138946 199792
rect 138664 199776 138716 199782
rect 138538 199702 138612 199730
rect 138998 199730 139026 200124
rect 139090 199918 139118 200124
rect 139078 199912 139130 199918
rect 139078 199854 139130 199860
rect 139182 199850 139210 200124
rect 139274 199923 139302 200124
rect 139260 199914 139316 199923
rect 139170 199844 139222 199850
rect 139260 199849 139316 199858
rect 139366 199850 139394 200124
rect 139170 199786 139222 199792
rect 139354 199844 139406 199850
rect 139354 199786 139406 199792
rect 138664 199718 138716 199724
rect 138216 199600 138290 199628
rect 138110 199336 138166 199345
rect 138110 199271 138166 199280
rect 138020 198484 138072 198490
rect 138020 198426 138072 198432
rect 138124 198336 138152 199271
rect 138032 198308 138152 198336
rect 137926 194440 137982 194449
rect 137926 194375 137982 194384
rect 138032 193594 138060 198308
rect 138216 196110 138244 199600
rect 138388 199572 138440 199578
rect 138388 199514 138440 199520
rect 138400 198665 138428 199514
rect 138386 198656 138442 198665
rect 138386 198591 138442 198600
rect 138294 198248 138350 198257
rect 138294 198183 138350 198192
rect 138204 196104 138256 196110
rect 138204 196046 138256 196052
rect 138112 196036 138164 196042
rect 138112 195978 138164 195984
rect 138124 195838 138152 195978
rect 138112 195832 138164 195838
rect 138112 195774 138164 195780
rect 138020 193588 138072 193594
rect 138020 193530 138072 193536
rect 138308 192914 138336 198183
rect 138388 198008 138440 198014
rect 138388 197950 138440 197956
rect 138296 192908 138348 192914
rect 138296 192850 138348 192856
rect 138400 191834 138428 197950
rect 138584 196858 138612 199702
rect 138572 196852 138624 196858
rect 138572 196794 138624 196800
rect 138570 196752 138626 196761
rect 138570 196687 138626 196696
rect 138584 196654 138612 196687
rect 138572 196648 138624 196654
rect 138572 196590 138624 196596
rect 138478 196344 138534 196353
rect 138478 196279 138534 196288
rect 138216 191806 138428 191834
rect 137928 191412 137980 191418
rect 137928 191354 137980 191360
rect 138112 191412 138164 191418
rect 138112 191354 138164 191360
rect 137836 191004 137888 191010
rect 137836 190946 137888 190952
rect 137940 190534 137968 191354
rect 138124 191214 138152 191354
rect 138112 191208 138164 191214
rect 138112 191150 138164 191156
rect 137928 190528 137980 190534
rect 137928 190470 137980 190476
rect 138018 184920 138074 184929
rect 138018 184855 138074 184864
rect 137744 181688 137796 181694
rect 137744 181630 137796 181636
rect 138032 181393 138060 184855
rect 138018 181384 138074 181393
rect 138018 181319 138074 181328
rect 137650 174992 137706 175001
rect 137650 174927 137706 174936
rect 137664 174729 137692 174927
rect 137650 174720 137706 174729
rect 137650 174655 137706 174664
rect 138216 151230 138244 191806
rect 138296 191208 138348 191214
rect 138296 191150 138348 191156
rect 138308 184278 138336 191150
rect 138492 186314 138520 196279
rect 138584 189825 138612 196590
rect 138676 195945 138704 199718
rect 138952 199714 139026 199730
rect 138756 199708 138808 199714
rect 138756 199650 138808 199656
rect 138940 199708 139026 199714
rect 138992 199702 139026 199708
rect 139124 199708 139176 199714
rect 138940 199650 138992 199656
rect 139124 199650 139176 199656
rect 139216 199708 139268 199714
rect 139216 199650 139268 199656
rect 138768 198801 138796 199650
rect 138848 199640 138900 199646
rect 138848 199582 138900 199588
rect 139032 199640 139084 199646
rect 139032 199582 139084 199588
rect 138754 198792 138810 198801
rect 138754 198727 138810 198736
rect 138754 198112 138810 198121
rect 138754 198047 138810 198056
rect 138662 195936 138718 195945
rect 138662 195871 138718 195880
rect 138664 195288 138716 195294
rect 138664 195230 138716 195236
rect 138570 189816 138626 189825
rect 138570 189751 138626 189760
rect 138492 186286 138612 186314
rect 138296 184272 138348 184278
rect 138296 184214 138348 184220
rect 138204 151224 138256 151230
rect 138204 151166 138256 151172
rect 137560 148436 137612 148442
rect 137560 148378 137612 148384
rect 137466 144256 137522 144265
rect 137466 144191 137522 144200
rect 138480 143336 138532 143342
rect 138480 143278 138532 143284
rect 137282 140584 137338 140593
rect 137282 140519 137338 140528
rect 137204 140134 137600 140162
rect 137572 139890 137600 140134
rect 138492 139890 138520 143278
rect 138584 141506 138612 186286
rect 138676 147014 138704 195230
rect 138768 180470 138796 198047
rect 138860 191185 138888 199582
rect 138940 193588 138992 193594
rect 138940 193530 138992 193536
rect 138846 191176 138902 191185
rect 138846 191111 138902 191120
rect 138952 191026 138980 193530
rect 139044 191214 139072 199582
rect 139136 197849 139164 199650
rect 139122 197840 139178 197849
rect 139122 197775 139178 197784
rect 139228 197169 139256 199650
rect 139308 199640 139360 199646
rect 139458 199628 139486 200124
rect 139550 199923 139578 200124
rect 139536 199914 139592 199923
rect 139536 199849 139592 199858
rect 139642 199850 139670 200124
rect 139630 199844 139682 199850
rect 139630 199786 139682 199792
rect 139584 199708 139636 199714
rect 139584 199650 139636 199656
rect 139458 199600 139532 199628
rect 139308 199582 139360 199588
rect 139320 198014 139348 199582
rect 139308 198008 139360 198014
rect 139308 197950 139360 197956
rect 139504 197554 139532 199600
rect 139596 197878 139624 199650
rect 139734 199628 139762 200124
rect 139826 199730 139854 200124
rect 139918 199923 139946 200124
rect 139904 199914 139960 199923
rect 140010 199918 140038 200124
rect 139904 199849 139960 199858
rect 139998 199912 140050 199918
rect 139998 199854 140050 199860
rect 140102 199730 140130 200124
rect 140194 199850 140222 200124
rect 140286 199923 140314 200124
rect 140272 199914 140328 199923
rect 140182 199844 140234 199850
rect 140272 199849 140328 199858
rect 140182 199786 140234 199792
rect 139826 199702 139900 199730
rect 139688 199600 139762 199628
rect 139688 198218 139716 199600
rect 139676 198212 139728 198218
rect 139676 198154 139728 198160
rect 139872 198082 139900 199702
rect 139952 199708 140004 199714
rect 139952 199650 140004 199656
rect 140056 199702 140130 199730
rect 139860 198076 139912 198082
rect 139860 198018 139912 198024
rect 139964 198014 139992 199650
rect 140056 198218 140084 199702
rect 140378 199696 140406 200124
rect 140470 199850 140498 200124
rect 140458 199844 140510 199850
rect 140458 199786 140510 199792
rect 140562 199730 140590 200124
rect 140654 199923 140682 200124
rect 140640 199914 140696 199923
rect 140640 199849 140696 199858
rect 140516 199714 140590 199730
rect 140504 199708 140590 199714
rect 140378 199668 140452 199696
rect 140136 199640 140188 199646
rect 140136 199582 140188 199588
rect 140044 198212 140096 198218
rect 140044 198154 140096 198160
rect 140148 198064 140176 199582
rect 140320 199572 140372 199578
rect 140320 199514 140372 199520
rect 140228 199504 140280 199510
rect 140228 199446 140280 199452
rect 140240 198121 140268 199446
rect 140332 199209 140360 199514
rect 140318 199200 140374 199209
rect 140318 199135 140374 199144
rect 140320 198212 140372 198218
rect 140320 198154 140372 198160
rect 140056 198036 140176 198064
rect 140226 198112 140282 198121
rect 140226 198047 140282 198056
rect 139952 198008 140004 198014
rect 139952 197950 140004 197956
rect 139768 197940 139820 197946
rect 139768 197882 139820 197888
rect 139584 197872 139636 197878
rect 139584 197814 139636 197820
rect 139504 197526 139716 197554
rect 139582 197432 139638 197441
rect 139492 197396 139544 197402
rect 139582 197367 139638 197376
rect 139492 197338 139544 197344
rect 139308 197328 139360 197334
rect 139308 197270 139360 197276
rect 139214 197160 139270 197169
rect 139214 197095 139270 197104
rect 139320 196382 139348 197270
rect 139308 196376 139360 196382
rect 139308 196318 139360 196324
rect 139504 192846 139532 197338
rect 139492 192840 139544 192846
rect 139492 192782 139544 192788
rect 139032 191208 139084 191214
rect 139032 191150 139084 191156
rect 138952 190998 139072 191026
rect 138938 189000 138994 189009
rect 138938 188935 138994 188944
rect 138952 188737 138980 188935
rect 138938 188728 138994 188737
rect 138938 188663 138994 188672
rect 138952 181626 138980 188663
rect 138940 181620 138992 181626
rect 138940 181562 138992 181568
rect 138756 180464 138808 180470
rect 138756 180406 138808 180412
rect 138664 147008 138716 147014
rect 138664 146950 138716 146956
rect 139044 146946 139072 190998
rect 139490 190224 139546 190233
rect 139490 190159 139546 190168
rect 139504 189825 139532 190159
rect 139490 189816 139546 189825
rect 139490 189751 139546 189760
rect 139596 182034 139624 197367
rect 139688 182850 139716 197526
rect 139780 184550 139808 197882
rect 139952 197872 140004 197878
rect 139952 197814 140004 197820
rect 139860 194608 139912 194614
rect 139860 194550 139912 194556
rect 139872 192574 139900 194550
rect 139964 194410 139992 197814
rect 140056 197674 140084 198036
rect 140332 197996 140360 198154
rect 140148 197968 140360 197996
rect 140044 197668 140096 197674
rect 140044 197610 140096 197616
rect 140044 196376 140096 196382
rect 140044 196318 140096 196324
rect 139952 194404 140004 194410
rect 139952 194346 140004 194352
rect 139964 194138 139992 194346
rect 139952 194132 140004 194138
rect 139952 194074 140004 194080
rect 139860 192568 139912 192574
rect 139860 192510 139912 192516
rect 139768 184544 139820 184550
rect 139768 184486 139820 184492
rect 139676 182844 139728 182850
rect 139676 182786 139728 182792
rect 139584 182028 139636 182034
rect 139584 181970 139636 181976
rect 140056 180606 140084 196318
rect 140148 191214 140176 197968
rect 140320 197872 140372 197878
rect 140320 197814 140372 197820
rect 140226 197568 140282 197577
rect 140226 197503 140282 197512
rect 140136 191208 140188 191214
rect 140136 191150 140188 191156
rect 140134 190224 140190 190233
rect 140134 190159 140190 190168
rect 140044 180600 140096 180606
rect 140044 180542 140096 180548
rect 140148 177750 140176 190159
rect 140240 181966 140268 197503
rect 140332 197402 140360 197814
rect 140320 197396 140372 197402
rect 140320 197338 140372 197344
rect 140228 181960 140280 181966
rect 140228 181902 140280 181908
rect 140136 177744 140188 177750
rect 140136 177686 140188 177692
rect 140424 151094 140452 199668
rect 140556 199702 140590 199708
rect 140746 199696 140774 200124
rect 140838 199918 140866 200124
rect 140826 199912 140878 199918
rect 140826 199854 140878 199860
rect 140930 199764 140958 200124
rect 140884 199736 140958 199764
rect 140746 199668 140820 199696
rect 140504 199650 140556 199656
rect 140688 199572 140740 199578
rect 140688 199514 140740 199520
rect 140596 199504 140648 199510
rect 140596 199446 140648 199452
rect 140504 199300 140556 199306
rect 140504 199242 140556 199248
rect 140516 199209 140544 199242
rect 140502 199200 140558 199209
rect 140502 199135 140558 199144
rect 140608 195974 140636 199446
rect 140700 198082 140728 199514
rect 140688 198076 140740 198082
rect 140688 198018 140740 198024
rect 140792 197946 140820 199668
rect 140884 198354 140912 199736
rect 141022 199696 141050 200124
rect 141114 199918 141142 200124
rect 141102 199912 141154 199918
rect 141102 199854 141154 199860
rect 141206 199730 141234 200124
rect 140976 199668 141050 199696
rect 141114 199702 141234 199730
rect 140976 198558 141004 199668
rect 141114 199628 141142 199702
rect 141298 199628 141326 200124
rect 141390 199918 141418 200124
rect 141378 199912 141430 199918
rect 141378 199854 141430 199860
rect 141482 199850 141510 200124
rect 141470 199844 141522 199850
rect 141470 199786 141522 199792
rect 141574 199696 141602 200124
rect 141114 199600 141188 199628
rect 140964 198552 141016 198558
rect 140964 198494 141016 198500
rect 140872 198348 140924 198354
rect 140872 198290 140924 198296
rect 140964 198280 141016 198286
rect 140964 198222 141016 198228
rect 140780 197940 140832 197946
rect 140780 197882 140832 197888
rect 140780 197804 140832 197810
rect 140780 197746 140832 197752
rect 140688 197668 140740 197674
rect 140688 197610 140740 197616
rect 140516 195946 140636 195974
rect 140516 184414 140544 195946
rect 140700 193934 140728 197610
rect 140792 195294 140820 197746
rect 140780 195288 140832 195294
rect 140780 195230 140832 195236
rect 140688 193928 140740 193934
rect 140688 193870 140740 193876
rect 140688 191208 140740 191214
rect 140688 191150 140740 191156
rect 140504 184408 140556 184414
rect 140504 184350 140556 184356
rect 140700 151162 140728 191150
rect 140976 182918 141004 198222
rect 141056 198008 141108 198014
rect 141056 197950 141108 197956
rect 141068 186314 141096 197950
rect 141160 197810 141188 199600
rect 141252 199600 141326 199628
rect 141528 199668 141602 199696
rect 141252 198422 141280 199600
rect 141424 199504 141476 199510
rect 141424 199446 141476 199452
rect 141240 198416 141292 198422
rect 141240 198358 141292 198364
rect 141148 197804 141200 197810
rect 141148 197746 141200 197752
rect 141332 196784 141384 196790
rect 141332 196726 141384 196732
rect 141344 193050 141372 196726
rect 141436 195673 141464 199446
rect 141528 197810 141556 199668
rect 141666 199594 141694 200124
rect 141758 199850 141786 200124
rect 141746 199844 141798 199850
rect 141746 199786 141798 199792
rect 141850 199594 141878 200124
rect 141942 199850 141970 200124
rect 142034 199918 142062 200124
rect 142022 199912 142074 199918
rect 142022 199854 142074 199860
rect 141930 199844 141982 199850
rect 141930 199786 141982 199792
rect 142126 199764 142154 200124
rect 142218 199923 142246 200124
rect 142204 199914 142260 199923
rect 142204 199849 142260 199858
rect 142080 199736 142154 199764
rect 142080 199730 142108 199736
rect 142310 199730 142338 200124
rect 141620 199566 141694 199594
rect 141804 199566 141878 199594
rect 141988 199702 142108 199730
rect 142264 199702 142338 199730
rect 142402 199730 142430 200124
rect 142494 199923 142522 200124
rect 142480 199914 142536 199923
rect 142586 199918 142614 200124
rect 142678 199918 142706 200124
rect 142770 199918 142798 200124
rect 142862 199923 142890 200124
rect 142480 199849 142536 199858
rect 142574 199912 142626 199918
rect 142574 199854 142626 199860
rect 142666 199912 142718 199918
rect 142666 199854 142718 199860
rect 142758 199912 142810 199918
rect 142758 199854 142810 199860
rect 142848 199914 142904 199923
rect 142848 199849 142904 199858
rect 142954 199850 142982 200124
rect 142942 199844 142994 199850
rect 142942 199786 142994 199792
rect 143046 199730 143074 200124
rect 143138 199782 143166 200124
rect 142402 199702 142476 199730
rect 143000 199714 143074 199730
rect 143126 199776 143178 199782
rect 143126 199718 143178 199724
rect 143230 199730 143258 200124
rect 143322 199918 143350 200124
rect 143310 199912 143362 199918
rect 143310 199854 143362 199860
rect 141516 197804 141568 197810
rect 141516 197746 141568 197752
rect 141516 197328 141568 197334
rect 141516 197270 141568 197276
rect 141422 195664 141478 195673
rect 141422 195599 141478 195608
rect 141528 194478 141556 197270
rect 141516 194472 141568 194478
rect 141516 194414 141568 194420
rect 141332 193044 141384 193050
rect 141332 192986 141384 192992
rect 141068 186286 141188 186314
rect 140964 182912 141016 182918
rect 140964 182854 141016 182860
rect 141160 177818 141188 186286
rect 141620 180794 141648 199566
rect 141700 199504 141752 199510
rect 141700 199446 141752 199452
rect 141712 198801 141740 199446
rect 141698 198792 141754 198801
rect 141698 198727 141754 198736
rect 141700 198076 141752 198082
rect 141700 198018 141752 198024
rect 141712 195974 141740 198018
rect 141804 196382 141832 199566
rect 141884 199504 141936 199510
rect 141884 199446 141936 199452
rect 141896 198286 141924 199446
rect 141884 198280 141936 198286
rect 141884 198222 141936 198228
rect 141884 198144 141936 198150
rect 141884 198086 141936 198092
rect 141896 197062 141924 198086
rect 141988 197305 142016 199702
rect 142160 199640 142212 199646
rect 142160 199582 142212 199588
rect 142172 199034 142200 199582
rect 142160 199028 142212 199034
rect 142160 198970 142212 198976
rect 142264 198966 142292 199702
rect 142344 199640 142396 199646
rect 142344 199582 142396 199588
rect 142252 198960 142304 198966
rect 142252 198902 142304 198908
rect 142068 198824 142120 198830
rect 142068 198766 142120 198772
rect 142080 198014 142108 198766
rect 142252 198552 142304 198558
rect 142250 198520 142252 198529
rect 142304 198520 142306 198529
rect 142250 198455 142306 198464
rect 142356 198336 142384 199582
rect 142264 198308 142384 198336
rect 142068 198008 142120 198014
rect 142068 197950 142120 197956
rect 142068 197804 142120 197810
rect 142068 197746 142120 197752
rect 141974 197296 142030 197305
rect 141974 197231 142030 197240
rect 141884 197056 141936 197062
rect 141884 196998 141936 197004
rect 141792 196376 141844 196382
rect 141792 196318 141844 196324
rect 142080 195974 142108 197746
rect 142264 197674 142292 198308
rect 142344 198212 142396 198218
rect 142344 198154 142396 198160
rect 142252 197668 142304 197674
rect 142252 197610 142304 197616
rect 141712 195946 141924 195974
rect 141896 182102 141924 195946
rect 141988 195946 142108 195974
rect 141988 195838 142016 195946
rect 142356 195906 142384 198154
rect 142344 195900 142396 195906
rect 142344 195842 142396 195848
rect 141976 195832 142028 195838
rect 141976 195774 142028 195780
rect 141988 194177 142016 195774
rect 142448 194614 142476 199702
rect 142528 199708 142580 199714
rect 142528 199650 142580 199656
rect 142988 199708 143074 199714
rect 143040 199702 143074 199708
rect 143230 199702 143350 199730
rect 143414 199714 143442 200124
rect 143506 199782 143534 200124
rect 143598 199918 143626 200124
rect 143586 199912 143638 199918
rect 143586 199854 143638 199860
rect 143494 199776 143546 199782
rect 143494 199718 143546 199724
rect 142988 199650 143040 199656
rect 142540 197305 142568 199650
rect 142804 199640 142856 199646
rect 142804 199582 142856 199588
rect 143080 199640 143132 199646
rect 143080 199582 143132 199588
rect 143172 199640 143224 199646
rect 143172 199582 143224 199588
rect 143322 199594 143350 199702
rect 143402 199708 143454 199714
rect 143402 199650 143454 199656
rect 143540 199640 143592 199646
rect 142620 199572 142672 199578
rect 142620 199514 142672 199520
rect 142712 199572 142764 199578
rect 142712 199514 142764 199520
rect 142632 198665 142660 199514
rect 142618 198656 142674 198665
rect 142618 198591 142674 198600
rect 142724 198200 142752 199514
rect 142632 198172 142752 198200
rect 142526 197296 142582 197305
rect 142526 197231 142582 197240
rect 142540 196382 142568 197231
rect 142528 196376 142580 196382
rect 142528 196318 142580 196324
rect 142436 194608 142488 194614
rect 142436 194550 142488 194556
rect 142632 194478 142660 198172
rect 142710 198112 142766 198121
rect 142710 198047 142766 198056
rect 142620 194472 142672 194478
rect 142620 194414 142672 194420
rect 141974 194168 142030 194177
rect 141974 194103 142030 194112
rect 142632 189689 142660 194414
rect 142618 189680 142674 189689
rect 142618 189615 142674 189624
rect 142724 187406 142752 198047
rect 142816 196790 142844 199582
rect 142896 198348 142948 198354
rect 142896 198290 142948 198296
rect 142804 196784 142856 196790
rect 142804 196726 142856 196732
rect 142804 195628 142856 195634
rect 142804 195570 142856 195576
rect 142816 195022 142844 195570
rect 142804 195016 142856 195022
rect 142804 194958 142856 194964
rect 142804 191208 142856 191214
rect 142804 191150 142856 191156
rect 142712 187400 142764 187406
rect 142712 187342 142764 187348
rect 141884 182096 141936 182102
rect 141884 182038 141936 182044
rect 141344 180766 141648 180794
rect 140780 177812 140832 177818
rect 140780 177754 140832 177760
rect 141148 177812 141200 177818
rect 141148 177754 141200 177760
rect 140792 177342 140820 177754
rect 141344 177342 141372 180766
rect 140780 177336 140832 177342
rect 140780 177278 140832 177284
rect 141332 177336 141384 177342
rect 141332 177278 141384 177284
rect 142160 177336 142212 177342
rect 142160 177278 142212 177284
rect 140778 176624 140834 176633
rect 140778 176559 140834 176568
rect 140792 175098 140820 176559
rect 140870 175264 140926 175273
rect 140870 175199 140926 175208
rect 140884 175166 140912 175199
rect 140872 175160 140924 175166
rect 140872 175102 140924 175108
rect 140780 175092 140832 175098
rect 140780 175034 140832 175040
rect 140792 174554 140820 175034
rect 140780 174548 140832 174554
rect 140780 174490 140832 174496
rect 140884 173942 140912 175102
rect 140872 173936 140924 173942
rect 140872 173878 140924 173884
rect 140688 151156 140740 151162
rect 140688 151098 140740 151104
rect 140412 151088 140464 151094
rect 140412 151030 140464 151036
rect 139032 146940 139084 146946
rect 139032 146882 139084 146888
rect 139400 145920 139452 145926
rect 139400 145862 139452 145868
rect 138572 141500 138624 141506
rect 138572 141442 138624 141448
rect 139412 139890 139440 145862
rect 139768 144832 139820 144838
rect 139768 144774 139820 144780
rect 139780 143750 139808 144774
rect 141792 144764 141844 144770
rect 141792 144706 141844 144712
rect 139768 143744 139820 143750
rect 139768 143686 139820 143692
rect 140412 143744 140464 143750
rect 140412 143686 140464 143692
rect 135364 139862 135516 139890
rect 136008 139862 136344 139890
rect 136836 139862 137172 139890
rect 137572 139862 138000 139890
rect 138492 139862 138828 139890
rect 139412 139862 139656 139890
rect 140424 139754 140452 143686
rect 141240 143200 141292 143206
rect 141240 143142 141292 143148
rect 141252 141438 141280 143142
rect 141240 141432 141292 141438
rect 141240 141374 141292 141380
rect 141252 139890 141280 141374
rect 141804 139890 141832 144706
rect 142172 144634 142200 177278
rect 142160 144628 142212 144634
rect 142160 144570 142212 144576
rect 142620 143064 142672 143070
rect 142620 143006 142672 143012
rect 142632 139890 142660 143006
rect 142816 140282 142844 191150
rect 142908 183326 142936 198290
rect 142988 197396 143040 197402
rect 142988 197338 143040 197344
rect 143000 191214 143028 197338
rect 143092 196489 143120 199582
rect 143078 196480 143134 196489
rect 143078 196415 143134 196424
rect 143080 196376 143132 196382
rect 143080 196318 143132 196324
rect 142988 191208 143040 191214
rect 142988 191150 143040 191156
rect 143092 186969 143120 196318
rect 143184 191350 143212 199582
rect 143322 199566 143488 199594
rect 143540 199582 143592 199588
rect 143264 199504 143316 199510
rect 143264 199446 143316 199452
rect 143356 199504 143408 199510
rect 143356 199446 143408 199452
rect 143276 195226 143304 199446
rect 143264 195220 143316 195226
rect 143264 195162 143316 195168
rect 143172 191344 143224 191350
rect 143172 191286 143224 191292
rect 143368 187338 143396 199446
rect 143460 198218 143488 199566
rect 143448 198212 143500 198218
rect 143448 198154 143500 198160
rect 143552 198064 143580 199582
rect 143690 199492 143718 200124
rect 143782 199850 143810 200124
rect 143770 199844 143822 199850
rect 143770 199786 143822 199792
rect 143874 199782 143902 200124
rect 143862 199776 143914 199782
rect 143862 199718 143914 199724
rect 143966 199696 143994 200124
rect 144058 199764 144086 200124
rect 144150 199918 144178 200124
rect 144138 199912 144190 199918
rect 144138 199854 144190 199860
rect 144058 199736 144132 199764
rect 143966 199668 144040 199696
rect 143908 199572 143960 199578
rect 143908 199514 143960 199520
rect 143816 199504 143868 199510
rect 143690 199464 143764 199492
rect 143460 198036 143580 198064
rect 143356 187332 143408 187338
rect 143356 187274 143408 187280
rect 143078 186960 143134 186969
rect 143078 186895 143134 186904
rect 143460 186182 143488 198036
rect 143736 187134 143764 199464
rect 143816 199446 143868 199452
rect 143828 196110 143856 199446
rect 143920 198354 143948 199514
rect 144012 199170 144040 199668
rect 144104 199306 144132 199736
rect 144242 199730 144270 200124
rect 144334 199923 144362 200124
rect 144320 199914 144376 199923
rect 144426 199918 144454 200124
rect 144320 199849 144376 199858
rect 144414 199912 144466 199918
rect 144414 199854 144466 199860
rect 144196 199702 144270 199730
rect 144368 199776 144420 199782
rect 144518 199764 144546 200124
rect 144610 199923 144638 200124
rect 144596 199914 144652 199923
rect 144596 199849 144652 199858
rect 144420 199736 144546 199764
rect 144368 199718 144420 199724
rect 144092 199300 144144 199306
rect 144092 199242 144144 199248
rect 144000 199164 144052 199170
rect 144000 199106 144052 199112
rect 143908 198348 143960 198354
rect 143908 198290 143960 198296
rect 143906 198248 143962 198257
rect 143906 198183 143962 198192
rect 143816 196104 143868 196110
rect 143816 196046 143868 196052
rect 143920 191418 143948 198183
rect 144104 196518 144132 199242
rect 144196 197470 144224 199702
rect 144702 199696 144730 200124
rect 144794 199850 144822 200124
rect 144886 199918 144914 200124
rect 144978 199918 145006 200124
rect 145070 199923 145098 200124
rect 144874 199912 144926 199918
rect 144874 199854 144926 199860
rect 144966 199912 145018 199918
rect 144966 199854 145018 199860
rect 145056 199914 145112 199923
rect 145162 199918 145190 200124
rect 145254 199918 145282 200124
rect 145346 199918 145374 200124
rect 145438 199918 145466 200124
rect 145530 199918 145558 200124
rect 145622 199923 145650 200124
rect 144782 199844 144834 199850
rect 145056 199849 145112 199858
rect 145150 199912 145202 199918
rect 145150 199854 145202 199860
rect 145242 199912 145294 199918
rect 145242 199854 145294 199860
rect 145334 199912 145386 199918
rect 145334 199854 145386 199860
rect 145426 199912 145478 199918
rect 145426 199854 145478 199860
rect 145518 199912 145570 199918
rect 145518 199854 145570 199860
rect 145608 199914 145664 199923
rect 145714 199918 145742 200124
rect 145608 199849 145664 199858
rect 145702 199912 145754 199918
rect 145702 199854 145754 199860
rect 144782 199786 144834 199792
rect 145196 199776 145248 199782
rect 145806 199764 145834 200124
rect 145898 199918 145926 200124
rect 145990 199918 146018 200124
rect 146082 199918 146110 200124
rect 146174 199923 146202 200124
rect 145886 199912 145938 199918
rect 145886 199854 145938 199860
rect 145978 199912 146030 199918
rect 145978 199854 146030 199860
rect 146070 199912 146122 199918
rect 146070 199854 146122 199860
rect 146160 199914 146216 199923
rect 146266 199918 146294 200124
rect 146358 199918 146386 200124
rect 146450 199918 146478 200124
rect 146542 199918 146570 200124
rect 146160 199849 146216 199858
rect 146254 199912 146306 199918
rect 146254 199854 146306 199860
rect 146346 199912 146398 199918
rect 146346 199854 146398 199860
rect 146438 199912 146490 199918
rect 146438 199854 146490 199860
rect 146530 199912 146582 199918
rect 146530 199854 146582 199860
rect 145196 199718 145248 199724
rect 145760 199736 145834 199764
rect 146208 199776 146260 199782
rect 144828 199708 144880 199714
rect 144702 199668 144776 199696
rect 144276 199640 144328 199646
rect 144276 199582 144328 199588
rect 144288 198665 144316 199582
rect 144368 199572 144420 199578
rect 144368 199514 144420 199520
rect 144460 199572 144512 199578
rect 144460 199514 144512 199520
rect 144380 199209 144408 199514
rect 144366 199200 144422 199209
rect 144366 199135 144422 199144
rect 144366 198792 144422 198801
rect 144366 198727 144422 198736
rect 144274 198656 144330 198665
rect 144274 198591 144330 198600
rect 144276 197940 144328 197946
rect 144276 197882 144328 197888
rect 144184 197464 144236 197470
rect 144184 197406 144236 197412
rect 144288 197130 144316 197882
rect 144276 197124 144328 197130
rect 144276 197066 144328 197072
rect 144092 196512 144144 196518
rect 144092 196454 144144 196460
rect 144184 193588 144236 193594
rect 144184 193530 144236 193536
rect 143908 191412 143960 191418
rect 143908 191354 143960 191360
rect 143724 187128 143776 187134
rect 143724 187070 143776 187076
rect 143448 186176 143500 186182
rect 143448 186118 143500 186124
rect 142896 183320 142948 183326
rect 142896 183262 142948 183268
rect 143632 143268 143684 143274
rect 143632 143210 143684 143216
rect 143540 142248 143592 142254
rect 143540 142190 143592 142196
rect 143552 142050 143580 142190
rect 143540 142044 143592 142050
rect 143540 141986 143592 141992
rect 142804 140276 142856 140282
rect 142804 140218 142856 140224
rect 143644 139890 143672 143210
rect 144196 140418 144224 193530
rect 144380 189990 144408 198727
rect 144368 189984 144420 189990
rect 144368 189926 144420 189932
rect 144472 189825 144500 199514
rect 144748 198937 144776 199668
rect 144828 199650 144880 199656
rect 144920 199708 144972 199714
rect 144920 199650 144972 199656
rect 144734 198928 144790 198937
rect 144734 198863 144790 198872
rect 144550 198112 144606 198121
rect 144550 198047 144606 198056
rect 144736 198076 144788 198082
rect 144564 189854 144592 198047
rect 144736 198018 144788 198024
rect 144644 197464 144696 197470
rect 144644 197406 144696 197412
rect 144552 189848 144604 189854
rect 144458 189816 144514 189825
rect 144552 189790 144604 189796
rect 144458 189751 144514 189760
rect 144656 188426 144684 197406
rect 144644 188420 144696 188426
rect 144644 188362 144696 188368
rect 144748 186314 144776 198018
rect 144840 197334 144868 199650
rect 144828 197328 144880 197334
rect 144828 197270 144880 197276
rect 144828 196240 144880 196246
rect 144828 196182 144880 196188
rect 144840 192642 144868 196182
rect 144932 193594 144960 199650
rect 145012 199572 145064 199578
rect 145012 199514 145064 199520
rect 145024 198082 145052 199514
rect 145102 198520 145158 198529
rect 145102 198455 145158 198464
rect 145012 198076 145064 198082
rect 145012 198018 145064 198024
rect 145012 197668 145064 197674
rect 145012 197610 145064 197616
rect 144920 193588 144972 193594
rect 144920 193530 144972 193536
rect 144828 192636 144880 192642
rect 144828 192578 144880 192584
rect 145024 191826 145052 197610
rect 145116 193118 145144 198455
rect 145208 197402 145236 199718
rect 145564 199708 145616 199714
rect 145484 199668 145564 199696
rect 145380 199640 145432 199646
rect 145380 199582 145432 199588
rect 145288 199572 145340 199578
rect 145288 199514 145340 199520
rect 145300 197946 145328 199514
rect 145288 197940 145340 197946
rect 145288 197882 145340 197888
rect 145286 197840 145342 197849
rect 145286 197775 145288 197784
rect 145340 197775 145342 197784
rect 145288 197746 145340 197752
rect 145196 197396 145248 197402
rect 145196 197338 145248 197344
rect 145392 196586 145420 199582
rect 145380 196580 145432 196586
rect 145380 196522 145432 196528
rect 145104 193112 145156 193118
rect 145104 193054 145156 193060
rect 145012 191820 145064 191826
rect 145012 191762 145064 191768
rect 144918 187504 144974 187513
rect 144918 187439 144974 187448
rect 144932 187202 144960 187439
rect 144920 187196 144972 187202
rect 144920 187138 144972 187144
rect 145116 187105 145144 193054
rect 145484 192370 145512 199668
rect 145564 199650 145616 199656
rect 145656 199708 145708 199714
rect 145656 199650 145708 199656
rect 145668 199288 145696 199650
rect 145576 199260 145696 199288
rect 145576 196246 145604 199260
rect 145656 199164 145708 199170
rect 145656 199106 145708 199112
rect 145668 197062 145696 199106
rect 145656 197056 145708 197062
rect 145656 196998 145708 197004
rect 145760 196704 145788 199736
rect 146208 199718 146260 199724
rect 146300 199776 146352 199782
rect 146300 199718 146352 199724
rect 146392 199776 146444 199782
rect 146634 199764 146662 200124
rect 146392 199718 146444 199724
rect 146588 199736 146662 199764
rect 146024 199708 146076 199714
rect 146024 199650 146076 199656
rect 145840 199640 145892 199646
rect 145840 199582 145892 199588
rect 145932 199640 145984 199646
rect 145932 199582 145984 199588
rect 145668 196676 145788 196704
rect 145564 196240 145616 196246
rect 145564 196182 145616 196188
rect 145564 196036 145616 196042
rect 145564 195978 145616 195984
rect 145472 192364 145524 192370
rect 145472 192306 145524 192312
rect 145472 191208 145524 191214
rect 145472 191150 145524 191156
rect 145102 187096 145158 187105
rect 145102 187031 145158 187040
rect 144472 186286 144776 186314
rect 144472 184346 144500 186286
rect 145378 186280 145434 186289
rect 145378 186215 145434 186224
rect 145392 184890 145420 186215
rect 145380 184884 145432 184890
rect 145380 184826 145432 184832
rect 144460 184340 144512 184346
rect 144460 184282 144512 184288
rect 144920 145852 144972 145858
rect 144920 145794 144972 145800
rect 144932 142322 144960 145794
rect 144920 142316 144972 142322
rect 144920 142258 144972 142264
rect 145380 142316 145432 142322
rect 145380 142258 145432 142264
rect 144276 141840 144328 141846
rect 144276 141782 144328 141788
rect 144184 140412 144236 140418
rect 144184 140354 144236 140360
rect 144288 139890 144316 141782
rect 145392 139890 145420 142258
rect 145484 140214 145512 191150
rect 145576 187678 145604 195978
rect 145564 187672 145616 187678
rect 145564 187614 145616 187620
rect 145668 187513 145696 196676
rect 145748 196580 145800 196586
rect 145748 196522 145800 196528
rect 145654 187504 145710 187513
rect 145654 187439 145710 187448
rect 145760 186289 145788 196522
rect 145852 189922 145880 199582
rect 145944 195537 145972 199582
rect 145930 195528 145986 195537
rect 145930 195463 145986 195472
rect 146036 191214 146064 199650
rect 146114 198112 146170 198121
rect 146114 198047 146170 198056
rect 146128 197878 146156 198047
rect 146116 197872 146168 197878
rect 146116 197814 146168 197820
rect 146220 197130 146248 199718
rect 146208 197124 146260 197130
rect 146208 197066 146260 197072
rect 146312 196042 146340 199718
rect 146404 199209 146432 199718
rect 146484 199572 146536 199578
rect 146484 199514 146536 199520
rect 146390 199200 146446 199209
rect 146390 199135 146446 199144
rect 146392 198824 146444 198830
rect 146392 198766 146444 198772
rect 146404 197674 146432 198766
rect 146392 197668 146444 197674
rect 146392 197610 146444 197616
rect 146392 197464 146444 197470
rect 146392 197406 146444 197412
rect 146300 196036 146352 196042
rect 146300 195978 146352 195984
rect 146024 191208 146076 191214
rect 146024 191150 146076 191156
rect 145840 189916 145892 189922
rect 145840 189858 145892 189864
rect 145562 186280 145618 186289
rect 145562 186215 145618 186224
rect 145746 186280 145802 186289
rect 145746 186215 145802 186224
rect 145576 185609 145604 186215
rect 145562 185600 145618 185609
rect 145562 185535 145618 185544
rect 146404 144498 146432 197406
rect 146496 195401 146524 199514
rect 146588 197538 146616 199736
rect 146726 199696 146754 200124
rect 146818 199923 146846 200124
rect 146804 199914 146860 199923
rect 146804 199849 146860 199858
rect 146680 199668 146754 199696
rect 146910 199696 146938 200124
rect 147002 199764 147030 200124
rect 147094 199918 147122 200124
rect 147082 199912 147134 199918
rect 147082 199854 147134 199860
rect 147186 199764 147214 200124
rect 147002 199736 147076 199764
rect 146910 199668 146984 199696
rect 146576 197532 146628 197538
rect 146576 197474 146628 197480
rect 146482 195392 146538 195401
rect 146482 195327 146538 195336
rect 146484 191208 146536 191214
rect 146484 191150 146536 191156
rect 146496 145790 146524 191150
rect 146576 191072 146628 191078
rect 146576 191014 146628 191020
rect 146588 163538 146616 191014
rect 146680 181830 146708 199668
rect 146760 199572 146812 199578
rect 146760 199514 146812 199520
rect 146772 192642 146800 199514
rect 146852 199504 146904 199510
rect 146852 199446 146904 199452
rect 146864 198830 146892 199446
rect 146852 198824 146904 198830
rect 146852 198766 146904 198772
rect 146956 198734 146984 199668
rect 146864 198706 146984 198734
rect 146760 192636 146812 192642
rect 146760 192578 146812 192584
rect 146668 181824 146720 181830
rect 146668 181766 146720 181772
rect 146576 163532 146628 163538
rect 146576 163474 146628 163480
rect 146772 151814 146800 192578
rect 146588 151786 146800 151814
rect 146484 145784 146536 145790
rect 146484 145726 146536 145732
rect 146588 145654 146616 151786
rect 146864 147674 146892 198706
rect 147048 198558 147076 199736
rect 147140 199736 147214 199764
rect 147036 198552 147088 198558
rect 147036 198494 147088 198500
rect 146944 196648 146996 196654
rect 146944 196590 146996 196596
rect 146680 147646 146892 147674
rect 146576 145648 146628 145654
rect 146576 145590 146628 145596
rect 146392 144492 146444 144498
rect 146392 144434 146444 144440
rect 146680 143426 146708 147646
rect 146956 143426 146984 196590
rect 147140 191214 147168 199736
rect 147278 199696 147306 200124
rect 147232 199668 147306 199696
rect 147232 191834 147260 199668
rect 147370 199628 147398 200124
rect 147462 199764 147490 200124
rect 147554 199918 147582 200124
rect 147542 199912 147594 199918
rect 147542 199854 147594 199860
rect 147462 199736 147536 199764
rect 147324 199600 147398 199628
rect 147324 193186 147352 199600
rect 147404 199504 147456 199510
rect 147404 199446 147456 199452
rect 147416 199209 147444 199446
rect 147402 199200 147458 199209
rect 147402 199135 147458 199144
rect 147508 199073 147536 199736
rect 147646 199730 147674 200124
rect 147738 199918 147766 200124
rect 147830 199923 147858 200124
rect 147726 199912 147778 199918
rect 147726 199854 147778 199860
rect 147816 199914 147872 199923
rect 147922 199918 147950 200124
rect 148014 199918 148042 200124
rect 147816 199849 147872 199858
rect 147910 199912 147962 199918
rect 147910 199854 147962 199860
rect 148002 199912 148054 199918
rect 148002 199854 148054 199860
rect 147600 199702 147674 199730
rect 147772 199776 147824 199782
rect 148106 199764 148134 200124
rect 147772 199718 147824 199724
rect 147876 199736 148134 199764
rect 148198 199764 148226 200124
rect 148290 199923 148318 200124
rect 148276 199914 148332 199923
rect 148382 199918 148410 200124
rect 148276 199849 148332 199858
rect 148370 199912 148422 199918
rect 148370 199854 148422 199860
rect 148474 199764 148502 200124
rect 148566 199923 148594 200124
rect 148552 199914 148608 199923
rect 148552 199849 148608 199858
rect 148198 199736 148272 199764
rect 147494 199064 147550 199073
rect 147494 198999 147550 199008
rect 147494 195936 147550 195945
rect 147494 195871 147550 195880
rect 147508 195537 147536 195871
rect 147494 195528 147550 195537
rect 147494 195463 147550 195472
rect 147312 193180 147364 193186
rect 147312 193122 147364 193128
rect 147232 191806 147352 191834
rect 147128 191208 147180 191214
rect 147128 191150 147180 191156
rect 147324 186930 147352 191806
rect 147600 191078 147628 199702
rect 147680 199640 147732 199646
rect 147680 199582 147732 199588
rect 147692 198762 147720 199582
rect 147680 198756 147732 198762
rect 147680 198698 147732 198704
rect 147692 197470 147720 198698
rect 147680 197464 147732 197470
rect 147680 197406 147732 197412
rect 147784 196042 147812 199718
rect 147876 199170 147904 199736
rect 148140 199640 148192 199646
rect 148140 199582 148192 199588
rect 147956 199436 148008 199442
rect 147956 199378 148008 199384
rect 147968 199170 147996 199378
rect 147864 199164 147916 199170
rect 147864 199106 147916 199112
rect 147956 199164 148008 199170
rect 147956 199106 148008 199112
rect 147862 197432 147918 197441
rect 147862 197367 147918 197376
rect 147772 196036 147824 196042
rect 147772 195978 147824 195984
rect 147588 191072 147640 191078
rect 147588 191014 147640 191020
rect 147312 186924 147364 186930
rect 147312 186866 147364 186872
rect 147876 182170 147904 197367
rect 148048 196036 148100 196042
rect 148048 195978 148100 195984
rect 148060 184521 148088 195978
rect 148152 191078 148180 199582
rect 148244 197742 148272 199736
rect 148336 199736 148502 199764
rect 148658 199764 148686 200124
rect 148750 199918 148778 200124
rect 148738 199912 148790 199918
rect 148738 199854 148790 199860
rect 148842 199764 148870 200124
rect 148934 199923 148962 200124
rect 148920 199914 148976 199923
rect 149026 199918 149054 200124
rect 149118 199923 149146 200124
rect 148920 199849 148976 199858
rect 149014 199912 149066 199918
rect 149014 199854 149066 199860
rect 149104 199914 149160 199923
rect 149104 199849 149160 199858
rect 148658 199736 148732 199764
rect 148232 197736 148284 197742
rect 148232 197678 148284 197684
rect 148336 193798 148364 199736
rect 148416 199640 148468 199646
rect 148416 199582 148468 199588
rect 148600 199640 148652 199646
rect 148600 199582 148652 199588
rect 148324 193792 148376 193798
rect 148324 193734 148376 193740
rect 148322 192128 148378 192137
rect 148322 192063 148378 192072
rect 148140 191072 148192 191078
rect 148140 191014 148192 191020
rect 148230 190496 148286 190505
rect 148230 190431 148286 190440
rect 148244 187882 148272 190431
rect 148232 187876 148284 187882
rect 148232 187818 148284 187824
rect 148046 184512 148102 184521
rect 148046 184447 148102 184456
rect 147864 182164 147916 182170
rect 147864 182106 147916 182112
rect 146588 143398 146708 143426
rect 146772 143398 146984 143426
rect 145930 143032 145986 143041
rect 145930 142967 145986 142976
rect 145472 140208 145524 140214
rect 145472 140150 145524 140156
rect 145944 139890 145972 142967
rect 146588 140457 146616 143398
rect 146772 143290 146800 143398
rect 146680 143262 146800 143290
rect 146574 140448 146630 140457
rect 146574 140383 146630 140392
rect 141252 139862 141312 139890
rect 141804 139862 142140 139890
rect 142632 139862 142968 139890
rect 143644 139862 143796 139890
rect 144288 139862 144624 139890
rect 145392 139862 145452 139890
rect 145944 139862 146280 139890
rect 140424 139726 140484 139754
rect 133696 139528 133748 139534
rect 130842 139496 130898 139505
rect 133748 139476 133860 139482
rect 133696 139470 133860 139476
rect 133708 139454 133860 139470
rect 130842 139431 130898 139440
rect 146680 139369 146708 143262
rect 146760 143132 146812 143138
rect 146760 143074 146812 143080
rect 146772 139890 146800 143074
rect 147680 142996 147732 143002
rect 147680 142938 147732 142944
rect 147692 139890 147720 142938
rect 148336 142866 148364 192063
rect 148428 187066 148456 199582
rect 148508 199436 148560 199442
rect 148508 199378 148560 199384
rect 148520 199102 148548 199378
rect 148508 199096 148560 199102
rect 148508 199038 148560 199044
rect 148508 196512 148560 196518
rect 148508 196454 148560 196460
rect 148520 190126 148548 196454
rect 148612 193730 148640 199582
rect 148600 193724 148652 193730
rect 148600 193666 148652 193672
rect 148600 193044 148652 193050
rect 148600 192986 148652 192992
rect 148612 192506 148640 192986
rect 148600 192500 148652 192506
rect 148600 192442 148652 192448
rect 148704 191418 148732 199736
rect 148796 199736 148870 199764
rect 148692 191412 148744 191418
rect 148692 191354 148744 191360
rect 148796 191298 148824 199736
rect 149210 199696 149238 200124
rect 149302 199850 149330 200124
rect 149394 199850 149422 200124
rect 149290 199844 149342 199850
rect 149290 199786 149342 199792
rect 149382 199844 149434 199850
rect 149382 199786 149434 199792
rect 149486 199730 149514 200124
rect 149440 199714 149514 199730
rect 149164 199668 149238 199696
rect 149428 199708 149514 199714
rect 148876 199640 148928 199646
rect 148876 199582 148928 199588
rect 148888 198529 148916 199582
rect 148968 199368 149020 199374
rect 148968 199310 149020 199316
rect 148980 198694 149008 199310
rect 148968 198688 149020 198694
rect 148968 198630 149020 198636
rect 148874 198520 148930 198529
rect 148874 198455 148930 198464
rect 149060 197124 149112 197130
rect 149060 197066 149112 197072
rect 149072 196625 149100 197066
rect 149164 196654 149192 199668
rect 149480 199702 149514 199708
rect 149578 199696 149606 200124
rect 149670 199923 149698 200124
rect 149656 199914 149712 199923
rect 149762 199918 149790 200124
rect 149656 199849 149712 199858
rect 149750 199912 149802 199918
rect 149750 199854 149802 199860
rect 149854 199730 149882 200124
rect 149808 199702 149882 199730
rect 149578 199668 149744 199696
rect 149428 199650 149480 199656
rect 149336 199640 149388 199646
rect 149256 199588 149336 199594
rect 149256 199582 149388 199588
rect 149256 199566 149376 199582
rect 149612 199572 149664 199578
rect 149152 196648 149204 196654
rect 149058 196616 149114 196625
rect 149152 196590 149204 196596
rect 149058 196551 149114 196560
rect 149256 194546 149284 199566
rect 149612 199514 149664 199520
rect 149336 199504 149388 199510
rect 149336 199446 149388 199452
rect 149348 195022 149376 199446
rect 149520 199164 149572 199170
rect 149520 199106 149572 199112
rect 149428 198824 149480 198830
rect 149532 198801 149560 199106
rect 149428 198766 149480 198772
rect 149518 198792 149574 198801
rect 149440 198626 149468 198766
rect 149518 198727 149574 198736
rect 149624 198676 149652 199514
rect 149532 198648 149652 198676
rect 149428 198620 149480 198626
rect 149428 198562 149480 198568
rect 149336 195016 149388 195022
rect 149336 194958 149388 194964
rect 149244 194540 149296 194546
rect 149244 194482 149296 194488
rect 148876 191412 148928 191418
rect 148876 191354 148928 191360
rect 148612 191270 148824 191298
rect 148508 190120 148560 190126
rect 148508 190062 148560 190068
rect 148416 187060 148468 187066
rect 148416 187002 148468 187008
rect 148416 182164 148468 182170
rect 148416 182106 148468 182112
rect 148428 182034 148456 182106
rect 148416 182028 148468 182034
rect 148416 181970 148468 181976
rect 148324 142860 148376 142866
rect 148324 142802 148376 142808
rect 148428 141681 148456 181970
rect 148612 141778 148640 191270
rect 148692 191072 148744 191078
rect 148692 191014 148744 191020
rect 148704 144566 148732 191014
rect 148888 144702 148916 191354
rect 149152 191208 149204 191214
rect 149152 191150 149204 191156
rect 148968 187876 149020 187882
rect 148968 187818 149020 187824
rect 148980 187649 149008 187818
rect 148966 187640 149022 187649
rect 148966 187575 149022 187584
rect 148876 144696 148928 144702
rect 148876 144638 148928 144644
rect 148692 144560 148744 144566
rect 148692 144502 148744 144508
rect 148968 142180 149020 142186
rect 148968 142122 149020 142128
rect 148600 141772 148652 141778
rect 148600 141714 148652 141720
rect 148414 141672 148470 141681
rect 148414 141607 148470 141616
rect 148980 139890 149008 142122
rect 149164 141642 149192 191150
rect 149336 191072 149388 191078
rect 149336 191014 149388 191020
rect 149348 182170 149376 191014
rect 149532 189938 149560 198648
rect 149716 197354 149744 199668
rect 149808 199016 149836 199702
rect 149946 199628 149974 200124
rect 150038 199782 150066 200124
rect 150026 199776 150078 199782
rect 150130 199764 150158 200124
rect 150222 199923 150250 200124
rect 150208 199914 150264 199923
rect 150208 199849 150264 199858
rect 150314 199764 150342 200124
rect 150130 199736 150204 199764
rect 150026 199718 150078 199724
rect 149946 199600 150112 199628
rect 149888 199504 149940 199510
rect 149888 199446 149940 199452
rect 149980 199504 150032 199510
rect 149980 199446 150032 199452
rect 149900 199170 149928 199446
rect 149888 199164 149940 199170
rect 149888 199106 149940 199112
rect 149808 198988 149928 199016
rect 149794 198928 149850 198937
rect 149794 198863 149850 198872
rect 149624 197326 149744 197354
rect 149624 190097 149652 197326
rect 149808 196722 149836 198863
rect 149900 198626 149928 198988
rect 149992 198801 150020 199446
rect 149978 198792 150034 198801
rect 149978 198727 150034 198736
rect 149888 198620 149940 198626
rect 149888 198562 149940 198568
rect 150084 197354 150112 199600
rect 150176 199209 150204 199736
rect 150268 199736 150342 199764
rect 150162 199200 150218 199209
rect 150162 199135 150218 199144
rect 150162 199064 150218 199073
rect 150162 198999 150218 199008
rect 149992 197326 150112 197354
rect 149796 196716 149848 196722
rect 149796 196658 149848 196664
rect 149796 194540 149848 194546
rect 149796 194482 149848 194488
rect 149808 194002 149836 194482
rect 149796 193996 149848 194002
rect 149796 193938 149848 193944
rect 149992 191834 150020 197326
rect 150072 196716 150124 196722
rect 150072 196658 150124 196664
rect 149900 191806 150020 191834
rect 149900 191214 149928 191806
rect 149888 191208 149940 191214
rect 149888 191150 149940 191156
rect 149610 190088 149666 190097
rect 149610 190023 149666 190032
rect 149532 189910 149836 189938
rect 149704 189032 149756 189038
rect 149704 188974 149756 188980
rect 149716 188018 149744 188974
rect 149704 188012 149756 188018
rect 149704 187954 149756 187960
rect 149336 182164 149388 182170
rect 149336 182106 149388 182112
rect 149242 142760 149298 142769
rect 149242 142695 149298 142704
rect 149152 141636 149204 141642
rect 149152 141578 149204 141584
rect 146772 139862 147108 139890
rect 147692 139862 147936 139890
rect 148764 139862 149008 139890
rect 149256 139890 149284 142695
rect 149716 141817 149744 187954
rect 149808 186314 149836 189910
rect 150084 186314 150112 196658
rect 150176 189038 150204 198999
rect 150268 191078 150296 199736
rect 150406 199696 150434 200124
rect 150498 199850 150526 200124
rect 150486 199844 150538 199850
rect 150486 199786 150538 199792
rect 150590 199730 150618 200124
rect 150360 199668 150434 199696
rect 150544 199702 150618 199730
rect 150360 199578 150388 199668
rect 150348 199572 150400 199578
rect 150348 199514 150400 199520
rect 150440 199572 150492 199578
rect 150440 199514 150492 199520
rect 150348 199368 150400 199374
rect 150348 199310 150400 199316
rect 150360 199209 150388 199310
rect 150346 199200 150402 199209
rect 150346 199135 150402 199144
rect 150348 192500 150400 192506
rect 150348 192442 150400 192448
rect 150360 192137 150388 192442
rect 150346 192128 150402 192137
rect 150346 192063 150402 192072
rect 150452 191834 150480 199514
rect 150544 199442 150572 199702
rect 150682 199560 150710 200124
rect 150636 199532 150710 199560
rect 150774 199560 150802 200124
rect 150866 199628 150894 200124
rect 150958 199730 150986 200124
rect 151050 199850 151078 200124
rect 151142 199923 151170 200124
rect 151128 199914 151184 199923
rect 151038 199844 151090 199850
rect 151128 199849 151184 199858
rect 151038 199786 151090 199792
rect 150958 199702 151124 199730
rect 150992 199640 151044 199646
rect 150866 199600 150940 199628
rect 150774 199532 150848 199560
rect 150532 199436 150584 199442
rect 150532 199378 150584 199384
rect 150636 195265 150664 199532
rect 150716 199436 150768 199442
rect 150716 199378 150768 199384
rect 150728 197946 150756 199378
rect 150820 198150 150848 199532
rect 150808 198144 150860 198150
rect 150808 198086 150860 198092
rect 150716 197940 150768 197946
rect 150716 197882 150768 197888
rect 150808 196716 150860 196722
rect 150808 196658 150860 196664
rect 150622 195256 150678 195265
rect 150622 195191 150678 195200
rect 150820 192710 150848 196658
rect 150808 192704 150860 192710
rect 150808 192646 150860 192652
rect 150360 191806 150480 191834
rect 150256 191072 150308 191078
rect 150256 191014 150308 191020
rect 150164 189032 150216 189038
rect 150164 188974 150216 188980
rect 150360 187610 150388 191806
rect 150624 191208 150676 191214
rect 150624 191150 150676 191156
rect 150348 187604 150400 187610
rect 150348 187546 150400 187552
rect 149808 186286 150020 186314
rect 150084 186286 150296 186314
rect 149796 182164 149848 182170
rect 149796 182106 149848 182112
rect 149888 182164 149940 182170
rect 149888 182106 149940 182112
rect 149808 144129 149836 182106
rect 149900 181830 149928 182106
rect 149888 181824 149940 181830
rect 149888 181766 149940 181772
rect 149992 151814 150020 186286
rect 149992 151786 150112 151814
rect 149980 145716 150032 145722
rect 149980 145658 150032 145664
rect 149794 144120 149850 144129
rect 149794 144055 149850 144064
rect 149992 142390 150020 145658
rect 149980 142384 150032 142390
rect 149980 142326 150032 142332
rect 149702 141808 149758 141817
rect 149702 141743 149758 141752
rect 149992 139890 150020 142326
rect 150084 140350 150112 151786
rect 150268 148782 150296 186286
rect 150636 181626 150664 191150
rect 150624 181620 150676 181626
rect 150624 181562 150676 181568
rect 150912 178702 150940 199600
rect 150992 199582 151044 199588
rect 150900 178696 150952 178702
rect 150900 178638 150952 178644
rect 150256 148776 150308 148782
rect 150256 148718 150308 148724
rect 150900 142248 150952 142254
rect 150900 142190 150952 142196
rect 150072 140344 150124 140350
rect 150072 140286 150124 140292
rect 150912 139890 150940 142190
rect 151004 140078 151032 199582
rect 151096 198422 151124 199702
rect 151234 199696 151262 200124
rect 151188 199668 151262 199696
rect 151084 198416 151136 198422
rect 151084 198358 151136 198364
rect 151188 198268 151216 199668
rect 151326 199594 151354 200124
rect 151418 199850 151446 200124
rect 151510 199850 151538 200124
rect 151406 199844 151458 199850
rect 151406 199786 151458 199792
rect 151498 199844 151550 199850
rect 151498 199786 151550 199792
rect 151602 199730 151630 200124
rect 151694 199918 151722 200124
rect 151786 199923 151814 200124
rect 151682 199912 151734 199918
rect 151682 199854 151734 199860
rect 151772 199914 151828 199923
rect 151772 199849 151828 199858
rect 151878 199764 151906 200124
rect 151970 199918 151998 200124
rect 152062 199923 152090 200124
rect 151958 199912 152010 199918
rect 151958 199854 152010 199860
rect 152048 199914 152104 199923
rect 152048 199849 152104 199858
rect 151452 199708 151504 199714
rect 151452 199650 151504 199656
rect 151556 199702 151630 199730
rect 151832 199736 151906 199764
rect 151280 199566 151354 199594
rect 151280 199345 151308 199566
rect 151360 199504 151412 199510
rect 151360 199446 151412 199452
rect 151266 199336 151322 199345
rect 151266 199271 151322 199280
rect 151268 198892 151320 198898
rect 151268 198834 151320 198840
rect 151096 198240 151216 198268
rect 151096 193050 151124 198240
rect 151174 198112 151230 198121
rect 151174 198047 151230 198056
rect 151084 193044 151136 193050
rect 151084 192986 151136 192992
rect 151188 186314 151216 198047
rect 151096 186286 151216 186314
rect 151096 144430 151124 186286
rect 151280 180794 151308 198834
rect 151372 191214 151400 199446
rect 151464 198558 151492 199650
rect 151452 198552 151504 198558
rect 151452 198494 151504 198500
rect 151360 191208 151412 191214
rect 151360 191150 151412 191156
rect 151556 188986 151584 199702
rect 151728 199640 151780 199646
rect 151728 199582 151780 199588
rect 151740 199073 151768 199582
rect 151726 199064 151782 199073
rect 151726 198999 151782 199008
rect 151726 198384 151782 198393
rect 151726 198319 151782 198328
rect 151636 197940 151688 197946
rect 151636 197882 151688 197888
rect 151648 196654 151676 197882
rect 151636 196648 151688 196654
rect 151636 196590 151688 196596
rect 151740 191834 151768 198319
rect 151648 191806 151768 191834
rect 151832 191834 151860 199736
rect 152154 199696 152182 200124
rect 152246 199918 152274 200124
rect 152338 199918 152366 200124
rect 152430 199923 152458 200124
rect 152234 199912 152286 199918
rect 152234 199854 152286 199860
rect 152326 199912 152378 199918
rect 152326 199854 152378 199860
rect 152416 199914 152472 199923
rect 152522 199918 152550 200124
rect 152614 199918 152642 200124
rect 152706 199918 152734 200124
rect 152416 199849 152472 199858
rect 152510 199912 152562 199918
rect 152510 199854 152562 199860
rect 152602 199912 152654 199918
rect 152602 199854 152654 199860
rect 152694 199912 152746 199918
rect 152694 199854 152746 199860
rect 152464 199776 152516 199782
rect 152798 199764 152826 200124
rect 152890 199918 152918 200124
rect 152878 199912 152930 199918
rect 152878 199854 152930 199860
rect 152982 199764 153010 200124
rect 152464 199718 152516 199724
rect 152752 199736 152826 199764
rect 152936 199736 153010 199764
rect 153074 199764 153102 200124
rect 153166 199923 153194 200124
rect 153152 199914 153208 199923
rect 153152 199849 153208 199858
rect 153258 199764 153286 200124
rect 153350 199850 153378 200124
rect 153442 199918 153470 200124
rect 153534 199923 153562 200124
rect 153430 199912 153482 199918
rect 153430 199854 153482 199860
rect 153520 199914 153576 199923
rect 153626 199918 153654 200124
rect 153718 199918 153746 200124
rect 153810 199918 153838 200124
rect 153902 199918 153930 200124
rect 153338 199844 153390 199850
rect 153520 199849 153576 199858
rect 153614 199912 153666 199918
rect 153614 199854 153666 199860
rect 153706 199912 153758 199918
rect 153706 199854 153758 199860
rect 153798 199912 153850 199918
rect 153798 199854 153850 199860
rect 153890 199912 153942 199918
rect 153890 199854 153942 199860
rect 153338 199786 153390 199792
rect 153074 199736 153148 199764
rect 152280 199708 152332 199714
rect 152154 199668 152228 199696
rect 151912 199572 151964 199578
rect 151912 199514 151964 199520
rect 151924 196858 151952 199514
rect 152004 199504 152056 199510
rect 152004 199446 152056 199452
rect 151912 196852 151964 196858
rect 151912 196794 151964 196800
rect 152016 196353 152044 199446
rect 152200 198744 152228 199668
rect 152280 199650 152332 199656
rect 152292 199073 152320 199650
rect 152372 199640 152424 199646
rect 152372 199582 152424 199588
rect 152384 199510 152412 199582
rect 152372 199504 152424 199510
rect 152372 199446 152424 199452
rect 152372 199368 152424 199374
rect 152372 199310 152424 199316
rect 152278 199064 152334 199073
rect 152278 198999 152334 199008
rect 152292 198801 152320 198999
rect 152108 198716 152228 198744
rect 152278 198792 152334 198801
rect 152278 198727 152334 198736
rect 152002 196344 152058 196353
rect 152002 196279 152058 196288
rect 151832 191806 151952 191834
rect 151648 191010 151676 191806
rect 151636 191004 151688 191010
rect 151636 190946 151688 190952
rect 151924 190058 151952 191806
rect 151912 190052 151964 190058
rect 151912 189994 151964 190000
rect 152108 189038 152136 198716
rect 152384 197354 152412 199310
rect 152200 197326 152412 197354
rect 152096 189032 152148 189038
rect 151726 189000 151782 189009
rect 151556 188958 151726 188986
rect 152096 188974 152148 188980
rect 152200 188970 152228 197326
rect 152280 196852 152332 196858
rect 152280 196794 152332 196800
rect 152292 190262 152320 196794
rect 152476 195786 152504 199718
rect 152556 199640 152608 199646
rect 152556 199582 152608 199588
rect 152568 196246 152596 199582
rect 152648 199436 152700 199442
rect 152648 199378 152700 199384
rect 152556 196240 152608 196246
rect 152556 196182 152608 196188
rect 152384 195758 152504 195786
rect 152384 191834 152412 195758
rect 152556 195560 152608 195566
rect 152556 195502 152608 195508
rect 152464 195492 152516 195498
rect 152464 195434 152516 195440
rect 152476 195158 152504 195434
rect 152464 195152 152516 195158
rect 152464 195094 152516 195100
rect 152568 194818 152596 195502
rect 152556 194812 152608 194818
rect 152556 194754 152608 194760
rect 152556 193588 152608 193594
rect 152556 193530 152608 193536
rect 152384 191806 152504 191834
rect 152476 190346 152504 191806
rect 152384 190318 152504 190346
rect 152280 190256 152332 190262
rect 152280 190198 152332 190204
rect 151726 188935 151782 188944
rect 152188 188964 152240 188970
rect 151740 188465 151768 188935
rect 152188 188906 152240 188912
rect 151726 188456 151782 188465
rect 151726 188391 151782 188400
rect 152384 181558 152412 190318
rect 152464 190256 152516 190262
rect 152464 190198 152516 190204
rect 152372 181552 152424 181558
rect 152372 181494 152424 181500
rect 151188 180766 151308 180794
rect 151188 145586 151216 180766
rect 152278 145752 152334 145761
rect 152278 145687 152334 145696
rect 151176 145580 151228 145586
rect 151176 145522 151228 145528
rect 151084 144424 151136 144430
rect 151084 144366 151136 144372
rect 152004 141704 152056 141710
rect 152004 141646 152056 141652
rect 150992 140072 151044 140078
rect 150992 140014 151044 140020
rect 149256 139862 149592 139890
rect 149992 139862 150420 139890
rect 150912 139862 151248 139890
rect 152016 139754 152044 141646
rect 152292 140026 152320 145687
rect 152476 142154 152504 190198
rect 152568 144362 152596 193530
rect 152660 181762 152688 199378
rect 152752 196489 152780 199736
rect 152832 199640 152884 199646
rect 152832 199582 152884 199588
rect 152844 196994 152872 199582
rect 152832 196988 152884 196994
rect 152832 196930 152884 196936
rect 152738 196480 152794 196489
rect 152738 196415 152794 196424
rect 152740 196240 152792 196246
rect 152740 196182 152792 196188
rect 152752 194546 152780 196182
rect 152740 194540 152792 194546
rect 152740 194482 152792 194488
rect 152936 193594 152964 199736
rect 153014 199336 153070 199345
rect 153014 199271 153070 199280
rect 153028 198490 153056 199271
rect 153120 199238 153148 199736
rect 153212 199736 153286 199764
rect 153752 199776 153804 199782
rect 153108 199232 153160 199238
rect 153108 199174 153160 199180
rect 153106 198792 153162 198801
rect 153106 198727 153108 198736
rect 153160 198727 153162 198736
rect 153108 198698 153160 198704
rect 153016 198484 153068 198490
rect 153016 198426 153068 198432
rect 153028 196858 153056 198426
rect 153016 196852 153068 196858
rect 153016 196794 153068 196800
rect 152924 193588 152976 193594
rect 152924 193530 152976 193536
rect 152936 193390 152964 193530
rect 152924 193384 152976 193390
rect 152924 193326 152976 193332
rect 153212 193214 153240 199736
rect 153752 199718 153804 199724
rect 153994 199730 154022 200124
rect 154086 199918 154114 200124
rect 154074 199912 154126 199918
rect 154074 199854 154126 199860
rect 154178 199764 154206 200124
rect 154270 199923 154298 200124
rect 154256 199914 154312 199923
rect 154362 199918 154390 200124
rect 154454 199918 154482 200124
rect 154546 199918 154574 200124
rect 154638 199918 154666 200124
rect 154256 199849 154312 199858
rect 154350 199912 154402 199918
rect 154350 199854 154402 199860
rect 154442 199912 154494 199918
rect 154442 199854 154494 199860
rect 154534 199912 154586 199918
rect 154534 199854 154586 199860
rect 154626 199912 154678 199918
rect 154626 199854 154678 199860
rect 154178 199736 154252 199764
rect 153568 199708 153620 199714
rect 153568 199650 153620 199656
rect 153292 199640 153344 199646
rect 153292 199582 153344 199588
rect 153476 199640 153528 199646
rect 153476 199582 153528 199588
rect 153120 193186 153240 193214
rect 153304 193214 153332 199582
rect 153384 199572 153436 199578
rect 153384 199514 153436 199520
rect 153396 199345 153424 199514
rect 153382 199336 153438 199345
rect 153382 199271 153438 199280
rect 153488 196722 153516 199582
rect 153476 196716 153528 196722
rect 153476 196658 153528 196664
rect 153474 196072 153530 196081
rect 153474 196007 153530 196016
rect 153304 193186 153424 193214
rect 152648 181756 152700 181762
rect 152648 181698 152700 181704
rect 152556 144356 152608 144362
rect 152556 144298 152608 144304
rect 152384 142126 152504 142154
rect 152384 141545 152412 142126
rect 153016 141704 153068 141710
rect 153016 141646 153068 141652
rect 152370 141536 152426 141545
rect 152370 141471 152426 141480
rect 153028 140894 153056 141646
rect 153120 141642 153148 193186
rect 153292 191276 153344 191282
rect 153292 191218 153344 191224
rect 153304 181898 153332 191218
rect 153396 191078 153424 193186
rect 153488 191214 153516 196007
rect 153476 191208 153528 191214
rect 153476 191150 153528 191156
rect 153384 191072 153436 191078
rect 153384 191014 153436 191020
rect 153580 186314 153608 199650
rect 153660 199504 153712 199510
rect 153660 199446 153712 199452
rect 153672 196217 153700 199446
rect 153764 199374 153792 199718
rect 153994 199702 154068 199730
rect 153844 199640 153896 199646
rect 153844 199582 153896 199588
rect 153752 199368 153804 199374
rect 153752 199310 153804 199316
rect 153750 198792 153806 198801
rect 153856 198762 153884 199582
rect 153936 199572 153988 199578
rect 153936 199514 153988 199520
rect 153750 198727 153806 198736
rect 153844 198756 153896 198762
rect 153658 196208 153714 196217
rect 153658 196143 153714 196152
rect 153764 192778 153792 198727
rect 153844 198698 153896 198704
rect 153752 192772 153804 192778
rect 153752 192714 153804 192720
rect 153948 188766 153976 199514
rect 154040 199492 154068 199702
rect 154040 199464 154160 199492
rect 154028 198756 154080 198762
rect 154028 198698 154080 198704
rect 154040 192710 154068 198698
rect 154132 196518 154160 199464
rect 154120 196512 154172 196518
rect 154120 196454 154172 196460
rect 154224 195974 154252 199736
rect 154730 199730 154758 200124
rect 154822 199923 154850 200124
rect 154808 199914 154864 199923
rect 154808 199849 154864 199858
rect 154914 199764 154942 200124
rect 155006 199918 155034 200124
rect 154994 199912 155046 199918
rect 154994 199854 155046 199860
rect 154914 199736 154988 199764
rect 154304 199708 154356 199714
rect 154304 199650 154356 199656
rect 154488 199708 154540 199714
rect 154488 199650 154540 199656
rect 154580 199708 154632 199714
rect 154580 199650 154632 199656
rect 154684 199702 154758 199730
rect 154132 195946 154252 195974
rect 154028 192704 154080 192710
rect 154028 192646 154080 192652
rect 154132 191282 154160 195946
rect 154212 195628 154264 195634
rect 154212 195570 154264 195576
rect 154120 191276 154172 191282
rect 154120 191218 154172 191224
rect 154224 191162 154252 195570
rect 154040 191134 154252 191162
rect 153936 188760 153988 188766
rect 153936 188702 153988 188708
rect 153488 186286 153608 186314
rect 153488 182918 153516 186286
rect 153476 182912 153528 182918
rect 153476 182854 153528 182860
rect 153292 181892 153344 181898
rect 153292 181834 153344 181840
rect 153934 145752 153990 145761
rect 153934 145687 153990 145696
rect 153382 142896 153438 142905
rect 153382 142831 153438 142840
rect 153108 141636 153160 141642
rect 153108 141578 153160 141584
rect 153016 140888 153068 140894
rect 153016 140830 153068 140836
rect 152292 139998 152504 140026
rect 152476 139890 152504 139998
rect 153396 139890 153424 142831
rect 153948 140026 153976 145687
rect 154040 141506 154068 191134
rect 154120 191072 154172 191078
rect 154120 191014 154172 191020
rect 154132 147014 154160 191014
rect 154316 188358 154344 199650
rect 154396 199232 154448 199238
rect 154396 199174 154448 199180
rect 154408 198694 154436 199174
rect 154396 198688 154448 198694
rect 154396 198630 154448 198636
rect 154396 191208 154448 191214
rect 154396 191150 154448 191156
rect 154304 188352 154356 188358
rect 154304 188294 154356 188300
rect 154408 180794 154436 191150
rect 154500 188465 154528 199650
rect 154592 198898 154620 199650
rect 154580 198892 154632 198898
rect 154580 198834 154632 198840
rect 154684 191834 154712 199702
rect 154856 199640 154908 199646
rect 154856 199582 154908 199588
rect 154764 199572 154816 199578
rect 154764 199514 154816 199520
rect 154592 191806 154712 191834
rect 154486 188456 154542 188465
rect 154486 188391 154542 188400
rect 154592 186726 154620 191806
rect 154672 191072 154724 191078
rect 154672 191014 154724 191020
rect 154580 186720 154632 186726
rect 154580 186662 154632 186668
rect 154316 180766 154436 180794
rect 154316 151094 154344 180766
rect 154684 178838 154712 191014
rect 154776 181830 154804 199514
rect 154868 198801 154896 199582
rect 154854 198792 154910 198801
rect 154854 198727 154910 198736
rect 154856 198416 154908 198422
rect 154856 198358 154908 198364
rect 154868 198014 154896 198358
rect 154856 198008 154908 198014
rect 154856 197950 154908 197956
rect 154960 191834 154988 199736
rect 155098 199730 155126 200124
rect 155190 199764 155218 200124
rect 155282 199918 155310 200124
rect 155374 199918 155402 200124
rect 155466 199918 155494 200124
rect 155558 199918 155586 200124
rect 155650 199918 155678 200124
rect 155270 199912 155322 199918
rect 155270 199854 155322 199860
rect 155362 199912 155414 199918
rect 155362 199854 155414 199860
rect 155454 199912 155506 199918
rect 155454 199854 155506 199860
rect 155546 199912 155598 199918
rect 155546 199854 155598 199860
rect 155638 199912 155690 199918
rect 155638 199854 155690 199860
rect 155316 199776 155368 199782
rect 155190 199736 155264 199764
rect 155052 199702 155126 199730
rect 155052 197538 155080 199702
rect 155040 197532 155092 197538
rect 155040 197474 155092 197480
rect 155236 197354 155264 199736
rect 155316 199718 155368 199724
rect 155408 199776 155460 199782
rect 155742 199764 155770 200124
rect 155408 199718 155460 199724
rect 155696 199736 155770 199764
rect 155144 197326 155264 197354
rect 154960 191806 155080 191834
rect 154948 191208 155000 191214
rect 154948 191150 155000 191156
rect 154856 189644 154908 189650
rect 154856 189586 154908 189592
rect 154868 183161 154896 189586
rect 154854 183152 154910 183161
rect 154854 183087 154910 183096
rect 154960 182986 154988 191150
rect 155052 185638 155080 191806
rect 155144 189786 155172 197326
rect 155328 191834 155356 199718
rect 155420 195634 155448 199718
rect 155592 199708 155644 199714
rect 155592 199650 155644 199656
rect 155500 199640 155552 199646
rect 155500 199582 155552 199588
rect 155408 195628 155460 195634
rect 155408 195570 155460 195576
rect 155236 191806 155356 191834
rect 155132 189780 155184 189786
rect 155132 189722 155184 189728
rect 155236 189650 155264 191806
rect 155512 191214 155540 199582
rect 155500 191208 155552 191214
rect 155500 191150 155552 191156
rect 155604 191078 155632 199650
rect 155592 191072 155644 191078
rect 155592 191014 155644 191020
rect 155406 190360 155462 190369
rect 155406 190295 155462 190304
rect 155224 189644 155276 189650
rect 155224 189586 155276 189592
rect 155040 185632 155092 185638
rect 155040 185574 155092 185580
rect 154948 182980 155000 182986
rect 154948 182922 155000 182928
rect 154764 181824 154816 181830
rect 154764 181766 154816 181772
rect 154672 178832 154724 178838
rect 154672 178774 154724 178780
rect 154304 151088 154356 151094
rect 154304 151030 154356 151036
rect 154120 147008 154172 147014
rect 154120 146950 154172 146956
rect 154948 145580 155000 145586
rect 154948 145522 155000 145528
rect 154028 141500 154080 141506
rect 154028 141442 154080 141448
rect 153948 139998 154160 140026
rect 154132 139890 154160 139998
rect 154960 139890 154988 145522
rect 155420 141545 155448 190295
rect 155696 186314 155724 199736
rect 155834 199696 155862 200124
rect 155926 199918 155954 200124
rect 155914 199912 155966 199918
rect 155914 199854 155966 199860
rect 156018 199764 156046 200124
rect 155788 199668 155862 199696
rect 155972 199736 156046 199764
rect 155788 190194 155816 199668
rect 155868 199572 155920 199578
rect 155868 199514 155920 199520
rect 155776 190188 155828 190194
rect 155776 190130 155828 190136
rect 155880 190126 155908 199514
rect 155972 198121 156000 199736
rect 156110 199594 156138 200124
rect 156064 199566 156138 199594
rect 155958 198112 156014 198121
rect 155958 198047 156014 198056
rect 155958 195528 156014 195537
rect 155958 195463 156014 195472
rect 155972 195430 156000 195463
rect 155960 195424 156012 195430
rect 155960 195366 156012 195372
rect 155868 190120 155920 190126
rect 155868 190062 155920 190068
rect 155960 187264 156012 187270
rect 155960 187206 156012 187212
rect 155972 186794 156000 187206
rect 155960 186788 156012 186794
rect 155960 186730 156012 186736
rect 155604 186286 155724 186314
rect 155604 141710 155632 186286
rect 156064 179081 156092 199566
rect 156202 199560 156230 200124
rect 156294 199628 156322 200124
rect 156386 199730 156414 200124
rect 156478 199918 156506 200124
rect 156570 199918 156598 200124
rect 156466 199912 156518 199918
rect 156466 199854 156518 199860
rect 156558 199912 156610 199918
rect 156558 199854 156610 199860
rect 156512 199776 156564 199782
rect 156386 199702 156460 199730
rect 156662 199764 156690 200124
rect 156754 199918 156782 200124
rect 156846 199923 156874 200124
rect 156742 199912 156794 199918
rect 156742 199854 156794 199860
rect 156832 199914 156888 199923
rect 156832 199849 156888 199858
rect 156938 199764 156966 200124
rect 156662 199736 156736 199764
rect 156512 199718 156564 199724
rect 156294 199600 156368 199628
rect 156202 199532 156276 199560
rect 156248 198257 156276 199532
rect 156234 198248 156290 198257
rect 156234 198183 156290 198192
rect 156144 191208 156196 191214
rect 156144 191150 156196 191156
rect 156050 179072 156106 179081
rect 156156 179042 156184 191150
rect 156340 187270 156368 199600
rect 156432 199560 156460 199702
rect 156524 199628 156552 199718
rect 156524 199600 156644 199628
rect 156432 199532 156552 199560
rect 156420 199436 156472 199442
rect 156420 199378 156472 199384
rect 156432 191350 156460 199378
rect 156420 191344 156472 191350
rect 156420 191286 156472 191292
rect 156524 191162 156552 199532
rect 156616 197266 156644 199600
rect 156604 197260 156656 197266
rect 156604 197202 156656 197208
rect 156604 196172 156656 196178
rect 156604 196114 156656 196120
rect 156616 195158 156644 196114
rect 156604 195152 156656 195158
rect 156604 195094 156656 195100
rect 156708 195090 156736 199736
rect 156892 199736 156966 199764
rect 157030 199764 157058 200124
rect 157122 199918 157150 200124
rect 157214 199918 157242 200124
rect 157110 199912 157162 199918
rect 157110 199854 157162 199860
rect 157202 199912 157254 199918
rect 157202 199854 157254 199860
rect 157306 199764 157334 200124
rect 157398 199918 157426 200124
rect 157386 199912 157438 199918
rect 157386 199854 157438 199860
rect 157490 199764 157518 200124
rect 157582 199918 157610 200124
rect 157570 199912 157622 199918
rect 157570 199854 157622 199860
rect 157674 199764 157702 200124
rect 157766 199918 157794 200124
rect 157858 199923 157886 200124
rect 157754 199912 157806 199918
rect 157754 199854 157806 199860
rect 157844 199914 157900 199923
rect 157950 199918 157978 200124
rect 158042 199918 158070 200124
rect 158134 199918 158162 200124
rect 158226 199918 158254 200124
rect 158318 199918 158346 200124
rect 157844 199849 157900 199858
rect 157938 199912 157990 199918
rect 157938 199854 157990 199860
rect 158030 199912 158082 199918
rect 158030 199854 158082 199860
rect 158122 199912 158174 199918
rect 158122 199854 158174 199860
rect 158214 199912 158266 199918
rect 158214 199854 158266 199860
rect 158306 199912 158358 199918
rect 158306 199854 158358 199860
rect 157800 199776 157852 199782
rect 157030 199736 157104 199764
rect 157306 199736 157380 199764
rect 157490 199736 157564 199764
rect 157674 199736 157748 199764
rect 156788 199640 156840 199646
rect 156788 199582 156840 199588
rect 156696 195084 156748 195090
rect 156696 195026 156748 195032
rect 156524 191134 156736 191162
rect 156604 191072 156656 191078
rect 156604 191014 156656 191020
rect 156328 187264 156380 187270
rect 156328 187206 156380 187212
rect 156050 179007 156106 179016
rect 156144 179036 156196 179042
rect 156144 178978 156196 178984
rect 156616 176118 156644 191014
rect 156604 176112 156656 176118
rect 156604 176054 156656 176060
rect 156708 146946 156736 191134
rect 156800 189990 156828 199582
rect 156892 198966 156920 199736
rect 156972 199640 157024 199646
rect 156972 199582 157024 199588
rect 156984 199345 157012 199582
rect 156970 199336 157026 199345
rect 156970 199271 157026 199280
rect 156970 199200 157026 199209
rect 156970 199135 157026 199144
rect 156984 198966 157012 199135
rect 156880 198960 156932 198966
rect 156880 198902 156932 198908
rect 156972 198960 157024 198966
rect 156972 198902 157024 198908
rect 156878 198384 156934 198393
rect 156878 198319 156934 198328
rect 156892 198082 156920 198319
rect 156880 198076 156932 198082
rect 156880 198018 156932 198024
rect 156880 197260 156932 197266
rect 156880 197202 156932 197208
rect 156892 191078 156920 197202
rect 157076 196217 157104 199736
rect 157156 199708 157208 199714
rect 157156 199650 157208 199656
rect 157062 196208 157118 196217
rect 157062 196143 157118 196152
rect 156972 196036 157024 196042
rect 156972 195978 157024 195984
rect 156984 191214 157012 195978
rect 156972 191208 157024 191214
rect 156972 191150 157024 191156
rect 156880 191072 156932 191078
rect 156880 191014 156932 191020
rect 156788 189984 156840 189990
rect 156788 189926 156840 189932
rect 157168 186998 157196 199650
rect 157248 199640 157300 199646
rect 157248 199582 157300 199588
rect 157260 196042 157288 199582
rect 157352 196081 157380 199736
rect 157432 199572 157484 199578
rect 157432 199514 157484 199520
rect 157338 196072 157394 196081
rect 157248 196036 157300 196042
rect 157338 196007 157394 196016
rect 157248 195978 157300 195984
rect 157444 193934 157472 199514
rect 157432 193928 157484 193934
rect 157432 193870 157484 193876
rect 157156 186992 157208 186998
rect 157156 186934 157208 186940
rect 157536 186314 157564 199736
rect 157616 199640 157668 199646
rect 157616 199582 157668 199588
rect 157628 194818 157656 199582
rect 157616 194812 157668 194818
rect 157616 194754 157668 194760
rect 157720 194138 157748 199736
rect 157800 199718 157852 199724
rect 157892 199776 157944 199782
rect 157892 199718 157944 199724
rect 158076 199776 158128 199782
rect 158410 199764 158438 200124
rect 158502 199918 158530 200124
rect 158490 199912 158542 199918
rect 158490 199854 158542 199860
rect 158594 199764 158622 200124
rect 158686 199918 158714 200124
rect 158674 199912 158726 199918
rect 158674 199854 158726 199860
rect 158778 199764 158806 200124
rect 158870 199923 158898 200124
rect 158856 199914 158912 199923
rect 158962 199918 158990 200124
rect 159054 199923 159082 200124
rect 158856 199849 158912 199858
rect 158950 199912 159002 199918
rect 158950 199854 159002 199860
rect 159040 199914 159096 199923
rect 159146 199918 159174 200124
rect 159238 199918 159266 200124
rect 159040 199849 159096 199858
rect 159134 199912 159186 199918
rect 159134 199854 159186 199860
rect 159226 199912 159278 199918
rect 159226 199854 159278 199860
rect 158410 199736 158484 199764
rect 158594 199736 158668 199764
rect 158076 199718 158128 199724
rect 157812 199209 157840 199718
rect 157798 199200 157854 199209
rect 157798 199135 157854 199144
rect 157800 198756 157852 198762
rect 157800 198698 157852 198704
rect 157812 196110 157840 198698
rect 157904 196489 157932 199718
rect 157984 199708 158036 199714
rect 157984 199650 158036 199656
rect 157890 196480 157946 196489
rect 157890 196415 157946 196424
rect 157800 196104 157852 196110
rect 157800 196046 157852 196052
rect 157708 194132 157760 194138
rect 157708 194074 157760 194080
rect 157996 186810 158024 199650
rect 158088 189854 158116 199718
rect 158168 199640 158220 199646
rect 158168 199582 158220 199588
rect 158180 198370 158208 199582
rect 158260 199572 158312 199578
rect 158260 199514 158312 199520
rect 158272 198734 158300 199514
rect 158456 198762 158484 199736
rect 158444 198756 158496 198762
rect 158272 198706 158392 198734
rect 158180 198342 158300 198370
rect 158168 198280 158220 198286
rect 158168 198222 158220 198228
rect 158180 197198 158208 198222
rect 158272 197810 158300 198342
rect 158260 197804 158312 197810
rect 158260 197746 158312 197752
rect 158168 197192 158220 197198
rect 158168 197134 158220 197140
rect 158076 189848 158128 189854
rect 158076 189790 158128 189796
rect 158180 186998 158208 197134
rect 158364 196330 158392 198706
rect 158444 198698 158496 198704
rect 158364 196302 158576 196330
rect 158352 196104 158404 196110
rect 158352 196046 158404 196052
rect 158364 189922 158392 196046
rect 158444 194132 158496 194138
rect 158444 194074 158496 194080
rect 158352 189916 158404 189922
rect 158352 189858 158404 189864
rect 158168 186992 158220 186998
rect 158168 186934 158220 186940
rect 157996 186782 158300 186810
rect 158272 186314 158300 186782
rect 157536 186286 158208 186314
rect 158272 186286 158392 186314
rect 158180 182850 158208 186286
rect 158364 183190 158392 186286
rect 158352 183184 158404 183190
rect 158352 183126 158404 183132
rect 158168 182844 158220 182850
rect 158168 182786 158220 182792
rect 156696 146940 156748 146946
rect 156696 146882 156748 146888
rect 156604 145784 156656 145790
rect 156604 145726 156656 145732
rect 156510 142760 156566 142769
rect 156510 142695 156566 142704
rect 155592 141704 155644 141710
rect 155592 141646 155644 141652
rect 155406 141536 155462 141545
rect 155406 141471 155462 141480
rect 156524 139890 156552 142695
rect 152476 139862 152904 139890
rect 153396 139862 153732 139890
rect 154132 139862 154560 139890
rect 154960 139862 155388 139890
rect 156216 139862 156552 139890
rect 156616 139890 156644 145726
rect 157432 145648 157484 145654
rect 157432 145590 157484 145596
rect 157444 139890 157472 145590
rect 158456 141574 158484 194074
rect 158548 188834 158576 196302
rect 158640 193866 158668 199736
rect 158732 199736 158806 199764
rect 158996 199776 159048 199782
rect 158732 194138 158760 199736
rect 158996 199718 159048 199724
rect 159088 199776 159140 199782
rect 159330 199730 159358 200124
rect 159422 199923 159450 200124
rect 159408 199914 159464 199923
rect 159408 199849 159464 199858
rect 159088 199718 159140 199724
rect 158812 199436 158864 199442
rect 158812 199378 158864 199384
rect 158720 194132 158772 194138
rect 158720 194074 158772 194080
rect 158628 193860 158680 193866
rect 158628 193802 158680 193808
rect 158824 191834 158852 199378
rect 158902 198792 158958 198801
rect 158902 198727 158958 198736
rect 158640 191806 158852 191834
rect 158640 191758 158668 191806
rect 158628 191752 158680 191758
rect 158628 191694 158680 191700
rect 158916 191214 158944 198727
rect 159008 196081 159036 199718
rect 159100 199424 159128 199718
rect 159284 199702 159358 199730
rect 159100 199396 159220 199424
rect 159086 198792 159142 198801
rect 159086 198727 159142 198736
rect 159100 197062 159128 198727
rect 159088 197056 159140 197062
rect 159088 196998 159140 197004
rect 159192 196790 159220 199396
rect 159180 196784 159232 196790
rect 159180 196726 159232 196732
rect 158994 196072 159050 196081
rect 158994 196007 159050 196016
rect 158996 191276 159048 191282
rect 158996 191218 159048 191224
rect 158904 191208 158956 191214
rect 158904 191150 158956 191156
rect 158626 191040 158682 191049
rect 158626 190975 158682 190984
rect 158536 188828 158588 188834
rect 158536 188770 158588 188776
rect 158640 151814 158668 190975
rect 159008 186314 159036 191218
rect 159284 189786 159312 199702
rect 159364 199640 159416 199646
rect 159364 199582 159416 199588
rect 159376 197742 159404 199582
rect 159514 199560 159542 200124
rect 159606 199764 159634 200124
rect 159698 199918 159726 200124
rect 159686 199912 159738 199918
rect 159686 199854 159738 199860
rect 159790 199764 159818 200124
rect 159882 199918 159910 200124
rect 159870 199912 159922 199918
rect 159870 199854 159922 199860
rect 159606 199736 159680 199764
rect 159468 199532 159542 199560
rect 159468 198286 159496 199532
rect 159548 199436 159600 199442
rect 159548 199378 159600 199384
rect 159456 198280 159508 198286
rect 159456 198222 159508 198228
rect 159456 198144 159508 198150
rect 159456 198086 159508 198092
rect 159364 197736 159416 197742
rect 159364 197678 159416 197684
rect 159468 191554 159496 198086
rect 159560 196178 159588 199378
rect 159548 196172 159600 196178
rect 159548 196114 159600 196120
rect 159546 196072 159602 196081
rect 159546 196007 159602 196016
rect 159456 191548 159508 191554
rect 159456 191490 159508 191496
rect 159560 191049 159588 196007
rect 159546 191040 159602 191049
rect 159546 190975 159602 190984
rect 159272 189780 159324 189786
rect 159272 189722 159324 189728
rect 158916 186286 159036 186314
rect 158916 185706 158944 186286
rect 158904 185700 158956 185706
rect 158904 185642 158956 185648
rect 158548 151786 158668 151814
rect 158444 141568 158496 141574
rect 158444 141510 158496 141516
rect 158548 140214 158576 151786
rect 158628 142860 158680 142866
rect 158628 142802 158680 142808
rect 158536 140208 158588 140214
rect 158536 140150 158588 140156
rect 158640 139890 158668 142802
rect 159652 140078 159680 199736
rect 159744 199736 159818 199764
rect 159744 198150 159772 199736
rect 159824 199640 159876 199646
rect 159974 199628 160002 200124
rect 160066 199918 160094 200124
rect 160054 199912 160106 199918
rect 160054 199854 160106 199860
rect 160158 199764 160186 200124
rect 160250 199923 160278 200124
rect 160236 199914 160292 199923
rect 160236 199849 160292 199858
rect 160342 199850 160370 200124
rect 160434 199850 160462 200124
rect 160330 199844 160382 199850
rect 160330 199786 160382 199792
rect 160422 199844 160474 199850
rect 160422 199786 160474 199792
rect 159824 199582 159876 199588
rect 159928 199600 160002 199628
rect 160112 199736 160186 199764
rect 159836 198422 159864 199582
rect 159824 198416 159876 198422
rect 159824 198358 159876 198364
rect 159824 198212 159876 198218
rect 159824 198154 159876 198160
rect 159732 198144 159784 198150
rect 159732 198086 159784 198092
rect 159732 191208 159784 191214
rect 159732 191150 159784 191156
rect 159836 191162 159864 198154
rect 159928 191282 159956 199600
rect 160008 195696 160060 195702
rect 160008 195638 160060 195644
rect 160020 191298 160048 195638
rect 160112 191418 160140 199736
rect 160526 199730 160554 200124
rect 160480 199702 160554 199730
rect 160284 199640 160336 199646
rect 160284 199582 160336 199588
rect 160192 199368 160244 199374
rect 160192 199310 160244 199316
rect 160204 195702 160232 199310
rect 160192 195696 160244 195702
rect 160192 195638 160244 195644
rect 160100 191412 160152 191418
rect 160100 191354 160152 191360
rect 160296 191350 160324 199582
rect 160376 199436 160428 199442
rect 160376 199378 160428 199384
rect 160388 195566 160416 199378
rect 160376 195560 160428 195566
rect 160376 195502 160428 195508
rect 160376 195356 160428 195362
rect 160376 195298 160428 195304
rect 160284 191344 160336 191350
rect 159916 191276 159968 191282
rect 160020 191270 160140 191298
rect 160284 191286 160336 191292
rect 159916 191218 159968 191224
rect 159744 182889 159772 191150
rect 159836 191134 160048 191162
rect 159916 191072 159968 191078
rect 159916 191014 159968 191020
rect 159928 183122 159956 191014
rect 160020 183394 160048 191134
rect 160112 191078 160140 191270
rect 160192 191208 160244 191214
rect 160192 191150 160244 191156
rect 160100 191072 160152 191078
rect 160100 191014 160152 191020
rect 160008 183388 160060 183394
rect 160008 183330 160060 183336
rect 159916 183116 159968 183122
rect 159916 183058 159968 183064
rect 159730 182880 159786 182889
rect 159730 182815 159786 182824
rect 160204 178770 160232 191150
rect 160284 191072 160336 191078
rect 160284 191014 160336 191020
rect 160296 181694 160324 191014
rect 160388 183054 160416 195298
rect 160480 191214 160508 199702
rect 160618 199696 160646 200124
rect 160710 199918 160738 200124
rect 160802 199918 160830 200124
rect 160894 199918 160922 200124
rect 160698 199912 160750 199918
rect 160698 199854 160750 199860
rect 160790 199912 160842 199918
rect 160790 199854 160842 199860
rect 160882 199912 160934 199918
rect 160882 199854 160934 199860
rect 160744 199776 160796 199782
rect 160986 199764 161014 200124
rect 161078 199918 161106 200124
rect 161170 199918 161198 200124
rect 161262 199923 161290 200124
rect 161066 199912 161118 199918
rect 161066 199854 161118 199860
rect 161158 199912 161210 199918
rect 161158 199854 161210 199860
rect 161248 199914 161304 199923
rect 161248 199849 161304 199858
rect 161354 199850 161382 200124
rect 161446 199918 161474 200124
rect 161434 199912 161486 199918
rect 161434 199854 161486 199860
rect 161342 199844 161394 199850
rect 161342 199786 161394 199792
rect 161204 199776 161256 199782
rect 160986 199736 161060 199764
rect 160744 199718 160796 199724
rect 160618 199668 160692 199696
rect 160558 199336 160614 199345
rect 160558 199271 160614 199280
rect 160572 195362 160600 199271
rect 160664 199238 160692 199668
rect 160652 199232 160704 199238
rect 160652 199174 160704 199180
rect 160756 198694 160784 199718
rect 160836 199572 160888 199578
rect 160836 199514 160888 199520
rect 160744 198688 160796 198694
rect 160744 198630 160796 198636
rect 160560 195356 160612 195362
rect 160560 195298 160612 195304
rect 160744 194812 160796 194818
rect 160744 194754 160796 194760
rect 160560 191412 160612 191418
rect 160560 191354 160612 191360
rect 160468 191208 160520 191214
rect 160468 191150 160520 191156
rect 160572 186969 160600 191354
rect 160756 189825 160784 194754
rect 160848 191078 160876 199514
rect 160928 199368 160980 199374
rect 160928 199310 160980 199316
rect 160940 199050 160968 199310
rect 161032 199170 161060 199736
rect 161204 199718 161256 199724
rect 161112 199708 161164 199714
rect 161112 199650 161164 199656
rect 161020 199164 161072 199170
rect 161020 199106 161072 199112
rect 160940 199022 161060 199050
rect 160928 198892 160980 198898
rect 160928 198834 160980 198840
rect 160940 198218 160968 198834
rect 161032 198490 161060 199022
rect 161020 198484 161072 198490
rect 161020 198426 161072 198432
rect 160928 198212 160980 198218
rect 160928 198154 160980 198160
rect 161124 196081 161152 199650
rect 161216 199424 161244 199718
rect 161296 199708 161348 199714
rect 161296 199650 161348 199656
rect 161308 199617 161336 199650
rect 161388 199640 161440 199646
rect 161294 199608 161350 199617
rect 161538 199628 161566 200124
rect 161630 199850 161658 200124
rect 161722 199923 161750 200124
rect 161708 199914 161764 199923
rect 161814 199918 161842 200124
rect 161618 199844 161670 199850
rect 161708 199849 161764 199858
rect 161802 199912 161854 199918
rect 161802 199854 161854 199860
rect 161618 199786 161670 199792
rect 161906 199696 161934 200124
rect 161860 199668 161934 199696
rect 161538 199600 161612 199628
rect 161388 199582 161440 199588
rect 161294 199543 161350 199552
rect 161400 199492 161428 199582
rect 161400 199464 161520 199492
rect 161216 199396 161428 199424
rect 161294 199336 161350 199345
rect 161204 199300 161256 199306
rect 161294 199271 161350 199280
rect 161204 199242 161256 199248
rect 161110 196072 161166 196081
rect 161110 196007 161166 196016
rect 161216 193662 161244 199242
rect 161308 198218 161336 199271
rect 161296 198212 161348 198218
rect 161296 198154 161348 198160
rect 161294 196480 161350 196489
rect 161294 196415 161350 196424
rect 161204 193656 161256 193662
rect 161204 193598 161256 193604
rect 160928 191752 160980 191758
rect 160928 191694 160980 191700
rect 160940 191418 160968 191694
rect 160928 191412 160980 191418
rect 160928 191354 160980 191360
rect 160836 191072 160888 191078
rect 160836 191014 160888 191020
rect 160742 189816 160798 189825
rect 160742 189751 160798 189760
rect 160558 186960 160614 186969
rect 160558 186895 160614 186904
rect 160376 183048 160428 183054
rect 160376 182990 160428 182996
rect 160284 181688 160336 181694
rect 160284 181630 160336 181636
rect 160192 178764 160244 178770
rect 160192 178706 160244 178712
rect 161308 178702 161336 196415
rect 161400 191049 161428 199396
rect 161492 199306 161520 199464
rect 161480 199300 161532 199306
rect 161480 199242 161532 199248
rect 161584 199170 161612 199600
rect 161662 199608 161718 199617
rect 161662 199543 161718 199552
rect 161676 199442 161704 199543
rect 161664 199436 161716 199442
rect 161664 199378 161716 199384
rect 161480 199164 161532 199170
rect 161480 199106 161532 199112
rect 161572 199164 161624 199170
rect 161572 199106 161624 199112
rect 161492 197878 161520 199106
rect 161860 198830 161888 199668
rect 161998 199628 162026 200124
rect 162090 199730 162118 200124
rect 162182 199918 162210 200124
rect 162274 199923 162302 200124
rect 162170 199912 162222 199918
rect 162170 199854 162222 199860
rect 162260 199914 162316 199923
rect 162366 199918 162394 200124
rect 162458 199918 162486 200124
rect 162550 199918 162578 200124
rect 162260 199849 162316 199858
rect 162354 199912 162406 199918
rect 162354 199854 162406 199860
rect 162446 199912 162498 199918
rect 162446 199854 162498 199860
rect 162538 199912 162590 199918
rect 162538 199854 162590 199860
rect 162642 199850 162670 200124
rect 162630 199844 162682 199850
rect 162630 199786 162682 199792
rect 162400 199776 162452 199782
rect 162090 199702 162348 199730
rect 162400 199718 162452 199724
rect 161952 199600 162026 199628
rect 162216 199640 162268 199646
rect 161848 198824 161900 198830
rect 161848 198766 161900 198772
rect 161480 197872 161532 197878
rect 161480 197814 161532 197820
rect 161848 196036 161900 196042
rect 161848 195978 161900 195984
rect 161664 195560 161716 195566
rect 161664 195502 161716 195508
rect 161676 193798 161704 195502
rect 161664 193792 161716 193798
rect 161664 193734 161716 193740
rect 161756 191208 161808 191214
rect 161756 191150 161808 191156
rect 161386 191040 161442 191049
rect 161386 190975 161442 190984
rect 161768 185502 161796 191150
rect 161860 185570 161888 195978
rect 161952 194274 161980 199600
rect 162216 199582 162268 199588
rect 162124 199572 162176 199578
rect 162124 199514 162176 199520
rect 162032 199436 162084 199442
rect 162032 199378 162084 199384
rect 161940 194268 161992 194274
rect 161940 194210 161992 194216
rect 161952 186862 161980 194210
rect 162044 191214 162072 199378
rect 162136 199345 162164 199514
rect 162122 199336 162178 199345
rect 162122 199271 162178 199280
rect 162124 199164 162176 199170
rect 162124 199106 162176 199112
rect 162136 196042 162164 199106
rect 162228 198734 162256 199582
rect 162320 199442 162348 199702
rect 162308 199436 162360 199442
rect 162308 199378 162360 199384
rect 162228 198706 162348 198734
rect 162124 196036 162176 196042
rect 162124 195978 162176 195984
rect 162032 191208 162084 191214
rect 162032 191150 162084 191156
rect 161940 186856 161992 186862
rect 161940 186798 161992 186804
rect 161848 185564 161900 185570
rect 161848 185506 161900 185512
rect 161756 185496 161808 185502
rect 161756 185438 161808 185444
rect 161296 178696 161348 178702
rect 161296 178638 161348 178644
rect 160100 145716 160152 145722
rect 160100 145658 160152 145664
rect 159824 143200 159876 143206
rect 159824 143142 159876 143148
rect 159640 140072 159692 140078
rect 159640 140014 159692 140020
rect 159836 139890 159864 143142
rect 156616 139862 157044 139890
rect 157444 139862 157872 139890
rect 158640 139862 158700 139890
rect 159528 139862 159864 139890
rect 160112 139890 160140 145658
rect 162320 144498 162348 198706
rect 162412 194070 162440 199718
rect 162492 199708 162544 199714
rect 162492 199650 162544 199656
rect 162584 199708 162636 199714
rect 162584 199650 162636 199656
rect 162504 199617 162532 199650
rect 162490 199608 162546 199617
rect 162490 199543 162546 199552
rect 162490 199336 162546 199345
rect 162490 199271 162546 199280
rect 162400 194064 162452 194070
rect 162400 194006 162452 194012
rect 162504 193225 162532 199271
rect 162490 193216 162546 193225
rect 162490 193151 162546 193160
rect 162504 192778 162532 193151
rect 162492 192772 162544 192778
rect 162492 192714 162544 192720
rect 162596 186314 162624 199650
rect 162734 199628 162762 200124
rect 162412 186286 162624 186314
rect 162688 199600 162762 199628
rect 162412 151814 162440 186286
rect 162688 180794 162716 199600
rect 162826 199560 162854 200124
rect 162918 199923 162946 200124
rect 162904 199914 162960 199923
rect 163010 199918 163038 200124
rect 163102 199918 163130 200124
rect 163194 199918 163222 200124
rect 162904 199849 162960 199858
rect 162998 199912 163050 199918
rect 162998 199854 163050 199860
rect 163090 199912 163142 199918
rect 163090 199854 163142 199860
rect 163182 199912 163234 199918
rect 163182 199854 163234 199860
rect 163286 199764 163314 200124
rect 163378 199918 163406 200124
rect 163470 199918 163498 200124
rect 163366 199912 163418 199918
rect 163366 199854 163418 199860
rect 163458 199912 163510 199918
rect 163458 199854 163510 199860
rect 163562 199764 163590 200124
rect 163240 199736 163314 199764
rect 163516 199736 163590 199764
rect 163044 199708 163096 199714
rect 163044 199650 163096 199656
rect 162780 199532 162854 199560
rect 162780 196926 162808 199532
rect 162860 199436 162912 199442
rect 162860 199378 162912 199384
rect 162768 196920 162820 196926
rect 162768 196862 162820 196868
rect 162872 196489 162900 199378
rect 162950 199336 163006 199345
rect 162950 199271 163006 199280
rect 162858 196480 162914 196489
rect 162858 196415 162914 196424
rect 162768 191276 162820 191282
rect 162768 191218 162820 191224
rect 162780 190602 162808 191218
rect 162768 190596 162820 190602
rect 162768 190538 162820 190544
rect 162504 180766 162716 180794
rect 162504 179217 162532 180766
rect 162490 179208 162546 179217
rect 162490 179143 162546 179152
rect 162412 151786 162532 151814
rect 162400 145920 162452 145926
rect 162400 145862 162452 145868
rect 162308 144492 162360 144498
rect 162308 144434 162360 144440
rect 162308 143064 162360 143070
rect 162308 143006 162360 143012
rect 161388 142248 161440 142254
rect 161388 142190 161440 142196
rect 161400 139890 161428 142190
rect 162320 139890 162348 143006
rect 160112 139862 160356 139890
rect 161184 139862 161428 139890
rect 162012 139862 162348 139890
rect 162412 139890 162440 145862
rect 162504 144430 162532 151786
rect 162780 148986 162808 190538
rect 162768 148980 162820 148986
rect 162768 148922 162820 148928
rect 162964 144566 162992 199271
rect 163056 195129 163084 199650
rect 163136 199572 163188 199578
rect 163136 199514 163188 199520
rect 163148 196081 163176 199514
rect 163240 198490 163268 199736
rect 163412 199708 163464 199714
rect 163412 199650 163464 199656
rect 163320 199640 163372 199646
rect 163320 199582 163372 199588
rect 163228 198484 163280 198490
rect 163228 198426 163280 198432
rect 163134 196072 163190 196081
rect 163134 196007 163190 196016
rect 163042 195120 163098 195129
rect 163042 195055 163098 195064
rect 163332 194206 163360 199582
rect 163320 194200 163372 194206
rect 163320 194142 163372 194148
rect 163424 191214 163452 199650
rect 163412 191208 163464 191214
rect 163412 191150 163464 191156
rect 163516 186314 163544 199736
rect 163654 199696 163682 200124
rect 163746 199918 163774 200124
rect 163734 199912 163786 199918
rect 163734 199854 163786 199860
rect 163608 199668 163682 199696
rect 163838 199696 163866 200124
rect 163930 199923 163958 200124
rect 163916 199914 163972 199923
rect 164022 199918 164050 200124
rect 163916 199849 163972 199858
rect 164010 199912 164062 199918
rect 164010 199854 164062 199860
rect 163964 199776 164016 199782
rect 164114 199764 164142 200124
rect 164206 199923 164234 200124
rect 164192 199914 164248 199923
rect 164298 199918 164326 200124
rect 164390 199923 164418 200124
rect 164192 199849 164248 199858
rect 164286 199912 164338 199918
rect 164286 199854 164338 199860
rect 164376 199914 164432 199923
rect 164482 199918 164510 200124
rect 164376 199849 164432 199858
rect 164470 199912 164522 199918
rect 164574 199889 164602 200124
rect 164666 199918 164694 200124
rect 164654 199912 164706 199918
rect 164470 199854 164522 199860
rect 164560 199880 164616 199889
rect 164654 199854 164706 199860
rect 164560 199815 164616 199824
rect 164516 199776 164568 199782
rect 164114 199736 164188 199764
rect 163964 199718 164016 199724
rect 163838 199668 163912 199696
rect 163608 195702 163636 199668
rect 163688 199572 163740 199578
rect 163688 199514 163740 199520
rect 163700 198966 163728 199514
rect 163778 199200 163834 199209
rect 163778 199135 163834 199144
rect 163688 198960 163740 198966
rect 163688 198902 163740 198908
rect 163688 198212 163740 198218
rect 163688 198154 163740 198160
rect 163596 195696 163648 195702
rect 163596 195638 163648 195644
rect 163596 194200 163648 194206
rect 163596 194142 163648 194148
rect 163608 190058 163636 194142
rect 163596 190052 163648 190058
rect 163596 189994 163648 190000
rect 163056 186286 163544 186314
rect 163056 178673 163084 186286
rect 163042 178664 163098 178673
rect 163042 178599 163098 178608
rect 162952 144560 163004 144566
rect 162952 144502 163004 144508
rect 162492 144424 162544 144430
rect 162492 144366 162544 144372
rect 163700 140321 163728 198154
rect 163792 197282 163820 199135
rect 163884 198354 163912 199668
rect 163872 198348 163924 198354
rect 163872 198290 163924 198296
rect 163976 197849 164004 199718
rect 163962 197840 164018 197849
rect 163962 197775 164018 197784
rect 163792 197254 163912 197282
rect 163780 197192 163832 197198
rect 163780 197134 163832 197140
rect 163792 179110 163820 197134
rect 163884 189718 163912 197254
rect 164054 196344 164110 196353
rect 164054 196279 164110 196288
rect 163964 191208 164016 191214
rect 163964 191150 164016 191156
rect 163872 189712 163924 189718
rect 163872 189654 163924 189660
rect 163780 179104 163832 179110
rect 163780 179046 163832 179052
rect 163870 142896 163926 142905
rect 163870 142831 163926 142840
rect 163686 140312 163742 140321
rect 163686 140247 163742 140256
rect 163884 139890 163912 142831
rect 163976 141574 164004 191150
rect 164068 191010 164096 196279
rect 164160 195566 164188 199736
rect 164422 199744 164478 199753
rect 164240 199708 164292 199714
rect 164292 199668 164372 199696
rect 164516 199718 164568 199724
rect 164606 199744 164662 199753
rect 164422 199679 164478 199688
rect 164240 199650 164292 199656
rect 164240 199504 164292 199510
rect 164240 199446 164292 199452
rect 164252 197470 164280 199446
rect 164240 197464 164292 197470
rect 164240 197406 164292 197412
rect 164240 196716 164292 196722
rect 164240 196658 164292 196664
rect 164148 195560 164200 195566
rect 164148 195502 164200 195508
rect 164056 191004 164108 191010
rect 164056 190946 164108 190952
rect 164252 190913 164280 196658
rect 164344 196081 164372 199668
rect 164330 196072 164386 196081
rect 164330 196007 164386 196016
rect 164436 191282 164464 199679
rect 164528 196722 164556 199718
rect 164758 199730 164786 200124
rect 164850 199764 164878 200124
rect 164942 199918 164970 200124
rect 164930 199912 164982 199918
rect 164930 199854 164982 199860
rect 165034 199764 165062 200124
rect 165126 199889 165154 200124
rect 165218 199918 165246 200124
rect 165206 199912 165258 199918
rect 165112 199880 165168 199889
rect 165310 199889 165338 200124
rect 165206 199854 165258 199860
rect 165296 199880 165352 199889
rect 165112 199815 165168 199824
rect 165296 199815 165352 199824
rect 164850 199736 164924 199764
rect 164606 199679 164662 199688
rect 164712 199702 164786 199730
rect 164516 196716 164568 196722
rect 164516 196658 164568 196664
rect 164516 196580 164568 196586
rect 164516 196522 164568 196528
rect 164528 191282 164556 196522
rect 164620 193458 164648 199679
rect 164712 198150 164740 199702
rect 164792 199504 164844 199510
rect 164792 199446 164844 199452
rect 164700 198144 164752 198150
rect 164700 198086 164752 198092
rect 164608 193452 164660 193458
rect 164608 193394 164660 193400
rect 164804 193214 164832 199446
rect 164896 197130 164924 199736
rect 164988 199736 165062 199764
rect 164884 197124 164936 197130
rect 164884 197066 164936 197072
rect 164712 193186 164832 193214
rect 164424 191276 164476 191282
rect 164424 191218 164476 191224
rect 164516 191276 164568 191282
rect 164516 191218 164568 191224
rect 164712 191162 164740 193186
rect 164436 191134 164740 191162
rect 164238 190904 164294 190913
rect 164238 190839 164294 190848
rect 164436 179178 164464 191134
rect 164516 191072 164568 191078
rect 164516 191014 164568 191020
rect 164528 184754 164556 191014
rect 164988 187202 165016 199736
rect 165402 199730 165430 200124
rect 165494 199918 165522 200124
rect 165482 199912 165534 199918
rect 165482 199854 165534 199860
rect 165586 199764 165614 200124
rect 165356 199702 165430 199730
rect 165540 199736 165614 199764
rect 165678 199764 165706 200124
rect 165770 199918 165798 200124
rect 165758 199912 165810 199918
rect 165758 199854 165810 199860
rect 165862 199764 165890 200124
rect 165954 199918 165982 200124
rect 166046 199918 166074 200124
rect 165942 199912 165994 199918
rect 165942 199854 165994 199860
rect 166034 199912 166086 199918
rect 166034 199854 166086 199860
rect 165678 199736 165752 199764
rect 165862 199736 165936 199764
rect 165068 199640 165120 199646
rect 165068 199582 165120 199588
rect 165160 199640 165212 199646
rect 165160 199582 165212 199588
rect 165252 199640 165304 199646
rect 165252 199582 165304 199588
rect 165080 198121 165108 199582
rect 165066 198112 165122 198121
rect 165066 198047 165122 198056
rect 165068 198008 165120 198014
rect 165068 197950 165120 197956
rect 165080 197334 165108 197950
rect 165068 197328 165120 197334
rect 165068 197270 165120 197276
rect 165172 196586 165200 199582
rect 165264 196704 165292 199582
rect 165356 198966 165384 199702
rect 165436 199028 165488 199034
rect 165436 198970 165488 198976
rect 165344 198960 165396 198966
rect 165344 198902 165396 198908
rect 165448 198830 165476 198970
rect 165344 198824 165396 198830
rect 165344 198766 165396 198772
rect 165436 198824 165488 198830
rect 165436 198766 165488 198772
rect 165356 197402 165384 198766
rect 165344 197396 165396 197402
rect 165344 197338 165396 197344
rect 165264 196676 165384 196704
rect 165160 196580 165212 196586
rect 165160 196522 165212 196528
rect 165252 196580 165304 196586
rect 165252 196522 165304 196528
rect 165158 196208 165214 196217
rect 165158 196143 165214 196152
rect 164976 187196 165028 187202
rect 164976 187138 165028 187144
rect 165172 186314 165200 196143
rect 165264 191622 165292 196522
rect 165252 191616 165304 191622
rect 165252 191558 165304 191564
rect 165264 187338 165292 191558
rect 165356 191078 165384 196676
rect 165540 196586 165568 199736
rect 165618 199336 165674 199345
rect 165618 199271 165674 199280
rect 165632 198694 165660 199271
rect 165620 198688 165672 198694
rect 165620 198630 165672 198636
rect 165620 198348 165672 198354
rect 165620 198290 165672 198296
rect 165632 197674 165660 198290
rect 165620 197668 165672 197674
rect 165620 197610 165672 197616
rect 165528 196580 165580 196586
rect 165528 196522 165580 196528
rect 165436 193452 165488 193458
rect 165436 193394 165488 193400
rect 165344 191072 165396 191078
rect 165344 191014 165396 191020
rect 165252 187332 165304 187338
rect 165252 187274 165304 187280
rect 165172 186286 165384 186314
rect 164516 184748 164568 184754
rect 164516 184690 164568 184696
rect 164424 179172 164476 179178
rect 164424 179114 164476 179120
rect 164424 146124 164476 146130
rect 164424 146066 164476 146072
rect 164436 143682 164464 146066
rect 164884 145852 164936 145858
rect 164884 145794 164936 145800
rect 164424 143676 164476 143682
rect 164424 143618 164476 143624
rect 163964 141568 164016 141574
rect 163964 141510 164016 141516
rect 162412 139862 162840 139890
rect 163668 139862 163912 139890
rect 164436 139890 164464 143618
rect 164896 139890 164924 145794
rect 165356 141778 165384 186286
rect 165448 148510 165476 193394
rect 165724 191842 165752 199736
rect 165804 199640 165856 199646
rect 165804 199582 165856 199588
rect 165816 196353 165844 199582
rect 165908 199442 165936 199736
rect 166138 199730 166166 200124
rect 166230 199918 166258 200124
rect 166322 199918 166350 200124
rect 166414 199918 166442 200124
rect 166218 199912 166270 199918
rect 166218 199854 166270 199860
rect 166310 199912 166362 199918
rect 166310 199854 166362 199860
rect 166402 199912 166454 199918
rect 166402 199854 166454 199860
rect 166092 199702 166166 199730
rect 166264 199776 166316 199782
rect 166264 199718 166316 199724
rect 166356 199776 166408 199782
rect 166506 199764 166534 200124
rect 166598 199918 166626 200124
rect 166586 199912 166638 199918
rect 166586 199854 166638 199860
rect 166690 199764 166718 200124
rect 166782 199889 166810 200124
rect 166874 199918 166902 200124
rect 166966 199918 166994 200124
rect 166862 199912 166914 199918
rect 166768 199880 166824 199889
rect 166862 199854 166914 199860
rect 166954 199912 167006 199918
rect 166954 199854 167006 199860
rect 166768 199815 166824 199824
rect 166356 199718 166408 199724
rect 166460 199736 166534 199764
rect 166644 199736 166718 199764
rect 166908 199776 166960 199782
rect 165988 199504 166040 199510
rect 165988 199446 166040 199452
rect 165896 199436 165948 199442
rect 165896 199378 165948 199384
rect 165896 197736 165948 197742
rect 165896 197678 165948 197684
rect 165908 196586 165936 197678
rect 165896 196580 165948 196586
rect 165896 196522 165948 196528
rect 165802 196344 165858 196353
rect 165802 196279 165858 196288
rect 165632 191814 165752 191842
rect 166000 191834 166028 199446
rect 166092 196994 166120 199702
rect 166172 199640 166224 199646
rect 166172 199582 166224 199588
rect 166080 196988 166132 196994
rect 166080 196930 166132 196936
rect 166184 194002 166212 199582
rect 166172 193996 166224 194002
rect 166172 193938 166224 193944
rect 165632 190466 165660 191814
rect 165816 191806 166028 191834
rect 165712 191208 165764 191214
rect 165712 191150 165764 191156
rect 165620 190460 165672 190466
rect 165620 190402 165672 190408
rect 165632 189106 165660 190402
rect 165620 189100 165672 189106
rect 165620 189042 165672 189048
rect 165528 184748 165580 184754
rect 165528 184690 165580 184696
rect 165540 184278 165568 184690
rect 165528 184272 165580 184278
rect 165528 184214 165580 184220
rect 165436 148504 165488 148510
rect 165436 148446 165488 148452
rect 165724 147218 165752 191150
rect 165816 148578 165844 191806
rect 166276 191214 166304 199718
rect 166368 196722 166396 199718
rect 166356 196716 166408 196722
rect 166356 196658 166408 196664
rect 166460 193214 166488 199736
rect 166540 199640 166592 199646
rect 166540 199582 166592 199588
rect 166552 198898 166580 199582
rect 166540 198892 166592 198898
rect 166540 198834 166592 198840
rect 166540 198416 166592 198422
rect 166540 198358 166592 198364
rect 166552 197878 166580 198358
rect 166540 197872 166592 197878
rect 166540 197814 166592 197820
rect 166368 193186 166488 193214
rect 166264 191208 166316 191214
rect 166264 191150 166316 191156
rect 166368 189156 166396 193186
rect 165908 189128 166396 189156
rect 165908 148646 165936 189128
rect 166644 188290 166672 199736
rect 167058 199764 167086 200124
rect 167150 199918 167178 200124
rect 167138 199912 167190 199918
rect 167138 199854 167190 199860
rect 167242 199764 167270 200124
rect 166908 199718 166960 199724
rect 167012 199736 167086 199764
rect 167196 199736 167270 199764
rect 166724 199572 166776 199578
rect 166724 199514 166776 199520
rect 166816 199572 166868 199578
rect 166816 199514 166868 199520
rect 166736 198529 166764 199514
rect 166722 198520 166778 198529
rect 166722 198455 166778 198464
rect 166724 198348 166776 198354
rect 166724 198290 166776 198296
rect 166736 197810 166764 198290
rect 166724 197804 166776 197810
rect 166724 197746 166776 197752
rect 166632 188284 166684 188290
rect 166632 188226 166684 188232
rect 166264 186720 166316 186726
rect 166264 186662 166316 186668
rect 166276 181354 166304 186662
rect 166264 181348 166316 181354
rect 166264 181290 166316 181296
rect 166828 180794 166856 199514
rect 166920 198422 166948 199718
rect 166908 198416 166960 198422
rect 166908 198358 166960 198364
rect 166908 198212 166960 198218
rect 166908 198154 166960 198160
rect 166920 198014 166948 198154
rect 166908 198008 166960 198014
rect 166908 197950 166960 197956
rect 166908 196716 166960 196722
rect 166908 196658 166960 196664
rect 166920 191282 166948 196658
rect 166908 191276 166960 191282
rect 166908 191218 166960 191224
rect 167012 190398 167040 199736
rect 167092 199368 167144 199374
rect 167092 199310 167144 199316
rect 167104 198966 167132 199310
rect 167092 198960 167144 198966
rect 167092 198902 167144 198908
rect 167092 197940 167144 197946
rect 167092 197882 167144 197888
rect 167104 197334 167132 197882
rect 167092 197328 167144 197334
rect 167092 197270 167144 197276
rect 167196 196246 167224 199736
rect 167334 199696 167362 200124
rect 167426 199889 167454 200124
rect 167412 199880 167468 199889
rect 167412 199815 167468 199824
rect 167518 199764 167546 200124
rect 167610 199850 167638 200124
rect 167702 199918 167730 200124
rect 167690 199912 167742 199918
rect 167690 199854 167742 199860
rect 167598 199844 167650 199850
rect 167598 199786 167650 199792
rect 167794 199764 167822 200124
rect 167288 199668 167362 199696
rect 167472 199736 167546 199764
rect 167748 199736 167822 199764
rect 167288 197266 167316 199668
rect 167368 199572 167420 199578
rect 167368 199514 167420 199520
rect 167380 199374 167408 199514
rect 167368 199368 167420 199374
rect 167368 199310 167420 199316
rect 167276 197260 167328 197266
rect 167276 197202 167328 197208
rect 167184 196240 167236 196246
rect 167184 196182 167236 196188
rect 167472 196058 167500 199736
rect 167748 199696 167776 199736
rect 167886 199696 167914 200124
rect 167978 199764 168006 200124
rect 168070 199918 168098 200124
rect 168162 199918 168190 200124
rect 168058 199912 168110 199918
rect 168058 199854 168110 199860
rect 168150 199912 168202 199918
rect 168254 199889 168282 200124
rect 168346 199918 168374 200124
rect 168438 199918 168466 200124
rect 168530 199918 168558 200124
rect 168622 199918 168650 200124
rect 168334 199912 168386 199918
rect 168150 199854 168202 199860
rect 168240 199880 168296 199889
rect 168334 199854 168386 199860
rect 168426 199912 168478 199918
rect 168426 199854 168478 199860
rect 168518 199912 168570 199918
rect 168518 199854 168570 199860
rect 168610 199912 168662 199918
rect 168610 199854 168662 199860
rect 168240 199815 168296 199824
rect 168196 199776 168248 199782
rect 167978 199736 168144 199764
rect 167656 199668 167776 199696
rect 167840 199668 167914 199696
rect 167552 199640 167604 199646
rect 167552 199582 167604 199588
rect 167196 196030 167500 196058
rect 167000 190392 167052 190398
rect 167000 190334 167052 190340
rect 167012 189174 167040 190334
rect 167000 189168 167052 189174
rect 167000 189110 167052 189116
rect 167092 189100 167144 189106
rect 167092 189042 167144 189048
rect 167000 188420 167052 188426
rect 167000 188362 167052 188368
rect 167012 188154 167040 188362
rect 167000 188148 167052 188154
rect 167000 188090 167052 188096
rect 167104 184754 167132 189042
rect 167196 187134 167224 196030
rect 167276 195628 167328 195634
rect 167276 195570 167328 195576
rect 167184 187128 167236 187134
rect 167184 187070 167236 187076
rect 167288 186930 167316 195570
rect 167564 192438 167592 199582
rect 167656 198506 167684 199668
rect 167736 199572 167788 199578
rect 167736 199514 167788 199520
rect 167748 199481 167776 199514
rect 167734 199472 167790 199481
rect 167734 199407 167790 199416
rect 167736 199368 167788 199374
rect 167736 199310 167788 199316
rect 167748 198676 167776 199310
rect 167840 198801 167868 199668
rect 168012 199640 168064 199646
rect 168012 199582 168064 199588
rect 167920 199436 167972 199442
rect 167920 199378 167972 199384
rect 167932 198898 167960 199378
rect 167920 198892 167972 198898
rect 167920 198834 167972 198840
rect 167826 198792 167882 198801
rect 167826 198727 167882 198736
rect 167748 198648 167960 198676
rect 167656 198478 167868 198506
rect 167736 198416 167788 198422
rect 167736 198358 167788 198364
rect 167644 196240 167696 196246
rect 167644 196182 167696 196188
rect 167656 195294 167684 196182
rect 167644 195288 167696 195294
rect 167644 195230 167696 195236
rect 167552 192432 167604 192438
rect 167552 192374 167604 192380
rect 167368 189168 167420 189174
rect 167368 189110 167420 189116
rect 167458 189136 167514 189145
rect 167276 186924 167328 186930
rect 167276 186866 167328 186872
rect 167092 184748 167144 184754
rect 167092 184690 167144 184696
rect 167380 184618 167408 189110
rect 167458 189071 167514 189080
rect 167472 188426 167500 189071
rect 167460 188420 167512 188426
rect 167460 188362 167512 188368
rect 167368 184612 167420 184618
rect 167368 184554 167420 184560
rect 166736 180766 166856 180794
rect 165896 148640 165948 148646
rect 165896 148582 165948 148588
rect 165804 148572 165856 148578
rect 165804 148514 165856 148520
rect 165712 147212 165764 147218
rect 165712 147154 165764 147160
rect 166540 146056 166592 146062
rect 166540 145998 166592 146004
rect 166448 142996 166500 143002
rect 166448 142938 166500 142944
rect 165344 141772 165396 141778
rect 165344 141714 165396 141720
rect 166460 139890 166488 142938
rect 164436 139862 164496 139890
rect 164896 139862 165324 139890
rect 166152 139862 166488 139890
rect 166552 139890 166580 145998
rect 166736 144294 166764 180766
rect 167656 175982 167684 195230
rect 167748 195090 167776 198358
rect 167840 195634 167868 198478
rect 167828 195628 167880 195634
rect 167828 195570 167880 195576
rect 167736 195084 167788 195090
rect 167736 195026 167788 195032
rect 167932 194449 167960 198648
rect 167918 194440 167974 194449
rect 167918 194375 167974 194384
rect 167644 175976 167696 175982
rect 167644 175918 167696 175924
rect 167368 145988 167420 145994
rect 167368 145930 167420 145936
rect 166724 144288 166776 144294
rect 166724 144230 166776 144236
rect 167380 139890 167408 145930
rect 168024 144362 168052 199582
rect 168116 196314 168144 199736
rect 168196 199718 168248 199724
rect 168288 199776 168340 199782
rect 168714 199764 168742 200124
rect 168806 199889 168834 200124
rect 168898 199918 168926 200124
rect 168990 199918 169018 200124
rect 169082 199918 169110 200124
rect 168886 199912 168938 199918
rect 168792 199880 168848 199889
rect 168886 199854 168938 199860
rect 168978 199912 169030 199918
rect 168978 199854 169030 199860
rect 169070 199912 169122 199918
rect 169070 199854 169122 199860
rect 168792 199815 168848 199824
rect 169174 199764 169202 200124
rect 168714 199753 168788 199764
rect 168714 199744 168802 199753
rect 168714 199736 168746 199744
rect 168288 199718 168340 199724
rect 168208 198121 168236 199718
rect 168194 198112 168250 198121
rect 168194 198047 168250 198056
rect 168194 197976 168250 197985
rect 168194 197911 168250 197920
rect 168208 197878 168236 197911
rect 168196 197872 168248 197878
rect 168196 197814 168248 197820
rect 168196 197532 168248 197538
rect 168196 197474 168248 197480
rect 168104 196308 168156 196314
rect 168104 196250 168156 196256
rect 168102 196208 168158 196217
rect 168102 196143 168158 196152
rect 168116 147082 168144 196143
rect 168208 190454 168236 197474
rect 168300 195158 168328 199718
rect 168472 199708 168524 199714
rect 168746 199679 168802 199688
rect 169036 199736 169202 199764
rect 168472 199650 168524 199656
rect 168378 199608 168434 199617
rect 168378 199543 168434 199552
rect 168392 199442 168420 199543
rect 168380 199436 168432 199442
rect 168380 199378 168432 199384
rect 168484 198694 168512 199650
rect 168656 199640 168708 199646
rect 168748 199640 168800 199646
rect 168656 199582 168708 199588
rect 168746 199608 168748 199617
rect 168800 199608 168802 199617
rect 168564 199572 168616 199578
rect 168564 199514 168616 199520
rect 168472 198688 168524 198694
rect 168472 198630 168524 198636
rect 168576 198370 168604 199514
rect 168668 198801 168696 199582
rect 168930 199608 168986 199617
rect 168746 199543 168802 199552
rect 168840 199572 168892 199578
rect 168930 199543 168986 199552
rect 168840 199514 168892 199520
rect 168852 199209 168880 199514
rect 168838 199200 168894 199209
rect 168838 199135 168894 199144
rect 168654 198792 168710 198801
rect 168654 198727 168710 198736
rect 168748 198688 168800 198694
rect 168748 198630 168800 198636
rect 168576 198342 168696 198370
rect 168564 198280 168616 198286
rect 168564 198222 168616 198228
rect 168576 196926 168604 198222
rect 168668 198014 168696 198342
rect 168656 198008 168708 198014
rect 168656 197950 168708 197956
rect 168760 197010 168788 198630
rect 168852 197538 168880 199135
rect 168840 197532 168892 197538
rect 168840 197474 168892 197480
rect 168668 196982 168788 197010
rect 168564 196920 168616 196926
rect 168564 196862 168616 196868
rect 168564 196512 168616 196518
rect 168564 196454 168616 196460
rect 168378 195392 168434 195401
rect 168378 195327 168434 195336
rect 168288 195152 168340 195158
rect 168288 195094 168340 195100
rect 168392 193186 168420 195327
rect 168472 193452 168524 193458
rect 168472 193394 168524 193400
rect 168380 193180 168432 193186
rect 168380 193122 168432 193128
rect 168208 190426 168328 190454
rect 168300 148442 168328 190426
rect 168378 186144 168434 186153
rect 168378 186079 168434 186088
rect 168392 185842 168420 186079
rect 168380 185836 168432 185842
rect 168380 185778 168432 185784
rect 168392 185026 168420 185778
rect 168380 185020 168432 185026
rect 168380 184962 168432 184968
rect 168484 148481 168512 193394
rect 168576 148714 168604 196454
rect 168668 148782 168696 196982
rect 168748 196920 168800 196926
rect 168748 196862 168800 196868
rect 168760 184686 168788 196862
rect 168838 196344 168894 196353
rect 168838 196279 168894 196288
rect 168852 187406 168880 196279
rect 168944 191486 168972 199543
rect 169036 196858 169064 199736
rect 169266 199696 169294 200124
rect 169358 199764 169386 200124
rect 169450 199889 169478 200124
rect 169436 199880 169492 199889
rect 169436 199815 169492 199824
rect 169542 199764 169570 200124
rect 169634 199918 169662 200124
rect 169622 199912 169674 199918
rect 169726 199889 169754 200124
rect 169818 199918 169846 200124
rect 169910 199918 169938 200124
rect 170002 199918 170030 200124
rect 170094 199918 170122 200124
rect 170186 199918 170214 200124
rect 169806 199912 169858 199918
rect 169622 199854 169674 199860
rect 169712 199880 169768 199889
rect 169806 199854 169858 199860
rect 169898 199912 169950 199918
rect 169898 199854 169950 199860
rect 169990 199912 170042 199918
rect 169990 199854 170042 199860
rect 170082 199912 170134 199918
rect 170082 199854 170134 199860
rect 170174 199912 170226 199918
rect 170174 199854 170226 199860
rect 169712 199815 169768 199824
rect 169358 199736 169432 199764
rect 169220 199668 169294 199696
rect 169116 199504 169168 199510
rect 169116 199446 169168 199452
rect 169128 196926 169156 199446
rect 169116 196920 169168 196926
rect 169116 196862 169168 196868
rect 169024 196852 169076 196858
rect 169024 196794 169076 196800
rect 169220 196518 169248 199668
rect 169298 199472 169354 199481
rect 169298 199407 169354 199416
rect 169312 198694 169340 199407
rect 169300 198688 169352 198694
rect 169300 198630 169352 198636
rect 169300 196852 169352 196858
rect 169300 196794 169352 196800
rect 169208 196512 169260 196518
rect 169208 196454 169260 196460
rect 169208 196308 169260 196314
rect 169208 196250 169260 196256
rect 168932 191480 168984 191486
rect 168932 191422 168984 191428
rect 168944 190454 168972 191422
rect 168944 190426 169156 190454
rect 168840 187400 168892 187406
rect 168840 187342 168892 187348
rect 168748 184680 168800 184686
rect 168748 184622 168800 184628
rect 168760 180794 168788 184622
rect 168760 180766 169064 180794
rect 168656 148776 168708 148782
rect 168656 148718 168708 148724
rect 168564 148708 168616 148714
rect 168564 148650 168616 148656
rect 168470 148472 168526 148481
rect 168288 148436 168340 148442
rect 168470 148407 168526 148416
rect 168288 148378 168340 148384
rect 169036 147150 169064 180766
rect 169128 176050 169156 190426
rect 169220 180305 169248 196250
rect 169312 192846 169340 196794
rect 169300 192840 169352 192846
rect 169300 192782 169352 192788
rect 169206 180296 169262 180305
rect 169206 180231 169262 180240
rect 169116 176044 169168 176050
rect 169116 175986 169168 175992
rect 169404 148170 169432 199736
rect 169496 199736 169570 199764
rect 169760 199776 169812 199782
rect 169496 193458 169524 199736
rect 169760 199718 169812 199724
rect 170128 199776 170180 199782
rect 170128 199718 170180 199724
rect 169668 199708 169720 199714
rect 169668 199650 169720 199656
rect 169576 199640 169628 199646
rect 169576 199582 169628 199588
rect 169588 196897 169616 199582
rect 169680 199209 169708 199650
rect 169666 199200 169722 199209
rect 169666 199135 169722 199144
rect 169772 198608 169800 199718
rect 169852 199708 169904 199714
rect 169852 199650 169904 199656
rect 169864 199617 169892 199650
rect 169850 199608 169906 199617
rect 169850 199543 169906 199552
rect 170034 199472 170090 199481
rect 170034 199407 170090 199416
rect 169772 198580 169892 198608
rect 169760 198484 169812 198490
rect 169760 198426 169812 198432
rect 169772 198393 169800 198426
rect 169758 198384 169814 198393
rect 169758 198319 169814 198328
rect 169760 197940 169812 197946
rect 169760 197882 169812 197888
rect 169574 196888 169630 196897
rect 169574 196823 169576 196832
rect 169628 196823 169630 196832
rect 169576 196794 169628 196800
rect 169588 196763 169616 196794
rect 169484 193452 169536 193458
rect 169484 193394 169536 193400
rect 169772 192370 169800 197882
rect 169864 196722 169892 198580
rect 170048 198490 170076 199407
rect 170036 198484 170088 198490
rect 170036 198426 170088 198432
rect 169944 197328 169996 197334
rect 169944 197270 169996 197276
rect 169956 197033 169984 197270
rect 169942 197024 169998 197033
rect 169942 196959 169998 196968
rect 169852 196716 169904 196722
rect 169852 196658 169904 196664
rect 170140 196602 170168 199718
rect 170278 199696 170306 200124
rect 170232 199668 170306 199696
rect 170232 199374 170260 199668
rect 170370 199628 170398 200124
rect 170462 199923 170490 200124
rect 170448 199914 170504 199923
rect 170448 199849 170504 199858
rect 170554 199696 170582 200124
rect 170646 199918 170674 200124
rect 170738 199923 170766 200124
rect 170634 199912 170686 199918
rect 170634 199854 170686 199860
rect 170724 199914 170780 199923
rect 170830 199918 170858 200124
rect 170724 199849 170780 199858
rect 170818 199912 170870 199918
rect 170818 199854 170870 199860
rect 170772 199776 170824 199782
rect 170922 199764 170950 200124
rect 171014 199918 171042 200124
rect 171106 199918 171134 200124
rect 171198 199918 171226 200124
rect 171002 199912 171054 199918
rect 171002 199854 171054 199860
rect 171094 199912 171146 199918
rect 171094 199854 171146 199860
rect 171186 199912 171238 199918
rect 171186 199854 171238 199860
rect 170772 199718 170824 199724
rect 170876 199736 170950 199764
rect 171048 199776 171100 199782
rect 170324 199600 170398 199628
rect 170508 199668 170582 199696
rect 170220 199368 170272 199374
rect 170220 199310 170272 199316
rect 169864 196574 170168 196602
rect 169760 192364 169812 192370
rect 169760 192306 169812 192312
rect 169864 184414 169892 196574
rect 169944 193656 169996 193662
rect 169944 193598 169996 193604
rect 169956 192953 169984 193598
rect 169942 192944 169998 192953
rect 169942 192879 169998 192888
rect 170218 187776 170274 187785
rect 170218 187711 170274 187720
rect 170232 185774 170260 187711
rect 170324 187066 170352 199600
rect 170404 199504 170456 199510
rect 170404 199446 170456 199452
rect 170416 196926 170444 199446
rect 170404 196920 170456 196926
rect 170404 196862 170456 196868
rect 170404 196580 170456 196586
rect 170404 196522 170456 196528
rect 170416 190398 170444 196522
rect 170508 195922 170536 199668
rect 170588 199368 170640 199374
rect 170588 199310 170640 199316
rect 170600 196382 170628 199310
rect 170680 198552 170732 198558
rect 170680 198494 170732 198500
rect 170692 197334 170720 198494
rect 170680 197328 170732 197334
rect 170680 197270 170732 197276
rect 170680 196716 170732 196722
rect 170680 196658 170732 196664
rect 170588 196376 170640 196382
rect 170588 196318 170640 196324
rect 170508 195894 170628 195922
rect 170494 195800 170550 195809
rect 170494 195735 170550 195744
rect 170508 195634 170536 195735
rect 170496 195628 170548 195634
rect 170496 195570 170548 195576
rect 170600 195401 170628 195894
rect 170586 195392 170642 195401
rect 170586 195327 170642 195336
rect 170404 190392 170456 190398
rect 170404 190334 170456 190340
rect 170404 187264 170456 187270
rect 170404 187206 170456 187212
rect 170312 187060 170364 187066
rect 170312 187002 170364 187008
rect 170220 185768 170272 185774
rect 170220 185710 170272 185716
rect 169852 184408 169904 184414
rect 169852 184350 169904 184356
rect 169392 148164 169444 148170
rect 169392 148106 169444 148112
rect 169024 147144 169076 147150
rect 169024 147086 169076 147092
rect 168104 147076 168156 147082
rect 168104 147018 168156 147024
rect 170416 146962 170444 187206
rect 170692 148850 170720 196658
rect 170784 195702 170812 199718
rect 170772 195696 170824 195702
rect 170772 195638 170824 195644
rect 170770 195528 170826 195537
rect 170770 195463 170826 195472
rect 170784 191729 170812 195463
rect 170876 193662 170904 199736
rect 171048 199718 171100 199724
rect 171140 199776 171192 199782
rect 171290 199764 171318 200124
rect 171382 199923 171410 200124
rect 171368 199914 171424 199923
rect 171368 199849 171424 199858
rect 171474 199764 171502 200124
rect 171140 199718 171192 199724
rect 171244 199736 171318 199764
rect 171428 199736 171502 199764
rect 170956 199232 171008 199238
rect 170956 199174 171008 199180
rect 170968 198830 170996 199174
rect 171060 198830 171088 199718
rect 170956 198824 171008 198830
rect 170956 198766 171008 198772
rect 171048 198824 171100 198830
rect 171048 198766 171100 198772
rect 171152 197062 171180 199718
rect 171140 197056 171192 197062
rect 171140 196998 171192 197004
rect 171244 196330 171272 199736
rect 171324 199504 171376 199510
rect 171324 199446 171376 199452
rect 171336 196704 171364 199446
rect 171428 197713 171456 199736
rect 171566 199696 171594 200124
rect 171520 199668 171594 199696
rect 171658 199696 171686 200124
rect 171750 199918 171778 200124
rect 171738 199912 171790 199918
rect 171738 199854 171790 199860
rect 171842 199764 171870 200124
rect 171934 199918 171962 200124
rect 171922 199912 171974 199918
rect 171922 199854 171974 199860
rect 172026 199764 172054 200124
rect 172118 199918 172146 200124
rect 172106 199912 172158 199918
rect 172106 199854 172158 199860
rect 171842 199736 171916 199764
rect 171658 199668 171732 199696
rect 171414 197704 171470 197713
rect 171414 197639 171470 197648
rect 171336 196676 171456 196704
rect 171324 196580 171376 196586
rect 171324 196522 171376 196528
rect 170968 196302 171272 196330
rect 170968 195430 170996 196302
rect 171232 196240 171284 196246
rect 171232 196182 171284 196188
rect 170956 195424 171008 195430
rect 170956 195366 171008 195372
rect 170864 193656 170916 193662
rect 170864 193598 170916 193604
rect 170876 193361 170904 193598
rect 170862 193352 170918 193361
rect 170862 193287 170918 193296
rect 170770 191720 170826 191729
rect 170770 191655 170826 191664
rect 170784 186794 170812 191655
rect 170968 189074 170996 195366
rect 170968 189046 171088 189074
rect 170772 186788 170824 186794
rect 170772 186730 170824 186736
rect 171060 184346 171088 189046
rect 171048 184340 171100 184346
rect 171048 184282 171100 184288
rect 171244 178906 171272 196182
rect 171336 184482 171364 196522
rect 171428 193866 171456 196676
rect 171416 193860 171468 193866
rect 171416 193802 171468 193808
rect 171520 193214 171548 199668
rect 171600 199436 171652 199442
rect 171600 199378 171652 199384
rect 171612 199209 171640 199378
rect 171598 199200 171654 199209
rect 171598 199135 171654 199144
rect 171704 198558 171732 199668
rect 171784 199640 171836 199646
rect 171784 199582 171836 199588
rect 171692 198552 171744 198558
rect 171692 198494 171744 198500
rect 171796 198404 171824 199582
rect 171428 193186 171548 193214
rect 171704 198376 171824 198404
rect 171428 184550 171456 193186
rect 171704 188601 171732 198376
rect 171784 198280 171836 198286
rect 171784 198222 171836 198228
rect 171796 197742 171824 198222
rect 171784 197736 171836 197742
rect 171784 197678 171836 197684
rect 171784 196784 171836 196790
rect 171784 196726 171836 196732
rect 171690 188592 171746 188601
rect 171690 188527 171746 188536
rect 171416 184544 171468 184550
rect 171416 184486 171468 184492
rect 171324 184476 171376 184482
rect 171324 184418 171376 184424
rect 171232 178900 171284 178906
rect 171232 178842 171284 178848
rect 170680 148844 170732 148850
rect 170680 148786 170732 148792
rect 170416 146934 170720 146962
rect 168012 144356 168064 144362
rect 168012 144298 168064 144304
rect 170586 144120 170642 144129
rect 170586 144055 170642 144064
rect 168932 143132 168984 143138
rect 168932 143074 168984 143080
rect 168840 142248 168892 142254
rect 168840 142190 168892 142196
rect 168852 140758 168880 142190
rect 168840 140752 168892 140758
rect 168840 140694 168892 140700
rect 168944 139890 168972 143074
rect 169668 142928 169720 142934
rect 169668 142870 169720 142876
rect 169680 139890 169708 142870
rect 170600 139890 170628 144055
rect 166552 139862 166980 139890
rect 167380 139862 167808 139890
rect 168636 139862 168972 139890
rect 169464 139862 169708 139890
rect 170292 139862 170628 139890
rect 152016 139726 152076 139754
rect 170692 139369 170720 146934
rect 171508 146260 171560 146266
rect 171508 146202 171560 146208
rect 171046 143032 171102 143041
rect 171046 142967 171102 142976
rect 171060 139890 171088 142967
rect 171520 139890 171548 146202
rect 171796 141370 171824 196726
rect 171888 196586 171916 199736
rect 171980 199736 172054 199764
rect 171980 198558 172008 199736
rect 172060 199640 172112 199646
rect 172060 199582 172112 199588
rect 172210 199594 172238 200124
rect 172302 199918 172330 200124
rect 172290 199912 172342 199918
rect 172290 199854 172342 199860
rect 172394 199696 172422 200124
rect 172348 199668 172422 199696
rect 171968 198552 172020 198558
rect 171968 198494 172020 198500
rect 172072 198506 172100 199582
rect 172210 199566 172284 199594
rect 172072 198478 172192 198506
rect 172060 197464 172112 197470
rect 172060 197406 172112 197412
rect 171968 196784 172020 196790
rect 171968 196726 172020 196732
rect 171876 196580 171928 196586
rect 171876 196522 171928 196528
rect 171980 184210 172008 196726
rect 171968 184204 172020 184210
rect 171968 184146 172020 184152
rect 171980 180794 172008 184146
rect 171888 180766 172008 180794
rect 171888 151162 171916 180766
rect 171876 151156 171928 151162
rect 171876 151098 171928 151104
rect 171784 141364 171836 141370
rect 171784 141306 171836 141312
rect 172072 140282 172100 197406
rect 172164 194177 172192 198478
rect 172256 196246 172284 199566
rect 172244 196240 172296 196246
rect 172244 196182 172296 196188
rect 172150 194168 172206 194177
rect 172150 194103 172206 194112
rect 172152 193996 172204 194002
rect 172152 193938 172204 193944
rect 172164 148238 172192 193938
rect 172348 180794 172376 199668
rect 172486 199628 172514 200124
rect 172440 199600 172514 199628
rect 172578 199628 172606 200124
rect 172670 199764 172698 200124
rect 172762 199923 172790 200124
rect 172748 199914 172804 199923
rect 172854 199918 172882 200124
rect 172946 199918 172974 200124
rect 173038 199918 173066 200124
rect 172748 199849 172804 199858
rect 172842 199912 172894 199918
rect 172842 199854 172894 199860
rect 172934 199912 172986 199918
rect 172934 199854 172986 199860
rect 173026 199912 173078 199918
rect 173026 199854 173078 199860
rect 172796 199776 172848 199782
rect 172670 199736 172744 199764
rect 172578 199600 172652 199628
rect 172440 198665 172468 199600
rect 172520 199504 172572 199510
rect 172520 199446 172572 199452
rect 172426 198656 172482 198665
rect 172532 198626 172560 199446
rect 172426 198591 172482 198600
rect 172520 198620 172572 198626
rect 172520 198562 172572 198568
rect 172428 198484 172480 198490
rect 172428 198426 172480 198432
rect 172440 198286 172468 198426
rect 172520 198348 172572 198354
rect 172520 198290 172572 198296
rect 172428 198280 172480 198286
rect 172428 198222 172480 198228
rect 172532 197810 172560 198290
rect 172520 197804 172572 197810
rect 172520 197746 172572 197752
rect 172624 188902 172652 199600
rect 172716 197878 172744 199736
rect 172796 199718 172848 199724
rect 172808 198665 172836 199718
rect 173130 199560 173158 200124
rect 173222 199923 173250 200124
rect 173208 199914 173264 199923
rect 173314 199918 173342 200124
rect 173406 199918 173434 200124
rect 173498 199918 173526 200124
rect 173590 199918 173618 200124
rect 173682 199918 173710 200124
rect 173774 199918 173802 200124
rect 173866 199918 173894 200124
rect 173958 199923 173986 200124
rect 173208 199849 173264 199858
rect 173302 199912 173354 199918
rect 173302 199854 173354 199860
rect 173394 199912 173446 199918
rect 173394 199854 173446 199860
rect 173486 199912 173538 199918
rect 173486 199854 173538 199860
rect 173578 199912 173630 199918
rect 173578 199854 173630 199860
rect 173670 199912 173722 199918
rect 173670 199854 173722 199860
rect 173762 199912 173814 199918
rect 173762 199854 173814 199860
rect 173854 199912 173906 199918
rect 173854 199854 173906 199860
rect 173944 199914 174000 199923
rect 173944 199849 174000 199858
rect 173256 199776 173308 199782
rect 173256 199718 173308 199724
rect 173348 199776 173400 199782
rect 173348 199718 173400 199724
rect 173532 199776 173584 199782
rect 173624 199776 173676 199782
rect 173532 199718 173584 199724
rect 173622 199744 173624 199753
rect 174050 199764 174078 200124
rect 174142 199923 174170 200124
rect 174128 199914 174184 199923
rect 174128 199849 174184 199858
rect 174234 199764 174262 200124
rect 174050 199753 174124 199764
rect 173676 199744 173678 199753
rect 174050 199744 174138 199753
rect 174050 199736 174082 199744
rect 173084 199532 173158 199560
rect 172980 199504 173032 199510
rect 172900 199464 172980 199492
rect 172794 198656 172850 198665
rect 172794 198591 172850 198600
rect 172796 198484 172848 198490
rect 172796 198426 172848 198432
rect 172704 197872 172756 197878
rect 172704 197814 172756 197820
rect 172808 194002 172836 198426
rect 172900 195634 172928 199464
rect 172980 199446 173032 199452
rect 172980 199368 173032 199374
rect 172980 199310 173032 199316
rect 172888 195628 172940 195634
rect 172888 195570 172940 195576
rect 172796 193996 172848 194002
rect 172796 193938 172848 193944
rect 172992 193730 173020 199310
rect 173084 198490 173112 199532
rect 173072 198484 173124 198490
rect 173072 198426 173124 198432
rect 173072 198280 173124 198286
rect 173072 198222 173124 198228
rect 173084 197606 173112 198222
rect 173164 197940 173216 197946
rect 173164 197882 173216 197888
rect 173072 197600 173124 197606
rect 173072 197542 173124 197548
rect 173176 196602 173204 197882
rect 173268 196790 173296 199718
rect 173360 197946 173388 199718
rect 173544 199617 173572 199718
rect 173622 199679 173678 199688
rect 174082 199679 174138 199688
rect 174188 199736 174262 199764
rect 173530 199608 173586 199617
rect 173530 199543 173586 199552
rect 173716 199572 173768 199578
rect 173716 199514 173768 199520
rect 173530 198656 173586 198665
rect 173530 198591 173586 198600
rect 173348 197940 173400 197946
rect 173348 197882 173400 197888
rect 173440 197396 173492 197402
rect 173440 197338 173492 197344
rect 173256 196784 173308 196790
rect 173256 196726 173308 196732
rect 173176 196574 173296 196602
rect 173164 193928 173216 193934
rect 173164 193870 173216 193876
rect 172980 193724 173032 193730
rect 172980 193666 173032 193672
rect 172612 188896 172664 188902
rect 172612 188838 172664 188844
rect 172256 180766 172376 180794
rect 172256 164898 172284 180766
rect 172244 164892 172296 164898
rect 172244 164834 172296 164840
rect 172152 148232 172204 148238
rect 172152 148174 172204 148180
rect 172520 146192 172572 146198
rect 172520 146134 172572 146140
rect 172060 140276 172112 140282
rect 172060 140218 172112 140224
rect 172532 139890 172560 146134
rect 173176 141914 173204 193870
rect 173268 192914 173296 196574
rect 173348 193724 173400 193730
rect 173348 193666 173400 193672
rect 173256 192908 173308 192914
rect 173256 192850 173308 192856
rect 173268 192302 173296 192850
rect 173256 192296 173308 192302
rect 173256 192238 173308 192244
rect 173360 151298 173388 193666
rect 173348 151292 173400 151298
rect 173348 151234 173400 151240
rect 173164 141908 173216 141914
rect 173164 141850 173216 141856
rect 173452 140593 173480 197338
rect 173544 188698 173572 198591
rect 173622 196888 173678 196897
rect 173622 196823 173678 196832
rect 173636 192982 173664 196823
rect 173624 192976 173676 192982
rect 173624 192918 173676 192924
rect 173728 190330 173756 199514
rect 173900 199504 173952 199510
rect 173820 199464 173900 199492
rect 173820 192545 173848 199464
rect 173900 199446 173952 199452
rect 174082 198656 174138 198665
rect 174082 198591 174138 198600
rect 174096 196364 174124 198591
rect 174188 196518 174216 199736
rect 174326 199696 174354 200124
rect 174280 199668 174354 199696
rect 174280 196897 174308 199668
rect 174418 199628 174446 200124
rect 174510 199764 174538 200124
rect 174602 199918 174630 200124
rect 174590 199912 174642 199918
rect 174590 199854 174642 199860
rect 174510 199736 174584 199764
rect 174372 199600 174446 199628
rect 174266 196888 174322 196897
rect 174266 196823 174322 196832
rect 174176 196512 174228 196518
rect 174176 196454 174228 196460
rect 173912 196336 174124 196364
rect 173806 192536 173862 192545
rect 173806 192471 173862 192480
rect 173912 191146 173940 196336
rect 173992 196036 174044 196042
rect 173992 195978 174044 195984
rect 173900 191140 173952 191146
rect 173900 191082 173952 191088
rect 173716 190324 173768 190330
rect 173716 190266 173768 190272
rect 173532 188692 173584 188698
rect 173532 188634 173584 188640
rect 173728 184686 173756 190266
rect 173716 184680 173768 184686
rect 173716 184622 173768 184628
rect 173808 144764 173860 144770
rect 173808 144706 173860 144712
rect 173820 143206 173848 144706
rect 174004 144702 174032 195978
rect 174372 194274 174400 199600
rect 174452 199436 174504 199442
rect 174452 199378 174504 199384
rect 174464 197033 174492 199378
rect 174556 198014 174584 199736
rect 174694 199730 174722 200124
rect 174786 199889 174814 200124
rect 174772 199880 174828 199889
rect 174772 199815 174828 199824
rect 174694 199702 174768 199730
rect 174636 199640 174688 199646
rect 174636 199582 174688 199588
rect 174544 198008 174596 198014
rect 174544 197950 174596 197956
rect 174544 197804 174596 197810
rect 174544 197746 174596 197752
rect 174556 197282 174584 197746
rect 174648 197354 174676 199582
rect 174740 197606 174768 199702
rect 174878 199594 174906 200124
rect 174970 199918 174998 200124
rect 175062 199923 175090 200124
rect 174958 199912 175010 199918
rect 174958 199854 175010 199860
rect 175048 199914 175104 199923
rect 175048 199849 175104 199858
rect 175154 199764 175182 200124
rect 175002 199744 175058 199753
rect 175002 199679 175058 199688
rect 175108 199736 175182 199764
rect 175246 199764 175274 200124
rect 175338 199889 175366 200124
rect 175324 199880 175380 199889
rect 175324 199815 175380 199824
rect 175430 199764 175458 200124
rect 175522 199918 175550 200124
rect 175614 199918 175642 200124
rect 175706 199918 175734 200124
rect 175798 199918 175826 200124
rect 175510 199912 175562 199918
rect 175510 199854 175562 199860
rect 175602 199912 175654 199918
rect 175602 199854 175654 199860
rect 175694 199912 175746 199918
rect 175694 199854 175746 199860
rect 175786 199912 175838 199918
rect 175786 199854 175838 199860
rect 175890 199764 175918 200124
rect 175246 199736 175320 199764
rect 175430 199736 175504 199764
rect 174832 199566 174906 199594
rect 174832 198121 174860 199566
rect 174912 199300 174964 199306
rect 174912 199242 174964 199248
rect 174924 199209 174952 199242
rect 174910 199200 174966 199209
rect 174910 199135 174966 199144
rect 174818 198112 174874 198121
rect 174818 198047 174874 198056
rect 174820 198008 174872 198014
rect 174820 197950 174872 197956
rect 174728 197600 174780 197606
rect 174728 197542 174780 197548
rect 174648 197326 174768 197354
rect 174556 197254 174676 197282
rect 174450 197024 174506 197033
rect 174450 196959 174506 196968
rect 174544 196716 174596 196722
rect 174544 196658 174596 196664
rect 174360 194268 174412 194274
rect 174360 194210 174412 194216
rect 174084 194200 174136 194206
rect 174084 194142 174136 194148
rect 174096 184210 174124 194142
rect 174176 191752 174228 191758
rect 174176 191694 174228 191700
rect 174188 190602 174216 191694
rect 174176 190596 174228 190602
rect 174176 190538 174228 190544
rect 174188 187474 174216 190538
rect 174176 187468 174228 187474
rect 174176 187410 174228 187416
rect 174084 184204 174136 184210
rect 174084 184146 174136 184152
rect 174556 148374 174584 196658
rect 174648 190454 174676 197254
rect 174740 191758 174768 197326
rect 174728 191752 174780 191758
rect 174728 191694 174780 191700
rect 174832 190454 174860 197950
rect 174912 197600 174964 197606
rect 174912 197542 174964 197548
rect 174924 194886 174952 197542
rect 175016 196042 175044 199679
rect 175004 196036 175056 196042
rect 175004 195978 175056 195984
rect 174912 194880 174964 194886
rect 174912 194822 174964 194828
rect 175108 194206 175136 199736
rect 175292 197606 175320 199736
rect 175280 197600 175332 197606
rect 175280 197542 175332 197548
rect 175476 197334 175504 199736
rect 175844 199736 175918 199764
rect 175648 199708 175700 199714
rect 175648 199650 175700 199656
rect 175556 199640 175608 199646
rect 175556 199582 175608 199588
rect 175568 198665 175596 199582
rect 175554 198656 175610 198665
rect 175554 198591 175610 198600
rect 175556 198484 175608 198490
rect 175556 198426 175608 198432
rect 175188 197328 175240 197334
rect 175188 197270 175240 197276
rect 175464 197328 175516 197334
rect 175464 197270 175516 197276
rect 175200 196722 175228 197270
rect 175188 196716 175240 196722
rect 175188 196658 175240 196664
rect 175280 196172 175332 196178
rect 175280 196114 175332 196120
rect 175188 195152 175240 195158
rect 175188 195094 175240 195100
rect 175200 194954 175228 195094
rect 175188 194948 175240 194954
rect 175188 194890 175240 194896
rect 175096 194200 175148 194206
rect 175096 194142 175148 194148
rect 175004 191888 175056 191894
rect 175004 191830 175056 191836
rect 175016 191146 175044 191830
rect 175004 191140 175056 191146
rect 175004 191082 175056 191088
rect 174648 190426 174768 190454
rect 174832 190426 175228 190454
rect 174544 148368 174596 148374
rect 174544 148310 174596 148316
rect 173992 144696 174044 144702
rect 173992 144638 174044 144644
rect 173808 143200 173860 143206
rect 173714 143168 173770 143177
rect 173808 143142 173860 143148
rect 173714 143103 173770 143112
rect 173438 140584 173494 140593
rect 173438 140519 173494 140528
rect 173728 139890 173756 143103
rect 174636 141840 174688 141846
rect 174636 141782 174688 141788
rect 174648 140826 174676 141782
rect 174740 141234 174768 190426
rect 175096 144832 175148 144838
rect 175096 144774 175148 144780
rect 174728 141228 174780 141234
rect 174728 141170 174780 141176
rect 174636 140820 174688 140826
rect 174636 140762 174688 140768
rect 174648 139890 174676 140762
rect 171060 139862 171120 139890
rect 171520 139862 171948 139890
rect 172532 139862 172776 139890
rect 173604 139862 173756 139890
rect 174432 139862 174676 139890
rect 175108 139890 175136 144774
rect 175200 144634 175228 190426
rect 175292 148306 175320 196114
rect 175464 196104 175516 196110
rect 175464 196046 175516 196052
rect 175476 181762 175504 196046
rect 175568 186114 175596 198426
rect 175660 187270 175688 199650
rect 175740 196036 175792 196042
rect 175740 195978 175792 195984
rect 175752 188086 175780 195978
rect 175844 195498 175872 199736
rect 175982 199696 176010 200124
rect 176074 199918 176102 200124
rect 176062 199912 176114 199918
rect 176062 199854 176114 199860
rect 176166 199850 176194 200124
rect 176154 199844 176206 199850
rect 176154 199786 176206 199792
rect 175936 199668 176010 199696
rect 176108 199708 176160 199714
rect 175936 198490 175964 199668
rect 176108 199650 176160 199656
rect 176120 199617 176148 199650
rect 176106 199608 176162 199617
rect 176258 199594 176286 200124
rect 176350 199696 176378 200124
rect 176442 199918 176470 200124
rect 176534 199918 176562 200124
rect 176430 199912 176482 199918
rect 176430 199854 176482 199860
rect 176522 199912 176574 199918
rect 176522 199854 176574 199860
rect 176626 199764 176654 200124
rect 176580 199736 176654 199764
rect 176718 199764 176746 200124
rect 176810 199889 176838 200124
rect 176796 199880 176852 199889
rect 176796 199815 176852 199824
rect 176902 199764 176930 200124
rect 176994 199918 177022 200124
rect 176982 199912 177034 199918
rect 177086 199889 177114 200124
rect 176982 199854 177034 199860
rect 177072 199880 177128 199889
rect 177072 199815 177128 199824
rect 177028 199776 177080 199782
rect 176718 199736 176792 199764
rect 176902 199736 176976 199764
rect 176350 199668 176424 199696
rect 176258 199566 176332 199594
rect 176106 199543 176162 199552
rect 176108 199504 176160 199510
rect 176108 199446 176160 199452
rect 175924 198484 175976 198490
rect 175924 198426 175976 198432
rect 176016 198484 176068 198490
rect 176016 198426 176068 198432
rect 176028 198354 176056 198426
rect 176016 198348 176068 198354
rect 176016 198290 176068 198296
rect 176120 197354 176148 199446
rect 176028 197326 176148 197354
rect 175924 197260 175976 197266
rect 175924 197202 175976 197208
rect 175832 195492 175884 195498
rect 175832 195434 175884 195440
rect 175936 195242 175964 197202
rect 176028 196042 176056 197326
rect 176304 196110 176332 199566
rect 176396 199442 176424 199668
rect 176384 199436 176436 199442
rect 176384 199378 176436 199384
rect 176476 199436 176528 199442
rect 176476 199378 176528 199384
rect 176384 199300 176436 199306
rect 176384 199242 176436 199248
rect 176396 196178 176424 199242
rect 176488 198762 176516 199378
rect 176476 198756 176528 198762
rect 176476 198698 176528 198704
rect 176580 197354 176608 199736
rect 176660 199572 176712 199578
rect 176660 199514 176712 199520
rect 176672 198490 176700 199514
rect 176764 198490 176792 199736
rect 176844 199640 176896 199646
rect 176842 199608 176844 199617
rect 176896 199608 176898 199617
rect 176842 199543 176898 199552
rect 176844 199504 176896 199510
rect 176844 199446 176896 199452
rect 176856 199209 176884 199446
rect 176842 199200 176898 199209
rect 176842 199135 176898 199144
rect 176948 198762 176976 199736
rect 177028 199718 177080 199724
rect 176936 198756 176988 198762
rect 176936 198698 176988 198704
rect 176660 198484 176712 198490
rect 176660 198426 176712 198432
rect 176752 198484 176804 198490
rect 176752 198426 176804 198432
rect 176488 197326 176608 197354
rect 176384 196172 176436 196178
rect 176384 196114 176436 196120
rect 176292 196104 176344 196110
rect 176292 196046 176344 196052
rect 176016 196036 176068 196042
rect 176016 195978 176068 195984
rect 176292 195492 176344 195498
rect 176292 195434 176344 195440
rect 175936 195214 176056 195242
rect 175922 194032 175978 194041
rect 175922 193967 175978 193976
rect 175936 191622 175964 193967
rect 175924 191616 175976 191622
rect 175924 191558 175976 191564
rect 175740 188080 175792 188086
rect 175740 188022 175792 188028
rect 175648 187264 175700 187270
rect 175648 187206 175700 187212
rect 175556 186108 175608 186114
rect 175556 186050 175608 186056
rect 175464 181756 175516 181762
rect 175464 181698 175516 181704
rect 176028 151230 176056 195214
rect 176016 151224 176068 151230
rect 176016 151166 176068 151172
rect 176304 149054 176332 195434
rect 176488 194206 176516 197326
rect 176568 197260 176620 197266
rect 176568 197202 176620 197208
rect 176580 196382 176608 197202
rect 176568 196376 176620 196382
rect 176568 196318 176620 196324
rect 176658 196072 176714 196081
rect 176658 196007 176714 196016
rect 176752 196036 176804 196042
rect 176476 194200 176528 194206
rect 176476 194142 176528 194148
rect 176672 185978 176700 196007
rect 176752 195978 176804 195984
rect 176764 186318 176792 195978
rect 176936 195764 176988 195770
rect 176936 195706 176988 195712
rect 176948 195498 176976 195706
rect 176936 195492 176988 195498
rect 176936 195434 176988 195440
rect 177040 191834 177068 199718
rect 177178 199696 177206 200124
rect 177270 199918 177298 200124
rect 177258 199912 177310 199918
rect 177258 199854 177310 199860
rect 177362 199764 177390 200124
rect 177454 199918 177482 200124
rect 177442 199912 177494 199918
rect 177442 199854 177494 199860
rect 177546 199832 177574 200124
rect 177652 200110 177896 200138
rect 177948 200126 178000 200132
rect 177764 199980 177816 199986
rect 177764 199922 177816 199928
rect 177546 199804 177620 199832
rect 177362 199736 177528 199764
rect 177178 199668 177252 199696
rect 177224 199238 177252 199668
rect 177304 199640 177356 199646
rect 177304 199582 177356 199588
rect 177316 199442 177344 199582
rect 177304 199436 177356 199442
rect 177304 199378 177356 199384
rect 177212 199232 177264 199238
rect 177212 199174 177264 199180
rect 177120 198756 177172 198762
rect 177500 198744 177528 199736
rect 177120 198698 177172 198704
rect 177316 198716 177528 198744
rect 177132 194342 177160 198698
rect 177316 196042 177344 198716
rect 177488 198620 177540 198626
rect 177488 198562 177540 198568
rect 177396 198348 177448 198354
rect 177396 198290 177448 198296
rect 177304 196036 177356 196042
rect 177304 195978 177356 195984
rect 177304 195356 177356 195362
rect 177304 195298 177356 195304
rect 177316 194886 177344 195298
rect 177304 194880 177356 194886
rect 177304 194822 177356 194828
rect 177302 194712 177358 194721
rect 177302 194647 177358 194656
rect 177120 194336 177172 194342
rect 177120 194278 177172 194284
rect 177132 193934 177160 194278
rect 177120 193928 177172 193934
rect 177120 193870 177172 193876
rect 177316 193322 177344 194647
rect 177304 193316 177356 193322
rect 177304 193258 177356 193264
rect 176948 191806 177068 191834
rect 176948 188630 176976 191806
rect 176936 188624 176988 188630
rect 176936 188566 176988 188572
rect 177316 187542 177344 193258
rect 177408 187542 177436 198290
rect 177304 187536 177356 187542
rect 177304 187478 177356 187484
rect 177396 187536 177448 187542
rect 177396 187478 177448 187484
rect 176752 186312 176804 186318
rect 176752 186254 176804 186260
rect 176660 185972 176712 185978
rect 176660 185914 176712 185920
rect 176672 185842 176700 185914
rect 176660 185836 176712 185842
rect 176660 185778 176712 185784
rect 176568 183116 176620 183122
rect 176568 183058 176620 183064
rect 176384 183048 176436 183054
rect 176384 182990 176436 182996
rect 176292 149048 176344 149054
rect 176292 148990 176344 148996
rect 175280 148300 175332 148306
rect 175280 148242 175332 148248
rect 175188 144628 175240 144634
rect 175188 144570 175240 144576
rect 176396 144401 176424 182990
rect 176474 180296 176530 180305
rect 176474 180231 176530 180240
rect 176382 144392 176438 144401
rect 176382 144327 176438 144336
rect 176384 142452 176436 142458
rect 176384 142394 176436 142400
rect 176396 139890 176424 142394
rect 175108 139862 175260 139890
rect 176088 139862 176424 139890
rect 176488 139369 176516 180231
rect 176580 140554 176608 183058
rect 176764 181422 176792 186254
rect 177304 184816 177356 184822
rect 177304 184758 177356 184764
rect 176752 181416 176804 181422
rect 176752 181358 176804 181364
rect 177316 178974 177344 184758
rect 177304 178968 177356 178974
rect 177304 178910 177356 178916
rect 177500 148918 177528 198562
rect 177592 197962 177620 199804
rect 177672 199436 177724 199442
rect 177672 199378 177724 199384
rect 177684 198529 177712 199378
rect 177670 198520 177726 198529
rect 177670 198455 177726 198464
rect 177776 198286 177804 199922
rect 177764 198280 177816 198286
rect 177764 198222 177816 198228
rect 177592 197934 177712 197962
rect 177580 197872 177632 197878
rect 177580 197814 177632 197820
rect 177592 190262 177620 197814
rect 177684 197810 177712 197934
rect 177868 197878 177896 200110
rect 177948 200048 178000 200054
rect 177948 199990 178000 199996
rect 177960 199782 177988 199990
rect 177948 199776 178000 199782
rect 177948 199718 178000 199724
rect 177948 198008 178000 198014
rect 177948 197950 178000 197956
rect 177856 197872 177908 197878
rect 177856 197814 177908 197820
rect 177672 197804 177724 197810
rect 177672 197746 177724 197752
rect 177764 197668 177816 197674
rect 177764 197610 177816 197616
rect 177580 190256 177632 190262
rect 177580 190198 177632 190204
rect 177776 184822 177804 197610
rect 177960 190454 177988 197950
rect 178052 195498 178080 200602
rect 178130 199608 178186 199617
rect 178130 199543 178186 199552
rect 178040 195492 178092 195498
rect 178040 195434 178092 195440
rect 178040 192364 178092 192370
rect 178040 192306 178092 192312
rect 177868 190426 177988 190454
rect 177764 184816 177816 184822
rect 177764 184758 177816 184764
rect 177764 182844 177816 182850
rect 177764 182786 177816 182792
rect 177488 148912 177540 148918
rect 177488 148854 177540 148860
rect 176660 145512 176712 145518
rect 176660 145454 176712 145460
rect 176568 140548 176620 140554
rect 176568 140490 176620 140496
rect 176672 139890 176700 145454
rect 177776 144158 177804 182786
rect 177764 144152 177816 144158
rect 177764 144094 177816 144100
rect 177868 140486 177896 190426
rect 177948 187536 178000 187542
rect 177948 187478 178000 187484
rect 177960 146985 177988 187478
rect 177946 146976 178002 146985
rect 177946 146911 178002 146920
rect 177946 144256 178002 144265
rect 178052 144226 178080 192306
rect 178144 186250 178172 199543
rect 178236 198014 178264 200670
rect 179144 200592 179196 200598
rect 178406 200560 178462 200569
rect 179144 200534 179196 200540
rect 178406 200495 178462 200504
rect 178224 198008 178276 198014
rect 178224 197950 178276 197956
rect 178420 196858 178448 200495
rect 178592 200456 178644 200462
rect 178592 200398 178644 200404
rect 178408 196852 178460 196858
rect 178408 196794 178460 196800
rect 178604 196790 178632 200398
rect 179052 200320 179104 200326
rect 179052 200262 179104 200268
rect 179064 200122 179092 200262
rect 179052 200116 179104 200122
rect 179052 200058 179104 200064
rect 178592 196784 178644 196790
rect 178592 196726 178644 196732
rect 178224 196512 178276 196518
rect 178224 196454 178276 196460
rect 178236 188562 178264 196454
rect 178684 195084 178736 195090
rect 178684 195026 178736 195032
rect 178224 188556 178276 188562
rect 178224 188498 178276 188504
rect 178132 186244 178184 186250
rect 178132 186186 178184 186192
rect 178144 185978 178172 186186
rect 178132 185972 178184 185978
rect 178132 185914 178184 185920
rect 177946 144191 178002 144200
rect 178040 144220 178092 144226
rect 177856 140480 177908 140486
rect 177856 140422 177908 140428
rect 177960 139890 177988 144191
rect 178040 144162 178092 144168
rect 178696 140350 178724 195026
rect 178960 193792 179012 193798
rect 178960 193734 179012 193740
rect 178868 191548 178920 191554
rect 178868 191490 178920 191496
rect 178776 191412 178828 191418
rect 178776 191354 178828 191360
rect 178788 140457 178816 191354
rect 178880 146962 178908 191490
rect 178972 151814 179000 193734
rect 179156 192681 179184 200534
rect 179236 200116 179288 200122
rect 179236 200058 179288 200064
rect 179248 199374 179276 200058
rect 179326 200016 179382 200025
rect 181916 199986 181944 200670
rect 179326 199951 179382 199960
rect 181904 199980 181956 199986
rect 179236 199368 179288 199374
rect 179236 199310 179288 199316
rect 179340 196897 179368 199951
rect 181904 199922 181956 199928
rect 181812 199912 181864 199918
rect 181812 199854 181864 199860
rect 180984 199776 181036 199782
rect 180984 199718 181036 199724
rect 180708 199708 180760 199714
rect 180708 199650 180760 199656
rect 179512 199640 179564 199646
rect 179512 199582 179564 199588
rect 180340 199640 180392 199646
rect 180524 199640 180576 199646
rect 180392 199588 180524 199594
rect 180340 199582 180576 199588
rect 179418 197976 179474 197985
rect 179418 197911 179474 197920
rect 179326 196888 179382 196897
rect 179326 196823 179382 196832
rect 179142 192672 179198 192681
rect 179142 192607 179198 192616
rect 179432 185745 179460 197911
rect 179418 185736 179474 185745
rect 179418 185671 179474 185680
rect 178972 151786 179092 151814
rect 178880 146934 179000 146962
rect 178868 143200 178920 143206
rect 178868 143142 178920 143148
rect 178774 140448 178830 140457
rect 178774 140383 178830 140392
rect 178684 140344 178736 140350
rect 178684 140286 178736 140292
rect 178880 139890 178908 143142
rect 178972 140418 179000 146934
rect 179064 144226 179092 151786
rect 179420 145444 179472 145450
rect 179420 145386 179472 145392
rect 179052 144220 179104 144226
rect 179052 144162 179104 144168
rect 179328 142520 179380 142526
rect 179328 142462 179380 142468
rect 178960 140412 179012 140418
rect 178960 140354 179012 140360
rect 176672 139862 176916 139890
rect 177744 139862 177988 139890
rect 178572 139862 178908 139890
rect 179340 139890 179368 142462
rect 179432 140826 179460 145386
rect 179420 140820 179472 140826
rect 179420 140762 179472 140768
rect 179524 140049 179552 199582
rect 180352 199566 180564 199582
rect 180720 199102 180748 199650
rect 179696 199096 179748 199102
rect 179696 199038 179748 199044
rect 180708 199096 180760 199102
rect 180708 199038 180760 199044
rect 179708 180794 179736 199038
rect 180800 198212 180852 198218
rect 180800 198154 180852 198160
rect 180156 198076 180208 198082
rect 180156 198018 180208 198024
rect 180064 194948 180116 194954
rect 180064 194890 180116 194896
rect 179616 180766 179736 180794
rect 179616 140185 179644 180766
rect 179696 146396 179748 146402
rect 179696 146338 179748 146344
rect 179708 144906 179736 146338
rect 179696 144900 179748 144906
rect 179696 144842 179748 144848
rect 180076 141982 180104 194890
rect 180168 146402 180196 198018
rect 180708 198008 180760 198014
rect 180708 197950 180760 197956
rect 180720 196761 180748 197950
rect 180706 196752 180762 196761
rect 180706 196687 180762 196696
rect 180248 188216 180300 188222
rect 180248 188158 180300 188164
rect 180260 155242 180288 188158
rect 180706 186960 180762 186969
rect 180706 186895 180762 186904
rect 180248 155236 180300 155242
rect 180248 155178 180300 155184
rect 180156 146396 180208 146402
rect 180156 146338 180208 146344
rect 180064 141976 180116 141982
rect 180064 141918 180116 141924
rect 180720 141681 180748 186895
rect 180812 186046 180840 198154
rect 180800 186040 180852 186046
rect 180800 185982 180852 185988
rect 180800 145376 180852 145382
rect 180800 145318 180852 145324
rect 180706 141672 180762 141681
rect 180706 141607 180762 141616
rect 180812 140826 180840 145318
rect 180996 141409 181024 199718
rect 181824 199209 181852 199854
rect 182836 199345 182864 200670
rect 187606 200631 187662 200640
rect 182916 200116 182968 200122
rect 182916 200058 182968 200064
rect 182822 199336 182878 199345
rect 182822 199271 182878 199280
rect 181810 199200 181866 199209
rect 181810 199135 181866 199144
rect 181076 198212 181128 198218
rect 181076 198154 181128 198160
rect 181088 194449 181116 198154
rect 182270 198112 182326 198121
rect 182270 198047 182326 198056
rect 182180 197940 182232 197946
rect 182180 197882 182232 197888
rect 182088 197736 182140 197742
rect 182088 197678 182140 197684
rect 182100 194449 182128 197678
rect 181074 194440 181130 194449
rect 181074 194375 181130 194384
rect 182086 194440 182142 194449
rect 182086 194375 182142 194384
rect 181994 189680 182050 189689
rect 181994 189615 182050 189624
rect 181904 185496 181956 185502
rect 181904 185438 181956 185444
rect 181916 184958 181944 185438
rect 181904 184952 181956 184958
rect 181904 184894 181956 184900
rect 181352 143472 181404 143478
rect 181352 143414 181404 143420
rect 180982 141400 181038 141409
rect 180982 141335 181038 141344
rect 179880 140820 179932 140826
rect 179880 140762 179932 140768
rect 180800 140820 180852 140826
rect 180800 140762 180852 140768
rect 179602 140176 179658 140185
rect 179602 140111 179658 140120
rect 179510 140040 179566 140049
rect 179510 139975 179566 139984
rect 179892 139890 179920 140762
rect 181364 139890 181392 143414
rect 181916 141302 181944 184894
rect 181904 141296 181956 141302
rect 181904 141238 181956 141244
rect 181536 140820 181588 140826
rect 181536 140762 181588 140768
rect 179340 139862 179400 139890
rect 179892 139862 180228 139890
rect 181056 139862 181392 139890
rect 181548 139890 181576 140762
rect 182008 140185 182036 189615
rect 181994 140176 182050 140185
rect 181994 140111 182050 140120
rect 182100 140049 182128 194375
rect 182192 183326 182220 197882
rect 182284 183530 182312 198047
rect 182640 197600 182692 197606
rect 182640 197542 182692 197548
rect 182652 195809 182680 197542
rect 182638 195800 182694 195809
rect 182638 195735 182694 195744
rect 182272 183524 182324 183530
rect 182272 183466 182324 183472
rect 182180 183320 182232 183326
rect 182180 183262 182232 183268
rect 182836 140690 182864 199271
rect 182928 198762 182956 200058
rect 184940 199640 184992 199646
rect 184940 199582 184992 199588
rect 186228 199640 186280 199646
rect 186228 199582 186280 199588
rect 184952 199170 184980 199582
rect 185400 199232 185452 199238
rect 185400 199174 185452 199180
rect 184940 199164 184992 199170
rect 184940 199106 184992 199112
rect 182916 198756 182968 198762
rect 182916 198698 182968 198704
rect 185412 198558 185440 199174
rect 185584 198756 185636 198762
rect 185584 198698 185636 198704
rect 185400 198552 185452 198558
rect 185400 198494 185452 198500
rect 184940 198144 184992 198150
rect 184940 198086 184992 198092
rect 184204 192432 184256 192438
rect 184204 192374 184256 192380
rect 182916 191888 182968 191894
rect 182916 191830 182968 191836
rect 182824 140684 182876 140690
rect 182824 140626 182876 140632
rect 182928 140622 182956 191830
rect 183282 190088 183338 190097
rect 183282 190023 183338 190032
rect 183296 142154 183324 190023
rect 183376 189780 183428 189786
rect 183376 189722 183428 189728
rect 183204 142126 183324 142154
rect 183008 142112 183060 142118
rect 183008 142054 183060 142060
rect 182916 140616 182968 140622
rect 182916 140558 182968 140564
rect 182086 140040 182142 140049
rect 182086 139975 182142 139984
rect 183020 139890 183048 142054
rect 183100 140684 183152 140690
rect 183100 140626 183152 140632
rect 181548 139862 181884 139890
rect 182560 139862 183048 139890
rect 182560 139466 182588 139862
rect 182548 139460 182600 139466
rect 182548 139402 182600 139408
rect 183112 139369 183140 140626
rect 183204 139505 183232 142126
rect 183388 141817 183416 189722
rect 183468 143336 183520 143342
rect 183468 143278 183520 143284
rect 183374 141808 183430 141817
rect 183374 141743 183430 141752
rect 183480 139890 183508 143278
rect 184216 142154 184244 192374
rect 184952 191690 184980 198086
rect 184940 191684 184992 191690
rect 184940 191626 184992 191632
rect 184848 191480 184900 191486
rect 184848 191422 184900 191428
rect 184860 185570 184888 191422
rect 184952 191418 184980 191626
rect 184940 191412 184992 191418
rect 184940 191354 184992 191360
rect 184296 185564 184348 185570
rect 184296 185506 184348 185512
rect 184848 185564 184900 185570
rect 184848 185506 184900 185512
rect 184308 145897 184336 185506
rect 184848 178764 184900 178770
rect 184848 178706 184900 178712
rect 184294 145888 184350 145897
rect 184294 145823 184350 145832
rect 184664 143268 184716 143274
rect 184664 143210 184716 143216
rect 184032 142126 184244 142154
rect 183480 139862 183540 139890
rect 183190 139496 183246 139505
rect 183190 139431 183246 139440
rect 184032 139369 184060 142126
rect 184676 139890 184704 143210
rect 184860 141409 184888 178706
rect 185492 143404 185544 143410
rect 185492 143346 185544 143352
rect 184846 141400 184902 141409
rect 184846 141335 184902 141344
rect 185504 139890 185532 143346
rect 185596 142066 185624 198698
rect 185676 197260 185728 197266
rect 185676 197202 185728 197208
rect 185688 151814 185716 197202
rect 185768 194132 185820 194138
rect 185768 194074 185820 194080
rect 185780 190454 185808 194074
rect 186136 190460 186188 190466
rect 185780 190426 186136 190454
rect 186136 190402 186188 190408
rect 186042 184648 186098 184657
rect 186042 184583 186098 184592
rect 185688 151786 185808 151814
rect 185676 147280 185728 147286
rect 185676 147222 185728 147228
rect 185688 143070 185716 147222
rect 185676 143064 185728 143070
rect 185676 143006 185728 143012
rect 185596 142038 185716 142066
rect 185584 141908 185636 141914
rect 185584 141850 185636 141856
rect 185596 141166 185624 141850
rect 185584 141160 185636 141166
rect 185584 141102 185636 141108
rect 185688 139942 185716 142038
rect 184368 139862 184704 139890
rect 185196 139862 185532 139890
rect 185676 139936 185728 139942
rect 185676 139878 185728 139884
rect 185780 139874 185808 151786
rect 186056 146033 186084 184583
rect 186042 146024 186098 146033
rect 186042 145959 186098 145968
rect 185950 143304 186006 143313
rect 185950 143239 186006 143248
rect 185964 142497 185992 143239
rect 186044 142656 186096 142662
rect 186044 142598 186096 142604
rect 185950 142488 186006 142497
rect 185950 142423 186006 142432
rect 186056 140593 186084 142598
rect 186148 141953 186176 190402
rect 186240 142662 186268 199582
rect 186412 197872 186464 197878
rect 186412 197814 186464 197820
rect 186320 197804 186372 197810
rect 186320 197746 186372 197752
rect 186332 180334 186360 197746
rect 186320 180328 186372 180334
rect 186320 180270 186372 180276
rect 186332 180130 186360 180270
rect 186424 180266 186452 197814
rect 186504 197192 186556 197198
rect 186504 197134 186556 197140
rect 186516 196042 186544 197134
rect 186504 196036 186556 196042
rect 186504 195978 186556 195984
rect 187516 196036 187568 196042
rect 187516 195978 187568 195984
rect 186412 180260 186464 180266
rect 186412 180202 186464 180208
rect 186320 180124 186372 180130
rect 186320 180066 186372 180072
rect 186504 179172 186556 179178
rect 186504 179114 186556 179120
rect 186516 151814 186544 179114
rect 186596 179036 186648 179042
rect 186596 178978 186648 178984
rect 186332 151786 186544 151814
rect 186228 142656 186280 142662
rect 186228 142598 186280 142604
rect 186226 142488 186282 142497
rect 186226 142423 186282 142432
rect 186134 141944 186190 141953
rect 186134 141879 186190 141888
rect 186042 140584 186098 140593
rect 186042 140519 186098 140528
rect 186240 139890 186268 142423
rect 186332 140729 186360 151786
rect 186608 142154 186636 178978
rect 187528 151814 187556 195978
rect 187344 151786 187556 151814
rect 186870 143440 186926 143449
rect 186870 143375 186926 143384
rect 186516 142126 186636 142154
rect 186412 141364 186464 141370
rect 186412 141306 186464 141312
rect 186318 140720 186374 140729
rect 186318 140655 186374 140664
rect 186320 140548 186372 140554
rect 186320 140490 186372 140496
rect 186332 140078 186360 140490
rect 186320 140072 186372 140078
rect 186320 140014 186372 140020
rect 185768 139868 185820 139874
rect 186024 139862 186268 139890
rect 185768 139810 185820 139816
rect 130842 139360 130898 139369
rect 130672 139318 130842 139346
rect 129186 139295 129242 139304
rect 130842 139295 130898 139304
rect 146666 139360 146722 139369
rect 146666 139295 146722 139304
rect 170678 139360 170734 139369
rect 170678 139295 170734 139304
rect 176474 139360 176530 139369
rect 176474 139295 176530 139304
rect 183098 139360 183154 139369
rect 183098 139295 183154 139304
rect 184018 139360 184074 139369
rect 186424 139330 186452 141306
rect 186516 139505 186544 142126
rect 186884 140162 186912 143375
rect 187344 140690 187372 151786
rect 187620 145466 187648 200631
rect 188988 200184 189040 200190
rect 188988 200126 189040 200132
rect 188896 198960 188948 198966
rect 188896 198902 188948 198908
rect 187792 190188 187844 190194
rect 187792 190130 187844 190136
rect 187700 147008 187752 147014
rect 187700 146950 187752 146956
rect 187712 146334 187740 146950
rect 187700 146328 187752 146334
rect 187700 146270 187752 146276
rect 187698 145616 187754 145625
rect 187698 145551 187754 145560
rect 187436 145438 187648 145466
rect 187436 142254 187464 145438
rect 187608 142520 187660 142526
rect 187608 142462 187660 142468
rect 187424 142248 187476 142254
rect 187424 142190 187476 142196
rect 187332 140684 187384 140690
rect 187332 140626 187384 140632
rect 186838 140134 186912 140162
rect 186838 139876 186866 140134
rect 187332 140072 187384 140078
rect 187332 140014 187384 140020
rect 187344 139641 187372 140014
rect 187436 139890 187464 142190
rect 187620 141914 187648 142462
rect 187608 141908 187660 141914
rect 187608 141850 187660 141856
rect 187712 140826 187740 145551
rect 187700 140820 187752 140826
rect 187700 140762 187752 140768
rect 187804 140486 187832 190130
rect 188620 182912 188672 182918
rect 188620 182854 188672 182860
rect 188342 179344 188398 179353
rect 188342 179279 188398 179288
rect 188356 151814 188384 179279
rect 187988 151786 188384 151814
rect 187792 140480 187844 140486
rect 187792 140422 187844 140428
rect 187436 139862 187680 139890
rect 187330 139632 187386 139641
rect 187330 139567 187386 139576
rect 187988 139505 188016 151786
rect 188160 147008 188212 147014
rect 188160 146950 188212 146956
rect 186502 139496 186558 139505
rect 186502 139431 186558 139440
rect 187974 139496 188030 139505
rect 187974 139431 188030 139440
rect 188172 139398 188200 146950
rect 188252 140820 188304 140826
rect 188252 140762 188304 140768
rect 188264 139890 188292 140762
rect 188264 139862 188508 139890
rect 188160 139392 188212 139398
rect 188160 139334 188212 139340
rect 184018 139295 184074 139304
rect 186412 139324 186464 139330
rect 123208 139266 123260 139272
rect 186412 139266 186464 139272
rect 131762 80744 131818 80753
rect 123772 80714 123984 80730
rect 123760 80708 123996 80714
rect 123812 80702 123944 80708
rect 123760 80650 123812 80656
rect 123944 80650 123996 80656
rect 128912 80708 128964 80714
rect 128912 80650 128964 80656
rect 131580 80708 131632 80714
rect 131580 80650 131632 80656
rect 131672 80708 131724 80714
rect 132222 80744 132278 80753
rect 131762 80679 131818 80688
rect 131948 80708 132000 80714
rect 131672 80650 131724 80656
rect 123482 80608 123538 80617
rect 123482 80543 123538 80552
rect 122378 80336 122434 80345
rect 122378 80271 122434 80280
rect 122392 74497 122420 80271
rect 122378 74488 122434 74497
rect 122378 74423 122434 74432
rect 123496 71602 123524 80543
rect 124496 80504 124548 80510
rect 124496 80446 124548 80452
rect 124508 75886 124536 80446
rect 128176 80368 128228 80374
rect 128176 80310 128228 80316
rect 126334 79928 126390 79937
rect 126334 79863 126390 79872
rect 126244 79620 126296 79626
rect 126244 79562 126296 79568
rect 124496 75880 124548 75886
rect 124496 75822 124548 75828
rect 126256 72894 126284 79562
rect 126348 78033 126376 79863
rect 127624 79552 127676 79558
rect 127624 79494 127676 79500
rect 126334 78024 126390 78033
rect 126334 77959 126390 77968
rect 126336 75948 126388 75954
rect 126336 75890 126388 75896
rect 126348 75274 126376 75890
rect 126336 75268 126388 75274
rect 126336 75210 126388 75216
rect 126244 72888 126296 72894
rect 126244 72830 126296 72836
rect 124220 72480 124272 72486
rect 124220 72422 124272 72428
rect 123484 71596 123536 71602
rect 123484 71538 123536 71544
rect 122104 48272 122156 48278
rect 122104 48214 122156 48220
rect 124232 16574 124260 72422
rect 127636 70786 127664 79494
rect 128188 77926 128216 80310
rect 128176 77920 128228 77926
rect 128176 77862 128228 77868
rect 128924 74798 128952 80650
rect 131592 80442 131620 80650
rect 131684 80578 131712 80650
rect 131672 80572 131724 80578
rect 131672 80514 131724 80520
rect 131580 80436 131632 80442
rect 131580 80378 131632 80384
rect 129924 80232 129976 80238
rect 129924 80174 129976 80180
rect 129188 78940 129240 78946
rect 129188 78882 129240 78888
rect 129200 78305 129228 78882
rect 129186 78296 129242 78305
rect 129186 78231 129242 78240
rect 129936 78198 129964 80174
rect 131776 80170 131804 80679
rect 131948 80650 132000 80656
rect 132132 80708 132184 80714
rect 132222 80679 132278 80688
rect 177856 80708 177908 80714
rect 132132 80650 132184 80656
rect 131960 80442 131988 80650
rect 132144 80510 132172 80650
rect 132236 80646 132264 80679
rect 177856 80650 177908 80656
rect 178040 80708 178092 80714
rect 178040 80650 178092 80656
rect 178408 80708 178460 80714
rect 178408 80650 178460 80656
rect 132224 80640 132276 80646
rect 177762 80608 177818 80617
rect 132224 80582 132276 80588
rect 177652 80566 177762 80594
rect 177762 80543 177818 80552
rect 132132 80504 132184 80510
rect 132132 80446 132184 80452
rect 177868 80442 177896 80650
rect 178052 80578 178080 80650
rect 178040 80572 178092 80578
rect 178040 80514 178092 80520
rect 131948 80436 132000 80442
rect 131948 80378 132000 80384
rect 177856 80436 177908 80442
rect 177856 80378 177908 80384
rect 177764 80368 177816 80374
rect 131946 80336 132002 80345
rect 177764 80310 177816 80316
rect 131946 80271 132002 80280
rect 131856 80232 131908 80238
rect 131856 80174 131908 80180
rect 131764 80164 131816 80170
rect 131764 80106 131816 80112
rect 130108 80096 130160 80102
rect 130108 80038 130160 80044
rect 131672 80096 131724 80102
rect 131868 80073 131896 80174
rect 131672 80038 131724 80044
rect 131854 80064 131910 80073
rect 130120 79490 130148 80038
rect 131684 79966 131712 80038
rect 131960 80034 131988 80271
rect 132052 80158 132388 80186
rect 131854 79999 131910 80008
rect 131948 80028 132000 80034
rect 131948 79970 132000 79976
rect 131672 79960 131724 79966
rect 131672 79902 131724 79908
rect 131580 79824 131632 79830
rect 131580 79766 131632 79772
rect 130108 79484 130160 79490
rect 130108 79426 130160 79432
rect 131028 78804 131080 78810
rect 131028 78746 131080 78752
rect 130384 78328 130436 78334
rect 130384 78270 130436 78276
rect 129924 78192 129976 78198
rect 129924 78134 129976 78140
rect 128912 74792 128964 74798
rect 128912 74734 128964 74740
rect 127624 70780 127676 70786
rect 127624 70722 127676 70728
rect 126244 69760 126296 69766
rect 126244 69702 126296 69708
rect 126256 40050 126284 69702
rect 130396 66910 130424 78270
rect 131040 78130 131068 78746
rect 131592 78402 131620 79766
rect 132052 78674 132080 80158
rect 132132 79960 132184 79966
rect 132132 79902 132184 79908
rect 132144 79801 132172 79902
rect 132130 79792 132186 79801
rect 132466 79744 132494 80036
rect 132558 79966 132586 80036
rect 132650 79966 132678 80036
rect 132546 79960 132598 79966
rect 132546 79902 132598 79908
rect 132638 79960 132690 79966
rect 132638 79902 132690 79908
rect 132130 79727 132186 79736
rect 132420 79716 132494 79744
rect 132040 78668 132092 78674
rect 132040 78610 132092 78616
rect 132132 78668 132184 78674
rect 132132 78610 132184 78616
rect 131580 78396 131632 78402
rect 131580 78338 131632 78344
rect 132144 78334 132172 78610
rect 132132 78328 132184 78334
rect 132132 78270 132184 78276
rect 131028 78124 131080 78130
rect 131028 78066 131080 78072
rect 132040 78124 132092 78130
rect 132040 78066 132092 78072
rect 131856 76492 131908 76498
rect 131856 76434 131908 76440
rect 130844 75812 130896 75818
rect 130844 75754 130896 75760
rect 130856 71262 130884 75754
rect 131764 73500 131816 73506
rect 131764 73442 131816 73448
rect 130844 71256 130896 71262
rect 130844 71198 130896 71204
rect 129740 66904 129792 66910
rect 129740 66846 129792 66852
rect 130384 66904 130436 66910
rect 130384 66846 130436 66852
rect 129752 66706 129780 66846
rect 129740 66700 129792 66706
rect 129740 66642 129792 66648
rect 126244 40044 126296 40050
rect 126244 39986 126296 39992
rect 120092 16546 120672 16574
rect 124232 16546 124536 16574
rect 117228 3596 117280 3602
rect 117228 3538 117280 3544
rect 117240 480 117268 3538
rect 113334 354 113446 480
rect 113192 326 113446 354
rect 113334 -960 113446 326
rect 117198 -960 117310 480
rect 120644 354 120672 16546
rect 121062 354 121174 480
rect 120644 326 121174 354
rect 124508 354 124536 16546
rect 129752 12442 129780 66642
rect 131120 63164 131172 63170
rect 131120 63106 131172 63112
rect 131132 62490 131160 63106
rect 131120 62484 131172 62490
rect 131120 62426 131172 62432
rect 131132 16590 131160 62426
rect 131776 44130 131804 73442
rect 131868 62490 131896 76434
rect 132052 75954 132080 78066
rect 132040 75948 132092 75954
rect 132040 75890 132092 75896
rect 132420 70854 132448 79716
rect 132742 79676 132770 80036
rect 132834 79778 132862 80036
rect 132926 79966 132954 80036
rect 133018 79966 133046 80036
rect 132914 79960 132966 79966
rect 132914 79902 132966 79908
rect 133006 79960 133058 79966
rect 133110 79937 133138 80036
rect 133202 79966 133230 80036
rect 133190 79960 133242 79966
rect 133006 79902 133058 79908
rect 133096 79928 133152 79937
rect 133190 79902 133242 79908
rect 133096 79863 133152 79872
rect 133144 79824 133196 79830
rect 132834 79762 132908 79778
rect 133294 79812 133322 80036
rect 133386 79966 133414 80036
rect 133374 79960 133426 79966
rect 133478 79937 133506 80036
rect 133374 79902 133426 79908
rect 133464 79928 133520 79937
rect 133464 79863 133520 79872
rect 133570 79812 133598 80036
rect 133662 79937 133690 80036
rect 133648 79928 133704 79937
rect 133648 79863 133704 79872
rect 133754 79812 133782 80036
rect 133846 79966 133874 80036
rect 133938 79966 133966 80036
rect 133834 79960 133886 79966
rect 133834 79902 133886 79908
rect 133926 79960 133978 79966
rect 134030 79937 134058 80036
rect 133926 79902 133978 79908
rect 134016 79928 134072 79937
rect 134016 79863 134072 79872
rect 134122 79812 134150 80036
rect 133294 79784 133368 79812
rect 133144 79766 133196 79772
rect 132834 79756 132920 79762
rect 132834 79750 132868 79756
rect 132868 79698 132920 79704
rect 133052 79688 133104 79694
rect 132742 79648 132816 79676
rect 132408 70848 132460 70854
rect 132408 70790 132460 70796
rect 132500 68332 132552 68338
rect 132500 68274 132552 68280
rect 131856 62484 131908 62490
rect 131856 62426 131908 62432
rect 131764 44124 131816 44130
rect 131764 44066 131816 44072
rect 131120 16584 131172 16590
rect 131120 16526 131172 16532
rect 129740 12436 129792 12442
rect 129740 12378 129792 12384
rect 128820 3528 128872 3534
rect 128820 3470 128872 3476
rect 128832 480 128860 3470
rect 124926 354 125038 480
rect 124508 326 125038 354
rect 121062 -960 121174 326
rect 124926 -960 125038 326
rect 128790 -960 128902 480
rect 132512 354 132540 68274
rect 132788 67153 132816 79648
rect 133156 79665 133184 79766
rect 133052 79630 133104 79636
rect 133142 79656 133198 79665
rect 132960 79620 133012 79626
rect 132960 79562 133012 79568
rect 132866 78432 132922 78441
rect 132866 78367 132922 78376
rect 132880 78198 132908 78367
rect 132868 78192 132920 78198
rect 132868 78134 132920 78140
rect 132774 67144 132830 67153
rect 132774 67079 132830 67088
rect 132972 64258 133000 79562
rect 133064 78577 133092 79630
rect 133142 79591 133198 79600
rect 133142 78704 133198 78713
rect 133142 78639 133198 78648
rect 133050 78568 133106 78577
rect 133050 78503 133106 78512
rect 133052 75268 133104 75274
rect 133052 75210 133104 75216
rect 133064 68490 133092 75210
rect 133156 72350 133184 78639
rect 133236 76832 133288 76838
rect 133236 76774 133288 76780
rect 133248 75154 133276 76774
rect 133340 75818 133368 79784
rect 133418 79792 133474 79801
rect 133570 79784 133644 79812
rect 133418 79727 133474 79736
rect 133328 75812 133380 75818
rect 133328 75754 133380 75760
rect 133326 75168 133382 75177
rect 133248 75126 133326 75154
rect 133326 75103 133382 75112
rect 133144 72344 133196 72350
rect 133144 72286 133196 72292
rect 133144 72208 133196 72214
rect 133144 72150 133196 72156
rect 133156 68678 133184 72150
rect 133144 68672 133196 68678
rect 133144 68614 133196 68620
rect 133064 68462 133276 68490
rect 133144 66020 133196 66026
rect 133144 65962 133196 65968
rect 132960 64252 133012 64258
rect 132960 64194 133012 64200
rect 133156 42158 133184 65962
rect 133248 64666 133276 68462
rect 133236 64660 133288 64666
rect 133236 64602 133288 64608
rect 133248 51746 133276 64602
rect 133340 64258 133368 75103
rect 133432 66026 133460 79727
rect 133616 72214 133644 79784
rect 133708 79784 133782 79812
rect 133984 79801 134150 79812
rect 133970 79792 134150 79801
rect 133708 79744 133736 79784
rect 133880 79756 133932 79762
rect 133708 79716 133828 79744
rect 133696 79620 133748 79626
rect 133696 79562 133748 79568
rect 133708 73154 133736 79562
rect 133800 75274 133828 79716
rect 134026 79784 134150 79792
rect 134214 79744 134242 80036
rect 134306 79898 134334 80036
rect 134398 79971 134426 80036
rect 134384 79962 134440 79971
rect 134294 79892 134346 79898
rect 134384 79897 134440 79906
rect 134294 79834 134346 79840
rect 133970 79727 134026 79736
rect 133880 79698 133932 79704
rect 134168 79716 134242 79744
rect 134340 79756 134392 79762
rect 133788 75268 133840 75274
rect 133788 75210 133840 75216
rect 133708 73126 133828 73154
rect 133604 72208 133656 72214
rect 133604 72150 133656 72156
rect 133800 69970 133828 73126
rect 133892 72282 133920 79698
rect 134062 79656 134118 79665
rect 134062 79591 134118 79600
rect 134076 77994 134104 79591
rect 134064 77988 134116 77994
rect 134064 77930 134116 77936
rect 134076 76158 134104 77930
rect 134064 76152 134116 76158
rect 134064 76094 134116 76100
rect 133880 72276 133932 72282
rect 133880 72218 133932 72224
rect 133788 69964 133840 69970
rect 133788 69906 133840 69912
rect 133420 66020 133472 66026
rect 133420 65962 133472 65968
rect 134168 65822 134196 79716
rect 134490 79744 134518 80036
rect 134582 79898 134610 80036
rect 134674 79898 134702 80036
rect 134766 79971 134794 80036
rect 134752 79962 134808 79971
rect 134570 79892 134622 79898
rect 134570 79834 134622 79840
rect 134662 79892 134714 79898
rect 134752 79897 134808 79906
rect 134858 79898 134886 80036
rect 134950 79898 134978 80036
rect 135042 79966 135070 80036
rect 135134 79966 135162 80036
rect 135226 79966 135254 80036
rect 135318 79966 135346 80036
rect 135030 79960 135082 79966
rect 135030 79902 135082 79908
rect 135122 79960 135174 79966
rect 135122 79902 135174 79908
rect 135214 79960 135266 79966
rect 135214 79902 135266 79908
rect 135306 79960 135358 79966
rect 135306 79902 135358 79908
rect 134662 79834 134714 79840
rect 134846 79892 134898 79898
rect 134846 79834 134898 79840
rect 134938 79892 134990 79898
rect 134938 79834 134990 79840
rect 135168 79824 135220 79830
rect 134614 79792 134670 79801
rect 135168 79766 135220 79772
rect 134490 79716 134564 79744
rect 134614 79727 134616 79736
rect 134340 79698 134392 79704
rect 134248 79620 134300 79626
rect 134248 79562 134300 79568
rect 134260 70394 134288 79562
rect 134352 76838 134380 79698
rect 134432 79620 134484 79626
rect 134432 79562 134484 79568
rect 134340 76832 134392 76838
rect 134340 76774 134392 76780
rect 134260 70366 134380 70394
rect 134352 66094 134380 70366
rect 134340 66088 134392 66094
rect 134340 66030 134392 66036
rect 134156 65816 134208 65822
rect 134156 65758 134208 65764
rect 134352 64874 134380 66030
rect 134260 64846 134380 64874
rect 133328 64252 133380 64258
rect 133328 64194 133380 64200
rect 133880 63912 133932 63918
rect 133880 63854 133932 63860
rect 133236 51740 133288 51746
rect 133236 51682 133288 51688
rect 133144 42152 133196 42158
rect 133144 42094 133196 42100
rect 133892 37262 133920 63854
rect 134260 60042 134288 64846
rect 134444 64530 134472 79562
rect 134536 78130 134564 79716
rect 134668 79727 134670 79736
rect 135076 79756 135128 79762
rect 134616 79698 134668 79704
rect 135076 79698 135128 79704
rect 134708 79688 134760 79694
rect 134614 79656 134670 79665
rect 134708 79630 134760 79636
rect 134614 79591 134670 79600
rect 134524 78124 134576 78130
rect 134524 78066 134576 78072
rect 134524 76152 134576 76158
rect 134524 76094 134576 76100
rect 134432 64524 134484 64530
rect 134432 64466 134484 64472
rect 134444 63918 134472 64466
rect 134432 63912 134484 63918
rect 134432 63854 134484 63860
rect 134248 60036 134300 60042
rect 134248 59978 134300 59984
rect 133880 37256 133932 37262
rect 133880 37198 133932 37204
rect 134536 13122 134564 76094
rect 134628 64598 134656 79591
rect 134720 65346 134748 79630
rect 134892 79552 134944 79558
rect 134892 79494 134944 79500
rect 134904 67114 134932 79494
rect 134984 79416 135036 79422
rect 134984 79358 135036 79364
rect 134996 78577 135024 79358
rect 134982 78568 135038 78577
rect 134982 78503 135038 78512
rect 134982 78024 135038 78033
rect 134982 77959 135038 77968
rect 134996 77790 135024 77959
rect 134984 77784 135036 77790
rect 134984 77726 135036 77732
rect 134984 76832 135036 76838
rect 134984 76774 135036 76780
rect 134892 67108 134944 67114
rect 134892 67050 134944 67056
rect 134708 65340 134760 65346
rect 134708 65282 134760 65288
rect 134616 64592 134668 64598
rect 134616 64534 134668 64540
rect 134524 13116 134576 13122
rect 134524 13058 134576 13064
rect 134628 8974 134656 64534
rect 134720 24138 134748 65282
rect 134904 58818 134932 67050
rect 134996 65278 135024 76774
rect 135088 76537 135116 79698
rect 135074 76528 135130 76537
rect 135074 76463 135130 76472
rect 135180 73642 135208 79766
rect 135260 79756 135312 79762
rect 135260 79698 135312 79704
rect 135272 77897 135300 79698
rect 135410 79676 135438 80036
rect 135502 79898 135530 80036
rect 135594 79971 135622 80036
rect 135580 79962 135636 79971
rect 135490 79892 135542 79898
rect 135580 79897 135636 79906
rect 135490 79834 135542 79840
rect 135686 79812 135714 80036
rect 135640 79784 135714 79812
rect 135536 79756 135588 79762
rect 135536 79698 135588 79704
rect 135410 79648 135484 79676
rect 135352 79416 135404 79422
rect 135352 79358 135404 79364
rect 135364 79082 135392 79358
rect 135352 79076 135404 79082
rect 135352 79018 135404 79024
rect 135352 78736 135404 78742
rect 135352 78678 135404 78684
rect 135258 77888 135314 77897
rect 135258 77823 135314 77832
rect 135364 74534 135392 78678
rect 135456 75698 135484 79648
rect 135548 76265 135576 79698
rect 135640 77926 135668 79784
rect 135778 79744 135806 80036
rect 135870 79971 135898 80036
rect 135856 79962 135912 79971
rect 135856 79897 135912 79906
rect 135962 79898 135990 80036
rect 136054 79898 136082 80036
rect 136146 79937 136174 80036
rect 136238 79966 136266 80036
rect 136226 79960 136278 79966
rect 136132 79928 136188 79937
rect 135950 79892 136002 79898
rect 135950 79834 136002 79840
rect 136042 79892 136094 79898
rect 136226 79902 136278 79908
rect 136330 79898 136358 80036
rect 136132 79863 136188 79872
rect 136318 79892 136370 79898
rect 136042 79834 136094 79840
rect 136318 79834 136370 79840
rect 136422 79812 136450 80036
rect 136514 79966 136542 80036
rect 136502 79960 136554 79966
rect 136502 79902 136554 79908
rect 136606 79898 136634 80036
rect 136698 79898 136726 80036
rect 136790 79971 136818 80036
rect 136776 79962 136832 79971
rect 136594 79892 136646 79898
rect 136594 79834 136646 79840
rect 136686 79892 136738 79898
rect 136776 79897 136832 79906
rect 136882 79898 136910 80036
rect 136686 79834 136738 79840
rect 136870 79892 136922 79898
rect 136870 79834 136922 79840
rect 136422 79784 136496 79812
rect 135732 79716 135806 79744
rect 136088 79756 136140 79762
rect 135732 78169 135760 79716
rect 136088 79698 136140 79704
rect 136180 79756 136232 79762
rect 136180 79698 136232 79704
rect 135996 79688 136048 79694
rect 135996 79630 136048 79636
rect 135812 79620 135864 79626
rect 135812 79562 135864 79568
rect 135824 78742 135852 79562
rect 135812 78736 135864 78742
rect 135812 78678 135864 78684
rect 136008 78248 136036 79630
rect 135824 78220 136036 78248
rect 135718 78160 135774 78169
rect 135718 78095 135774 78104
rect 135628 77920 135680 77926
rect 135628 77862 135680 77868
rect 135720 77852 135772 77858
rect 135720 77794 135772 77800
rect 135534 76256 135590 76265
rect 135534 76191 135590 76200
rect 135732 75886 135760 77794
rect 135720 75880 135772 75886
rect 135720 75822 135772 75828
rect 135456 75670 135760 75698
rect 135536 75268 135588 75274
rect 135536 75210 135588 75216
rect 135364 74506 135484 74534
rect 135168 73636 135220 73642
rect 135168 73578 135220 73584
rect 135456 65618 135484 74506
rect 135548 68270 135576 75210
rect 135628 75132 135680 75138
rect 135628 75074 135680 75080
rect 135536 68264 135588 68270
rect 135536 68206 135588 68212
rect 135444 65612 135496 65618
rect 135444 65554 135496 65560
rect 134984 65272 135036 65278
rect 134984 65214 135036 65220
rect 134892 58812 134944 58818
rect 134892 58754 134944 58760
rect 134708 24132 134760 24138
rect 134708 24074 134760 24080
rect 134616 8968 134668 8974
rect 134616 8910 134668 8916
rect 135456 3466 135484 65554
rect 135640 64870 135668 75074
rect 135732 70394 135760 75670
rect 135824 74050 135852 78220
rect 135904 78124 135956 78130
rect 135904 78066 135956 78072
rect 135812 74044 135864 74050
rect 135812 73986 135864 73992
rect 135732 70366 135852 70394
rect 135916 70378 135944 78066
rect 136100 77466 136128 79698
rect 136192 79665 136220 79698
rect 136364 79688 136416 79694
rect 136178 79656 136234 79665
rect 136364 79630 136416 79636
rect 136178 79591 136234 79600
rect 136272 79552 136324 79558
rect 136272 79494 136324 79500
rect 136008 77438 136128 77466
rect 136008 75274 136036 77438
rect 136088 77308 136140 77314
rect 136088 77250 136140 77256
rect 135996 75268 136048 75274
rect 135996 75210 136048 75216
rect 135824 68490 135852 70366
rect 135904 70372 135956 70378
rect 135904 70314 135956 70320
rect 135824 68462 136036 68490
rect 136008 66230 136036 68462
rect 135996 66224 136048 66230
rect 135996 66166 136048 66172
rect 135904 65816 135956 65822
rect 135904 65758 135956 65764
rect 135628 64864 135680 64870
rect 135628 64806 135680 64812
rect 135444 3460 135496 3466
rect 135444 3402 135496 3408
rect 135916 3330 135944 65758
rect 136008 51066 136036 66166
rect 136100 64734 136128 77250
rect 136284 76566 136312 79494
rect 136272 76560 136324 76566
rect 136272 76502 136324 76508
rect 136376 70394 136404 79630
rect 136468 79422 136496 79784
rect 136822 79792 136878 79801
rect 136744 79750 136822 79778
rect 136548 79688 136600 79694
rect 136548 79630 136600 79636
rect 136640 79688 136692 79694
rect 136640 79630 136692 79636
rect 136456 79416 136508 79422
rect 136456 79358 136508 79364
rect 136456 79076 136508 79082
rect 136456 79018 136508 79024
rect 136468 78606 136496 79018
rect 136456 78600 136508 78606
rect 136456 78542 136508 78548
rect 136560 75138 136588 79630
rect 136652 78470 136680 79630
rect 136744 79082 136772 79750
rect 136974 79744 137002 80036
rect 137066 79966 137094 80036
rect 137054 79960 137106 79966
rect 137158 79937 137186 80036
rect 137054 79902 137106 79908
rect 137144 79928 137200 79937
rect 137250 79898 137278 80036
rect 137342 79971 137370 80036
rect 137328 79962 137384 79971
rect 137144 79863 137200 79872
rect 137238 79892 137290 79898
rect 137328 79897 137384 79906
rect 137434 79898 137462 80036
rect 137526 79966 137554 80036
rect 137618 79966 137646 80036
rect 137710 79966 137738 80036
rect 137514 79960 137566 79966
rect 137514 79902 137566 79908
rect 137606 79960 137658 79966
rect 137606 79902 137658 79908
rect 137698 79960 137750 79966
rect 137698 79902 137750 79908
rect 137238 79834 137290 79840
rect 137422 79892 137474 79898
rect 137422 79834 137474 79840
rect 137560 79824 137612 79830
rect 137190 79792 137246 79801
rect 136822 79727 136878 79736
rect 136928 79716 137002 79744
rect 137100 79756 137152 79762
rect 136824 79688 136876 79694
rect 136822 79656 136824 79665
rect 136876 79656 136878 79665
rect 136822 79591 136878 79600
rect 136732 79076 136784 79082
rect 136732 79018 136784 79024
rect 136732 78736 136784 78742
rect 136732 78678 136784 78684
rect 136640 78464 136692 78470
rect 136640 78406 136692 78412
rect 136640 78328 136692 78334
rect 136640 78270 136692 78276
rect 136652 76945 136680 78270
rect 136638 76936 136694 76945
rect 136638 76871 136694 76880
rect 136548 75132 136600 75138
rect 136548 75074 136600 75080
rect 136376 70366 136496 70394
rect 136468 69018 136496 70366
rect 136456 69012 136508 69018
rect 136456 68954 136508 68960
rect 136640 67516 136692 67522
rect 136640 67458 136692 67464
rect 136652 67114 136680 67458
rect 136744 67182 136772 78678
rect 136824 77716 136876 77722
rect 136824 77658 136876 77664
rect 136836 76702 136864 77658
rect 136824 76696 136876 76702
rect 136824 76638 136876 76644
rect 136824 76560 136876 76566
rect 136824 76502 136876 76508
rect 136836 67522 136864 76502
rect 136824 67516 136876 67522
rect 136824 67458 136876 67464
rect 136836 67318 136864 67458
rect 136824 67312 136876 67318
rect 136824 67254 136876 67260
rect 136928 67250 136956 79716
rect 137560 79766 137612 79772
rect 137190 79727 137246 79736
rect 137100 79698 137152 79704
rect 137008 79620 137060 79626
rect 137008 79562 137060 79568
rect 137020 78742 137048 79562
rect 137008 78736 137060 78742
rect 137008 78678 137060 78684
rect 137008 77920 137060 77926
rect 137008 77862 137060 77868
rect 137020 76809 137048 77862
rect 137006 76800 137062 76809
rect 137006 76735 137062 76744
rect 137112 75313 137140 79698
rect 137204 77353 137232 79727
rect 137466 79656 137522 79665
rect 137284 79620 137336 79626
rect 137284 79562 137336 79568
rect 137376 79620 137428 79626
rect 137466 79591 137522 79600
rect 137376 79562 137428 79568
rect 137190 77344 137246 77353
rect 137190 77279 137246 77288
rect 137192 76084 137244 76090
rect 137192 76026 137244 76032
rect 137098 75304 137154 75313
rect 137098 75239 137154 75248
rect 137204 71194 137232 76026
rect 137296 74662 137324 79562
rect 137388 79257 137416 79562
rect 137374 79248 137430 79257
rect 137374 79183 137430 79192
rect 137480 78062 137508 79591
rect 137572 79393 137600 79766
rect 137652 79756 137704 79762
rect 137802 79744 137830 80036
rect 137652 79698 137704 79704
rect 137756 79716 137830 79744
rect 137558 79384 137614 79393
rect 137558 79319 137614 79328
rect 137468 78056 137520 78062
rect 137468 77998 137520 78004
rect 137664 76566 137692 79698
rect 137652 76560 137704 76566
rect 137652 76502 137704 76508
rect 137284 74656 137336 74662
rect 137284 74598 137336 74604
rect 137756 73506 137784 79716
rect 137894 79676 137922 80036
rect 137986 79966 138014 80036
rect 138078 79971 138106 80036
rect 137974 79960 138026 79966
rect 137974 79902 138026 79908
rect 138064 79962 138120 79971
rect 138170 79966 138198 80036
rect 138262 79966 138290 80036
rect 138064 79897 138120 79906
rect 138158 79960 138210 79966
rect 138158 79902 138210 79908
rect 138250 79960 138302 79966
rect 138250 79902 138302 79908
rect 138020 79824 138072 79830
rect 138354 79778 138382 80036
rect 138446 79937 138474 80036
rect 138432 79928 138488 79937
rect 138432 79863 138488 79872
rect 138020 79766 138072 79772
rect 137848 79648 137922 79676
rect 137744 73500 137796 73506
rect 137744 73442 137796 73448
rect 137192 71188 137244 71194
rect 137192 71130 137244 71136
rect 137848 70394 137876 79648
rect 138032 76362 138060 79766
rect 138308 79750 138382 79778
rect 138112 79688 138164 79694
rect 138112 79630 138164 79636
rect 138124 78033 138152 79630
rect 138308 79529 138336 79750
rect 138388 79688 138440 79694
rect 138538 79642 138566 80036
rect 138630 79744 138658 80036
rect 138722 79898 138750 80036
rect 138814 79898 138842 80036
rect 138906 79971 138934 80036
rect 138892 79962 138948 79971
rect 138710 79892 138762 79898
rect 138710 79834 138762 79840
rect 138802 79892 138854 79898
rect 138892 79897 138948 79906
rect 138998 79898 139026 80036
rect 139090 79898 139118 80036
rect 139182 79966 139210 80036
rect 139170 79960 139222 79966
rect 139170 79902 139222 79908
rect 138802 79834 138854 79840
rect 138986 79892 139038 79898
rect 138986 79834 139038 79840
rect 139078 79892 139130 79898
rect 139078 79834 139130 79840
rect 139274 79812 139302 80036
rect 139228 79784 139302 79812
rect 138940 79756 138992 79762
rect 138630 79716 138704 79744
rect 138388 79630 138440 79636
rect 138294 79520 138350 79529
rect 138294 79455 138350 79464
rect 138400 78198 138428 79630
rect 138492 79614 138566 79642
rect 138388 78192 138440 78198
rect 138388 78134 138440 78140
rect 138110 78024 138166 78033
rect 138110 77959 138166 77968
rect 138492 76566 138520 79614
rect 138572 79552 138624 79558
rect 138572 79494 138624 79500
rect 138296 76560 138348 76566
rect 138480 76560 138532 76566
rect 138296 76502 138348 76508
rect 138386 76528 138442 76537
rect 138020 76356 138072 76362
rect 138020 76298 138072 76304
rect 138204 75880 138256 75886
rect 138204 75822 138256 75828
rect 137928 75812 137980 75818
rect 137928 75754 137980 75760
rect 137940 74798 137968 75754
rect 138216 75342 138244 75822
rect 138204 75336 138256 75342
rect 138204 75278 138256 75284
rect 137928 74792 137980 74798
rect 137928 74734 137980 74740
rect 138204 73772 138256 73778
rect 138204 73714 138256 73720
rect 137112 70366 137876 70394
rect 136916 67244 136968 67250
rect 136916 67186 136968 67192
rect 136732 67176 136784 67182
rect 136732 67118 136784 67124
rect 136640 67108 136692 67114
rect 136640 67050 136692 67056
rect 136088 64728 136140 64734
rect 136088 64670 136140 64676
rect 137112 64054 137140 70366
rect 137284 67516 137336 67522
rect 137284 67458 137336 67464
rect 137100 64048 137152 64054
rect 137100 63990 137152 63996
rect 137112 63578 137140 63990
rect 137100 63572 137152 63578
rect 137100 63514 137152 63520
rect 135996 51060 136048 51066
rect 135996 51002 136048 51008
rect 137296 37942 137324 67458
rect 137376 63572 137428 63578
rect 137376 63514 137428 63520
rect 137388 44878 137416 63514
rect 137376 44872 137428 44878
rect 137376 44814 137428 44820
rect 137284 37936 137336 37942
rect 137284 37878 137336 37884
rect 138216 28966 138244 73714
rect 138308 67289 138336 76502
rect 138480 76502 138532 76508
rect 138386 76463 138442 76472
rect 138294 67280 138350 67289
rect 138294 67215 138350 67224
rect 138308 64870 138336 67215
rect 138400 64874 138428 76463
rect 138480 76356 138532 76362
rect 138480 76298 138532 76304
rect 138492 65958 138520 76298
rect 138584 76090 138612 79494
rect 138676 77081 138704 79716
rect 139228 79744 139256 79784
rect 139366 79744 139394 80036
rect 139458 79830 139486 80036
rect 139550 79937 139578 80036
rect 139536 79928 139592 79937
rect 139536 79863 139592 79872
rect 139446 79824 139498 79830
rect 139642 79778 139670 80036
rect 139734 79937 139762 80036
rect 139826 79966 139854 80036
rect 139918 79966 139946 80036
rect 140010 79966 140038 80036
rect 139814 79960 139866 79966
rect 139720 79928 139776 79937
rect 139814 79902 139866 79908
rect 139906 79960 139958 79966
rect 139906 79902 139958 79908
rect 139998 79960 140050 79966
rect 139998 79902 140050 79908
rect 139720 79863 139776 79872
rect 139952 79824 140004 79830
rect 139446 79766 139498 79772
rect 138940 79698 138992 79704
rect 139136 79716 139256 79744
rect 139320 79716 139394 79744
rect 139596 79750 139670 79778
rect 139858 79792 139914 79801
rect 139952 79766 140004 79772
rect 140102 79778 140130 80036
rect 140194 79966 140222 80036
rect 140286 79966 140314 80036
rect 140182 79960 140234 79966
rect 140182 79902 140234 79908
rect 140274 79960 140326 79966
rect 140274 79902 140326 79908
rect 140378 79812 140406 80036
rect 140470 79966 140498 80036
rect 140458 79960 140510 79966
rect 140562 79937 140590 80036
rect 140654 79966 140682 80036
rect 140746 79966 140774 80036
rect 140642 79960 140694 79966
rect 140458 79902 140510 79908
rect 140548 79928 140604 79937
rect 140642 79902 140694 79908
rect 140734 79960 140786 79966
rect 140838 79937 140866 80036
rect 140930 79966 140958 80036
rect 141022 79966 141050 80036
rect 140918 79960 140970 79966
rect 140734 79902 140786 79908
rect 140824 79928 140880 79937
rect 140548 79863 140604 79872
rect 140918 79902 140970 79908
rect 141010 79960 141062 79966
rect 141114 79937 141142 80036
rect 141206 79966 141234 80036
rect 141194 79960 141246 79966
rect 141010 79902 141062 79908
rect 141100 79928 141156 79937
rect 140824 79863 140880 79872
rect 141298 79937 141326 80036
rect 141390 79966 141418 80036
rect 141378 79960 141430 79966
rect 141194 79902 141246 79908
rect 141284 79928 141340 79937
rect 141100 79863 141156 79872
rect 141378 79902 141430 79908
rect 141284 79863 141340 79872
rect 140240 79784 140406 79812
rect 140780 79824 140832 79830
rect 138756 79688 138808 79694
rect 138756 79630 138808 79636
rect 138768 78946 138796 79630
rect 138756 78940 138808 78946
rect 138756 78882 138808 78888
rect 138848 78260 138900 78266
rect 138848 78202 138900 78208
rect 138662 77072 138718 77081
rect 138662 77007 138718 77016
rect 138572 76084 138624 76090
rect 138572 76026 138624 76032
rect 138664 75336 138716 75342
rect 138664 75278 138716 75284
rect 138572 75268 138624 75274
rect 138572 75210 138624 75216
rect 138584 68814 138612 75210
rect 138676 68950 138704 75278
rect 138860 73778 138888 78202
rect 138952 77314 138980 79698
rect 139032 79688 139084 79694
rect 139032 79630 139084 79636
rect 138940 77308 138992 77314
rect 138940 77250 138992 77256
rect 138848 73772 138900 73778
rect 138848 73714 138900 73720
rect 139044 70394 139072 79630
rect 139136 78577 139164 79716
rect 139216 79620 139268 79626
rect 139216 79562 139268 79568
rect 139122 78568 139178 78577
rect 139122 78503 139178 78512
rect 139122 78296 139178 78305
rect 139122 78231 139178 78240
rect 139136 71330 139164 78231
rect 139124 71324 139176 71330
rect 139124 71266 139176 71272
rect 138952 70366 139072 70394
rect 138664 68944 138716 68950
rect 138664 68886 138716 68892
rect 138572 68808 138624 68814
rect 138624 68756 138888 68762
rect 138572 68750 138888 68756
rect 138584 68734 138888 68750
rect 138584 68685 138612 68734
rect 138756 67516 138808 67522
rect 138756 67458 138808 67464
rect 138768 67114 138796 67458
rect 138756 67108 138808 67114
rect 138756 67050 138808 67056
rect 138480 65952 138532 65958
rect 138480 65894 138532 65900
rect 138296 64864 138348 64870
rect 138400 64846 138704 64874
rect 138296 64806 138348 64812
rect 138676 64122 138704 64846
rect 138664 64116 138716 64122
rect 138664 64058 138716 64064
rect 138204 28960 138256 28966
rect 138204 28902 138256 28908
rect 138676 6186 138704 64058
rect 138768 40730 138796 67050
rect 138860 43450 138888 68734
rect 138952 67522 138980 70366
rect 139228 69562 139256 79562
rect 139320 75274 139348 79716
rect 139400 79620 139452 79626
rect 139400 79562 139452 79568
rect 139412 78402 139440 79562
rect 139596 78656 139624 79750
rect 139858 79727 139860 79736
rect 139912 79727 139914 79736
rect 139860 79698 139912 79704
rect 139676 79688 139728 79694
rect 139676 79630 139728 79636
rect 139504 78628 139624 78656
rect 139400 78396 139452 78402
rect 139400 78338 139452 78344
rect 139504 77110 139532 78628
rect 139582 78568 139638 78577
rect 139582 78503 139638 78512
rect 139492 77104 139544 77110
rect 139492 77046 139544 77052
rect 139308 75268 139360 75274
rect 139308 75210 139360 75216
rect 139596 75138 139624 78503
rect 139584 75132 139636 75138
rect 139584 75074 139636 75080
rect 139584 74996 139636 75002
rect 139584 74938 139636 74944
rect 139216 69556 139268 69562
rect 139216 69498 139268 69504
rect 138940 67516 138992 67522
rect 138940 67458 138992 67464
rect 139596 64190 139624 74938
rect 139688 64326 139716 79630
rect 139768 79620 139820 79626
rect 139768 79562 139820 79568
rect 139780 64394 139808 79562
rect 139964 78538 139992 79766
rect 140102 79750 140176 79778
rect 139952 78532 140004 78538
rect 139952 78474 140004 78480
rect 140148 78384 140176 79750
rect 139872 78356 140176 78384
rect 139872 68338 139900 78356
rect 140240 78282 140268 79784
rect 140780 79766 140832 79772
rect 140962 79792 141018 79801
rect 140688 79756 140740 79762
rect 140688 79698 140740 79704
rect 140412 79688 140464 79694
rect 139964 78254 140268 78282
rect 140332 79648 140412 79676
rect 139860 68332 139912 68338
rect 139860 68274 139912 68280
rect 139768 64388 139820 64394
rect 139768 64330 139820 64336
rect 139676 64320 139728 64326
rect 139676 64262 139728 64268
rect 139584 64184 139636 64190
rect 139584 64126 139636 64132
rect 138848 43444 138900 43450
rect 138848 43386 138900 43392
rect 138756 40724 138808 40730
rect 138756 40666 138808 40672
rect 139596 20670 139624 64126
rect 139688 63646 139716 64262
rect 139676 63640 139728 63646
rect 139676 63582 139728 63588
rect 139780 63578 139808 64330
rect 139768 63572 139820 63578
rect 139768 63514 139820 63520
rect 139964 55214 139992 78254
rect 140044 78192 140096 78198
rect 140044 78134 140096 78140
rect 140056 73817 140084 78134
rect 140332 77294 140360 79648
rect 140412 79630 140464 79636
rect 140502 79656 140558 79665
rect 140502 79591 140558 79600
rect 140596 79620 140648 79626
rect 140412 78056 140464 78062
rect 140412 77998 140464 78004
rect 140240 77266 140360 77294
rect 140042 73808 140098 73817
rect 140042 73743 140098 73752
rect 140136 63640 140188 63646
rect 140136 63582 140188 63588
rect 140044 63572 140096 63578
rect 140044 63514 140096 63520
rect 139952 55208 140004 55214
rect 139952 55150 140004 55156
rect 139584 20664 139636 20670
rect 139584 20606 139636 20612
rect 140056 14482 140084 63514
rect 140148 49026 140176 63582
rect 140240 57934 140268 77266
rect 140320 75132 140372 75138
rect 140320 75074 140372 75080
rect 140332 65890 140360 75074
rect 140424 74526 140452 77998
rect 140516 77217 140544 79591
rect 140596 79562 140648 79568
rect 140502 77208 140558 77217
rect 140502 77143 140558 77152
rect 140504 75472 140556 75478
rect 140504 75414 140556 75420
rect 140516 74866 140544 75414
rect 140504 74860 140556 74866
rect 140504 74802 140556 74808
rect 140412 74520 140464 74526
rect 140412 74462 140464 74468
rect 140320 65884 140372 65890
rect 140320 65826 140372 65832
rect 140608 65414 140636 79562
rect 140700 75002 140728 79698
rect 140792 76566 140820 79766
rect 141482 79778 141510 80036
rect 141574 79898 141602 80036
rect 141562 79892 141614 79898
rect 141562 79834 141614 79840
rect 140962 79727 141018 79736
rect 141436 79750 141510 79778
rect 140976 79642 141004 79727
rect 141332 79688 141384 79694
rect 141238 79656 141294 79665
rect 140976 79614 141096 79642
rect 140964 79552 141016 79558
rect 140964 79494 141016 79500
rect 140870 79384 140926 79393
rect 140870 79319 140926 79328
rect 140780 76560 140832 76566
rect 140780 76502 140832 76508
rect 140884 76226 140912 79319
rect 140872 76220 140924 76226
rect 140872 76162 140924 76168
rect 140688 74996 140740 75002
rect 140688 74938 140740 74944
rect 140976 70394 141004 79494
rect 141068 75410 141096 79614
rect 141332 79630 141384 79636
rect 141238 79591 141294 79600
rect 141252 78826 141280 79591
rect 141160 78798 141280 78826
rect 141160 76673 141188 78798
rect 141240 78736 141292 78742
rect 141240 78678 141292 78684
rect 141146 76664 141202 76673
rect 141146 76599 141202 76608
rect 141148 76220 141200 76226
rect 141148 76162 141200 76168
rect 141056 75404 141108 75410
rect 141056 75346 141108 75352
rect 141056 75132 141108 75138
rect 141056 75074 141108 75080
rect 140884 70366 141004 70394
rect 140884 65482 140912 70366
rect 141068 66162 141096 75074
rect 141056 66156 141108 66162
rect 141056 66098 141108 66104
rect 141160 65754 141188 76162
rect 141252 66065 141280 78678
rect 141344 77761 141372 79630
rect 141436 78441 141464 79750
rect 141666 79744 141694 80036
rect 141758 79966 141786 80036
rect 141850 79966 141878 80036
rect 141746 79960 141798 79966
rect 141746 79902 141798 79908
rect 141838 79960 141890 79966
rect 141942 79937 141970 80036
rect 142034 79966 142062 80036
rect 142022 79960 142074 79966
rect 141838 79902 141890 79908
rect 141928 79928 141984 79937
rect 142022 79902 142074 79908
rect 141928 79863 141984 79872
rect 141746 79824 141798 79830
rect 141798 79784 141878 79812
rect 141746 79766 141798 79772
rect 141620 79716 141694 79744
rect 141514 79520 141570 79529
rect 141514 79455 141570 79464
rect 141528 78810 141556 79455
rect 141620 79354 141648 79716
rect 141698 79656 141754 79665
rect 141850 79642 141878 79784
rect 141976 79756 142028 79762
rect 142126 79744 142154 80036
rect 142218 79898 142246 80036
rect 142310 79937 142338 80036
rect 142296 79928 142352 79937
rect 142206 79892 142258 79898
rect 142402 79898 142430 80036
rect 142494 79966 142522 80036
rect 142482 79960 142534 79966
rect 142482 79902 142534 79908
rect 142296 79863 142352 79872
rect 142390 79892 142442 79898
rect 142206 79834 142258 79840
rect 142390 79834 142442 79840
rect 142586 79778 142614 80036
rect 142540 79750 142614 79778
rect 142126 79716 142200 79744
rect 141976 79698 142028 79704
rect 141698 79591 141700 79600
rect 141752 79591 141754 79600
rect 141804 79614 141878 79642
rect 141700 79562 141752 79568
rect 141698 79520 141754 79529
rect 141698 79455 141754 79464
rect 141608 79348 141660 79354
rect 141608 79290 141660 79296
rect 141516 78804 141568 78810
rect 141516 78746 141568 78752
rect 141422 78432 141478 78441
rect 141422 78367 141478 78376
rect 141330 77752 141386 77761
rect 141330 77687 141386 77696
rect 141422 76664 141478 76673
rect 141422 76599 141478 76608
rect 141332 76560 141384 76566
rect 141332 76502 141384 76508
rect 141238 66056 141294 66065
rect 141238 65991 141294 66000
rect 141148 65748 141200 65754
rect 141148 65690 141200 65696
rect 140872 65476 140924 65482
rect 140872 65418 140924 65424
rect 140596 65408 140648 65414
rect 140596 65350 140648 65356
rect 141344 64802 141372 76502
rect 141436 68474 141464 76599
rect 141516 76560 141568 76566
rect 141516 76502 141568 76508
rect 141528 69902 141556 76502
rect 141712 71534 141740 79455
rect 141804 75070 141832 79614
rect 141884 79484 141936 79490
rect 141884 79426 141936 79432
rect 141896 78742 141924 79426
rect 141884 78736 141936 78742
rect 141884 78678 141936 78684
rect 141882 78568 141938 78577
rect 141882 78503 141938 78512
rect 141896 75138 141924 78503
rect 141884 75132 141936 75138
rect 141884 75074 141936 75080
rect 141792 75064 141844 75070
rect 141792 75006 141844 75012
rect 141988 73154 142016 79698
rect 142068 79620 142120 79626
rect 142068 79562 142120 79568
rect 142080 78334 142108 79562
rect 142172 78713 142200 79716
rect 142540 79694 142568 79750
rect 142528 79688 142580 79694
rect 142678 79676 142706 80036
rect 142770 79971 142798 80036
rect 142756 79962 142812 79971
rect 142756 79897 142812 79906
rect 142862 79812 142890 80036
rect 142954 79966 142982 80036
rect 143046 79971 143074 80036
rect 142942 79960 142994 79966
rect 142942 79902 142994 79908
rect 143032 79962 143088 79971
rect 143032 79897 143088 79906
rect 143138 79898 143166 80036
rect 143230 79966 143258 80036
rect 143218 79960 143270 79966
rect 143218 79902 143270 79908
rect 143126 79892 143178 79898
rect 143126 79834 143178 79840
rect 142862 79784 142936 79812
rect 142528 79630 142580 79636
rect 142632 79648 142706 79676
rect 142344 79552 142396 79558
rect 142344 79494 142396 79500
rect 142528 79552 142580 79558
rect 142528 79494 142580 79500
rect 142252 79484 142304 79490
rect 142252 79426 142304 79432
rect 142158 78704 142214 78713
rect 142158 78639 142214 78648
rect 142068 78328 142120 78334
rect 142068 78270 142120 78276
rect 142066 77752 142122 77761
rect 142066 77687 142122 77696
rect 142080 75682 142108 77687
rect 142068 75676 142120 75682
rect 142068 75618 142120 75624
rect 142068 75404 142120 75410
rect 142068 75346 142120 75352
rect 141896 73126 142016 73154
rect 141700 71528 141752 71534
rect 141700 71470 141752 71476
rect 141896 70394 141924 73126
rect 141620 70366 141924 70394
rect 141974 70408 142030 70417
rect 141516 69896 141568 69902
rect 141516 69838 141568 69844
rect 141424 68468 141476 68474
rect 141424 68410 141476 68416
rect 141516 65476 141568 65482
rect 141516 65418 141568 65424
rect 141332 64796 141384 64802
rect 141332 64738 141384 64744
rect 141424 64456 141476 64462
rect 141424 64398 141476 64404
rect 140228 57928 140280 57934
rect 140228 57870 140280 57876
rect 140136 49020 140188 49026
rect 140136 48962 140188 48968
rect 141436 28286 141464 64398
rect 141528 55894 141556 65418
rect 141620 64705 141648 70366
rect 141974 70343 142030 70352
rect 141988 69737 142016 70343
rect 141974 69728 142030 69737
rect 141974 69663 142030 69672
rect 141606 64696 141662 64705
rect 141606 64631 141662 64640
rect 142080 64462 142108 75346
rect 142264 74186 142292 79426
rect 142356 75478 142384 79494
rect 142344 75472 142396 75478
rect 142344 75414 142396 75420
rect 142252 74180 142304 74186
rect 142252 74122 142304 74128
rect 142068 64456 142120 64462
rect 142068 64398 142120 64404
rect 142540 63374 142568 79494
rect 142632 73982 142660 79648
rect 142804 79620 142856 79626
rect 142908 79608 142936 79784
rect 143080 79756 143132 79762
rect 143080 79698 143132 79704
rect 143172 79756 143224 79762
rect 143322 79744 143350 80036
rect 143414 79830 143442 80036
rect 143506 79966 143534 80036
rect 143598 79966 143626 80036
rect 143494 79960 143546 79966
rect 143494 79902 143546 79908
rect 143586 79960 143638 79966
rect 143586 79902 143638 79908
rect 143402 79824 143454 79830
rect 143402 79766 143454 79772
rect 143690 79744 143718 80036
rect 143782 79966 143810 80036
rect 143770 79960 143822 79966
rect 143770 79902 143822 79908
rect 143874 79812 143902 80036
rect 143966 79966 143994 80036
rect 143954 79960 144006 79966
rect 143954 79902 144006 79908
rect 144058 79898 144086 80036
rect 144046 79892 144098 79898
rect 144046 79834 144098 79840
rect 143172 79698 143224 79704
rect 143276 79716 143350 79744
rect 143644 79716 143718 79744
rect 143828 79784 143902 79812
rect 142908 79580 143028 79608
rect 142804 79562 142856 79568
rect 142712 78736 142764 78742
rect 142712 78678 142764 78684
rect 142620 73976 142672 73982
rect 142620 73918 142672 73924
rect 142724 65550 142752 78678
rect 142816 78577 142844 79562
rect 142896 79484 142948 79490
rect 142896 79426 142948 79432
rect 142908 78713 142936 79426
rect 143000 78742 143028 79580
rect 142988 78736 143040 78742
rect 142894 78704 142950 78713
rect 142988 78678 143040 78684
rect 142894 78639 142950 78648
rect 142802 78568 142858 78577
rect 142802 78503 142858 78512
rect 142988 78532 143040 78538
rect 142988 78474 143040 78480
rect 142896 77648 142948 77654
rect 142896 77590 142948 77596
rect 142804 74656 142856 74662
rect 142804 74598 142856 74604
rect 142712 65544 142764 65550
rect 142712 65486 142764 65492
rect 142528 63368 142580 63374
rect 142528 63310 142580 63316
rect 141516 55888 141568 55894
rect 141516 55830 141568 55836
rect 141424 28280 141476 28286
rect 141424 28222 141476 28228
rect 140044 14476 140096 14482
rect 140044 14418 140096 14424
rect 138664 6180 138716 6186
rect 138664 6122 138716 6128
rect 136548 3528 136600 3534
rect 136548 3470 136600 3476
rect 135904 3324 135956 3330
rect 135904 3266 135956 3272
rect 136560 480 136588 3470
rect 142816 3466 142844 74598
rect 142908 71602 142936 77590
rect 143000 71738 143028 78474
rect 143092 76566 143120 79698
rect 143080 76560 143132 76566
rect 143080 76502 143132 76508
rect 143080 75472 143132 75478
rect 143184 75449 143212 79698
rect 143276 78130 143304 79716
rect 143540 79688 143592 79694
rect 143540 79630 143592 79636
rect 143356 79620 143408 79626
rect 143356 79562 143408 79568
rect 143448 79620 143500 79626
rect 143448 79562 143500 79568
rect 143368 78674 143396 79562
rect 143356 78668 143408 78674
rect 143356 78610 143408 78616
rect 143264 78124 143316 78130
rect 143264 78066 143316 78072
rect 143460 77294 143488 79562
rect 143552 78713 143580 79630
rect 143538 78704 143594 78713
rect 143538 78639 143594 78648
rect 143460 77266 143580 77294
rect 143552 75954 143580 77266
rect 143540 75948 143592 75954
rect 143540 75890 143592 75896
rect 143080 75414 143132 75420
rect 143170 75440 143226 75449
rect 142988 71732 143040 71738
rect 142988 71674 143040 71680
rect 142896 71596 142948 71602
rect 142896 71538 142948 71544
rect 143092 70394 143120 75414
rect 143170 75375 143226 75384
rect 143552 72690 143580 75890
rect 143540 72684 143592 72690
rect 143540 72626 143592 72632
rect 142908 70366 143120 70394
rect 142908 64190 142936 70366
rect 143644 67454 143672 79716
rect 143828 79665 143856 79784
rect 144150 79778 144178 80036
rect 144242 79937 144270 80036
rect 144334 79966 144362 80036
rect 144426 79966 144454 80036
rect 144518 79971 144546 80036
rect 144322 79960 144374 79966
rect 144228 79928 144284 79937
rect 144322 79902 144374 79908
rect 144414 79960 144466 79966
rect 144414 79902 144466 79908
rect 144504 79962 144560 79971
rect 144610 79966 144638 80036
rect 144702 79966 144730 80036
rect 144794 79966 144822 80036
rect 144886 79971 144914 80036
rect 144504 79897 144560 79906
rect 144598 79960 144650 79966
rect 144598 79902 144650 79908
rect 144690 79960 144742 79966
rect 144690 79902 144742 79908
rect 144782 79960 144834 79966
rect 144782 79902 144834 79908
rect 144872 79962 144928 79971
rect 144872 79897 144928 79906
rect 144978 79898 145006 80036
rect 144228 79863 144284 79872
rect 144966 79892 145018 79898
rect 144966 79834 145018 79840
rect 144690 79824 144742 79830
rect 144742 79801 144776 79812
rect 144742 79792 144790 79801
rect 144150 79750 144500 79778
rect 144690 79766 144734 79772
rect 144000 79688 144052 79694
rect 143814 79656 143870 79665
rect 144276 79688 144328 79694
rect 144000 79630 144052 79636
rect 144182 79656 144238 79665
rect 143814 79591 143870 79600
rect 143908 79620 143960 79626
rect 143908 79562 143960 79568
rect 143816 79484 143868 79490
rect 143816 79426 143868 79432
rect 143828 74390 143856 79426
rect 143920 75342 143948 79562
rect 143908 75336 143960 75342
rect 143908 75278 143960 75284
rect 143816 74384 143868 74390
rect 143816 74326 143868 74332
rect 144012 72729 144040 79630
rect 144092 79620 144144 79626
rect 144276 79630 144328 79636
rect 144182 79591 144238 79600
rect 144092 79562 144144 79568
rect 144104 76634 144132 79562
rect 144092 76628 144144 76634
rect 144092 76570 144144 76576
rect 144196 74361 144224 79591
rect 144182 74352 144238 74361
rect 144182 74287 144238 74296
rect 143998 72720 144054 72729
rect 143998 72655 144054 72664
rect 144288 70394 144316 79630
rect 144472 71233 144500 79750
rect 145070 79744 145098 80036
rect 145162 79898 145190 80036
rect 145254 79966 145282 80036
rect 145242 79960 145294 79966
rect 145346 79937 145374 80036
rect 145438 79966 145466 80036
rect 145530 79966 145558 80036
rect 145622 79966 145650 80036
rect 145426 79960 145478 79966
rect 145242 79902 145294 79908
rect 145332 79928 145388 79937
rect 145150 79892 145202 79898
rect 145426 79902 145478 79908
rect 145518 79960 145570 79966
rect 145518 79902 145570 79908
rect 145610 79960 145662 79966
rect 145610 79902 145662 79908
rect 145332 79863 145388 79872
rect 145150 79834 145202 79840
rect 145380 79824 145432 79830
rect 145380 79766 145432 79772
rect 144734 79727 144790 79736
rect 145024 79716 145098 79744
rect 144552 79688 144604 79694
rect 144552 79630 144604 79636
rect 144736 79688 144788 79694
rect 144736 79630 144788 79636
rect 144564 77722 144592 79630
rect 144552 77716 144604 77722
rect 144552 77658 144604 77664
rect 144458 71224 144514 71233
rect 144458 71159 144514 71168
rect 144748 71074 144776 79630
rect 144826 76664 144882 76673
rect 144826 76599 144882 76608
rect 143920 70366 144316 70394
rect 144380 71046 144776 71074
rect 143920 69873 143948 70366
rect 143906 69864 143962 69873
rect 143906 69799 143962 69808
rect 144380 67590 144408 71046
rect 144840 70394 144868 76599
rect 145024 71641 145052 79716
rect 145196 79688 145248 79694
rect 145196 79630 145248 79636
rect 145104 79620 145156 79626
rect 145104 79562 145156 79568
rect 145116 74050 145144 79562
rect 145208 75834 145236 79630
rect 145288 79620 145340 79626
rect 145288 79562 145340 79568
rect 145300 78674 145328 79562
rect 145288 78668 145340 78674
rect 145288 78610 145340 78616
rect 145286 75848 145342 75857
rect 145208 75806 145286 75834
rect 145286 75783 145342 75792
rect 145300 75177 145328 75783
rect 145286 75168 145342 75177
rect 145286 75103 145342 75112
rect 145392 74934 145420 79766
rect 145472 79756 145524 79762
rect 145472 79698 145524 79704
rect 145564 79756 145616 79762
rect 145714 79744 145742 80036
rect 145806 79898 145834 80036
rect 145898 79966 145926 80036
rect 145990 79971 146018 80036
rect 145886 79960 145938 79966
rect 145886 79902 145938 79908
rect 145976 79962 146032 79971
rect 146082 79966 146110 80036
rect 146174 79966 146202 80036
rect 146266 79971 146294 80036
rect 145794 79892 145846 79898
rect 145976 79897 146032 79906
rect 146070 79960 146122 79966
rect 146070 79902 146122 79908
rect 146162 79960 146214 79966
rect 146162 79902 146214 79908
rect 146252 79962 146308 79971
rect 146358 79966 146386 80036
rect 146252 79897 146308 79906
rect 146346 79960 146398 79966
rect 146346 79902 146398 79908
rect 146450 79898 146478 80036
rect 146542 79971 146570 80036
rect 146528 79962 146584 79971
rect 145794 79834 145846 79840
rect 146438 79892 146490 79898
rect 146528 79897 146584 79906
rect 146634 79898 146662 80036
rect 146726 79903 146754 80036
rect 146818 79966 146846 80036
rect 146806 79960 146858 79966
rect 146438 79834 146490 79840
rect 146622 79892 146674 79898
rect 146622 79834 146674 79840
rect 146712 79894 146768 79903
rect 146806 79902 146858 79908
rect 146910 79898 146938 80036
rect 147002 79898 147030 80036
rect 147094 79937 147122 80036
rect 147080 79928 147136 79937
rect 145932 79824 145984 79830
rect 145932 79766 145984 79772
rect 146070 79824 146122 79830
rect 146712 79829 146768 79838
rect 146898 79892 146950 79898
rect 146898 79834 146950 79840
rect 146990 79892 147042 79898
rect 147186 79898 147214 80036
rect 147278 79898 147306 80036
rect 147370 79966 147398 80036
rect 147462 79966 147490 80036
rect 147554 79966 147582 80036
rect 147358 79960 147410 79966
rect 147358 79902 147410 79908
rect 147450 79960 147502 79966
rect 147450 79902 147502 79908
rect 147542 79960 147594 79966
rect 147542 79902 147594 79908
rect 147646 79898 147674 80036
rect 147738 79937 147766 80036
rect 147724 79928 147780 79937
rect 147080 79863 147136 79872
rect 147174 79892 147226 79898
rect 146990 79834 147042 79840
rect 147174 79834 147226 79840
rect 147266 79892 147318 79898
rect 147266 79834 147318 79840
rect 147634 79892 147686 79898
rect 147724 79863 147780 79872
rect 147634 79834 147686 79840
rect 147404 79824 147456 79830
rect 146122 79772 146202 79778
rect 146070 79766 146202 79772
rect 147404 79766 147456 79772
rect 147496 79824 147548 79830
rect 147830 79812 147858 80036
rect 147784 79784 147858 79812
rect 147784 79778 147812 79784
rect 147496 79766 147548 79772
rect 145564 79698 145616 79704
rect 145668 79716 145742 79744
rect 145840 79756 145892 79762
rect 145484 78792 145512 79698
rect 145576 79218 145604 79698
rect 145564 79212 145616 79218
rect 145564 79154 145616 79160
rect 145484 78764 145604 78792
rect 145472 78668 145524 78674
rect 145472 78610 145524 78616
rect 145380 74928 145432 74934
rect 145380 74870 145432 74876
rect 145104 74044 145156 74050
rect 145104 73986 145156 73992
rect 145116 73846 145144 73986
rect 145104 73840 145156 73846
rect 145104 73782 145156 73788
rect 145010 71632 145066 71641
rect 145010 71567 145066 71576
rect 144472 70366 144868 70394
rect 144368 67584 144420 67590
rect 144368 67526 144420 67532
rect 143632 67448 143684 67454
rect 143632 67390 143684 67396
rect 144276 67448 144328 67454
rect 144276 67390 144328 67396
rect 142896 64184 142948 64190
rect 142896 64126 142948 64132
rect 143448 63368 143500 63374
rect 143448 63310 143500 63316
rect 143460 58682 143488 63310
rect 143448 58676 143500 58682
rect 143448 58618 143500 58624
rect 144184 51060 144236 51066
rect 144184 51002 144236 51008
rect 142804 3460 142856 3466
rect 142804 3402 142856 3408
rect 144196 3398 144224 51002
rect 144288 36582 144316 67390
rect 144380 50454 144408 67526
rect 144368 50448 144420 50454
rect 144368 50390 144420 50396
rect 144472 48278 144500 70366
rect 145484 67590 145512 78610
rect 145576 75002 145604 78764
rect 145668 75886 145696 79716
rect 145840 79698 145892 79704
rect 145852 78169 145880 79698
rect 145944 79014 145972 79766
rect 146082 79750 146202 79766
rect 146024 79620 146076 79626
rect 146174 79608 146202 79750
rect 147220 79756 147272 79762
rect 147220 79698 147272 79704
rect 147312 79756 147364 79762
rect 147312 79698 147364 79704
rect 146944 79688 146996 79694
rect 146574 79656 146630 79665
rect 146024 79562 146076 79568
rect 146128 79580 146202 79608
rect 146484 79620 146536 79626
rect 145932 79008 145984 79014
rect 145932 78950 145984 78956
rect 145838 78160 145894 78169
rect 145838 78095 145894 78104
rect 145932 78124 145984 78130
rect 145932 78066 145984 78072
rect 145656 75880 145708 75886
rect 145656 75822 145708 75828
rect 145564 74996 145616 75002
rect 145564 74938 145616 74944
rect 145668 74050 145696 75822
rect 145944 74202 145972 78066
rect 146036 77994 146064 79562
rect 146128 78266 146156 79580
rect 146944 79630 146996 79636
rect 146574 79591 146630 79600
rect 146852 79620 146904 79626
rect 146484 79562 146536 79568
rect 146392 79552 146444 79558
rect 146392 79494 146444 79500
rect 146404 79150 146432 79494
rect 146392 79144 146444 79150
rect 146392 79086 146444 79092
rect 146300 78328 146352 78334
rect 146300 78270 146352 78276
rect 146116 78260 146168 78266
rect 146116 78202 146168 78208
rect 146024 77988 146076 77994
rect 146024 77930 146076 77936
rect 146116 74996 146168 75002
rect 146116 74938 146168 74944
rect 145760 74174 145972 74202
rect 145564 74044 145616 74050
rect 145564 73986 145616 73992
rect 145656 74044 145708 74050
rect 145656 73986 145708 73992
rect 145472 67584 145524 67590
rect 145472 67526 145524 67532
rect 144460 48272 144512 48278
rect 144460 48214 144512 48220
rect 144276 36576 144328 36582
rect 144276 36518 144328 36524
rect 145576 4826 145604 73986
rect 145656 67584 145708 67590
rect 145760 67561 145788 74174
rect 146128 74118 146156 74938
rect 146116 74112 146168 74118
rect 146116 74054 146168 74060
rect 145932 74044 145984 74050
rect 145932 73986 145984 73992
rect 145656 67526 145708 67532
rect 145746 67552 145802 67561
rect 145668 67386 145696 67526
rect 145746 67487 145802 67496
rect 145656 67380 145708 67386
rect 145656 67322 145708 67328
rect 145668 54602 145696 67322
rect 145944 66910 145972 73986
rect 146128 70394 146156 74054
rect 146312 71777 146340 78270
rect 146496 76673 146524 79562
rect 146482 76664 146538 76673
rect 146482 76599 146538 76608
rect 146588 75478 146616 79591
rect 146852 79562 146904 79568
rect 146760 79552 146812 79558
rect 146760 79494 146812 79500
rect 146668 76832 146720 76838
rect 146668 76774 146720 76780
rect 146576 75472 146628 75478
rect 146576 75414 146628 75420
rect 146298 71768 146354 71777
rect 146298 71703 146354 71712
rect 146680 70394 146708 76774
rect 146772 76634 146800 79494
rect 146760 76628 146812 76634
rect 146760 76570 146812 76576
rect 146760 76356 146812 76362
rect 146760 76298 146812 76304
rect 146036 70366 146156 70394
rect 146496 70366 146708 70394
rect 145932 66904 145984 66910
rect 145932 66846 145984 66852
rect 146036 65550 146064 70366
rect 146496 68746 146524 70366
rect 146484 68740 146536 68746
rect 146484 68682 146536 68688
rect 146772 67561 146800 76298
rect 146864 76022 146892 79562
rect 146852 76016 146904 76022
rect 146852 75958 146904 75964
rect 146852 75268 146904 75274
rect 146852 75210 146904 75216
rect 146864 68610 146892 75210
rect 146956 73953 146984 79630
rect 147036 79552 147088 79558
rect 147232 79506 147260 79698
rect 147036 79494 147088 79500
rect 147048 76838 147076 79494
rect 147140 79478 147260 79506
rect 147036 76832 147088 76838
rect 147036 76774 147088 76780
rect 147036 76628 147088 76634
rect 147036 76570 147088 76576
rect 146942 73944 146998 73953
rect 146942 73879 146998 73888
rect 147048 73154 147076 76570
rect 146956 73126 147076 73154
rect 146956 72554 146984 73126
rect 146944 72548 146996 72554
rect 146944 72490 146996 72496
rect 146852 68604 146904 68610
rect 146852 68546 146904 68552
rect 146758 67552 146814 67561
rect 146758 67487 146814 67496
rect 146024 65544 146076 65550
rect 146024 65486 146076 65492
rect 146300 62960 146352 62966
rect 146300 62902 146352 62908
rect 145656 54596 145708 54602
rect 145656 54538 145708 54544
rect 145564 4820 145616 4826
rect 145564 4762 145616 4768
rect 146312 3466 146340 62902
rect 146956 18698 146984 72490
rect 147140 70922 147168 79478
rect 147324 76362 147352 79698
rect 147312 76356 147364 76362
rect 147312 76298 147364 76304
rect 147220 76016 147272 76022
rect 147220 75958 147272 75964
rect 147232 74866 147260 75958
rect 147416 75585 147444 79766
rect 147402 75576 147458 75585
rect 147402 75511 147458 75520
rect 147404 75472 147456 75478
rect 147404 75414 147456 75420
rect 147220 74860 147272 74866
rect 147220 74802 147272 74808
rect 147128 70916 147180 70922
rect 147128 70858 147180 70864
rect 147140 70394 147168 70858
rect 147048 70366 147168 70394
rect 147048 43518 147076 70366
rect 147126 67552 147182 67561
rect 147126 67487 147182 67496
rect 147140 67017 147168 67487
rect 147126 67008 147182 67017
rect 147126 66943 147182 66952
rect 147140 53106 147168 66943
rect 147232 65618 147260 74802
rect 147416 69834 147444 75414
rect 147508 75274 147536 79766
rect 147588 79756 147640 79762
rect 147738 79750 147812 79778
rect 147922 79778 147950 80036
rect 148014 79903 148042 80036
rect 148106 79966 148134 80036
rect 148198 79971 148226 80036
rect 148094 79960 148146 79966
rect 148000 79894 148056 79903
rect 148094 79902 148146 79908
rect 148184 79962 148240 79971
rect 148184 79897 148240 79906
rect 148000 79829 148056 79838
rect 147922 79750 147996 79778
rect 147738 79744 147766 79750
rect 147588 79698 147640 79704
rect 147692 79716 147766 79744
rect 147600 75750 147628 79698
rect 147588 75744 147640 75750
rect 147588 75686 147640 75692
rect 147496 75268 147548 75274
rect 147496 75210 147548 75216
rect 147692 74497 147720 79716
rect 147968 77110 147996 79750
rect 148290 79744 148318 80036
rect 148382 79971 148410 80036
rect 148368 79962 148424 79971
rect 148368 79897 148424 79906
rect 148474 79744 148502 80036
rect 148566 79898 148594 80036
rect 148554 79892 148606 79898
rect 148554 79834 148606 79840
rect 148658 79778 148686 80036
rect 148750 79937 148778 80036
rect 148842 79966 148870 80036
rect 148934 79966 148962 80036
rect 149026 79966 149054 80036
rect 148830 79960 148882 79966
rect 148736 79928 148792 79937
rect 148830 79902 148882 79908
rect 148922 79960 148974 79966
rect 148922 79902 148974 79908
rect 149014 79960 149066 79966
rect 149014 79902 149066 79908
rect 148736 79863 148792 79872
rect 148612 79750 148686 79778
rect 148968 79824 149020 79830
rect 148968 79766 149020 79772
rect 148876 79756 148928 79762
rect 148290 79716 148364 79744
rect 148474 79716 148548 79744
rect 148230 79656 148286 79665
rect 148230 79591 148286 79600
rect 148140 79552 148192 79558
rect 148140 79494 148192 79500
rect 147956 77104 148008 77110
rect 147956 77046 148008 77052
rect 148152 76566 148180 79494
rect 148244 76786 148272 79591
rect 148336 79121 148364 79716
rect 148414 79656 148470 79665
rect 148414 79591 148470 79600
rect 148322 79112 148378 79121
rect 148322 79047 148378 79056
rect 148244 76758 148364 76786
rect 148232 76696 148284 76702
rect 148232 76638 148284 76644
rect 148140 76560 148192 76566
rect 148140 76502 148192 76508
rect 148140 75472 148192 75478
rect 148140 75414 148192 75420
rect 147678 74488 147734 74497
rect 147678 74423 147734 74432
rect 147680 71460 147732 71466
rect 147680 71402 147732 71408
rect 147404 69828 147456 69834
rect 147404 69770 147456 69776
rect 147220 65612 147272 65618
rect 147220 65554 147272 65560
rect 147128 53100 147180 53106
rect 147128 53042 147180 53048
rect 147036 43512 147088 43518
rect 147036 43454 147088 43460
rect 146944 18692 146996 18698
rect 146944 18634 146996 18640
rect 147692 6254 147720 71402
rect 148152 66978 148180 75414
rect 148140 66972 148192 66978
rect 148140 66914 148192 66920
rect 148152 55214 148180 66914
rect 148244 66842 148272 76638
rect 148336 71466 148364 76758
rect 148428 75478 148456 79591
rect 148520 75546 148548 79716
rect 148612 76702 148640 79750
rect 148876 79698 148928 79704
rect 148692 79688 148744 79694
rect 148692 79630 148744 79636
rect 148600 76696 148652 76702
rect 148600 76638 148652 76644
rect 148600 76560 148652 76566
rect 148600 76502 148652 76508
rect 148508 75540 148560 75546
rect 148508 75482 148560 75488
rect 148416 75472 148468 75478
rect 148416 75414 148468 75420
rect 148416 71732 148468 71738
rect 148416 71674 148468 71680
rect 148324 71460 148376 71466
rect 148324 71402 148376 71408
rect 148428 71398 148456 71674
rect 148416 71392 148468 71398
rect 148416 71334 148468 71340
rect 148232 66836 148284 66842
rect 148232 66778 148284 66784
rect 148244 64326 148272 66778
rect 148232 64320 148284 64326
rect 148232 64262 148284 64268
rect 148152 55186 148364 55214
rect 148336 26926 148364 55186
rect 148428 42090 148456 71334
rect 148520 62898 148548 75482
rect 148612 68542 148640 76502
rect 148704 71738 148732 79630
rect 148784 79620 148836 79626
rect 148784 79562 148836 79568
rect 148796 72826 148824 79562
rect 148888 77858 148916 79698
rect 148876 77852 148928 77858
rect 148876 77794 148928 77800
rect 148980 76770 149008 79766
rect 149118 79744 149146 80036
rect 149210 79830 149238 80036
rect 149302 79835 149330 80036
rect 149198 79824 149250 79830
rect 149198 79766 149250 79772
rect 149288 79826 149344 79835
rect 149288 79761 149344 79770
rect 149072 79716 149146 79744
rect 149394 79744 149422 80036
rect 149486 79966 149514 80036
rect 149578 79966 149606 80036
rect 149670 79966 149698 80036
rect 149474 79960 149526 79966
rect 149474 79902 149526 79908
rect 149566 79960 149618 79966
rect 149566 79902 149618 79908
rect 149658 79960 149710 79966
rect 149658 79902 149710 79908
rect 149762 79898 149790 80036
rect 149854 79898 149882 80036
rect 149946 79898 149974 80036
rect 149750 79892 149802 79898
rect 149750 79834 149802 79840
rect 149842 79892 149894 79898
rect 149842 79834 149894 79840
rect 149934 79892 149986 79898
rect 149934 79834 149986 79840
rect 149612 79756 149664 79762
rect 149394 79716 149468 79744
rect 148968 76764 149020 76770
rect 148968 76706 149020 76712
rect 148784 72820 148836 72826
rect 148784 72762 148836 72768
rect 149072 72758 149100 79716
rect 149440 79665 149468 79716
rect 149612 79698 149664 79704
rect 149704 79756 149756 79762
rect 149704 79698 149756 79704
rect 149796 79756 149848 79762
rect 149796 79698 149848 79704
rect 149520 79688 149572 79694
rect 149426 79656 149482 79665
rect 149152 79620 149204 79626
rect 149520 79630 149572 79636
rect 149426 79591 149482 79600
rect 149152 79562 149204 79568
rect 149164 75614 149192 79562
rect 149244 79552 149296 79558
rect 149244 79494 149296 79500
rect 149334 79520 149390 79529
rect 149256 79286 149284 79494
rect 149334 79455 149390 79464
rect 149244 79280 149296 79286
rect 149244 79222 149296 79228
rect 149348 77294 149376 79455
rect 149428 79416 149480 79422
rect 149428 79358 149480 79364
rect 149440 79082 149468 79358
rect 149428 79076 149480 79082
rect 149428 79018 149480 79024
rect 149256 77266 149376 77294
rect 149152 75608 149204 75614
rect 149152 75550 149204 75556
rect 149256 73030 149284 77266
rect 149336 74044 149388 74050
rect 149336 73986 149388 73992
rect 149348 73234 149376 73986
rect 149336 73228 149388 73234
rect 149336 73170 149388 73176
rect 149244 73024 149296 73030
rect 149244 72966 149296 72972
rect 149060 72752 149112 72758
rect 149060 72694 149112 72700
rect 148692 71732 148744 71738
rect 148692 71674 148744 71680
rect 148600 68536 148652 68542
rect 148600 68478 148652 68484
rect 149256 68338 149284 72966
rect 149348 70174 149376 73170
rect 149532 70394 149560 79630
rect 149624 78033 149652 79698
rect 149610 78024 149666 78033
rect 149610 77959 149666 77968
rect 149716 73778 149744 79698
rect 149808 75041 149836 79698
rect 149888 79688 149940 79694
rect 150038 79676 150066 80036
rect 150130 79898 150158 80036
rect 150118 79892 150170 79898
rect 150118 79834 150170 79840
rect 150222 79744 150250 80036
rect 150314 79898 150342 80036
rect 150302 79892 150354 79898
rect 150302 79834 150354 79840
rect 150406 79778 150434 80036
rect 149888 79630 149940 79636
rect 149992 79648 150066 79676
rect 150176 79716 150250 79744
rect 150360 79750 150434 79778
rect 149794 75032 149850 75041
rect 149794 74967 149850 74976
rect 149900 74050 149928 79630
rect 149992 77761 150020 79648
rect 149978 77752 150034 77761
rect 149978 77687 150034 77696
rect 150176 77625 150204 79716
rect 150256 79484 150308 79490
rect 150256 79426 150308 79432
rect 150162 77616 150218 77625
rect 150162 77551 150218 77560
rect 149980 77104 150032 77110
rect 149980 77046 150032 77052
rect 149888 74044 149940 74050
rect 149888 73986 149940 73992
rect 149704 73772 149756 73778
rect 149704 73714 149756 73720
rect 149796 73092 149848 73098
rect 149796 73034 149848 73040
rect 149808 72418 149836 73034
rect 149796 72412 149848 72418
rect 149796 72354 149848 72360
rect 149532 70366 149652 70394
rect 149336 70168 149388 70174
rect 149336 70110 149388 70116
rect 149244 68332 149296 68338
rect 149244 68274 149296 68280
rect 149624 66774 149652 70366
rect 149612 66768 149664 66774
rect 149612 66710 149664 66716
rect 149624 64874 149652 66710
rect 149624 64846 149744 64874
rect 148508 62892 148560 62898
rect 148508 62834 148560 62840
rect 148416 42084 148468 42090
rect 148416 42026 148468 42032
rect 148324 26920 148376 26926
rect 148324 26862 148376 26868
rect 149716 11762 149744 64846
rect 149808 61470 149836 72354
rect 149992 70394 150020 77046
rect 150268 70394 150296 79426
rect 150360 73098 150388 79750
rect 150498 79676 150526 80036
rect 150590 79971 150618 80036
rect 150576 79962 150632 79971
rect 150576 79897 150632 79906
rect 150682 79830 150710 80036
rect 150774 79966 150802 80036
rect 150762 79960 150814 79966
rect 150762 79902 150814 79908
rect 150670 79824 150722 79830
rect 150866 79812 150894 80036
rect 150958 79971 150986 80036
rect 150944 79962 151000 79971
rect 151050 79966 151078 80036
rect 150944 79897 151000 79906
rect 151038 79960 151090 79966
rect 151038 79902 151090 79908
rect 150820 79784 150894 79812
rect 150820 79778 150848 79784
rect 150670 79766 150722 79772
rect 150452 79648 150526 79676
rect 150774 79750 150848 79778
rect 150774 79676 150802 79750
rect 151142 79744 151170 80036
rect 151096 79716 151170 79744
rect 151234 79744 151262 80036
rect 151326 79898 151354 80036
rect 151418 79966 151446 80036
rect 151510 79971 151538 80036
rect 151406 79960 151458 79966
rect 151406 79902 151458 79908
rect 151496 79962 151552 79971
rect 151602 79966 151630 80036
rect 151694 79966 151722 80036
rect 151314 79892 151366 79898
rect 151496 79897 151552 79906
rect 151590 79960 151642 79966
rect 151590 79902 151642 79908
rect 151682 79960 151734 79966
rect 151682 79902 151734 79908
rect 151314 79834 151366 79840
rect 151498 79824 151550 79830
rect 151786 79812 151814 80036
rect 151878 79966 151906 80036
rect 151970 79966 151998 80036
rect 151866 79960 151918 79966
rect 151866 79902 151918 79908
rect 151958 79960 152010 79966
rect 151958 79902 152010 79908
rect 152062 79898 152090 80036
rect 152050 79892 152102 79898
rect 152050 79834 152102 79840
rect 152154 79830 152182 80036
rect 151550 79784 151676 79812
rect 151498 79766 151550 79772
rect 151234 79716 151308 79744
rect 150774 79648 150848 79676
rect 150452 75274 150480 79648
rect 150716 79552 150768 79558
rect 150622 79520 150678 79529
rect 150532 79484 150584 79490
rect 150716 79494 150768 79500
rect 150622 79455 150678 79464
rect 150532 79426 150584 79432
rect 150440 75268 150492 75274
rect 150440 75210 150492 75216
rect 150348 73092 150400 73098
rect 150348 73034 150400 73040
rect 150544 70786 150572 79426
rect 150532 70780 150584 70786
rect 150532 70722 150584 70728
rect 150544 70394 150572 70722
rect 149900 70366 150020 70394
rect 150084 70366 150296 70394
rect 150452 70366 150572 70394
rect 150636 70394 150664 79455
rect 150728 78198 150756 79494
rect 150716 78192 150768 78198
rect 150716 78134 150768 78140
rect 150716 76696 150768 76702
rect 150716 76638 150768 76644
rect 150728 74254 150756 76638
rect 150820 76498 150848 79648
rect 150898 79656 150954 79665
rect 150898 79591 150954 79600
rect 150912 76702 150940 79591
rect 150992 79552 151044 79558
rect 150992 79494 151044 79500
rect 150900 76696 150952 76702
rect 150900 76638 150952 76644
rect 150900 76560 150952 76566
rect 150900 76502 150952 76508
rect 150808 76492 150860 76498
rect 150808 76434 150860 76440
rect 150716 74248 150768 74254
rect 150716 74190 150768 74196
rect 150636 70366 150848 70394
rect 149900 66201 149928 70366
rect 150084 68406 150112 70366
rect 150452 68406 150480 70366
rect 150072 68400 150124 68406
rect 150072 68342 150124 68348
rect 150440 68400 150492 68406
rect 150440 68342 150492 68348
rect 149886 66192 149942 66201
rect 149886 66127 149942 66136
rect 150820 63442 150848 70366
rect 150808 63436 150860 63442
rect 150808 63378 150860 63384
rect 149796 61464 149848 61470
rect 149796 61406 149848 61412
rect 150440 56636 150492 56642
rect 150440 56578 150492 56584
rect 150452 16574 150480 56578
rect 150912 48278 150940 76502
rect 151004 70310 151032 79494
rect 151096 76401 151124 79716
rect 151082 76392 151138 76401
rect 151082 76327 151138 76336
rect 151176 75268 151228 75274
rect 151176 75210 151228 75216
rect 150992 70304 151044 70310
rect 150992 70246 151044 70252
rect 151188 70242 151216 75210
rect 151280 73710 151308 79716
rect 151544 79688 151596 79694
rect 151450 79656 151506 79665
rect 151360 79620 151412 79626
rect 151544 79630 151596 79636
rect 151450 79591 151506 79600
rect 151360 79562 151412 79568
rect 151268 73704 151320 73710
rect 151268 73646 151320 73652
rect 151372 71670 151400 79562
rect 151464 73681 151492 79591
rect 151556 77897 151584 79630
rect 151542 77888 151598 77897
rect 151542 77823 151598 77832
rect 151648 76566 151676 79784
rect 151740 79784 151814 79812
rect 152142 79824 152194 79830
rect 151740 78062 151768 79784
rect 152142 79766 152194 79772
rect 152246 79778 152274 80036
rect 152338 79937 152366 80036
rect 152430 79966 152458 80036
rect 152418 79960 152470 79966
rect 152324 79928 152380 79937
rect 152522 79937 152550 80036
rect 152418 79902 152470 79908
rect 152508 79928 152564 79937
rect 152324 79863 152380 79872
rect 152508 79863 152564 79872
rect 151912 79756 151964 79762
rect 151912 79698 151964 79704
rect 152004 79756 152056 79762
rect 152246 79750 152320 79778
rect 152004 79698 152056 79704
rect 151924 78538 151952 79698
rect 151912 78532 151964 78538
rect 151912 78474 151964 78480
rect 151728 78056 151780 78062
rect 151728 77998 151780 78004
rect 151636 76560 151688 76566
rect 151636 76502 151688 76508
rect 152016 75449 152044 79698
rect 152096 79688 152148 79694
rect 152096 79630 152148 79636
rect 152002 75440 152058 75449
rect 152002 75375 152058 75384
rect 151820 74792 151872 74798
rect 151820 74734 151872 74740
rect 151450 73672 151506 73681
rect 151450 73607 151506 73616
rect 151832 72622 151860 74734
rect 151820 72616 151872 72622
rect 151820 72558 151872 72564
rect 151360 71664 151412 71670
rect 151360 71606 151412 71612
rect 151728 71664 151780 71670
rect 151728 71606 151780 71612
rect 151740 71126 151768 71606
rect 151728 71120 151780 71126
rect 151728 71062 151780 71068
rect 151176 70236 151228 70242
rect 151176 70178 151228 70184
rect 150900 48272 150952 48278
rect 150900 48214 150952 48220
rect 150452 16546 151400 16574
rect 149704 11756 149756 11762
rect 149704 11698 149756 11704
rect 147680 6248 147732 6254
rect 147680 6190 147732 6196
rect 144276 3460 144328 3466
rect 144276 3402 144328 3408
rect 146300 3460 146352 3466
rect 146300 3402 146352 3408
rect 147496 3460 147548 3466
rect 147496 3402 147548 3408
rect 144184 3392 144236 3398
rect 144184 3334 144236 3340
rect 140412 3324 140464 3330
rect 140412 3266 140464 3272
rect 140424 480 140452 3266
rect 144288 480 144316 3402
rect 147508 480 147536 3402
rect 151372 480 151400 16546
rect 151832 8294 151860 72558
rect 152108 71774 152136 79630
rect 152188 79620 152240 79626
rect 152188 79562 152240 79568
rect 152200 79529 152228 79562
rect 152186 79520 152242 79529
rect 152186 79455 152242 79464
rect 152292 78878 152320 79750
rect 152464 79756 152516 79762
rect 152464 79698 152516 79704
rect 152280 78872 152332 78878
rect 152280 78814 152332 78820
rect 152372 78260 152424 78266
rect 152372 78202 152424 78208
rect 152384 76072 152412 78202
rect 152292 76044 152412 76072
rect 152292 72962 152320 76044
rect 152476 75993 152504 79698
rect 152614 79676 152642 80036
rect 152706 79744 152734 80036
rect 152798 79898 152826 80036
rect 152786 79892 152838 79898
rect 152786 79834 152838 79840
rect 152890 79812 152918 80036
rect 152982 79966 153010 80036
rect 152970 79960 153022 79966
rect 152970 79902 153022 79908
rect 153074 79830 153102 80036
rect 153166 79971 153194 80036
rect 153152 79962 153208 79971
rect 153152 79897 153208 79906
rect 153258 79898 153286 80036
rect 153246 79892 153298 79898
rect 153246 79834 153298 79840
rect 153062 79824 153114 79830
rect 152890 79784 152964 79812
rect 152706 79716 152780 79744
rect 152614 79648 152688 79676
rect 152554 79384 152610 79393
rect 152554 79319 152610 79328
rect 152462 75984 152518 75993
rect 152372 75948 152424 75954
rect 152462 75919 152518 75928
rect 152372 75890 152424 75896
rect 152280 72956 152332 72962
rect 152280 72898 152332 72904
rect 152108 71746 152228 71774
rect 152200 69630 152228 71746
rect 152384 70394 152412 75890
rect 152464 73908 152516 73914
rect 152464 73850 152516 73856
rect 152476 73166 152504 73850
rect 152464 73160 152516 73166
rect 152464 73102 152516 73108
rect 152384 70366 152504 70394
rect 152188 69624 152240 69630
rect 152188 69566 152240 69572
rect 151912 63232 151964 63238
rect 151912 63174 151964 63180
rect 151924 56642 151952 63174
rect 151912 56636 151964 56642
rect 151912 56578 151964 56584
rect 152476 33114 152504 70366
rect 152568 63238 152596 79319
rect 152660 74322 152688 79648
rect 152648 74316 152700 74322
rect 152648 74258 152700 74264
rect 152752 70394 152780 79716
rect 152832 79688 152884 79694
rect 152832 79630 152884 79636
rect 152844 78033 152872 79630
rect 152936 78266 152964 79784
rect 153062 79766 153114 79772
rect 153350 79744 153378 80036
rect 153442 79898 153470 80036
rect 153430 79892 153482 79898
rect 153430 79834 153482 79840
rect 153534 79778 153562 80036
rect 153626 79966 153654 80036
rect 153614 79960 153666 79966
rect 153614 79902 153666 79908
rect 153488 79750 153562 79778
rect 153350 79716 153424 79744
rect 153016 79620 153068 79626
rect 153016 79562 153068 79568
rect 153292 79620 153344 79626
rect 153292 79562 153344 79568
rect 152924 78260 152976 78266
rect 152924 78202 152976 78208
rect 152830 78024 152886 78033
rect 152830 77959 152886 77968
rect 153028 72894 153056 79562
rect 153108 79552 153160 79558
rect 153108 79494 153160 79500
rect 153200 79552 153252 79558
rect 153200 79494 153252 79500
rect 153120 75818 153148 79494
rect 153212 76906 153240 79494
rect 153304 78742 153332 79562
rect 153292 78736 153344 78742
rect 153292 78678 153344 78684
rect 153396 77294 153424 79716
rect 153488 79558 153516 79750
rect 153718 79744 153746 80036
rect 153810 79801 153838 80036
rect 153902 79830 153930 80036
rect 153994 79971 154022 80036
rect 153980 79962 154036 79971
rect 153980 79897 154036 79906
rect 154086 79830 154114 80036
rect 154178 79937 154206 80036
rect 154270 79966 154298 80036
rect 154362 79966 154390 80036
rect 154454 79966 154482 80036
rect 154258 79960 154310 79966
rect 154164 79928 154220 79937
rect 154258 79902 154310 79908
rect 154350 79960 154402 79966
rect 154350 79902 154402 79908
rect 154442 79960 154494 79966
rect 154442 79902 154494 79908
rect 154164 79863 154220 79872
rect 153890 79824 153942 79830
rect 153672 79716 153746 79744
rect 153796 79792 153852 79801
rect 153890 79766 153942 79772
rect 154074 79824 154126 79830
rect 154074 79766 154126 79772
rect 154212 79824 154264 79830
rect 154442 79824 154494 79830
rect 154212 79766 154264 79772
rect 154362 79772 154442 79778
rect 154362 79766 154494 79772
rect 153796 79727 153852 79736
rect 153568 79688 153620 79694
rect 153568 79630 153620 79636
rect 153476 79552 153528 79558
rect 153476 79494 153528 79500
rect 153396 77266 153516 77294
rect 153200 76900 153252 76906
rect 153200 76842 153252 76848
rect 153108 75812 153160 75818
rect 153108 75754 153160 75760
rect 153384 73364 153436 73370
rect 153384 73306 153436 73312
rect 153016 72888 153068 72894
rect 153016 72830 153068 72836
rect 153108 71256 153160 71262
rect 153108 71198 153160 71204
rect 152752 70366 152964 70394
rect 152936 70106 152964 70366
rect 152924 70100 152976 70106
rect 152924 70042 152976 70048
rect 153120 68202 153148 71198
rect 153108 68196 153160 68202
rect 153108 68138 153160 68144
rect 153396 63306 153424 73306
rect 153488 67386 153516 77266
rect 153580 72690 153608 79630
rect 153672 74225 153700 79716
rect 154120 79688 154172 79694
rect 153750 79656 153806 79665
rect 153934 79656 153990 79665
rect 153750 79591 153806 79600
rect 153844 79620 153896 79626
rect 153764 75138 153792 79591
rect 154120 79630 154172 79636
rect 153934 79591 153990 79600
rect 153844 79562 153896 79568
rect 153856 75857 153884 79562
rect 153948 76430 153976 79591
rect 154028 78668 154080 78674
rect 154028 78610 154080 78616
rect 153936 76424 153988 76430
rect 153936 76366 153988 76372
rect 153842 75848 153898 75857
rect 153842 75783 153898 75792
rect 153752 75132 153804 75138
rect 153752 75074 153804 75080
rect 153658 74216 153714 74225
rect 153658 74151 153714 74160
rect 153934 73944 153990 73953
rect 153934 73879 153990 73888
rect 153568 72684 153620 72690
rect 153568 72626 153620 72632
rect 153476 67380 153528 67386
rect 153476 67322 153528 67328
rect 153384 63300 153436 63306
rect 153384 63242 153436 63248
rect 152556 63232 152608 63238
rect 152556 63174 152608 63180
rect 153396 62150 153424 63242
rect 153384 62144 153436 62150
rect 153384 62086 153436 62092
rect 153844 62144 153896 62150
rect 153844 62086 153896 62092
rect 152464 33108 152516 33114
rect 152464 33050 152516 33056
rect 153856 14618 153884 62086
rect 153948 45558 153976 73879
rect 154040 73370 154068 78610
rect 154132 77654 154160 79630
rect 154120 77648 154172 77654
rect 154120 77590 154172 77596
rect 154224 74798 154252 79766
rect 154362 79750 154482 79766
rect 154362 79676 154390 79750
rect 154316 79648 154390 79676
rect 154212 74792 154264 74798
rect 154212 74734 154264 74740
rect 154028 73364 154080 73370
rect 154028 73306 154080 73312
rect 154316 70394 154344 79648
rect 154546 79642 154574 80036
rect 154638 79744 154666 80036
rect 154730 79971 154758 80036
rect 154716 79962 154772 79971
rect 154716 79897 154772 79906
rect 154822 79744 154850 80036
rect 154914 79971 154942 80036
rect 154900 79962 154956 79971
rect 155006 79966 155034 80036
rect 154900 79897 154956 79906
rect 154994 79960 155046 79966
rect 155098 79937 155126 80036
rect 155190 79966 155218 80036
rect 155178 79960 155230 79966
rect 154994 79902 155046 79908
rect 155084 79928 155140 79937
rect 155178 79902 155230 79908
rect 155282 79898 155310 80036
rect 155374 79937 155402 80036
rect 155360 79928 155416 79937
rect 155084 79863 155140 79872
rect 155270 79892 155322 79898
rect 155360 79863 155416 79872
rect 155270 79834 155322 79840
rect 155222 79792 155278 79801
rect 154948 79756 155000 79762
rect 154638 79716 154712 79744
rect 154822 79716 154896 79744
rect 154684 79665 154712 79716
rect 154500 79614 154574 79642
rect 154670 79656 154726 79665
rect 154396 78736 154448 78742
rect 154396 78678 154448 78684
rect 154040 70366 154344 70394
rect 153936 45552 153988 45558
rect 153936 45494 153988 45500
rect 154040 30326 154068 70366
rect 154408 51814 154436 78678
rect 154500 78674 154528 79614
rect 154670 79591 154726 79600
rect 154672 79484 154724 79490
rect 154592 79444 154672 79472
rect 154592 79150 154620 79444
rect 154868 79472 154896 79716
rect 155466 79778 155494 80036
rect 155222 79727 155278 79736
rect 155316 79756 155368 79762
rect 154948 79698 155000 79704
rect 154672 79426 154724 79432
rect 154776 79444 154896 79472
rect 154672 79280 154724 79286
rect 154672 79222 154724 79228
rect 154580 79144 154632 79150
rect 154580 79086 154632 79092
rect 154488 78668 154540 78674
rect 154488 78610 154540 78616
rect 154578 78568 154634 78577
rect 154578 78503 154634 78512
rect 154592 73710 154620 78503
rect 154684 75993 154712 79222
rect 154670 75984 154726 75993
rect 154670 75919 154726 75928
rect 154672 74248 154724 74254
rect 154672 74190 154724 74196
rect 154580 73704 154632 73710
rect 154580 73646 154632 73652
rect 154684 57934 154712 74190
rect 154776 64802 154804 79444
rect 154854 78568 154910 78577
rect 154854 78503 154910 78512
rect 154868 66094 154896 78503
rect 154960 76786 154988 79698
rect 155132 79688 155184 79694
rect 155132 79630 155184 79636
rect 155144 78334 155172 79630
rect 155132 78328 155184 78334
rect 155132 78270 155184 78276
rect 154960 76758 155080 76786
rect 154948 76696 155000 76702
rect 154948 76638 155000 76644
rect 154856 66088 154908 66094
rect 154856 66030 154908 66036
rect 154960 65793 154988 76638
rect 155052 68134 155080 76758
rect 155132 76492 155184 76498
rect 155132 76434 155184 76440
rect 155144 69601 155172 76434
rect 155236 75954 155264 79727
rect 155316 79698 155368 79704
rect 155420 79750 155494 79778
rect 155328 75993 155356 79698
rect 155314 75984 155370 75993
rect 155224 75948 155276 75954
rect 155314 75919 155370 75928
rect 155224 75890 155276 75896
rect 155420 74254 155448 79750
rect 155558 79676 155586 80036
rect 155650 79898 155678 80036
rect 155742 79903 155770 80036
rect 155834 79966 155862 80036
rect 155822 79960 155874 79966
rect 155638 79892 155690 79898
rect 155638 79834 155690 79840
rect 155728 79894 155784 79903
rect 155822 79902 155874 79908
rect 155926 79898 155954 80036
rect 156018 79898 156046 80036
rect 156110 79971 156138 80036
rect 156096 79962 156152 79971
rect 156202 79966 156230 80036
rect 155728 79829 155784 79838
rect 155914 79892 155966 79898
rect 155914 79834 155966 79840
rect 156006 79892 156058 79898
rect 156096 79897 156152 79906
rect 156190 79960 156242 79966
rect 156294 79937 156322 80036
rect 156190 79902 156242 79908
rect 156280 79928 156336 79937
rect 156280 79863 156336 79872
rect 156006 79834 156058 79840
rect 156236 79824 156288 79830
rect 156236 79766 156288 79772
rect 155776 79756 155828 79762
rect 155776 79698 155828 79704
rect 156144 79756 156196 79762
rect 156144 79698 156196 79704
rect 155512 79648 155586 79676
rect 155682 79656 155738 79665
rect 155512 79393 155540 79648
rect 155682 79591 155738 79600
rect 155498 79384 155554 79393
rect 155498 79319 155554 79328
rect 155592 79144 155644 79150
rect 155592 79086 155644 79092
rect 155498 77888 155554 77897
rect 155498 77823 155554 77832
rect 155512 77654 155540 77823
rect 155500 77648 155552 77654
rect 155500 77590 155552 77596
rect 155408 74248 155460 74254
rect 155408 74190 155460 74196
rect 155604 72418 155632 79086
rect 155592 72412 155644 72418
rect 155592 72354 155644 72360
rect 155696 70394 155724 79591
rect 155788 76702 155816 79698
rect 155868 79688 155920 79694
rect 155868 79630 155920 79636
rect 156050 79656 156106 79665
rect 155776 76696 155828 76702
rect 155776 76638 155828 76644
rect 155880 76498 155908 79630
rect 155960 79620 156012 79626
rect 156050 79591 156106 79600
rect 155960 79562 156012 79568
rect 155972 76566 156000 79562
rect 155960 76560 156012 76566
rect 155960 76502 156012 76508
rect 155868 76492 155920 76498
rect 155868 76434 155920 76440
rect 156064 75682 156092 79591
rect 156156 76673 156184 79698
rect 156142 76664 156198 76673
rect 156142 76599 156198 76608
rect 156248 76401 156276 79766
rect 156386 79744 156414 80036
rect 156340 79716 156414 79744
rect 156234 76392 156290 76401
rect 156234 76327 156290 76336
rect 156340 76242 156368 79716
rect 156478 79676 156506 80036
rect 156570 79812 156598 80036
rect 156662 79966 156690 80036
rect 156650 79960 156702 79966
rect 156650 79902 156702 79908
rect 156754 79898 156782 80036
rect 156846 79898 156874 80036
rect 156938 79966 156966 80036
rect 157030 79966 157058 80036
rect 157122 79966 157150 80036
rect 157214 79966 157242 80036
rect 157306 79971 157334 80036
rect 156926 79960 156978 79966
rect 156926 79902 156978 79908
rect 157018 79960 157070 79966
rect 157018 79902 157070 79908
rect 157110 79960 157162 79966
rect 157110 79902 157162 79908
rect 157202 79960 157254 79966
rect 157202 79902 157254 79908
rect 157292 79962 157348 79971
rect 157398 79966 157426 80036
rect 157490 79966 157518 80036
rect 156742 79892 156794 79898
rect 156742 79834 156794 79840
rect 156834 79892 156886 79898
rect 157292 79897 157348 79906
rect 157386 79960 157438 79966
rect 157386 79902 157438 79908
rect 157478 79960 157530 79966
rect 157478 79902 157530 79908
rect 157582 79898 157610 80036
rect 157674 79966 157702 80036
rect 157662 79960 157714 79966
rect 157766 79937 157794 80036
rect 157662 79902 157714 79908
rect 157752 79928 157808 79937
rect 156834 79834 156886 79840
rect 157570 79892 157622 79898
rect 157752 79863 157808 79872
rect 157016 79826 157072 79835
rect 157570 79834 157622 79840
rect 156570 79784 156690 79812
rect 156662 79676 156690 79784
rect 157016 79761 157072 79770
rect 157708 79824 157760 79830
rect 157708 79766 157760 79772
rect 157340 79756 157392 79762
rect 157340 79698 157392 79704
rect 157524 79756 157576 79762
rect 157524 79698 157576 79704
rect 156478 79648 156552 79676
rect 156420 79552 156472 79558
rect 156420 79494 156472 79500
rect 156156 76214 156368 76242
rect 156052 75676 156104 75682
rect 156052 75618 156104 75624
rect 155604 70366 155724 70394
rect 155130 69592 155186 69601
rect 155130 69527 155186 69536
rect 155040 68128 155092 68134
rect 155040 68070 155092 68076
rect 154946 65784 155002 65793
rect 154946 65719 155002 65728
rect 154764 64796 154816 64802
rect 154764 64738 154816 64744
rect 154672 57928 154724 57934
rect 154672 57870 154724 57876
rect 154396 51808 154448 51814
rect 154396 51750 154448 51756
rect 155604 38622 155632 70366
rect 155868 68808 155920 68814
rect 155868 68750 155920 68756
rect 155880 68134 155908 68750
rect 155868 68128 155920 68134
rect 155868 68070 155920 68076
rect 156156 66774 156184 76214
rect 156236 76152 156288 76158
rect 156236 76094 156288 76100
rect 156248 68882 156276 76094
rect 156432 73154 156460 79494
rect 156340 73126 156460 73154
rect 156340 70922 156368 73126
rect 156524 72962 156552 79648
rect 156616 79648 156690 79676
rect 156972 79688 157024 79694
rect 156512 72956 156564 72962
rect 156512 72898 156564 72904
rect 156328 70916 156380 70922
rect 156328 70858 156380 70864
rect 156236 68876 156288 68882
rect 156236 68818 156288 68824
rect 156248 68066 156276 68818
rect 156236 68060 156288 68066
rect 156236 68002 156288 68008
rect 156144 66768 156196 66774
rect 156144 66710 156196 66716
rect 156340 64874 156368 70858
rect 156616 70394 156644 79648
rect 156972 79630 157024 79636
rect 157064 79688 157116 79694
rect 157064 79630 157116 79636
rect 157156 79688 157208 79694
rect 157156 79630 157208 79636
rect 156880 79620 156932 79626
rect 156880 79562 156932 79568
rect 156788 79552 156840 79558
rect 156788 79494 156840 79500
rect 156696 77240 156748 77246
rect 156696 77182 156748 77188
rect 156708 76974 156736 77182
rect 156696 76968 156748 76974
rect 156696 76910 156748 76916
rect 156800 76838 156828 79494
rect 156788 76832 156840 76838
rect 156788 76774 156840 76780
rect 156788 76696 156840 76702
rect 156788 76638 156840 76644
rect 156616 70366 156736 70394
rect 156708 70038 156736 70366
rect 156696 70032 156748 70038
rect 156696 69974 156748 69980
rect 156696 68060 156748 68066
rect 156696 68002 156748 68008
rect 156340 64846 156644 64874
rect 155592 38616 155644 38622
rect 155592 38558 155644 38564
rect 154028 30320 154080 30326
rect 154028 30262 154080 30268
rect 153844 14612 153896 14618
rect 153844 14554 153896 14560
rect 151820 8288 151872 8294
rect 151820 8230 151872 8236
rect 155224 4820 155276 4826
rect 155224 4762 155276 4768
rect 155236 480 155264 4762
rect 156616 3602 156644 64846
rect 156708 15910 156736 68002
rect 156800 60654 156828 76638
rect 156892 75970 156920 79562
rect 156984 76158 157012 79630
rect 156972 76152 157024 76158
rect 156972 76094 157024 76100
rect 156892 75942 157012 75970
rect 156880 75676 156932 75682
rect 156880 75618 156932 75624
rect 156892 66026 156920 75618
rect 156984 70990 157012 75942
rect 157076 73154 157104 79630
rect 157168 76702 157196 79630
rect 157156 76696 157208 76702
rect 157156 76638 157208 76644
rect 157352 75886 157380 79698
rect 157432 78804 157484 78810
rect 157432 78746 157484 78752
rect 157340 75880 157392 75886
rect 157340 75822 157392 75828
rect 157340 75676 157392 75682
rect 157340 75618 157392 75624
rect 157076 73126 157196 73154
rect 157168 73030 157196 73126
rect 157156 73024 157208 73030
rect 157156 72966 157208 72972
rect 156972 70984 157024 70990
rect 156972 70926 157024 70932
rect 157352 66162 157380 75618
rect 157444 72282 157472 78746
rect 157536 77994 157564 79698
rect 157616 79688 157668 79694
rect 157616 79630 157668 79636
rect 157524 77988 157576 77994
rect 157524 77930 157576 77936
rect 157628 76616 157656 79630
rect 157536 76588 157656 76616
rect 157432 72276 157484 72282
rect 157432 72218 157484 72224
rect 157444 71058 157472 72218
rect 157432 71052 157484 71058
rect 157432 70994 157484 71000
rect 157536 67522 157564 76588
rect 157616 75880 157668 75886
rect 157616 75822 157668 75828
rect 157628 70106 157656 75822
rect 157720 74458 157748 79766
rect 157858 79744 157886 80036
rect 157950 79971 157978 80036
rect 157936 79962 157992 79971
rect 157936 79897 157992 79906
rect 157812 79716 157886 79744
rect 158042 79744 158070 80036
rect 158134 79812 158162 80036
rect 158226 79966 158254 80036
rect 158318 79966 158346 80036
rect 158214 79960 158266 79966
rect 158214 79902 158266 79908
rect 158306 79960 158358 79966
rect 158306 79902 158358 79908
rect 158134 79784 158208 79812
rect 158180 79778 158208 79784
rect 158180 79750 158254 79778
rect 158042 79716 158116 79744
rect 157812 76702 157840 79716
rect 157982 79656 158038 79665
rect 157892 79620 157944 79626
rect 157982 79591 158038 79600
rect 157892 79562 157944 79568
rect 157904 78198 157932 79562
rect 157892 78192 157944 78198
rect 157892 78134 157944 78140
rect 157996 77926 158024 79591
rect 157984 77920 158036 77926
rect 157984 77862 158036 77868
rect 157800 76696 157852 76702
rect 157800 76638 157852 76644
rect 158088 75682 158116 79716
rect 158226 79676 158254 79750
rect 158410 79744 158438 80036
rect 158502 79898 158530 80036
rect 158594 79898 158622 80036
rect 158686 79937 158714 80036
rect 158672 79928 158728 79937
rect 158490 79892 158542 79898
rect 158490 79834 158542 79840
rect 158582 79892 158634 79898
rect 158672 79863 158728 79872
rect 158582 79834 158634 79840
rect 158536 79756 158588 79762
rect 158410 79716 158484 79744
rect 158180 79648 158254 79676
rect 158180 78810 158208 79648
rect 158260 79552 158312 79558
rect 158260 79494 158312 79500
rect 158168 78804 158220 78810
rect 158168 78746 158220 78752
rect 158272 76072 158300 79494
rect 158456 77294 158484 79716
rect 158778 79744 158806 80036
rect 158870 79778 158898 80036
rect 158962 79898 158990 80036
rect 158950 79892 159002 79898
rect 158950 79834 159002 79840
rect 159054 79778 159082 80036
rect 159146 79966 159174 80036
rect 159238 79966 159266 80172
rect 177776 80102 177804 80310
rect 178316 80300 178368 80306
rect 178316 80242 178368 80248
rect 178040 80164 178092 80170
rect 178040 80106 178092 80112
rect 178132 80164 178184 80170
rect 178132 80106 178184 80112
rect 177764 80096 177816 80102
rect 177764 80038 177816 80044
rect 177946 80064 178002 80073
rect 159330 79966 159358 80036
rect 159134 79960 159186 79966
rect 159134 79902 159186 79908
rect 159226 79960 159278 79966
rect 159226 79902 159278 79908
rect 159318 79960 159370 79966
rect 159318 79902 159370 79908
rect 159422 79812 159450 80036
rect 159514 79966 159542 80036
rect 159606 79971 159634 80036
rect 159502 79960 159554 79966
rect 159502 79902 159554 79908
rect 159592 79962 159648 79971
rect 159592 79897 159648 79906
rect 159376 79784 159450 79812
rect 158870 79750 158944 79778
rect 159054 79750 159128 79778
rect 158536 79698 158588 79704
rect 158732 79716 158806 79744
rect 158548 78130 158576 79698
rect 158536 78124 158588 78130
rect 158536 78066 158588 78072
rect 158626 77752 158682 77761
rect 158626 77687 158682 77696
rect 158456 77266 158576 77294
rect 158444 76696 158496 76702
rect 158444 76638 158496 76644
rect 158180 76044 158300 76072
rect 158076 75676 158128 75682
rect 158076 75618 158128 75624
rect 157708 74452 157760 74458
rect 157708 74394 157760 74400
rect 158180 70394 158208 76044
rect 158260 75948 158312 75954
rect 158260 75890 158312 75896
rect 157720 70366 158208 70394
rect 157616 70100 157668 70106
rect 157616 70042 157668 70048
rect 157720 69834 157748 70366
rect 157708 69828 157760 69834
rect 157708 69770 157760 69776
rect 157524 67516 157576 67522
rect 157524 67458 157576 67464
rect 157340 66156 157392 66162
rect 157340 66098 157392 66104
rect 156880 66020 156932 66026
rect 156880 65962 156932 65968
rect 156892 64874 156920 65962
rect 156892 64846 157288 64874
rect 156788 60648 156840 60654
rect 156788 60590 156840 60596
rect 156696 15904 156748 15910
rect 156696 15846 156748 15852
rect 157260 10334 157288 64846
rect 158272 41410 158300 75890
rect 158352 72684 158404 72690
rect 158352 72626 158404 72632
rect 158364 65414 158392 72626
rect 158352 65408 158404 65414
rect 158352 65350 158404 65356
rect 158456 57866 158484 76638
rect 158548 76498 158576 77266
rect 158536 76492 158588 76498
rect 158536 76434 158588 76440
rect 158640 71738 158668 77687
rect 158732 75410 158760 79716
rect 158916 79540 158944 79750
rect 158994 79656 159050 79665
rect 158994 79591 159050 79600
rect 158824 79512 158944 79540
rect 158824 75478 158852 79512
rect 158904 79416 158956 79422
rect 158904 79358 158956 79364
rect 158812 75472 158864 75478
rect 158812 75414 158864 75420
rect 158720 75404 158772 75410
rect 158720 75346 158772 75352
rect 158812 75336 158864 75342
rect 158812 75278 158864 75284
rect 158720 75268 158772 75274
rect 158720 75210 158772 75216
rect 158628 71732 158680 71738
rect 158628 71674 158680 71680
rect 158536 70100 158588 70106
rect 158536 70042 158588 70048
rect 158444 57860 158496 57866
rect 158444 57802 158496 57808
rect 158260 41404 158312 41410
rect 158260 41346 158312 41352
rect 158548 35290 158576 70042
rect 158628 69828 158680 69834
rect 158628 69770 158680 69776
rect 158536 35284 158588 35290
rect 158536 35226 158588 35232
rect 157248 10328 157300 10334
rect 157248 10270 157300 10276
rect 158640 6254 158668 69770
rect 158732 34474 158760 75210
rect 158824 63510 158852 75278
rect 158916 64598 158944 79358
rect 159008 75274 159036 79591
rect 159100 77518 159128 79750
rect 159376 79744 159404 79784
rect 159548 79756 159600 79762
rect 159376 79716 159496 79744
rect 159272 79688 159324 79694
rect 159272 79630 159324 79636
rect 159180 79620 159232 79626
rect 159180 79562 159232 79568
rect 159088 77512 159140 77518
rect 159088 77454 159140 77460
rect 159088 75472 159140 75478
rect 159088 75414 159140 75420
rect 158996 75268 159048 75274
rect 158996 75210 159048 75216
rect 158996 75064 159048 75070
rect 158996 75006 159048 75012
rect 159008 66230 159036 75006
rect 159100 67425 159128 75414
rect 159192 68610 159220 79562
rect 159284 76974 159312 79630
rect 159364 79416 159416 79422
rect 159364 79358 159416 79364
rect 159376 79218 159404 79358
rect 159364 79212 159416 79218
rect 159364 79154 159416 79160
rect 159468 78985 159496 79716
rect 159548 79698 159600 79704
rect 159454 78976 159510 78985
rect 159454 78911 159510 78920
rect 159560 78674 159588 79698
rect 159698 79642 159726 80036
rect 159790 79971 159818 80036
rect 159776 79962 159832 79971
rect 159882 79966 159910 80036
rect 159776 79897 159832 79906
rect 159870 79960 159922 79966
rect 159870 79902 159922 79908
rect 159974 79898 160002 80036
rect 160066 79898 160094 80036
rect 160158 79971 160186 80036
rect 160144 79962 160200 79971
rect 160250 79966 160278 80036
rect 159962 79892 160014 79898
rect 159962 79834 160014 79840
rect 160054 79892 160106 79898
rect 160144 79897 160200 79906
rect 160238 79960 160290 79966
rect 160342 79937 160370 80036
rect 160434 79966 160462 80036
rect 160422 79960 160474 79966
rect 160238 79902 160290 79908
rect 160328 79928 160384 79937
rect 160422 79902 160474 79908
rect 160526 79898 160554 80036
rect 160618 79937 160646 80036
rect 160710 79966 160738 80036
rect 160802 79971 160830 80036
rect 160698 79960 160750 79966
rect 160604 79928 160660 79937
rect 160328 79863 160384 79872
rect 160514 79892 160566 79898
rect 160054 79834 160106 79840
rect 160698 79902 160750 79908
rect 160788 79962 160844 79971
rect 160788 79897 160844 79906
rect 160604 79863 160660 79872
rect 160514 79834 160566 79840
rect 160652 79824 160704 79830
rect 160894 79812 160922 80036
rect 160986 79966 161014 80036
rect 161078 79971 161106 80036
rect 160974 79960 161026 79966
rect 160974 79902 161026 79908
rect 161064 79962 161120 79971
rect 161064 79897 161120 79906
rect 161170 79898 161198 80036
rect 161158 79892 161210 79898
rect 161158 79834 161210 79840
rect 161262 79830 161290 80036
rect 161354 79971 161382 80036
rect 161340 79962 161396 79971
rect 161340 79897 161396 79906
rect 160652 79766 160704 79772
rect 160756 79784 160922 79812
rect 161250 79824 161302 79830
rect 161018 79792 161074 79801
rect 160008 79756 160060 79762
rect 160008 79698 160060 79704
rect 160560 79756 160612 79762
rect 160560 79698 160612 79704
rect 159914 79656 159970 79665
rect 159698 79614 159772 79642
rect 159548 78668 159600 78674
rect 159548 78610 159600 78616
rect 159272 76968 159324 76974
rect 159272 76910 159324 76916
rect 159272 75404 159324 75410
rect 159272 75346 159324 75352
rect 159180 68604 159232 68610
rect 159180 68546 159232 68552
rect 159284 68542 159312 75346
rect 159744 75342 159772 79614
rect 159824 79620 159876 79626
rect 159914 79591 159970 79600
rect 159824 79562 159876 79568
rect 159732 75336 159784 75342
rect 159732 75278 159784 75284
rect 159836 75041 159864 79562
rect 159822 75032 159878 75041
rect 159822 74967 159878 74976
rect 159928 72554 159956 79591
rect 160020 75070 160048 79698
rect 160100 79688 160152 79694
rect 160284 79688 160336 79694
rect 160100 79630 160152 79636
rect 160190 79656 160246 79665
rect 160112 76906 160140 79630
rect 160284 79630 160336 79636
rect 160190 79591 160246 79600
rect 160100 76900 160152 76906
rect 160100 76842 160152 76848
rect 160100 76696 160152 76702
rect 160100 76638 160152 76644
rect 160008 75064 160060 75070
rect 160008 75006 160060 75012
rect 159916 72548 159968 72554
rect 159916 72490 159968 72496
rect 159272 68536 159324 68542
rect 159272 68478 159324 68484
rect 159086 67416 159142 67425
rect 159086 67351 159142 67360
rect 158996 66224 159048 66230
rect 158996 66166 159048 66172
rect 160112 65754 160140 76638
rect 160204 68950 160232 79591
rect 160296 70038 160324 79630
rect 160376 79484 160428 79490
rect 160376 79426 160428 79432
rect 160388 76702 160416 79426
rect 160572 79354 160600 79698
rect 160468 79348 160520 79354
rect 160468 79290 160520 79296
rect 160560 79348 160612 79354
rect 160560 79290 160612 79296
rect 160376 76696 160428 76702
rect 160376 76638 160428 76644
rect 160376 75676 160428 75682
rect 160376 75618 160428 75624
rect 160284 70032 160336 70038
rect 160284 69974 160336 69980
rect 160388 69630 160416 75618
rect 160480 73681 160508 79290
rect 160664 77217 160692 79766
rect 160756 79558 160784 79784
rect 161446 79778 161474 80036
rect 161538 79830 161566 80036
rect 161630 79966 161658 80036
rect 161722 79966 161750 80036
rect 161814 79971 161842 80036
rect 161618 79960 161670 79966
rect 161618 79902 161670 79908
rect 161710 79960 161762 79966
rect 161710 79902 161762 79908
rect 161800 79962 161856 79971
rect 161906 79966 161934 80036
rect 161998 79971 162026 80036
rect 161800 79897 161856 79906
rect 161894 79960 161946 79966
rect 161894 79902 161946 79908
rect 161984 79962 162040 79971
rect 162090 79966 162118 80036
rect 162182 79966 162210 80036
rect 162274 79966 162302 80036
rect 161984 79897 162040 79906
rect 162078 79960 162130 79966
rect 162078 79902 162130 79908
rect 162170 79960 162222 79966
rect 162170 79902 162222 79908
rect 162262 79960 162314 79966
rect 162262 79902 162314 79908
rect 161250 79766 161302 79772
rect 161018 79727 161074 79736
rect 161400 79750 161474 79778
rect 161526 79824 161578 79830
rect 161940 79824 161992 79830
rect 161526 79766 161578 79772
rect 161846 79792 161902 79801
rect 161756 79756 161808 79762
rect 160928 79688 160980 79694
rect 160928 79630 160980 79636
rect 160744 79552 160796 79558
rect 160744 79494 160796 79500
rect 160940 78946 160968 79630
rect 160928 78940 160980 78946
rect 160928 78882 160980 78888
rect 160650 77208 160706 77217
rect 160650 77143 160706 77152
rect 161032 76809 161060 79727
rect 161204 79688 161256 79694
rect 161204 79630 161256 79636
rect 161294 79656 161350 79665
rect 161112 79552 161164 79558
rect 161112 79494 161164 79500
rect 161018 76800 161074 76809
rect 161018 76735 161074 76744
rect 160466 73672 160522 73681
rect 160466 73607 160522 73616
rect 161124 72350 161152 79494
rect 161216 75682 161244 79630
rect 161294 79591 161350 79600
rect 161204 75676 161256 75682
rect 161204 75618 161256 75624
rect 161308 73846 161336 79591
rect 161296 73840 161348 73846
rect 161296 73782 161348 73788
rect 161400 72894 161428 79750
rect 162366 79812 162394 80036
rect 161940 79766 161992 79772
rect 162122 79792 162178 79801
rect 161846 79727 161902 79736
rect 161756 79698 161808 79704
rect 161480 79688 161532 79694
rect 161480 79630 161532 79636
rect 161492 74361 161520 79630
rect 161664 79620 161716 79626
rect 161664 79562 161716 79568
rect 161572 75268 161624 75274
rect 161572 75210 161624 75216
rect 161478 74352 161534 74361
rect 161478 74287 161534 74296
rect 161480 74248 161532 74254
rect 161480 74190 161532 74196
rect 161388 72888 161440 72894
rect 161388 72830 161440 72836
rect 161112 72344 161164 72350
rect 161112 72286 161164 72292
rect 161400 70786 161428 72830
rect 160468 70780 160520 70786
rect 160468 70722 160520 70728
rect 161388 70780 161440 70786
rect 161388 70722 161440 70728
rect 160480 69698 160508 70722
rect 161204 70032 161256 70038
rect 161204 69974 161256 69980
rect 160468 69692 160520 69698
rect 160468 69634 160520 69640
rect 160376 69624 160428 69630
rect 160376 69566 160428 69572
rect 160192 68944 160244 68950
rect 160192 68886 160244 68892
rect 160100 65748 160152 65754
rect 160100 65690 160152 65696
rect 158904 64592 158956 64598
rect 158904 64534 158956 64540
rect 158812 63504 158864 63510
rect 158812 63446 158864 63452
rect 158720 34468 158772 34474
rect 158720 34410 158772 34416
rect 161216 31142 161244 69974
rect 161388 69624 161440 69630
rect 161388 69566 161440 69572
rect 161294 65784 161350 65793
rect 161294 65719 161350 65728
rect 161308 65521 161336 65719
rect 161294 65512 161350 65521
rect 161294 65447 161350 65456
rect 161204 31136 161256 31142
rect 161204 31078 161256 31084
rect 161308 20670 161336 65447
rect 161296 20664 161348 20670
rect 161296 20606 161348 20612
rect 161400 17270 161428 69566
rect 161492 34406 161520 74190
rect 161584 62082 161612 75210
rect 161676 64569 161704 79562
rect 161768 78878 161796 79698
rect 161756 78872 161808 78878
rect 161756 78814 161808 78820
rect 161754 78568 161810 78577
rect 161754 78503 161810 78512
rect 161768 66978 161796 78503
rect 161860 68678 161888 79727
rect 161952 79665 161980 79766
rect 162320 79784 162394 79812
rect 162122 79727 162178 79736
rect 162216 79756 162268 79762
rect 162032 79688 162084 79694
rect 161938 79656 161994 79665
rect 162032 79630 162084 79636
rect 161938 79591 161994 79600
rect 161940 79552 161992 79558
rect 161940 79494 161992 79500
rect 161848 68672 161900 68678
rect 161848 68614 161900 68620
rect 161952 68513 161980 79494
rect 162044 69018 162072 79630
rect 162136 75750 162164 79727
rect 162216 79698 162268 79704
rect 162124 75744 162176 75750
rect 162124 75686 162176 75692
rect 162228 75274 162256 79698
rect 162216 75268 162268 75274
rect 162216 75210 162268 75216
rect 162320 70394 162348 79784
rect 162458 79778 162486 80036
rect 162550 79971 162578 80036
rect 162536 79962 162592 79971
rect 162536 79897 162592 79906
rect 162642 79898 162670 80036
rect 162734 79971 162762 80036
rect 162720 79962 162776 79971
rect 162630 79892 162682 79898
rect 162720 79897 162776 79906
rect 162630 79834 162682 79840
rect 162826 79830 162854 80036
rect 162918 79937 162946 80036
rect 163010 79966 163038 80036
rect 162998 79960 163050 79966
rect 162904 79928 162960 79937
rect 162998 79902 163050 79908
rect 162904 79863 162960 79872
rect 162814 79824 162866 79830
rect 162458 79750 162532 79778
rect 163102 79801 163130 80036
rect 163194 79898 163222 80036
rect 163286 79937 163314 80036
rect 163272 79928 163328 79937
rect 163182 79892 163234 79898
rect 163272 79863 163328 79872
rect 163182 79834 163234 79840
rect 162814 79766 162866 79772
rect 163088 79792 163144 79801
rect 162504 74254 162532 79750
rect 163088 79727 163144 79736
rect 163378 79744 163406 80036
rect 163470 79966 163498 80036
rect 163458 79960 163510 79966
rect 163458 79902 163510 79908
rect 163562 79898 163590 80036
rect 163550 79892 163602 79898
rect 163550 79834 163602 79840
rect 163502 79792 163558 79801
rect 163378 79716 163452 79744
rect 163502 79727 163558 79736
rect 162860 79688 162912 79694
rect 162766 79656 162822 79665
rect 162676 79620 162728 79626
rect 162860 79630 162912 79636
rect 162952 79688 163004 79694
rect 162952 79630 163004 79636
rect 163318 79656 163374 79665
rect 162766 79591 162822 79600
rect 162676 79562 162728 79568
rect 162584 77512 162636 77518
rect 162584 77454 162636 77460
rect 162596 74934 162624 77454
rect 162688 75954 162716 79562
rect 162676 75948 162728 75954
rect 162676 75890 162728 75896
rect 162676 75676 162728 75682
rect 162676 75618 162728 75624
rect 162584 74928 162636 74934
rect 162584 74870 162636 74876
rect 162492 74248 162544 74254
rect 162492 74190 162544 74196
rect 162688 73914 162716 75618
rect 162780 75313 162808 79591
rect 162766 75304 162822 75313
rect 162766 75239 162822 75248
rect 162872 75188 162900 79630
rect 162780 75160 162900 75188
rect 162676 73908 162728 73914
rect 162676 73850 162728 73856
rect 162780 73001 162808 75160
rect 162860 75064 162912 75070
rect 162860 75006 162912 75012
rect 162766 72992 162822 73001
rect 162766 72927 162822 72936
rect 162768 72820 162820 72826
rect 162768 72762 162820 72768
rect 162136 70366 162348 70394
rect 162136 69562 162164 70366
rect 162124 69556 162176 69562
rect 162124 69498 162176 69504
rect 162584 69556 162636 69562
rect 162584 69498 162636 69504
rect 162596 69426 162624 69498
rect 162584 69420 162636 69426
rect 162584 69362 162636 69368
rect 162032 69012 162084 69018
rect 162032 68954 162084 68960
rect 161938 68504 161994 68513
rect 161938 68439 161994 68448
rect 161848 67312 161900 67318
rect 161848 67254 161900 67260
rect 161756 66972 161808 66978
rect 161756 66914 161808 66920
rect 161662 64560 161718 64569
rect 161662 64495 161718 64504
rect 161572 62076 161624 62082
rect 161572 62018 161624 62024
rect 161860 60722 161888 67254
rect 161848 60716 161900 60722
rect 161848 60658 161900 60664
rect 161480 34400 161532 34406
rect 161480 34342 161532 34348
rect 161388 17264 161440 17270
rect 161388 17206 161440 17212
rect 162596 7682 162624 69362
rect 162676 69012 162728 69018
rect 162676 68954 162728 68960
rect 162688 68270 162716 68954
rect 162676 68264 162728 68270
rect 162676 68206 162728 68212
rect 162688 25566 162716 68206
rect 162780 63510 162808 72762
rect 162768 63504 162820 63510
rect 162768 63446 162820 63452
rect 162872 63374 162900 75006
rect 162860 63368 162912 63374
rect 162860 63310 162912 63316
rect 162872 58750 162900 63310
rect 162964 62762 162992 79630
rect 163228 79620 163280 79626
rect 163318 79591 163374 79600
rect 163228 79562 163280 79568
rect 163042 79384 163098 79393
rect 163042 79319 163098 79328
rect 163056 64462 163084 79319
rect 163134 79112 163190 79121
rect 163134 79047 163190 79056
rect 163148 69018 163176 79047
rect 163136 69012 163188 69018
rect 163136 68954 163188 68960
rect 163240 68649 163268 79562
rect 163332 74458 163360 79591
rect 163320 74452 163372 74458
rect 163320 74394 163372 74400
rect 163424 72758 163452 79716
rect 163516 79608 163544 79727
rect 163654 79676 163682 80036
rect 163746 79801 163774 80036
rect 163838 79830 163866 80036
rect 163930 79830 163958 80036
rect 164022 79971 164050 80036
rect 164008 79962 164064 79971
rect 164114 79966 164142 80036
rect 164206 79971 164234 80036
rect 164008 79897 164064 79906
rect 164102 79960 164154 79966
rect 164102 79902 164154 79908
rect 164192 79962 164248 79971
rect 164192 79897 164248 79906
rect 163826 79824 163878 79830
rect 163732 79792 163788 79801
rect 163826 79766 163878 79772
rect 163918 79824 163970 79830
rect 164298 79801 164326 80036
rect 163918 79766 163970 79772
rect 164284 79792 164340 79801
rect 163732 79727 163788 79736
rect 164284 79727 164340 79736
rect 163872 79688 163924 79694
rect 163654 79648 163820 79676
rect 163516 79580 163636 79608
rect 163504 77240 163556 77246
rect 163504 77182 163556 77188
rect 163516 75070 163544 77182
rect 163504 75064 163556 75070
rect 163504 75006 163556 75012
rect 163412 72752 163464 72758
rect 163412 72694 163464 72700
rect 163608 70394 163636 79580
rect 163688 79552 163740 79558
rect 163688 79494 163740 79500
rect 163700 76158 163728 79494
rect 163688 76152 163740 76158
rect 163688 76094 163740 76100
rect 163792 74118 163820 79648
rect 164390 79676 164418 80036
rect 164482 79898 164510 80036
rect 164574 79966 164602 80036
rect 164666 79971 164694 80036
rect 164562 79960 164614 79966
rect 164562 79902 164614 79908
rect 164652 79962 164708 79971
rect 164470 79892 164522 79898
rect 164652 79897 164708 79906
rect 164470 79834 164522 79840
rect 164758 79778 164786 80036
rect 164850 79966 164878 80036
rect 164942 79971 164970 80036
rect 164838 79960 164890 79966
rect 164838 79902 164890 79908
rect 164928 79962 164984 79971
rect 164928 79897 164984 79906
rect 164608 79756 164660 79762
rect 163872 79630 163924 79636
rect 164344 79648 164418 79676
rect 164528 79716 164608 79744
rect 163780 74112 163832 74118
rect 163780 74054 163832 74060
rect 163884 72865 163912 79630
rect 163964 79620 164016 79626
rect 163964 79562 164016 79568
rect 164148 79620 164200 79626
rect 164148 79562 164200 79568
rect 163870 72856 163926 72865
rect 163976 72826 164004 79562
rect 164056 79484 164108 79490
rect 164056 79426 164108 79432
rect 163870 72791 163926 72800
rect 163964 72820 164016 72826
rect 163964 72762 164016 72768
rect 163332 70366 163636 70394
rect 164068 70394 164096 79426
rect 164160 77246 164188 79562
rect 164238 79520 164294 79529
rect 164238 79455 164294 79464
rect 164148 77240 164200 77246
rect 164148 77182 164200 77188
rect 164148 76900 164200 76906
rect 164148 76842 164200 76848
rect 164160 73953 164188 76842
rect 164146 73944 164202 73953
rect 164146 73879 164202 73888
rect 164068 70366 164188 70394
rect 163226 68640 163282 68649
rect 163226 68575 163282 68584
rect 163332 68202 163360 70366
rect 164160 69494 164188 70366
rect 164148 69488 164200 69494
rect 164148 69430 164200 69436
rect 164056 69012 164108 69018
rect 164056 68954 164108 68960
rect 164068 68746 164096 68954
rect 164056 68740 164108 68746
rect 164056 68682 164108 68688
rect 163320 68196 163372 68202
rect 163320 68138 163372 68144
rect 163044 64456 163096 64462
rect 163044 64398 163096 64404
rect 162952 62756 163004 62762
rect 162952 62698 163004 62704
rect 162860 58744 162912 58750
rect 162860 58686 162912 58692
rect 164068 39438 164096 68682
rect 164056 39432 164108 39438
rect 164056 39374 164108 39380
rect 162676 25560 162728 25566
rect 162676 25502 162728 25508
rect 162952 13252 163004 13258
rect 162952 13194 163004 13200
rect 162584 7676 162636 7682
rect 162584 7618 162636 7624
rect 158628 6248 158680 6254
rect 158628 6190 158680 6196
rect 156604 3596 156656 3602
rect 156604 3538 156656 3544
rect 162964 480 162992 13194
rect 164160 7614 164188 69430
rect 164252 56030 164280 79455
rect 164344 63170 164372 79648
rect 164528 79642 164556 79716
rect 164608 79698 164660 79704
rect 164712 79750 164786 79778
rect 164482 79614 164556 79642
rect 164606 79656 164662 79665
rect 164482 79540 164510 79614
rect 164606 79591 164662 79600
rect 164482 79512 164556 79540
rect 164424 78260 164476 78266
rect 164424 78202 164476 78208
rect 164332 63164 164384 63170
rect 164332 63106 164384 63112
rect 164436 62558 164464 78202
rect 164528 67590 164556 79512
rect 164620 77450 164648 79591
rect 164608 77444 164660 77450
rect 164608 77386 164660 77392
rect 164712 77330 164740 79750
rect 165034 79744 165062 80036
rect 165126 79966 165154 80036
rect 165218 79966 165246 80036
rect 165310 79966 165338 80036
rect 165402 79966 165430 80036
rect 165494 79971 165522 80036
rect 165114 79960 165166 79966
rect 165114 79902 165166 79908
rect 165206 79960 165258 79966
rect 165206 79902 165258 79908
rect 165298 79960 165350 79966
rect 165298 79902 165350 79908
rect 165390 79960 165442 79966
rect 165390 79902 165442 79908
rect 165480 79962 165536 79971
rect 165480 79897 165536 79906
rect 165586 79812 165614 80036
rect 165678 79971 165706 80036
rect 165664 79962 165720 79971
rect 165664 79897 165720 79906
rect 165770 79898 165798 80036
rect 165862 79898 165890 80036
rect 165954 79966 165982 80036
rect 165942 79960 165994 79966
rect 165942 79902 165994 79908
rect 165758 79892 165810 79898
rect 165758 79834 165810 79840
rect 165850 79892 165902 79898
rect 165850 79834 165902 79840
rect 165586 79784 165660 79812
rect 165632 79778 165660 79784
rect 166046 79778 166074 80036
rect 166138 79966 166166 80036
rect 166230 79971 166258 80036
rect 166126 79960 166178 79966
rect 166126 79902 166178 79908
rect 166216 79962 166272 79971
rect 166216 79897 166272 79906
rect 166322 79898 166350 80036
rect 166414 79966 166442 80036
rect 166402 79960 166454 79966
rect 166402 79902 166454 79908
rect 166310 79892 166362 79898
rect 166310 79834 166362 79840
rect 166506 79830 166534 80036
rect 166598 79971 166626 80036
rect 166584 79962 166640 79971
rect 166690 79966 166718 80036
rect 166782 79966 166810 80036
rect 166584 79897 166640 79906
rect 166678 79960 166730 79966
rect 166678 79902 166730 79908
rect 166770 79960 166822 79966
rect 166770 79902 166822 79908
rect 166874 79835 166902 80036
rect 166966 79966 166994 80036
rect 166954 79960 167006 79966
rect 166954 79902 167006 79908
rect 166494 79824 166546 79830
rect 166170 79792 166226 79801
rect 164988 79716 165062 79744
rect 165252 79756 165304 79762
rect 164792 79688 164844 79694
rect 164792 79630 164844 79636
rect 164620 77302 164740 77330
rect 164620 74322 164648 77302
rect 164608 74316 164660 74322
rect 164608 74258 164660 74264
rect 164804 70394 164832 79630
rect 164884 79552 164936 79558
rect 164884 79494 164936 79500
rect 164896 72729 164924 79494
rect 164988 75682 165016 79716
rect 165252 79698 165304 79704
rect 165344 79756 165396 79762
rect 165632 79750 165752 79778
rect 165344 79698 165396 79704
rect 165160 79688 165212 79694
rect 165160 79630 165212 79636
rect 165068 76152 165120 76158
rect 165068 76094 165120 76100
rect 164976 75676 165028 75682
rect 164976 75618 165028 75624
rect 164882 72720 164938 72729
rect 164882 72655 164938 72664
rect 164712 70366 164832 70394
rect 164712 70310 164740 70366
rect 164700 70304 164752 70310
rect 164700 70246 164752 70252
rect 164516 67584 164568 67590
rect 164516 67526 164568 67532
rect 165080 64530 165108 76094
rect 165172 69562 165200 79630
rect 165264 78266 165292 79698
rect 165252 78260 165304 78266
rect 165252 78202 165304 78208
rect 165356 72457 165384 79698
rect 165436 79620 165488 79626
rect 165436 79562 165488 79568
rect 165448 78538 165476 79562
rect 165436 78532 165488 78538
rect 165436 78474 165488 78480
rect 165620 78464 165672 78470
rect 165620 78406 165672 78412
rect 165528 77444 165580 77450
rect 165528 77386 165580 77392
rect 165342 72448 165398 72457
rect 165342 72383 165398 72392
rect 165540 72214 165568 77386
rect 165528 72208 165580 72214
rect 165528 72150 165580 72156
rect 165160 69556 165212 69562
rect 165160 69498 165212 69504
rect 165436 67584 165488 67590
rect 165436 67526 165488 67532
rect 165448 67114 165476 67526
rect 165632 67318 165660 78406
rect 165724 76702 165752 79750
rect 165896 79756 165948 79762
rect 166046 79750 166120 79778
rect 165896 79698 165948 79704
rect 165804 79688 165856 79694
rect 165804 79630 165856 79636
rect 165816 78985 165844 79630
rect 165802 78976 165858 78985
rect 165802 78911 165858 78920
rect 165908 77246 165936 79698
rect 165988 79688 166040 79694
rect 165988 79630 166040 79636
rect 165896 77240 165948 77246
rect 165896 77182 165948 77188
rect 165712 76696 165764 76702
rect 165712 76638 165764 76644
rect 165804 75404 165856 75410
rect 165804 75346 165856 75352
rect 165712 75336 165764 75342
rect 165712 75278 165764 75284
rect 165620 67312 165672 67318
rect 165620 67254 165672 67260
rect 165436 67108 165488 67114
rect 165436 67050 165488 67056
rect 165068 64524 165120 64530
rect 165068 64466 165120 64472
rect 164424 62552 164476 62558
rect 164424 62494 164476 62500
rect 164240 56024 164292 56030
rect 164240 55966 164292 55972
rect 165448 29714 165476 67050
rect 165528 63300 165580 63306
rect 165528 63242 165580 63248
rect 165540 62558 165568 63242
rect 165620 63028 165672 63034
rect 165620 62970 165672 62976
rect 165528 62552 165580 62558
rect 165528 62494 165580 62500
rect 165436 29708 165488 29714
rect 165436 29650 165488 29656
rect 164148 7608 164200 7614
rect 164148 7550 164200 7556
rect 165540 4826 165568 62494
rect 165528 4820 165580 4826
rect 165528 4762 165580 4768
rect 165632 3602 165660 62970
rect 165724 55214 165752 75278
rect 165816 62422 165844 75346
rect 165896 75268 165948 75274
rect 165896 75210 165948 75216
rect 165908 67454 165936 75210
rect 166000 67590 166028 79630
rect 166092 78441 166120 79750
rect 166494 79766 166546 79772
rect 166860 79826 166916 79835
rect 167058 79812 167086 80036
rect 167150 79971 167178 80036
rect 167136 79962 167192 79971
rect 167136 79897 167192 79906
rect 167242 79898 167270 80036
rect 167230 79892 167282 79898
rect 167230 79834 167282 79840
rect 166170 79727 166226 79736
rect 166264 79756 166316 79762
rect 166860 79761 166916 79770
rect 167012 79784 167086 79812
rect 166184 78470 166212 79727
rect 166264 79698 166316 79704
rect 166172 78464 166224 78470
rect 166078 78432 166134 78441
rect 166172 78406 166224 78412
rect 166078 78367 166134 78376
rect 166172 77240 166224 77246
rect 166172 77182 166224 77188
rect 166184 74089 166212 77182
rect 166276 75410 166304 79698
rect 166540 79688 166592 79694
rect 166540 79630 166592 79636
rect 166448 79620 166500 79626
rect 166448 79562 166500 79568
rect 166356 79552 166408 79558
rect 166356 79494 166408 79500
rect 166264 75404 166316 75410
rect 166264 75346 166316 75352
rect 166170 74080 166226 74089
rect 166170 74015 166226 74024
rect 166368 73930 166396 79494
rect 166460 75274 166488 79562
rect 166552 75342 166580 79630
rect 166724 79620 166776 79626
rect 166644 79580 166724 79608
rect 166644 77790 166672 79580
rect 166724 79562 166776 79568
rect 166816 79620 166868 79626
rect 166816 79562 166868 79568
rect 166722 79520 166778 79529
rect 166722 79455 166778 79464
rect 166632 77784 166684 77790
rect 166632 77726 166684 77732
rect 166736 77722 166764 79455
rect 166828 78849 166856 79562
rect 166814 78840 166870 78849
rect 166814 78775 166870 78784
rect 166816 77920 166868 77926
rect 166816 77862 166868 77868
rect 166724 77716 166776 77722
rect 166724 77658 166776 77664
rect 166540 75336 166592 75342
rect 166540 75278 166592 75284
rect 166448 75268 166500 75274
rect 166448 75210 166500 75216
rect 166092 73902 166396 73930
rect 166092 70258 166120 73902
rect 166170 73808 166226 73817
rect 166170 73743 166226 73752
rect 166184 70378 166212 73743
rect 166828 70394 166856 77862
rect 167012 77294 167040 79784
rect 167334 79778 167362 80036
rect 167288 79750 167362 79778
rect 167288 79422 167316 79750
rect 167426 79744 167454 80036
rect 167518 79966 167546 80036
rect 167610 79966 167638 80036
rect 167506 79960 167558 79966
rect 167506 79902 167558 79908
rect 167598 79960 167650 79966
rect 167598 79902 167650 79908
rect 167702 79778 167730 80036
rect 167656 79750 167730 79778
rect 167426 79716 167500 79744
rect 167184 79416 167236 79422
rect 167184 79358 167236 79364
rect 167276 79416 167328 79422
rect 167276 79358 167328 79364
rect 167196 79286 167224 79358
rect 167184 79280 167236 79286
rect 167184 79222 167236 79228
rect 167012 77266 167132 77294
rect 167104 76922 167132 77266
rect 167288 77042 167316 79358
rect 167276 77036 167328 77042
rect 167276 76978 167328 76984
rect 167104 76894 167408 76922
rect 167092 75812 167144 75818
rect 167092 75754 167144 75760
rect 167000 75336 167052 75342
rect 167000 75278 167052 75284
rect 166172 70372 166224 70378
rect 166172 70314 166224 70320
rect 166644 70366 166856 70394
rect 166092 70230 166212 70258
rect 166184 69698 166212 70230
rect 166172 69692 166224 69698
rect 166172 69634 166224 69640
rect 165988 67584 166040 67590
rect 165988 67526 166040 67532
rect 165896 67448 165948 67454
rect 165896 67390 165948 67396
rect 166184 67046 166212 69634
rect 166644 69018 166672 70366
rect 166632 69012 166684 69018
rect 166632 68954 166684 68960
rect 166816 67584 166868 67590
rect 166816 67526 166868 67532
rect 166172 67040 166224 67046
rect 166172 66982 166224 66988
rect 166828 66842 166856 67526
rect 166908 67448 166960 67454
rect 166908 67390 166960 67396
rect 166920 67182 166948 67390
rect 166908 67176 166960 67182
rect 166908 67118 166960 67124
rect 166816 66836 166868 66842
rect 166816 66778 166868 66784
rect 166724 62620 166776 62626
rect 166724 62562 166776 62568
rect 166736 62422 166764 62562
rect 165804 62416 165856 62422
rect 165804 62358 165856 62364
rect 166724 62416 166776 62422
rect 166724 62358 166776 62364
rect 165712 55208 165764 55214
rect 165712 55150 165764 55156
rect 166736 31074 166764 62358
rect 166724 31068 166776 31074
rect 166724 31010 166776 31016
rect 166828 26994 166856 66778
rect 166816 26988 166868 26994
rect 166816 26930 166868 26936
rect 166920 21418 166948 67118
rect 167012 51066 167040 75278
rect 167104 75206 167132 75754
rect 167184 75268 167236 75274
rect 167184 75210 167236 75216
rect 167092 75200 167144 75206
rect 167092 75142 167144 75148
rect 167092 70168 167144 70174
rect 167092 70110 167144 70116
rect 167104 69766 167132 70110
rect 167092 69760 167144 69766
rect 167092 69702 167144 69708
rect 167196 64874 167224 75210
rect 167276 75200 167328 75206
rect 167276 75142 167328 75148
rect 167288 65686 167316 75142
rect 167380 68882 167408 76894
rect 167472 70174 167500 79716
rect 167550 79656 167606 79665
rect 167550 79591 167606 79600
rect 167564 78538 167592 79591
rect 167552 78532 167604 78538
rect 167552 78474 167604 78480
rect 167552 78056 167604 78062
rect 167552 77998 167604 78004
rect 167564 70394 167592 77998
rect 167656 75154 167684 79750
rect 167794 79676 167822 80036
rect 167748 79648 167822 79676
rect 167886 79676 167914 80036
rect 167978 79744 168006 80036
rect 168070 79971 168098 80036
rect 168056 79962 168112 79971
rect 168056 79897 168112 79906
rect 168162 79778 168190 80036
rect 168254 79903 168282 80036
rect 168240 79894 168296 79903
rect 168240 79829 168296 79838
rect 168346 79778 168374 80036
rect 168438 79830 168466 80036
rect 168530 79830 168558 80036
rect 168116 79750 168190 79778
rect 168300 79750 168374 79778
rect 168426 79824 168478 79830
rect 168426 79766 168478 79772
rect 168518 79824 168570 79830
rect 168622 79801 168650 80036
rect 168518 79766 168570 79772
rect 168608 79792 168664 79801
rect 167978 79716 168052 79744
rect 167886 79648 167960 79676
rect 167748 75274 167776 79648
rect 167828 79552 167880 79558
rect 167828 79494 167880 79500
rect 167840 76650 167868 79494
rect 167932 76945 167960 79648
rect 168024 78985 168052 79716
rect 168010 78976 168066 78985
rect 168010 78911 168066 78920
rect 167918 76936 167974 76945
rect 167918 76871 167974 76880
rect 167840 76622 167960 76650
rect 167736 75268 167788 75274
rect 167736 75210 167788 75216
rect 167656 75126 167868 75154
rect 167840 70394 167868 75126
rect 167932 72826 167960 76622
rect 168116 75206 168144 79750
rect 168194 79656 168250 79665
rect 168194 79591 168250 79600
rect 168208 75206 168236 79591
rect 168300 75342 168328 79750
rect 168714 79778 168742 80036
rect 168806 79898 168834 80036
rect 168794 79892 168846 79898
rect 168794 79834 168846 79840
rect 168714 79750 168834 79778
rect 168608 79727 168664 79736
rect 168656 79688 168708 79694
rect 168378 79656 168434 79665
rect 168806 79676 168834 79750
rect 168898 79744 168926 80036
rect 168990 79898 169018 80036
rect 168978 79892 169030 79898
rect 168978 79834 169030 79840
rect 169082 79778 169110 80036
rect 169174 79966 169202 80036
rect 169162 79960 169214 79966
rect 169162 79902 169214 79908
rect 169266 79812 169294 80036
rect 169220 79784 169294 79812
rect 169082 79750 169156 79778
rect 168898 79716 168972 79744
rect 168806 79648 168880 79676
rect 168656 79630 168708 79636
rect 168378 79591 168434 79600
rect 168288 75336 168340 75342
rect 168288 75278 168340 75284
rect 168104 75200 168156 75206
rect 168104 75142 168156 75148
rect 168196 75200 168248 75206
rect 168196 75142 168248 75148
rect 167920 72820 167972 72826
rect 167920 72762 167972 72768
rect 167564 70366 167776 70394
rect 167840 70366 168328 70394
rect 167460 70168 167512 70174
rect 167460 70110 167512 70116
rect 167368 68876 167420 68882
rect 167368 68818 167420 68824
rect 167748 67590 167776 70366
rect 167736 67584 167788 67590
rect 167736 67526 167788 67532
rect 167276 65680 167328 65686
rect 167276 65622 167328 65628
rect 167104 64846 167224 64874
rect 167104 53786 167132 64846
rect 168300 63102 168328 70366
rect 168288 63096 168340 63102
rect 168288 63038 168340 63044
rect 167092 53780 167144 53786
rect 167092 53722 167144 53728
rect 167000 51060 167052 51066
rect 167000 51002 167052 51008
rect 168300 35222 168328 63038
rect 168392 46918 168420 79591
rect 168564 79552 168616 79558
rect 168564 79494 168616 79500
rect 168472 79484 168524 79490
rect 168472 79426 168524 79432
rect 168484 77178 168512 79426
rect 168472 77172 168524 77178
rect 168472 77114 168524 77120
rect 168484 76770 168512 77114
rect 168472 76764 168524 76770
rect 168472 76706 168524 76712
rect 168472 75268 168524 75274
rect 168472 75210 168524 75216
rect 168484 62082 168512 75210
rect 168576 62830 168604 79494
rect 168668 63442 168696 79630
rect 168748 79552 168800 79558
rect 168748 79494 168800 79500
rect 168760 64734 168788 79494
rect 168852 77382 168880 79648
rect 168944 78062 168972 79716
rect 169024 79688 169076 79694
rect 169024 79630 169076 79636
rect 169036 78402 169064 79630
rect 169024 78396 169076 78402
rect 169024 78338 169076 78344
rect 168932 78056 168984 78062
rect 168932 77998 168984 78004
rect 169128 77518 169156 79750
rect 169116 77512 169168 77518
rect 169116 77454 169168 77460
rect 168840 77376 168892 77382
rect 168840 77318 168892 77324
rect 169022 76800 169078 76809
rect 169022 76735 169078 76744
rect 169036 74186 169064 76735
rect 169220 75274 169248 79784
rect 169358 79744 169386 80036
rect 169450 79830 169478 80036
rect 169542 79971 169570 80036
rect 169528 79962 169584 79971
rect 169528 79897 169584 79906
rect 169634 79898 169662 80036
rect 169622 79892 169674 79898
rect 169622 79834 169674 79840
rect 169438 79824 169490 79830
rect 169438 79766 169490 79772
rect 169312 79716 169386 79744
rect 169208 75268 169260 75274
rect 169208 75210 169260 75216
rect 169024 74180 169076 74186
rect 169024 74122 169076 74128
rect 169312 70394 169340 79716
rect 169726 79676 169754 80036
rect 169818 79778 169846 80036
rect 169910 79937 169938 80036
rect 169896 79928 169952 79937
rect 170002 79898 170030 80036
rect 170094 79898 170122 80036
rect 170186 79937 170214 80036
rect 170172 79928 170228 79937
rect 169896 79863 169952 79872
rect 169990 79892 170042 79898
rect 169990 79834 170042 79840
rect 170082 79892 170134 79898
rect 170172 79863 170228 79872
rect 170082 79834 170134 79840
rect 169818 79750 169892 79778
rect 169726 79648 169800 79676
rect 169484 79552 169536 79558
rect 169484 79494 169536 79500
rect 169496 78690 169524 79494
rect 169772 79121 169800 79648
rect 169758 79112 169814 79121
rect 169758 79047 169814 79056
rect 169404 78662 169524 78690
rect 169404 76809 169432 78662
rect 169484 78600 169536 78606
rect 169484 78542 169536 78548
rect 169390 76800 169446 76809
rect 169390 76735 169446 76744
rect 169496 74526 169524 78542
rect 169576 78532 169628 78538
rect 169576 78474 169628 78480
rect 169484 74520 169536 74526
rect 169484 74462 169536 74468
rect 169220 70366 169340 70394
rect 169220 67250 169248 70366
rect 168840 67244 168892 67250
rect 168840 67186 168892 67192
rect 169208 67244 169260 67250
rect 169208 67186 169260 67192
rect 168852 66638 168880 67186
rect 168840 66632 168892 66638
rect 168840 66574 168892 66580
rect 168748 64728 168800 64734
rect 168748 64670 168800 64676
rect 168656 63436 168708 63442
rect 168656 63378 168708 63384
rect 169588 63238 169616 78474
rect 169668 77988 169720 77994
rect 169668 77930 169720 77936
rect 169680 75857 169708 77930
rect 169758 75984 169814 75993
rect 169758 75919 169814 75928
rect 169666 75848 169722 75857
rect 169666 75783 169722 75792
rect 169772 65958 169800 75919
rect 169760 65952 169812 65958
rect 169760 65894 169812 65900
rect 169576 63232 169628 63238
rect 169576 63174 169628 63180
rect 168564 62824 168616 62830
rect 168564 62766 168616 62772
rect 168472 62076 168524 62082
rect 168472 62018 168524 62024
rect 169760 49700 169812 49706
rect 169760 49642 169812 49648
rect 168380 46912 168432 46918
rect 168380 46854 168432 46860
rect 168288 35216 168340 35222
rect 168288 35158 168340 35164
rect 166908 21412 166960 21418
rect 166908 21354 166960 21360
rect 169772 16574 169800 49642
rect 169864 48210 169892 79750
rect 169944 79756 169996 79762
rect 169944 79698 169996 79704
rect 170036 79756 170088 79762
rect 170036 79698 170088 79704
rect 169956 67454 169984 79698
rect 170048 74866 170076 79698
rect 170278 79676 170306 80036
rect 170232 79648 170306 79676
rect 170232 75410 170260 79648
rect 170370 79608 170398 80036
rect 170462 79676 170490 80036
rect 170554 79744 170582 80036
rect 170646 79812 170674 80036
rect 170738 79966 170766 80036
rect 170830 79971 170858 80036
rect 170726 79960 170778 79966
rect 170726 79902 170778 79908
rect 170816 79962 170872 79971
rect 170816 79897 170872 79906
rect 170646 79784 170720 79812
rect 170554 79716 170628 79744
rect 170462 79648 170536 79676
rect 170324 79580 170398 79608
rect 170220 75404 170272 75410
rect 170220 75346 170272 75352
rect 170036 74860 170088 74866
rect 170036 74802 170088 74808
rect 170324 70394 170352 79580
rect 170404 79484 170456 79490
rect 170404 79426 170456 79432
rect 170416 78606 170444 79426
rect 170508 79082 170536 79648
rect 170496 79076 170548 79082
rect 170496 79018 170548 79024
rect 170600 78674 170628 79716
rect 170588 78668 170640 78674
rect 170588 78610 170640 78616
rect 170404 78600 170456 78606
rect 170404 78542 170456 78548
rect 170588 78532 170640 78538
rect 170588 78474 170640 78480
rect 170600 75070 170628 78474
rect 170692 78441 170720 79784
rect 170922 79778 170950 80036
rect 171014 79801 171042 80036
rect 170876 79750 170950 79778
rect 171000 79792 171056 79801
rect 170678 78432 170734 78441
rect 170678 78367 170734 78376
rect 170876 78305 170904 79750
rect 171000 79727 171056 79736
rect 171106 79676 171134 80036
rect 171060 79648 171134 79676
rect 170956 79552 171008 79558
rect 170956 79494 171008 79500
rect 170862 78296 170918 78305
rect 170862 78231 170918 78240
rect 170968 78033 170996 79494
rect 171060 78538 171088 79648
rect 171198 79608 171226 80036
rect 171290 79744 171318 80036
rect 171382 79898 171410 80036
rect 171370 79892 171422 79898
rect 171370 79834 171422 79840
rect 171474 79778 171502 80036
rect 171566 79830 171594 80036
rect 171658 79971 171686 80036
rect 171644 79962 171700 79971
rect 171644 79897 171700 79906
rect 171750 79898 171778 80036
rect 171842 79898 171870 80036
rect 171738 79892 171790 79898
rect 171738 79834 171790 79840
rect 171830 79892 171882 79898
rect 171830 79834 171882 79840
rect 171428 79750 171502 79778
rect 171554 79824 171606 79830
rect 171554 79766 171606 79772
rect 171290 79716 171364 79744
rect 171152 79580 171226 79608
rect 171048 78532 171100 78538
rect 171048 78474 171100 78480
rect 170954 78024 171010 78033
rect 170954 77959 171010 77968
rect 170680 77512 170732 77518
rect 170680 77454 170732 77460
rect 170588 75064 170640 75070
rect 170588 75006 170640 75012
rect 170232 70366 170352 70394
rect 170232 70281 170260 70366
rect 170218 70272 170274 70281
rect 170218 70207 170274 70216
rect 169944 67448 169996 67454
rect 169944 67390 169996 67396
rect 170692 62694 170720 77454
rect 170864 75948 170916 75954
rect 170864 75890 170916 75896
rect 170876 72593 170904 75890
rect 171048 75744 171100 75750
rect 171048 75686 171100 75692
rect 171060 73098 171088 75686
rect 171048 73092 171100 73098
rect 171048 73034 171100 73040
rect 170862 72584 170918 72593
rect 170862 72519 170918 72528
rect 171048 65952 171100 65958
rect 171048 65894 171100 65900
rect 170680 62688 170732 62694
rect 170680 62630 170732 62636
rect 169852 48204 169904 48210
rect 169852 48146 169904 48152
rect 171060 22778 171088 65894
rect 171152 46850 171180 79580
rect 171232 78736 171284 78742
rect 171232 78678 171284 78684
rect 171244 65482 171272 78678
rect 171336 78470 171364 79716
rect 171324 78464 171376 78470
rect 171324 78406 171376 78412
rect 171324 76424 171376 76430
rect 171324 76366 171376 76372
rect 171336 65890 171364 76366
rect 171428 70009 171456 79750
rect 171508 79688 171560 79694
rect 171692 79688 171744 79694
rect 171508 79630 171560 79636
rect 171598 79656 171654 79665
rect 171520 78742 171548 79630
rect 171692 79630 171744 79636
rect 171784 79688 171836 79694
rect 171934 79676 171962 80036
rect 172026 79801 172054 80036
rect 172118 79812 172146 80036
rect 172210 79966 172238 80036
rect 172198 79960 172250 79966
rect 172198 79902 172250 79908
rect 172302 79898 172330 80036
rect 172394 79898 172422 80036
rect 172486 79971 172514 80036
rect 172472 79962 172528 79971
rect 172578 79966 172606 80036
rect 172290 79892 172342 79898
rect 172290 79834 172342 79840
rect 172382 79892 172434 79898
rect 172472 79897 172528 79906
rect 172566 79960 172618 79966
rect 172670 79937 172698 80036
rect 172566 79902 172618 79908
rect 172656 79928 172712 79937
rect 172762 79898 172790 80036
rect 172854 79966 172882 80036
rect 172946 79966 172974 80036
rect 172842 79960 172894 79966
rect 172842 79902 172894 79908
rect 172934 79960 172986 79966
rect 172934 79902 172986 79908
rect 172656 79863 172712 79872
rect 172750 79892 172802 79898
rect 172382 79834 172434 79840
rect 172750 79834 172802 79840
rect 172566 79824 172618 79830
rect 172012 79792 172068 79801
rect 172118 79784 172192 79812
rect 172164 79778 172192 79784
rect 172618 79792 172666 79801
rect 172164 79750 172284 79778
rect 172566 79766 172610 79772
rect 172578 79750 172610 79766
rect 172012 79727 172068 79736
rect 171934 79648 172008 79676
rect 171784 79630 171836 79636
rect 171598 79591 171654 79600
rect 171508 78736 171560 78742
rect 171508 78678 171560 78684
rect 171508 78600 171560 78606
rect 171508 78542 171560 78548
rect 171520 71194 171548 78542
rect 171612 77858 171640 79591
rect 171600 77852 171652 77858
rect 171600 77794 171652 77800
rect 171704 75342 171732 79630
rect 171796 76430 171824 79630
rect 171876 79552 171928 79558
rect 171876 79494 171928 79500
rect 171888 78985 171916 79494
rect 171980 79286 172008 79648
rect 172060 79484 172112 79490
rect 172060 79426 172112 79432
rect 171968 79280 172020 79286
rect 171968 79222 172020 79228
rect 171874 78976 171930 78985
rect 171874 78911 171930 78920
rect 171876 77784 171928 77790
rect 171876 77726 171928 77732
rect 171784 76424 171836 76430
rect 171784 76366 171836 76372
rect 171692 75336 171744 75342
rect 171692 75278 171744 75284
rect 171888 73166 171916 77726
rect 171968 75336 172020 75342
rect 171968 75278 172020 75284
rect 171876 73160 171928 73166
rect 171876 73102 171928 73108
rect 171980 71233 172008 75278
rect 172072 74390 172100 79426
rect 172256 78742 172284 79750
rect 172610 79727 172666 79736
rect 173038 79744 173066 80036
rect 173130 79937 173158 80036
rect 173116 79928 173172 79937
rect 173116 79863 173172 79872
rect 173222 79744 173250 80036
rect 173314 79898 173342 80036
rect 173406 79898 173434 80036
rect 173498 79966 173526 80036
rect 173590 79966 173618 80036
rect 173682 79966 173710 80036
rect 173774 79971 173802 80036
rect 173486 79960 173538 79966
rect 173486 79902 173538 79908
rect 173578 79960 173630 79966
rect 173578 79902 173630 79908
rect 173670 79960 173722 79966
rect 173670 79902 173722 79908
rect 173760 79962 173816 79971
rect 173866 79966 173894 80036
rect 173958 79971 173986 80036
rect 173302 79892 173354 79898
rect 173302 79834 173354 79840
rect 173394 79892 173446 79898
rect 173760 79897 173816 79906
rect 173854 79960 173906 79966
rect 173854 79902 173906 79908
rect 173944 79962 174000 79971
rect 174050 79966 174078 80036
rect 173944 79897 174000 79906
rect 174038 79960 174090 79966
rect 174038 79902 174090 79908
rect 173394 79834 173446 79840
rect 174038 79824 174090 79830
rect 174036 79792 174038 79801
rect 174142 79812 174170 80036
rect 174234 79966 174262 80036
rect 174326 79966 174354 80036
rect 174222 79960 174274 79966
rect 174222 79902 174274 79908
rect 174314 79960 174366 79966
rect 174314 79902 174366 79908
rect 174268 79824 174320 79830
rect 174090 79792 174092 79801
rect 174142 79784 174216 79812
rect 173038 79716 173112 79744
rect 172796 79688 172848 79694
rect 172796 79630 172848 79636
rect 172704 79620 172756 79626
rect 172704 79562 172756 79568
rect 172520 79552 172572 79558
rect 172520 79494 172572 79500
rect 172336 79484 172388 79490
rect 172336 79426 172388 79432
rect 172244 78736 172296 78742
rect 172244 78678 172296 78684
rect 172348 77294 172376 79426
rect 172532 78606 172560 79494
rect 172520 78600 172572 78606
rect 172426 78568 172482 78577
rect 172520 78542 172572 78548
rect 172610 78568 172666 78577
rect 172426 78503 172482 78512
rect 172610 78503 172666 78512
rect 172256 77266 172376 77294
rect 172152 74860 172204 74866
rect 172152 74802 172204 74808
rect 172060 74384 172112 74390
rect 172060 74326 172112 74332
rect 172164 71330 172192 74802
rect 172256 71670 172284 77266
rect 172440 76537 172468 78503
rect 172426 76528 172482 76537
rect 172426 76463 172482 76472
rect 172520 75948 172572 75954
rect 172520 75890 172572 75896
rect 172244 71664 172296 71670
rect 172244 71606 172296 71612
rect 172152 71324 172204 71330
rect 172152 71266 172204 71272
rect 171966 71224 172022 71233
rect 171508 71188 171560 71194
rect 171966 71159 172022 71168
rect 171508 71130 171560 71136
rect 171414 70000 171470 70009
rect 172532 69970 172560 75890
rect 171414 69935 171470 69944
rect 172520 69964 172572 69970
rect 172520 69906 172572 69912
rect 172624 69902 172652 78503
rect 172716 71534 172744 79562
rect 172808 78062 172836 79630
rect 172980 79620 173032 79626
rect 172980 79562 173032 79568
rect 172796 78056 172848 78062
rect 172796 77998 172848 78004
rect 172992 75954 173020 79562
rect 172980 75948 173032 75954
rect 172980 75890 173032 75896
rect 173084 75002 173112 79716
rect 173176 79716 173250 79744
rect 173716 79756 173768 79762
rect 173176 79665 173204 79716
rect 173716 79698 173768 79704
rect 173900 79756 173952 79762
rect 174036 79727 174092 79736
rect 173900 79698 173952 79704
rect 173348 79688 173400 79694
rect 173162 79656 173218 79665
rect 173348 79630 173400 79636
rect 173440 79688 173492 79694
rect 173440 79630 173492 79636
rect 173162 79591 173218 79600
rect 173256 79620 173308 79626
rect 173256 79562 173308 79568
rect 173164 79552 173216 79558
rect 173164 79494 173216 79500
rect 173176 77654 173204 79494
rect 173268 78441 173296 79562
rect 173254 78432 173310 78441
rect 173254 78367 173310 78376
rect 173164 77648 173216 77654
rect 173164 77590 173216 77596
rect 173360 77042 173388 79630
rect 173348 77036 173400 77042
rect 173348 76978 173400 76984
rect 173072 74996 173124 75002
rect 173072 74938 173124 74944
rect 173452 74050 173480 79630
rect 173624 79620 173676 79626
rect 173624 79562 173676 79568
rect 173636 78690 173664 79562
rect 173544 78662 173664 78690
rect 173440 74044 173492 74050
rect 173440 73986 173492 73992
rect 172704 71528 172756 71534
rect 172704 71470 172756 71476
rect 173544 70394 173572 78662
rect 173624 78600 173676 78606
rect 173624 78542 173676 78548
rect 172716 70366 173572 70394
rect 172612 69896 172664 69902
rect 172612 69838 172664 69844
rect 172716 69766 172744 70366
rect 173636 70145 173664 78542
rect 173728 78130 173756 79698
rect 173806 79656 173862 79665
rect 173806 79591 173862 79600
rect 173912 79608 173940 79698
rect 173716 78124 173768 78130
rect 173716 78066 173768 78072
rect 173714 77888 173770 77897
rect 173714 77823 173770 77832
rect 173728 72622 173756 77823
rect 173820 77654 173848 79591
rect 173912 79580 174032 79608
rect 173900 79484 173952 79490
rect 173900 79426 173952 79432
rect 173912 78674 173940 79426
rect 173900 78668 173952 78674
rect 173900 78610 173952 78616
rect 173900 77716 173952 77722
rect 173900 77658 173952 77664
rect 173808 77648 173860 77654
rect 173808 77590 173860 77596
rect 173912 73030 173940 77658
rect 174004 76673 174032 79580
rect 174188 77926 174216 79784
rect 174418 79778 174446 80036
rect 174268 79766 174320 79772
rect 174280 79014 174308 79766
rect 174372 79750 174446 79778
rect 174510 79778 174538 80036
rect 174602 79966 174630 80036
rect 174590 79960 174642 79966
rect 174694 79937 174722 80036
rect 174786 79966 174814 80036
rect 174878 79966 174906 80036
rect 174774 79960 174826 79966
rect 174590 79902 174642 79908
rect 174680 79928 174736 79937
rect 174774 79902 174826 79908
rect 174866 79960 174918 79966
rect 174866 79902 174918 79908
rect 174680 79863 174736 79872
rect 174636 79824 174688 79830
rect 174510 79750 174584 79778
rect 174636 79766 174688 79772
rect 174728 79824 174780 79830
rect 174970 79778 174998 80036
rect 175062 79898 175090 80036
rect 175154 79966 175182 80036
rect 175246 79971 175274 80036
rect 175142 79960 175194 79966
rect 175142 79902 175194 79908
rect 175232 79962 175288 79971
rect 175050 79892 175102 79898
rect 175232 79897 175288 79906
rect 175050 79834 175102 79840
rect 174728 79766 174780 79772
rect 174268 79008 174320 79014
rect 174268 78950 174320 78956
rect 174176 77920 174228 77926
rect 174176 77862 174228 77868
rect 173990 76664 174046 76673
rect 173990 76599 174046 76608
rect 173992 75948 174044 75954
rect 173992 75890 174044 75896
rect 173900 73024 173952 73030
rect 173900 72966 173952 72972
rect 173716 72616 173768 72622
rect 173716 72558 173768 72564
rect 173622 70136 173678 70145
rect 173622 70071 173678 70080
rect 173164 69896 173216 69902
rect 173164 69838 173216 69844
rect 172704 69760 172756 69766
rect 172704 69702 172756 69708
rect 171324 65884 171376 65890
rect 171324 65826 171376 65832
rect 172336 65884 172388 65890
rect 172336 65826 172388 65832
rect 171232 65476 171284 65482
rect 171232 65418 171284 65424
rect 171140 46844 171192 46850
rect 171140 46786 171192 46792
rect 171048 22772 171100 22778
rect 171048 22714 171100 22720
rect 169772 16546 170720 16574
rect 165620 3596 165672 3602
rect 165620 3538 165672 3544
rect 166816 3596 166868 3602
rect 166816 3538 166868 3544
rect 166828 480 166856 3538
rect 170692 480 170720 16546
rect 172348 14550 172376 65826
rect 172428 65476 172480 65482
rect 172428 65418 172480 65424
rect 172440 65278 172468 65418
rect 172428 65272 172480 65278
rect 172428 65214 172480 65220
rect 172336 14544 172388 14550
rect 172336 14486 172388 14492
rect 172440 10402 172468 65214
rect 173176 49706 173204 69838
rect 174004 63646 174032 75890
rect 174268 75880 174320 75886
rect 174268 75822 174320 75828
rect 174280 70394 174308 75822
rect 174372 75818 174400 79750
rect 174452 77920 174504 77926
rect 174452 77862 174504 77868
rect 174360 75812 174412 75818
rect 174360 75754 174412 75760
rect 174464 75342 174492 77862
rect 174452 75336 174504 75342
rect 174452 75278 174504 75284
rect 174556 71774 174584 79750
rect 174648 77790 174676 79766
rect 174636 77784 174688 77790
rect 174636 77726 174688 77732
rect 174636 77376 174688 77382
rect 174636 77318 174688 77324
rect 174096 70366 174308 70394
rect 174464 71746 174584 71774
rect 174096 65890 174124 70366
rect 174084 65884 174136 65890
rect 174084 65826 174136 65832
rect 173992 63640 174044 63646
rect 173992 63582 174044 63588
rect 174464 60722 174492 71746
rect 174544 69556 174596 69562
rect 174544 69498 174596 69504
rect 174452 60716 174504 60722
rect 174452 60658 174504 60664
rect 174556 49706 174584 69498
rect 174648 68474 174676 77318
rect 174740 73982 174768 79766
rect 174832 79750 174998 79778
rect 174832 75954 174860 79750
rect 175338 79744 175366 80036
rect 175292 79716 175366 79744
rect 175188 79688 175240 79694
rect 175002 79656 175058 79665
rect 175188 79630 175240 79636
rect 175002 79591 175058 79600
rect 175096 79620 175148 79626
rect 175016 76362 175044 79591
rect 175096 79562 175148 79568
rect 175004 76356 175056 76362
rect 175004 76298 175056 76304
rect 174820 75948 174872 75954
rect 174820 75890 174872 75896
rect 175108 75886 175136 79562
rect 175096 75880 175148 75886
rect 175096 75822 175148 75828
rect 174728 73976 174780 73982
rect 174728 73918 174780 73924
rect 175200 71602 175228 79630
rect 175292 78985 175320 79716
rect 175430 79676 175458 80036
rect 175522 79744 175550 80036
rect 175614 79966 175642 80036
rect 175602 79960 175654 79966
rect 175602 79902 175654 79908
rect 175706 79898 175734 80036
rect 175798 79966 175826 80036
rect 175786 79960 175838 79966
rect 175786 79902 175838 79908
rect 175694 79892 175746 79898
rect 175694 79834 175746 79840
rect 175648 79756 175700 79762
rect 175522 79716 175596 79744
rect 175430 79648 175504 79676
rect 175278 78976 175334 78985
rect 175278 78911 175334 78920
rect 175476 78266 175504 79648
rect 175464 78260 175516 78266
rect 175464 78202 175516 78208
rect 175372 75540 175424 75546
rect 175372 75482 175424 75488
rect 175280 75268 175332 75274
rect 175280 75210 175332 75216
rect 175188 71596 175240 71602
rect 175188 71538 175240 71544
rect 174636 68468 174688 68474
rect 174636 68410 174688 68416
rect 175292 65890 175320 75210
rect 175384 67046 175412 75482
rect 175476 72486 175504 78202
rect 175568 77897 175596 79716
rect 175890 79744 175918 80036
rect 175982 79937 176010 80036
rect 176074 79966 176102 80036
rect 176062 79960 176114 79966
rect 175968 79928 176024 79937
rect 176062 79902 176114 79908
rect 176166 79898 176194 80036
rect 175968 79863 176024 79872
rect 176154 79892 176206 79898
rect 176154 79834 176206 79840
rect 176016 79824 176068 79830
rect 176258 79778 176286 80036
rect 176350 79966 176378 80036
rect 176338 79960 176390 79966
rect 176338 79902 176390 79908
rect 176442 79830 176470 80036
rect 176534 79966 176562 80036
rect 176626 79971 176654 80036
rect 176522 79960 176574 79966
rect 176522 79902 176574 79908
rect 176612 79962 176668 79971
rect 176612 79897 176668 79906
rect 176016 79766 176068 79772
rect 175648 79698 175700 79704
rect 175752 79716 175918 79744
rect 175660 79150 175688 79698
rect 175648 79144 175700 79150
rect 175648 79086 175700 79092
rect 175554 77888 175610 77897
rect 175554 77823 175610 77832
rect 175464 72480 175516 72486
rect 175464 72422 175516 72428
rect 175660 70394 175688 79086
rect 175752 78810 175780 79716
rect 175832 79620 175884 79626
rect 175832 79562 175884 79568
rect 175740 78804 175792 78810
rect 175740 78746 175792 78752
rect 175844 75750 175872 79562
rect 175922 78568 175978 78577
rect 175922 78503 175978 78512
rect 175832 75744 175884 75750
rect 175832 75686 175884 75692
rect 175936 75546 175964 78503
rect 176028 76265 176056 79766
rect 176108 79756 176160 79762
rect 176108 79698 176160 79704
rect 176212 79750 176286 79778
rect 176430 79824 176482 79830
rect 176430 79766 176482 79772
rect 176718 79778 176746 80036
rect 176810 79898 176838 80036
rect 176902 79971 176930 80036
rect 176888 79962 176944 79971
rect 176994 79966 177022 80036
rect 176798 79892 176850 79898
rect 176888 79897 176944 79906
rect 176982 79960 177034 79966
rect 176982 79902 177034 79908
rect 176798 79834 176850 79840
rect 176936 79824 176988 79830
rect 176718 79750 176792 79778
rect 177086 79812 177114 80036
rect 177178 79966 177206 80036
rect 177166 79960 177218 79966
rect 177166 79902 177218 79908
rect 177270 79898 177298 80036
rect 177362 79898 177390 80036
rect 177454 79937 177482 80036
rect 177546 79948 177574 80036
rect 177946 79999 177948 80008
rect 178000 79999 178002 80008
rect 177948 79970 178000 79976
rect 177440 79928 177496 79937
rect 177258 79892 177310 79898
rect 177258 79834 177310 79840
rect 177350 79892 177402 79898
rect 177546 79920 177620 79948
rect 177440 79863 177496 79872
rect 177350 79834 177402 79840
rect 177086 79784 177160 79812
rect 176936 79766 176988 79772
rect 177132 79778 177160 79784
rect 176014 76256 176070 76265
rect 176014 76191 176070 76200
rect 175924 75540 175976 75546
rect 175924 75482 175976 75488
rect 175832 75472 175884 75478
rect 175832 75414 175884 75420
rect 175568 70366 175688 70394
rect 175568 70242 175596 70366
rect 175556 70236 175608 70242
rect 175556 70178 175608 70184
rect 175372 67040 175424 67046
rect 175372 66982 175424 66988
rect 175096 65884 175148 65890
rect 175096 65826 175148 65832
rect 175280 65884 175332 65890
rect 175280 65826 175332 65832
rect 175108 65482 175136 65826
rect 175096 65476 175148 65482
rect 175096 65418 175148 65424
rect 173164 49700 173216 49706
rect 173164 49642 173216 49648
rect 174544 49700 174596 49706
rect 174544 49642 174596 49648
rect 175108 18630 175136 65418
rect 175844 64874 175872 75414
rect 176120 71262 176148 79698
rect 176212 75274 176240 79750
rect 176292 79688 176344 79694
rect 176292 79630 176344 79636
rect 176200 75268 176252 75274
rect 176200 75210 176252 75216
rect 176108 71256 176160 71262
rect 176108 71198 176160 71204
rect 176304 71058 176332 79630
rect 176568 79620 176620 79626
rect 176568 79562 176620 79568
rect 176474 78568 176530 78577
rect 176474 78503 176530 78512
rect 176488 75478 176516 78503
rect 176476 75472 176528 75478
rect 176476 75414 176528 75420
rect 176580 75041 176608 79562
rect 176566 75032 176622 75041
rect 176566 74967 176622 74976
rect 176764 71398 176792 79750
rect 176948 71466 176976 79766
rect 177132 79750 177206 79778
rect 177178 79676 177206 79750
rect 177304 79756 177356 79762
rect 177304 79698 177356 79704
rect 177178 79648 177252 79676
rect 177224 78402 177252 79648
rect 177212 78396 177264 78402
rect 177212 78338 177264 78344
rect 177316 77178 177344 79698
rect 177592 78674 177620 79920
rect 177672 79824 177724 79830
rect 177672 79766 177724 79772
rect 177580 78668 177632 78674
rect 177580 78610 177632 78616
rect 177684 77246 177712 79766
rect 178052 78606 178080 80106
rect 178144 80034 178172 80106
rect 178132 80028 178184 80034
rect 178132 79970 178184 79976
rect 178040 78600 178092 78606
rect 178040 78542 178092 78548
rect 177856 77988 177908 77994
rect 177856 77930 177908 77936
rect 177672 77240 177724 77246
rect 177672 77182 177724 77188
rect 177304 77172 177356 77178
rect 177304 77114 177356 77120
rect 177868 74254 177896 77930
rect 177948 75200 178000 75206
rect 177948 75142 178000 75148
rect 177856 74248 177908 74254
rect 177856 74190 177908 74196
rect 177960 72690 177988 75142
rect 178328 74225 178356 80242
rect 178420 80238 178448 80650
rect 178592 80640 178644 80646
rect 178592 80582 178644 80588
rect 187700 80640 187752 80646
rect 187700 80582 187752 80588
rect 178604 80481 178632 80582
rect 184204 80504 184256 80510
rect 178590 80472 178646 80481
rect 184204 80446 184256 80452
rect 187054 80472 187110 80481
rect 178590 80407 178646 80416
rect 178408 80232 178460 80238
rect 178408 80174 178460 80180
rect 181168 80164 181220 80170
rect 181168 80106 181220 80112
rect 179604 80096 179656 80102
rect 179604 80038 179656 80044
rect 178500 79892 178552 79898
rect 178500 79834 178552 79840
rect 178512 76906 178540 79834
rect 179616 79150 179644 80038
rect 179604 79144 179656 79150
rect 179604 79086 179656 79092
rect 181180 78810 181208 80106
rect 181626 79928 181682 79937
rect 181626 79863 181682 79872
rect 182916 79892 182968 79898
rect 181534 79792 181590 79801
rect 181534 79727 181590 79736
rect 181444 79620 181496 79626
rect 181444 79562 181496 79568
rect 181456 79218 181484 79562
rect 181548 79218 181576 79727
rect 181444 79212 181496 79218
rect 181444 79154 181496 79160
rect 181536 79212 181588 79218
rect 181536 79154 181588 79160
rect 180248 78804 180300 78810
rect 180248 78746 180300 78752
rect 181168 78804 181220 78810
rect 181168 78746 181220 78752
rect 179696 78124 179748 78130
rect 179696 78066 179748 78072
rect 178500 76900 178552 76906
rect 178500 76842 178552 76848
rect 179708 75546 179736 78066
rect 179696 75540 179748 75546
rect 179696 75482 179748 75488
rect 178314 74216 178370 74225
rect 178314 74151 178370 74160
rect 177948 72684 178000 72690
rect 177948 72626 178000 72632
rect 176936 71460 176988 71466
rect 176936 71402 176988 71408
rect 176752 71392 176804 71398
rect 176752 71334 176804 71340
rect 176016 71052 176068 71058
rect 176016 70994 176068 71000
rect 176292 71052 176344 71058
rect 176292 70994 176344 71000
rect 175844 64846 175964 64874
rect 175188 64660 175240 64666
rect 175188 64602 175240 64608
rect 175200 63646 175228 64602
rect 175188 63640 175240 63646
rect 175188 63582 175240 63588
rect 175096 18624 175148 18630
rect 175096 18566 175148 18572
rect 175200 13190 175228 63582
rect 175936 13258 175964 64846
rect 176028 55962 176056 70994
rect 180260 70990 180288 78746
rect 180616 78736 180668 78742
rect 180616 78678 180668 78684
rect 180340 77988 180392 77994
rect 180340 77930 180392 77936
rect 180352 76945 180380 77930
rect 180628 77081 180656 78678
rect 181640 78305 181668 79863
rect 182916 79834 182968 79840
rect 181626 78296 181682 78305
rect 181626 78231 181682 78240
rect 181720 78192 181772 78198
rect 181720 78134 181772 78140
rect 181536 78124 181588 78130
rect 181536 78066 181588 78072
rect 181260 78056 181312 78062
rect 180706 78024 180762 78033
rect 181260 77998 181312 78004
rect 180706 77959 180762 77968
rect 180720 77217 180748 77959
rect 180706 77208 180762 77217
rect 180706 77143 180762 77152
rect 180614 77072 180670 77081
rect 180614 77007 180670 77016
rect 180338 76936 180394 76945
rect 180338 76871 180394 76880
rect 181272 75614 181300 77998
rect 181352 77920 181404 77926
rect 181352 77862 181404 77868
rect 181260 75608 181312 75614
rect 181260 75550 181312 75556
rect 181364 74934 181392 77862
rect 181444 77852 181496 77858
rect 181444 77794 181496 77800
rect 181456 77217 181484 77794
rect 181442 77208 181498 77217
rect 181442 77143 181498 77152
rect 181352 74928 181404 74934
rect 181352 74870 181404 74876
rect 181548 74202 181576 78066
rect 181456 74174 181576 74202
rect 180248 70984 180300 70990
rect 180248 70926 180300 70932
rect 181456 68270 181484 74174
rect 181732 73930 181760 78134
rect 181812 78056 181864 78062
rect 181812 77998 181864 78004
rect 181548 73902 181760 73930
rect 181548 69426 181576 73902
rect 181824 70394 181852 77998
rect 182928 77897 182956 79834
rect 182914 77888 182970 77897
rect 182914 77823 182970 77832
rect 182916 76628 182968 76634
rect 182916 76570 182968 76576
rect 182088 75608 182140 75614
rect 182088 75550 182140 75556
rect 181640 70366 181852 70394
rect 181640 69494 181668 70366
rect 181628 69488 181680 69494
rect 181628 69430 181680 69436
rect 181536 69420 181588 69426
rect 181536 69362 181588 69368
rect 181444 68264 181496 68270
rect 181444 68206 181496 68212
rect 176568 65884 176620 65890
rect 176568 65826 176620 65832
rect 176660 65884 176712 65890
rect 176660 65826 176712 65832
rect 176580 65346 176608 65826
rect 176568 65340 176620 65346
rect 176568 65282 176620 65288
rect 176016 55956 176068 55962
rect 176016 55898 176068 55904
rect 176580 39370 176608 65282
rect 176672 65278 176700 65826
rect 176660 65272 176712 65278
rect 176660 65214 176712 65220
rect 176568 39364 176620 39370
rect 176568 39306 176620 39312
rect 182100 24818 182128 75550
rect 182824 73228 182876 73234
rect 182824 73170 182876 73176
rect 182180 68264 182232 68270
rect 182180 68206 182232 68212
rect 182088 24812 182140 24818
rect 182088 24754 182140 24760
rect 182192 16574 182220 68206
rect 182836 16590 182864 73170
rect 182928 52426 182956 76570
rect 184216 72214 184244 80446
rect 187054 80407 187110 80416
rect 184938 80200 184994 80209
rect 184938 80135 184994 80144
rect 184952 80034 184980 80135
rect 184940 80028 184992 80034
rect 184940 79970 184992 79976
rect 186962 79384 187018 79393
rect 186962 79319 187018 79328
rect 184940 73840 184992 73846
rect 184940 73782 184992 73788
rect 184952 72486 184980 73782
rect 184940 72480 184992 72486
rect 184940 72422 184992 72428
rect 186228 72480 186280 72486
rect 186228 72422 186280 72428
rect 184204 72208 184256 72214
rect 184204 72150 184256 72156
rect 184940 64320 184992 64326
rect 184940 64262 184992 64268
rect 184848 56024 184900 56030
rect 184848 55966 184900 55972
rect 184860 55146 184888 55966
rect 184848 55140 184900 55146
rect 184848 55082 184900 55088
rect 182916 52420 182968 52426
rect 182916 52362 182968 52368
rect 182824 16584 182876 16590
rect 182192 16546 182312 16574
rect 178408 15904 178460 15910
rect 178408 15846 178460 15852
rect 175924 13252 175976 13258
rect 175924 13194 175976 13200
rect 175188 13184 175240 13190
rect 175188 13126 175240 13132
rect 172428 10396 172480 10402
rect 172428 10338 172480 10344
rect 174544 3596 174596 3602
rect 174544 3538 174596 3544
rect 174556 480 174584 3538
rect 178420 480 178448 15846
rect 182284 480 182312 16546
rect 182824 16526 182876 16532
rect 184860 5506 184888 55082
rect 184952 16574 184980 64262
rect 186240 56574 186268 72422
rect 186976 67017 187004 79319
rect 187068 73137 187096 80407
rect 187712 79422 187740 80582
rect 188344 80572 188396 80578
rect 188344 80514 188396 80520
rect 187700 79416 187752 79422
rect 187700 79358 187752 79364
rect 187054 73128 187110 73137
rect 187054 73063 187110 73072
rect 186962 67008 187018 67017
rect 186962 66943 187018 66952
rect 188356 64598 188384 80514
rect 188632 65414 188660 182854
rect 188804 146328 188856 146334
rect 188804 146270 188856 146276
rect 188712 140480 188764 140486
rect 188712 140422 188764 140428
rect 188724 133793 188752 140422
rect 188710 133784 188766 133793
rect 188816 133770 188844 146270
rect 188908 143546 188936 198902
rect 189000 147014 189028 200126
rect 189080 197328 189132 197334
rect 189080 197270 189132 197276
rect 188988 147008 189040 147014
rect 188988 146950 189040 146956
rect 188896 143540 188948 143546
rect 188896 143482 188948 143488
rect 188988 142384 189040 142390
rect 188988 142326 189040 142332
rect 188896 141636 188948 141642
rect 188896 141578 188948 141584
rect 188908 133890 188936 141578
rect 189000 138718 189028 142326
rect 188988 138712 189040 138718
rect 188988 138654 189040 138660
rect 188896 133884 188948 133890
rect 188896 133826 188948 133832
rect 188816 133742 189028 133770
rect 188710 133719 188766 133728
rect 188896 133680 188948 133686
rect 188896 133622 188948 133628
rect 188908 133498 188936 133622
rect 188724 133470 188936 133498
rect 188620 65408 188672 65414
rect 188620 65350 188672 65356
rect 188344 64592 188396 64598
rect 188344 64534 188396 64540
rect 186228 56568 186280 56574
rect 186228 56510 186280 56516
rect 188724 51814 188752 133470
rect 189000 132546 189028 133742
rect 188816 132518 189028 132546
rect 188816 67386 188844 132518
rect 188894 104136 188950 104145
rect 188894 104071 188950 104080
rect 188804 67380 188856 67386
rect 188804 67322 188856 67328
rect 188908 64462 188936 104071
rect 189092 84930 189120 197270
rect 189356 193316 189408 193322
rect 189356 193258 189408 193264
rect 189172 190120 189224 190126
rect 189172 190062 189224 190068
rect 189184 86494 189212 190062
rect 189264 181348 189316 181354
rect 189264 181290 189316 181296
rect 189172 86488 189224 86494
rect 189172 86430 189224 86436
rect 189080 84924 189132 84930
rect 189080 84866 189132 84872
rect 188988 81116 189040 81122
rect 188988 81058 189040 81064
rect 189000 81002 189028 81058
rect 189000 80974 189120 81002
rect 188988 80912 189040 80918
rect 188988 80854 189040 80860
rect 189000 79558 189028 80854
rect 189092 80646 189120 80974
rect 189080 80640 189132 80646
rect 189080 80582 189132 80588
rect 189080 79688 189132 79694
rect 189080 79630 189132 79636
rect 188988 79552 189040 79558
rect 188988 79494 189040 79500
rect 189092 79370 189120 79630
rect 189000 79342 189120 79370
rect 189000 77761 189028 79342
rect 188986 77752 189042 77761
rect 188986 77687 189042 77696
rect 189000 74534 189028 77687
rect 189000 74506 189120 74534
rect 188988 70984 189040 70990
rect 188988 70926 189040 70932
rect 188896 64456 188948 64462
rect 188896 64398 188948 64404
rect 186228 51808 186280 51814
rect 186228 51750 186280 51756
rect 188712 51808 188764 51814
rect 188712 51750 188764 51756
rect 184952 16546 185072 16574
rect 184848 5500 184900 5506
rect 184848 5442 184900 5448
rect 132654 354 132766 480
rect 132512 326 132766 354
rect 132654 -960 132766 326
rect 136518 -960 136630 480
rect 140382 -960 140494 480
rect 144246 -960 144358 480
rect 147466 -960 147578 480
rect 151330 -960 151442 480
rect 155194 -960 155306 480
rect 159058 -960 159170 480
rect 162922 -960 163034 480
rect 166786 -960 166898 480
rect 170650 -960 170762 480
rect 174514 -960 174626 480
rect 178378 -960 178490 480
rect 182242 -960 182354 480
rect 185044 354 185072 16546
rect 186240 12442 186268 51750
rect 189000 28966 189028 70926
rect 188988 28960 189040 28966
rect 188988 28902 189040 28908
rect 186228 12436 186280 12442
rect 186228 12378 186280 12384
rect 185462 354 185574 480
rect 185044 326 185574 354
rect 189092 354 189120 74506
rect 189172 73908 189224 73914
rect 189172 73850 189224 73856
rect 189184 73710 189212 73850
rect 189172 73704 189224 73710
rect 189172 73646 189224 73652
rect 189276 66094 189304 181290
rect 189368 86630 189396 193258
rect 189460 193050 189488 700334
rect 189552 198490 189580 700538
rect 189724 700392 189776 700398
rect 189724 700334 189776 700340
rect 189632 259548 189684 259554
rect 189632 259490 189684 259496
rect 189540 198484 189592 198490
rect 189540 198426 189592 198432
rect 189552 194138 189580 198426
rect 189540 194132 189592 194138
rect 189540 194074 189592 194080
rect 189448 193044 189500 193050
rect 189448 192986 189500 192992
rect 189540 190596 189592 190602
rect 189540 190538 189592 190544
rect 189448 181824 189500 181830
rect 189448 181766 189500 181772
rect 189356 86624 189408 86630
rect 189356 86566 189408 86572
rect 189356 86488 189408 86494
rect 189356 86430 189408 86436
rect 189368 69601 189396 86430
rect 189354 69592 189410 69601
rect 189354 69527 189410 69536
rect 189460 68814 189488 181766
rect 189552 86766 189580 190538
rect 189644 142458 189672 259490
rect 189736 198762 189764 700334
rect 190656 699786 190684 703520
rect 191840 700528 191892 700534
rect 191840 700470 191892 700476
rect 190644 699780 190696 699786
rect 190644 699722 190696 699728
rect 189816 520328 189868 520334
rect 189816 520270 189868 520276
rect 189828 199073 189856 520270
rect 191748 400240 191800 400246
rect 191748 400182 191800 400188
rect 191104 364404 191156 364410
rect 191104 364346 191156 364352
rect 190552 266416 190604 266422
rect 190552 266358 190604 266364
rect 190460 265804 190512 265810
rect 190460 265746 190512 265752
rect 189906 263120 189962 263129
rect 189906 263055 189962 263064
rect 189920 262585 189948 263055
rect 189906 262576 189962 262585
rect 189906 262511 189962 262520
rect 189814 199064 189870 199073
rect 189814 198999 189870 199008
rect 189724 198756 189776 198762
rect 189724 198698 189776 198704
rect 189724 194064 189776 194070
rect 189724 194006 189776 194012
rect 189632 142452 189684 142458
rect 189632 142394 189684 142400
rect 189632 141704 189684 141710
rect 189632 141646 189684 141652
rect 189540 86760 189592 86766
rect 189540 86702 189592 86708
rect 189540 86624 189592 86630
rect 189540 86566 189592 86572
rect 189552 78606 189580 86566
rect 189540 78600 189592 78606
rect 189540 78542 189592 78548
rect 189448 68808 189500 68814
rect 189448 68750 189500 68756
rect 189264 66088 189316 66094
rect 189264 66030 189316 66036
rect 189644 38622 189672 141646
rect 189736 88398 189764 194006
rect 189920 145586 189948 262511
rect 189998 260128 190054 260137
rect 189998 260063 190054 260072
rect 190012 198257 190040 260063
rect 190092 244316 190144 244322
rect 190092 244258 190144 244264
rect 190104 198966 190132 244258
rect 190472 208962 190500 265746
rect 190460 208956 190512 208962
rect 190460 208898 190512 208904
rect 190460 200388 190512 200394
rect 190460 200330 190512 200336
rect 190472 199034 190500 200330
rect 190460 199028 190512 199034
rect 190460 198970 190512 198976
rect 190092 198960 190144 198966
rect 190092 198902 190144 198908
rect 189998 198248 190054 198257
rect 189998 198183 190054 198192
rect 190012 191146 190040 198183
rect 190000 191140 190052 191146
rect 190000 191082 190052 191088
rect 190460 179104 190512 179110
rect 190460 179046 190512 179052
rect 189908 145580 189960 145586
rect 189908 145522 189960 145528
rect 190000 142452 190052 142458
rect 190000 142394 190052 142400
rect 189816 140548 189868 140554
rect 189816 140490 189868 140496
rect 189724 88392 189776 88398
rect 189724 88334 189776 88340
rect 189724 84924 189776 84930
rect 189724 84866 189776 84872
rect 189736 78266 189764 84866
rect 189724 78260 189776 78266
rect 189724 78202 189776 78208
rect 189828 73914 189856 140490
rect 189908 139392 189960 139398
rect 189908 139334 189960 139340
rect 189920 138786 189948 139334
rect 189908 138780 189960 138786
rect 189908 138722 189960 138728
rect 190012 137290 190040 142394
rect 190000 137284 190052 137290
rect 190000 137226 190052 137232
rect 189908 88392 189960 88398
rect 189908 88334 189960 88340
rect 190090 88360 190146 88369
rect 189920 81433 189948 88334
rect 190090 88295 190146 88304
rect 189906 81424 189962 81433
rect 189906 81359 189962 81368
rect 190104 81138 190132 88295
rect 190184 86760 190236 86766
rect 190184 86702 190236 86708
rect 189920 81110 190132 81138
rect 189816 73908 189868 73914
rect 189816 73850 189868 73856
rect 189172 38616 189224 38622
rect 189172 38558 189224 38564
rect 189632 38616 189684 38622
rect 189632 38558 189684 38564
rect 189184 38010 189212 38558
rect 189172 38004 189224 38010
rect 189172 37946 189224 37952
rect 189172 30320 189224 30326
rect 189172 30262 189224 30268
rect 189184 29646 189212 30262
rect 189920 29646 189948 81110
rect 190196 80054 190224 86702
rect 190012 80026 190224 80054
rect 190012 77790 190040 80026
rect 190000 77784 190052 77790
rect 190000 77726 190052 77732
rect 190472 41410 190500 179046
rect 190564 142769 190592 266358
rect 190644 262404 190696 262410
rect 190644 262346 190696 262352
rect 190656 143478 190684 262346
rect 190736 260296 190788 260302
rect 190736 260238 190788 260244
rect 190748 145790 190776 260238
rect 190828 208956 190880 208962
rect 190828 208898 190880 208904
rect 190840 198626 190868 208898
rect 191116 199714 191144 364346
rect 191656 267028 191708 267034
rect 191656 266970 191708 266976
rect 191668 266422 191696 266970
rect 191656 266416 191708 266422
rect 191656 266358 191708 266364
rect 191196 260364 191248 260370
rect 191196 260306 191248 260312
rect 191208 217326 191236 260306
rect 191288 248464 191340 248470
rect 191288 248406 191340 248412
rect 191196 217320 191248 217326
rect 191196 217262 191248 217268
rect 191104 199708 191156 199714
rect 191104 199650 191156 199656
rect 190828 198620 190880 198626
rect 190828 198562 190880 198568
rect 190828 189984 190880 189990
rect 190828 189926 190880 189932
rect 190736 145784 190788 145790
rect 190736 145726 190788 145732
rect 190644 143472 190696 143478
rect 190644 143414 190696 143420
rect 190550 142760 190606 142769
rect 190550 142695 190606 142704
rect 190736 141228 190788 141234
rect 190736 141170 190788 141176
rect 190552 140004 190604 140010
rect 190552 139946 190604 139952
rect 190460 41404 190512 41410
rect 190460 41346 190512 41352
rect 190564 34474 190592 139946
rect 190642 138000 190698 138009
rect 190642 137935 190698 137944
rect 190656 60654 190684 137935
rect 190748 69834 190776 141170
rect 190840 76838 190868 189926
rect 190920 176112 190972 176118
rect 190920 176054 190972 176060
rect 190828 76832 190880 76838
rect 190828 76774 190880 76780
rect 190932 72962 190960 176054
rect 191208 142866 191236 217262
rect 191300 200666 191328 248406
rect 191656 237448 191708 237454
rect 191656 237390 191708 237396
rect 191380 205692 191432 205698
rect 191380 205634 191432 205640
rect 191288 200660 191340 200666
rect 191288 200602 191340 200608
rect 191392 198558 191420 205634
rect 191668 200394 191696 237390
rect 191760 200870 191788 400182
rect 191748 200864 191800 200870
rect 191748 200806 191800 200812
rect 191760 200598 191788 200806
rect 191748 200592 191800 200598
rect 191748 200534 191800 200540
rect 191656 200388 191708 200394
rect 191656 200330 191708 200336
rect 191748 198620 191800 198626
rect 191748 198562 191800 198568
rect 191380 198552 191432 198558
rect 191380 198494 191432 198500
rect 191760 198082 191788 198562
rect 191748 198076 191800 198082
rect 191748 198018 191800 198024
rect 191852 192642 191880 700470
rect 193220 700460 193272 700466
rect 193220 700402 193272 700408
rect 192484 699712 192536 699718
rect 192484 699654 192536 699660
rect 192116 262608 192168 262614
rect 192116 262550 192168 262556
rect 192024 195220 192076 195226
rect 192024 195162 192076 195168
rect 191840 192636 191892 192642
rect 191840 192578 191892 192584
rect 191932 189712 191984 189718
rect 191932 189654 191984 189660
rect 191380 148164 191432 148170
rect 191380 148106 191432 148112
rect 191196 142860 191248 142866
rect 191196 142802 191248 142808
rect 191286 140176 191342 140185
rect 191286 140111 191342 140120
rect 191196 139936 191248 139942
rect 191196 139878 191248 139884
rect 191102 138816 191158 138825
rect 191102 138751 191158 138760
rect 191010 136640 191066 136649
rect 191010 136575 191066 136584
rect 190920 72956 190972 72962
rect 190920 72898 190972 72904
rect 190736 69828 190788 69834
rect 190736 69770 190788 69776
rect 191024 66026 191052 136575
rect 191116 69018 191144 138751
rect 191208 77178 191236 139878
rect 191300 81025 191328 140111
rect 191392 137358 191420 148106
rect 191840 143744 191892 143750
rect 191840 143686 191892 143692
rect 191380 137352 191432 137358
rect 191380 137294 191432 137300
rect 191380 81184 191432 81190
rect 191380 81126 191432 81132
rect 191286 81016 191342 81025
rect 191286 80951 191342 80960
rect 191286 80880 191342 80889
rect 191286 80815 191342 80824
rect 191300 80617 191328 80815
rect 191286 80608 191342 80617
rect 191286 80543 191342 80552
rect 191392 80510 191420 81126
rect 191380 80504 191432 80510
rect 191380 80446 191432 80452
rect 191380 80096 191432 80102
rect 191380 80038 191432 80044
rect 191196 77172 191248 77178
rect 191196 77114 191248 77120
rect 191104 69012 191156 69018
rect 191104 68954 191156 68960
rect 191012 66020 191064 66026
rect 191012 65962 191064 65968
rect 191392 64530 191420 80038
rect 191380 64524 191432 64530
rect 191380 64466 191432 64472
rect 190644 60648 190696 60654
rect 190644 60590 190696 60596
rect 190552 34468 190604 34474
rect 190552 34410 190604 34416
rect 191748 34468 191800 34474
rect 191748 34410 191800 34416
rect 191760 33794 191788 34410
rect 191748 33788 191800 33794
rect 191748 33730 191800 33736
rect 189172 29640 189224 29646
rect 189172 29582 189224 29588
rect 189908 29640 189960 29646
rect 189908 29582 189960 29588
rect 191852 3602 191880 143686
rect 191944 57866 191972 189654
rect 192036 70922 192064 195162
rect 192128 143002 192156 262550
rect 192208 262268 192260 262274
rect 192208 262210 192260 262216
rect 192220 143206 192248 262210
rect 192496 199306 192524 699654
rect 192576 356108 192628 356114
rect 192576 356050 192628 356056
rect 192588 264246 192616 356050
rect 192576 264240 192628 264246
rect 192576 264182 192628 264188
rect 192576 262880 192628 262886
rect 192576 262822 192628 262828
rect 192484 199300 192536 199306
rect 192484 199242 192536 199248
rect 192484 197124 192536 197130
rect 192484 197066 192536 197072
rect 192300 194268 192352 194274
rect 192300 194210 192352 194216
rect 192208 143200 192260 143206
rect 192208 143142 192260 143148
rect 192116 142996 192168 143002
rect 192116 142938 192168 142944
rect 192208 141160 192260 141166
rect 192208 141102 192260 141108
rect 192024 70916 192076 70922
rect 192024 70858 192076 70864
rect 192220 70106 192248 141102
rect 192312 75818 192340 194210
rect 192392 189848 192444 189854
rect 192392 189790 192444 189796
rect 192300 75812 192352 75818
rect 192300 75754 192352 75760
rect 192404 72282 192432 189790
rect 192496 153202 192524 197066
rect 192484 153196 192536 153202
rect 192484 153138 192536 153144
rect 192588 145654 192616 262822
rect 192760 260908 192812 260914
rect 192760 260850 192812 260856
rect 192668 259956 192720 259962
rect 192668 259898 192720 259904
rect 192576 145648 192628 145654
rect 192576 145590 192628 145596
rect 192680 143138 192708 259898
rect 192772 252618 192800 260850
rect 192760 252612 192812 252618
rect 192760 252554 192812 252560
rect 193232 198286 193260 700402
rect 194520 699718 194548 703520
rect 198384 700330 198412 703520
rect 198372 700324 198424 700330
rect 198372 700266 198424 700272
rect 195980 699780 196032 699786
rect 195980 699722 196032 699728
rect 194508 699712 194560 699718
rect 194508 699654 194560 699660
rect 194600 372632 194652 372638
rect 194600 372574 194652 372580
rect 194508 349172 194560 349178
rect 194508 349114 194560 349120
rect 193496 265124 193548 265130
rect 193496 265066 193548 265072
rect 193312 265056 193364 265062
rect 193312 264998 193364 265004
rect 193220 198280 193272 198286
rect 193220 198222 193272 198228
rect 193232 197713 193260 198222
rect 193218 197704 193274 197713
rect 193218 197639 193274 197648
rect 192760 196648 192812 196654
rect 192760 196590 192812 196596
rect 192772 177410 192800 196590
rect 193220 195628 193272 195634
rect 193220 195570 193272 195576
rect 192760 177404 192812 177410
rect 192760 177346 192812 177352
rect 192760 147212 192812 147218
rect 192760 147154 192812 147160
rect 192668 143132 192720 143138
rect 192668 143074 192720 143080
rect 192484 140616 192536 140622
rect 192484 140558 192536 140564
rect 192496 75342 192524 140558
rect 192576 139868 192628 139874
rect 192576 139810 192628 139816
rect 192588 75410 192616 139810
rect 192772 138854 192800 147154
rect 192852 144152 192904 144158
rect 192852 144094 192904 144100
rect 192760 138848 192812 138854
rect 192760 138790 192812 138796
rect 192666 91896 192722 91905
rect 192666 91831 192722 91840
rect 192576 75404 192628 75410
rect 192576 75346 192628 75352
rect 192484 75336 192536 75342
rect 192484 75278 192536 75284
rect 192392 72276 192444 72282
rect 192392 72218 192444 72224
rect 192208 70100 192260 70106
rect 192208 70042 192260 70048
rect 192680 69630 192708 91831
rect 192668 69624 192720 69630
rect 192668 69566 192720 69572
rect 192864 67590 192892 144094
rect 193232 75002 193260 195570
rect 193324 142905 193352 264998
rect 193404 263220 193456 263226
rect 193404 263162 193456 263168
rect 193310 142896 193366 142905
rect 193310 142831 193366 142840
rect 193310 141808 193366 141817
rect 193310 141743 193366 141752
rect 193220 74996 193272 75002
rect 193220 74938 193272 74944
rect 193324 68610 193352 141743
rect 193416 140758 193444 263162
rect 193508 144838 193536 265066
rect 193680 260160 193732 260166
rect 193680 260102 193732 260108
rect 193588 195696 193640 195702
rect 193588 195638 193640 195644
rect 193496 144832 193548 144838
rect 193496 144774 193548 144780
rect 193404 140752 193456 140758
rect 193404 140694 193456 140700
rect 193416 140078 193444 140694
rect 193496 140412 193548 140418
rect 193496 140354 193548 140360
rect 193404 140072 193456 140078
rect 193404 140014 193456 140020
rect 193508 72554 193536 140354
rect 193600 77217 193628 195638
rect 193692 144770 193720 260102
rect 193772 259752 193824 259758
rect 193772 259694 193824 259700
rect 193784 146130 193812 259694
rect 194520 200462 194548 349114
rect 194508 200456 194560 200462
rect 194508 200398 194560 200404
rect 194520 198898 194548 200398
rect 194508 198892 194560 198898
rect 194508 198834 194560 198840
rect 194612 198694 194640 372574
rect 194784 264988 194836 264994
rect 194784 264930 194836 264936
rect 194692 263696 194744 263702
rect 194692 263638 194744 263644
rect 194600 198688 194652 198694
rect 194600 198630 194652 198636
rect 194612 198150 194640 198630
rect 194600 198144 194652 198150
rect 194600 198086 194652 198092
rect 194600 191344 194652 191350
rect 194600 191286 194652 191292
rect 193956 190392 194008 190398
rect 193956 190334 194008 190340
rect 193864 186992 193916 186998
rect 193864 186934 193916 186940
rect 193772 146124 193824 146130
rect 193772 146066 193824 146072
rect 193680 144764 193732 144770
rect 193680 144706 193732 144712
rect 193772 140684 193824 140690
rect 193772 140626 193824 140632
rect 193680 140208 193732 140214
rect 193680 140150 193732 140156
rect 193586 77208 193642 77217
rect 193586 77143 193642 77152
rect 193692 73953 193720 140150
rect 193784 77926 193812 140626
rect 193772 77920 193824 77926
rect 193772 77862 193824 77868
rect 193876 74526 193904 186934
rect 193968 76974 193996 190334
rect 194230 141944 194286 141953
rect 194230 141879 194286 141888
rect 194048 139324 194100 139330
rect 194048 139266 194100 139272
rect 194060 80578 194088 139266
rect 194048 80572 194100 80578
rect 194048 80514 194100 80520
rect 194048 79892 194100 79898
rect 194048 79834 194100 79840
rect 193956 76968 194008 76974
rect 193956 76910 194008 76916
rect 193864 74520 193916 74526
rect 193864 74462 193916 74468
rect 193678 73944 193734 73953
rect 193678 73879 193734 73888
rect 193496 72548 193548 72554
rect 193496 72490 193548 72496
rect 193312 68604 193364 68610
rect 193312 68546 193364 68552
rect 192852 67584 192904 67590
rect 192852 67526 192904 67532
rect 194060 62626 194088 79834
rect 194244 68542 194272 141879
rect 194506 77208 194562 77217
rect 194506 77143 194562 77152
rect 194520 75206 194548 77143
rect 194508 75200 194560 75206
rect 194508 75142 194560 75148
rect 194612 72486 194640 191286
rect 194704 143313 194732 263638
rect 194796 145926 194824 264930
rect 195060 264240 195112 264246
rect 195060 264182 195112 264188
rect 195072 263702 195100 264182
rect 195060 263696 195112 263702
rect 195060 263638 195112 263644
rect 194968 263628 195020 263634
rect 194968 263570 195020 263576
rect 194876 259480 194928 259486
rect 194876 259422 194928 259428
rect 194784 145920 194836 145926
rect 194784 145862 194836 145868
rect 194784 144220 194836 144226
rect 194784 144162 194836 144168
rect 194690 143304 194746 143313
rect 194690 143239 194746 143248
rect 194600 72480 194652 72486
rect 194600 72422 194652 72428
rect 194796 70038 194824 144162
rect 194888 141846 194916 259422
rect 194980 145722 195008 263570
rect 195060 260092 195112 260098
rect 195060 260034 195112 260040
rect 194968 145716 195020 145722
rect 194968 145658 195020 145664
rect 195072 143342 195100 260034
rect 195992 191486 196020 699722
rect 199384 698352 199436 698358
rect 199384 698294 199436 698300
rect 196624 380928 196676 380934
rect 196624 380870 196676 380876
rect 196072 265736 196124 265742
rect 196072 265678 196124 265684
rect 196084 198218 196112 265678
rect 196636 265062 196664 380870
rect 199396 267102 199424 698294
rect 200764 673532 200816 673538
rect 200764 673474 200816 673480
rect 199384 267096 199436 267102
rect 199384 267038 199436 267044
rect 197544 265192 197596 265198
rect 197544 265134 197596 265140
rect 196624 265056 196676 265062
rect 196624 264998 196676 265004
rect 196624 262472 196676 262478
rect 196624 262414 196676 262420
rect 196440 260228 196492 260234
rect 196440 260170 196492 260176
rect 196256 259888 196308 259894
rect 196256 259830 196308 259836
rect 196164 259684 196216 259690
rect 196164 259626 196216 259632
rect 196072 198212 196124 198218
rect 196072 198154 196124 198160
rect 196072 192772 196124 192778
rect 196072 192714 196124 192720
rect 195980 191480 196032 191486
rect 195980 191422 196032 191428
rect 195980 186856 196032 186862
rect 195980 186798 196032 186804
rect 195152 181688 195204 181694
rect 195152 181630 195204 181636
rect 195164 180878 195192 181630
rect 195152 180872 195204 180878
rect 195152 180814 195204 180820
rect 195060 143336 195112 143342
rect 195060 143278 195112 143284
rect 194876 141840 194928 141846
rect 194876 141782 194928 141788
rect 194874 141672 194930 141681
rect 194874 141607 194930 141616
rect 194784 70032 194836 70038
rect 194784 69974 194836 69980
rect 194888 68950 194916 141607
rect 195058 140584 195114 140593
rect 195058 140519 195114 140528
rect 194968 140140 195020 140146
rect 194968 140082 195020 140088
rect 194980 72894 195008 140082
rect 195072 74186 195100 140519
rect 195060 74180 195112 74186
rect 195060 74122 195112 74128
rect 194968 72888 195020 72894
rect 194968 72830 195020 72836
rect 195164 72350 195192 180814
rect 195428 148980 195480 148986
rect 195428 148922 195480 148928
rect 195242 141400 195298 141409
rect 195242 141335 195298 141344
rect 195256 79354 195284 141335
rect 195334 139088 195390 139097
rect 195334 139023 195390 139032
rect 195244 79348 195296 79354
rect 195244 79290 195296 79296
rect 195348 78033 195376 139023
rect 195440 137698 195468 148922
rect 195518 144392 195574 144401
rect 195518 144327 195574 144336
rect 195428 137692 195480 137698
rect 195428 137634 195480 137640
rect 195334 78024 195390 78033
rect 195334 77959 195390 77968
rect 195152 72344 195204 72350
rect 195152 72286 195204 72292
rect 194876 68944 194928 68950
rect 194876 68886 194928 68892
rect 194232 68536 194284 68542
rect 194232 68478 194284 68484
rect 195532 65754 195560 144327
rect 195992 73098 196020 186798
rect 195980 73092 196032 73098
rect 195980 73034 196032 73040
rect 196084 72593 196112 192714
rect 196176 143410 196204 259626
rect 196268 146266 196296 259830
rect 196348 259820 196400 259826
rect 196348 259762 196400 259768
rect 196256 146260 196308 146266
rect 196256 146202 196308 146208
rect 196360 146062 196388 259762
rect 196452 147286 196480 260170
rect 196532 252612 196584 252618
rect 196532 252554 196584 252560
rect 196440 147280 196492 147286
rect 196440 147222 196492 147228
rect 196348 146056 196400 146062
rect 196348 145998 196400 146004
rect 196544 145518 196572 252554
rect 196532 145512 196584 145518
rect 196532 145454 196584 145460
rect 196532 144492 196584 144498
rect 196532 144434 196584 144440
rect 196440 144424 196492 144430
rect 196440 144366 196492 144372
rect 196348 143676 196400 143682
rect 196348 143618 196400 143624
rect 196256 143540 196308 143546
rect 196256 143482 196308 143488
rect 196164 143404 196216 143410
rect 196164 143346 196216 143352
rect 196164 141976 196216 141982
rect 196164 141918 196216 141924
rect 196070 72584 196126 72593
rect 196070 72519 196126 72528
rect 195520 65748 195572 65754
rect 195520 65690 195572 65696
rect 194048 62620 194100 62626
rect 194048 62562 194100 62568
rect 192484 60648 192536 60654
rect 192484 60590 192536 60596
rect 191932 57860 191984 57866
rect 191932 57802 191984 57808
rect 192496 37262 192524 60590
rect 193128 57860 193180 57866
rect 193128 57802 193180 57808
rect 193140 57322 193168 57802
rect 193128 57316 193180 57322
rect 193128 57258 193180 57264
rect 196176 51066 196204 141918
rect 196268 68678 196296 143482
rect 196360 142934 196388 143618
rect 196348 142928 196400 142934
rect 196348 142870 196400 142876
rect 196346 137456 196402 137465
rect 196346 137391 196402 137400
rect 196256 68672 196308 68678
rect 196256 68614 196308 68620
rect 196360 66978 196388 137391
rect 196452 78130 196480 144366
rect 196544 78198 196572 144434
rect 196636 143682 196664 262414
rect 197452 261044 197504 261050
rect 197452 260986 197504 260992
rect 197358 195120 197414 195129
rect 197358 195055 197414 195064
rect 196716 192704 196768 192710
rect 196716 192646 196768 192652
rect 196624 143676 196676 143682
rect 196624 143618 196676 143624
rect 196624 141296 196676 141302
rect 196624 141238 196676 141244
rect 196636 80850 196664 141238
rect 196728 133210 196756 192646
rect 197372 191350 197400 195055
rect 197360 191344 197412 191350
rect 197360 191286 197412 191292
rect 197360 191072 197412 191078
rect 197360 191014 197412 191020
rect 197372 190913 197400 191014
rect 197082 190904 197138 190913
rect 197082 190839 197138 190848
rect 197358 190904 197414 190913
rect 197358 190839 197414 190848
rect 197096 190641 197124 190839
rect 197082 190632 197138 190641
rect 197082 190567 197138 190576
rect 197360 155236 197412 155242
rect 197360 155178 197412 155184
rect 196806 134464 196862 134473
rect 196806 134399 196862 134408
rect 196716 133204 196768 133210
rect 196716 133146 196768 133152
rect 196820 83473 196848 134399
rect 196806 83464 196862 83473
rect 196806 83399 196862 83408
rect 196624 80844 196676 80850
rect 196624 80786 196676 80792
rect 196532 78192 196584 78198
rect 196532 78134 196584 78140
rect 196440 78124 196492 78130
rect 196440 78066 196492 78072
rect 196440 76560 196492 76566
rect 196440 76502 196492 76508
rect 196452 75886 196480 76502
rect 196440 75880 196492 75886
rect 196440 75822 196492 75828
rect 196348 66972 196400 66978
rect 196348 66914 196400 66920
rect 196164 51060 196216 51066
rect 196164 51002 196216 51008
rect 196176 50386 196204 51002
rect 196164 50380 196216 50386
rect 196164 50322 196216 50328
rect 192484 37256 192536 37262
rect 192484 37198 192536 37204
rect 191930 34504 191986 34513
rect 191930 34439 191986 34448
rect 191944 34406 191972 34439
rect 191932 34400 191984 34406
rect 191932 34342 191984 34348
rect 193128 34400 193180 34406
rect 193128 34342 193180 34348
rect 193140 33182 193168 34342
rect 193128 33176 193180 33182
rect 193128 33118 193180 33124
rect 196452 16574 196480 75822
rect 197372 73166 197400 155178
rect 197464 142118 197492 260986
rect 197556 145450 197584 265134
rect 200776 263634 200804 673474
rect 200764 263628 200816 263634
rect 200764 263570 200816 263576
rect 198924 263152 198976 263158
rect 198924 263094 198976 263100
rect 198740 263084 198792 263090
rect 198740 263026 198792 263032
rect 197820 262812 197872 262818
rect 197820 262754 197872 262760
rect 197728 191684 197780 191690
rect 197728 191626 197780 191632
rect 197740 191078 197768 191626
rect 197728 191072 197780 191078
rect 197728 191014 197780 191020
rect 197728 190052 197780 190058
rect 197728 189994 197780 190000
rect 197544 145444 197596 145450
rect 197544 145386 197596 145392
rect 197636 144696 197688 144702
rect 197636 144638 197688 144644
rect 197544 144560 197596 144566
rect 197544 144502 197596 144508
rect 197452 142112 197504 142118
rect 197452 142054 197504 142060
rect 197452 138780 197504 138786
rect 197452 138722 197504 138728
rect 197360 73160 197412 73166
rect 197360 73102 197412 73108
rect 197464 62762 197492 138722
rect 197556 68746 197584 144502
rect 197648 71602 197676 144638
rect 197740 72758 197768 189994
rect 197832 145858 197860 262754
rect 198372 262744 198424 262750
rect 198372 262686 198424 262692
rect 197912 260024 197964 260030
rect 197912 259966 197964 259972
rect 197820 145852 197872 145858
rect 197820 145794 197872 145800
rect 197924 145382 197952 259966
rect 198004 195560 198056 195566
rect 198004 195502 198056 195508
rect 198016 191758 198044 195502
rect 198096 193248 198148 193254
rect 198096 193190 198148 193196
rect 198004 191752 198056 191758
rect 198004 191694 198056 191700
rect 197912 145376 197964 145382
rect 197912 145318 197964 145324
rect 197820 143268 197872 143274
rect 197820 143210 197872 143216
rect 197832 142866 197860 143210
rect 197820 142860 197872 142866
rect 197820 142802 197872 142808
rect 197912 141568 197964 141574
rect 197912 141510 197964 141516
rect 197820 140344 197872 140350
rect 197820 140286 197872 140292
rect 197728 72752 197780 72758
rect 197728 72694 197780 72700
rect 197636 71596 197688 71602
rect 197636 71538 197688 71544
rect 197832 69698 197860 140286
rect 197924 78062 197952 141510
rect 197912 78056 197964 78062
rect 197912 77998 197964 78004
rect 198016 74118 198044 191694
rect 198108 157350 198136 193190
rect 198096 157344 198148 157350
rect 198096 157286 198148 157292
rect 198384 142866 198412 262686
rect 198464 262676 198516 262682
rect 198464 262618 198516 262624
rect 198476 144265 198504 262618
rect 198752 262546 198780 263026
rect 198830 262984 198886 262993
rect 198830 262919 198886 262928
rect 198740 262540 198792 262546
rect 198740 262482 198792 262488
rect 198844 262449 198872 262919
rect 198936 262886 198964 263094
rect 198924 262880 198976 262886
rect 198924 262822 198976 262828
rect 199568 262880 199620 262886
rect 199568 262822 199620 262828
rect 199200 262540 199252 262546
rect 199200 262482 199252 262488
rect 198830 262440 198886 262449
rect 198830 262375 198886 262384
rect 199106 262440 199162 262449
rect 199106 262375 199162 262384
rect 198924 259616 198976 259622
rect 198924 259558 198976 259564
rect 198832 194200 198884 194206
rect 198832 194142 198884 194148
rect 198740 192976 198792 192982
rect 198740 192918 198792 192924
rect 198462 144256 198518 144265
rect 198462 144191 198518 144200
rect 198372 142860 198424 142866
rect 198372 142802 198424 142808
rect 198096 140276 198148 140282
rect 198096 140218 198148 140224
rect 198108 81190 198136 140218
rect 198186 135960 198242 135969
rect 198186 135895 198242 135904
rect 198096 81184 198148 81190
rect 198096 81126 198148 81132
rect 198200 80102 198228 135895
rect 198188 80096 198240 80102
rect 198188 80038 198240 80044
rect 198004 74112 198056 74118
rect 198004 74054 198056 74060
rect 198752 69766 198780 192918
rect 198844 75478 198872 194142
rect 198936 141914 198964 259558
rect 199120 145994 199148 262375
rect 199212 146198 199240 262482
rect 199384 187332 199436 187338
rect 199384 187274 199436 187280
rect 199292 187196 199344 187202
rect 199292 187138 199344 187144
rect 199200 146192 199252 146198
rect 199200 146134 199252 146140
rect 199108 145988 199160 145994
rect 199108 145930 199160 145936
rect 199016 144628 199068 144634
rect 199016 144570 199068 144576
rect 198924 141908 198976 141914
rect 198924 141850 198976 141856
rect 198936 141574 198964 141850
rect 198924 141568 198976 141574
rect 198924 141510 198976 141516
rect 198832 75472 198884 75478
rect 198832 75414 198884 75420
rect 198740 69760 198792 69766
rect 198740 69702 198792 69708
rect 197820 69692 197872 69698
rect 197820 69634 197872 69640
rect 197544 68740 197596 68746
rect 197544 68682 197596 68688
rect 197452 62756 197504 62762
rect 197452 62698 197504 62704
rect 199028 60722 199056 144570
rect 199200 141772 199252 141778
rect 199200 141714 199252 141720
rect 199106 137320 199162 137329
rect 199106 137255 199162 137264
rect 198740 60716 198792 60722
rect 198740 60658 198792 60664
rect 199016 60716 199068 60722
rect 199016 60658 199068 60664
rect 198752 59906 198780 60658
rect 198740 59900 198792 59906
rect 198740 59842 198792 59848
rect 199120 55146 199148 137255
rect 199108 55140 199160 55146
rect 199108 55082 199160 55088
rect 199212 49706 199240 141714
rect 199304 75682 199332 187138
rect 199396 76702 199424 187274
rect 199476 153196 199528 153202
rect 199476 153138 199528 153144
rect 199488 151842 199516 153138
rect 199476 151836 199528 151842
rect 199476 151778 199528 151784
rect 199384 76696 199436 76702
rect 199384 76638 199436 76644
rect 199292 75676 199344 75682
rect 199292 75618 199344 75624
rect 199488 70310 199516 151778
rect 199580 144129 199608 262822
rect 200120 200456 200172 200462
rect 200120 200398 200172 200404
rect 199660 148504 199712 148510
rect 199660 148446 199712 148452
rect 199566 144120 199622 144129
rect 199566 144055 199622 144064
rect 199568 137692 199620 137698
rect 199568 137634 199620 137640
rect 199476 70304 199528 70310
rect 199476 70246 199528 70252
rect 199580 63170 199608 137634
rect 199672 67114 199700 148446
rect 200132 74089 200160 200398
rect 200764 197056 200816 197062
rect 200764 196998 200816 197004
rect 200304 196988 200356 196994
rect 200304 196930 200356 196936
rect 200212 191276 200264 191282
rect 200212 191218 200264 191224
rect 200118 74080 200174 74089
rect 200118 74015 200174 74024
rect 199660 67108 199712 67114
rect 199660 67050 199712 67056
rect 199568 63164 199620 63170
rect 199568 63106 199620 63112
rect 200120 59900 200172 59906
rect 200120 59842 200172 59848
rect 199200 49700 199252 49706
rect 199200 49642 199252 49648
rect 200132 16574 200160 59842
rect 200224 55214 200252 191218
rect 200316 76770 200344 196930
rect 200486 195664 200542 195673
rect 200486 195599 200542 195608
rect 200396 191412 200448 191418
rect 200396 191354 200448 191360
rect 200304 76764 200356 76770
rect 200304 76706 200356 76712
rect 200408 74322 200436 191354
rect 200500 187377 200528 195599
rect 200776 195294 200804 196998
rect 200764 195288 200816 195294
rect 200764 195230 200816 195236
rect 201512 188834 201540 703582
rect 202064 703474 202092 703582
rect 202206 703520 202318 704960
rect 205652 703582 205956 703610
rect 202248 703474 202276 703520
rect 202064 703446 202276 703474
rect 202788 206304 202840 206310
rect 202788 206246 202840 206252
rect 202800 205698 202828 206246
rect 201684 205692 201736 205698
rect 201684 205634 201736 205640
rect 202788 205692 202840 205698
rect 202788 205634 202840 205640
rect 201592 198212 201644 198218
rect 201592 198154 201644 198160
rect 201500 188828 201552 188834
rect 201500 188770 201552 188776
rect 201512 187746 201540 188770
rect 201500 187740 201552 187746
rect 201500 187682 201552 187688
rect 200486 187368 200542 187377
rect 200486 187303 200542 187312
rect 201500 186924 201552 186930
rect 201500 186866 201552 186872
rect 200488 184748 200540 184754
rect 200488 184690 200540 184696
rect 200396 74316 200448 74322
rect 200396 74258 200448 74264
rect 200500 73030 200528 184690
rect 200672 148640 200724 148646
rect 200672 148582 200724 148588
rect 200580 148572 200632 148578
rect 200580 148514 200632 148520
rect 200488 73024 200540 73030
rect 200488 72966 200540 72972
rect 200592 66842 200620 148514
rect 200684 67182 200712 148582
rect 200764 148232 200816 148238
rect 200764 148174 200816 148180
rect 200776 67318 200804 148174
rect 200856 138848 200908 138854
rect 200856 138790 200908 138796
rect 200868 79898 200896 138790
rect 200948 107704 201000 107710
rect 200948 107646 201000 107652
rect 200856 79892 200908 79898
rect 200856 79834 200908 79840
rect 200960 77110 200988 107646
rect 200948 77104 201000 77110
rect 200948 77046 201000 77052
rect 200764 67312 200816 67318
rect 200764 67254 200816 67260
rect 200672 67176 200724 67182
rect 200672 67118 200724 67124
rect 200580 66836 200632 66842
rect 200580 66778 200632 66784
rect 200212 55208 200264 55214
rect 200212 55150 200264 55156
rect 201408 55208 201460 55214
rect 201408 55150 201460 55156
rect 201420 54534 201448 55150
rect 201408 54528 201460 54534
rect 201408 54470 201460 54476
rect 201512 53786 201540 186866
rect 201604 64297 201632 198154
rect 201696 77246 201724 205634
rect 204536 200864 204588 200870
rect 204536 200806 204588 200812
rect 204352 198280 204404 198286
rect 204352 198222 204404 198228
rect 204260 195424 204312 195430
rect 204260 195366 204312 195372
rect 202880 192840 202932 192846
rect 202880 192782 202932 192788
rect 202892 192642 202920 192782
rect 202880 192636 202932 192642
rect 202880 192578 202932 192584
rect 201774 190904 201830 190913
rect 201774 190839 201830 190848
rect 201684 77240 201736 77246
rect 201684 77182 201736 77188
rect 201788 65686 201816 190839
rect 201960 187128 202012 187134
rect 201960 187070 202012 187076
rect 201868 184612 201920 184618
rect 201868 184554 201920 184560
rect 201880 68882 201908 184554
rect 201972 72826 202000 187070
rect 202234 148336 202290 148345
rect 202234 148271 202290 148280
rect 202144 147076 202196 147082
rect 202144 147018 202196 147024
rect 202052 144356 202104 144362
rect 202052 144298 202104 144304
rect 201960 72820 202012 72826
rect 201960 72762 202012 72768
rect 201868 68876 201920 68882
rect 201868 68818 201920 68824
rect 201776 65680 201828 65686
rect 201776 65622 201828 65628
rect 201590 64288 201646 64297
rect 201590 64223 201646 64232
rect 202064 63102 202092 144298
rect 202156 70174 202184 147018
rect 202248 77994 202276 148271
rect 202326 138952 202382 138961
rect 202326 138887 202382 138896
rect 202340 93854 202368 138887
rect 202340 93826 202460 93854
rect 202432 81054 202460 93826
rect 202420 81048 202472 81054
rect 202420 80990 202472 80996
rect 202236 77988 202288 77994
rect 202236 77930 202288 77936
rect 202892 71194 202920 192578
rect 203064 187400 203116 187406
rect 203064 187342 203116 187348
rect 202972 186788 203024 186794
rect 202972 186730 203024 186736
rect 202880 71188 202932 71194
rect 202880 71130 202932 71136
rect 202144 70168 202196 70174
rect 202144 70110 202196 70116
rect 202984 69737 203012 186730
rect 203076 79694 203104 187342
rect 203248 148844 203300 148850
rect 203248 148786 203300 148792
rect 203154 148472 203210 148481
rect 203154 148407 203210 148416
rect 203064 79688 203116 79694
rect 203064 79630 203116 79636
rect 202970 69728 203026 69737
rect 202970 69663 203026 69672
rect 202052 63096 202104 63102
rect 202052 63038 202104 63044
rect 201500 53780 201552 53786
rect 201500 53722 201552 53728
rect 202788 53780 202840 53786
rect 202788 53722 202840 53728
rect 202800 53174 202828 53722
rect 202788 53168 202840 53174
rect 202788 53110 202840 53116
rect 203168 46918 203196 148407
rect 203260 48210 203288 148786
rect 203432 148776 203484 148782
rect 203432 148718 203484 148724
rect 203340 148708 203392 148714
rect 203340 148650 203392 148656
rect 203352 62082 203380 148650
rect 203444 62830 203472 148718
rect 203616 148436 203668 148442
rect 203616 148378 203668 148384
rect 203524 147144 203576 147150
rect 203524 147086 203576 147092
rect 203432 62824 203484 62830
rect 203432 62766 203484 62772
rect 203536 62694 203564 147086
rect 203628 78334 203656 148378
rect 203708 137352 203760 137358
rect 203708 137294 203760 137300
rect 203616 78328 203668 78334
rect 203616 78270 203668 78276
rect 203720 67250 203748 137294
rect 203708 67244 203760 67250
rect 203708 67186 203760 67192
rect 204272 63374 204300 195366
rect 204364 70009 204392 198222
rect 204444 196104 204496 196110
rect 204444 196046 204496 196052
rect 204456 71330 204484 196046
rect 204548 80986 204576 200806
rect 204720 196920 204772 196926
rect 204720 196862 204772 196868
rect 204732 196110 204760 196862
rect 204720 196104 204772 196110
rect 204720 196046 204772 196052
rect 204812 187060 204864 187066
rect 204812 187002 204864 187008
rect 204720 184408 204772 184414
rect 204626 184376 204682 184385
rect 204720 184350 204772 184356
rect 204626 184311 204682 184320
rect 204536 80980 204588 80986
rect 204536 80922 204588 80928
rect 204444 71324 204496 71330
rect 204444 71266 204496 71272
rect 204350 70000 204406 70009
rect 204350 69935 204406 69944
rect 204640 65793 204668 184311
rect 204732 65958 204760 184350
rect 204824 70281 204852 187002
rect 205652 185910 205680 703582
rect 205928 703474 205956 703582
rect 206070 703520 206182 704960
rect 209934 703520 210046 704960
rect 213798 703520 213910 704960
rect 217018 703520 217130 704960
rect 220882 703520 220994 704960
rect 224746 703520 224858 704960
rect 228610 703520 228722 704960
rect 232474 703520 232586 704960
rect 236338 703520 236450 704960
rect 240202 703520 240314 704960
rect 244066 703520 244178 704960
rect 247930 703520 248042 704960
rect 251794 703520 251906 704960
rect 253952 703582 254900 703610
rect 206112 703474 206140 703520
rect 205928 703446 206140 703474
rect 209976 702434 210004 703520
rect 209976 702406 210648 702434
rect 208398 220960 208454 220969
rect 208398 220895 208454 220904
rect 208412 220862 208440 220895
rect 208400 220856 208452 220862
rect 208400 220798 208452 220804
rect 207018 197024 207074 197033
rect 207018 196959 207074 196968
rect 207032 196761 207060 196959
rect 207018 196752 207074 196761
rect 207018 196687 207074 196696
rect 207202 196752 207258 196761
rect 207202 196687 207258 196696
rect 206284 195016 206336 195022
rect 206284 194958 206336 194964
rect 205732 193860 205784 193866
rect 205732 193802 205784 193808
rect 205640 185904 205692 185910
rect 205640 185846 205692 185852
rect 204904 184680 204956 184686
rect 204904 184622 204956 184628
rect 204916 72622 204944 184622
rect 204996 164892 205048 164898
rect 204996 164834 205048 164840
rect 205008 164286 205036 164834
rect 204996 164280 205048 164286
rect 204996 164222 205048 164228
rect 205008 81977 205036 164222
rect 205088 151292 205140 151298
rect 205088 151234 205140 151240
rect 204994 81968 205050 81977
rect 204994 81903 205050 81912
rect 205100 75546 205128 151234
rect 205088 75540 205140 75546
rect 205088 75482 205140 75488
rect 204904 72616 204956 72622
rect 204904 72558 204956 72564
rect 204810 70272 204866 70281
rect 204810 70207 204866 70216
rect 204720 65952 204772 65958
rect 204720 65894 204772 65900
rect 204626 65784 204682 65793
rect 204626 65719 204682 65728
rect 204260 63368 204312 63374
rect 204260 63310 204312 63316
rect 203524 62688 203576 62694
rect 203524 62630 203576 62636
rect 203340 62076 203392 62082
rect 203340 62018 203392 62024
rect 203352 61402 203380 62018
rect 203340 61396 203392 61402
rect 203340 61338 203392 61344
rect 205744 55214 205772 193802
rect 206192 192908 206244 192914
rect 206192 192850 206244 192856
rect 205824 190256 205876 190262
rect 205824 190198 205876 190204
rect 205836 69902 205864 190198
rect 206100 188692 206152 188698
rect 206100 188634 206152 188640
rect 205916 184544 205968 184550
rect 205916 184486 205968 184492
rect 205824 69896 205876 69902
rect 205824 69838 205876 69844
rect 205928 65890 205956 184486
rect 206008 184476 206060 184482
rect 206008 184418 206060 184424
rect 205916 65884 205968 65890
rect 205916 65826 205968 65832
rect 206020 65822 206048 184418
rect 206112 69970 206140 188634
rect 206204 74050 206232 192850
rect 206296 190398 206324 194958
rect 207020 193996 207072 194002
rect 207020 193938 207072 193944
rect 207032 193866 207060 193938
rect 207020 193860 207072 193866
rect 207020 193802 207072 193808
rect 206560 191208 206612 191214
rect 206560 191150 206612 191156
rect 206284 190392 206336 190398
rect 206284 190334 206336 190340
rect 206284 184340 206336 184346
rect 206284 184282 206336 184288
rect 206296 78470 206324 184282
rect 206376 184272 206428 184278
rect 206376 184214 206428 184220
rect 206388 81705 206416 184214
rect 206468 148300 206520 148306
rect 206468 148242 206520 148248
rect 206374 81696 206430 81705
rect 206374 81631 206430 81640
rect 206284 78464 206336 78470
rect 206284 78406 206336 78412
rect 206192 74044 206244 74050
rect 206192 73986 206244 73992
rect 206480 71058 206508 148242
rect 206468 71052 206520 71058
rect 206468 70994 206520 71000
rect 206100 69964 206152 69970
rect 206100 69906 206152 69912
rect 206008 65816 206060 65822
rect 206008 65758 206060 65764
rect 206572 63306 206600 191150
rect 207032 74202 207060 193802
rect 207112 187740 207164 187746
rect 207112 187682 207164 187688
rect 207124 74534 207152 187682
rect 207216 78441 207244 196687
rect 207664 191208 207716 191214
rect 207664 191150 207716 191156
rect 207676 190454 207704 191150
rect 207584 190426 207704 190454
rect 207388 188896 207440 188902
rect 207388 188838 207440 188844
rect 207296 188284 207348 188290
rect 207296 188226 207348 188232
rect 207202 78432 207258 78441
rect 207202 78367 207258 78376
rect 207124 74506 207244 74534
rect 207032 74174 207152 74202
rect 207018 74080 207074 74089
rect 207018 74015 207074 74024
rect 207032 73982 207060 74015
rect 207020 73976 207072 73982
rect 207020 73918 207072 73924
rect 207124 71369 207152 74174
rect 207110 71360 207166 71369
rect 207110 71295 207166 71304
rect 207216 67522 207244 74506
rect 207308 71262 207336 188226
rect 207400 71534 207428 188838
rect 207584 186017 207612 190426
rect 207756 189848 207808 189854
rect 207756 189790 207808 189796
rect 207768 188902 207796 189790
rect 207756 188896 207808 188902
rect 207756 188838 207808 188844
rect 207570 186008 207626 186017
rect 207570 185943 207626 185952
rect 207480 185020 207532 185026
rect 207480 184962 207532 184968
rect 207388 71528 207440 71534
rect 207388 71470 207440 71476
rect 207296 71256 207348 71262
rect 207296 71198 207348 71204
rect 207492 68474 207520 184962
rect 207584 81326 207612 185943
rect 207664 175976 207716 175982
rect 207664 175918 207716 175924
rect 207572 81320 207624 81326
rect 207572 81262 207624 81268
rect 207676 80714 207704 175918
rect 207756 149048 207808 149054
rect 207756 148990 207808 148996
rect 207664 80708 207716 80714
rect 207664 80650 207716 80656
rect 207768 70990 207796 148990
rect 207848 144288 207900 144294
rect 207848 144230 207900 144236
rect 207756 70984 207808 70990
rect 207756 70926 207808 70932
rect 207860 70378 207888 144230
rect 208412 72690 208440 220798
rect 209318 202192 209374 202201
rect 209318 202127 209374 202136
rect 209332 201521 209360 202127
rect 208490 201512 208546 201521
rect 208490 201447 208546 201456
rect 209318 201512 209374 201521
rect 209318 201447 209374 201456
rect 208400 72684 208452 72690
rect 208400 72626 208452 72632
rect 207848 70372 207900 70378
rect 207848 70314 207900 70320
rect 207480 68468 207532 68474
rect 207480 68410 207532 68416
rect 207204 67516 207256 67522
rect 207204 67458 207256 67464
rect 208504 67153 208532 201447
rect 209964 200320 210016 200326
rect 209964 200262 210016 200268
rect 209872 194064 209924 194070
rect 209872 194006 209924 194012
rect 208676 185972 208728 185978
rect 208676 185914 208728 185920
rect 208584 184204 208636 184210
rect 208584 184146 208636 184152
rect 208490 67144 208546 67153
rect 208490 67079 208546 67088
rect 208596 65482 208624 184146
rect 208688 67289 208716 185914
rect 208858 185600 208914 185609
rect 208858 185535 208914 185544
rect 208768 183388 208820 183394
rect 208768 183330 208820 183336
rect 208780 68202 208808 183330
rect 208872 74225 208900 185535
rect 209780 183252 209832 183258
rect 209780 183194 209832 183200
rect 208952 176044 209004 176050
rect 208952 175986 209004 175992
rect 208964 74254 208992 175986
rect 209136 151224 209188 151230
rect 209136 151166 209188 151172
rect 209044 151156 209096 151162
rect 209044 151098 209096 151104
rect 209056 77042 209084 151098
rect 209148 81122 209176 151166
rect 209136 81116 209188 81122
rect 209136 81058 209188 81064
rect 209044 77036 209096 77042
rect 209044 76978 209096 76984
rect 208952 74248 209004 74254
rect 208858 74216 208914 74225
rect 208952 74190 209004 74196
rect 208858 74151 208914 74160
rect 208768 68196 208820 68202
rect 208768 68138 208820 68144
rect 208674 67280 208730 67289
rect 208674 67215 208730 67224
rect 208584 65476 208636 65482
rect 208584 65418 208636 65424
rect 206560 63300 206612 63306
rect 206560 63242 206612 63248
rect 209792 63238 209820 183194
rect 209884 71398 209912 194006
rect 209976 77897 210004 200262
rect 210424 191140 210476 191146
rect 210424 191082 210476 191088
rect 210148 188624 210200 188630
rect 210148 188566 210200 188572
rect 210056 186108 210108 186114
rect 210056 186050 210108 186056
rect 209962 77888 210018 77897
rect 209962 77823 210018 77832
rect 209872 71392 209924 71398
rect 209872 71334 209924 71340
rect 210068 67046 210096 186050
rect 210160 71466 210188 188566
rect 210240 187264 210292 187270
rect 210240 187206 210292 187212
rect 210148 71460 210200 71466
rect 210148 71402 210200 71408
rect 210252 70242 210280 187206
rect 210332 181756 210384 181762
rect 210332 181698 210384 181704
rect 210240 70236 210292 70242
rect 210240 70178 210292 70184
rect 210056 67040 210108 67046
rect 210056 66982 210108 66988
rect 210344 65346 210372 181698
rect 210436 77654 210464 191082
rect 210516 186040 210568 186046
rect 210516 185982 210568 185988
rect 210528 78946 210556 185982
rect 210620 181898 210648 702406
rect 220924 683114 220952 703520
rect 228652 702434 228680 703520
rect 232516 702434 232544 703520
rect 236380 702434 236408 703520
rect 220832 683086 220952 683114
rect 227732 702406 228680 702434
rect 231872 702406 232544 702434
rect 236012 702406 236408 702434
rect 215944 484424 215996 484430
rect 215944 484366 215996 484372
rect 215956 264246 215984 484366
rect 215944 264240 215996 264246
rect 215944 264182 215996 264188
rect 211160 262336 211212 262342
rect 211160 262278 211212 262284
rect 211068 200932 211120 200938
rect 211068 200874 211120 200880
rect 211080 200326 211108 200874
rect 211068 200320 211120 200326
rect 211068 200262 211120 200268
rect 210608 181892 210660 181898
rect 210608 181834 210660 181840
rect 210608 148912 210660 148918
rect 210608 148854 210660 148860
rect 210620 79286 210648 148854
rect 210608 79280 210660 79286
rect 210608 79222 210660 79228
rect 210516 78940 210568 78946
rect 210516 78882 210568 78888
rect 210424 77648 210476 77654
rect 210424 77590 210476 77596
rect 211172 68270 211200 262278
rect 214104 200388 214156 200394
rect 214104 200330 214156 200336
rect 212540 198144 212592 198150
rect 212540 198086 212592 198092
rect 211436 198076 211488 198082
rect 211436 198018 211488 198024
rect 211344 183184 211396 183190
rect 211344 183126 211396 183132
rect 211252 143064 211304 143070
rect 211252 143006 211304 143012
rect 211160 68264 211212 68270
rect 211160 68206 211212 68212
rect 210332 65340 210384 65346
rect 210332 65282 210384 65288
rect 209780 63232 209832 63238
rect 209780 63174 209832 63180
rect 205652 55186 205772 55214
rect 203248 48204 203300 48210
rect 203248 48146 203300 48152
rect 204168 48204 204220 48210
rect 204168 48146 204220 48152
rect 204180 47666 204208 48146
rect 204168 47660 204220 47666
rect 204168 47602 204220 47608
rect 203156 46912 203208 46918
rect 203156 46854 203208 46860
rect 204168 46912 204220 46918
rect 204168 46854 204220 46860
rect 204180 46238 204208 46854
rect 205652 46850 205680 55186
rect 205640 46844 205692 46850
rect 205640 46786 205692 46792
rect 205652 46306 205680 46786
rect 205640 46300 205692 46306
rect 205640 46242 205692 46248
rect 204168 46232 204220 46238
rect 204168 46174 204220 46180
rect 207664 28280 207716 28286
rect 207664 28222 207716 28228
rect 196452 16546 196664 16574
rect 200132 16546 200528 16574
rect 193220 11756 193272 11762
rect 193220 11698 193272 11704
rect 191840 3596 191892 3602
rect 191840 3538 191892 3544
rect 193232 480 193260 11698
rect 189326 354 189438 480
rect 189092 326 189438 354
rect 185462 -960 185574 326
rect 189326 -960 189438 326
rect 193190 -960 193302 480
rect 196636 354 196664 16546
rect 197054 354 197166 480
rect 196636 326 197166 354
rect 200500 354 200528 16546
rect 204352 14612 204404 14618
rect 204352 14554 204404 14560
rect 200918 354 201030 480
rect 200500 326 201030 354
rect 204364 354 204392 14554
rect 207676 3602 207704 28222
rect 210424 24132 210476 24138
rect 210424 24074 210476 24080
rect 210436 3602 210464 24074
rect 207664 3596 207716 3602
rect 207664 3538 207716 3544
rect 208676 3596 208728 3602
rect 208676 3538 208728 3544
rect 210424 3596 210476 3602
rect 210424 3538 210476 3544
rect 208688 480 208716 3538
rect 211264 3534 211292 143006
rect 211356 66162 211384 183126
rect 211448 80782 211476 198018
rect 211618 195256 211674 195265
rect 211618 195191 211674 195200
rect 211528 178968 211580 178974
rect 211528 178910 211580 178916
rect 211436 80776 211488 80782
rect 211436 80718 211488 80724
rect 211344 66156 211396 66162
rect 211344 66098 211396 66104
rect 211540 63510 211568 178910
rect 211632 79121 211660 195191
rect 211712 185836 211764 185842
rect 211712 185778 211764 185784
rect 211618 79112 211674 79121
rect 211618 79047 211674 79056
rect 211724 78402 211752 185778
rect 211896 181416 211948 181422
rect 211896 181358 211948 181364
rect 211804 140888 211856 140894
rect 211804 140830 211856 140836
rect 211712 78396 211764 78402
rect 211712 78338 211764 78344
rect 211528 63504 211580 63510
rect 211528 63446 211580 63452
rect 211816 3534 211844 140830
rect 211908 76906 211936 181358
rect 211988 148368 212040 148374
rect 211988 148310 212040 148316
rect 211896 76900 211948 76906
rect 211896 76842 211948 76848
rect 212000 67454 212028 148310
rect 211988 67448 212040 67454
rect 211988 67390 212040 67396
rect 212552 64734 212580 198086
rect 213920 196784 213972 196790
rect 213920 196726 213972 196732
rect 212724 193928 212776 193934
rect 212724 193870 212776 193876
rect 212632 183320 212684 183326
rect 212632 183262 212684 183268
rect 212540 64728 212592 64734
rect 212540 64670 212592 64676
rect 212644 63442 212672 183262
rect 212736 78810 212764 193870
rect 212816 185768 212868 185774
rect 212816 185710 212868 185716
rect 212828 79082 212856 185710
rect 213000 180192 213052 180198
rect 213000 180134 213052 180140
rect 212906 178800 212962 178809
rect 212906 178735 212962 178744
rect 212816 79076 212868 79082
rect 212816 79018 212868 79024
rect 212724 78804 212776 78810
rect 212724 78746 212776 78752
rect 212920 75585 212948 178735
rect 213012 80889 213040 180134
rect 213092 142996 213144 143002
rect 213092 142938 213144 142944
rect 212998 80880 213054 80889
rect 212998 80815 213054 80824
rect 212906 75576 212962 75585
rect 212906 75511 212962 75520
rect 212632 63436 212684 63442
rect 212632 63378 212684 63384
rect 213104 62966 213132 142938
rect 213184 141568 213236 141574
rect 213184 141510 213236 141516
rect 213196 63034 213224 141510
rect 213932 64666 213960 196726
rect 214012 196716 214064 196722
rect 214012 196658 214064 196664
rect 214024 64841 214052 196658
rect 214116 78538 214144 200330
rect 218428 199708 218480 199714
rect 218428 199650 218480 199656
rect 217230 199608 217286 199617
rect 217230 199543 217286 199552
rect 216678 199472 216734 199481
rect 216678 199407 216734 199416
rect 214196 196852 214248 196858
rect 214196 196794 214248 196800
rect 214104 78532 214156 78538
rect 214104 78474 214156 78480
rect 214208 75614 214236 196794
rect 215298 195800 215354 195809
rect 215298 195735 215354 195744
rect 214654 195664 214710 195673
rect 214654 195599 214710 195608
rect 214288 195492 214340 195498
rect 214288 195434 214340 195440
rect 214300 75750 214328 195434
rect 214470 195392 214526 195401
rect 214470 195327 214526 195336
rect 214564 195356 214616 195362
rect 214380 195288 214432 195294
rect 214380 195230 214432 195236
rect 214288 75744 214340 75750
rect 214288 75686 214340 75692
rect 214196 75608 214248 75614
rect 214196 75550 214248 75556
rect 214392 75070 214420 195230
rect 214484 76537 214512 195327
rect 214564 195298 214616 195304
rect 214470 76528 214526 76537
rect 214470 76463 214526 76472
rect 214576 76430 214604 195298
rect 214668 79490 214696 195599
rect 215312 195537 215340 195735
rect 215298 195528 215354 195537
rect 215298 195463 215354 195472
rect 215482 195528 215538 195537
rect 215482 195463 215538 195472
rect 215298 192808 215354 192817
rect 215298 192743 215354 192752
rect 214748 178696 214800 178702
rect 214748 178638 214800 178644
rect 214656 79484 214708 79490
rect 214656 79426 214708 79432
rect 214760 77353 214788 178638
rect 214746 77344 214802 77353
rect 214746 77279 214802 77288
rect 214564 76424 214616 76430
rect 214564 76366 214616 76372
rect 214380 75064 214432 75070
rect 214380 75006 214432 75012
rect 214010 64832 214066 64841
rect 214010 64767 214066 64776
rect 215312 64705 215340 192743
rect 215390 189544 215446 189553
rect 215390 189479 215446 189488
rect 215404 74390 215432 189479
rect 215496 79218 215524 195463
rect 215574 192672 215630 192681
rect 215574 192607 215630 192616
rect 215484 79212 215536 79218
rect 215484 79154 215536 79160
rect 215588 76265 215616 192607
rect 215666 190360 215722 190369
rect 215666 190295 215722 190304
rect 215680 80034 215708 190295
rect 215760 188488 215812 188494
rect 215760 188430 215812 188436
rect 215668 80028 215720 80034
rect 215668 79970 215720 79976
rect 215772 79150 215800 188430
rect 215852 178900 215904 178906
rect 215852 178842 215904 178848
rect 215760 79144 215812 79150
rect 215760 79086 215812 79092
rect 215574 76256 215630 76265
rect 215574 76191 215630 76200
rect 215392 74384 215444 74390
rect 215392 74326 215444 74332
rect 215404 73846 215432 74326
rect 215392 73840 215444 73846
rect 215392 73782 215444 73788
rect 215864 71670 215892 178842
rect 216036 146940 216088 146946
rect 216036 146882 216088 146888
rect 216048 146402 216076 146882
rect 215944 146396 215996 146402
rect 215944 146338 215996 146344
rect 216036 146396 216088 146402
rect 216036 146338 216088 146344
rect 215852 71664 215904 71670
rect 215852 71606 215904 71612
rect 215864 71058 215892 71606
rect 215852 71052 215904 71058
rect 215852 70994 215904 71000
rect 215956 64802 215984 146338
rect 216048 66774 216076 146338
rect 216128 133204 216180 133210
rect 216128 133146 216180 133152
rect 216140 132530 216168 133146
rect 216128 132524 216180 132530
rect 216128 132466 216180 132472
rect 216140 75138 216168 132466
rect 216128 75132 216180 75138
rect 216128 75074 216180 75080
rect 216692 74905 216720 199407
rect 217244 198801 217272 199543
rect 218440 198830 218468 199650
rect 218060 198824 218112 198830
rect 217046 198792 217102 198801
rect 217046 198727 217102 198736
rect 217230 198792 217286 198801
rect 218060 198766 218112 198772
rect 218428 198824 218480 198830
rect 218428 198766 218480 198772
rect 217230 198727 217286 198736
rect 216864 191344 216916 191350
rect 216864 191286 216916 191292
rect 216876 191146 216904 191286
rect 216864 191140 216916 191146
rect 216864 191082 216916 191088
rect 216770 183016 216826 183025
rect 216770 182951 216826 182960
rect 216678 74896 216734 74905
rect 216678 74831 216734 74840
rect 216036 66768 216088 66774
rect 216036 66710 216088 66716
rect 216784 66065 216812 182951
rect 216876 74458 216904 191082
rect 216956 188420 217008 188426
rect 216956 188362 217008 188368
rect 216864 74452 216916 74458
rect 216864 74394 216916 74400
rect 216968 71505 216996 188362
rect 217060 82249 217088 198727
rect 217138 193896 217194 193905
rect 217138 193831 217194 193840
rect 217046 82240 217102 82249
rect 217046 82175 217102 82184
rect 217152 78878 217180 193831
rect 217232 189916 217284 189922
rect 217232 189858 217284 189864
rect 217140 78872 217192 78878
rect 217140 78814 217192 78820
rect 217244 76498 217272 189858
rect 217416 181892 217468 181898
rect 217416 181834 217468 181840
rect 217324 178832 217376 178838
rect 217324 178774 217376 178780
rect 217232 76492 217284 76498
rect 217232 76434 217284 76440
rect 217336 75886 217364 178774
rect 217428 82113 217456 181834
rect 217414 82104 217470 82113
rect 217414 82039 217470 82048
rect 217324 75880 217376 75886
rect 217324 75822 217376 75828
rect 218072 73250 218100 198766
rect 218242 196888 218298 196897
rect 218242 196823 218298 196832
rect 218152 185768 218204 185774
rect 218152 185710 218204 185716
rect 218164 185638 218192 185710
rect 218152 185632 218204 185638
rect 218152 185574 218204 185580
rect 218152 185496 218204 185502
rect 218152 185438 218204 185444
rect 218164 74534 218192 185438
rect 218256 78985 218284 196823
rect 219622 191448 219678 191457
rect 219622 191383 219678 191392
rect 218428 188352 218480 188358
rect 218428 188294 218480 188300
rect 218336 185768 218388 185774
rect 218336 185710 218388 185716
rect 218242 78976 218298 78985
rect 218242 78911 218298 78920
rect 218164 74506 218284 74534
rect 218072 73222 218192 73250
rect 218060 73160 218112 73166
rect 218060 73102 218112 73108
rect 218072 72418 218100 73102
rect 218060 72412 218112 72418
rect 218060 72354 218112 72360
rect 216954 71496 217010 71505
rect 216954 71431 217010 71440
rect 218164 68921 218192 73222
rect 218150 68912 218206 68921
rect 218150 68847 218206 68856
rect 218256 66201 218284 74506
rect 218348 71777 218376 185710
rect 218440 185502 218468 188294
rect 218428 185496 218480 185502
rect 218428 185438 218480 185444
rect 218426 184512 218482 184521
rect 218426 184447 218482 184456
rect 218440 78849 218468 184447
rect 219530 183560 219586 183569
rect 219530 183495 219586 183504
rect 219438 181656 219494 181665
rect 219438 181591 219494 181600
rect 218612 151088 218664 151094
rect 218612 151030 218664 151036
rect 218520 141500 218572 141506
rect 218520 141442 218572 141448
rect 218426 78840 218482 78849
rect 218426 78775 218482 78784
rect 218334 71768 218390 71777
rect 218334 71703 218390 71712
rect 218242 66192 218298 66201
rect 218242 66127 218298 66136
rect 216770 66056 216826 66065
rect 216770 65991 216826 66000
rect 215944 64796 215996 64802
rect 215944 64738 215996 64744
rect 215298 64696 215354 64705
rect 213920 64660 213972 64666
rect 215298 64631 215354 64640
rect 213920 64602 213972 64608
rect 213184 63028 213236 63034
rect 213184 62970 213236 62976
rect 213092 62960 213144 62966
rect 213092 62902 213144 62908
rect 215300 58812 215352 58818
rect 215300 58754 215352 58760
rect 215312 16574 215340 58754
rect 218532 57934 218560 141442
rect 218624 73166 218652 151030
rect 218612 73160 218664 73166
rect 218612 73102 218664 73108
rect 219452 67561 219480 181591
rect 219544 71641 219572 183495
rect 219636 79014 219664 191383
rect 220832 190913 220860 683086
rect 221004 200864 221056 200870
rect 221004 200806 221056 200812
rect 221016 200258 221044 200806
rect 221004 200252 221056 200258
rect 221004 200194 221056 200200
rect 220818 190904 220874 190913
rect 220818 190839 220874 190848
rect 221016 190454 221044 200194
rect 220924 190426 221044 190454
rect 220174 183560 220230 183569
rect 220174 183495 220230 183504
rect 219806 183288 219862 183297
rect 219806 183223 219862 183232
rect 219714 181384 219770 181393
rect 219714 181319 219770 181328
rect 219624 79008 219676 79014
rect 219624 78950 219676 78956
rect 219728 71738 219756 181319
rect 219820 75721 219848 183223
rect 220188 183025 220216 183495
rect 220174 183016 220230 183025
rect 220174 182951 220230 182960
rect 220820 181620 220872 181626
rect 220820 181562 220872 181568
rect 219992 181552 220044 181558
rect 219992 181494 220044 181500
rect 220082 181520 220138 181529
rect 219900 180124 219952 180130
rect 219900 180066 219952 180072
rect 219912 78674 219940 180066
rect 220004 80918 220032 181494
rect 220082 181455 220138 181464
rect 219992 80912 220044 80918
rect 219992 80854 220044 80860
rect 220096 80753 220124 181455
rect 220082 80744 220138 80753
rect 220082 80679 220138 80688
rect 219900 78668 219952 78674
rect 219900 78610 219952 78616
rect 219806 75712 219862 75721
rect 219806 75647 219862 75656
rect 219716 71732 219768 71738
rect 219716 71674 219768 71680
rect 219530 71632 219586 71641
rect 219530 71567 219586 71576
rect 219438 67552 219494 67561
rect 219438 67487 219494 67496
rect 218060 57928 218112 57934
rect 218060 57870 218112 57876
rect 218520 57928 218572 57934
rect 218520 57870 218572 57876
rect 218072 57254 218100 57870
rect 218060 57248 218112 57254
rect 218060 57190 218112 57196
rect 220832 48278 220860 181562
rect 220924 77081 220952 190426
rect 221004 185632 221056 185638
rect 221004 185574 221056 185580
rect 220910 77072 220966 77081
rect 220910 77007 220966 77016
rect 221016 66230 221044 185574
rect 227732 183190 227760 702406
rect 231872 191729 231900 702406
rect 231858 191720 231914 191729
rect 231858 191655 231914 191664
rect 227720 183184 227772 183190
rect 227720 183126 227772 183132
rect 221096 182980 221148 182986
rect 221096 182922 221148 182928
rect 221004 66224 221056 66230
rect 221004 66166 221056 66172
rect 221108 65929 221136 182922
rect 236012 179081 236040 702406
rect 239404 700324 239456 700330
rect 239404 700266 239456 700272
rect 239416 199617 239444 700266
rect 240244 683114 240272 703520
rect 244108 700398 244136 703520
rect 247972 702434 248000 703520
rect 251836 702434 251864 703520
rect 247052 702406 248000 702434
rect 251192 702406 251864 702434
rect 244096 700392 244148 700398
rect 244096 700334 244148 700340
rect 240152 683086 240272 683114
rect 239402 199608 239458 199617
rect 239402 199543 239458 199552
rect 240152 185774 240180 683086
rect 240140 185768 240192 185774
rect 240140 185710 240192 185716
rect 247052 183122 247080 702406
rect 251192 188766 251220 702406
rect 251180 188760 251232 188766
rect 251180 188702 251232 188708
rect 247040 183116 247092 183122
rect 247040 183058 247092 183064
rect 253952 181966 253980 703582
rect 254872 703474 254900 703582
rect 255014 703520 255126 704960
rect 258878 703520 258990 704960
rect 262742 703520 262854 704960
rect 266606 703520 266718 704960
rect 270470 703520 270582 704960
rect 273272 703582 274220 703610
rect 255056 703474 255084 703520
rect 254872 703446 255084 703474
rect 262784 699718 262812 703520
rect 266648 702434 266676 703520
rect 266372 702406 266676 702434
rect 260104 699712 260156 699718
rect 260104 699654 260156 699660
rect 262772 699712 262824 699718
rect 262772 699654 262824 699660
rect 260116 190369 260144 699654
rect 260102 190360 260158 190369
rect 260102 190295 260158 190304
rect 266372 190233 266400 702406
rect 266358 190224 266414 190233
rect 266358 190159 266414 190168
rect 273272 186182 273300 703582
rect 274192 703474 274220 703582
rect 274334 703520 274446 704960
rect 277412 703582 278084 703610
rect 274376 703474 274404 703520
rect 274192 703446 274404 703474
rect 273260 186176 273312 186182
rect 273260 186118 273312 186124
rect 277412 182034 277440 703582
rect 278056 703474 278084 703582
rect 278198 703520 278310 704960
rect 281552 703582 281948 703610
rect 278240 703474 278268 703520
rect 278056 703446 278268 703474
rect 281552 193118 281580 703582
rect 281920 703474 281948 703582
rect 282062 703520 282174 704960
rect 285926 703520 286038 704960
rect 289146 703520 289258 704960
rect 293010 703520 293122 704960
rect 296874 703520 296986 704960
rect 300738 703520 300850 704960
rect 304602 703520 304714 704960
rect 308466 703520 308578 704960
rect 312330 703520 312442 704960
rect 316194 703520 316306 704960
rect 320058 703520 320170 704960
rect 323922 703520 324034 704960
rect 327142 703520 327254 704960
rect 331006 703520 331118 704960
rect 333992 703582 334756 703610
rect 282104 703474 282132 703520
rect 281920 703446 282132 703474
rect 285968 702434 285996 703520
rect 289188 702434 289216 703520
rect 293052 702434 293080 703520
rect 285692 702406 285996 702434
rect 288452 702406 289216 702434
rect 292592 702406 293080 702434
rect 285692 263090 285720 702406
rect 288452 269890 288480 702406
rect 288440 269884 288492 269890
rect 288440 269826 288492 269832
rect 285680 263084 285732 263090
rect 285680 263026 285732 263032
rect 281540 193112 281592 193118
rect 281540 193054 281592 193060
rect 277400 182028 277452 182034
rect 277400 181970 277452 181976
rect 253940 181960 253992 181966
rect 253940 181902 253992 181908
rect 292592 181490 292620 702406
rect 300780 696658 300808 703520
rect 304644 702434 304672 703520
rect 303632 702406 304672 702434
rect 299480 696652 299532 696658
rect 299480 696594 299532 696600
rect 300768 696652 300820 696658
rect 300768 696594 300820 696600
rect 299492 181558 299520 696594
rect 303632 199782 303660 702406
rect 308508 699718 308536 703520
rect 312372 699718 312400 703520
rect 316236 699718 316264 703520
rect 323964 702434 323992 703520
rect 322952 702406 323992 702434
rect 305644 699712 305696 699718
rect 305644 699654 305696 699660
rect 308496 699712 308548 699718
rect 308496 699654 308548 699660
rect 309784 699712 309836 699718
rect 309784 699654 309836 699660
rect 312360 699712 312412 699718
rect 312360 699654 312412 699660
rect 313924 699712 313976 699718
rect 313924 699654 313976 699660
rect 316224 699712 316276 699718
rect 316224 699654 316276 699660
rect 303620 199776 303672 199782
rect 303620 199718 303672 199724
rect 299480 181552 299532 181558
rect 299480 181494 299532 181500
rect 292580 181484 292632 181490
rect 292580 181426 292632 181432
rect 305656 180441 305684 699654
rect 305642 180432 305698 180441
rect 305642 180367 305698 180376
rect 235998 179072 236054 179081
rect 235998 179007 236054 179016
rect 221186 178936 221242 178945
rect 221186 178871 221242 178880
rect 221094 65920 221150 65929
rect 221094 65855 221150 65864
rect 221200 63345 221228 178871
rect 309796 178770 309824 699654
rect 313936 187542 313964 699654
rect 313924 187536 313976 187542
rect 313924 187478 313976 187484
rect 322952 180402 322980 702406
rect 327184 683114 327212 703520
rect 331048 699718 331076 703520
rect 327724 699712 327776 699718
rect 327724 699654 327776 699660
rect 331036 699712 331088 699718
rect 331036 699654 331088 699660
rect 327092 683086 327212 683114
rect 327092 263022 327120 683086
rect 327080 263016 327132 263022
rect 327080 262958 327132 262964
rect 327736 195838 327764 699654
rect 333992 197169 334020 703582
rect 334728 703474 334756 703582
rect 334870 703520 334982 704960
rect 338734 703520 338846 704960
rect 342272 703582 342484 703610
rect 334912 703474 334940 703520
rect 334728 703446 334940 703474
rect 333978 197160 334034 197169
rect 333978 197095 334034 197104
rect 327724 195832 327776 195838
rect 327724 195774 327776 195780
rect 342272 192817 342300 703582
rect 342456 703474 342484 703582
rect 342598 703520 342710 704960
rect 346462 703520 346574 704960
rect 349172 703582 350212 703610
rect 342640 703474 342668 703520
rect 342456 703446 342668 703474
rect 342258 192808 342314 192817
rect 342258 192743 342314 192752
rect 349172 183054 349200 703582
rect 350184 703474 350212 703582
rect 350326 703520 350438 704960
rect 353312 703582 354076 703610
rect 350368 703474 350396 703520
rect 350184 703446 350396 703474
rect 349160 183048 349212 183054
rect 349160 182990 349212 182996
rect 322940 180396 322992 180402
rect 322940 180338 322992 180344
rect 309784 178764 309836 178770
rect 309784 178706 309836 178712
rect 221740 177404 221792 177410
rect 221740 177346 221792 177352
rect 221752 176730 221780 177346
rect 221280 176724 221332 176730
rect 221280 176666 221332 176672
rect 221740 176724 221792 176730
rect 221740 176666 221792 176672
rect 221292 73778 221320 176666
rect 353312 174962 353340 703582
rect 354048 703474 354076 703582
rect 354190 703520 354302 704960
rect 357452 703582 357940 703610
rect 354232 703474 354260 703520
rect 354048 703446 354260 703474
rect 357452 175030 357480 703582
rect 357912 703474 357940 703582
rect 358054 703520 358166 704960
rect 361918 703520 362030 704960
rect 365138 703520 365250 704960
rect 369002 703520 369114 704960
rect 372866 703520 372978 704960
rect 376730 703520 376842 704960
rect 380594 703520 380706 704960
rect 384458 703520 384570 704960
rect 388322 703520 388434 704960
rect 392186 703520 392298 704960
rect 396050 703520 396162 704960
rect 399914 703520 400026 704960
rect 403134 703520 403246 704960
rect 406998 703520 407110 704960
rect 409892 703582 410748 703610
rect 358096 703474 358124 703520
rect 357912 703446 358124 703474
rect 361960 699718 361988 703520
rect 365180 702434 365208 703520
rect 369044 702434 369072 703520
rect 364352 702406 365208 702434
rect 368492 702406 369072 702434
rect 359464 699712 359516 699718
rect 359464 699654 359516 699660
rect 361948 699712 362000 699718
rect 361948 699654 362000 699660
rect 359476 336054 359504 699654
rect 359464 336048 359516 336054
rect 359464 335990 359516 335996
rect 364352 177682 364380 702406
rect 364340 177676 364392 177682
rect 364340 177618 364392 177624
rect 368492 175098 368520 702406
rect 376772 195673 376800 703520
rect 380636 699718 380664 703520
rect 384500 699718 384528 703520
rect 392228 702434 392256 703520
rect 391952 702406 392256 702434
rect 377404 699712 377456 699718
rect 377404 699654 377456 699660
rect 380624 699712 380676 699718
rect 380624 699654 380676 699660
rect 381544 699712 381596 699718
rect 381544 699654 381596 699660
rect 384488 699712 384540 699718
rect 384488 699654 384540 699660
rect 376758 195664 376814 195673
rect 376758 195599 376814 195608
rect 377416 191457 377444 699654
rect 377402 191448 377458 191457
rect 377402 191383 377458 191392
rect 368480 175092 368532 175098
rect 368480 175034 368532 175040
rect 357440 175024 357492 175030
rect 381556 175001 381584 699654
rect 391952 194449 391980 702406
rect 396092 275330 396120 703520
rect 399956 702434 399984 703520
rect 398852 702406 399984 702434
rect 396080 275324 396132 275330
rect 396080 275266 396132 275272
rect 391938 194440 391994 194449
rect 391938 194375 391994 194384
rect 398852 191622 398880 702406
rect 403176 683114 403204 703520
rect 407040 703050 407068 703520
rect 405740 703044 405792 703050
rect 405740 702986 405792 702992
rect 407028 703044 407080 703050
rect 407028 702986 407080 702992
rect 402992 683086 403204 683114
rect 402992 199714 403020 683086
rect 402980 199708 403032 199714
rect 402980 199650 403032 199656
rect 398840 191616 398892 191622
rect 398840 191558 398892 191564
rect 405752 180470 405780 702986
rect 405740 180464 405792 180470
rect 405740 180406 405792 180412
rect 409892 177750 409920 703582
rect 410720 703474 410748 703582
rect 410862 703520 410974 704960
rect 414726 703520 414838 704960
rect 418172 703582 418476 703610
rect 410904 703474 410932 703520
rect 410720 703446 410932 703474
rect 418172 184890 418200 703582
rect 418448 703474 418476 703582
rect 418590 703520 418702 704960
rect 422454 703520 422566 704960
rect 426318 703520 426430 704960
rect 430182 703520 430294 704960
rect 434046 703520 434158 704960
rect 437266 703520 437378 704960
rect 441130 703520 441242 704960
rect 444994 703520 445106 704960
rect 448858 703520 448970 704960
rect 452722 703520 452834 704960
rect 456586 703520 456698 704960
rect 460450 703520 460562 704960
rect 464314 703520 464426 704960
rect 468178 703520 468290 704960
rect 472042 703520 472154 704960
rect 474752 703582 475148 703610
rect 418632 703474 418660 703520
rect 418448 703446 418660 703474
rect 422496 683114 422524 703520
rect 426360 703050 426388 703520
rect 425060 703044 425112 703050
rect 425060 702986 425112 702992
rect 426348 703044 426400 703050
rect 426348 702986 426400 702992
rect 422312 683086 422524 683114
rect 422312 200841 422340 683086
rect 422298 200832 422354 200841
rect 422298 200767 422354 200776
rect 418160 184884 418212 184890
rect 418160 184826 418212 184832
rect 425072 178702 425100 702986
rect 430224 699718 430252 703520
rect 434088 699718 434116 703520
rect 437308 703050 437336 703520
rect 436100 703044 436152 703050
rect 436100 702986 436152 702992
rect 437296 703044 437348 703050
rect 437296 702986 437348 702992
rect 428464 699712 428516 699718
rect 428464 699654 428516 699660
rect 430212 699712 430264 699718
rect 430212 699654 430264 699660
rect 431224 699712 431276 699718
rect 431224 699654 431276 699660
rect 434076 699712 434128 699718
rect 434076 699654 434128 699660
rect 428476 200734 428504 699654
rect 428464 200728 428516 200734
rect 428464 200670 428516 200676
rect 431236 190097 431264 699654
rect 431222 190088 431278 190097
rect 431222 190023 431278 190032
rect 436112 184657 436140 702986
rect 441172 702434 441200 703520
rect 445036 702434 445064 703520
rect 448900 702434 448928 703520
rect 440252 702406 441200 702434
rect 444392 702406 445064 702434
rect 448532 702406 448928 702434
rect 440252 267034 440280 702406
rect 440240 267028 440292 267034
rect 440240 266970 440292 266976
rect 444392 262954 444420 702406
rect 444380 262948 444432 262954
rect 444380 262890 444432 262896
rect 448532 199646 448560 702406
rect 452764 683114 452792 703520
rect 456628 703050 456656 703520
rect 455420 703044 455472 703050
rect 455420 702986 455472 702992
rect 456616 703044 456668 703050
rect 456616 702986 456668 702992
rect 452672 683086 452792 683114
rect 448520 199640 448572 199646
rect 448520 199582 448572 199588
rect 452672 186969 452700 683086
rect 455432 188737 455460 702986
rect 460492 702434 460520 703520
rect 464356 702434 464384 703520
rect 468220 702434 468248 703520
rect 459572 702406 460520 702434
rect 463712 702406 464384 702434
rect 467852 702406 468248 702434
rect 455418 188728 455474 188737
rect 455418 188663 455474 188672
rect 452658 186960 452714 186969
rect 452658 186895 452714 186904
rect 436098 184648 436154 184657
rect 436098 184583 436154 184592
rect 459572 178945 459600 702406
rect 459558 178936 459614 178945
rect 459558 178871 459614 178880
rect 463712 178809 463740 702406
rect 467852 262886 467880 702406
rect 472084 683114 472112 703520
rect 471992 683086 472112 683114
rect 467840 262880 467892 262886
rect 467840 262822 467892 262828
rect 471992 188018 472020 683086
rect 474752 200938 474780 703582
rect 475120 703474 475148 703582
rect 475262 703520 475374 704960
rect 479126 703520 479238 704960
rect 482990 703520 483102 704960
rect 485792 703582 486740 703610
rect 475304 703474 475332 703520
rect 475120 703446 475332 703474
rect 479168 699718 479196 703520
rect 476764 699712 476816 699718
rect 476764 699654 476816 699660
rect 479156 699712 479208 699718
rect 479156 699654 479208 699660
rect 474740 200932 474792 200938
rect 474740 200874 474792 200880
rect 471980 188012 472032 188018
rect 471980 187954 472032 187960
rect 463698 178800 463754 178809
rect 463698 178735 463754 178744
rect 425060 178696 425112 178702
rect 425060 178638 425112 178644
rect 409880 177744 409932 177750
rect 476776 177721 476804 699654
rect 483032 263129 483060 703520
rect 483018 263120 483074 263129
rect 483018 263055 483074 263064
rect 485792 183433 485820 703582
rect 486712 703474 486740 703582
rect 486854 703520 486966 704960
rect 489932 703582 490604 703610
rect 486896 703474 486924 703520
rect 486712 703446 486924 703474
rect 489932 187377 489960 703582
rect 490576 703474 490604 703582
rect 490718 703520 490830 704960
rect 494072 703582 494468 703610
rect 490760 703474 490788 703520
rect 490576 703446 490788 703474
rect 494072 191321 494100 703582
rect 494440 703474 494468 703582
rect 494582 703520 494694 704960
rect 498446 703520 498558 704960
rect 502310 703520 502422 704960
rect 506174 703520 506286 704960
rect 509252 703582 509924 703610
rect 494624 703474 494652 703520
rect 494440 703446 494652 703474
rect 498488 702434 498516 703520
rect 498212 702406 498516 702434
rect 494058 191312 494114 191321
rect 494058 191247 494114 191256
rect 490564 190528 490616 190534
rect 490564 190470 490616 190476
rect 489918 187368 489974 187377
rect 489918 187303 489974 187312
rect 485778 183424 485834 183433
rect 485778 183359 485834 183368
rect 409880 177686 409932 177692
rect 476762 177712 476818 177721
rect 476762 177647 476818 177656
rect 357440 174966 357492 174972
rect 381542 174992 381598 175001
rect 353300 174956 353352 174962
rect 381542 174927 381598 174936
rect 353300 174898 353352 174904
rect 490576 146266 490604 190470
rect 498212 180538 498240 702406
rect 502352 193866 502380 703520
rect 502340 193860 502392 193866
rect 502340 193802 502392 193808
rect 509252 191214 509280 703582
rect 509896 703474 509924 703582
rect 510038 703520 510150 704960
rect 513258 703520 513370 704960
rect 517122 703520 517234 704960
rect 520986 703520 521098 704960
rect 524850 703520 524962 704960
rect 528714 703520 528826 704960
rect 532578 703520 532690 704960
rect 536442 703520 536554 704960
rect 540306 703520 540418 704960
rect 544170 703520 544282 704960
rect 546512 703582 547276 703610
rect 510080 703474 510108 703520
rect 509896 703446 510108 703474
rect 513300 696658 513328 703520
rect 517164 702434 517192 703520
rect 521028 702434 521056 703520
rect 524892 702434 524920 703520
rect 516152 702406 517192 702434
rect 520292 702406 521056 702434
rect 524432 702406 524920 702434
rect 514024 700392 514076 700398
rect 514024 700334 514076 700340
rect 512000 696652 512052 696658
rect 512000 696594 512052 696600
rect 513288 696652 513340 696658
rect 513288 696594 513340 696600
rect 509240 191208 509292 191214
rect 509240 191150 509292 191156
rect 512012 184521 512040 696594
rect 514036 200705 514064 700334
rect 514022 200696 514078 200705
rect 514022 200631 514078 200640
rect 516152 199481 516180 702406
rect 516138 199472 516194 199481
rect 516138 199407 516194 199416
rect 520292 191146 520320 702406
rect 520280 191140 520332 191146
rect 520280 191082 520332 191088
rect 524432 188873 524460 702406
rect 528756 683114 528784 703520
rect 532620 697610 532648 703520
rect 536484 702434 536512 703520
rect 540348 702434 540376 703520
rect 544212 702434 544240 703520
rect 544384 702500 544436 702506
rect 544384 702442 544436 702448
rect 535472 702406 536512 702434
rect 539612 702406 540376 702434
rect 543752 702406 544240 702434
rect 531320 697604 531372 697610
rect 531320 697546 531372 697552
rect 532608 697604 532660 697610
rect 532608 697546 532660 697552
rect 528572 683086 528784 683114
rect 528572 199578 528600 683086
rect 531332 200870 531360 697546
rect 531320 200864 531372 200870
rect 531320 200806 531372 200812
rect 528560 199572 528612 199578
rect 528560 199514 528612 199520
rect 524418 188864 524474 188873
rect 524418 188799 524474 188808
rect 511998 184512 512054 184521
rect 511998 184447 512054 184456
rect 535472 181665 535500 702406
rect 539612 199510 539640 702406
rect 543004 700460 543056 700466
rect 543004 700402 543056 700408
rect 541624 661088 541676 661094
rect 541624 661030 541676 661036
rect 539600 199504 539652 199510
rect 539600 199446 539652 199452
rect 535458 181656 535514 181665
rect 535458 181591 535514 181600
rect 541636 180674 541664 661030
rect 541624 180668 541676 180674
rect 541624 180610 541676 180616
rect 498200 180532 498252 180538
rect 498200 180474 498252 180480
rect 543016 177993 543044 700402
rect 543752 183297 543780 702406
rect 544396 199345 544424 702442
rect 546512 262857 546540 703582
rect 547248 703474 547276 703582
rect 547390 703520 547502 704960
rect 551254 703520 551366 704960
rect 555118 703520 555230 704960
rect 558982 703520 559094 704960
rect 561692 703582 562732 703610
rect 547432 703474 547460 703520
rect 547248 703446 547460 703474
rect 551296 699718 551324 703520
rect 555160 700330 555188 703520
rect 555148 700324 555200 700330
rect 555148 700266 555200 700272
rect 559024 699718 559052 703520
rect 548524 699712 548576 699718
rect 548524 699654 548576 699660
rect 551284 699712 551336 699718
rect 551284 699654 551336 699660
rect 558184 699712 558236 699718
rect 558184 699654 558236 699660
rect 559012 699712 559064 699718
rect 559012 699654 559064 699660
rect 546498 262848 546554 262857
rect 546498 262783 546554 262792
rect 544382 199336 544438 199345
rect 544382 199271 544438 199280
rect 544384 192568 544436 192574
rect 544384 192510 544436 192516
rect 543738 183288 543794 183297
rect 543738 183223 543794 183232
rect 543002 177984 543058 177993
rect 543002 177919 543058 177928
rect 490564 146260 490616 146266
rect 490564 146202 490616 146208
rect 329840 142860 329892 142866
rect 329840 142802 329892 142808
rect 288440 139528 288492 139534
rect 288440 139470 288492 139476
rect 269120 75200 269172 75206
rect 269120 75142 269172 75148
rect 221280 73772 221332 73778
rect 221280 73714 221332 73720
rect 253940 72480 253992 72486
rect 253940 72422 253992 72428
rect 221186 63336 221242 63345
rect 221186 63271 221242 63280
rect 234620 54596 234672 54602
rect 234620 54538 234672 54544
rect 220820 48272 220872 48278
rect 220820 48214 220872 48220
rect 222108 48272 222160 48278
rect 222108 48214 222160 48220
rect 222120 47598 222148 48214
rect 222108 47592 222160 47598
rect 222108 47534 222160 47540
rect 230480 46300 230532 46306
rect 230480 46242 230532 46248
rect 219440 36576 219492 36582
rect 219440 36518 219492 36524
rect 219452 16574 219480 36518
rect 226340 18692 226392 18698
rect 226340 18634 226392 18640
rect 226352 16574 226380 18634
rect 230492 16574 230520 46242
rect 234632 16574 234660 54538
rect 245660 39432 245712 39438
rect 245660 39374 245712 39380
rect 245672 16574 245700 39374
rect 249800 26988 249852 26994
rect 249800 26930 249852 26936
rect 249812 16574 249840 26930
rect 253952 16574 253980 72422
rect 260840 65612 260892 65618
rect 260840 65554 260892 65560
rect 256700 57316 256752 57322
rect 256700 57258 256752 57264
rect 256712 16574 256740 57258
rect 260852 16574 260880 65554
rect 264980 64252 265032 64258
rect 264980 64194 265032 64200
rect 215312 16546 215984 16574
rect 219452 16546 219848 16574
rect 226352 16546 227392 16574
rect 230492 16546 231256 16574
rect 234632 16546 235120 16574
rect 245672 16546 246712 16574
rect 249812 16546 250576 16574
rect 253952 16546 254440 16574
rect 256712 16546 257200 16574
rect 260852 16546 261064 16574
rect 211252 3528 211304 3534
rect 211252 3470 211304 3476
rect 211804 3528 211856 3534
rect 211804 3470 211856 3476
rect 212540 3528 212592 3534
rect 212540 3470 212592 3476
rect 212552 480 212580 3470
rect 204782 354 204894 480
rect 204364 326 204894 354
rect 197054 -960 197166 326
rect 200918 -960 201030 326
rect 204782 -960 204894 326
rect 208646 -960 208758 480
rect 212510 -960 212622 480
rect 215956 354 215984 16546
rect 216374 354 216486 480
rect 215956 326 216486 354
rect 219820 354 219848 16546
rect 227364 480 227392 16546
rect 231228 480 231256 16546
rect 235092 480 235120 16546
rect 241704 8968 241756 8974
rect 241704 8910 241756 8916
rect 241716 3534 241744 8910
rect 242808 3596 242860 3602
rect 242808 3538 242860 3544
rect 241704 3528 241756 3534
rect 241704 3470 241756 3476
rect 242820 480 242848 3538
rect 246684 480 246712 16546
rect 250548 480 250576 16546
rect 254412 480 254440 16546
rect 220238 354 220350 480
rect 219820 326 220350 354
rect 216374 -960 216486 326
rect 220238 -960 220350 326
rect 223458 -960 223570 480
rect 227322 -960 227434 480
rect 231186 -960 231298 480
rect 235050 -960 235162 480
rect 238914 -960 239026 480
rect 242778 -960 242890 480
rect 246642 -960 246754 480
rect 250506 -960 250618 480
rect 254370 -960 254482 480
rect 257172 354 257200 16546
rect 257590 354 257702 480
rect 257172 326 257702 354
rect 261036 354 261064 16546
rect 261454 354 261566 480
rect 261036 326 261566 354
rect 264992 354 265020 64194
rect 269132 16574 269160 75142
rect 276020 53168 276072 53174
rect 276020 53110 276072 53116
rect 276032 16574 276060 53110
rect 284300 47660 284352 47666
rect 284300 47602 284352 47608
rect 269132 16546 269252 16574
rect 276032 16546 276520 16574
rect 269224 480 269252 16546
rect 265318 354 265430 480
rect 264992 326 265430 354
rect 257590 -960 257702 326
rect 261454 -960 261566 326
rect 265318 -960 265430 326
rect 269182 -960 269294 480
rect 273046 -960 273158 480
rect 276492 354 276520 16546
rect 280804 4820 280856 4826
rect 280804 4762 280856 4768
rect 280816 480 280844 4762
rect 276910 354 277022 480
rect 276492 326 277022 354
rect 276910 -960 277022 326
rect 280774 -960 280886 480
rect 284312 354 284340 47602
rect 288452 16574 288480 139470
rect 321560 73908 321612 73914
rect 321560 73850 321612 73856
rect 306380 71120 306432 71126
rect 306380 71062 306432 71068
rect 302240 62892 302292 62898
rect 302240 62834 302292 62840
rect 295340 61464 295392 61470
rect 295340 61406 295392 61412
rect 295352 16574 295380 61406
rect 302252 16574 302280 62834
rect 306392 16574 306420 71062
rect 314660 69692 314712 69698
rect 314660 69634 314712 69640
rect 310520 68400 310572 68406
rect 310520 68342 310572 68348
rect 310532 16574 310560 68342
rect 314672 16574 314700 69634
rect 321572 16574 321600 73850
rect 329852 16574 329880 142802
rect 518900 142316 518952 142322
rect 518900 142258 518952 142264
rect 492680 140072 492732 140078
rect 492680 140014 492732 140020
rect 416780 137284 416832 137290
rect 416780 137226 416832 137232
rect 386420 66972 386472 66978
rect 386420 66914 386472 66920
rect 345020 55888 345072 55894
rect 345020 55830 345072 55836
rect 340880 39364 340932 39370
rect 340880 39306 340932 39312
rect 332600 29708 332652 29714
rect 332600 29650 332652 29656
rect 332612 16574 332640 29650
rect 288452 16546 288572 16574
rect 295352 16546 295656 16574
rect 302252 16546 303384 16574
rect 306392 16546 307248 16574
rect 310532 16546 311112 16574
rect 314672 16546 314976 16574
rect 321572 16546 322704 16574
rect 329852 16546 330432 16574
rect 332612 16546 333192 16574
rect 288544 480 288572 16546
rect 295628 480 295656 16546
rect 299480 10396 299532 10402
rect 299480 10338 299532 10344
rect 299492 480 299520 10338
rect 303356 480 303384 16546
rect 307220 480 307248 16546
rect 311084 480 311112 16546
rect 314948 480 314976 16546
rect 318800 7676 318852 7682
rect 318800 7618 318852 7624
rect 318812 480 318840 7618
rect 322676 480 322704 16546
rect 326528 3528 326580 3534
rect 326528 3470 326580 3476
rect 326540 480 326568 3470
rect 330404 480 330432 16546
rect 284638 354 284750 480
rect 284312 326 284750 354
rect 284638 -960 284750 326
rect 288502 -960 288614 480
rect 292366 -960 292478 480
rect 295586 -960 295698 480
rect 299450 -960 299562 480
rect 303314 -960 303426 480
rect 307178 -960 307290 480
rect 311042 -960 311154 480
rect 314906 -960 315018 480
rect 318770 -960 318882 480
rect 322634 -960 322746 480
rect 326498 -960 326610 480
rect 330362 -960 330474 480
rect 333164 354 333192 16546
rect 333582 354 333694 480
rect 333164 326 333694 354
rect 333582 -960 333694 326
rect 337446 -960 337558 480
rect 340892 354 340920 39306
rect 341310 354 341422 480
rect 340892 326 341422 354
rect 345032 354 345060 55830
rect 374644 49020 374696 49026
rect 374644 48962 374696 48968
rect 371240 35284 371292 35290
rect 371240 35226 371292 35232
rect 356060 33788 356112 33794
rect 356060 33730 356112 33736
rect 347780 26920 347832 26926
rect 347780 26862 347832 26868
rect 347792 16574 347820 26862
rect 356072 16574 356100 33730
rect 364340 31136 364392 31142
rect 364340 31078 364392 31084
rect 347792 16546 348648 16574
rect 356072 16546 356376 16574
rect 345174 354 345286 480
rect 345032 326 345286 354
rect 348620 354 348648 16546
rect 352472 14544 352524 14550
rect 352472 14486 352524 14492
rect 349038 354 349150 480
rect 348620 326 349150 354
rect 352484 354 352512 14486
rect 352902 354 353014 480
rect 352484 326 353014 354
rect 356348 354 356376 16546
rect 360660 7608 360712 7614
rect 360660 7550 360712 7556
rect 360672 480 360700 7550
rect 356766 354 356878 480
rect 356348 326 356878 354
rect 341310 -960 341422 326
rect 345174 -960 345286 326
rect 349038 -960 349150 326
rect 352902 -960 353014 326
rect 356766 -960 356878 326
rect 360630 -960 360742 480
rect 364352 354 364380 31078
rect 371252 16574 371280 35226
rect 371252 16546 371648 16574
rect 371620 480 371648 16546
rect 374656 3534 374684 48962
rect 377404 42152 377456 42158
rect 377404 42094 377456 42100
rect 377416 3602 377444 42094
rect 378140 38004 378192 38010
rect 378140 37946 378192 37952
rect 377404 3596 377456 3602
rect 377404 3538 377456 3544
rect 378152 3534 378180 37946
rect 386432 16574 386460 66914
rect 408500 65544 408552 65550
rect 408500 65486 408552 65492
rect 400864 50448 400916 50454
rect 400864 50390 400916 50396
rect 394700 43512 394752 43518
rect 394700 43454 394752 43460
rect 390560 40724 390612 40730
rect 390560 40666 390612 40672
rect 390572 16574 390600 40666
rect 394712 16574 394740 43454
rect 386432 16546 387104 16574
rect 390572 16546 390968 16574
rect 394712 16546 394832 16574
rect 374644 3528 374696 3534
rect 374644 3470 374696 3476
rect 375472 3528 375524 3534
rect 375472 3470 375524 3476
rect 378140 3528 378192 3534
rect 378140 3470 378192 3476
rect 379336 3528 379388 3534
rect 379336 3470 379388 3476
rect 375484 480 375512 3470
rect 379348 480 379376 3470
rect 383200 3460 383252 3466
rect 383200 3402 383252 3408
rect 383212 480 383240 3402
rect 387076 480 387104 16546
rect 390940 480 390968 16546
rect 394804 480 394832 16546
rect 398656 6248 398708 6254
rect 398656 6190 398708 6196
rect 398668 480 398696 6190
rect 400876 3466 400904 50390
rect 408512 16574 408540 65486
rect 416792 16574 416820 137226
rect 484400 71052 484452 71058
rect 484400 70994 484452 71000
rect 462320 68332 462372 68338
rect 462320 68274 462372 68280
rect 425060 62824 425112 62830
rect 425060 62766 425112 62772
rect 420920 47592 420972 47598
rect 420920 47534 420972 47540
rect 408512 16546 409184 16574
rect 416792 16546 416912 16574
rect 400864 3460 400916 3466
rect 400864 3402 400916 3408
rect 402520 3460 402572 3466
rect 402520 3402 402572 3408
rect 402532 480 402560 3402
rect 364494 354 364606 480
rect 364352 326 364606 354
rect 364494 -960 364606 326
rect 367714 -960 367826 480
rect 371578 -960 371690 480
rect 375442 -960 375554 480
rect 379306 -960 379418 480
rect 383170 -960 383282 480
rect 387034 -960 387146 480
rect 390898 -960 391010 480
rect 394762 -960 394874 480
rect 398626 -960 398738 480
rect 402490 -960 402602 480
rect 405710 -960 405822 480
rect 409156 354 409184 16546
rect 409574 354 409686 480
rect 409156 326 409686 354
rect 409574 -960 409686 326
rect 413438 -960 413550 480
rect 416884 354 416912 16546
rect 417302 354 417414 480
rect 416884 326 417414 354
rect 420932 354 420960 47534
rect 425072 480 425100 62766
rect 454040 60036 454092 60042
rect 454040 59978 454092 59984
rect 436100 44872 436152 44878
rect 436100 44814 436152 44820
rect 436112 16574 436140 44814
rect 442264 37936 442316 37942
rect 442264 37878 442316 37884
rect 436112 16546 436232 16574
rect 432788 6180 432840 6186
rect 432788 6122 432840 6128
rect 432800 480 432828 6122
rect 421166 354 421278 480
rect 420932 326 421278 354
rect 417302 -960 417414 326
rect 421166 -960 421278 326
rect 425030 -960 425142 480
rect 428894 -960 429006 480
rect 432758 -960 432870 480
rect 436204 354 436232 16546
rect 442276 3466 442304 37878
rect 447600 13184 447652 13190
rect 447600 13126 447652 13132
rect 442264 3460 442316 3466
rect 442264 3402 442316 3408
rect 443736 3460 443788 3466
rect 443736 3402 443788 3408
rect 443748 480 443776 3402
rect 447612 480 447640 13126
rect 454052 3466 454080 59978
rect 462332 16574 462360 68274
rect 477500 64184 477552 64190
rect 477500 64126 477552 64132
rect 470600 57248 470652 57254
rect 470600 57190 470652 57196
rect 466460 21412 466512 21418
rect 466460 21354 466512 21360
rect 466472 16574 466500 21354
rect 470612 16574 470640 57190
rect 473360 25560 473412 25566
rect 473360 25502 473412 25508
rect 462332 16546 463096 16574
rect 466472 16546 466960 16574
rect 470612 16546 470824 16574
rect 459192 14476 459244 14482
rect 459192 14418 459244 14424
rect 454040 3460 454092 3466
rect 454040 3402 454092 3408
rect 455328 3460 455380 3466
rect 455328 3402 455380 3408
rect 455340 480 455368 3402
rect 459204 480 459232 14418
rect 463068 480 463096 16546
rect 466932 480 466960 16546
rect 470796 480 470824 16546
rect 473372 3466 473400 25502
rect 473360 3460 473412 3466
rect 473360 3402 473412 3408
rect 474648 3460 474700 3466
rect 474648 3402 474700 3408
rect 474660 480 474688 3402
rect 436622 354 436734 480
rect 436204 326 436734 354
rect 436622 -960 436734 326
rect 440486 -960 440598 480
rect 443706 -960 443818 480
rect 447570 -960 447682 480
rect 451434 -960 451546 480
rect 455298 -960 455410 480
rect 459162 -960 459274 480
rect 463026 -960 463138 480
rect 466890 -960 467002 480
rect 470754 -960 470866 480
rect 474618 -960 474730 480
rect 477512 354 477540 64126
rect 481640 18624 481692 18630
rect 481640 18566 481692 18572
rect 481652 16574 481680 18566
rect 484412 16574 484440 70994
rect 488540 66904 488592 66910
rect 488540 66846 488592 66852
rect 488552 16574 488580 66846
rect 492692 16574 492720 140014
rect 512000 138712 512052 138718
rect 512000 138654 512052 138660
rect 496084 61396 496136 61402
rect 496084 61338 496136 61344
rect 481652 16546 481772 16574
rect 484412 16546 485176 16574
rect 488552 16546 489040 16574
rect 492692 16546 492904 16574
rect 481744 480 481772 16546
rect 477838 354 477950 480
rect 477512 326 477950 354
rect 477838 -960 477950 326
rect 481702 -960 481814 480
rect 485148 354 485176 16546
rect 485566 354 485678 480
rect 485148 326 485678 354
rect 489012 354 489040 16546
rect 489430 354 489542 480
rect 489012 326 489542 354
rect 492876 354 492904 16546
rect 496096 3466 496124 61338
rect 502984 51740 503036 51746
rect 502984 51682 503036 51688
rect 500224 29640 500276 29646
rect 500224 29582 500276 29588
rect 496084 3460 496136 3466
rect 496084 3402 496136 3408
rect 497188 3460 497240 3466
rect 497188 3402 497240 3408
rect 497200 480 497228 3402
rect 500236 2922 500264 29582
rect 502996 3466 503024 51682
rect 503720 42084 503772 42090
rect 503720 42026 503772 42032
rect 503732 16574 503760 42026
rect 512012 16574 512040 138654
rect 514024 22772 514076 22778
rect 514024 22714 514076 22720
rect 503732 16546 504496 16574
rect 512012 16546 512224 16574
rect 502984 3460 503036 3466
rect 502984 3402 503036 3408
rect 500224 2916 500276 2922
rect 500224 2858 500276 2864
rect 501052 2916 501104 2922
rect 501052 2858 501104 2864
rect 501064 480 501092 2858
rect 493294 354 493406 480
rect 492876 326 493406 354
rect 485566 -960 485678 326
rect 489430 -960 489542 326
rect 493294 -960 493406 326
rect 497158 -960 497270 480
rect 501022 -960 501134 480
rect 504468 354 504496 16546
rect 508780 3528 508832 3534
rect 508780 3470 508832 3476
rect 508792 480 508820 3470
rect 504886 354 504998 480
rect 504468 326 504998 354
rect 504886 -960 504998 326
rect 508750 -960 508862 480
rect 512196 354 512224 16546
rect 514036 3058 514064 22714
rect 518912 16574 518940 142258
rect 544396 142118 544424 192510
rect 548536 184385 548564 699654
rect 552664 690056 552716 690062
rect 552664 689998 552716 690004
rect 548616 669384 548668 669390
rect 548616 669326 548668 669332
rect 548522 184376 548578 184385
rect 548522 184311 548578 184320
rect 548628 180305 548656 669326
rect 552676 182889 552704 689998
rect 556804 685908 556856 685914
rect 556804 685850 556856 685856
rect 552756 681760 552808 681766
rect 552756 681702 552808 681708
rect 552768 182986 552796 681702
rect 555424 524476 555476 524482
rect 555424 524418 555476 524424
rect 554044 505164 554096 505170
rect 554044 505106 554096 505112
rect 552848 404388 552900 404394
rect 552848 404330 552900 404336
rect 552756 182980 552808 182986
rect 552756 182922 552808 182928
rect 552662 182880 552718 182889
rect 552662 182815 552718 182824
rect 552860 180606 552888 404330
rect 554056 184929 554084 505106
rect 554136 496868 554188 496874
rect 554136 496810 554188 496816
rect 554042 184920 554098 184929
rect 554042 184855 554098 184864
rect 552848 180600 552900 180606
rect 552848 180542 552900 180548
rect 548614 180296 548670 180305
rect 548614 180231 548670 180240
rect 554148 177857 554176 496810
rect 555436 180810 555464 524418
rect 555516 309188 555568 309194
rect 555516 309130 555568 309136
rect 555424 180804 555476 180810
rect 555424 180746 555476 180752
rect 554134 177848 554190 177857
rect 555528 177818 555556 309130
rect 554134 177783 554190 177792
rect 555516 177812 555568 177818
rect 555516 177754 555568 177760
rect 556816 174865 556844 685850
rect 556896 460964 556948 460970
rect 556896 460906 556948 460912
rect 556908 193089 556936 460906
rect 556988 372632 557040 372638
rect 556988 372574 557040 372580
rect 556894 193080 556950 193089
rect 556894 193015 556950 193024
rect 557000 177886 557028 372574
rect 558196 202201 558224 699654
rect 559564 694204 559616 694210
rect 559564 694146 559616 694152
rect 558276 641776 558328 641782
rect 558276 641718 558328 641724
rect 558182 202192 558238 202201
rect 558182 202127 558238 202136
rect 558288 184793 558316 641718
rect 558368 545148 558420 545154
rect 558368 545090 558420 545096
rect 558380 197305 558408 545090
rect 558460 345092 558512 345098
rect 558460 345034 558512 345040
rect 558366 197296 558422 197305
rect 558366 197231 558422 197240
rect 558274 184784 558330 184793
rect 558274 184719 558330 184728
rect 558472 180742 558500 345034
rect 558552 280220 558604 280226
rect 558552 280162 558604 280168
rect 558460 180736 558512 180742
rect 558460 180678 558512 180684
rect 556988 177880 557040 177886
rect 556988 177822 557040 177828
rect 558564 177342 558592 280162
rect 558552 177336 558604 177342
rect 558552 177278 558604 177284
rect 559576 175137 559604 694146
rect 560944 601724 560996 601730
rect 560944 601666 560996 601672
rect 559656 368552 559708 368558
rect 559656 368494 559708 368500
rect 559668 176662 559696 368494
rect 560956 185609 560984 601666
rect 561036 480276 561088 480282
rect 561036 480218 561088 480224
rect 560942 185600 560998 185609
rect 560942 185535 560998 185544
rect 561048 184249 561076 480218
rect 561128 473408 561180 473414
rect 561128 473350 561180 473356
rect 561140 196761 561168 473350
rect 561220 360256 561272 360262
rect 561220 360198 561272 360204
rect 561126 196752 561182 196761
rect 561126 196687 561182 196696
rect 561034 184240 561090 184249
rect 561034 184175 561090 184184
rect 561232 182102 561260 360198
rect 561312 288448 561364 288454
rect 561312 288390 561364 288396
rect 561220 182096 561272 182102
rect 561220 182038 561272 182044
rect 561324 177954 561352 288390
rect 561692 189961 561720 703582
rect 562704 703474 562732 703582
rect 562846 703520 562958 704960
rect 566710 703520 566822 704960
rect 569972 703582 570460 703610
rect 562888 703474 562916 703520
rect 562704 703446 562916 703474
rect 566752 700398 566780 703520
rect 566740 700392 566792 700398
rect 566740 700334 566792 700340
rect 566464 677612 566516 677618
rect 566464 677554 566516 677560
rect 562324 568608 562376 568614
rect 562324 568550 562376 568556
rect 561678 189952 561734 189961
rect 561678 189887 561734 189896
rect 561312 177948 561364 177954
rect 561312 177890 561364 177896
rect 559656 176656 559708 176662
rect 559656 176598 559708 176604
rect 562336 175166 562364 568550
rect 565084 541000 565136 541006
rect 565084 540942 565136 540948
rect 563704 448588 563756 448594
rect 563704 448530 563756 448536
rect 563716 190466 563744 448530
rect 563796 431996 563848 432002
rect 563796 431938 563848 431944
rect 563704 190460 563756 190466
rect 563704 190402 563756 190408
rect 563808 189009 563836 431938
rect 563888 429208 563940 429214
rect 563888 429150 563940 429156
rect 563900 189786 563928 429150
rect 563980 353320 564032 353326
rect 563980 353262 564032 353268
rect 563888 189780 563940 189786
rect 563888 189722 563940 189728
rect 563794 189000 563850 189009
rect 563794 188935 563850 188944
rect 563992 188358 564020 353262
rect 564072 276072 564124 276078
rect 564072 276014 564124 276020
rect 564084 194410 564112 276014
rect 564072 194404 564124 194410
rect 564072 194346 564124 194352
rect 563980 188352 564032 188358
rect 563980 188294 564032 188300
rect 565096 175234 565124 540942
rect 566476 191690 566504 677554
rect 566556 654152 566608 654158
rect 566556 654094 566608 654100
rect 566568 196897 566596 654094
rect 566648 488572 566700 488578
rect 566648 488514 566700 488520
rect 566554 196888 566610 196897
rect 566554 196823 566610 196832
rect 566464 191684 566516 191690
rect 566464 191626 566516 191632
rect 566660 187513 566688 488514
rect 567844 476128 567896 476134
rect 567844 476070 567896 476076
rect 566740 316056 566792 316062
rect 566740 315998 566792 316004
rect 566752 189038 566780 315998
rect 566832 264988 566884 264994
rect 566832 264930 566884 264936
rect 566740 189032 566792 189038
rect 566740 188974 566792 188980
rect 566646 187504 566702 187513
rect 566646 187439 566702 187448
rect 566844 178673 566872 264930
rect 567856 194478 567884 476070
rect 567936 436144 567988 436150
rect 567936 436086 567988 436092
rect 567844 194472 567896 194478
rect 567844 194414 567896 194420
rect 567948 186289 567976 436086
rect 569224 392012 569276 392018
rect 569224 391954 569276 391960
rect 569236 189854 569264 391954
rect 569316 376780 569368 376786
rect 569316 376722 569368 376728
rect 569224 189848 569276 189854
rect 569224 189790 569276 189796
rect 569328 187610 569356 376722
rect 569408 292596 569460 292602
rect 569408 292538 569460 292544
rect 569316 187604 569368 187610
rect 569316 187546 569368 187552
rect 567934 186280 567990 186289
rect 567934 186215 567990 186224
rect 569420 182918 569448 292538
rect 569972 262993 570000 703582
rect 570432 703474 570460 703582
rect 570574 703520 570686 704960
rect 574438 703520 574550 704960
rect 578302 703520 578414 704960
rect 581012 703582 582052 703610
rect 570616 703474 570644 703520
rect 570432 703446 570644 703474
rect 574480 700466 574508 703520
rect 574468 700460 574520 700466
rect 574468 700402 574520 700408
rect 578344 683114 578372 703520
rect 580170 702536 580226 702545
rect 580170 702471 580172 702480
rect 580224 702471 580226 702480
rect 580172 702442 580224 702448
rect 580170 698456 580226 698465
rect 580170 698391 580226 698400
rect 580184 698358 580212 698391
rect 580172 698352 580224 698358
rect 580172 698294 580224 698300
rect 580170 694376 580226 694385
rect 580170 694311 580226 694320
rect 580184 694210 580212 694311
rect 580172 694204 580224 694210
rect 580172 694146 580224 694152
rect 580170 690296 580226 690305
rect 580170 690231 580226 690240
rect 580184 690062 580212 690231
rect 580172 690056 580224 690062
rect 580172 689998 580224 690004
rect 579802 686216 579858 686225
rect 579802 686151 579858 686160
rect 579816 685914 579844 686151
rect 579804 685908 579856 685914
rect 579804 685850 579856 685856
rect 578252 683086 578372 683114
rect 570604 625184 570656 625190
rect 570604 625126 570656 625132
rect 569958 262984 570014 262993
rect 569958 262919 570014 262928
rect 570616 196625 570644 625126
rect 576124 621036 576176 621042
rect 576124 620978 576176 620984
rect 574744 589348 574796 589354
rect 574744 589290 574796 589296
rect 571984 549296 572036 549302
rect 571984 549238 572036 549244
rect 570696 444440 570748 444446
rect 570696 444382 570748 444388
rect 570602 196616 570658 196625
rect 570602 196551 570658 196560
rect 569408 182912 569460 182918
rect 569408 182854 569460 182860
rect 570708 181529 570736 444382
rect 571996 194585 572024 549238
rect 573364 465112 573416 465118
rect 573364 465054 573416 465060
rect 572076 440292 572128 440298
rect 572076 440234 572128 440240
rect 571982 194576 572038 194585
rect 571982 194511 572038 194520
rect 572088 189922 572116 440234
rect 572168 412684 572220 412690
rect 572168 412626 572220 412632
rect 572076 189916 572128 189922
rect 572076 189858 572128 189864
rect 572180 186998 572208 412626
rect 572260 332648 572312 332654
rect 572260 332590 572312 332596
rect 572272 191758 572300 332590
rect 572352 305040 572404 305046
rect 572352 304982 572404 304988
rect 572260 191752 572312 191758
rect 572260 191694 572312 191700
rect 572168 186992 572220 186998
rect 572168 186934 572220 186940
rect 572364 182170 572392 304982
rect 573376 183161 573404 465054
rect 574756 195945 574784 589290
rect 574836 509312 574888 509318
rect 574836 509254 574888 509260
rect 574742 195936 574798 195945
rect 574742 195871 574798 195880
rect 574848 189689 574876 509254
rect 574928 492720 574980 492726
rect 574928 492662 574980 492668
rect 574940 192681 574968 492662
rect 575020 340944 575072 340950
rect 575020 340886 575072 340892
rect 574926 192672 574982 192681
rect 574926 192607 574982 192616
rect 575032 191826 575060 340886
rect 575112 320204 575164 320210
rect 575112 320146 575164 320152
rect 575124 192642 575152 320146
rect 575204 273284 575256 273290
rect 575204 273226 575256 273232
rect 575112 192636 575164 192642
rect 575112 192578 575164 192584
rect 575020 191820 575072 191826
rect 575020 191762 575072 191768
rect 574834 189680 574890 189689
rect 574834 189615 574890 189624
rect 573362 183152 573418 183161
rect 573362 183087 573418 183096
rect 575216 182850 575244 273226
rect 576136 183025 576164 620978
rect 576216 553444 576268 553450
rect 576216 553386 576268 553392
rect 576228 192409 576256 553386
rect 577504 529100 577556 529106
rect 577504 529042 577556 529048
rect 576308 501016 576360 501022
rect 576308 500958 576360 500964
rect 576214 192400 576270 192409
rect 576214 192335 576270 192344
rect 576320 191185 576348 500958
rect 576398 259584 576454 259593
rect 576398 259519 576454 259528
rect 576412 205630 576440 259519
rect 576400 205624 576452 205630
rect 576400 205566 576452 205572
rect 577516 195401 577544 529042
rect 577596 425128 577648 425134
rect 577596 425070 577648 425076
rect 577502 195392 577558 195401
rect 577502 195327 577558 195336
rect 577608 193186 577636 425070
rect 577688 313336 577740 313342
rect 577688 313278 577740 313284
rect 577700 195906 577728 313278
rect 577780 300892 577832 300898
rect 577780 300834 577832 300840
rect 577688 195900 577740 195906
rect 577688 195842 577740 195848
rect 577792 195537 577820 300834
rect 577872 260908 577924 260914
rect 577872 260850 577924 260856
rect 577778 195528 577834 195537
rect 577778 195463 577834 195472
rect 577596 193180 577648 193186
rect 577596 193122 577648 193128
rect 576306 191176 576362 191185
rect 576306 191111 576362 191120
rect 577884 189825 577912 260850
rect 577870 189816 577926 189825
rect 577870 189751 577926 189760
rect 576122 183016 576178 183025
rect 576122 182951 576178 182960
rect 575204 182844 575256 182850
rect 575204 182786 575256 182792
rect 572352 182164 572404 182170
rect 572352 182106 572404 182112
rect 570694 181520 570750 181529
rect 570694 181455 570750 181464
rect 578252 181393 578280 683086
rect 580170 682136 580226 682145
rect 580170 682071 580226 682080
rect 580184 681766 580212 682071
rect 580172 681760 580224 681766
rect 580172 681702 580224 681708
rect 580170 678056 580226 678065
rect 580170 677991 580226 678000
rect 580184 677618 580212 677991
rect 580172 677612 580224 677618
rect 580172 677554 580224 677560
rect 580170 673976 580226 673985
rect 580170 673911 580226 673920
rect 580184 673538 580212 673911
rect 580172 673532 580224 673538
rect 580172 673474 580224 673480
rect 580170 669896 580226 669905
rect 580170 669831 580226 669840
rect 580184 669390 580212 669831
rect 580172 669384 580224 669390
rect 580172 669326 580224 669332
rect 580170 662416 580226 662425
rect 580170 662351 580226 662360
rect 580184 661094 580212 662351
rect 580172 661088 580224 661094
rect 580172 661030 580224 661036
rect 580170 658336 580226 658345
rect 580170 658271 580172 658280
rect 580224 658271 580226 658280
rect 580172 658242 580224 658248
rect 580170 654256 580226 654265
rect 580170 654191 580226 654200
rect 580184 654158 580212 654191
rect 580172 654152 580224 654158
rect 580172 654094 580224 654100
rect 580170 646096 580226 646105
rect 580170 646031 580226 646040
rect 580184 645930 580212 646031
rect 580172 645924 580224 645930
rect 580172 645866 580224 645872
rect 580170 642016 580226 642025
rect 580170 641951 580226 641960
rect 580184 641782 580212 641951
rect 580172 641776 580224 641782
rect 580172 641718 580224 641724
rect 580170 626376 580226 626385
rect 580170 626311 580226 626320
rect 580184 625190 580212 626311
rect 580172 625184 580224 625190
rect 580172 625126 580224 625132
rect 579802 622296 579858 622305
rect 579802 622231 579858 622240
rect 579816 621042 579844 622231
rect 579804 621036 579856 621042
rect 579804 620978 579856 620984
rect 580170 605976 580226 605985
rect 580170 605911 580226 605920
rect 580184 605878 580212 605911
rect 580172 605872 580224 605878
rect 580172 605814 580224 605820
rect 580170 601896 580226 601905
rect 580170 601831 580226 601840
rect 580184 601730 580212 601831
rect 580172 601724 580224 601730
rect 580172 601666 580224 601672
rect 580354 597816 580410 597825
rect 580354 597751 580410 597760
rect 580170 589656 580226 589665
rect 580170 589591 580226 589600
rect 580184 589354 580212 589591
rect 580172 589348 580224 589354
rect 580172 589290 580224 589296
rect 578882 586256 578938 586265
rect 578882 586191 578938 586200
rect 578896 191049 578924 586191
rect 580170 569936 580226 569945
rect 580170 569871 580226 569880
rect 580184 568614 580212 569871
rect 580172 568608 580224 568614
rect 580172 568550 580224 568556
rect 580172 565888 580224 565894
rect 580170 565856 580172 565865
rect 580224 565856 580226 565865
rect 580170 565791 580226 565800
rect 580170 553616 580226 553625
rect 580170 553551 580226 553560
rect 580184 553450 580212 553551
rect 580172 553444 580224 553450
rect 580172 553386 580224 553392
rect 580170 549536 580226 549545
rect 580170 549471 580226 549480
rect 580184 549302 580212 549471
rect 580172 549296 580224 549302
rect 580172 549238 580224 549244
rect 579894 546136 579950 546145
rect 579894 546071 579950 546080
rect 579908 545154 579936 546071
rect 579896 545148 579948 545154
rect 579896 545090 579948 545096
rect 580170 542056 580226 542065
rect 580170 541991 580226 542000
rect 580184 541006 580212 541991
rect 580172 541000 580224 541006
rect 580172 540942 580224 540948
rect 580170 537976 580226 537985
rect 580170 537911 580226 537920
rect 580184 536858 580212 537911
rect 580172 536852 580224 536858
rect 580172 536794 580224 536800
rect 579802 529816 579858 529825
rect 579802 529751 579858 529760
rect 579816 529106 579844 529751
rect 579804 529100 579856 529106
rect 579804 529042 579856 529048
rect 580170 525736 580226 525745
rect 580170 525671 580226 525680
rect 580184 524482 580212 525671
rect 580172 524476 580224 524482
rect 580172 524418 580224 524424
rect 580170 521656 580226 521665
rect 580170 521591 580226 521600
rect 580184 520334 580212 521591
rect 580172 520328 580224 520334
rect 580172 520270 580224 520276
rect 580170 510096 580226 510105
rect 580170 510031 580226 510040
rect 580184 509318 580212 510031
rect 580172 509312 580224 509318
rect 580172 509254 580224 509260
rect 580078 506016 580134 506025
rect 580078 505951 580134 505960
rect 580092 505170 580120 505951
rect 580080 505164 580132 505170
rect 580080 505106 580132 505112
rect 580078 501936 580134 501945
rect 580078 501871 580134 501880
rect 580092 501022 580120 501871
rect 580080 501016 580132 501022
rect 580080 500958 580132 500964
rect 579894 497856 579950 497865
rect 579894 497791 579950 497800
rect 579908 496874 579936 497791
rect 579896 496868 579948 496874
rect 579896 496810 579948 496816
rect 580170 493776 580226 493785
rect 580170 493711 580226 493720
rect 580184 492726 580212 493711
rect 580172 492720 580224 492726
rect 580172 492662 580224 492668
rect 580170 489696 580226 489705
rect 580170 489631 580226 489640
rect 580184 488578 580212 489631
rect 580172 488572 580224 488578
rect 580172 488514 580224 488520
rect 580170 485616 580226 485625
rect 580170 485551 580226 485560
rect 580184 484430 580212 485551
rect 580172 484424 580224 484430
rect 580172 484366 580224 484372
rect 580170 481536 580226 481545
rect 580170 481471 580226 481480
rect 580184 480282 580212 481471
rect 580172 480276 580224 480282
rect 580172 480218 580224 480224
rect 580170 477456 580226 477465
rect 580170 477391 580226 477400
rect 580184 476134 580212 477391
rect 580172 476128 580224 476134
rect 580172 476070 580224 476076
rect 580172 473408 580224 473414
rect 580170 473376 580172 473385
rect 580224 473376 580226 473385
rect 580170 473311 580226 473320
rect 580170 465896 580226 465905
rect 580170 465831 580226 465840
rect 580184 465118 580212 465831
rect 580172 465112 580224 465118
rect 580172 465054 580224 465060
rect 580078 461816 580134 461825
rect 580078 461751 580134 461760
rect 580092 460970 580120 461751
rect 580080 460964 580132 460970
rect 580080 460906 580132 460912
rect 580078 457736 580134 457745
rect 580078 457671 580134 457680
rect 580092 456822 580120 457671
rect 580080 456816 580132 456822
rect 580080 456758 580132 456764
rect 578974 453656 579030 453665
rect 578974 453591 579030 453600
rect 578988 194546 579016 453591
rect 579710 449576 579766 449585
rect 579710 449511 579766 449520
rect 579724 448594 579752 449511
rect 579712 448588 579764 448594
rect 579712 448530 579764 448536
rect 580170 445496 580226 445505
rect 580170 445431 580226 445440
rect 580184 444446 580212 445431
rect 580172 444440 580224 444446
rect 580172 444382 580224 444388
rect 580170 441416 580226 441425
rect 580170 441351 580226 441360
rect 580184 440298 580212 441351
rect 580172 440292 580224 440298
rect 580172 440234 580224 440240
rect 579618 437336 579674 437345
rect 579618 437271 579674 437280
rect 579632 436150 579660 437271
rect 579620 436144 579672 436150
rect 579620 436086 579672 436092
rect 580170 433256 580226 433265
rect 580170 433191 580226 433200
rect 580184 432002 580212 433191
rect 580172 431996 580224 432002
rect 580172 431938 580224 431944
rect 579986 429856 580042 429865
rect 579986 429791 580042 429800
rect 580000 429214 580028 429791
rect 579988 429208 580040 429214
rect 579988 429150 580040 429156
rect 579618 425776 579674 425785
rect 579618 425711 579674 425720
rect 579632 425134 579660 425711
rect 579620 425128 579672 425134
rect 579620 425070 579672 425076
rect 580170 413536 580226 413545
rect 580170 413471 580226 413480
rect 580184 412690 580212 413471
rect 580172 412684 580224 412690
rect 580172 412626 580224 412632
rect 580170 405376 580226 405385
rect 580170 405311 580226 405320
rect 580184 404394 580212 405311
rect 580172 404388 580224 404394
rect 580172 404330 580224 404336
rect 580170 401296 580226 401305
rect 580170 401231 580226 401240
rect 580184 400246 580212 401231
rect 580172 400240 580224 400246
rect 580172 400182 580224 400188
rect 580170 393136 580226 393145
rect 580170 393071 580226 393080
rect 580184 392018 580212 393071
rect 580172 392012 580224 392018
rect 580172 391954 580224 391960
rect 579802 385656 579858 385665
rect 579802 385591 579858 385600
rect 579816 385082 579844 385591
rect 579804 385076 579856 385082
rect 579804 385018 579856 385024
rect 579986 381576 580042 381585
rect 579986 381511 580042 381520
rect 580000 380934 580028 381511
rect 579988 380928 580040 380934
rect 579988 380870 580040 380876
rect 580170 377496 580226 377505
rect 580170 377431 580226 377440
rect 580184 376786 580212 377431
rect 580172 376780 580224 376786
rect 580172 376722 580224 376728
rect 580170 373416 580226 373425
rect 580170 373351 580226 373360
rect 580184 372638 580212 373351
rect 580172 372632 580224 372638
rect 580172 372574 580224 372580
rect 580170 369336 580226 369345
rect 580170 369271 580226 369280
rect 580184 368558 580212 369271
rect 580172 368552 580224 368558
rect 580172 368494 580224 368500
rect 579618 365256 579674 365265
rect 579618 365191 579674 365200
rect 579632 364410 579660 365191
rect 579620 364404 579672 364410
rect 579620 364346 579672 364352
rect 579618 361176 579674 361185
rect 579618 361111 579674 361120
rect 579632 360262 579660 361111
rect 579620 360256 579672 360262
rect 579620 360198 579672 360204
rect 580170 357096 580226 357105
rect 580170 357031 580226 357040
rect 580184 356114 580212 357031
rect 580172 356108 580224 356114
rect 580172 356050 580224 356056
rect 579618 353696 579674 353705
rect 579618 353631 579674 353640
rect 579632 353326 579660 353631
rect 579620 353320 579672 353326
rect 579620 353262 579672 353268
rect 580170 349616 580226 349625
rect 580170 349551 580226 349560
rect 580184 349178 580212 349551
rect 580172 349172 580224 349178
rect 580172 349114 580224 349120
rect 580170 345536 580226 345545
rect 580170 345471 580226 345480
rect 580184 345098 580212 345471
rect 580172 345092 580224 345098
rect 580172 345034 580224 345040
rect 580170 341456 580226 341465
rect 580170 341391 580226 341400
rect 580184 340950 580212 341391
rect 580172 340944 580224 340950
rect 580172 340886 580224 340892
rect 579986 337376 580042 337385
rect 579986 337311 580042 337320
rect 580000 336802 580028 337311
rect 579988 336796 580040 336802
rect 579988 336738 580040 336744
rect 579986 333296 580042 333305
rect 579986 333231 580042 333240
rect 580000 332654 580028 333231
rect 579988 332648 580040 332654
rect 579988 332590 580040 332596
rect 579618 321056 579674 321065
rect 579618 320991 579674 321000
rect 579632 320210 579660 320991
rect 579620 320204 579672 320210
rect 579620 320146 579672 320152
rect 579618 316976 579674 316985
rect 579618 316911 579674 316920
rect 579632 316062 579660 316911
rect 579620 316056 579672 316062
rect 579620 315998 579672 316004
rect 580170 309496 580226 309505
rect 580170 309431 580226 309440
rect 580184 309194 580212 309431
rect 580172 309188 580224 309194
rect 580172 309130 580224 309136
rect 579618 305416 579674 305425
rect 579618 305351 579674 305360
rect 579632 305046 579660 305351
rect 579620 305040 579672 305046
rect 579620 304982 579672 304988
rect 580170 297256 580226 297265
rect 580170 297191 580226 297200
rect 580184 296750 580212 297191
rect 580172 296744 580224 296750
rect 580172 296686 580224 296692
rect 579986 293176 580042 293185
rect 579986 293111 580042 293120
rect 580000 292602 580028 293111
rect 579988 292596 580040 292602
rect 579988 292538 580040 292544
rect 579986 289096 580042 289105
rect 579986 289031 580042 289040
rect 580000 288454 580028 289031
rect 579988 288448 580040 288454
rect 579988 288390 580040 288396
rect 579066 285016 579122 285025
rect 579066 284951 579122 284960
rect 578976 194540 579028 194546
rect 578976 194482 579028 194488
rect 578882 191040 578938 191049
rect 578882 190975 578938 190984
rect 579080 187678 579108 284951
rect 580170 280936 580226 280945
rect 580170 280871 580226 280880
rect 580184 280226 580212 280871
rect 580172 280220 580224 280226
rect 580172 280162 580224 280168
rect 580170 276856 580226 276865
rect 580170 276791 580226 276800
rect 580184 276078 580212 276791
rect 580172 276072 580224 276078
rect 580172 276014 580224 276020
rect 580170 273456 580226 273465
rect 580170 273391 580226 273400
rect 580184 273290 580212 273391
rect 580172 273284 580224 273290
rect 580172 273226 580224 273232
rect 580170 265296 580226 265305
rect 580170 265231 580226 265240
rect 580184 264994 580212 265231
rect 580172 264988 580224 264994
rect 580172 264930 580224 264936
rect 580262 257136 580318 257145
rect 580262 257071 580318 257080
rect 579802 253056 579858 253065
rect 579802 252991 579858 253000
rect 579816 252618 579844 252991
rect 579804 252612 579856 252618
rect 579804 252554 579856 252560
rect 579802 248976 579858 248985
rect 579802 248911 579858 248920
rect 579816 248470 579844 248911
rect 579804 248464 579856 248470
rect 579804 248406 579856 248412
rect 580170 244896 580226 244905
rect 580170 244831 580226 244840
rect 580184 244322 580212 244831
rect 580172 244316 580224 244322
rect 580172 244258 580224 244264
rect 580172 237448 580224 237454
rect 580170 237416 580172 237425
rect 580224 237416 580226 237425
rect 580170 237351 580226 237360
rect 580170 221096 580226 221105
rect 580170 221031 580226 221040
rect 580184 220862 580212 221031
rect 580172 220856 580224 220862
rect 580172 220798 580224 220804
rect 580172 217320 580224 217326
rect 580172 217262 580224 217268
rect 580184 217025 580212 217262
rect 580170 217016 580226 217025
rect 580170 216951 580226 216960
rect 579988 205624 580040 205630
rect 579988 205566 580040 205572
rect 580000 204785 580028 205566
rect 579986 204776 580042 204785
rect 579986 204711 580042 204720
rect 580170 200696 580226 200705
rect 580170 200631 580226 200640
rect 580184 200190 580212 200631
rect 580172 200184 580224 200190
rect 580172 200126 580224 200132
rect 580170 197296 580226 197305
rect 580170 197231 580226 197240
rect 580184 196110 580212 197231
rect 580172 196104 580224 196110
rect 580172 196046 580224 196052
rect 580276 195974 580304 257071
rect 580264 195968 580316 195974
rect 580264 195910 580316 195916
rect 580368 195265 580396 597751
rect 580446 469976 580502 469985
rect 580446 469911 580502 469920
rect 580354 195256 580410 195265
rect 580354 195191 580410 195200
rect 579618 193216 579674 193225
rect 579618 193151 579674 193160
rect 579632 192506 579660 193151
rect 579620 192500 579672 192506
rect 579620 192442 579672 192448
rect 579988 190392 580040 190398
rect 579988 190334 580040 190340
rect 580000 189145 580028 190334
rect 579986 189136 580042 189145
rect 579986 189071 580042 189080
rect 579068 187672 579120 187678
rect 580460 187649 580488 469911
rect 580538 389736 580594 389745
rect 580538 389671 580594 389680
rect 580552 192545 580580 389671
rect 580630 313576 580686 313585
rect 580630 313511 580686 313520
rect 580644 313342 580672 313511
rect 580632 313336 580684 313342
rect 580632 313278 580684 313284
rect 580630 301336 580686 301345
rect 580630 301271 580686 301280
rect 580644 300898 580672 301271
rect 580632 300892 580684 300898
rect 580632 300834 580684 300840
rect 580630 269376 580686 269385
rect 580630 269311 580686 269320
rect 580644 206310 580672 269311
rect 580722 261216 580778 261225
rect 580722 261151 580778 261160
rect 580736 260914 580764 261151
rect 580724 260908 580776 260914
rect 580724 260850 580776 260856
rect 580722 240816 580778 240825
rect 580722 240751 580778 240760
rect 580632 206304 580684 206310
rect 580632 206246 580684 206252
rect 580736 200802 580764 240751
rect 580814 225176 580870 225185
rect 580814 225111 580870 225120
rect 580724 200796 580776 200802
rect 580724 200738 580776 200744
rect 580632 196036 580684 196042
rect 580632 195978 580684 195984
rect 580538 192536 580594 192545
rect 580538 192471 580594 192480
rect 579068 187614 579120 187620
rect 580446 187640 580502 187649
rect 580446 187575 580502 187584
rect 580170 185056 580226 185065
rect 580170 184991 580226 185000
rect 580184 184958 580212 184991
rect 580172 184952 580224 184958
rect 580172 184894 580224 184900
rect 578238 181384 578294 181393
rect 578238 181319 578294 181328
rect 580170 180976 580226 180985
rect 580170 180911 580226 180920
rect 580184 180878 580212 180911
rect 580172 180872 580224 180878
rect 580172 180814 580224 180820
rect 566830 178664 566886 178673
rect 566830 178599 566886 178608
rect 579802 176896 579858 176905
rect 579802 176831 579858 176840
rect 579816 176730 579844 176831
rect 579804 176724 579856 176730
rect 579804 176666 579856 176672
rect 565084 175228 565136 175234
rect 565084 175170 565136 175176
rect 562324 175160 562376 175166
rect 559562 175128 559618 175137
rect 562324 175102 562376 175108
rect 559562 175063 559618 175072
rect 556802 174856 556858 174865
rect 556802 174791 556858 174800
rect 580262 172816 580318 172825
rect 580262 172751 580318 172760
rect 580170 164656 580226 164665
rect 580170 164591 580226 164600
rect 580184 164286 580212 164591
rect 580172 164280 580224 164286
rect 580172 164222 580224 164228
rect 580172 157344 580224 157350
rect 580172 157286 580224 157292
rect 580184 157185 580212 157286
rect 580170 157176 580226 157185
rect 580170 157111 580226 157120
rect 579802 153096 579858 153105
rect 579802 153031 579858 153040
rect 579816 151842 579844 153031
rect 579804 151836 579856 151842
rect 579804 151778 579856 151784
rect 580172 146260 580224 146266
rect 580172 146202 580224 146208
rect 580184 144945 580212 146202
rect 580170 144936 580226 144945
rect 580276 144906 580304 172751
rect 580354 168736 580410 168745
rect 580354 168671 580410 168680
rect 580368 147626 580396 168671
rect 580356 147620 580408 147626
rect 580356 147562 580408 147568
rect 580170 144871 580226 144880
rect 580264 144900 580316 144906
rect 580264 144842 580316 144848
rect 580540 143676 580592 143682
rect 580540 143618 580592 143624
rect 580448 143608 580500 143614
rect 580448 143550 580500 143556
rect 580264 142248 580316 142254
rect 580264 142190 580316 142196
rect 544384 142112 544436 142118
rect 544384 142054 544436 142060
rect 580172 142112 580224 142118
rect 580172 142054 580224 142060
rect 580184 140865 580212 142054
rect 580170 140856 580226 140865
rect 580170 140791 580226 140800
rect 579802 132696 579858 132705
rect 579802 132631 579858 132640
rect 579816 132530 579844 132631
rect 579804 132524 579856 132530
rect 579804 132466 579856 132472
rect 580170 108896 580226 108905
rect 580170 108831 580226 108840
rect 580184 107710 580212 108831
rect 580172 107704 580224 107710
rect 580172 107646 580224 107652
rect 580172 81388 580224 81394
rect 580172 81330 580224 81336
rect 580184 81025 580212 81330
rect 580170 81016 580226 81025
rect 580170 80951 580226 80960
rect 534078 75168 534134 75177
rect 534078 75103 534134 75112
rect 527180 17264 527232 17270
rect 527180 17206 527232 17212
rect 527192 16574 527220 17206
rect 534092 16574 534120 75103
rect 560944 73840 560996 73846
rect 560944 73782 560996 73788
rect 545764 58676 545816 58682
rect 545764 58618 545816 58624
rect 542360 53100 542412 53106
rect 542360 53042 542412 53048
rect 542372 16574 542400 53042
rect 518912 16546 519768 16574
rect 527192 16546 527496 16574
rect 534092 16546 535224 16574
rect 542372 16546 542952 16574
rect 514024 3052 514076 3058
rect 514024 2994 514076 3000
rect 515864 3052 515916 3058
rect 515864 2994 515916 3000
rect 515876 480 515904 2994
rect 519740 480 519768 16546
rect 527468 480 527496 16546
rect 531320 13116 531372 13122
rect 531320 13058 531372 13064
rect 531332 480 531360 13058
rect 535196 480 535224 16546
rect 539048 3460 539100 3466
rect 539048 3402 539100 3408
rect 539060 480 539088 3402
rect 542924 480 542952 16546
rect 545776 3534 545804 58618
rect 553400 50380 553452 50386
rect 553400 50322 553452 50328
rect 548524 35216 548576 35222
rect 548524 35158 548576 35164
rect 545764 3528 545816 3534
rect 545764 3470 545816 3476
rect 546776 3528 546828 3534
rect 546776 3470 546828 3476
rect 546788 480 546816 3470
rect 548536 3126 548564 35158
rect 548524 3120 548576 3126
rect 548524 3062 548576 3068
rect 550640 3120 550692 3126
rect 550640 3062 550692 3068
rect 550652 480 550680 3062
rect 512614 354 512726 480
rect 512196 326 512726 354
rect 512614 -960 512726 326
rect 515834 -960 515946 480
rect 519698 -960 519810 480
rect 523562 -960 523674 480
rect 527426 -960 527538 480
rect 531290 -960 531402 480
rect 535154 -960 535266 480
rect 539018 -960 539130 480
rect 542882 -960 542994 480
rect 546746 -960 546858 480
rect 550610 -960 550722 480
rect 553412 354 553440 50322
rect 556804 46232 556856 46238
rect 556804 46174 556856 46180
rect 556816 3466 556844 46174
rect 557540 43444 557592 43450
rect 557540 43386 557592 43392
rect 556804 3460 556856 3466
rect 556804 3402 556856 3408
rect 553830 354 553942 480
rect 553412 326 553942 354
rect 557552 354 557580 43386
rect 560956 8294 560984 73782
rect 580172 73160 580224 73166
rect 580172 73102 580224 73108
rect 580184 72865 580212 73102
rect 580170 72856 580226 72865
rect 580170 72791 580226 72800
rect 579618 69592 579674 69601
rect 579618 69527 579674 69536
rect 578884 54528 578936 54534
rect 578884 54470 578936 54476
rect 571984 33176 572036 33182
rect 571984 33118 572036 33124
rect 563704 31068 563756 31074
rect 563704 31010 563756 31016
rect 562324 10328 562376 10334
rect 562324 10270 562376 10276
rect 560944 8288 560996 8294
rect 560944 8230 560996 8236
rect 562336 3466 562364 10270
rect 561588 3460 561640 3466
rect 561588 3402 561640 3408
rect 562324 3460 562376 3466
rect 562324 3402 562376 3408
rect 561600 480 561628 3402
rect 563716 3058 563744 31010
rect 571996 3534 572024 33118
rect 571984 3528 572036 3534
rect 571984 3470 572036 3476
rect 573180 3528 573232 3534
rect 573180 3470 573232 3476
rect 563704 3052 563756 3058
rect 563704 2994 563756 3000
rect 565452 3052 565504 3058
rect 565452 2994 565504 3000
rect 565464 480 565492 2994
rect 573192 480 573220 3470
rect 577044 3392 577096 3398
rect 577044 3334 577096 3340
rect 577056 480 577084 3334
rect 578896 785 578924 54470
rect 579632 6914 579660 69527
rect 580276 60625 580304 142190
rect 580356 141432 580408 141438
rect 580356 141374 580408 141380
rect 580368 68785 580396 141374
rect 580460 76945 580488 143550
rect 580552 84425 580580 143618
rect 580644 128625 580672 195978
rect 580828 195294 580856 225111
rect 580816 195288 580868 195294
rect 580816 195230 580868 195236
rect 581012 188329 581040 703582
rect 582024 703474 582052 703582
rect 582166 703520 582278 704960
rect 582208 703474 582236 703520
rect 582024 703446 582236 703474
rect 582470 637936 582526 637945
rect 582470 637871 582526 637880
rect 582378 629776 582434 629785
rect 582378 629711 582434 629720
rect 581642 610056 581698 610065
rect 581642 609991 581698 610000
rect 580998 188320 581054 188329
rect 580998 188255 581054 188264
rect 581656 185638 581684 609991
rect 581734 574016 581790 574025
rect 581734 573951 581790 573960
rect 581748 193905 581776 573951
rect 581734 193896 581790 193905
rect 581734 193831 581790 193840
rect 581644 185632 581696 185638
rect 581644 185574 581696 185580
rect 582392 178022 582420 629711
rect 582484 199442 582512 637871
rect 582562 614136 582618 614145
rect 582562 614071 582618 614080
rect 582472 199436 582524 199442
rect 582472 199378 582524 199384
rect 582576 198014 582604 614071
rect 582654 557696 582710 557705
rect 582654 557631 582710 557640
rect 582564 198008 582616 198014
rect 582564 197950 582616 197956
rect 582668 179382 582696 557631
rect 582746 533896 582802 533905
rect 582746 533831 582802 533840
rect 582760 180033 582788 533831
rect 582838 517576 582894 517585
rect 582838 517511 582894 517520
rect 582852 180169 582880 517511
rect 582838 180160 582894 180169
rect 582838 180095 582894 180104
rect 582746 180024 582802 180033
rect 582746 179959 582802 179968
rect 582656 179376 582708 179382
rect 582656 179318 582708 179324
rect 582380 178016 582432 178022
rect 582380 177958 582432 177964
rect 580816 146396 580868 146402
rect 580816 146338 580868 146344
rect 580724 142180 580776 142186
rect 580724 142122 580776 142128
rect 580630 128616 580686 128625
rect 580630 128551 580686 128560
rect 580630 96656 580686 96665
rect 580630 96591 580686 96600
rect 580538 84416 580594 84425
rect 580538 84351 580594 84360
rect 580446 76936 580502 76945
rect 580446 76871 580502 76880
rect 580354 68776 580410 68785
rect 580354 68711 580410 68720
rect 580644 63481 580672 96591
rect 580736 92585 580764 142122
rect 580828 112985 580856 146338
rect 580908 146328 580960 146334
rect 580908 146270 580960 146276
rect 580920 117065 580948 146270
rect 580906 117056 580962 117065
rect 580906 116991 580962 117000
rect 580814 112976 580870 112985
rect 580814 112911 580870 112920
rect 580814 104816 580870 104825
rect 580814 104751 580870 104760
rect 580722 92576 580778 92585
rect 580722 92511 580778 92520
rect 580722 88496 580778 88505
rect 580722 88431 580778 88440
rect 580736 64870 580764 88431
rect 580828 79626 580856 104751
rect 580906 100736 580962 100745
rect 580906 100671 580962 100680
rect 580816 79620 580868 79626
rect 580816 79562 580868 79568
rect 580920 78713 580948 100671
rect 580906 78704 580962 78713
rect 580906 78639 580962 78648
rect 580724 64864 580776 64870
rect 580724 64806 580776 64812
rect 580630 63472 580686 63481
rect 580630 63407 580686 63416
rect 580262 60616 580318 60625
rect 580262 60551 580318 60560
rect 579896 56568 579948 56574
rect 579894 56536 579896 56545
rect 579948 56536 579950 56545
rect 579894 56471 579950 56480
rect 579894 52456 579950 52465
rect 579894 52391 579896 52400
rect 579948 52391 579950 52400
rect 579896 52362 579948 52368
rect 580172 49700 580224 49706
rect 580172 49642 580224 49648
rect 580184 48385 580212 49642
rect 580170 48376 580226 48385
rect 580170 48311 580226 48320
rect 579988 45552 580040 45558
rect 579988 45494 580040 45500
rect 580000 44305 580028 45494
rect 579986 44296 580042 44305
rect 579986 44231 580042 44240
rect 580172 41404 580224 41410
rect 580172 41346 580224 41352
rect 580184 40905 580212 41346
rect 580170 40896 580226 40905
rect 580170 40831 580226 40840
rect 580172 37256 580224 37262
rect 580172 37198 580224 37204
rect 580184 36825 580212 37198
rect 580170 36816 580226 36825
rect 580170 36751 580226 36760
rect 580172 33108 580224 33114
rect 580172 33050 580224 33056
rect 580184 32745 580212 33050
rect 580170 32736 580226 32745
rect 580170 32671 580226 32680
rect 580172 28960 580224 28966
rect 580172 28902 580224 28908
rect 580184 28665 580212 28902
rect 580170 28656 580226 28665
rect 580170 28591 580226 28600
rect 580172 24812 580224 24818
rect 580172 24754 580224 24760
rect 580184 24585 580212 24754
rect 580170 24576 580226 24585
rect 580170 24511 580226 24520
rect 580172 20664 580224 20670
rect 580172 20606 580224 20612
rect 580184 20505 580212 20606
rect 580170 20496 580226 20505
rect 580170 20431 580226 20440
rect 580172 16584 580224 16590
rect 580172 16526 580224 16532
rect 580184 16425 580212 16526
rect 580170 16416 580226 16425
rect 580170 16351 580226 16360
rect 580172 12436 580224 12442
rect 580172 12378 580224 12384
rect 580184 12345 580212 12378
rect 580170 12336 580226 12345
rect 580170 12271 580226 12280
rect 580172 8288 580224 8294
rect 580170 8256 580172 8265
rect 580224 8256 580226 8265
rect 580170 8191 580226 8200
rect 579632 6886 580488 6914
rect 580172 5500 580224 5506
rect 580172 5442 580224 5448
rect 580184 4865 580212 5442
rect 580170 4856 580226 4865
rect 580170 4791 580226 4800
rect 578882 776 578938 785
rect 578882 711 578938 720
rect 557694 354 557806 480
rect 557552 326 557806 354
rect 553830 -960 553942 326
rect 557694 -960 557806 326
rect 561558 -960 561670 480
rect 565422 -960 565534 480
rect 569286 -960 569398 480
rect 573150 -960 573262 480
rect 577014 -960 577126 480
rect 580460 354 580488 6886
rect 580878 354 580990 480
rect 580460 326 580990 354
rect 580878 -960 580990 326
<< via2 >>
rect 3422 701120 3478 701176
rect 3054 697720 3110 697776
rect 3422 689560 3478 689616
rect 3146 685480 3202 685536
rect 3422 681400 3478 681456
rect 3422 677320 3478 677376
rect 3238 665080 3294 665136
rect 3422 661036 3424 661056
rect 3424 661036 3476 661056
rect 3476 661036 3478 661056
rect 3422 661000 3478 661036
rect 3054 653520 3110 653576
rect 3422 645360 3478 645416
rect 3146 641280 3202 641336
rect 3146 637200 3202 637256
rect 3422 633120 3478 633176
rect 3238 624960 3294 625016
rect 3422 621560 3478 621616
rect 3146 617480 3202 617536
rect 3146 613400 3202 613456
rect 3422 609320 3478 609376
rect 3054 605240 3110 605296
rect 3054 597080 3110 597136
rect 3146 593000 3202 593056
rect 3238 588920 3294 588976
rect 3146 584840 3202 584896
rect 3330 581440 3386 581496
rect 2870 569200 2926 569256
rect 3054 561040 3110 561096
rect 3054 556960 3110 557016
rect 3054 548800 3110 548856
rect 3146 544720 3202 544776
rect 3330 537240 3386 537296
rect 3330 533160 3386 533216
rect 2870 520920 2926 520976
rect 2962 516840 3018 516896
rect 3054 512760 3110 512816
rect 3054 504600 3110 504656
rect 3330 497120 3386 497176
rect 3330 488960 3386 489016
rect 2870 476720 2926 476776
rect 2870 472640 2926 472696
rect 2962 468560 3018 468616
rect 3238 457000 3294 457056
rect 3330 452920 3386 452976
rect 3330 448840 3386 448896
rect 3330 440680 3386 440736
rect 2870 428440 2926 428496
rect 3238 400560 3294 400616
rect 2962 388320 3018 388376
rect 3146 384920 3202 384976
rect 3330 380840 3386 380896
rect 3330 376780 3386 376816
rect 3330 376760 3332 376780
rect 3332 376760 3384 376780
rect 3384 376760 3386 376780
rect 3330 372680 3386 372736
rect 3330 368600 3386 368656
rect 3330 364540 3386 364576
rect 3330 364520 3332 364540
rect 3332 364520 3384 364540
rect 3384 364520 3386 364540
rect 3330 360440 3386 360496
rect 3330 356360 3386 356416
rect 3238 352280 3294 352336
rect 3146 348880 3202 348936
rect 3330 344800 3386 344856
rect 3146 340720 3202 340776
rect 3330 336640 3386 336696
rect 3330 332596 3332 332616
rect 3332 332596 3384 332616
rect 3384 332596 3386 332616
rect 3330 332560 3386 332596
rect 3330 328500 3386 328536
rect 3330 328480 3332 328500
rect 3332 328480 3384 328500
rect 3384 328480 3386 328500
rect 3330 324400 3386 324456
rect 3146 320320 3202 320376
rect 3330 316240 3386 316296
rect 3330 308760 3386 308816
rect 3054 304680 3110 304736
rect 3146 300600 3202 300656
rect 3330 296520 3386 296576
rect 3146 292440 3202 292496
rect 3330 288360 3386 288416
rect 3330 284316 3332 284336
rect 3332 284316 3384 284336
rect 3384 284316 3386 284336
rect 3330 284280 3386 284316
rect 3330 280220 3386 280256
rect 3330 280200 3332 280220
rect 3332 280200 3384 280220
rect 3384 280200 3386 280220
rect 3146 272040 3202 272096
rect 3330 264560 3386 264616
rect 3054 260480 3110 260536
rect 3146 256400 3202 256456
rect 3146 252320 3202 252376
rect 3330 248240 3386 248296
rect 3146 244160 3202 244216
rect 3330 240100 3386 240136
rect 3330 240080 3332 240100
rect 3332 240080 3384 240100
rect 3384 240080 3386 240100
rect 3330 236020 3386 236056
rect 3330 236000 3332 236020
rect 3332 236000 3384 236020
rect 3384 236000 3386 236020
rect 3330 232600 3386 232656
rect 3330 228520 3386 228576
rect 3330 224440 3386 224496
rect 3238 220360 3294 220416
rect 3330 216280 3386 216336
rect 3514 601160 3570 601216
rect 3514 577360 3570 577416
rect 3514 552880 3570 552936
rect 3514 541320 3570 541376
rect 3514 529080 3570 529136
rect 3514 525000 3570 525056
rect 3514 508680 3570 508736
rect 3514 493040 3570 493096
rect 3514 484880 3570 484936
rect 3514 480800 3570 480856
rect 3514 465160 3570 465216
rect 3514 461080 3570 461136
rect 3514 444760 3570 444816
rect 3514 436600 3570 436656
rect 3514 432520 3570 432576
rect 3514 416880 3570 416936
rect 3514 412800 3570 412856
rect 3514 408720 3570 408776
rect 3514 404640 3570 404696
rect 3606 396480 3662 396536
rect 3514 199960 3570 200016
rect 3422 195880 3478 195936
rect 3422 192480 3478 192536
rect 3238 188400 3294 188456
rect 3146 184320 3202 184376
rect 3238 180240 3294 180296
rect 3238 172080 3294 172136
rect 3330 168000 3386 168056
rect 3054 163920 3110 163976
rect 3606 159840 3662 159896
rect 3514 155760 3570 155816
rect 3606 152360 3662 152416
rect 3146 144200 3202 144256
rect 2778 140120 2834 140176
rect 3514 136040 3570 136096
rect 3330 131960 3386 132016
rect 3422 127880 3478 127936
rect 3422 123800 3478 123856
rect 26882 199416 26938 199472
rect 48962 200640 49018 200696
rect 43442 199688 43498 199744
rect 60738 190304 60794 190360
rect 79322 200776 79378 200832
rect 84198 194520 84254 194576
rect 80794 191120 80850 191176
rect 89074 192888 89130 192944
rect 92478 227740 92480 227760
rect 92480 227740 92532 227760
rect 92532 227740 92534 227760
rect 92478 227704 92534 227740
rect 91098 195880 91154 195936
rect 93122 191664 93178 191720
rect 93306 190984 93362 191040
rect 93766 227704 93822 227760
rect 64142 145560 64198 145616
rect 3330 119720 3386 119776
rect 3330 112240 3386 112296
rect 3054 108160 3110 108216
rect 2962 104080 3018 104136
rect 2870 100000 2926 100056
rect 2962 95920 3018 95976
rect 3054 91840 3110 91896
rect 2870 76200 2926 76256
rect 3146 72120 3202 72176
rect 3146 36080 3202 36136
rect 3146 27920 3202 27976
rect 3514 116320 3570 116376
rect 3514 87760 3570 87816
rect 3514 83680 3570 83736
rect 3514 79636 3516 79656
rect 3516 79636 3568 79656
rect 3568 79636 3570 79656
rect 3514 79600 3570 79636
rect 3514 68040 3570 68096
rect 3514 59880 3570 59936
rect 3514 51720 3570 51776
rect 3514 47640 3570 47696
rect 3514 43560 3570 43616
rect 3514 39480 3570 39536
rect 3422 23840 3478 23896
rect 3146 19760 3202 19816
rect 3054 11600 3110 11656
rect 2962 7520 3018 7576
rect 2778 3440 2834 3496
rect 3330 15680 3386 15736
rect 94502 186088 94558 186144
rect 95146 76472 95202 76528
rect 96986 81912 97042 81968
rect 97078 71712 97134 71768
rect 97722 67360 97778 67416
rect 98734 200912 98790 200968
rect 98642 191256 98698 191312
rect 99838 148416 99894 148472
rect 99838 69536 99894 69592
rect 99286 67088 99342 67144
rect 102782 199552 102838 199608
rect 102874 196968 102930 197024
rect 101218 81776 101274 81832
rect 101494 80960 101550 81016
rect 102046 64776 102102 64832
rect 103150 68584 103206 68640
rect 104162 195744 104218 195800
rect 104346 192480 104402 192536
rect 103334 67496 103390 67552
rect 104530 77152 104586 77208
rect 104714 75792 104770 75848
rect 105542 195200 105598 195256
rect 105450 135904 105506 135960
rect 104806 67224 104862 67280
rect 105542 80824 105598 80880
rect 105634 79464 105690 79520
rect 106922 196832 106978 196888
rect 105818 71032 105874 71088
rect 106922 70216 106978 70272
rect 107106 69400 107162 69456
rect 107566 200640 107622 200696
rect 107566 200232 107622 200288
rect 109038 197240 109094 197296
rect 109866 75384 109922 75440
rect 110234 145832 110290 145888
rect 110418 190168 110474 190224
rect 111798 200912 111854 200968
rect 111798 200368 111854 200424
rect 112442 189896 112498 189952
rect 112534 145968 112590 146024
rect 112810 262384 112866 262440
rect 112442 72528 112498 72584
rect 113086 200368 113142 200424
rect 112994 189896 113050 189952
rect 112718 72392 112774 72448
rect 113638 142160 113694 142216
rect 112994 71168 113050 71224
rect 115386 262792 115442 262848
rect 115110 143248 115166 143304
rect 115018 142704 115074 142760
rect 116582 199144 116638 199200
rect 117318 193160 117374 193216
rect 116766 138624 116822 138680
rect 116674 81640 116730 81696
rect 117778 200640 117834 200696
rect 117686 142976 117742 143032
rect 117686 141888 117742 141944
rect 118054 192480 118110 192536
rect 119250 144880 119306 144936
rect 119066 142840 119122 142896
rect 118606 139304 118662 139360
rect 119342 138896 119398 138952
rect 119250 95104 119306 95160
rect 119434 89800 119490 89856
rect 119250 74840 119306 74896
rect 115478 66952 115534 67008
rect 119802 78512 119858 78568
rect 119802 72800 119858 72856
rect 120262 198600 120318 198656
rect 120262 197920 120318 197976
rect 120630 223488 120686 223544
rect 122562 259528 122618 259584
rect 126978 262792 127034 262848
rect 130382 263608 130438 263664
rect 141238 262384 141294 262440
rect 154486 262520 154542 262576
rect 166906 262384 166962 262440
rect 170586 263608 170642 263664
rect 171046 263608 171102 263664
rect 173070 263744 173126 263800
rect 171138 260072 171194 260128
rect 154026 259664 154082 259720
rect 184938 259936 184994 259992
rect 185858 259936 185914 259992
rect 187146 259528 187202 259584
rect 120998 223488 121054 223544
rect 131670 200504 131726 200560
rect 121274 198600 121330 198656
rect 120446 145696 120502 145752
rect 120722 80144 120778 80200
rect 120906 139304 120962 139360
rect 121734 138760 121790 138816
rect 121734 138488 121790 138544
rect 121734 138080 121790 138136
rect 121734 135904 121790 135960
rect 121734 89800 121790 89856
rect 129738 199960 129794 200016
rect 128358 199824 128414 199880
rect 122838 197784 122894 197840
rect 122470 197376 122526 197432
rect 122470 195880 122526 195936
rect 122838 195880 122894 195936
rect 122470 190440 122526 190496
rect 122746 189488 122802 189544
rect 122746 181464 122802 181520
rect 122746 180648 122802 180704
rect 122746 171128 122802 171184
rect 122746 170992 122802 171048
rect 122746 161472 122802 161528
rect 122746 161336 122802 161392
rect 122746 151816 122802 151872
rect 122746 151680 122802 151736
rect 122746 147600 122802 147656
rect 123482 197784 123538 197840
rect 123574 194248 123630 194304
rect 124954 199144 125010 199200
rect 124402 143248 124458 143304
rect 125598 148552 125654 148608
rect 125782 148416 125838 148472
rect 125230 144880 125286 144936
rect 126426 197920 126482 197976
rect 126794 197920 126850 197976
rect 126702 194384 126758 194440
rect 126610 178064 126666 178120
rect 124218 139576 124274 139632
rect 127990 181192 128046 181248
rect 128174 180784 128230 180840
rect 128542 193976 128598 194032
rect 129094 188944 129150 189000
rect 128726 181056 128782 181112
rect 130934 199144 130990 199200
rect 129646 196424 129702 196480
rect 129646 188944 129702 189000
rect 129186 180920 129242 180976
rect 129094 148688 129150 148744
rect 123574 139304 123630 139360
rect 124126 139304 124182 139360
rect 127622 139304 127678 139360
rect 129186 139304 129242 139360
rect 131118 185000 131174 185056
rect 131118 143112 131174 143168
rect 131762 199280 131818 199336
rect 177762 200368 177818 200424
rect 131854 198736 131910 198792
rect 132038 199144 132094 199200
rect 132130 198600 132186 198656
rect 131854 145968 131910 146024
rect 131210 141888 131266 141944
rect 132728 199824 132784 199880
rect 132498 199280 132554 199336
rect 133096 199824 133152 199880
rect 133142 199280 133198 199336
rect 133556 199824 133612 199880
rect 134108 199824 134164 199880
rect 134384 199824 134440 199880
rect 134752 199858 134808 199914
rect 133510 199280 133566 199336
rect 133510 199144 133566 199200
rect 133418 198736 133474 198792
rect 133510 195880 133566 195936
rect 133786 199144 133842 199200
rect 133786 194248 133842 194304
rect 134154 199280 134210 199336
rect 134338 198736 134394 198792
rect 134798 198736 134854 198792
rect 134982 199280 135038 199336
rect 135074 198736 135130 198792
rect 135074 197104 135130 197160
rect 134798 193840 134854 193896
rect 134522 190712 134578 190768
rect 136224 199858 136280 199914
rect 135626 198736 135682 198792
rect 135534 198328 135590 198384
rect 135258 193976 135314 194032
rect 134522 178880 134578 178936
rect 135994 199280 136050 199336
rect 135994 193024 136050 193080
rect 136178 198464 136234 198520
rect 136546 199280 136602 199336
rect 136362 195880 136418 195936
rect 136730 199280 136786 199336
rect 136822 196016 136878 196072
rect 137006 198464 137062 198520
rect 136914 192752 136970 192808
rect 137328 199858 137384 199914
rect 137374 199280 137430 199336
rect 137282 199144 137338 199200
rect 137190 198328 137246 198384
rect 137880 199858 137936 199914
rect 136546 176568 136602 176624
rect 135350 145832 135406 145888
rect 136822 142160 136878 142216
rect 137650 198736 137706 198792
rect 137834 199280 137890 199336
rect 137834 199144 137890 199200
rect 138432 199858 138488 199914
rect 138800 199858 138856 199914
rect 139260 199858 139316 199914
rect 138110 199280 138166 199336
rect 137926 194384 137982 194440
rect 138386 198600 138442 198656
rect 138294 198192 138350 198248
rect 138570 196696 138626 196752
rect 138478 196288 138534 196344
rect 138018 184864 138074 184920
rect 138018 181328 138074 181384
rect 137650 174936 137706 174992
rect 137650 174664 137706 174720
rect 138754 198736 138810 198792
rect 138754 198056 138810 198112
rect 138662 195880 138718 195936
rect 138570 189760 138626 189816
rect 137466 144200 137522 144256
rect 137282 140528 137338 140584
rect 138846 191120 138902 191176
rect 139122 197784 139178 197840
rect 139536 199858 139592 199914
rect 139904 199858 139960 199914
rect 140272 199858 140328 199914
rect 140640 199858 140696 199914
rect 140318 199144 140374 199200
rect 140226 198056 140282 198112
rect 139582 197376 139638 197432
rect 139214 197104 139270 197160
rect 138938 188944 138994 189000
rect 138938 188672 138994 188728
rect 139490 190168 139546 190224
rect 139490 189760 139546 189816
rect 140226 197512 140282 197568
rect 140134 190168 140190 190224
rect 140502 199144 140558 199200
rect 142204 199858 142260 199914
rect 142480 199858 142536 199914
rect 142848 199858 142904 199914
rect 141422 195608 141478 195664
rect 141698 198736 141754 198792
rect 142250 198500 142252 198520
rect 142252 198500 142304 198520
rect 142304 198500 142306 198520
rect 142250 198464 142306 198500
rect 141974 197240 142030 197296
rect 142618 198600 142674 198656
rect 142526 197240 142582 197296
rect 142710 198056 142766 198112
rect 141974 194112 142030 194168
rect 142618 189624 142674 189680
rect 140778 176568 140834 176624
rect 140870 175208 140926 175264
rect 143078 196424 143134 196480
rect 143078 186904 143134 186960
rect 144320 199858 144376 199914
rect 144596 199858 144652 199914
rect 143906 198192 143962 198248
rect 145056 199858 145112 199914
rect 145608 199858 145664 199914
rect 146160 199858 146216 199914
rect 144366 199144 144422 199200
rect 144366 198736 144422 198792
rect 144274 198600 144330 198656
rect 144734 198872 144790 198928
rect 144550 198056 144606 198112
rect 144458 189760 144514 189816
rect 145102 198464 145158 198520
rect 145286 197804 145342 197840
rect 145286 197784 145288 197804
rect 145288 197784 145340 197804
rect 145340 197784 145342 197804
rect 144918 187448 144974 187504
rect 145102 187040 145158 187096
rect 145378 186224 145434 186280
rect 145654 187448 145710 187504
rect 145930 195472 145986 195528
rect 146114 198056 146170 198112
rect 146390 199144 146446 199200
rect 145562 186224 145618 186280
rect 145746 186224 145802 186280
rect 145562 185544 145618 185600
rect 146804 199858 146860 199914
rect 146482 195336 146538 195392
rect 147402 199144 147458 199200
rect 147816 199858 147872 199914
rect 148276 199858 148332 199914
rect 148552 199858 148608 199914
rect 147494 199008 147550 199064
rect 147494 195880 147550 195936
rect 147494 195472 147550 195528
rect 147862 197376 147918 197432
rect 148920 199858 148976 199914
rect 149104 199858 149160 199914
rect 148322 192072 148378 192128
rect 148230 190440 148286 190496
rect 148046 184456 148102 184512
rect 145930 142976 145986 143032
rect 146574 140392 146630 140448
rect 130842 139440 130898 139496
rect 148874 198464 148930 198520
rect 149656 199858 149712 199914
rect 149058 196560 149114 196616
rect 149518 198736 149574 198792
rect 148966 187584 149022 187640
rect 148414 141616 148470 141672
rect 150208 199858 150264 199914
rect 149794 198872 149850 198928
rect 149978 198736 150034 198792
rect 150162 199144 150218 199200
rect 150162 199008 150218 199064
rect 149610 190032 149666 190088
rect 149242 142704 149298 142760
rect 150346 199144 150402 199200
rect 150346 192072 150402 192128
rect 151128 199858 151184 199914
rect 150622 195200 150678 195256
rect 149794 144064 149850 144120
rect 149702 141752 149758 141808
rect 151772 199858 151828 199914
rect 152048 199858 152104 199914
rect 151266 199280 151322 199336
rect 151174 198056 151230 198112
rect 151726 199008 151782 199064
rect 151726 198328 151782 198384
rect 152416 199858 152472 199914
rect 153152 199858 153208 199914
rect 153520 199858 153576 199914
rect 152278 199008 152334 199064
rect 152278 198736 152334 198792
rect 152002 196288 152058 196344
rect 151726 188944 151782 189000
rect 151726 188400 151782 188456
rect 152278 145696 152334 145752
rect 152738 196424 152794 196480
rect 153014 199280 153070 199336
rect 153106 198756 153162 198792
rect 153106 198736 153108 198756
rect 153108 198736 153160 198756
rect 153160 198736 153162 198756
rect 154256 199858 154312 199914
rect 153382 199280 153438 199336
rect 153474 196016 153530 196072
rect 152370 141480 152426 141536
rect 153750 198736 153806 198792
rect 153658 196152 153714 196208
rect 154808 199858 154864 199914
rect 153934 145696 153990 145752
rect 153382 142840 153438 142896
rect 154486 188400 154542 188456
rect 154854 198736 154910 198792
rect 154854 183096 154910 183152
rect 155406 190304 155462 190360
rect 155958 198056 156014 198112
rect 155958 195472 156014 195528
rect 156832 199858 156888 199914
rect 156234 198192 156290 198248
rect 156050 179016 156106 179072
rect 157844 199858 157900 199914
rect 156970 199280 157026 199336
rect 156970 199144 157026 199200
rect 156878 198328 156934 198384
rect 157062 196152 157118 196208
rect 157338 196016 157394 196072
rect 158856 199858 158912 199914
rect 159040 199858 159096 199914
rect 157798 199144 157854 199200
rect 157890 196424 157946 196480
rect 156510 142704 156566 142760
rect 155406 141480 155462 141536
rect 159408 199858 159464 199914
rect 158902 198736 158958 198792
rect 159086 198736 159142 198792
rect 158994 196016 159050 196072
rect 158626 190984 158682 191040
rect 159546 196016 159602 196072
rect 159546 190984 159602 191040
rect 160236 199858 160292 199914
rect 159730 182824 159786 182880
rect 161248 199858 161304 199914
rect 160558 199280 160614 199336
rect 161294 199552 161350 199608
rect 161708 199858 161764 199914
rect 161294 199280 161350 199336
rect 161110 196016 161166 196072
rect 161294 196424 161350 196480
rect 160742 189760 160798 189816
rect 160558 186904 160614 186960
rect 161662 199552 161718 199608
rect 162260 199858 162316 199914
rect 161386 190984 161442 191040
rect 162122 199280 162178 199336
rect 162490 199552 162546 199608
rect 162490 199280 162546 199336
rect 162490 193160 162546 193216
rect 162904 199858 162960 199914
rect 162950 199280 163006 199336
rect 162858 196424 162914 196480
rect 162490 179152 162546 179208
rect 163134 196016 163190 196072
rect 163042 195064 163098 195120
rect 163916 199858 163972 199914
rect 164192 199858 164248 199914
rect 164376 199858 164432 199914
rect 164560 199824 164616 199880
rect 163778 199144 163834 199200
rect 163042 178608 163098 178664
rect 163962 197784 164018 197840
rect 164054 196288 164110 196344
rect 163870 142840 163926 142896
rect 163686 140256 163742 140312
rect 164422 199688 164478 199744
rect 164330 196016 164386 196072
rect 164606 199688 164662 199744
rect 165112 199824 165168 199880
rect 165296 199824 165352 199880
rect 164238 190848 164294 190904
rect 165066 198056 165122 198112
rect 165158 196152 165214 196208
rect 165618 199280 165674 199336
rect 166768 199824 166824 199880
rect 165802 196288 165858 196344
rect 166722 198464 166778 198520
rect 167412 199824 167468 199880
rect 168240 199824 168296 199880
rect 167734 199416 167790 199472
rect 167826 198736 167882 198792
rect 167458 189080 167514 189136
rect 167918 194384 167974 194440
rect 168792 199824 168848 199880
rect 168194 198056 168250 198112
rect 168194 197920 168250 197976
rect 168102 196152 168158 196208
rect 168746 199688 168802 199744
rect 168378 199552 168434 199608
rect 168746 199588 168748 199608
rect 168748 199588 168800 199608
rect 168800 199588 168802 199608
rect 168746 199552 168802 199588
rect 168930 199552 168986 199608
rect 168838 199144 168894 199200
rect 168654 198736 168710 198792
rect 168378 195336 168434 195392
rect 168378 186088 168434 186144
rect 168838 196288 168894 196344
rect 169436 199824 169492 199880
rect 169712 199824 169768 199880
rect 169298 199416 169354 199472
rect 168470 148416 168526 148472
rect 169206 180240 169262 180296
rect 169666 199144 169722 199200
rect 169850 199552 169906 199608
rect 170034 199416 170090 199472
rect 169758 198328 169814 198384
rect 169574 196852 169630 196888
rect 169574 196832 169576 196852
rect 169576 196832 169628 196852
rect 169628 196832 169630 196852
rect 169942 196968 169998 197024
rect 170448 199858 170504 199914
rect 170724 199858 170780 199914
rect 169942 192888 169998 192944
rect 170218 187720 170274 187776
rect 170494 195744 170550 195800
rect 170586 195336 170642 195392
rect 170770 195472 170826 195528
rect 171368 199858 171424 199914
rect 171414 197648 171470 197704
rect 170862 193296 170918 193352
rect 170770 191664 170826 191720
rect 171598 199144 171654 199200
rect 171690 188536 171746 188592
rect 170586 144064 170642 144120
rect 171046 142976 171102 143032
rect 172150 194112 172206 194168
rect 172748 199858 172804 199914
rect 172426 198600 172482 198656
rect 173208 199858 173264 199914
rect 173944 199858 174000 199914
rect 174128 199858 174184 199914
rect 173622 199724 173624 199744
rect 173624 199724 173676 199744
rect 173676 199724 173678 199744
rect 172794 198600 172850 198656
rect 173622 199688 173678 199724
rect 174082 199688 174138 199744
rect 173530 199552 173586 199608
rect 173530 198600 173586 198656
rect 173622 196832 173678 196888
rect 174082 198600 174138 198656
rect 174266 196832 174322 196888
rect 173806 192480 173862 192536
rect 174772 199824 174828 199880
rect 175048 199858 175104 199914
rect 175002 199688 175058 199744
rect 175324 199824 175380 199880
rect 174910 199144 174966 199200
rect 174818 198056 174874 198112
rect 174450 196968 174506 197024
rect 175554 198600 175610 198656
rect 173714 143112 173770 143168
rect 173438 140528 173494 140584
rect 176106 199552 176162 199608
rect 176796 199824 176852 199880
rect 177072 199824 177128 199880
rect 176842 199588 176844 199608
rect 176844 199588 176896 199608
rect 176896 199588 176898 199608
rect 176842 199552 176898 199588
rect 176842 199144 176898 199200
rect 175922 193976 175978 194032
rect 176658 196016 176714 196072
rect 177302 194656 177358 194712
rect 176474 180240 176530 180296
rect 176382 144336 176438 144392
rect 177670 198464 177726 198520
rect 178130 199552 178186 199608
rect 177946 146920 178002 146976
rect 177946 144200 178002 144256
rect 178406 200504 178462 200560
rect 179326 199960 179382 200016
rect 179418 197920 179474 197976
rect 179326 196832 179382 196888
rect 179142 192616 179198 192672
rect 179418 185680 179474 185736
rect 178774 140392 178830 140448
rect 180706 196696 180762 196752
rect 180706 186904 180762 186960
rect 180706 141616 180762 141672
rect 187606 200640 187662 200696
rect 182822 199280 182878 199336
rect 181810 199144 181866 199200
rect 182270 198056 182326 198112
rect 181074 194384 181130 194440
rect 182086 194384 182142 194440
rect 181994 189624 182050 189680
rect 180982 141344 181038 141400
rect 179602 140120 179658 140176
rect 179510 139984 179566 140040
rect 181994 140120 182050 140176
rect 182638 195744 182694 195800
rect 183282 190032 183338 190088
rect 182086 139984 182142 140040
rect 183374 141752 183430 141808
rect 184294 145832 184350 145888
rect 183190 139440 183246 139496
rect 184846 141344 184902 141400
rect 186042 184592 186098 184648
rect 186042 145968 186098 146024
rect 185950 143248 186006 143304
rect 185950 142432 186006 142488
rect 186226 142432 186282 142488
rect 186134 141888 186190 141944
rect 186042 140528 186098 140584
rect 186870 143384 186926 143440
rect 186318 140664 186374 140720
rect 130842 139304 130898 139360
rect 146666 139304 146722 139360
rect 170678 139304 170734 139360
rect 176474 139304 176530 139360
rect 183098 139304 183154 139360
rect 184018 139304 184074 139360
rect 187698 145560 187754 145616
rect 188342 179288 188398 179344
rect 187330 139576 187386 139632
rect 186502 139440 186558 139496
rect 187974 139440 188030 139496
rect 131762 80688 131818 80744
rect 123482 80552 123538 80608
rect 122378 80280 122434 80336
rect 122378 74432 122434 74488
rect 126334 79872 126390 79928
rect 126334 77968 126390 78024
rect 129186 78240 129242 78296
rect 132222 80688 132278 80744
rect 177762 80552 177818 80608
rect 131946 80280 132002 80336
rect 131854 80008 131910 80064
rect 132130 79736 132186 79792
rect 133096 79872 133152 79928
rect 133464 79872 133520 79928
rect 133648 79872 133704 79928
rect 134016 79872 134072 79928
rect 132866 78376 132922 78432
rect 132774 67088 132830 67144
rect 133142 79600 133198 79656
rect 133142 78648 133198 78704
rect 133050 78512 133106 78568
rect 133418 79736 133474 79792
rect 133326 75112 133382 75168
rect 133970 79736 134026 79792
rect 134384 79906 134440 79962
rect 134062 79600 134118 79656
rect 134752 79906 134808 79962
rect 134614 79756 134670 79792
rect 134614 79736 134616 79756
rect 134616 79736 134668 79756
rect 134668 79736 134670 79756
rect 134614 79600 134670 79656
rect 134982 78512 135038 78568
rect 134982 77968 135038 78024
rect 135074 76472 135130 76528
rect 135580 79906 135636 79962
rect 135258 77832 135314 77888
rect 135856 79906 135912 79962
rect 136132 79872 136188 79928
rect 136776 79906 136832 79962
rect 135718 78104 135774 78160
rect 135534 76200 135590 76256
rect 136178 79600 136234 79656
rect 136822 79736 136878 79792
rect 137144 79872 137200 79928
rect 137328 79906 137384 79962
rect 136822 79636 136824 79656
rect 136824 79636 136876 79656
rect 136876 79636 136878 79656
rect 136822 79600 136878 79636
rect 136638 76880 136694 76936
rect 137190 79736 137246 79792
rect 137006 76744 137062 76800
rect 137466 79600 137522 79656
rect 137190 77288 137246 77344
rect 137098 75248 137154 75304
rect 137374 79192 137430 79248
rect 137558 79328 137614 79384
rect 138064 79906 138120 79962
rect 138432 79872 138488 79928
rect 138892 79906 138948 79962
rect 138294 79464 138350 79520
rect 138110 77968 138166 78024
rect 138386 76472 138442 76528
rect 138294 67224 138350 67280
rect 139536 79872 139592 79928
rect 139720 79872 139776 79928
rect 139858 79756 139914 79792
rect 140548 79872 140604 79928
rect 140824 79872 140880 79928
rect 141100 79872 141156 79928
rect 141284 79872 141340 79928
rect 138662 77016 138718 77072
rect 139122 78512 139178 78568
rect 139122 78240 139178 78296
rect 139858 79736 139860 79756
rect 139860 79736 139912 79756
rect 139912 79736 139914 79756
rect 139582 78512 139638 78568
rect 140502 79600 140558 79656
rect 140042 73752 140098 73808
rect 140502 77152 140558 77208
rect 140962 79736 141018 79792
rect 140870 79328 140926 79384
rect 141238 79600 141294 79656
rect 141146 76608 141202 76664
rect 141928 79872 141984 79928
rect 141514 79464 141570 79520
rect 141698 79620 141754 79656
rect 142296 79872 142352 79928
rect 141698 79600 141700 79620
rect 141700 79600 141752 79620
rect 141752 79600 141754 79620
rect 141698 79464 141754 79520
rect 141422 78376 141478 78432
rect 141330 77696 141386 77752
rect 141422 76608 141478 76664
rect 141238 66000 141294 66056
rect 141882 78512 141938 78568
rect 142756 79906 142812 79962
rect 143032 79906 143088 79962
rect 142158 78648 142214 78704
rect 142066 77696 142122 77752
rect 141974 70352 142030 70408
rect 141974 69672 142030 69728
rect 141606 64640 141662 64696
rect 142894 78648 142950 78704
rect 142802 78512 142858 78568
rect 143538 78648 143594 78704
rect 143170 75384 143226 75440
rect 144228 79872 144284 79928
rect 144504 79906 144560 79962
rect 144872 79906 144928 79962
rect 144734 79772 144742 79792
rect 144742 79772 144790 79792
rect 143814 79600 143870 79656
rect 144182 79600 144238 79656
rect 144182 74296 144238 74352
rect 143998 72664 144054 72720
rect 144734 79736 144790 79772
rect 145332 79872 145388 79928
rect 144458 71168 144514 71224
rect 144826 76608 144882 76664
rect 143906 69808 143962 69864
rect 145286 75792 145342 75848
rect 145286 75112 145342 75168
rect 145976 79906 146032 79962
rect 146252 79906 146308 79962
rect 146528 79906 146584 79962
rect 146712 79838 146768 79894
rect 147080 79872 147136 79928
rect 147724 79872 147780 79928
rect 145010 71576 145066 71632
rect 145838 78104 145894 78160
rect 146574 79600 146630 79656
rect 145746 67496 145802 67552
rect 146482 76608 146538 76664
rect 146298 71712 146354 71768
rect 146942 73888 146998 73944
rect 146758 67496 146814 67552
rect 147402 75520 147458 75576
rect 147126 67496 147182 67552
rect 147126 66952 147182 67008
rect 148184 79906 148240 79962
rect 148000 79838 148056 79894
rect 148368 79906 148424 79962
rect 148736 79872 148792 79928
rect 148230 79600 148286 79656
rect 148414 79600 148470 79656
rect 148322 79056 148378 79112
rect 147678 74432 147734 74488
rect 149288 79770 149344 79826
rect 149426 79600 149482 79656
rect 149334 79464 149390 79520
rect 149610 77968 149666 78024
rect 149794 74976 149850 75032
rect 149978 77696 150034 77752
rect 150162 77560 150218 77616
rect 150576 79906 150632 79962
rect 150944 79906 151000 79962
rect 151496 79906 151552 79962
rect 150622 79464 150678 79520
rect 150898 79600 150954 79656
rect 149886 66136 149942 66192
rect 151082 76336 151138 76392
rect 151450 79600 151506 79656
rect 151542 77832 151598 77888
rect 152324 79872 152380 79928
rect 152508 79872 152564 79928
rect 152002 75384 152058 75440
rect 151450 73616 151506 73672
rect 152186 79464 152242 79520
rect 153152 79906 153208 79962
rect 152554 79328 152610 79384
rect 152462 75928 152518 75984
rect 152830 77968 152886 78024
rect 153980 79906 154036 79962
rect 154164 79872 154220 79928
rect 153796 79736 153852 79792
rect 153750 79600 153806 79656
rect 153934 79600 153990 79656
rect 153842 75792 153898 75848
rect 153658 74160 153714 74216
rect 153934 73888 153990 73944
rect 154716 79906 154772 79962
rect 154900 79906 154956 79962
rect 155084 79872 155140 79928
rect 155360 79872 155416 79928
rect 154670 79600 154726 79656
rect 155222 79736 155278 79792
rect 154578 78512 154634 78568
rect 154670 75928 154726 75984
rect 154854 78512 154910 78568
rect 155314 75928 155370 75984
rect 156096 79906 156152 79962
rect 155728 79838 155784 79894
rect 156280 79872 156336 79928
rect 155682 79600 155738 79656
rect 155498 79328 155554 79384
rect 155498 77832 155554 77888
rect 156050 79600 156106 79656
rect 156142 76608 156198 76664
rect 156234 76336 156290 76392
rect 157292 79906 157348 79962
rect 157752 79872 157808 79928
rect 157016 79824 157072 79826
rect 157016 79772 157018 79824
rect 157018 79772 157070 79824
rect 157070 79772 157072 79824
rect 157016 79770 157072 79772
rect 155130 69536 155186 69592
rect 154946 65728 155002 65784
rect 157936 79906 157992 79962
rect 157982 79600 158038 79656
rect 158672 79872 158728 79928
rect 159592 79906 159648 79962
rect 158626 77696 158682 77752
rect 158994 79600 159050 79656
rect 159454 78920 159510 78976
rect 159776 79906 159832 79962
rect 160144 79906 160200 79962
rect 160328 79872 160384 79928
rect 160604 79872 160660 79928
rect 160788 79906 160844 79962
rect 161064 79906 161120 79962
rect 161340 79906 161396 79962
rect 159914 79600 159970 79656
rect 159822 74976 159878 75032
rect 160190 79600 160246 79656
rect 159086 67360 159142 67416
rect 161018 79736 161074 79792
rect 161800 79906 161856 79962
rect 161984 79906 162040 79962
rect 160650 77152 160706 77208
rect 161018 76744 161074 76800
rect 160466 73616 160522 73672
rect 161294 79600 161350 79656
rect 161846 79736 161902 79792
rect 161478 74296 161534 74352
rect 161294 65728 161350 65784
rect 161294 65456 161350 65512
rect 161754 78512 161810 78568
rect 162122 79736 162178 79792
rect 161938 79600 161994 79656
rect 162536 79906 162592 79962
rect 162720 79906 162776 79962
rect 162904 79872 162960 79928
rect 163272 79872 163328 79928
rect 163088 79736 163144 79792
rect 163502 79736 163558 79792
rect 162766 79600 162822 79656
rect 162766 75248 162822 75304
rect 162766 72936 162822 72992
rect 161938 68448 161994 68504
rect 161662 64504 161718 64560
rect 163318 79600 163374 79656
rect 163042 79328 163098 79384
rect 163134 79056 163190 79112
rect 164008 79906 164064 79962
rect 164192 79906 164248 79962
rect 163732 79736 163788 79792
rect 164284 79736 164340 79792
rect 164652 79906 164708 79962
rect 164928 79906 164984 79962
rect 163870 72800 163926 72856
rect 164238 79464 164294 79520
rect 164146 73888 164202 73944
rect 163226 68584 163282 68640
rect 164606 79600 164662 79656
rect 165480 79906 165536 79962
rect 165664 79906 165720 79962
rect 166216 79906 166272 79962
rect 166584 79906 166640 79962
rect 164882 72664 164938 72720
rect 165342 72392 165398 72448
rect 165802 78920 165858 78976
rect 166170 79736 166226 79792
rect 166860 79770 166916 79826
rect 167136 79906 167192 79962
rect 166078 78376 166134 78432
rect 166170 74024 166226 74080
rect 166722 79464 166778 79520
rect 166814 78784 166870 78840
rect 166170 73752 166226 73808
rect 167550 79600 167606 79656
rect 168056 79906 168112 79962
rect 168240 79838 168296 79894
rect 168010 78920 168066 78976
rect 167918 76880 167974 76936
rect 168194 79600 168250 79656
rect 168608 79736 168664 79792
rect 168378 79600 168434 79656
rect 169022 76744 169078 76800
rect 169528 79906 169584 79962
rect 169896 79872 169952 79928
rect 170172 79872 170228 79928
rect 169758 79056 169814 79112
rect 169390 76744 169446 76800
rect 169758 75928 169814 75984
rect 169666 75792 169722 75848
rect 170816 79906 170872 79962
rect 170678 78376 170734 78432
rect 171000 79736 171056 79792
rect 170862 78240 170918 78296
rect 171644 79906 171700 79962
rect 170954 77968 171010 78024
rect 170218 70216 170274 70272
rect 170862 72528 170918 72584
rect 171598 79600 171654 79656
rect 172472 79906 172528 79962
rect 172656 79872 172712 79928
rect 172012 79736 172068 79792
rect 172610 79772 172618 79792
rect 172618 79772 172666 79792
rect 171874 78920 171930 78976
rect 172610 79736 172666 79772
rect 173116 79872 173172 79928
rect 173760 79906 173816 79962
rect 173944 79906 174000 79962
rect 174036 79772 174038 79792
rect 174038 79772 174090 79792
rect 174090 79772 174092 79792
rect 172426 78512 172482 78568
rect 172610 78512 172666 78568
rect 172426 76472 172482 76528
rect 171966 71168 172022 71224
rect 171414 69944 171470 70000
rect 174036 79736 174092 79772
rect 173162 79600 173218 79656
rect 173254 78376 173310 78432
rect 173806 79600 173862 79656
rect 173714 77832 173770 77888
rect 174680 79872 174736 79928
rect 175232 79906 175288 79962
rect 173990 76608 174046 76664
rect 173622 70080 173678 70136
rect 175002 79600 175058 79656
rect 175278 78920 175334 78976
rect 175968 79872 176024 79928
rect 176612 79906 176668 79962
rect 175554 77832 175610 77888
rect 175922 78512 175978 78568
rect 176888 79906 176944 79962
rect 177946 80028 178002 80064
rect 177946 80008 177948 80028
rect 177948 80008 178000 80028
rect 178000 80008 178002 80028
rect 177440 79872 177496 79928
rect 176014 76200 176070 76256
rect 176474 78512 176530 78568
rect 176566 74976 176622 75032
rect 178590 80416 178646 80472
rect 181626 79872 181682 79928
rect 181534 79736 181590 79792
rect 178314 74160 178370 74216
rect 181626 78240 181682 78296
rect 180706 77968 180762 78024
rect 180706 77152 180762 77208
rect 180614 77016 180670 77072
rect 180338 76880 180394 76936
rect 181442 77152 181498 77208
rect 182914 77832 182970 77888
rect 187054 80416 187110 80472
rect 184938 80144 184994 80200
rect 186962 79328 187018 79384
rect 187054 73072 187110 73128
rect 186962 66952 187018 67008
rect 188710 133728 188766 133784
rect 188894 104080 188950 104136
rect 188986 77696 189042 77752
rect 189354 69536 189410 69592
rect 189906 263064 189962 263120
rect 189906 262520 189962 262576
rect 189814 199008 189870 199064
rect 189998 260072 190054 260128
rect 189998 198192 190054 198248
rect 190090 88304 190146 88360
rect 189906 81368 189962 81424
rect 190550 142704 190606 142760
rect 190642 137944 190698 138000
rect 191286 140120 191342 140176
rect 191102 138760 191158 138816
rect 191010 136584 191066 136640
rect 191286 80960 191342 81016
rect 191286 80824 191342 80880
rect 191286 80552 191342 80608
rect 193218 197648 193274 197704
rect 192666 91840 192722 91896
rect 193310 142840 193366 142896
rect 193310 141752 193366 141808
rect 193586 77152 193642 77208
rect 194230 141888 194286 141944
rect 193678 73888 193734 73944
rect 194506 77152 194562 77208
rect 194690 143248 194746 143304
rect 194874 141616 194930 141672
rect 195058 140528 195114 140584
rect 195242 141344 195298 141400
rect 195334 139032 195390 139088
rect 195518 144336 195574 144392
rect 195334 77968 195390 78024
rect 196070 72528 196126 72584
rect 196346 137400 196402 137456
rect 197358 195064 197414 195120
rect 197082 190848 197138 190904
rect 197358 190848 197414 190904
rect 197082 190576 197138 190632
rect 196806 134408 196862 134464
rect 196806 83408 196862 83464
rect 191930 34448 191986 34504
rect 198830 262928 198886 262984
rect 198830 262384 198886 262440
rect 199106 262384 199162 262440
rect 198462 144200 198518 144256
rect 198186 135904 198242 135960
rect 199106 137264 199162 137320
rect 199566 144064 199622 144120
rect 200118 74024 200174 74080
rect 200486 195608 200542 195664
rect 200486 187312 200542 187368
rect 201774 190848 201830 190904
rect 202234 148280 202290 148336
rect 201590 64232 201646 64288
rect 202326 138896 202382 138952
rect 203154 148416 203210 148472
rect 202970 69672 203026 69728
rect 204626 184320 204682 184376
rect 204350 69944 204406 70000
rect 208398 220904 208454 220960
rect 207018 196968 207074 197024
rect 207018 196696 207074 196752
rect 207202 196696 207258 196752
rect 204994 81912 205050 81968
rect 204810 70216 204866 70272
rect 204626 65728 204682 65784
rect 206374 81640 206430 81696
rect 207202 78376 207258 78432
rect 207018 74024 207074 74080
rect 207110 71304 207166 71360
rect 207570 185952 207626 186008
rect 209318 202136 209374 202192
rect 208490 201456 208546 201512
rect 209318 201456 209374 201512
rect 208490 67088 208546 67144
rect 208858 185544 208914 185600
rect 208858 74160 208914 74216
rect 208674 67224 208730 67280
rect 209962 77832 210018 77888
rect 211618 195200 211674 195256
rect 211618 79056 211674 79112
rect 212906 178744 212962 178800
rect 212998 80824 213054 80880
rect 212906 75520 212962 75576
rect 217230 199552 217286 199608
rect 216678 199416 216734 199472
rect 215298 195744 215354 195800
rect 214654 195608 214710 195664
rect 214470 195336 214526 195392
rect 214470 76472 214526 76528
rect 215298 195472 215354 195528
rect 215482 195472 215538 195528
rect 215298 192752 215354 192808
rect 214746 77288 214802 77344
rect 214010 64776 214066 64832
rect 215390 189488 215446 189544
rect 215574 192616 215630 192672
rect 215666 190304 215722 190360
rect 215574 76200 215630 76256
rect 217046 198736 217102 198792
rect 217230 198736 217286 198792
rect 216770 182960 216826 183016
rect 216678 74840 216734 74896
rect 217138 193840 217194 193896
rect 217046 82184 217102 82240
rect 217414 82048 217470 82104
rect 218242 196832 218298 196888
rect 219622 191392 219678 191448
rect 218242 78920 218298 78976
rect 216954 71440 217010 71496
rect 218150 68856 218206 68912
rect 218426 184456 218482 184512
rect 219530 183504 219586 183560
rect 219438 181600 219494 181656
rect 218426 78784 218482 78840
rect 218334 71712 218390 71768
rect 218242 66136 218298 66192
rect 216770 66000 216826 66056
rect 215298 64640 215354 64696
rect 220818 190848 220874 190904
rect 220174 183504 220230 183560
rect 219806 183232 219862 183288
rect 219714 181328 219770 181384
rect 220174 182960 220230 183016
rect 220082 181464 220138 181520
rect 220082 80688 220138 80744
rect 219806 75656 219862 75712
rect 219530 71576 219586 71632
rect 219438 67496 219494 67552
rect 220910 77016 220966 77072
rect 231858 191664 231914 191720
rect 239402 199552 239458 199608
rect 260102 190304 260158 190360
rect 266358 190168 266414 190224
rect 305642 180376 305698 180432
rect 235998 179016 236054 179072
rect 221186 178880 221242 178936
rect 221094 65864 221150 65920
rect 333978 197104 334034 197160
rect 342258 192752 342314 192808
rect 376758 195608 376814 195664
rect 377402 191392 377458 191448
rect 391938 194384 391994 194440
rect 422298 200776 422354 200832
rect 431222 190032 431278 190088
rect 455418 188672 455474 188728
rect 452658 186904 452714 186960
rect 436098 184592 436154 184648
rect 459558 178880 459614 178936
rect 463698 178744 463754 178800
rect 483018 263064 483074 263120
rect 494058 191256 494114 191312
rect 489918 187312 489974 187368
rect 485778 183368 485834 183424
rect 476762 177656 476818 177712
rect 381542 174936 381598 174992
rect 514022 200640 514078 200696
rect 516138 199416 516194 199472
rect 524418 188808 524474 188864
rect 511998 184456 512054 184512
rect 535458 181600 535514 181656
rect 546498 262792 546554 262848
rect 544382 199280 544438 199336
rect 543738 183232 543794 183288
rect 543002 177928 543058 177984
rect 221186 63280 221242 63336
rect 548522 184320 548578 184376
rect 552662 182824 552718 182880
rect 554042 184864 554098 184920
rect 548614 180240 548670 180296
rect 554134 177792 554190 177848
rect 556894 193024 556950 193080
rect 558182 202136 558238 202192
rect 558366 197240 558422 197296
rect 558274 184728 558330 184784
rect 560942 185544 560998 185600
rect 561126 196696 561182 196752
rect 561034 184184 561090 184240
rect 561678 189896 561734 189952
rect 563794 188944 563850 189000
rect 566554 196832 566610 196888
rect 566646 187448 566702 187504
rect 567934 186224 567990 186280
rect 580170 702500 580226 702536
rect 580170 702480 580172 702500
rect 580172 702480 580224 702500
rect 580224 702480 580226 702500
rect 580170 698400 580226 698456
rect 580170 694320 580226 694376
rect 580170 690240 580226 690296
rect 579802 686160 579858 686216
rect 569958 262928 570014 262984
rect 570602 196560 570658 196616
rect 571982 194520 572038 194576
rect 574742 195880 574798 195936
rect 574926 192616 574982 192672
rect 574834 189624 574890 189680
rect 573362 183096 573418 183152
rect 576214 192344 576270 192400
rect 576398 259528 576454 259584
rect 577502 195336 577558 195392
rect 577778 195472 577834 195528
rect 576306 191120 576362 191176
rect 577870 189760 577926 189816
rect 576122 182960 576178 183016
rect 570694 181464 570750 181520
rect 580170 682080 580226 682136
rect 580170 678000 580226 678056
rect 580170 673920 580226 673976
rect 580170 669840 580226 669896
rect 580170 662360 580226 662416
rect 580170 658300 580226 658336
rect 580170 658280 580172 658300
rect 580172 658280 580224 658300
rect 580224 658280 580226 658300
rect 580170 654200 580226 654256
rect 580170 646040 580226 646096
rect 580170 641960 580226 642016
rect 580170 626320 580226 626376
rect 579802 622240 579858 622296
rect 580170 605920 580226 605976
rect 580170 601840 580226 601896
rect 580354 597760 580410 597816
rect 580170 589600 580226 589656
rect 578882 586200 578938 586256
rect 580170 569880 580226 569936
rect 580170 565836 580172 565856
rect 580172 565836 580224 565856
rect 580224 565836 580226 565856
rect 580170 565800 580226 565836
rect 580170 553560 580226 553616
rect 580170 549480 580226 549536
rect 579894 546080 579950 546136
rect 580170 542000 580226 542056
rect 580170 537920 580226 537976
rect 579802 529760 579858 529816
rect 580170 525680 580226 525736
rect 580170 521600 580226 521656
rect 580170 510040 580226 510096
rect 580078 505960 580134 506016
rect 580078 501880 580134 501936
rect 579894 497800 579950 497856
rect 580170 493720 580226 493776
rect 580170 489640 580226 489696
rect 580170 485560 580226 485616
rect 580170 481480 580226 481536
rect 580170 477400 580226 477456
rect 580170 473356 580172 473376
rect 580172 473356 580224 473376
rect 580224 473356 580226 473376
rect 580170 473320 580226 473356
rect 580170 465840 580226 465896
rect 580078 461760 580134 461816
rect 580078 457680 580134 457736
rect 578974 453600 579030 453656
rect 579710 449520 579766 449576
rect 580170 445440 580226 445496
rect 580170 441360 580226 441416
rect 579618 437280 579674 437336
rect 580170 433200 580226 433256
rect 579986 429800 580042 429856
rect 579618 425720 579674 425776
rect 580170 413480 580226 413536
rect 580170 405320 580226 405376
rect 580170 401240 580226 401296
rect 580170 393080 580226 393136
rect 579802 385600 579858 385656
rect 579986 381520 580042 381576
rect 580170 377440 580226 377496
rect 580170 373360 580226 373416
rect 580170 369280 580226 369336
rect 579618 365200 579674 365256
rect 579618 361120 579674 361176
rect 580170 357040 580226 357096
rect 579618 353640 579674 353696
rect 580170 349560 580226 349616
rect 580170 345480 580226 345536
rect 580170 341400 580226 341456
rect 579986 337320 580042 337376
rect 579986 333240 580042 333296
rect 579618 321000 579674 321056
rect 579618 316920 579674 316976
rect 580170 309440 580226 309496
rect 579618 305360 579674 305416
rect 580170 297200 580226 297256
rect 579986 293120 580042 293176
rect 579986 289040 580042 289096
rect 579066 284960 579122 285016
rect 578882 190984 578938 191040
rect 580170 280880 580226 280936
rect 580170 276800 580226 276856
rect 580170 273400 580226 273456
rect 580170 265240 580226 265296
rect 580262 257080 580318 257136
rect 579802 253000 579858 253056
rect 579802 248920 579858 248976
rect 580170 244840 580226 244896
rect 580170 237396 580172 237416
rect 580172 237396 580224 237416
rect 580224 237396 580226 237416
rect 580170 237360 580226 237396
rect 580170 221040 580226 221096
rect 580170 216960 580226 217016
rect 579986 204720 580042 204776
rect 580170 200640 580226 200696
rect 580170 197240 580226 197296
rect 580446 469920 580502 469976
rect 580354 195200 580410 195256
rect 579618 193160 579674 193216
rect 579986 189080 580042 189136
rect 580538 389680 580594 389736
rect 580630 313520 580686 313576
rect 580630 301280 580686 301336
rect 580630 269320 580686 269376
rect 580722 261160 580778 261216
rect 580722 240760 580778 240816
rect 580814 225120 580870 225176
rect 580538 192480 580594 192536
rect 580446 187584 580502 187640
rect 580170 185000 580226 185056
rect 578238 181328 578294 181384
rect 580170 180920 580226 180976
rect 566830 178608 566886 178664
rect 579802 176840 579858 176896
rect 559562 175072 559618 175128
rect 556802 174800 556858 174856
rect 580262 172760 580318 172816
rect 580170 164600 580226 164656
rect 580170 157120 580226 157176
rect 579802 153040 579858 153096
rect 580170 144880 580226 144936
rect 580354 168680 580410 168736
rect 580170 140800 580226 140856
rect 579802 132640 579858 132696
rect 580170 108840 580226 108896
rect 580170 80960 580226 81016
rect 534078 75112 534134 75168
rect 580170 72800 580226 72856
rect 579618 69536 579674 69592
rect 582470 637880 582526 637936
rect 582378 629720 582434 629776
rect 581642 610000 581698 610056
rect 580998 188264 581054 188320
rect 581734 573960 581790 574016
rect 581734 193840 581790 193896
rect 582562 614080 582618 614136
rect 582654 557640 582710 557696
rect 582746 533840 582802 533896
rect 582838 517520 582894 517576
rect 582838 180104 582894 180160
rect 582746 179968 582802 180024
rect 580630 128560 580686 128616
rect 580630 96600 580686 96656
rect 580538 84360 580594 84416
rect 580446 76880 580502 76936
rect 580354 68720 580410 68776
rect 580906 117000 580962 117056
rect 580814 112920 580870 112976
rect 580814 104760 580870 104816
rect 580722 92520 580778 92576
rect 580722 88440 580778 88496
rect 580906 100680 580962 100736
rect 580906 78648 580962 78704
rect 580630 63416 580686 63472
rect 580262 60560 580318 60616
rect 579894 56516 579896 56536
rect 579896 56516 579948 56536
rect 579948 56516 579950 56536
rect 579894 56480 579950 56516
rect 579894 52420 579950 52456
rect 579894 52400 579896 52420
rect 579896 52400 579948 52420
rect 579948 52400 579950 52420
rect 580170 48320 580226 48376
rect 579986 44240 580042 44296
rect 580170 40840 580226 40896
rect 580170 36760 580226 36816
rect 580170 32680 580226 32736
rect 580170 28600 580226 28656
rect 580170 24520 580226 24576
rect 580170 20440 580226 20496
rect 580170 16360 580226 16416
rect 580170 12280 580226 12336
rect 580170 8236 580172 8256
rect 580172 8236 580224 8256
rect 580224 8236 580226 8256
rect 580170 8200 580226 8236
rect 580170 4800 580226 4856
rect 578882 720 578938 776
<< metal3 >>
rect 580165 702538 580231 702541
rect 583520 702538 584960 702628
rect 580165 702536 584960 702538
rect 580165 702480 580170 702536
rect 580226 702480 584960 702536
rect 580165 702478 584960 702480
rect 580165 702475 580231 702478
rect 583520 702388 584960 702478
rect -960 701178 480 701268
rect 3417 701178 3483 701181
rect -960 701176 3483 701178
rect -960 701120 3422 701176
rect 3478 701120 3483 701176
rect -960 701118 3483 701120
rect -960 701028 480 701118
rect 3417 701115 3483 701118
rect 580165 698458 580231 698461
rect 583520 698458 584960 698548
rect 580165 698456 584960 698458
rect 580165 698400 580170 698456
rect 580226 698400 584960 698456
rect 580165 698398 584960 698400
rect 580165 698395 580231 698398
rect 583520 698308 584960 698398
rect -960 697778 480 697868
rect 3049 697778 3115 697781
rect -960 697776 3115 697778
rect -960 697720 3054 697776
rect 3110 697720 3115 697776
rect -960 697718 3115 697720
rect -960 697628 480 697718
rect 3049 697715 3115 697718
rect 580165 694378 580231 694381
rect 583520 694378 584960 694468
rect 580165 694376 584960 694378
rect 580165 694320 580170 694376
rect 580226 694320 584960 694376
rect 580165 694318 584960 694320
rect 580165 694315 580231 694318
rect 583520 694228 584960 694318
rect -960 693548 480 693788
rect 580165 690298 580231 690301
rect 583520 690298 584960 690388
rect 580165 690296 584960 690298
rect 580165 690240 580170 690296
rect 580226 690240 584960 690296
rect 580165 690238 584960 690240
rect 580165 690235 580231 690238
rect 583520 690148 584960 690238
rect -960 689618 480 689708
rect 3417 689618 3483 689621
rect -960 689616 3483 689618
rect -960 689560 3422 689616
rect 3478 689560 3483 689616
rect -960 689558 3483 689560
rect -960 689468 480 689558
rect 3417 689555 3483 689558
rect 579797 686218 579863 686221
rect 583520 686218 584960 686308
rect 579797 686216 584960 686218
rect 579797 686160 579802 686216
rect 579858 686160 584960 686216
rect 579797 686158 584960 686160
rect 579797 686155 579863 686158
rect 583520 686068 584960 686158
rect -960 685538 480 685628
rect 3141 685538 3207 685541
rect -960 685536 3207 685538
rect -960 685480 3146 685536
rect 3202 685480 3207 685536
rect -960 685478 3207 685480
rect -960 685388 480 685478
rect 3141 685475 3207 685478
rect 580165 682138 580231 682141
rect 583520 682138 584960 682228
rect 580165 682136 584960 682138
rect 580165 682080 580170 682136
rect 580226 682080 584960 682136
rect 580165 682078 584960 682080
rect 580165 682075 580231 682078
rect 583520 681988 584960 682078
rect -960 681458 480 681548
rect 3417 681458 3483 681461
rect -960 681456 3483 681458
rect -960 681400 3422 681456
rect 3478 681400 3483 681456
rect -960 681398 3483 681400
rect -960 681308 480 681398
rect 3417 681395 3483 681398
rect 580165 678058 580231 678061
rect 583520 678058 584960 678148
rect 580165 678056 584960 678058
rect 580165 678000 580170 678056
rect 580226 678000 584960 678056
rect 580165 677998 584960 678000
rect 580165 677995 580231 677998
rect 583520 677908 584960 677998
rect -960 677378 480 677468
rect 3417 677378 3483 677381
rect -960 677376 3483 677378
rect -960 677320 3422 677376
rect 3478 677320 3483 677376
rect -960 677318 3483 677320
rect -960 677228 480 677318
rect 3417 677315 3483 677318
rect 580165 673978 580231 673981
rect 583520 673978 584960 674068
rect 580165 673976 584960 673978
rect 580165 673920 580170 673976
rect 580226 673920 584960 673976
rect 580165 673918 584960 673920
rect 580165 673915 580231 673918
rect 583520 673828 584960 673918
rect -960 673148 480 673388
rect 580165 669898 580231 669901
rect 583520 669898 584960 669988
rect 580165 669896 584960 669898
rect 580165 669840 580170 669896
rect 580226 669840 584960 669896
rect 580165 669838 584960 669840
rect 580165 669835 580231 669838
rect 583520 669748 584960 669838
rect -960 669068 480 669308
rect 583520 665668 584960 665908
rect -960 665138 480 665228
rect 3233 665138 3299 665141
rect -960 665136 3299 665138
rect -960 665080 3238 665136
rect 3294 665080 3299 665136
rect -960 665078 3299 665080
rect -960 664988 480 665078
rect 3233 665075 3299 665078
rect 580165 662418 580231 662421
rect 583520 662418 584960 662508
rect 580165 662416 584960 662418
rect 580165 662360 580170 662416
rect 580226 662360 584960 662416
rect 580165 662358 584960 662360
rect 580165 662355 580231 662358
rect 583520 662268 584960 662358
rect -960 661058 480 661148
rect 3417 661058 3483 661061
rect -960 661056 3483 661058
rect -960 661000 3422 661056
rect 3478 661000 3483 661056
rect -960 660998 3483 661000
rect -960 660908 480 660998
rect 3417 660995 3483 660998
rect 580165 658338 580231 658341
rect 583520 658338 584960 658428
rect 580165 658336 584960 658338
rect 580165 658280 580170 658336
rect 580226 658280 584960 658336
rect 580165 658278 584960 658280
rect 580165 658275 580231 658278
rect 583520 658188 584960 658278
rect -960 657658 480 657748
rect -960 657598 674 657658
rect -960 657522 480 657598
rect 614 657522 674 657598
rect -960 657508 674 657522
rect 246 657462 674 657508
rect 246 656978 306 657462
rect 95734 656978 95740 656980
rect 246 656918 95740 656978
rect 95734 656916 95740 656918
rect 95804 656916 95810 656980
rect 580165 654258 580231 654261
rect 583520 654258 584960 654348
rect 580165 654256 584960 654258
rect 580165 654200 580170 654256
rect 580226 654200 584960 654256
rect 580165 654198 584960 654200
rect 580165 654195 580231 654198
rect 583520 654108 584960 654198
rect -960 653578 480 653668
rect 3049 653578 3115 653581
rect -960 653576 3115 653578
rect -960 653520 3054 653576
rect 3110 653520 3115 653576
rect -960 653518 3115 653520
rect -960 653428 480 653518
rect 3049 653515 3115 653518
rect 583520 650028 584960 650268
rect -960 649348 480 649588
rect 580165 646098 580231 646101
rect 583520 646098 584960 646188
rect 580165 646096 584960 646098
rect 580165 646040 580170 646096
rect 580226 646040 584960 646096
rect 580165 646038 584960 646040
rect 580165 646035 580231 646038
rect 583520 645948 584960 646038
rect -960 645418 480 645508
rect 3417 645418 3483 645421
rect -960 645416 3483 645418
rect -960 645360 3422 645416
rect 3478 645360 3483 645416
rect -960 645358 3483 645360
rect -960 645268 480 645358
rect 3417 645355 3483 645358
rect 580165 642018 580231 642021
rect 583520 642018 584960 642108
rect 580165 642016 584960 642018
rect 580165 641960 580170 642016
rect 580226 641960 584960 642016
rect 580165 641958 584960 641960
rect 580165 641955 580231 641958
rect 583520 641868 584960 641958
rect -960 641338 480 641428
rect 3141 641338 3207 641341
rect -960 641336 3207 641338
rect -960 641280 3146 641336
rect 3202 641280 3207 641336
rect -960 641278 3207 641280
rect -960 641188 480 641278
rect 3141 641275 3207 641278
rect 582465 637938 582531 637941
rect 583520 637938 584960 638028
rect 582465 637936 584960 637938
rect 582465 637880 582470 637936
rect 582526 637880 584960 637936
rect 582465 637878 584960 637880
rect 582465 637875 582531 637878
rect 583520 637788 584960 637878
rect -960 637258 480 637348
rect 3141 637258 3207 637261
rect -960 637256 3207 637258
rect -960 637200 3146 637256
rect 3202 637200 3207 637256
rect -960 637198 3207 637200
rect -960 637108 480 637198
rect 3141 637195 3207 637198
rect 583520 633708 584960 633948
rect -960 633178 480 633268
rect 3417 633178 3483 633181
rect -960 633176 3483 633178
rect -960 633120 3422 633176
rect 3478 633120 3483 633176
rect -960 633118 3483 633120
rect -960 633028 480 633118
rect 3417 633115 3483 633118
rect 582373 629778 582439 629781
rect 583520 629778 584960 629868
rect 582373 629776 584960 629778
rect 582373 629720 582378 629776
rect 582434 629720 584960 629776
rect 582373 629718 584960 629720
rect 582373 629715 582439 629718
rect 583520 629628 584960 629718
rect -960 628948 480 629188
rect 580165 626378 580231 626381
rect 583520 626378 584960 626468
rect 580165 626376 584960 626378
rect 580165 626320 580170 626376
rect 580226 626320 584960 626376
rect 580165 626318 584960 626320
rect 580165 626315 580231 626318
rect 583520 626228 584960 626318
rect -960 625018 480 625108
rect 3233 625018 3299 625021
rect -960 625016 3299 625018
rect -960 624960 3238 625016
rect 3294 624960 3299 625016
rect -960 624958 3299 624960
rect -960 624868 480 624958
rect 3233 624955 3299 624958
rect 579797 622298 579863 622301
rect 583520 622298 584960 622388
rect 579797 622296 584960 622298
rect 579797 622240 579802 622296
rect 579858 622240 584960 622296
rect 579797 622238 584960 622240
rect 579797 622235 579863 622238
rect 583520 622148 584960 622238
rect -960 621618 480 621708
rect 3417 621618 3483 621621
rect -960 621616 3483 621618
rect -960 621560 3422 621616
rect 3478 621560 3483 621616
rect -960 621558 3483 621560
rect -960 621468 480 621558
rect 3417 621555 3483 621558
rect 583520 618068 584960 618308
rect -960 617538 480 617628
rect 3141 617538 3207 617541
rect -960 617536 3207 617538
rect -960 617480 3146 617536
rect 3202 617480 3207 617536
rect -960 617478 3207 617480
rect -960 617388 480 617478
rect 3141 617475 3207 617478
rect 582557 614138 582623 614141
rect 583520 614138 584960 614228
rect 582557 614136 584960 614138
rect 582557 614080 582562 614136
rect 582618 614080 584960 614136
rect 582557 614078 584960 614080
rect 582557 614075 582623 614078
rect 583520 613988 584960 614078
rect -960 613458 480 613548
rect 3141 613458 3207 613461
rect -960 613456 3207 613458
rect -960 613400 3146 613456
rect 3202 613400 3207 613456
rect -960 613398 3207 613400
rect -960 613308 480 613398
rect 3141 613395 3207 613398
rect 581637 610058 581703 610061
rect 583520 610058 584960 610148
rect 581637 610056 584960 610058
rect 581637 610000 581642 610056
rect 581698 610000 584960 610056
rect 581637 609998 584960 610000
rect 581637 609995 581703 609998
rect 583520 609908 584960 609998
rect -960 609378 480 609468
rect 3417 609378 3483 609381
rect -960 609376 3483 609378
rect -960 609320 3422 609376
rect 3478 609320 3483 609376
rect -960 609318 3483 609320
rect -960 609228 480 609318
rect 3417 609315 3483 609318
rect 580165 605978 580231 605981
rect 583520 605978 584960 606068
rect 580165 605976 584960 605978
rect 580165 605920 580170 605976
rect 580226 605920 584960 605976
rect 580165 605918 584960 605920
rect 580165 605915 580231 605918
rect 583520 605828 584960 605918
rect -960 605298 480 605388
rect 3049 605298 3115 605301
rect -960 605296 3115 605298
rect -960 605240 3054 605296
rect 3110 605240 3115 605296
rect -960 605238 3115 605240
rect -960 605148 480 605238
rect 3049 605235 3115 605238
rect 580165 601898 580231 601901
rect 583520 601898 584960 601988
rect 580165 601896 584960 601898
rect 580165 601840 580170 601896
rect 580226 601840 584960 601896
rect 580165 601838 584960 601840
rect 580165 601835 580231 601838
rect 583520 601748 584960 601838
rect -960 601218 480 601308
rect 3509 601218 3575 601221
rect -960 601216 3575 601218
rect -960 601160 3514 601216
rect 3570 601160 3575 601216
rect -960 601158 3575 601160
rect -960 601068 480 601158
rect 3509 601155 3575 601158
rect 580349 597818 580415 597821
rect 583520 597818 584960 597908
rect 580349 597816 584960 597818
rect 580349 597760 580354 597816
rect 580410 597760 584960 597816
rect 580349 597758 584960 597760
rect 580349 597755 580415 597758
rect 583520 597668 584960 597758
rect -960 597138 480 597228
rect 3049 597138 3115 597141
rect -960 597136 3115 597138
rect -960 597080 3054 597136
rect 3110 597080 3115 597136
rect -960 597078 3115 597080
rect -960 596988 480 597078
rect 3049 597075 3115 597078
rect 583520 593588 584960 593828
rect -960 593058 480 593148
rect 3141 593058 3207 593061
rect -960 593056 3207 593058
rect -960 593000 3146 593056
rect 3202 593000 3207 593056
rect -960 592998 3207 593000
rect -960 592908 480 592998
rect 3141 592995 3207 592998
rect 580165 589658 580231 589661
rect 583520 589658 584960 589748
rect 580165 589656 584960 589658
rect 580165 589600 580170 589656
rect 580226 589600 584960 589656
rect 580165 589598 584960 589600
rect 580165 589595 580231 589598
rect 583520 589508 584960 589598
rect -960 588978 480 589068
rect 3233 588978 3299 588981
rect -960 588976 3299 588978
rect -960 588920 3238 588976
rect 3294 588920 3299 588976
rect -960 588918 3299 588920
rect -960 588828 480 588918
rect 3233 588915 3299 588918
rect 578877 586258 578943 586261
rect 583520 586258 584960 586348
rect 578877 586256 584960 586258
rect 578877 586200 578882 586256
rect 578938 586200 584960 586256
rect 578877 586198 584960 586200
rect 578877 586195 578943 586198
rect 583520 586108 584960 586198
rect -960 584898 480 584988
rect 3141 584898 3207 584901
rect -960 584896 3207 584898
rect -960 584840 3146 584896
rect 3202 584840 3207 584896
rect -960 584838 3207 584840
rect -960 584748 480 584838
rect 3141 584835 3207 584838
rect 583520 582028 584960 582268
rect -960 581498 480 581588
rect 3325 581498 3391 581501
rect -960 581496 3391 581498
rect -960 581440 3330 581496
rect 3386 581440 3391 581496
rect -960 581438 3391 581440
rect -960 581348 480 581438
rect 3325 581435 3391 581438
rect 583520 577948 584960 578188
rect -960 577418 480 577508
rect 3509 577418 3575 577421
rect -960 577416 3575 577418
rect -960 577360 3514 577416
rect 3570 577360 3575 577416
rect -960 577358 3575 577360
rect -960 577268 480 577358
rect 3509 577355 3575 577358
rect 581729 574018 581795 574021
rect 583520 574018 584960 574108
rect 581729 574016 584960 574018
rect 581729 573960 581734 574016
rect 581790 573960 584960 574016
rect 581729 573958 584960 573960
rect 581729 573955 581795 573958
rect 583520 573868 584960 573958
rect -960 573188 480 573428
rect 580165 569938 580231 569941
rect 583520 569938 584960 570028
rect 580165 569936 584960 569938
rect 580165 569880 580170 569936
rect 580226 569880 584960 569936
rect 580165 569878 584960 569880
rect 580165 569875 580231 569878
rect 583520 569788 584960 569878
rect -960 569258 480 569348
rect 2865 569258 2931 569261
rect -960 569256 2931 569258
rect -960 569200 2870 569256
rect 2926 569200 2931 569256
rect -960 569198 2931 569200
rect -960 569108 480 569198
rect 2865 569195 2931 569198
rect 580165 565858 580231 565861
rect 583520 565858 584960 565948
rect 580165 565856 584960 565858
rect 580165 565800 580170 565856
rect 580226 565800 584960 565856
rect 580165 565798 584960 565800
rect 580165 565795 580231 565798
rect 583520 565708 584960 565798
rect -960 565028 480 565268
rect 583520 561628 584960 561868
rect -960 561098 480 561188
rect 3049 561098 3115 561101
rect -960 561096 3115 561098
rect -960 561040 3054 561096
rect 3110 561040 3115 561096
rect -960 561038 3115 561040
rect -960 560948 480 561038
rect 3049 561035 3115 561038
rect 582649 557698 582715 557701
rect 583520 557698 584960 557788
rect 582649 557696 584960 557698
rect 582649 557640 582654 557696
rect 582710 557640 584960 557696
rect 582649 557638 584960 557640
rect 582649 557635 582715 557638
rect 583520 557548 584960 557638
rect -960 557018 480 557108
rect 3049 557018 3115 557021
rect -960 557016 3115 557018
rect -960 556960 3054 557016
rect 3110 556960 3115 557016
rect -960 556958 3115 556960
rect -960 556868 480 556958
rect 3049 556955 3115 556958
rect 580165 553618 580231 553621
rect 583520 553618 584960 553708
rect 580165 553616 584960 553618
rect 580165 553560 580170 553616
rect 580226 553560 584960 553616
rect 580165 553558 584960 553560
rect 580165 553555 580231 553558
rect 583520 553468 584960 553558
rect -960 552938 480 553028
rect 3509 552938 3575 552941
rect -960 552936 3575 552938
rect -960 552880 3514 552936
rect 3570 552880 3575 552936
rect -960 552878 3575 552880
rect -960 552788 480 552878
rect 3509 552875 3575 552878
rect 580165 549538 580231 549541
rect 583520 549538 584960 549628
rect 580165 549536 584960 549538
rect 580165 549480 580170 549536
rect 580226 549480 584960 549536
rect 580165 549478 584960 549480
rect 580165 549475 580231 549478
rect 583520 549388 584960 549478
rect -960 548858 480 548948
rect 3049 548858 3115 548861
rect -960 548856 3115 548858
rect -960 548800 3054 548856
rect 3110 548800 3115 548856
rect -960 548798 3115 548800
rect -960 548708 480 548798
rect 3049 548795 3115 548798
rect 579889 546138 579955 546141
rect 583520 546138 584960 546228
rect 579889 546136 584960 546138
rect 579889 546080 579894 546136
rect 579950 546080 584960 546136
rect 579889 546078 584960 546080
rect 579889 546075 579955 546078
rect 583520 545988 584960 546078
rect -960 544778 480 544868
rect 3141 544778 3207 544781
rect -960 544776 3207 544778
rect -960 544720 3146 544776
rect 3202 544720 3207 544776
rect -960 544718 3207 544720
rect -960 544628 480 544718
rect 3141 544715 3207 544718
rect 580165 542058 580231 542061
rect 583520 542058 584960 542148
rect 580165 542056 584960 542058
rect 580165 542000 580170 542056
rect 580226 542000 584960 542056
rect 580165 541998 584960 542000
rect 580165 541995 580231 541998
rect 583520 541908 584960 541998
rect -960 541378 480 541468
rect 3509 541378 3575 541381
rect -960 541376 3575 541378
rect -960 541320 3514 541376
rect 3570 541320 3575 541376
rect -960 541318 3575 541320
rect -960 541228 480 541318
rect 3509 541315 3575 541318
rect 580165 537978 580231 537981
rect 583520 537978 584960 538068
rect 580165 537976 584960 537978
rect 580165 537920 580170 537976
rect 580226 537920 584960 537976
rect 580165 537918 584960 537920
rect 580165 537915 580231 537918
rect 583520 537828 584960 537918
rect -960 537298 480 537388
rect 3325 537298 3391 537301
rect -960 537296 3391 537298
rect -960 537240 3330 537296
rect 3386 537240 3391 537296
rect -960 537238 3391 537240
rect -960 537148 480 537238
rect 3325 537235 3391 537238
rect 582741 533898 582807 533901
rect 583520 533898 584960 533988
rect 582741 533896 584960 533898
rect 582741 533840 582746 533896
rect 582802 533840 584960 533896
rect 582741 533838 584960 533840
rect 582741 533835 582807 533838
rect 583520 533748 584960 533838
rect -960 533218 480 533308
rect 3325 533218 3391 533221
rect -960 533216 3391 533218
rect -960 533160 3330 533216
rect 3386 533160 3391 533216
rect -960 533158 3391 533160
rect -960 533068 480 533158
rect 3325 533155 3391 533158
rect 579797 529818 579863 529821
rect 583520 529818 584960 529908
rect 579797 529816 584960 529818
rect 579797 529760 579802 529816
rect 579858 529760 584960 529816
rect 579797 529758 584960 529760
rect 579797 529755 579863 529758
rect 583520 529668 584960 529758
rect -960 529138 480 529228
rect 3509 529138 3575 529141
rect -960 529136 3575 529138
rect -960 529080 3514 529136
rect 3570 529080 3575 529136
rect -960 529078 3575 529080
rect -960 528988 480 529078
rect 3509 529075 3575 529078
rect 580165 525738 580231 525741
rect 583520 525738 584960 525828
rect 580165 525736 584960 525738
rect 580165 525680 580170 525736
rect 580226 525680 584960 525736
rect 580165 525678 584960 525680
rect 580165 525675 580231 525678
rect 583520 525588 584960 525678
rect -960 525058 480 525148
rect 3509 525058 3575 525061
rect -960 525056 3575 525058
rect -960 525000 3514 525056
rect 3570 525000 3575 525056
rect -960 524998 3575 525000
rect -960 524908 480 524998
rect 3509 524995 3575 524998
rect 580165 521658 580231 521661
rect 583520 521658 584960 521748
rect 580165 521656 584960 521658
rect 580165 521600 580170 521656
rect 580226 521600 584960 521656
rect 580165 521598 584960 521600
rect 580165 521595 580231 521598
rect 583520 521508 584960 521598
rect -960 520978 480 521068
rect 2865 520978 2931 520981
rect -960 520976 2931 520978
rect -960 520920 2870 520976
rect 2926 520920 2931 520976
rect -960 520918 2931 520920
rect -960 520828 480 520918
rect 2865 520915 2931 520918
rect 582833 517578 582899 517581
rect 583520 517578 584960 517668
rect 582833 517576 584960 517578
rect 582833 517520 582838 517576
rect 582894 517520 584960 517576
rect 582833 517518 584960 517520
rect 582833 517515 582899 517518
rect 583520 517428 584960 517518
rect -960 516898 480 516988
rect 2957 516898 3023 516901
rect -960 516896 3023 516898
rect -960 516840 2962 516896
rect 3018 516840 3023 516896
rect -960 516838 3023 516840
rect -960 516748 480 516838
rect 2957 516835 3023 516838
rect 583520 513348 584960 513588
rect -960 512818 480 512908
rect 3049 512818 3115 512821
rect -960 512816 3115 512818
rect -960 512760 3054 512816
rect 3110 512760 3115 512816
rect -960 512758 3115 512760
rect -960 512668 480 512758
rect 3049 512755 3115 512758
rect 580165 510098 580231 510101
rect 583520 510098 584960 510188
rect 580165 510096 584960 510098
rect 580165 510040 580170 510096
rect 580226 510040 584960 510096
rect 580165 510038 584960 510040
rect 580165 510035 580231 510038
rect 583520 509948 584960 510038
rect -960 508738 480 508828
rect 3509 508738 3575 508741
rect -960 508736 3575 508738
rect -960 508680 3514 508736
rect 3570 508680 3575 508736
rect -960 508678 3575 508680
rect -960 508588 480 508678
rect 3509 508675 3575 508678
rect 580073 506018 580139 506021
rect 583520 506018 584960 506108
rect 580073 506016 584960 506018
rect 580073 505960 580078 506016
rect 580134 505960 584960 506016
rect 580073 505958 584960 505960
rect 580073 505955 580139 505958
rect 583520 505868 584960 505958
rect -960 504658 480 504748
rect 3049 504658 3115 504661
rect -960 504656 3115 504658
rect -960 504600 3054 504656
rect 3110 504600 3115 504656
rect -960 504598 3115 504600
rect -960 504508 480 504598
rect 3049 504595 3115 504598
rect 580073 501938 580139 501941
rect 583520 501938 584960 502028
rect 580073 501936 584960 501938
rect 580073 501880 580078 501936
rect 580134 501880 584960 501936
rect 580073 501878 584960 501880
rect 580073 501875 580139 501878
rect 583520 501788 584960 501878
rect -960 501108 480 501348
rect 579889 497858 579955 497861
rect 583520 497858 584960 497948
rect 579889 497856 584960 497858
rect 579889 497800 579894 497856
rect 579950 497800 584960 497856
rect 579889 497798 584960 497800
rect 579889 497795 579955 497798
rect 583520 497708 584960 497798
rect -960 497178 480 497268
rect 3325 497178 3391 497181
rect -960 497176 3391 497178
rect -960 497120 3330 497176
rect 3386 497120 3391 497176
rect -960 497118 3391 497120
rect -960 497028 480 497118
rect 3325 497115 3391 497118
rect 580165 493778 580231 493781
rect 583520 493778 584960 493868
rect 580165 493776 584960 493778
rect 580165 493720 580170 493776
rect 580226 493720 584960 493776
rect 580165 493718 584960 493720
rect 580165 493715 580231 493718
rect 583520 493628 584960 493718
rect -960 493098 480 493188
rect 3509 493098 3575 493101
rect -960 493096 3575 493098
rect -960 493040 3514 493096
rect 3570 493040 3575 493096
rect -960 493038 3575 493040
rect -960 492948 480 493038
rect 3509 493035 3575 493038
rect 580165 489698 580231 489701
rect 583520 489698 584960 489788
rect 580165 489696 584960 489698
rect 580165 489640 580170 489696
rect 580226 489640 584960 489696
rect 580165 489638 584960 489640
rect 580165 489635 580231 489638
rect 583520 489548 584960 489638
rect -960 489018 480 489108
rect 3325 489018 3391 489021
rect -960 489016 3391 489018
rect -960 488960 3330 489016
rect 3386 488960 3391 489016
rect -960 488958 3391 488960
rect -960 488868 480 488958
rect 3325 488955 3391 488958
rect 580165 485618 580231 485621
rect 583520 485618 584960 485708
rect 580165 485616 584960 485618
rect 580165 485560 580170 485616
rect 580226 485560 584960 485616
rect 580165 485558 584960 485560
rect 580165 485555 580231 485558
rect 583520 485468 584960 485558
rect -960 484938 480 485028
rect 3509 484938 3575 484941
rect -960 484936 3575 484938
rect -960 484880 3514 484936
rect 3570 484880 3575 484936
rect -960 484878 3575 484880
rect -960 484788 480 484878
rect 3509 484875 3575 484878
rect 580165 481538 580231 481541
rect 583520 481538 584960 481628
rect 580165 481536 584960 481538
rect 580165 481480 580170 481536
rect 580226 481480 584960 481536
rect 580165 481478 584960 481480
rect 580165 481475 580231 481478
rect 583520 481388 584960 481478
rect -960 480858 480 480948
rect 3509 480858 3575 480861
rect -960 480856 3575 480858
rect -960 480800 3514 480856
rect 3570 480800 3575 480856
rect -960 480798 3575 480800
rect -960 480708 480 480798
rect 3509 480795 3575 480798
rect 580165 477458 580231 477461
rect 583520 477458 584960 477548
rect 580165 477456 584960 477458
rect 580165 477400 580170 477456
rect 580226 477400 584960 477456
rect 580165 477398 584960 477400
rect 580165 477395 580231 477398
rect 583520 477308 584960 477398
rect -960 476778 480 476868
rect 2865 476778 2931 476781
rect -960 476776 2931 476778
rect -960 476720 2870 476776
rect 2926 476720 2931 476776
rect -960 476718 2931 476720
rect -960 476628 480 476718
rect 2865 476715 2931 476718
rect 580165 473378 580231 473381
rect 583520 473378 584960 473468
rect 580165 473376 584960 473378
rect 580165 473320 580170 473376
rect 580226 473320 584960 473376
rect 580165 473318 584960 473320
rect 580165 473315 580231 473318
rect 583520 473228 584960 473318
rect -960 472698 480 472788
rect 2865 472698 2931 472701
rect -960 472696 2931 472698
rect -960 472640 2870 472696
rect 2926 472640 2931 472696
rect -960 472638 2931 472640
rect -960 472548 480 472638
rect 2865 472635 2931 472638
rect 580441 469978 580507 469981
rect 583520 469978 584960 470068
rect 580441 469976 584960 469978
rect 580441 469920 580446 469976
rect 580502 469920 584960 469976
rect 580441 469918 584960 469920
rect 580441 469915 580507 469918
rect 583520 469828 584960 469918
rect -960 468618 480 468708
rect 2957 468618 3023 468621
rect -960 468616 3023 468618
rect -960 468560 2962 468616
rect 3018 468560 3023 468616
rect -960 468558 3023 468560
rect -960 468468 480 468558
rect 2957 468555 3023 468558
rect 580165 465898 580231 465901
rect 583520 465898 584960 465988
rect 580165 465896 584960 465898
rect 580165 465840 580170 465896
rect 580226 465840 584960 465896
rect 580165 465838 584960 465840
rect 580165 465835 580231 465838
rect 583520 465748 584960 465838
rect -960 465218 480 465308
rect 3509 465218 3575 465221
rect -960 465216 3575 465218
rect -960 465160 3514 465216
rect 3570 465160 3575 465216
rect -960 465158 3575 465160
rect -960 465068 480 465158
rect 3509 465155 3575 465158
rect 580073 461818 580139 461821
rect 583520 461818 584960 461908
rect 580073 461816 584960 461818
rect 580073 461760 580078 461816
rect 580134 461760 584960 461816
rect 580073 461758 584960 461760
rect 580073 461755 580139 461758
rect 583520 461668 584960 461758
rect -960 461138 480 461228
rect 3509 461138 3575 461141
rect -960 461136 3575 461138
rect -960 461080 3514 461136
rect 3570 461080 3575 461136
rect -960 461078 3575 461080
rect -960 460988 480 461078
rect 3509 461075 3575 461078
rect 580073 457738 580139 457741
rect 583520 457738 584960 457828
rect 580073 457736 584960 457738
rect 580073 457680 580078 457736
rect 580134 457680 584960 457736
rect 580073 457678 584960 457680
rect 580073 457675 580139 457678
rect 583520 457588 584960 457678
rect -960 457058 480 457148
rect 3233 457058 3299 457061
rect -960 457056 3299 457058
rect -960 457000 3238 457056
rect 3294 457000 3299 457056
rect -960 456998 3299 457000
rect -960 456908 480 456998
rect 3233 456995 3299 456998
rect 578969 453658 579035 453661
rect 583520 453658 584960 453748
rect 578969 453656 584960 453658
rect 578969 453600 578974 453656
rect 579030 453600 584960 453656
rect 578969 453598 584960 453600
rect 578969 453595 579035 453598
rect 583520 453508 584960 453598
rect -960 452978 480 453068
rect 3325 452978 3391 452981
rect -960 452976 3391 452978
rect -960 452920 3330 452976
rect 3386 452920 3391 452976
rect -960 452918 3391 452920
rect -960 452828 480 452918
rect 3325 452915 3391 452918
rect 579705 449578 579771 449581
rect 583520 449578 584960 449668
rect 579705 449576 584960 449578
rect 579705 449520 579710 449576
rect 579766 449520 584960 449576
rect 579705 449518 584960 449520
rect 579705 449515 579771 449518
rect 583520 449428 584960 449518
rect -960 448898 480 448988
rect 3325 448898 3391 448901
rect -960 448896 3391 448898
rect -960 448840 3330 448896
rect 3386 448840 3391 448896
rect -960 448838 3391 448840
rect -960 448748 480 448838
rect 3325 448835 3391 448838
rect 580165 445498 580231 445501
rect 583520 445498 584960 445588
rect 580165 445496 584960 445498
rect 580165 445440 580170 445496
rect 580226 445440 584960 445496
rect 580165 445438 584960 445440
rect 580165 445435 580231 445438
rect 583520 445348 584960 445438
rect -960 444818 480 444908
rect 3509 444818 3575 444821
rect -960 444816 3575 444818
rect -960 444760 3514 444816
rect 3570 444760 3575 444816
rect -960 444758 3575 444760
rect -960 444668 480 444758
rect 3509 444755 3575 444758
rect 580165 441418 580231 441421
rect 583520 441418 584960 441508
rect 580165 441416 584960 441418
rect 580165 441360 580170 441416
rect 580226 441360 584960 441416
rect 580165 441358 584960 441360
rect 580165 441355 580231 441358
rect 583520 441268 584960 441358
rect -960 440738 480 440828
rect 3325 440738 3391 440741
rect -960 440736 3391 440738
rect -960 440680 3330 440736
rect 3386 440680 3391 440736
rect -960 440678 3391 440680
rect -960 440588 480 440678
rect 3325 440675 3391 440678
rect 579613 437338 579679 437341
rect 583520 437338 584960 437428
rect 579613 437336 584960 437338
rect 579613 437280 579618 437336
rect 579674 437280 584960 437336
rect 579613 437278 584960 437280
rect 579613 437275 579679 437278
rect 583520 437188 584960 437278
rect -960 436658 480 436748
rect 3509 436658 3575 436661
rect -960 436656 3575 436658
rect -960 436600 3514 436656
rect 3570 436600 3575 436656
rect -960 436598 3575 436600
rect -960 436508 480 436598
rect 3509 436595 3575 436598
rect 580165 433258 580231 433261
rect 583520 433258 584960 433348
rect 580165 433256 584960 433258
rect 580165 433200 580170 433256
rect 580226 433200 584960 433256
rect 580165 433198 584960 433200
rect 580165 433195 580231 433198
rect 583520 433108 584960 433198
rect -960 432578 480 432668
rect 3509 432578 3575 432581
rect -960 432576 3575 432578
rect -960 432520 3514 432576
rect 3570 432520 3575 432576
rect -960 432518 3575 432520
rect -960 432428 480 432518
rect 3509 432515 3575 432518
rect 579981 429858 580047 429861
rect 583520 429858 584960 429948
rect 579981 429856 584960 429858
rect 579981 429800 579986 429856
rect 580042 429800 584960 429856
rect 579981 429798 584960 429800
rect 579981 429795 580047 429798
rect 583520 429708 584960 429798
rect -960 428498 480 428588
rect 2865 428498 2931 428501
rect -960 428496 2931 428498
rect -960 428440 2870 428496
rect 2926 428440 2931 428496
rect -960 428438 2931 428440
rect -960 428348 480 428438
rect 2865 428435 2931 428438
rect 579613 425778 579679 425781
rect 583520 425778 584960 425868
rect 579613 425776 584960 425778
rect 579613 425720 579618 425776
rect 579674 425720 584960 425776
rect 579613 425718 584960 425720
rect 579613 425715 579679 425718
rect 583520 425628 584960 425718
rect -960 424948 480 425188
rect 583520 421548 584960 421788
rect -960 420868 480 421108
rect 583520 417468 584960 417708
rect -960 416938 480 417028
rect 3509 416938 3575 416941
rect -960 416936 3575 416938
rect -960 416880 3514 416936
rect 3570 416880 3575 416936
rect -960 416878 3575 416880
rect -960 416788 480 416878
rect 3509 416875 3575 416878
rect 580165 413538 580231 413541
rect 583520 413538 584960 413628
rect 580165 413536 584960 413538
rect 580165 413480 580170 413536
rect 580226 413480 584960 413536
rect 580165 413478 584960 413480
rect 580165 413475 580231 413478
rect 583520 413388 584960 413478
rect -960 412858 480 412948
rect 3509 412858 3575 412861
rect -960 412856 3575 412858
rect -960 412800 3514 412856
rect 3570 412800 3575 412856
rect -960 412798 3575 412800
rect -960 412708 480 412798
rect 3509 412795 3575 412798
rect 583520 409308 584960 409548
rect -960 408778 480 408868
rect 3509 408778 3575 408781
rect -960 408776 3575 408778
rect -960 408720 3514 408776
rect 3570 408720 3575 408776
rect -960 408718 3575 408720
rect -960 408628 480 408718
rect 3509 408715 3575 408718
rect 580165 405378 580231 405381
rect 583520 405378 584960 405468
rect 580165 405376 584960 405378
rect 580165 405320 580170 405376
rect 580226 405320 584960 405376
rect 580165 405318 584960 405320
rect 580165 405315 580231 405318
rect 583520 405228 584960 405318
rect -960 404698 480 404788
rect 3509 404698 3575 404701
rect -960 404696 3575 404698
rect -960 404640 3514 404696
rect 3570 404640 3575 404696
rect -960 404638 3575 404640
rect -960 404548 480 404638
rect 3509 404635 3575 404638
rect 580165 401298 580231 401301
rect 583520 401298 584960 401388
rect 580165 401296 584960 401298
rect 580165 401240 580170 401296
rect 580226 401240 584960 401296
rect 580165 401238 584960 401240
rect 580165 401235 580231 401238
rect 583520 401148 584960 401238
rect -960 400618 480 400708
rect 3233 400618 3299 400621
rect -960 400616 3299 400618
rect -960 400560 3238 400616
rect 3294 400560 3299 400616
rect -960 400558 3299 400560
rect -960 400468 480 400558
rect 3233 400555 3299 400558
rect 583520 397068 584960 397308
rect -960 396538 480 396628
rect 3601 396538 3667 396541
rect -960 396536 3667 396538
rect -960 396480 3606 396536
rect 3662 396480 3667 396536
rect -960 396478 3667 396480
rect -960 396388 480 396478
rect 3601 396475 3667 396478
rect 580165 393138 580231 393141
rect 583520 393138 584960 393228
rect 580165 393136 584960 393138
rect 580165 393080 580170 393136
rect 580226 393080 584960 393136
rect 580165 393078 584960 393080
rect 580165 393075 580231 393078
rect 583520 392988 584960 393078
rect -960 392308 480 392548
rect 580533 389738 580599 389741
rect 583520 389738 584960 389828
rect 580533 389736 584960 389738
rect 580533 389680 580538 389736
rect 580594 389680 584960 389736
rect 580533 389678 584960 389680
rect 580533 389675 580599 389678
rect 583520 389588 584960 389678
rect -960 388378 480 388468
rect 2957 388378 3023 388381
rect -960 388376 3023 388378
rect -960 388320 2962 388376
rect 3018 388320 3023 388376
rect -960 388318 3023 388320
rect -960 388228 480 388318
rect 2957 388315 3023 388318
rect 579797 385658 579863 385661
rect 583520 385658 584960 385748
rect 579797 385656 584960 385658
rect 579797 385600 579802 385656
rect 579858 385600 584960 385656
rect 579797 385598 584960 385600
rect 579797 385595 579863 385598
rect 583520 385508 584960 385598
rect -960 384978 480 385068
rect 3141 384978 3207 384981
rect -960 384976 3207 384978
rect -960 384920 3146 384976
rect 3202 384920 3207 384976
rect -960 384918 3207 384920
rect -960 384828 480 384918
rect 3141 384915 3207 384918
rect 579981 381578 580047 381581
rect 583520 381578 584960 381668
rect 579981 381576 584960 381578
rect 579981 381520 579986 381576
rect 580042 381520 584960 381576
rect 579981 381518 584960 381520
rect 579981 381515 580047 381518
rect 583520 381428 584960 381518
rect -960 380898 480 380988
rect 3325 380898 3391 380901
rect -960 380896 3391 380898
rect -960 380840 3330 380896
rect 3386 380840 3391 380896
rect -960 380838 3391 380840
rect -960 380748 480 380838
rect 3325 380835 3391 380838
rect 580165 377498 580231 377501
rect 583520 377498 584960 377588
rect 580165 377496 584960 377498
rect 580165 377440 580170 377496
rect 580226 377440 584960 377496
rect 580165 377438 584960 377440
rect 580165 377435 580231 377438
rect 583520 377348 584960 377438
rect -960 376818 480 376908
rect 3325 376818 3391 376821
rect -960 376816 3391 376818
rect -960 376760 3330 376816
rect 3386 376760 3391 376816
rect -960 376758 3391 376760
rect -960 376668 480 376758
rect 3325 376755 3391 376758
rect 580165 373418 580231 373421
rect 583520 373418 584960 373508
rect 580165 373416 584960 373418
rect 580165 373360 580170 373416
rect 580226 373360 584960 373416
rect 580165 373358 584960 373360
rect 580165 373355 580231 373358
rect 583520 373268 584960 373358
rect -960 372738 480 372828
rect 3325 372738 3391 372741
rect -960 372736 3391 372738
rect -960 372680 3330 372736
rect 3386 372680 3391 372736
rect -960 372678 3391 372680
rect -960 372588 480 372678
rect 3325 372675 3391 372678
rect 580165 369338 580231 369341
rect 583520 369338 584960 369428
rect 580165 369336 584960 369338
rect 580165 369280 580170 369336
rect 580226 369280 584960 369336
rect 580165 369278 584960 369280
rect 580165 369275 580231 369278
rect 583520 369188 584960 369278
rect -960 368658 480 368748
rect 3325 368658 3391 368661
rect -960 368656 3391 368658
rect -960 368600 3330 368656
rect 3386 368600 3391 368656
rect -960 368598 3391 368600
rect -960 368508 480 368598
rect 3325 368595 3391 368598
rect 579613 365258 579679 365261
rect 583520 365258 584960 365348
rect 579613 365256 584960 365258
rect 579613 365200 579618 365256
rect 579674 365200 584960 365256
rect 579613 365198 584960 365200
rect 579613 365195 579679 365198
rect 583520 365108 584960 365198
rect -960 364578 480 364668
rect 3325 364578 3391 364581
rect -960 364576 3391 364578
rect -960 364520 3330 364576
rect 3386 364520 3391 364576
rect -960 364518 3391 364520
rect -960 364428 480 364518
rect 3325 364515 3391 364518
rect 579613 361178 579679 361181
rect 583520 361178 584960 361268
rect 579613 361176 584960 361178
rect 579613 361120 579618 361176
rect 579674 361120 584960 361176
rect 579613 361118 584960 361120
rect 579613 361115 579679 361118
rect 583520 361028 584960 361118
rect -960 360498 480 360588
rect 3325 360498 3391 360501
rect -960 360496 3391 360498
rect -960 360440 3330 360496
rect 3386 360440 3391 360496
rect -960 360438 3391 360440
rect -960 360348 480 360438
rect 3325 360435 3391 360438
rect 580165 357098 580231 357101
rect 583520 357098 584960 357188
rect 580165 357096 584960 357098
rect 580165 357040 580170 357096
rect 580226 357040 584960 357096
rect 580165 357038 584960 357040
rect 580165 357035 580231 357038
rect 583520 356948 584960 357038
rect -960 356418 480 356508
rect 3325 356418 3391 356421
rect -960 356416 3391 356418
rect -960 356360 3330 356416
rect 3386 356360 3391 356416
rect -960 356358 3391 356360
rect -960 356268 480 356358
rect 3325 356355 3391 356358
rect 579613 353698 579679 353701
rect 583520 353698 584960 353788
rect 579613 353696 584960 353698
rect 579613 353640 579618 353696
rect 579674 353640 584960 353696
rect 579613 353638 584960 353640
rect 579613 353635 579679 353638
rect 583520 353548 584960 353638
rect -960 352338 480 352428
rect 3233 352338 3299 352341
rect -960 352336 3299 352338
rect -960 352280 3238 352336
rect 3294 352280 3299 352336
rect -960 352278 3299 352280
rect -960 352188 480 352278
rect 3233 352275 3299 352278
rect 580165 349618 580231 349621
rect 583520 349618 584960 349708
rect 580165 349616 584960 349618
rect 580165 349560 580170 349616
rect 580226 349560 584960 349616
rect 580165 349558 584960 349560
rect 580165 349555 580231 349558
rect 583520 349468 584960 349558
rect -960 348938 480 349028
rect 3141 348938 3207 348941
rect -960 348936 3207 348938
rect -960 348880 3146 348936
rect 3202 348880 3207 348936
rect -960 348878 3207 348880
rect -960 348788 480 348878
rect 3141 348875 3207 348878
rect 580165 345538 580231 345541
rect 583520 345538 584960 345628
rect 580165 345536 584960 345538
rect 580165 345480 580170 345536
rect 580226 345480 584960 345536
rect 580165 345478 584960 345480
rect 580165 345475 580231 345478
rect 583520 345388 584960 345478
rect -960 344858 480 344948
rect 3325 344858 3391 344861
rect -960 344856 3391 344858
rect -960 344800 3330 344856
rect 3386 344800 3391 344856
rect -960 344798 3391 344800
rect -960 344708 480 344798
rect 3325 344795 3391 344798
rect 580165 341458 580231 341461
rect 583520 341458 584960 341548
rect 580165 341456 584960 341458
rect 580165 341400 580170 341456
rect 580226 341400 584960 341456
rect 580165 341398 584960 341400
rect 580165 341395 580231 341398
rect 583520 341308 584960 341398
rect -960 340778 480 340868
rect 3141 340778 3207 340781
rect -960 340776 3207 340778
rect -960 340720 3146 340776
rect 3202 340720 3207 340776
rect -960 340718 3207 340720
rect -960 340628 480 340718
rect 3141 340715 3207 340718
rect 579981 337378 580047 337381
rect 583520 337378 584960 337468
rect 579981 337376 584960 337378
rect 579981 337320 579986 337376
rect 580042 337320 584960 337376
rect 579981 337318 584960 337320
rect 579981 337315 580047 337318
rect 583520 337228 584960 337318
rect -960 336698 480 336788
rect 3325 336698 3391 336701
rect -960 336696 3391 336698
rect -960 336640 3330 336696
rect 3386 336640 3391 336696
rect -960 336638 3391 336640
rect -960 336548 480 336638
rect 3325 336635 3391 336638
rect 579981 333298 580047 333301
rect 583520 333298 584960 333388
rect 579981 333296 584960 333298
rect 579981 333240 579986 333296
rect 580042 333240 584960 333296
rect 579981 333238 584960 333240
rect 579981 333235 580047 333238
rect 583520 333148 584960 333238
rect -960 332618 480 332708
rect 3325 332618 3391 332621
rect -960 332616 3391 332618
rect -960 332560 3330 332616
rect 3386 332560 3391 332616
rect -960 332558 3391 332560
rect -960 332468 480 332558
rect 3325 332555 3391 332558
rect 583520 329068 584960 329308
rect -960 328538 480 328628
rect 3325 328538 3391 328541
rect -960 328536 3391 328538
rect -960 328480 3330 328536
rect 3386 328480 3391 328536
rect -960 328478 3391 328480
rect -960 328388 480 328478
rect 3325 328475 3391 328478
rect 583520 324988 584960 325228
rect -960 324458 480 324548
rect 3325 324458 3391 324461
rect -960 324456 3391 324458
rect -960 324400 3330 324456
rect 3386 324400 3391 324456
rect -960 324398 3391 324400
rect -960 324308 480 324398
rect 3325 324395 3391 324398
rect 579613 321058 579679 321061
rect 583520 321058 584960 321148
rect 579613 321056 584960 321058
rect 579613 321000 579618 321056
rect 579674 321000 584960 321056
rect 579613 320998 584960 321000
rect 579613 320995 579679 320998
rect 583520 320908 584960 320998
rect -960 320378 480 320468
rect 3141 320378 3207 320381
rect -960 320376 3207 320378
rect -960 320320 3146 320376
rect 3202 320320 3207 320376
rect -960 320318 3207 320320
rect -960 320228 480 320318
rect 3141 320315 3207 320318
rect 579613 316978 579679 316981
rect 583520 316978 584960 317068
rect 579613 316976 584960 316978
rect 579613 316920 579618 316976
rect 579674 316920 584960 316976
rect 579613 316918 584960 316920
rect 579613 316915 579679 316918
rect 583520 316828 584960 316918
rect -960 316298 480 316388
rect 3325 316298 3391 316301
rect -960 316296 3391 316298
rect -960 316240 3330 316296
rect 3386 316240 3391 316296
rect -960 316238 3391 316240
rect -960 316148 480 316238
rect 3325 316235 3391 316238
rect 580625 313578 580691 313581
rect 583520 313578 584960 313668
rect 580625 313576 584960 313578
rect 580625 313520 580630 313576
rect 580686 313520 584960 313576
rect 580625 313518 584960 313520
rect 580625 313515 580691 313518
rect 583520 313428 584960 313518
rect -960 312068 480 312308
rect 580165 309498 580231 309501
rect 583520 309498 584960 309588
rect 580165 309496 584960 309498
rect 580165 309440 580170 309496
rect 580226 309440 584960 309496
rect 580165 309438 584960 309440
rect 580165 309435 580231 309438
rect 583520 309348 584960 309438
rect -960 308818 480 308908
rect 3325 308818 3391 308821
rect -960 308816 3391 308818
rect -960 308760 3330 308816
rect 3386 308760 3391 308816
rect -960 308758 3391 308760
rect -960 308668 480 308758
rect 3325 308755 3391 308758
rect 579613 305418 579679 305421
rect 583520 305418 584960 305508
rect 579613 305416 584960 305418
rect 579613 305360 579618 305416
rect 579674 305360 584960 305416
rect 579613 305358 584960 305360
rect 579613 305355 579679 305358
rect 583520 305268 584960 305358
rect -960 304738 480 304828
rect 3049 304738 3115 304741
rect -960 304736 3115 304738
rect -960 304680 3054 304736
rect 3110 304680 3115 304736
rect -960 304678 3115 304680
rect -960 304588 480 304678
rect 3049 304675 3115 304678
rect 580625 301338 580691 301341
rect 583520 301338 584960 301428
rect 580625 301336 584960 301338
rect 580625 301280 580630 301336
rect 580686 301280 584960 301336
rect 580625 301278 584960 301280
rect 580625 301275 580691 301278
rect 583520 301188 584960 301278
rect -960 300658 480 300748
rect 3141 300658 3207 300661
rect -960 300656 3207 300658
rect -960 300600 3146 300656
rect 3202 300600 3207 300656
rect -960 300598 3207 300600
rect -960 300508 480 300598
rect 3141 300595 3207 300598
rect 580165 297258 580231 297261
rect 583520 297258 584960 297348
rect 580165 297256 584960 297258
rect 580165 297200 580170 297256
rect 580226 297200 584960 297256
rect 580165 297198 584960 297200
rect 580165 297195 580231 297198
rect 583520 297108 584960 297198
rect -960 296578 480 296668
rect 3325 296578 3391 296581
rect -960 296576 3391 296578
rect -960 296520 3330 296576
rect 3386 296520 3391 296576
rect -960 296518 3391 296520
rect -960 296428 480 296518
rect 3325 296515 3391 296518
rect 579981 293178 580047 293181
rect 583520 293178 584960 293268
rect 579981 293176 584960 293178
rect 579981 293120 579986 293176
rect 580042 293120 584960 293176
rect 579981 293118 584960 293120
rect 579981 293115 580047 293118
rect 583520 293028 584960 293118
rect -960 292498 480 292588
rect 3141 292498 3207 292501
rect -960 292496 3207 292498
rect -960 292440 3146 292496
rect 3202 292440 3207 292496
rect -960 292438 3207 292440
rect -960 292348 480 292438
rect 3141 292435 3207 292438
rect 579981 289098 580047 289101
rect 583520 289098 584960 289188
rect 579981 289096 584960 289098
rect 579981 289040 579986 289096
rect 580042 289040 584960 289096
rect 579981 289038 584960 289040
rect 579981 289035 580047 289038
rect 583520 288948 584960 289038
rect -960 288418 480 288508
rect 3325 288418 3391 288421
rect -960 288416 3391 288418
rect -960 288360 3330 288416
rect 3386 288360 3391 288416
rect -960 288358 3391 288360
rect -960 288268 480 288358
rect 3325 288355 3391 288358
rect 579061 285018 579127 285021
rect 583520 285018 584960 285108
rect 579061 285016 584960 285018
rect 579061 284960 579066 285016
rect 579122 284960 584960 285016
rect 579061 284958 584960 284960
rect 579061 284955 579127 284958
rect 583520 284868 584960 284958
rect -960 284338 480 284428
rect 3325 284338 3391 284341
rect -960 284336 3391 284338
rect -960 284280 3330 284336
rect 3386 284280 3391 284336
rect -960 284278 3391 284280
rect -960 284188 480 284278
rect 3325 284275 3391 284278
rect 580165 280938 580231 280941
rect 583520 280938 584960 281028
rect 580165 280936 584960 280938
rect 580165 280880 580170 280936
rect 580226 280880 584960 280936
rect 580165 280878 584960 280880
rect 580165 280875 580231 280878
rect 583520 280788 584960 280878
rect -960 280258 480 280348
rect 3325 280258 3391 280261
rect -960 280256 3391 280258
rect -960 280200 3330 280256
rect 3386 280200 3391 280256
rect -960 280198 3391 280200
rect -960 280108 480 280198
rect 3325 280195 3391 280198
rect 580165 276858 580231 276861
rect 583520 276858 584960 276948
rect 580165 276856 584960 276858
rect 580165 276800 580170 276856
rect 580226 276800 584960 276856
rect 580165 276798 584960 276800
rect 580165 276795 580231 276798
rect 583520 276708 584960 276798
rect -960 276028 480 276268
rect 580165 273458 580231 273461
rect 583520 273458 584960 273548
rect 580165 273456 584960 273458
rect 580165 273400 580170 273456
rect 580226 273400 584960 273456
rect 580165 273398 584960 273400
rect 580165 273395 580231 273398
rect 583520 273308 584960 273398
rect -960 272098 480 272188
rect 3141 272098 3207 272101
rect -960 272096 3207 272098
rect -960 272040 3146 272096
rect 3202 272040 3207 272096
rect -960 272038 3207 272040
rect -960 271948 480 272038
rect 3141 272035 3207 272038
rect 580625 269378 580691 269381
rect 583520 269378 584960 269468
rect 580625 269376 584960 269378
rect 580625 269320 580630 269376
rect 580686 269320 584960 269376
rect 580625 269318 584960 269320
rect 580625 269315 580691 269318
rect 583520 269228 584960 269318
rect -960 268548 480 268788
rect 580165 265298 580231 265301
rect 583520 265298 584960 265388
rect 580165 265296 584960 265298
rect 580165 265240 580170 265296
rect 580226 265240 584960 265296
rect 580165 265238 584960 265240
rect 580165 265235 580231 265238
rect 583520 265148 584960 265238
rect -960 264618 480 264708
rect 3325 264618 3391 264621
rect -960 264616 3391 264618
rect -960 264560 3330 264616
rect 3386 264560 3391 264616
rect -960 264558 3391 264560
rect -960 264468 480 264558
rect 3325 264555 3391 264558
rect 173065 263802 173131 263805
rect 191966 263802 191972 263804
rect 173065 263800 191972 263802
rect 173065 263744 173070 263800
rect 173126 263744 191972 263800
rect 173065 263742 191972 263744
rect 173065 263739 173131 263742
rect 191966 263740 191972 263742
rect 192036 263740 192042 263804
rect 118550 263604 118556 263668
rect 118620 263666 118626 263668
rect 130377 263666 130443 263669
rect 118620 263664 130443 263666
rect 118620 263608 130382 263664
rect 130438 263608 130443 263664
rect 118620 263606 130443 263608
rect 118620 263604 118626 263606
rect 130377 263603 130443 263606
rect 170581 263666 170647 263669
rect 171041 263666 171107 263669
rect 191782 263666 191788 263668
rect 170581 263664 191788 263666
rect 170581 263608 170586 263664
rect 170642 263608 171046 263664
rect 171102 263608 191788 263664
rect 170581 263606 191788 263608
rect 170581 263603 170647 263606
rect 171041 263603 171107 263606
rect 191782 263604 191788 263606
rect 191852 263604 191858 263668
rect 189901 263122 189967 263125
rect 483013 263122 483079 263125
rect 189901 263120 483079 263122
rect 189901 263064 189906 263120
rect 189962 263064 483018 263120
rect 483074 263064 483079 263120
rect 189901 263062 483079 263064
rect 189901 263059 189967 263062
rect 483013 263059 483079 263062
rect 198825 262986 198891 262989
rect 569953 262986 570019 262989
rect 198825 262984 570019 262986
rect 198825 262928 198830 262984
rect 198886 262928 569958 262984
rect 570014 262928 570019 262984
rect 198825 262926 570019 262928
rect 198825 262923 198891 262926
rect 569953 262923 570019 262926
rect 115381 262850 115447 262853
rect 126973 262850 127039 262853
rect 546493 262850 546559 262853
rect 115381 262848 127039 262850
rect 115381 262792 115386 262848
rect 115442 262792 126978 262848
rect 127034 262792 127039 262848
rect 115381 262790 127039 262792
rect 115381 262787 115447 262790
rect 126973 262787 127039 262790
rect 142110 262848 546559 262850
rect 142110 262792 546498 262848
rect 546554 262792 546559 262848
rect 142110 262790 546559 262792
rect 112805 262442 112871 262445
rect 141233 262442 141299 262445
rect 142110 262442 142170 262790
rect 546493 262787 546559 262790
rect 154481 262578 154547 262581
rect 189901 262578 189967 262581
rect 154481 262576 189967 262578
rect 154481 262520 154486 262576
rect 154542 262520 189906 262576
rect 189962 262520 189967 262576
rect 154481 262518 189967 262520
rect 154481 262515 154547 262518
rect 189901 262515 189967 262518
rect 112805 262440 142170 262442
rect 112805 262384 112810 262440
rect 112866 262384 141238 262440
rect 141294 262384 142170 262440
rect 112805 262382 142170 262384
rect 166901 262442 166967 262445
rect 198825 262442 198891 262445
rect 199101 262442 199167 262445
rect 166901 262440 199167 262442
rect 166901 262384 166906 262440
rect 166962 262384 198830 262440
rect 198886 262384 199106 262440
rect 199162 262384 199167 262440
rect 166901 262382 199167 262384
rect 112805 262379 112871 262382
rect 141233 262379 141299 262382
rect 166901 262379 166967 262382
rect 198825 262379 198891 262382
rect 199101 262379 199167 262382
rect 580717 261218 580783 261221
rect 583520 261218 584960 261308
rect 580717 261216 584960 261218
rect 580717 261160 580722 261216
rect 580778 261160 584960 261216
rect 580717 261158 584960 261160
rect 580717 261155 580783 261158
rect 583520 261068 584960 261158
rect -960 260538 480 260628
rect 3049 260538 3115 260541
rect -960 260536 3115 260538
rect -960 260480 3054 260536
rect 3110 260480 3115 260536
rect -960 260478 3115 260480
rect -960 260388 480 260478
rect 3049 260475 3115 260478
rect 171133 260130 171199 260133
rect 189993 260130 190059 260133
rect 171133 260128 190059 260130
rect 171133 260072 171138 260128
rect 171194 260072 189998 260128
rect 190054 260072 190059 260128
rect 171133 260070 190059 260072
rect 171133 260067 171199 260070
rect 189993 260067 190059 260070
rect 184933 259994 184999 259997
rect 185853 259994 185919 259997
rect 186998 259994 187004 259996
rect 184933 259992 187004 259994
rect 184933 259936 184938 259992
rect 184994 259936 185858 259992
rect 185914 259936 187004 259992
rect 184933 259934 187004 259936
rect 184933 259931 184999 259934
rect 185853 259931 185919 259934
rect 186998 259932 187004 259934
rect 187068 259932 187074 259996
rect 154021 259722 154087 259725
rect 187918 259722 187924 259724
rect 154021 259720 187924 259722
rect 154021 259664 154026 259720
rect 154082 259664 187924 259720
rect 154021 259662 187924 259664
rect 154021 259659 154087 259662
rect 187918 259660 187924 259662
rect 187988 259722 187994 259724
rect 187988 259662 190470 259722
rect 187988 259660 187994 259662
rect 122557 259588 122623 259589
rect 187141 259588 187207 259589
rect 122557 259584 122604 259588
rect 122668 259586 122674 259588
rect 122557 259528 122562 259584
rect 122557 259524 122604 259528
rect 122668 259526 122714 259586
rect 187141 259584 187188 259588
rect 187252 259586 187258 259588
rect 190410 259586 190470 259662
rect 576393 259586 576459 259589
rect 187141 259528 187146 259584
rect 122668 259524 122674 259526
rect 187141 259524 187188 259528
rect 187252 259526 187298 259586
rect 190410 259584 576459 259586
rect 190410 259528 576398 259584
rect 576454 259528 576459 259584
rect 190410 259526 576459 259528
rect 187252 259524 187258 259526
rect 122557 259523 122623 259524
rect 187141 259523 187207 259524
rect 576393 259523 576459 259526
rect 580257 257138 580323 257141
rect 583520 257138 584960 257228
rect 580257 257136 584960 257138
rect 580257 257080 580262 257136
rect 580318 257080 584960 257136
rect 580257 257078 584960 257080
rect 580257 257075 580323 257078
rect 583520 256988 584960 257078
rect -960 256458 480 256548
rect 3141 256458 3207 256461
rect -960 256456 3207 256458
rect -960 256400 3146 256456
rect 3202 256400 3207 256456
rect -960 256398 3207 256400
rect -960 256308 480 256398
rect 3141 256395 3207 256398
rect 579797 253058 579863 253061
rect 583520 253058 584960 253148
rect 579797 253056 584960 253058
rect 579797 253000 579802 253056
rect 579858 253000 584960 253056
rect 579797 252998 584960 253000
rect 579797 252995 579863 252998
rect 583520 252908 584960 252998
rect -960 252378 480 252468
rect 3141 252378 3207 252381
rect -960 252376 3207 252378
rect -960 252320 3146 252376
rect 3202 252320 3207 252376
rect -960 252318 3207 252320
rect -960 252228 480 252318
rect 3141 252315 3207 252318
rect 579797 248978 579863 248981
rect 583520 248978 584960 249068
rect 579797 248976 584960 248978
rect 579797 248920 579802 248976
rect 579858 248920 584960 248976
rect 579797 248918 584960 248920
rect 579797 248915 579863 248918
rect 583520 248828 584960 248918
rect -960 248298 480 248388
rect 3325 248298 3391 248301
rect -960 248296 3391 248298
rect -960 248240 3330 248296
rect 3386 248240 3391 248296
rect -960 248238 3391 248240
rect -960 248148 480 248238
rect 3325 248235 3391 248238
rect 580165 244898 580231 244901
rect 583520 244898 584960 244988
rect 580165 244896 584960 244898
rect 580165 244840 580170 244896
rect 580226 244840 584960 244896
rect 580165 244838 584960 244840
rect 580165 244835 580231 244838
rect 583520 244748 584960 244838
rect -960 244218 480 244308
rect 3141 244218 3207 244221
rect -960 244216 3207 244218
rect -960 244160 3146 244216
rect 3202 244160 3207 244216
rect -960 244158 3207 244160
rect -960 244068 480 244158
rect 3141 244155 3207 244158
rect 580717 240818 580783 240821
rect 583520 240818 584960 240908
rect 580717 240816 584960 240818
rect 580717 240760 580722 240816
rect 580778 240760 584960 240816
rect 580717 240758 584960 240760
rect 580717 240755 580783 240758
rect 583520 240668 584960 240758
rect -960 240138 480 240228
rect 3325 240138 3391 240141
rect -960 240136 3391 240138
rect -960 240080 3330 240136
rect 3386 240080 3391 240136
rect -960 240078 3391 240080
rect -960 239988 480 240078
rect 3325 240075 3391 240078
rect 580165 237418 580231 237421
rect 583520 237418 584960 237508
rect 580165 237416 584960 237418
rect 580165 237360 580170 237416
rect 580226 237360 584960 237416
rect 580165 237358 584960 237360
rect 580165 237355 580231 237358
rect 583520 237268 584960 237358
rect -960 236058 480 236148
rect 3325 236058 3391 236061
rect -960 236056 3391 236058
rect -960 236000 3330 236056
rect 3386 236000 3391 236056
rect -960 235998 3391 236000
rect -960 235908 480 235998
rect 3325 235995 3391 235998
rect 188286 233276 188292 233340
rect 188356 233338 188362 233340
rect 583520 233338 584960 233428
rect 188356 233278 584960 233338
rect 188356 233276 188362 233278
rect 583520 233188 584960 233278
rect -960 232658 480 232748
rect 3325 232658 3391 232661
rect -960 232656 3391 232658
rect -960 232600 3330 232656
rect 3386 232600 3391 232656
rect -960 232598 3391 232600
rect -960 232508 480 232598
rect 3325 232595 3391 232598
rect 583520 229108 584960 229348
rect -960 228578 480 228668
rect 3325 228578 3391 228581
rect -960 228576 3391 228578
rect -960 228520 3330 228576
rect 3386 228520 3391 228576
rect -960 228518 3391 228520
rect -960 228428 480 228518
rect 3325 228515 3391 228518
rect 92473 227762 92539 227765
rect 93761 227762 93827 227765
rect 122046 227762 122052 227764
rect 92473 227760 122052 227762
rect 92473 227704 92478 227760
rect 92534 227704 93766 227760
rect 93822 227704 122052 227760
rect 92473 227702 122052 227704
rect 92473 227699 92539 227702
rect 93761 227699 93827 227702
rect 122046 227700 122052 227702
rect 122116 227700 122122 227764
rect 580809 225178 580875 225181
rect 583520 225178 584960 225268
rect 580809 225176 584960 225178
rect 580809 225120 580814 225176
rect 580870 225120 584960 225176
rect 580809 225118 584960 225120
rect 580809 225115 580875 225118
rect 583520 225028 584960 225118
rect -960 224498 480 224588
rect 3325 224498 3391 224501
rect -960 224496 3391 224498
rect -960 224440 3330 224496
rect 3386 224440 3391 224496
rect -960 224438 3391 224440
rect -960 224348 480 224438
rect 3325 224435 3391 224438
rect 120625 223546 120691 223549
rect 120993 223546 121059 223549
rect 120625 223544 121059 223546
rect 120625 223488 120630 223544
rect 120686 223488 120998 223544
rect 121054 223488 121059 223544
rect 120625 223486 121059 223488
rect 120625 223483 120691 223486
rect 120993 223483 121059 223486
rect 580165 221098 580231 221101
rect 583520 221098 584960 221188
rect 580165 221096 584960 221098
rect 580165 221040 580170 221096
rect 580226 221040 584960 221096
rect 580165 221038 584960 221040
rect 580165 221035 580231 221038
rect 186814 220900 186820 220964
rect 186884 220962 186890 220964
rect 208393 220962 208459 220965
rect 186884 220960 208459 220962
rect 186884 220904 208398 220960
rect 208454 220904 208459 220960
rect 583520 220948 584960 221038
rect 186884 220902 208459 220904
rect 186884 220900 186890 220902
rect 208393 220899 208459 220902
rect -960 220418 480 220508
rect 3233 220418 3299 220421
rect -960 220416 3299 220418
rect -960 220360 3238 220416
rect 3294 220360 3299 220416
rect -960 220358 3299 220360
rect -960 220268 480 220358
rect 3233 220355 3299 220358
rect 580165 217018 580231 217021
rect 583520 217018 584960 217108
rect 580165 217016 584960 217018
rect 580165 216960 580170 217016
rect 580226 216960 584960 217016
rect 580165 216958 584960 216960
rect 580165 216955 580231 216958
rect 583520 216868 584960 216958
rect -960 216338 480 216428
rect 3325 216338 3391 216341
rect -960 216336 3391 216338
rect -960 216280 3330 216336
rect 3386 216280 3391 216336
rect -960 216278 3391 216280
rect -960 216188 480 216278
rect 3325 216275 3391 216278
rect 583520 212788 584960 213028
rect -960 212258 480 212348
rect -960 212198 674 212258
rect -960 212122 480 212198
rect 614 212122 674 212198
rect -960 212108 674 212122
rect 246 212062 674 212108
rect 246 211578 306 212062
rect 246 211518 6930 211578
rect 6870 211170 6930 211518
rect 122230 211170 122236 211172
rect 6870 211110 122236 211170
rect 122230 211108 122236 211110
rect 122300 211108 122306 211172
rect 583520 208858 584960 208948
rect 583342 208798 584960 208858
rect 583342 208722 583402 208798
rect 583520 208722 584960 208798
rect 583342 208708 584960 208722
rect 583342 208662 583586 208708
rect 186262 208388 186268 208452
rect 186332 208450 186338 208452
rect 583526 208450 583586 208662
rect 186332 208390 583586 208450
rect 186332 208388 186338 208390
rect -960 208178 480 208268
rect -960 208118 674 208178
rect -960 208042 480 208118
rect 614 208042 674 208118
rect -960 208028 674 208042
rect 246 207982 674 208028
rect 246 207498 306 207982
rect 246 207438 6930 207498
rect 6870 207090 6930 207438
rect 121862 207090 121868 207092
rect 6870 207030 121868 207090
rect 121862 207028 121868 207030
rect 121932 207028 121938 207092
rect 579981 204778 580047 204781
rect 583520 204778 584960 204868
rect 579981 204776 584960 204778
rect 579981 204720 579986 204776
rect 580042 204720 584960 204776
rect 579981 204718 584960 204720
rect 579981 204715 580047 204718
rect 583520 204628 584960 204718
rect -960 203948 480 204188
rect 209313 202194 209379 202197
rect 558177 202194 558243 202197
rect 209313 202192 558243 202194
rect 209313 202136 209318 202192
rect 209374 202136 558182 202192
rect 558238 202136 558243 202192
rect 209313 202134 558243 202136
rect 209313 202131 209379 202134
rect 558177 202131 558243 202134
rect 176326 201452 176332 201516
rect 176396 201514 176402 201516
rect 208485 201514 208551 201517
rect 209313 201514 209379 201517
rect 176396 201512 209379 201514
rect 176396 201456 208490 201512
rect 208546 201456 209318 201512
rect 209374 201456 209379 201512
rect 176396 201454 209379 201456
rect 176396 201452 176402 201454
rect 208485 201451 208551 201454
rect 209313 201451 209379 201454
rect 98729 200970 98795 200973
rect 111793 200970 111859 200973
rect 98729 200968 111859 200970
rect 98729 200912 98734 200968
rect 98790 200912 111798 200968
rect 111854 200912 111859 200968
rect 98729 200910 111859 200912
rect 98729 200907 98795 200910
rect 111793 200907 111859 200910
rect 122046 200908 122052 200972
rect 122116 200970 122122 200972
rect 122116 200910 138030 200970
rect 122116 200908 122122 200910
rect 79317 200834 79383 200837
rect 121494 200834 121500 200836
rect 79317 200832 121500 200834
rect 79317 200776 79322 200832
rect 79378 200776 121500 200832
rect 79317 200774 121500 200776
rect 79317 200771 79383 200774
rect 121494 200772 121500 200774
rect 121564 200772 121570 200836
rect 137970 200834 138030 200910
rect 156822 200834 156828 200836
rect 137970 200774 156828 200834
rect 156822 200772 156828 200774
rect 156892 200772 156898 200836
rect 168230 200772 168236 200836
rect 168300 200834 168306 200836
rect 186814 200834 186820 200836
rect 168300 200774 186820 200834
rect 168300 200772 168306 200774
rect 186814 200772 186820 200774
rect 186884 200772 186890 200836
rect 203006 200772 203012 200836
rect 203076 200834 203082 200836
rect 422293 200834 422359 200837
rect 203076 200832 422359 200834
rect 203076 200776 422298 200832
rect 422354 200776 422359 200832
rect 203076 200774 422359 200776
rect 203076 200772 203082 200774
rect 422293 200771 422359 200774
rect 48957 200698 49023 200701
rect 107561 200698 107627 200701
rect 48957 200696 107627 200698
rect 48957 200640 48962 200696
rect 49018 200640 107566 200696
rect 107622 200640 107627 200696
rect 48957 200638 107627 200640
rect 48957 200635 49023 200638
rect 107561 200635 107627 200638
rect 117773 200698 117839 200701
rect 138606 200698 138612 200700
rect 117773 200696 138612 200698
rect 117773 200640 117778 200696
rect 117834 200640 138612 200696
rect 117773 200638 138612 200640
rect 117773 200635 117839 200638
rect 138606 200636 138612 200638
rect 138676 200636 138682 200700
rect 152406 200636 152412 200700
rect 152476 200698 152482 200700
rect 186078 200698 186084 200700
rect 152476 200638 186084 200698
rect 152476 200636 152482 200638
rect 186078 200636 186084 200638
rect 186148 200636 186154 200700
rect 187182 200636 187188 200700
rect 187252 200698 187258 200700
rect 187601 200698 187667 200701
rect 187252 200696 187667 200698
rect 187252 200640 187606 200696
rect 187662 200640 187667 200696
rect 187252 200638 187667 200640
rect 187252 200636 187258 200638
rect 187601 200635 187667 200638
rect 207054 200636 207060 200700
rect 207124 200698 207130 200700
rect 514017 200698 514083 200701
rect 207124 200696 514083 200698
rect 207124 200640 514022 200696
rect 514078 200640 514083 200696
rect 207124 200638 514083 200640
rect 207124 200636 207130 200638
rect 514017 200635 514083 200638
rect 580165 200698 580231 200701
rect 583520 200698 584960 200788
rect 580165 200696 584960 200698
rect 580165 200640 580170 200696
rect 580226 200640 584960 200696
rect 580165 200638 584960 200640
rect 580165 200635 580231 200638
rect 131665 200562 131731 200565
rect 138238 200562 138244 200564
rect 131665 200560 138244 200562
rect 131665 200504 131670 200560
rect 131726 200504 138244 200560
rect 131665 200502 138244 200504
rect 131665 200499 131731 200502
rect 138238 200500 138244 200502
rect 138308 200500 138314 200564
rect 173014 200500 173020 200564
rect 173084 200562 173090 200564
rect 178401 200562 178467 200565
rect 173084 200560 178467 200562
rect 173084 200504 178406 200560
rect 178462 200504 178467 200560
rect 583520 200548 584960 200638
rect 173084 200502 178467 200504
rect 173084 200500 173090 200502
rect 178401 200499 178467 200502
rect 111793 200426 111859 200429
rect 113081 200426 113147 200429
rect 145598 200426 145604 200428
rect 111793 200424 145604 200426
rect 111793 200368 111798 200424
rect 111854 200368 113086 200424
rect 113142 200368 145604 200424
rect 111793 200366 145604 200368
rect 111793 200363 111859 200366
rect 113081 200363 113147 200366
rect 145598 200364 145604 200366
rect 145668 200364 145674 200428
rect 176142 200364 176148 200428
rect 176212 200426 176218 200428
rect 177757 200426 177823 200429
rect 176212 200424 177823 200426
rect 176212 200368 177762 200424
rect 177818 200368 177823 200424
rect 176212 200366 177823 200368
rect 176212 200364 176218 200366
rect 177757 200363 177823 200366
rect 107561 200290 107627 200293
rect 139342 200290 139348 200292
rect 107561 200288 139348 200290
rect 107561 200232 107566 200288
rect 107622 200232 139348 200288
rect 107561 200230 139348 200232
rect 107561 200227 107627 200230
rect 139342 200228 139348 200230
rect 139412 200228 139418 200292
rect 147630 200230 159466 200290
rect -960 200018 480 200108
rect 121494 200092 121500 200156
rect 121564 200154 121570 200156
rect 122414 200154 122420 200156
rect 121564 200094 122420 200154
rect 121564 200092 121570 200094
rect 122414 200092 122420 200094
rect 122484 200154 122490 200156
rect 147630 200154 147690 200230
rect 122484 200094 147690 200154
rect 122484 200092 122490 200094
rect 147990 200092 147996 200156
rect 148060 200154 148066 200156
rect 149462 200154 149468 200156
rect 148060 200094 149468 200154
rect 148060 200092 148066 200094
rect 149462 200092 149468 200094
rect 149532 200092 149538 200156
rect 153326 200092 153332 200156
rect 153396 200154 153402 200156
rect 154430 200154 154436 200156
rect 153396 200094 154436 200154
rect 153396 200092 153402 200094
rect 154430 200092 154436 200094
rect 154500 200092 154506 200156
rect 3509 200018 3575 200021
rect -960 200016 3575 200018
rect -960 199960 3514 200016
rect 3570 199960 3575 200016
rect -960 199958 3575 199960
rect -960 199868 480 199958
rect 3509 199955 3575 199958
rect 129733 200018 129799 200021
rect 129733 200016 134626 200018
rect 129733 199960 129738 200016
rect 129794 199960 134626 200016
rect 129733 199958 134626 199960
rect 129733 199955 129799 199958
rect 128353 199882 128419 199885
rect 132723 199882 132789 199885
rect 133091 199884 133157 199885
rect 133086 199882 133092 199884
rect 128353 199880 132789 199882
rect 128353 199824 128358 199880
rect 128414 199824 132728 199880
rect 132784 199824 132789 199880
rect 128353 199822 132789 199824
rect 133000 199822 133092 199882
rect 128353 199819 128419 199822
rect 132723 199819 132789 199822
rect 133086 199820 133092 199822
rect 133156 199820 133162 199884
rect 133270 199820 133276 199884
rect 133340 199882 133346 199884
rect 133551 199882 133617 199885
rect 133340 199880 133617 199882
rect 133340 199824 133556 199880
rect 133612 199824 133617 199880
rect 133340 199822 133617 199824
rect 133340 199820 133346 199822
rect 133091 199819 133157 199820
rect 133551 199819 133617 199822
rect 133822 199820 133828 199884
rect 133892 199882 133898 199884
rect 134103 199882 134169 199885
rect 134379 199884 134445 199885
rect 134374 199882 134380 199884
rect 133892 199880 134169 199882
rect 133892 199824 134108 199880
rect 134164 199824 134169 199880
rect 133892 199822 134169 199824
rect 134288 199822 134380 199882
rect 133892 199820 133898 199822
rect 134103 199819 134169 199822
rect 134374 199820 134380 199822
rect 134444 199820 134450 199884
rect 134566 199882 134626 199958
rect 138054 199956 138060 200020
rect 138124 200018 138130 200020
rect 138124 199958 138306 200018
rect 138124 199956 138130 199958
rect 134747 199914 134813 199919
rect 134747 199882 134752 199914
rect 134566 199858 134752 199882
rect 134808 199858 134813 199914
rect 136219 199914 136285 199919
rect 134566 199853 134813 199858
rect 134566 199822 134810 199853
rect 136030 199820 136036 199884
rect 136100 199882 136106 199884
rect 136219 199882 136224 199914
rect 136100 199858 136224 199882
rect 136280 199858 136285 199914
rect 137323 199914 137389 199919
rect 137323 199884 137328 199914
rect 137384 199884 137389 199914
rect 137875 199914 137941 199919
rect 136100 199853 136285 199858
rect 136100 199822 136282 199853
rect 136100 199820 136106 199822
rect 137318 199820 137324 199884
rect 137388 199882 137394 199884
rect 137388 199822 137446 199882
rect 137875 199858 137880 199914
rect 137936 199882 137941 199914
rect 138054 199882 138060 199884
rect 137936 199858 138060 199882
rect 137875 199853 138060 199858
rect 137878 199822 138060 199853
rect 137388 199820 137394 199822
rect 138054 199820 138060 199822
rect 138124 199820 138130 199884
rect 138246 199882 138306 199958
rect 159406 199919 159466 200230
rect 160318 200228 160324 200292
rect 160388 200290 160394 200292
rect 161606 200290 161612 200292
rect 160388 200230 161612 200290
rect 160388 200228 160394 200230
rect 161606 200228 161612 200230
rect 161676 200228 161682 200292
rect 203006 200290 203012 200292
rect 170722 200230 203012 200290
rect 160502 200092 160508 200156
rect 160572 200154 160578 200156
rect 161422 200154 161428 200156
rect 160572 200094 161428 200154
rect 160572 200092 160578 200094
rect 161422 200092 161428 200094
rect 161492 200092 161498 200156
rect 170722 199919 170782 200230
rect 203006 200228 203012 200230
rect 203076 200228 203082 200292
rect 177062 200154 177068 200156
rect 174632 200094 177068 200154
rect 138427 199914 138493 199919
rect 138427 199882 138432 199914
rect 138246 199858 138432 199882
rect 138488 199858 138493 199914
rect 138246 199853 138493 199858
rect 138795 199914 138861 199919
rect 139255 199916 139321 199919
rect 138795 199858 138800 199914
rect 138856 199882 138861 199914
rect 139212 199914 139321 199916
rect 139212 199884 139260 199914
rect 138974 199882 138980 199884
rect 138856 199858 138980 199882
rect 138795 199853 138980 199858
rect 138246 199822 138490 199853
rect 138798 199822 138980 199853
rect 138974 199820 138980 199822
rect 139044 199820 139050 199884
rect 139158 199820 139164 199884
rect 139228 199858 139260 199884
rect 139316 199858 139321 199914
rect 139531 199914 139597 199919
rect 139531 199884 139536 199914
rect 139592 199884 139597 199914
rect 139899 199914 139965 199919
rect 139899 199884 139904 199914
rect 139960 199884 139965 199914
rect 140267 199914 140333 199919
rect 140267 199884 140272 199914
rect 140328 199884 140333 199914
rect 140635 199914 140701 199919
rect 140635 199884 140640 199914
rect 140696 199884 140701 199914
rect 142199 199916 142265 199919
rect 142475 199916 142541 199919
rect 142843 199916 142909 199919
rect 142199 199914 142308 199916
rect 139228 199853 139321 199858
rect 139228 199822 139272 199853
rect 139228 199820 139234 199822
rect 139526 199820 139532 199884
rect 139596 199882 139602 199884
rect 139596 199822 139654 199882
rect 139596 199820 139602 199822
rect 139894 199820 139900 199884
rect 139964 199882 139970 199884
rect 139964 199822 140022 199882
rect 139964 199820 139970 199822
rect 140262 199820 140268 199884
rect 140332 199882 140338 199884
rect 140332 199822 140390 199882
rect 140332 199820 140338 199822
rect 140630 199820 140636 199884
rect 140700 199882 140706 199884
rect 140700 199822 140758 199882
rect 140700 199820 140706 199822
rect 141182 199820 141188 199884
rect 141252 199882 141258 199884
rect 142199 199882 142204 199914
rect 141252 199858 142204 199882
rect 142260 199858 142308 199914
rect 142475 199914 142598 199916
rect 142475 199884 142480 199914
rect 142536 199884 142598 199914
rect 141252 199822 142308 199858
rect 141252 199820 141258 199822
rect 142470 199820 142476 199884
rect 142540 199856 142598 199884
rect 142843 199914 143090 199916
rect 142843 199858 142848 199914
rect 142904 199884 143090 199914
rect 144315 199914 144381 199919
rect 144315 199884 144320 199914
rect 144376 199884 144381 199914
rect 144591 199916 144657 199919
rect 144591 199914 144930 199916
rect 142904 199858 143028 199884
rect 142843 199856 143028 199858
rect 142540 199820 142546 199856
rect 142843 199853 142909 199856
rect 143022 199820 143028 199856
rect 143092 199820 143098 199884
rect 144310 199820 144316 199884
rect 144380 199882 144386 199884
rect 144380 199822 144438 199882
rect 144591 199858 144596 199914
rect 144652 199884 144930 199914
rect 145051 199914 145117 199919
rect 144652 199858 144868 199884
rect 144591 199856 144868 199858
rect 144591 199853 144657 199856
rect 144380 199820 144386 199822
rect 144862 199820 144868 199856
rect 144932 199820 144938 199884
rect 145051 199858 145056 199914
rect 145112 199882 145117 199914
rect 145603 199914 145669 199919
rect 145603 199884 145608 199914
rect 145664 199884 145669 199914
rect 146155 199914 146221 199919
rect 146155 199884 146160 199914
rect 146216 199884 146221 199914
rect 146799 199914 146865 199919
rect 145414 199882 145420 199884
rect 145112 199858 145420 199882
rect 145051 199853 145420 199858
rect 145054 199822 145420 199853
rect 145414 199820 145420 199822
rect 145484 199820 145490 199884
rect 145598 199820 145604 199884
rect 145668 199882 145674 199884
rect 145668 199822 145726 199882
rect 145668 199820 145674 199822
rect 146150 199820 146156 199884
rect 146220 199882 146226 199884
rect 146220 199822 146278 199882
rect 146220 199820 146226 199822
rect 146518 199820 146524 199884
rect 146588 199882 146594 199884
rect 146799 199882 146804 199914
rect 146588 199858 146804 199882
rect 146860 199858 146865 199914
rect 147811 199914 147877 199919
rect 147811 199884 147816 199914
rect 147872 199884 147877 199914
rect 148271 199916 148337 199919
rect 148271 199914 148380 199916
rect 146588 199853 146865 199858
rect 146588 199822 146862 199853
rect 146588 199820 146594 199822
rect 147806 199820 147812 199884
rect 147876 199882 147882 199884
rect 147876 199822 147934 199882
rect 148271 199858 148276 199914
rect 148332 199884 148380 199914
rect 148547 199914 148613 199919
rect 148547 199884 148552 199914
rect 148608 199884 148613 199914
rect 148915 199914 148981 199919
rect 148915 199884 148920 199914
rect 148976 199884 148981 199914
rect 149099 199914 149165 199919
rect 148332 199858 148364 199884
rect 148271 199853 148364 199858
rect 148320 199822 148364 199853
rect 147876 199820 147882 199822
rect 148358 199820 148364 199822
rect 148428 199820 148434 199884
rect 148542 199820 148548 199884
rect 148612 199882 148618 199884
rect 148612 199822 148670 199882
rect 148612 199820 148618 199822
rect 148910 199820 148916 199884
rect 148980 199882 148986 199884
rect 148980 199822 149038 199882
rect 149099 199858 149104 199914
rect 149160 199882 149165 199914
rect 149651 199914 149717 199919
rect 149651 199884 149656 199914
rect 149712 199884 149717 199914
rect 150203 199914 150269 199919
rect 150203 199884 150208 199914
rect 150264 199884 150269 199914
rect 151123 199914 151189 199919
rect 151767 199916 151833 199919
rect 149278 199882 149284 199884
rect 149160 199858 149284 199882
rect 149099 199853 149284 199858
rect 149102 199822 149284 199853
rect 148980 199820 148986 199822
rect 149278 199820 149284 199822
rect 149348 199820 149354 199884
rect 149646 199820 149652 199884
rect 149716 199882 149722 199884
rect 149716 199822 149774 199882
rect 149716 199820 149722 199822
rect 150198 199820 150204 199884
rect 150268 199882 150274 199884
rect 150268 199822 150326 199882
rect 150268 199820 150274 199822
rect 150566 199820 150572 199884
rect 150636 199882 150642 199884
rect 151123 199882 151128 199914
rect 150636 199858 151128 199882
rect 151184 199858 151189 199914
rect 151494 199914 151833 199916
rect 151494 199884 151772 199914
rect 150636 199853 151189 199858
rect 150636 199822 151186 199853
rect 150636 199820 150642 199822
rect 151486 199820 151492 199884
rect 151556 199858 151772 199884
rect 151828 199858 151833 199914
rect 152043 199914 152109 199919
rect 152043 199884 152048 199914
rect 152104 199884 152109 199914
rect 152411 199916 152477 199919
rect 153147 199916 153213 199919
rect 152411 199914 152534 199916
rect 152411 199884 152416 199914
rect 152472 199884 152534 199914
rect 153147 199914 153270 199916
rect 153147 199884 153152 199914
rect 153208 199884 153270 199914
rect 153515 199914 153581 199919
rect 153515 199884 153520 199914
rect 153576 199884 153581 199914
rect 154251 199914 154317 199919
rect 154251 199884 154256 199914
rect 154312 199884 154317 199914
rect 154803 199914 154869 199919
rect 154803 199884 154808 199914
rect 154864 199884 154869 199914
rect 156827 199916 156893 199919
rect 157839 199916 157905 199919
rect 156827 199914 156950 199916
rect 156827 199884 156832 199914
rect 156888 199884 156950 199914
rect 151556 199856 151833 199858
rect 151556 199820 151562 199856
rect 151767 199853 151833 199856
rect 152038 199820 152044 199884
rect 152108 199882 152114 199884
rect 152108 199822 152166 199882
rect 152108 199820 152114 199822
rect 152406 199820 152412 199884
rect 152476 199856 152534 199884
rect 152476 199820 152482 199856
rect 153142 199820 153148 199884
rect 153212 199856 153270 199884
rect 153212 199820 153218 199856
rect 153510 199820 153516 199884
rect 153580 199882 153586 199884
rect 153580 199822 153638 199882
rect 153580 199820 153586 199822
rect 154246 199820 154252 199884
rect 154316 199882 154322 199884
rect 154316 199822 154374 199882
rect 154316 199820 154322 199822
rect 154798 199820 154804 199884
rect 154868 199882 154874 199884
rect 154868 199822 154926 199882
rect 154868 199820 154874 199822
rect 156822 199820 156828 199884
rect 156892 199856 156950 199884
rect 157796 199914 157905 199916
rect 157796 199858 157844 199914
rect 157900 199882 157905 199914
rect 158851 199914 158917 199919
rect 158851 199884 158856 199914
rect 158912 199884 158917 199914
rect 159035 199914 159101 199919
rect 158294 199882 158300 199884
rect 157900 199858 158300 199882
rect 156892 199820 156898 199856
rect 157796 199822 158300 199858
rect 158294 199820 158300 199822
rect 158364 199820 158370 199884
rect 158846 199820 158852 199884
rect 158916 199882 158922 199884
rect 158916 199822 158974 199882
rect 159035 199858 159040 199914
rect 159096 199882 159101 199914
rect 159403 199914 159469 199919
rect 159214 199882 159220 199884
rect 159096 199858 159220 199882
rect 159035 199853 159220 199858
rect 159038 199822 159220 199853
rect 158916 199820 158922 199822
rect 159214 199820 159220 199822
rect 159284 199820 159290 199884
rect 159403 199858 159408 199914
rect 159464 199858 159469 199914
rect 159403 199853 159469 199858
rect 160231 199916 160297 199919
rect 160231 199914 160570 199916
rect 160231 199858 160236 199914
rect 160292 199882 160570 199914
rect 161243 199914 161309 199919
rect 161243 199884 161248 199914
rect 161304 199884 161309 199914
rect 161703 199914 161769 199919
rect 160870 199882 160876 199884
rect 160292 199858 160876 199882
rect 160231 199856 160876 199858
rect 160231 199853 160297 199856
rect 160510 199822 160876 199856
rect 160870 199820 160876 199822
rect 160940 199820 160946 199884
rect 161238 199820 161244 199884
rect 161308 199882 161314 199884
rect 161308 199822 161366 199882
rect 161703 199858 161708 199914
rect 161764 199882 161769 199914
rect 162255 199916 162321 199919
rect 162255 199914 162548 199916
rect 161974 199882 161980 199884
rect 161764 199858 161980 199882
rect 161703 199853 161980 199858
rect 161706 199822 161980 199853
rect 161308 199820 161314 199822
rect 161974 199820 161980 199822
rect 162044 199820 162050 199884
rect 162255 199858 162260 199914
rect 162316 199884 162548 199914
rect 162899 199914 162965 199919
rect 163911 199916 163977 199919
rect 162899 199884 162904 199914
rect 162960 199884 162965 199914
rect 163868 199914 163977 199916
rect 163868 199884 163916 199914
rect 162316 199858 162532 199884
rect 162255 199856 162532 199858
rect 162255 199853 162321 199856
rect 162488 199822 162532 199856
rect 162526 199820 162532 199822
rect 162596 199820 162602 199884
rect 162894 199820 162900 199884
rect 162964 199882 162970 199884
rect 162964 199822 163022 199882
rect 162964 199820 162970 199822
rect 163814 199820 163820 199884
rect 163884 199858 163916 199884
rect 163972 199858 163977 199914
rect 164187 199914 164253 199919
rect 164187 199884 164192 199914
rect 164248 199884 164253 199914
rect 164371 199914 164437 199919
rect 163884 199853 163977 199858
rect 163884 199822 163928 199853
rect 163884 199820 163890 199822
rect 164182 199820 164188 199884
rect 164252 199882 164258 199884
rect 164252 199822 164310 199882
rect 164371 199858 164376 199914
rect 164432 199858 164437 199914
rect 170443 199914 170509 199919
rect 164371 199853 164437 199858
rect 164555 199880 164621 199885
rect 165107 199884 165173 199885
rect 165102 199882 165108 199884
rect 164252 199820 164258 199822
rect 134379 199819 134445 199820
rect 164374 199749 164434 199853
rect 164555 199824 164560 199880
rect 164616 199824 164621 199880
rect 164555 199819 164621 199824
rect 165016 199822 165108 199882
rect 165102 199820 165108 199822
rect 165172 199820 165178 199884
rect 165291 199882 165357 199885
rect 166022 199882 166028 199884
rect 165291 199880 166028 199882
rect 165291 199824 165296 199880
rect 165352 199824 166028 199880
rect 165291 199822 166028 199824
rect 165107 199819 165173 199820
rect 165291 199819 165357 199822
rect 166022 199820 166028 199822
rect 166092 199820 166098 199884
rect 166763 199880 166829 199885
rect 166763 199824 166768 199880
rect 166824 199824 166829 199880
rect 166763 199819 166829 199824
rect 167407 199882 167473 199885
rect 168235 199884 168301 199885
rect 168046 199882 168052 199884
rect 167407 199880 168052 199882
rect 167407 199824 167412 199880
rect 167468 199824 168052 199880
rect 167407 199822 168052 199824
rect 167407 199819 167473 199822
rect 168046 199820 168052 199822
rect 168116 199820 168122 199884
rect 168230 199820 168236 199884
rect 168300 199882 168306 199884
rect 168787 199882 168853 199885
rect 168300 199822 168392 199882
rect 168606 199880 168853 199882
rect 168606 199824 168792 199880
rect 168848 199824 168853 199880
rect 168606 199822 168853 199824
rect 168300 199820 168306 199822
rect 168235 199819 168301 199820
rect 164558 199749 164618 199819
rect 43437 199746 43503 199749
rect 160686 199746 160692 199748
rect 43437 199744 160692 199746
rect 43437 199688 43442 199744
rect 43498 199688 160692 199744
rect 43437 199686 160692 199688
rect 43437 199683 43503 199686
rect 160686 199684 160692 199686
rect 160756 199684 160762 199748
rect 160878 199686 164250 199746
rect 164374 199744 164483 199749
rect 164374 199688 164422 199744
rect 164478 199688 164483 199744
rect 164374 199686 164483 199688
rect 164558 199744 164667 199749
rect 164558 199688 164606 199744
rect 164662 199688 164667 199744
rect 164558 199686 164667 199688
rect 102777 199610 102843 199613
rect 102777 199608 113190 199610
rect 102777 199552 102782 199608
rect 102838 199552 113190 199608
rect 102777 199550 113190 199552
rect 102777 199547 102843 199550
rect 26877 199474 26943 199477
rect 26877 199472 103530 199474
rect 26877 199416 26882 199472
rect 26938 199416 103530 199472
rect 26877 199414 103530 199416
rect 26877 199411 26943 199414
rect 103470 198930 103530 199414
rect 113130 199066 113190 199550
rect 122230 199548 122236 199612
rect 122300 199610 122306 199612
rect 160878 199610 160938 199686
rect 122300 199550 160938 199610
rect 122300 199548 122306 199550
rect 161054 199548 161060 199612
rect 161124 199610 161130 199612
rect 161289 199610 161355 199613
rect 161124 199608 161355 199610
rect 161124 199552 161294 199608
rect 161350 199552 161355 199608
rect 161124 199550 161355 199552
rect 161124 199548 161130 199550
rect 161289 199547 161355 199550
rect 161422 199548 161428 199612
rect 161492 199610 161498 199612
rect 161657 199610 161723 199613
rect 161492 199608 161723 199610
rect 161492 199552 161662 199608
rect 161718 199552 161723 199608
rect 161492 199550 161723 199552
rect 161492 199548 161498 199550
rect 161657 199547 161723 199550
rect 162158 199548 162164 199612
rect 162228 199610 162234 199612
rect 162485 199610 162551 199613
rect 162228 199608 162551 199610
rect 162228 199552 162490 199608
rect 162546 199552 162551 199608
rect 162228 199550 162551 199552
rect 164190 199610 164250 199686
rect 164417 199683 164483 199686
rect 164601 199683 164667 199686
rect 166390 199684 166396 199748
rect 166460 199746 166466 199748
rect 166766 199746 166826 199819
rect 166460 199686 166826 199746
rect 166460 199684 166466 199686
rect 168373 199610 168439 199613
rect 164190 199608 168439 199610
rect 164190 199552 168378 199608
rect 168434 199552 168439 199608
rect 164190 199550 168439 199552
rect 162228 199548 162234 199550
rect 162485 199547 162551 199550
rect 168373 199547 168439 199550
rect 121862 199412 121868 199476
rect 121932 199474 121938 199476
rect 121932 199414 164066 199474
rect 121932 199412 121938 199414
rect 131757 199338 131823 199341
rect 132493 199338 132559 199341
rect 133137 199340 133203 199341
rect 133505 199340 133571 199341
rect 131757 199336 132559 199338
rect 131757 199280 131762 199336
rect 131818 199280 132498 199336
rect 132554 199280 132559 199336
rect 131757 199278 132559 199280
rect 131757 199275 131823 199278
rect 132493 199275 132559 199278
rect 133086 199276 133092 199340
rect 133156 199338 133203 199340
rect 133454 199338 133460 199340
rect 133156 199336 133248 199338
rect 133198 199280 133248 199336
rect 133156 199278 133248 199280
rect 133414 199278 133460 199338
rect 133524 199336 133571 199340
rect 133566 199280 133571 199336
rect 133156 199276 133203 199278
rect 133454 199276 133460 199278
rect 133524 199276 133571 199280
rect 133822 199276 133828 199340
rect 133892 199338 133898 199340
rect 134149 199338 134215 199341
rect 133892 199336 134215 199338
rect 133892 199280 134154 199336
rect 134210 199280 134215 199336
rect 133892 199278 134215 199280
rect 133892 199276 133898 199278
rect 133137 199275 133203 199276
rect 133505 199275 133571 199276
rect 134149 199275 134215 199278
rect 134558 199276 134564 199340
rect 134628 199338 134634 199340
rect 134977 199338 135043 199341
rect 134628 199336 135043 199338
rect 134628 199280 134982 199336
rect 135038 199280 135043 199336
rect 134628 199278 135043 199280
rect 134628 199276 134634 199278
rect 134977 199275 135043 199278
rect 135846 199276 135852 199340
rect 135916 199338 135922 199340
rect 135989 199338 136055 199341
rect 135916 199336 136055 199338
rect 135916 199280 135994 199336
rect 136050 199280 136055 199336
rect 135916 199278 136055 199280
rect 135916 199276 135922 199278
rect 135989 199275 136055 199278
rect 136398 199276 136404 199340
rect 136468 199338 136474 199340
rect 136541 199338 136607 199341
rect 136468 199336 136607 199338
rect 136468 199280 136546 199336
rect 136602 199280 136607 199336
rect 136468 199278 136607 199280
rect 136468 199276 136474 199278
rect 136541 199275 136607 199278
rect 136725 199338 136791 199341
rect 137369 199340 137435 199341
rect 136950 199338 136956 199340
rect 136725 199336 136956 199338
rect 136725 199280 136730 199336
rect 136786 199280 136956 199336
rect 136725 199278 136956 199280
rect 136725 199275 136791 199278
rect 136950 199276 136956 199278
rect 137020 199276 137026 199340
rect 137318 199276 137324 199340
rect 137388 199338 137435 199340
rect 137829 199338 137895 199341
rect 138105 199338 138171 199341
rect 137388 199336 137480 199338
rect 137430 199280 137480 199336
rect 137388 199278 137480 199280
rect 137829 199336 138171 199338
rect 137829 199280 137834 199336
rect 137890 199280 138110 199336
rect 138166 199280 138171 199336
rect 137829 199278 138171 199280
rect 137388 199276 137435 199278
rect 137369 199275 137435 199276
rect 137829 199275 137895 199278
rect 138105 199275 138171 199278
rect 138238 199276 138244 199340
rect 138308 199338 138314 199340
rect 151261 199338 151327 199341
rect 138308 199336 151327 199338
rect 138308 199280 151266 199336
rect 151322 199280 151327 199336
rect 138308 199278 151327 199280
rect 138308 199276 138314 199278
rect 151261 199275 151327 199278
rect 153009 199338 153075 199341
rect 153142 199338 153148 199340
rect 153009 199336 153148 199338
rect 153009 199280 153014 199336
rect 153070 199280 153148 199336
rect 153009 199278 153148 199280
rect 153009 199275 153075 199278
rect 153142 199276 153148 199278
rect 153212 199276 153218 199340
rect 153377 199338 153443 199341
rect 156965 199338 157031 199341
rect 153377 199336 157031 199338
rect 153377 199280 153382 199336
rect 153438 199280 156970 199336
rect 157026 199280 157031 199336
rect 153377 199278 157031 199280
rect 153377 199275 153443 199278
rect 156965 199275 157031 199278
rect 160553 199338 160619 199341
rect 161289 199340 161355 199341
rect 160870 199338 160876 199340
rect 160553 199336 160876 199338
rect 160553 199280 160558 199336
rect 160614 199280 160876 199336
rect 160553 199278 160876 199280
rect 160553 199275 160619 199278
rect 160870 199276 160876 199278
rect 160940 199276 160946 199340
rect 161238 199276 161244 199340
rect 161308 199338 161355 199340
rect 161308 199336 161400 199338
rect 161350 199280 161400 199336
rect 161308 199278 161400 199280
rect 161308 199276 161355 199278
rect 161606 199276 161612 199340
rect 161676 199338 161682 199340
rect 162117 199338 162183 199341
rect 161676 199336 162183 199338
rect 161676 199280 162122 199336
rect 162178 199280 162183 199336
rect 161676 199278 162183 199280
rect 161676 199276 161682 199278
rect 161289 199275 161355 199276
rect 162117 199275 162183 199278
rect 162485 199340 162551 199341
rect 162945 199340 163011 199341
rect 162485 199336 162532 199340
rect 162596 199338 162602 199340
rect 162894 199338 162900 199340
rect 162485 199280 162490 199336
rect 162485 199276 162532 199280
rect 162596 199278 162642 199338
rect 162854 199278 162900 199338
rect 162964 199336 163011 199340
rect 163006 199280 163011 199336
rect 162596 199276 162602 199278
rect 162894 199276 162900 199278
rect 162964 199276 163011 199280
rect 162485 199275 162551 199276
rect 162945 199275 163011 199276
rect 116577 199202 116643 199205
rect 124949 199202 125015 199205
rect 116577 199200 125015 199202
rect 116577 199144 116582 199200
rect 116638 199144 124954 199200
rect 125010 199144 125015 199200
rect 116577 199142 125015 199144
rect 116577 199139 116643 199142
rect 124949 199139 125015 199142
rect 130929 199202 130995 199205
rect 132033 199202 132099 199205
rect 130929 199200 132099 199202
rect 130929 199144 130934 199200
rect 130990 199144 132038 199200
rect 132094 199144 132099 199200
rect 130929 199142 132099 199144
rect 130929 199139 130995 199142
rect 132033 199139 132099 199142
rect 133270 199140 133276 199204
rect 133340 199202 133346 199204
rect 133505 199202 133571 199205
rect 133340 199200 133571 199202
rect 133340 199144 133510 199200
rect 133566 199144 133571 199200
rect 133340 199142 133571 199144
rect 133340 199140 133346 199142
rect 133505 199139 133571 199142
rect 133781 199202 133847 199205
rect 134374 199202 134380 199204
rect 133781 199200 134380 199202
rect 133781 199144 133786 199200
rect 133842 199144 134380 199200
rect 133781 199142 134380 199144
rect 133781 199139 133847 199142
rect 134374 199140 134380 199142
rect 134444 199140 134450 199204
rect 136766 199140 136772 199204
rect 136836 199202 136842 199204
rect 137277 199202 137343 199205
rect 136836 199200 137343 199202
rect 136836 199144 137282 199200
rect 137338 199144 137343 199200
rect 136836 199142 137343 199144
rect 136836 199140 136842 199142
rect 137277 199139 137343 199142
rect 137829 199202 137895 199205
rect 138054 199202 138060 199204
rect 137829 199200 138060 199202
rect 137829 199144 137834 199200
rect 137890 199144 138060 199200
rect 137829 199142 138060 199144
rect 137829 199139 137895 199142
rect 138054 199140 138060 199142
rect 138124 199140 138130 199204
rect 139342 199140 139348 199204
rect 139412 199202 139418 199204
rect 140313 199202 140379 199205
rect 139412 199200 140379 199202
rect 139412 199144 140318 199200
rect 140374 199144 140379 199200
rect 139412 199142 140379 199144
rect 139412 199140 139418 199142
rect 140313 199139 140379 199142
rect 140497 199202 140563 199205
rect 141182 199202 141188 199204
rect 140497 199200 141188 199202
rect 140497 199144 140502 199200
rect 140558 199144 141188 199200
rect 140497 199142 141188 199144
rect 140497 199139 140563 199142
rect 141182 199140 141188 199142
rect 141252 199140 141258 199204
rect 143942 199140 143948 199204
rect 144012 199202 144018 199204
rect 144361 199202 144427 199205
rect 144012 199200 144427 199202
rect 144012 199144 144366 199200
rect 144422 199144 144427 199200
rect 144012 199142 144427 199144
rect 144012 199140 144018 199142
rect 144361 199139 144427 199142
rect 146385 199202 146451 199205
rect 146886 199202 146892 199204
rect 146385 199200 146892 199202
rect 146385 199144 146390 199200
rect 146446 199144 146892 199200
rect 146385 199142 146892 199144
rect 146385 199139 146451 199142
rect 146886 199140 146892 199142
rect 146956 199140 146962 199204
rect 147070 199140 147076 199204
rect 147140 199202 147146 199204
rect 147397 199202 147463 199205
rect 147140 199200 147463 199202
rect 147140 199144 147402 199200
rect 147458 199144 147463 199200
rect 147140 199142 147463 199144
rect 147140 199140 147146 199142
rect 147397 199139 147463 199142
rect 149462 199140 149468 199204
rect 149532 199202 149538 199204
rect 150157 199202 150223 199205
rect 149532 199200 150223 199202
rect 149532 199144 150162 199200
rect 150218 199144 150223 199200
rect 149532 199142 150223 199144
rect 149532 199140 149538 199142
rect 150157 199139 150223 199142
rect 150341 199202 150407 199205
rect 156965 199202 157031 199205
rect 150341 199200 157031 199202
rect 150341 199144 150346 199200
rect 150402 199144 156970 199200
rect 157026 199144 157031 199200
rect 150341 199142 157031 199144
rect 150341 199139 150407 199142
rect 156965 199139 157031 199142
rect 157793 199202 157859 199205
rect 158110 199202 158116 199204
rect 157793 199200 158116 199202
rect 157793 199144 157798 199200
rect 157854 199144 158116 199200
rect 157793 199142 158116 199144
rect 157793 199139 157859 199142
rect 158110 199140 158116 199142
rect 158180 199140 158186 199204
rect 158294 199140 158300 199204
rect 158364 199202 158370 199204
rect 163773 199202 163839 199205
rect 158364 199200 163839 199202
rect 158364 199144 163778 199200
rect 163834 199144 163839 199200
rect 158364 199142 163839 199144
rect 164006 199202 164066 199414
rect 167494 199412 167500 199476
rect 167564 199474 167570 199476
rect 167729 199474 167795 199477
rect 167564 199472 167795 199474
rect 167564 199416 167734 199472
rect 167790 199416 167795 199472
rect 167564 199414 167795 199416
rect 168606 199474 168666 199822
rect 168787 199819 168853 199822
rect 168966 199820 168972 199884
rect 169036 199882 169042 199884
rect 169431 199882 169497 199885
rect 169707 199884 169773 199885
rect 170443 199884 170448 199914
rect 170504 199884 170509 199914
rect 170719 199914 170785 199919
rect 169702 199882 169708 199884
rect 169036 199880 169497 199882
rect 169036 199824 169436 199880
rect 169492 199824 169497 199880
rect 169036 199822 169497 199824
rect 169616 199822 169708 199882
rect 169036 199820 169042 199822
rect 169431 199819 169497 199822
rect 169702 199820 169708 199822
rect 169772 199820 169778 199884
rect 170438 199820 170444 199884
rect 170508 199882 170514 199884
rect 170508 199822 170566 199882
rect 170719 199858 170724 199914
rect 170780 199858 170785 199914
rect 170719 199853 170785 199858
rect 171363 199914 171429 199919
rect 171363 199858 171368 199914
rect 171424 199882 171429 199914
rect 172743 199916 172809 199919
rect 172743 199914 172944 199916
rect 172278 199882 172284 199884
rect 171424 199858 172284 199882
rect 171363 199853 172284 199858
rect 171366 199822 172284 199853
rect 170508 199820 170514 199822
rect 172278 199820 172284 199822
rect 172348 199820 172354 199884
rect 172743 199858 172748 199914
rect 172804 199882 172944 199914
rect 173203 199914 173269 199919
rect 173203 199884 173208 199914
rect 173264 199884 173269 199914
rect 173939 199914 174005 199919
rect 173014 199882 173020 199884
rect 172804 199858 173020 199882
rect 172743 199856 173020 199858
rect 172743 199853 172809 199856
rect 172884 199822 173020 199856
rect 173014 199820 173020 199822
rect 173084 199820 173090 199884
rect 173198 199820 173204 199884
rect 173268 199882 173274 199884
rect 173268 199822 173326 199882
rect 173939 199858 173944 199914
rect 174000 199858 174005 199914
rect 174123 199914 174189 199919
rect 174123 199884 174128 199914
rect 174184 199884 174189 199914
rect 173939 199853 174005 199858
rect 173268 199820 173274 199822
rect 169707 199819 169773 199820
rect 168741 199746 168807 199749
rect 173617 199748 173683 199749
rect 169150 199746 169156 199748
rect 168741 199744 169156 199746
rect 168741 199688 168746 199744
rect 168802 199688 169156 199744
rect 168741 199686 169156 199688
rect 168741 199683 168807 199686
rect 169150 199684 169156 199686
rect 169220 199684 169226 199748
rect 173566 199746 173572 199748
rect 173526 199686 173572 199746
rect 173636 199744 173683 199748
rect 173678 199688 173683 199744
rect 173566 199684 173572 199686
rect 173636 199684 173683 199688
rect 173617 199683 173683 199684
rect 168741 199610 168807 199613
rect 168925 199610 168991 199613
rect 168741 199608 168991 199610
rect 168741 199552 168746 199608
rect 168802 199552 168930 199608
rect 168986 199552 168991 199608
rect 168741 199550 168991 199552
rect 168741 199547 168807 199550
rect 168925 199547 168991 199550
rect 169845 199610 169911 199613
rect 170990 199610 170996 199612
rect 169845 199608 170996 199610
rect 169845 199552 169850 199608
rect 169906 199552 170996 199608
rect 169845 199550 170996 199552
rect 169845 199547 169911 199550
rect 170990 199548 170996 199550
rect 171060 199548 171066 199612
rect 173525 199610 173591 199613
rect 173750 199610 173756 199612
rect 173525 199608 173756 199610
rect 173525 199552 173530 199608
rect 173586 199552 173756 199608
rect 173525 199550 173756 199552
rect 173525 199547 173591 199550
rect 173750 199548 173756 199550
rect 173820 199548 173826 199612
rect 173942 199610 174002 199853
rect 174118 199820 174124 199884
rect 174188 199882 174194 199884
rect 174188 199822 174246 199882
rect 174188 199820 174194 199822
rect 174077 199746 174143 199749
rect 174632 199746 174692 200094
rect 177062 200092 177068 200094
rect 177132 200092 177138 200156
rect 207054 200154 207060 200156
rect 183510 200094 207060 200154
rect 179321 200018 179387 200021
rect 176150 200016 179387 200018
rect 176150 199960 179326 200016
rect 179382 199960 179387 200016
rect 176150 199958 179387 199960
rect 175043 199914 175109 199919
rect 174767 199882 174833 199885
rect 174767 199880 174876 199882
rect 174767 199824 174772 199880
rect 174828 199824 174876 199880
rect 175043 199858 175048 199914
rect 175104 199858 175109 199914
rect 175043 199853 175109 199858
rect 175319 199882 175385 199885
rect 176150 199882 176210 199958
rect 179321 199955 179387 199958
rect 176791 199884 176857 199885
rect 176786 199882 176792 199884
rect 175319 199880 176210 199882
rect 174767 199819 174876 199824
rect 174077 199744 174692 199746
rect 174077 199688 174082 199744
rect 174138 199688 174692 199744
rect 174077 199686 174692 199688
rect 174816 199748 174876 199819
rect 175046 199749 175106 199853
rect 175319 199824 175324 199880
rect 175380 199824 176210 199880
rect 175319 199822 176210 199824
rect 176700 199822 176792 199882
rect 175319 199819 175385 199822
rect 176786 199820 176792 199822
rect 176856 199820 176862 199884
rect 177067 199882 177133 199885
rect 177246 199882 177252 199884
rect 177067 199880 177252 199882
rect 177067 199824 177072 199880
rect 177128 199824 177252 199880
rect 177067 199822 177252 199824
rect 176791 199819 176857 199820
rect 177067 199819 177133 199822
rect 177246 199820 177252 199822
rect 177316 199820 177322 199884
rect 174816 199686 174860 199748
rect 174077 199683 174143 199686
rect 174854 199684 174860 199686
rect 174924 199684 174930 199748
rect 174997 199744 175106 199749
rect 183510 199746 183570 200094
rect 207054 200092 207060 200094
rect 207124 200092 207130 200156
rect 174997 199688 175002 199744
rect 175058 199688 175106 199744
rect 174997 199686 175106 199688
rect 175966 199686 183570 199746
rect 174997 199683 175063 199686
rect 175966 199610 176026 199686
rect 173942 199550 176026 199610
rect 176101 199612 176167 199613
rect 176101 199608 176148 199612
rect 176212 199610 176218 199612
rect 176101 199552 176106 199608
rect 176101 199548 176148 199552
rect 176212 199550 176258 199610
rect 176212 199548 176218 199550
rect 176326 199548 176332 199612
rect 176396 199610 176402 199612
rect 176837 199610 176903 199613
rect 176396 199608 176903 199610
rect 176396 199552 176842 199608
rect 176898 199552 176903 199608
rect 176396 199550 176903 199552
rect 176396 199548 176402 199550
rect 176101 199547 176167 199548
rect 176837 199547 176903 199550
rect 177062 199548 177068 199612
rect 177132 199610 177138 199612
rect 178125 199610 178191 199613
rect 177132 199608 178191 199610
rect 177132 199552 178130 199608
rect 178186 199552 178191 199608
rect 177132 199550 178191 199552
rect 177132 199548 177138 199550
rect 178125 199547 178191 199550
rect 217225 199610 217291 199613
rect 239397 199610 239463 199613
rect 217225 199608 239463 199610
rect 217225 199552 217230 199608
rect 217286 199552 239402 199608
rect 239458 199552 239463 199608
rect 217225 199550 239463 199552
rect 217225 199547 217291 199550
rect 239397 199547 239463 199550
rect 169293 199474 169359 199477
rect 168606 199472 169359 199474
rect 168606 199416 169298 199472
rect 169354 199416 169359 199472
rect 168606 199414 169359 199416
rect 167564 199412 167570 199414
rect 167729 199411 167795 199414
rect 169293 199411 169359 199414
rect 170029 199474 170095 199477
rect 216673 199474 216739 199477
rect 516133 199474 516199 199477
rect 170029 199472 516199 199474
rect 170029 199416 170034 199472
rect 170090 199416 216678 199472
rect 216734 199416 516138 199472
rect 516194 199416 516199 199472
rect 170029 199414 516199 199416
rect 170029 199411 170095 199414
rect 216673 199411 216739 199414
rect 516133 199411 516199 199414
rect 165613 199338 165679 199341
rect 182817 199338 182883 199341
rect 211102 199338 211108 199340
rect 165613 199336 182883 199338
rect 165613 199280 165618 199336
rect 165674 199280 182822 199336
rect 182878 199280 182883 199336
rect 165613 199278 182883 199280
rect 165613 199275 165679 199278
rect 182817 199275 182883 199278
rect 200070 199278 211108 199338
rect 168833 199202 168899 199205
rect 164006 199200 168899 199202
rect 164006 199144 168838 199200
rect 168894 199144 168899 199200
rect 164006 199142 168899 199144
rect 158364 199140 158370 199142
rect 163773 199139 163839 199142
rect 168833 199139 168899 199142
rect 169334 199140 169340 199204
rect 169404 199202 169410 199204
rect 169661 199202 169727 199205
rect 169404 199200 169727 199202
rect 169404 199144 169666 199200
rect 169722 199144 169727 199200
rect 169404 199142 169727 199144
rect 169404 199140 169410 199142
rect 169661 199139 169727 199142
rect 170806 199140 170812 199204
rect 170876 199202 170882 199204
rect 171593 199202 171659 199205
rect 170876 199200 171659 199202
rect 170876 199144 171598 199200
rect 171654 199144 171659 199200
rect 170876 199142 171659 199144
rect 170876 199140 170882 199142
rect 171593 199139 171659 199142
rect 174905 199202 174971 199205
rect 176837 199202 176903 199205
rect 174905 199200 176903 199202
rect 174905 199144 174910 199200
rect 174966 199144 176842 199200
rect 176898 199144 176903 199200
rect 174905 199142 176903 199144
rect 174905 199139 174971 199142
rect 176837 199139 176903 199142
rect 181805 199202 181871 199205
rect 200070 199202 200130 199278
rect 211102 199276 211108 199278
rect 211172 199338 211178 199340
rect 544377 199338 544443 199341
rect 211172 199336 544443 199338
rect 211172 199280 544382 199336
rect 544438 199280 544443 199336
rect 211172 199278 544443 199280
rect 211172 199276 211178 199278
rect 544377 199275 544443 199278
rect 181805 199200 200130 199202
rect 181805 199144 181810 199200
rect 181866 199144 200130 199200
rect 181805 199142 200130 199144
rect 181805 199139 181871 199142
rect 114134 199066 114140 199068
rect 113130 199006 114140 199066
rect 114134 199004 114140 199006
rect 114204 199066 114210 199068
rect 147489 199066 147555 199069
rect 150157 199068 150223 199069
rect 151721 199068 151787 199069
rect 150157 199066 150204 199068
rect 114204 199064 147555 199066
rect 114204 199008 147494 199064
rect 147550 199008 147555 199064
rect 114204 199006 147555 199008
rect 150112 199064 150204 199066
rect 150112 199008 150162 199064
rect 150112 199006 150204 199008
rect 114204 199004 114210 199006
rect 147489 199003 147555 199006
rect 150157 199004 150204 199006
rect 150268 199004 150274 199068
rect 151670 199066 151676 199068
rect 151630 199006 151676 199066
rect 151740 199064 151787 199068
rect 151782 199008 151787 199064
rect 151670 199004 151676 199006
rect 151740 199004 151787 199008
rect 150157 199003 150223 199004
rect 151721 199003 151787 199004
rect 152273 199066 152339 199069
rect 189809 199066 189875 199069
rect 152273 199064 189875 199066
rect 152273 199008 152278 199064
rect 152334 199008 189814 199064
rect 189870 199008 189875 199064
rect 152273 199006 189875 199008
rect 152273 199003 152339 199006
rect 189809 199003 189875 199006
rect 109534 198930 109540 198932
rect 103470 198870 109540 198930
rect 109534 198868 109540 198870
rect 109604 198930 109610 198932
rect 144729 198930 144795 198933
rect 109604 198928 144795 198930
rect 109604 198872 144734 198928
rect 144790 198872 144795 198928
rect 109604 198870 144795 198872
rect 109604 198868 109610 198870
rect 144729 198867 144795 198870
rect 149278 198868 149284 198932
rect 149348 198930 149354 198932
rect 149789 198930 149855 198933
rect 188286 198930 188292 198932
rect 149348 198928 188292 198930
rect 149348 198872 149794 198928
rect 149850 198872 188292 198928
rect 149348 198870 188292 198872
rect 149348 198868 149354 198870
rect 149789 198867 149855 198870
rect 188286 198868 188292 198870
rect 188356 198868 188362 198932
rect 131849 198794 131915 198797
rect 133413 198794 133479 198797
rect 134333 198794 134399 198797
rect 131849 198792 132786 198794
rect 131849 198736 131854 198792
rect 131910 198736 132786 198792
rect 131849 198734 132786 198736
rect 131849 198731 131915 198734
rect 120257 198658 120323 198661
rect 121269 198658 121335 198661
rect 132125 198658 132191 198661
rect 120257 198656 132191 198658
rect 120257 198600 120262 198656
rect 120318 198600 121274 198656
rect 121330 198600 132130 198656
rect 132186 198600 132191 198656
rect 120257 198598 132191 198600
rect 132726 198658 132786 198734
rect 133413 198792 134399 198794
rect 133413 198736 133418 198792
rect 133474 198736 134338 198792
rect 134394 198736 134399 198792
rect 133413 198734 134399 198736
rect 133413 198731 133479 198734
rect 134333 198731 134399 198734
rect 134793 198794 134859 198797
rect 135069 198794 135135 198797
rect 134793 198792 135135 198794
rect 134793 198736 134798 198792
rect 134854 198736 135074 198792
rect 135130 198736 135135 198792
rect 134793 198734 135135 198736
rect 134793 198731 134859 198734
rect 135069 198731 135135 198734
rect 135621 198794 135687 198797
rect 137645 198794 137711 198797
rect 135621 198792 137711 198794
rect 135621 198736 135626 198792
rect 135682 198736 137650 198792
rect 137706 198736 137711 198792
rect 135621 198734 137711 198736
rect 135621 198731 135687 198734
rect 137645 198731 137711 198734
rect 138606 198732 138612 198796
rect 138676 198794 138682 198796
rect 138749 198794 138815 198797
rect 138676 198792 138815 198794
rect 138676 198736 138754 198792
rect 138810 198736 138815 198792
rect 138676 198734 138815 198736
rect 138676 198732 138682 198734
rect 138749 198731 138815 198734
rect 140814 198732 140820 198796
rect 140884 198794 140890 198796
rect 141693 198794 141759 198797
rect 144361 198796 144427 198797
rect 140884 198792 141759 198794
rect 140884 198736 141698 198792
rect 141754 198736 141759 198792
rect 140884 198734 141759 198736
rect 140884 198732 140890 198734
rect 141693 198731 141759 198734
rect 144310 198732 144316 198796
rect 144380 198794 144427 198796
rect 149513 198794 149579 198797
rect 149973 198796 150039 198797
rect 149830 198794 149836 198796
rect 144380 198792 144472 198794
rect 144422 198736 144472 198792
rect 144380 198734 144472 198736
rect 149513 198792 149836 198794
rect 149513 198736 149518 198792
rect 149574 198736 149836 198792
rect 149513 198734 149836 198736
rect 144380 198732 144427 198734
rect 144361 198731 144427 198732
rect 149513 198731 149579 198734
rect 149830 198732 149836 198734
rect 149900 198732 149906 198796
rect 149973 198792 150020 198796
rect 150084 198794 150090 198796
rect 149973 198736 149978 198792
rect 149973 198732 150020 198736
rect 150084 198734 150130 198794
rect 150084 198732 150090 198734
rect 151118 198732 151124 198796
rect 151188 198794 151194 198796
rect 152273 198794 152339 198797
rect 151188 198792 152339 198794
rect 151188 198736 152278 198792
rect 152334 198736 152339 198792
rect 151188 198734 152339 198736
rect 151188 198732 151194 198734
rect 149973 198731 150039 198732
rect 152273 198731 152339 198734
rect 153101 198794 153167 198797
rect 153326 198794 153332 198796
rect 153101 198792 153332 198794
rect 153101 198736 153106 198792
rect 153162 198736 153332 198792
rect 153101 198734 153332 198736
rect 153101 198731 153167 198734
rect 153326 198732 153332 198734
rect 153396 198732 153402 198796
rect 153745 198794 153811 198797
rect 154246 198794 154252 198796
rect 153745 198792 154252 198794
rect 153745 198736 153750 198792
rect 153806 198736 154252 198792
rect 153745 198734 154252 198736
rect 153745 198731 153811 198734
rect 154246 198732 154252 198734
rect 154316 198732 154322 198796
rect 154430 198732 154436 198796
rect 154500 198794 154506 198796
rect 154849 198794 154915 198797
rect 158897 198796 158963 198797
rect 154500 198792 154915 198794
rect 154500 198736 154854 198792
rect 154910 198736 154915 198792
rect 154500 198734 154915 198736
rect 154500 198732 154506 198734
rect 154849 198731 154915 198734
rect 158846 198732 158852 198796
rect 158916 198794 158963 198796
rect 159081 198794 159147 198797
rect 159214 198794 159220 198796
rect 158916 198792 159008 198794
rect 158958 198736 159008 198792
rect 158916 198734 159008 198736
rect 159081 198792 159220 198794
rect 159081 198736 159086 198792
rect 159142 198736 159220 198792
rect 159081 198734 159220 198736
rect 158916 198732 158963 198734
rect 158897 198731 158963 198732
rect 159081 198731 159147 198734
rect 159214 198732 159220 198734
rect 159284 198732 159290 198796
rect 160686 198732 160692 198796
rect 160756 198794 160762 198796
rect 165470 198794 165476 198796
rect 160756 198734 165476 198794
rect 160756 198732 160762 198734
rect 165470 198732 165476 198734
rect 165540 198794 165546 198796
rect 167821 198794 167887 198797
rect 165540 198792 167887 198794
rect 165540 198736 167826 198792
rect 167882 198736 167887 198792
rect 165540 198734 167887 198736
rect 165540 198732 165546 198734
rect 167821 198731 167887 198734
rect 168649 198794 168715 198797
rect 217041 198794 217107 198797
rect 217225 198794 217291 198797
rect 168649 198792 217291 198794
rect 168649 198736 168654 198792
rect 168710 198736 217046 198792
rect 217102 198736 217230 198792
rect 217286 198736 217291 198792
rect 168649 198734 217291 198736
rect 168649 198731 168715 198734
rect 217041 198731 217107 198734
rect 217225 198731 217291 198734
rect 138381 198658 138447 198661
rect 138790 198658 138796 198660
rect 132726 198598 138030 198658
rect 120257 198595 120323 198598
rect 121269 198595 121335 198598
rect 132125 198595 132191 198598
rect 136173 198524 136239 198525
rect 137001 198524 137067 198525
rect 124070 198460 124076 198524
rect 124140 198522 124146 198524
rect 136173 198522 136220 198524
rect 124140 198462 136052 198522
rect 136128 198520 136220 198522
rect 136128 198464 136178 198520
rect 136128 198462 136220 198464
rect 124140 198460 124146 198462
rect 122046 198324 122052 198388
rect 122116 198386 122122 198388
rect 135529 198386 135595 198389
rect 122116 198384 135595 198386
rect 122116 198328 135534 198384
rect 135590 198328 135595 198384
rect 122116 198326 135595 198328
rect 135992 198386 136052 198462
rect 136173 198460 136220 198462
rect 136284 198460 136290 198524
rect 136950 198460 136956 198524
rect 137020 198522 137067 198524
rect 137020 198520 137112 198522
rect 137062 198464 137112 198520
rect 137020 198462 137112 198464
rect 137020 198460 137067 198462
rect 136173 198459 136239 198460
rect 137001 198459 137067 198460
rect 137185 198386 137251 198389
rect 135992 198384 137251 198386
rect 135992 198328 137190 198384
rect 137246 198328 137251 198384
rect 135992 198326 137251 198328
rect 137970 198386 138030 198598
rect 138381 198656 138796 198658
rect 138381 198600 138386 198656
rect 138442 198600 138796 198656
rect 138381 198598 138796 198600
rect 138381 198595 138447 198598
rect 138790 198596 138796 198598
rect 138860 198596 138866 198660
rect 140998 198596 141004 198660
rect 141068 198658 141074 198660
rect 142613 198658 142679 198661
rect 144269 198660 144335 198661
rect 172421 198660 172487 198661
rect 144269 198658 144316 198660
rect 141068 198656 142679 198658
rect 141068 198600 142618 198656
rect 142674 198600 142679 198656
rect 141068 198598 142679 198600
rect 144188 198656 144316 198658
rect 144380 198658 144386 198660
rect 144188 198600 144274 198656
rect 144188 198598 144316 198600
rect 141068 198596 141074 198598
rect 142613 198595 142679 198598
rect 144269 198596 144316 198598
rect 144380 198598 168390 198658
rect 144380 198596 144386 198598
rect 144269 198595 144335 198596
rect 138606 198460 138612 198524
rect 138676 198522 138682 198524
rect 142245 198522 142311 198525
rect 138676 198520 142311 198522
rect 138676 198464 142250 198520
rect 142306 198464 142311 198520
rect 138676 198462 142311 198464
rect 138676 198460 138682 198462
rect 142245 198459 142311 198462
rect 145097 198522 145163 198525
rect 146150 198522 146156 198524
rect 145097 198520 146156 198522
rect 145097 198464 145102 198520
rect 145158 198464 146156 198520
rect 145097 198462 146156 198464
rect 145097 198459 145163 198462
rect 146150 198460 146156 198462
rect 146220 198460 146226 198524
rect 148869 198522 148935 198525
rect 148869 198520 157350 198522
rect 148869 198464 148874 198520
rect 148930 198464 157350 198520
rect 148869 198462 157350 198464
rect 148869 198459 148935 198462
rect 150566 198386 150572 198388
rect 137970 198326 150572 198386
rect 122116 198324 122122 198326
rect 135529 198323 135595 198326
rect 137185 198323 137251 198326
rect 150566 198324 150572 198326
rect 150636 198324 150642 198388
rect 151486 198324 151492 198388
rect 151556 198386 151562 198388
rect 151721 198386 151787 198389
rect 151556 198384 151787 198386
rect 151556 198328 151726 198384
rect 151782 198328 151787 198384
rect 151556 198326 151787 198328
rect 151556 198324 151562 198326
rect 151721 198323 151787 198326
rect 154798 198324 154804 198388
rect 154868 198386 154874 198388
rect 156873 198386 156939 198389
rect 154868 198384 156939 198386
rect 154868 198328 156878 198384
rect 156934 198328 156939 198384
rect 154868 198326 156939 198328
rect 157290 198386 157350 198462
rect 166574 198460 166580 198524
rect 166644 198522 166650 198524
rect 166717 198522 166783 198525
rect 166644 198520 166783 198522
rect 166644 198464 166722 198520
rect 166778 198464 166783 198520
rect 166644 198462 166783 198464
rect 168330 198522 168390 198598
rect 172421 198656 172468 198660
rect 172532 198658 172538 198660
rect 172789 198658 172855 198661
rect 173525 198658 173591 198661
rect 172421 198600 172426 198656
rect 172421 198596 172468 198600
rect 172532 198598 172578 198658
rect 172789 198656 173591 198658
rect 172789 198600 172794 198656
rect 172850 198600 173530 198656
rect 173586 198600 173591 198656
rect 172789 198598 173591 198600
rect 172532 198596 172538 198598
rect 172421 198595 172487 198596
rect 172789 198595 172855 198598
rect 173525 198595 173591 198598
rect 174077 198660 174143 198661
rect 175549 198660 175615 198661
rect 174077 198656 174124 198660
rect 174188 198658 174194 198660
rect 174077 198600 174082 198656
rect 174077 198596 174124 198600
rect 174188 198598 174234 198658
rect 175549 198656 175596 198660
rect 175660 198658 175666 198660
rect 175549 198600 175554 198656
rect 174188 198596 174194 198598
rect 175549 198596 175596 198600
rect 175660 198598 175706 198658
rect 175660 198596 175666 198598
rect 174077 198595 174143 198596
rect 175549 198595 175615 198596
rect 177665 198522 177731 198525
rect 168330 198520 177731 198522
rect 168330 198464 177670 198520
rect 177726 198464 177731 198520
rect 168330 198462 177731 198464
rect 166644 198460 166650 198462
rect 166717 198459 166783 198462
rect 177665 198459 177731 198462
rect 169753 198386 169819 198389
rect 157290 198384 169819 198386
rect 157290 198328 169758 198384
rect 169814 198328 169819 198384
rect 157290 198326 169819 198328
rect 154868 198324 154874 198326
rect 156873 198323 156939 198326
rect 169753 198323 169819 198326
rect 173198 198324 173204 198388
rect 173268 198386 173274 198388
rect 173268 198326 178050 198386
rect 173268 198324 173274 198326
rect 138289 198250 138355 198253
rect 139158 198250 139164 198252
rect 138289 198248 139164 198250
rect 138289 198192 138294 198248
rect 138350 198192 139164 198248
rect 138289 198190 139164 198192
rect 138289 198187 138355 198190
rect 139158 198188 139164 198190
rect 139228 198188 139234 198252
rect 139894 198188 139900 198252
rect 139964 198250 139970 198252
rect 143901 198250 143967 198253
rect 139964 198248 143967 198250
rect 139964 198192 143906 198248
rect 143962 198192 143967 198248
rect 139964 198190 143967 198192
rect 139964 198188 139970 198190
rect 143901 198187 143967 198190
rect 156229 198250 156295 198253
rect 177990 198250 178050 198326
rect 189993 198250 190059 198253
rect 156229 198248 165538 198250
rect 156229 198192 156234 198248
rect 156290 198192 165538 198248
rect 156229 198190 165538 198192
rect 156229 198187 156295 198190
rect 138606 198114 138612 198116
rect 126286 198054 138612 198114
rect 104750 197916 104756 197980
rect 104820 197978 104826 197980
rect 120257 197978 120323 197981
rect 104820 197976 120323 197978
rect 104820 197920 120262 197976
rect 120318 197920 120323 197976
rect 104820 197918 120323 197920
rect 104820 197916 104826 197918
rect 120257 197915 120323 197918
rect 122833 197842 122899 197845
rect 123477 197842 123543 197845
rect 126286 197842 126346 198054
rect 138606 198052 138612 198054
rect 138676 198052 138682 198116
rect 138749 198114 138815 198117
rect 138974 198114 138980 198116
rect 138749 198112 138980 198114
rect 138749 198056 138754 198112
rect 138810 198056 138980 198112
rect 138749 198054 138980 198056
rect 138749 198051 138815 198054
rect 138974 198052 138980 198054
rect 139044 198052 139050 198116
rect 139894 198052 139900 198116
rect 139964 198114 139970 198116
rect 140221 198114 140287 198117
rect 139964 198112 140287 198114
rect 139964 198056 140226 198112
rect 140282 198056 140287 198112
rect 139964 198054 140287 198056
rect 139964 198052 139970 198054
rect 140221 198051 140287 198054
rect 142705 198114 142771 198117
rect 143022 198114 143028 198116
rect 142705 198112 143028 198114
rect 142705 198056 142710 198112
rect 142766 198056 143028 198112
rect 142705 198054 143028 198056
rect 142705 198051 142771 198054
rect 143022 198052 143028 198054
rect 143092 198052 143098 198116
rect 144545 198114 144611 198117
rect 144862 198114 144868 198116
rect 144545 198112 144868 198114
rect 144545 198056 144550 198112
rect 144606 198056 144868 198112
rect 144545 198054 144868 198056
rect 144545 198051 144611 198054
rect 144862 198052 144868 198054
rect 144932 198052 144938 198116
rect 146109 198114 146175 198117
rect 148542 198114 148548 198116
rect 146109 198112 148548 198114
rect 146109 198056 146114 198112
rect 146170 198056 148548 198112
rect 146109 198054 148548 198056
rect 146109 198051 146175 198054
rect 148542 198052 148548 198054
rect 148612 198052 148618 198116
rect 151169 198114 151235 198117
rect 152406 198114 152412 198116
rect 151169 198112 152412 198114
rect 151169 198056 151174 198112
rect 151230 198056 152412 198112
rect 151169 198054 152412 198056
rect 151169 198051 151235 198054
rect 152406 198052 152412 198054
rect 152476 198052 152482 198116
rect 154614 198052 154620 198116
rect 154684 198114 154690 198116
rect 155953 198114 156019 198117
rect 154684 198112 156019 198114
rect 154684 198056 155958 198112
rect 156014 198056 156019 198112
rect 154684 198054 156019 198056
rect 154684 198052 154690 198054
rect 155953 198051 156019 198054
rect 165061 198114 165127 198117
rect 165286 198114 165292 198116
rect 165061 198112 165292 198114
rect 165061 198056 165066 198112
rect 165122 198056 165292 198112
rect 165061 198054 165292 198056
rect 165061 198051 165127 198054
rect 165286 198052 165292 198054
rect 165356 198052 165362 198116
rect 165478 198114 165538 198190
rect 166950 198190 176210 198250
rect 177990 198248 190059 198250
rect 177990 198192 189998 198248
rect 190054 198192 190059 198248
rect 177990 198190 190059 198192
rect 166206 198114 166212 198116
rect 165478 198054 166212 198114
rect 166206 198052 166212 198054
rect 166276 198052 166282 198116
rect 166950 198114 167010 198190
rect 166766 198054 167010 198114
rect 168189 198116 168255 198117
rect 168189 198112 168236 198116
rect 168300 198114 168306 198116
rect 168189 198056 168194 198112
rect 126421 197978 126487 197981
rect 126789 197978 126855 197981
rect 149646 197978 149652 197980
rect 126421 197976 149652 197978
rect 126421 197920 126426 197976
rect 126482 197920 126794 197976
rect 126850 197920 149652 197976
rect 126421 197918 149652 197920
rect 126421 197915 126487 197918
rect 126789 197915 126855 197918
rect 149646 197916 149652 197918
rect 149716 197916 149722 197980
rect 122833 197840 126346 197842
rect 122833 197784 122838 197840
rect 122894 197784 123482 197840
rect 123538 197784 126346 197840
rect 122833 197782 126346 197784
rect 122833 197779 122899 197782
rect 123477 197779 123543 197782
rect 138606 197780 138612 197844
rect 138676 197842 138682 197844
rect 139117 197842 139183 197845
rect 138676 197840 139183 197842
rect 138676 197784 139122 197840
rect 139178 197784 139183 197840
rect 138676 197782 139183 197784
rect 138676 197780 138682 197782
rect 139117 197779 139183 197782
rect 145281 197842 145347 197845
rect 146518 197842 146524 197844
rect 145281 197840 146524 197842
rect 145281 197784 145286 197840
rect 145342 197784 146524 197840
rect 145281 197782 146524 197784
rect 145281 197779 145347 197782
rect 146518 197780 146524 197782
rect 146588 197780 146594 197844
rect 163957 197842 164023 197845
rect 166766 197842 166826 198054
rect 168189 198052 168236 198056
rect 168300 198054 168346 198114
rect 168300 198052 168306 198054
rect 174486 198052 174492 198116
rect 174556 198114 174562 198116
rect 174813 198114 174879 198117
rect 174556 198112 174879 198114
rect 174556 198056 174818 198112
rect 174874 198056 174879 198112
rect 174556 198054 174879 198056
rect 176150 198114 176210 198190
rect 189993 198187 190059 198190
rect 182265 198114 182331 198117
rect 176150 198112 182331 198114
rect 176150 198056 182270 198112
rect 182326 198056 182331 198112
rect 176150 198054 182331 198056
rect 174556 198052 174562 198054
rect 168189 198051 168255 198052
rect 174813 198051 174879 198054
rect 182265 198051 182331 198054
rect 168189 197978 168255 197981
rect 179413 197978 179479 197981
rect 168189 197976 179479 197978
rect 168189 197920 168194 197976
rect 168250 197920 179418 197976
rect 179474 197920 179479 197976
rect 168189 197918 179479 197920
rect 168189 197915 168255 197918
rect 179413 197915 179479 197918
rect 163957 197840 166826 197842
rect 163957 197784 163962 197840
rect 164018 197784 166826 197840
rect 163957 197782 166826 197784
rect 163957 197779 164023 197782
rect 139526 197706 139532 197708
rect 122790 197646 139532 197706
rect 122465 197434 122531 197437
rect 122790 197434 122850 197646
rect 139526 197644 139532 197646
rect 139596 197644 139602 197708
rect 171409 197706 171475 197709
rect 193213 197706 193279 197709
rect 171409 197704 193279 197706
rect 171409 197648 171414 197704
rect 171470 197648 193218 197704
rect 193274 197648 193279 197704
rect 171409 197646 193279 197648
rect 171409 197643 171475 197646
rect 193213 197643 193279 197646
rect 140221 197570 140287 197573
rect 140630 197570 140636 197572
rect 140221 197568 140636 197570
rect 140221 197512 140226 197568
rect 140282 197512 140636 197568
rect 140221 197510 140636 197512
rect 140221 197507 140287 197510
rect 140630 197508 140636 197510
rect 140700 197508 140706 197572
rect 122465 197432 122850 197434
rect 122465 197376 122470 197432
rect 122526 197376 122850 197432
rect 122465 197374 122850 197376
rect 139577 197434 139643 197437
rect 147857 197436 147923 197437
rect 140262 197434 140268 197436
rect 139577 197432 140268 197434
rect 139577 197376 139582 197432
rect 139638 197376 140268 197432
rect 139577 197374 140268 197376
rect 122465 197371 122531 197374
rect 139577 197371 139643 197374
rect 140262 197372 140268 197374
rect 140332 197372 140338 197436
rect 147806 197372 147812 197436
rect 147876 197434 147923 197436
rect 147876 197432 147968 197434
rect 147918 197376 147968 197432
rect 147876 197374 147968 197376
rect 147876 197372 147923 197374
rect 147857 197371 147923 197372
rect 109033 197298 109099 197301
rect 141969 197298 142035 197301
rect 109033 197296 142035 197298
rect 109033 197240 109038 197296
rect 109094 197240 141974 197296
rect 142030 197240 142035 197296
rect 109033 197238 142035 197240
rect 109033 197235 109099 197238
rect 141969 197235 142035 197238
rect 142521 197298 142587 197301
rect 558361 197298 558427 197301
rect 142521 197296 558427 197298
rect 142521 197240 142526 197296
rect 142582 197240 558366 197296
rect 558422 197240 558427 197296
rect 142521 197238 558427 197240
rect 142521 197235 142587 197238
rect 558361 197235 558427 197238
rect 580165 197298 580231 197301
rect 583520 197298 584960 197388
rect 580165 197296 584960 197298
rect 580165 197240 580170 197296
rect 580226 197240 584960 197296
rect 580165 197238 584960 197240
rect 580165 197235 580231 197238
rect 135069 197162 135135 197165
rect 139209 197162 139275 197165
rect 135069 197160 139275 197162
rect 135069 197104 135074 197160
rect 135130 197104 139214 197160
rect 139270 197104 139275 197160
rect 135069 197102 139275 197104
rect 135069 197099 135135 197102
rect 139209 197099 139275 197102
rect 142470 197100 142476 197164
rect 142540 197162 142546 197164
rect 333973 197162 334039 197165
rect 142540 197160 334039 197162
rect 142540 197104 333978 197160
rect 334034 197104 334039 197160
rect 583520 197148 584960 197238
rect 142540 197102 334039 197104
rect 142540 197100 142546 197102
rect 333973 197099 334039 197102
rect 102869 197026 102935 197029
rect 169937 197026 170003 197029
rect 102869 197024 170003 197026
rect 102869 196968 102874 197024
rect 102930 196968 169942 197024
rect 169998 196968 170003 197024
rect 102869 196966 170003 196968
rect 102869 196963 102935 196966
rect 169937 196963 170003 196966
rect 174445 197026 174511 197029
rect 207013 197026 207079 197029
rect 174445 197024 207079 197026
rect 174445 196968 174450 197024
rect 174506 196968 207018 197024
rect 207074 196968 207079 197024
rect 174445 196966 207079 196968
rect 174445 196963 174511 196966
rect 207013 196963 207079 196966
rect 106917 196890 106983 196893
rect 169569 196890 169635 196893
rect 173617 196892 173683 196893
rect 106917 196888 169635 196890
rect 106917 196832 106922 196888
rect 106978 196832 169574 196888
rect 169630 196832 169635 196888
rect 106917 196830 169635 196832
rect 106917 196827 106983 196830
rect 169569 196827 169635 196830
rect 173566 196828 173572 196892
rect 173636 196890 173683 196892
rect 174261 196892 174327 196893
rect 173636 196888 173728 196890
rect 173678 196832 173728 196888
rect 173636 196830 173728 196832
rect 174261 196888 174308 196892
rect 174372 196890 174378 196892
rect 179321 196890 179387 196893
rect 218237 196890 218303 196893
rect 566549 196890 566615 196893
rect 174261 196832 174266 196888
rect 173636 196828 173683 196830
rect 173617 196827 173683 196828
rect 174261 196828 174308 196832
rect 174372 196830 174418 196890
rect 179321 196888 566615 196890
rect 179321 196832 179326 196888
rect 179382 196832 218242 196888
rect 218298 196832 566554 196888
rect 566610 196832 566615 196888
rect 179321 196830 566615 196832
rect 174372 196828 174378 196830
rect 174261 196827 174327 196828
rect 179321 196827 179387 196830
rect 218237 196827 218303 196830
rect 566549 196827 566615 196830
rect 138565 196754 138631 196757
rect 180701 196754 180767 196757
rect 138565 196752 180767 196754
rect 138565 196696 138570 196752
rect 138626 196696 180706 196752
rect 180762 196696 180767 196752
rect 138565 196694 180767 196696
rect 138565 196691 138631 196694
rect 180701 196691 180767 196694
rect 207013 196754 207079 196757
rect 207197 196754 207263 196757
rect 561121 196754 561187 196757
rect 207013 196752 561187 196754
rect 207013 196696 207018 196752
rect 207074 196696 207202 196752
rect 207258 196696 561126 196752
rect 561182 196696 561187 196752
rect 207013 196694 561187 196696
rect 207013 196691 207079 196694
rect 207197 196691 207263 196694
rect 561121 196691 561187 196694
rect 108798 196556 108804 196620
rect 108868 196618 108874 196620
rect 142470 196618 142476 196620
rect 108868 196558 142476 196618
rect 108868 196556 108874 196558
rect 142470 196556 142476 196558
rect 142540 196556 142546 196620
rect 147806 196556 147812 196620
rect 147876 196618 147882 196620
rect 149053 196618 149119 196621
rect 570597 196618 570663 196621
rect 147876 196616 570663 196618
rect 147876 196560 149058 196616
rect 149114 196560 570602 196616
rect 570658 196560 570663 196616
rect 147876 196558 570663 196560
rect 147876 196556 147882 196558
rect 149053 196555 149119 196558
rect 570597 196555 570663 196558
rect 129641 196482 129707 196485
rect 143073 196482 143139 196485
rect 129641 196480 143139 196482
rect 129641 196424 129646 196480
rect 129702 196424 143078 196480
rect 143134 196424 143139 196480
rect 129641 196422 143139 196424
rect 129641 196419 129707 196422
rect 143073 196419 143139 196422
rect 152733 196484 152799 196485
rect 152733 196480 152780 196484
rect 152844 196482 152850 196484
rect 157885 196482 157951 196485
rect 158294 196482 158300 196484
rect 152733 196424 152738 196480
rect 152733 196420 152780 196424
rect 152844 196422 152890 196482
rect 157885 196480 158300 196482
rect 157885 196424 157890 196480
rect 157946 196424 158300 196480
rect 157885 196422 158300 196424
rect 152844 196420 152850 196422
rect 152733 196419 152799 196420
rect 157885 196419 157951 196422
rect 158294 196420 158300 196422
rect 158364 196420 158370 196484
rect 160502 196420 160508 196484
rect 160572 196482 160578 196484
rect 161289 196482 161355 196485
rect 160572 196480 161355 196482
rect 160572 196424 161294 196480
rect 161350 196424 161355 196480
rect 160572 196422 161355 196424
rect 160572 196420 160578 196422
rect 161289 196419 161355 196422
rect 162853 196482 162919 196485
rect 196014 196482 196020 196484
rect 162853 196480 196020 196482
rect 162853 196424 162858 196480
rect 162914 196424 196020 196480
rect 162853 196422 196020 196424
rect 162853 196419 162919 196422
rect 196014 196420 196020 196422
rect 196084 196420 196090 196484
rect 138473 196348 138539 196349
rect 138422 196284 138428 196348
rect 138492 196346 138539 196348
rect 151997 196346 152063 196349
rect 152958 196346 152964 196348
rect 138492 196344 138584 196346
rect 138534 196288 138584 196344
rect 138492 196286 138584 196288
rect 151997 196344 152964 196346
rect 151997 196288 152002 196344
rect 152058 196288 152964 196344
rect 151997 196286 152964 196288
rect 138492 196284 138539 196286
rect 138473 196283 138539 196284
rect 151997 196283 152063 196286
rect 152958 196284 152964 196286
rect 153028 196284 153034 196348
rect 163814 196284 163820 196348
rect 163884 196346 163890 196348
rect 164049 196346 164115 196349
rect 163884 196344 164115 196346
rect 163884 196288 164054 196344
rect 164110 196288 164115 196344
rect 163884 196286 164115 196288
rect 163884 196284 163890 196286
rect 164049 196283 164115 196286
rect 165797 196346 165863 196349
rect 166758 196346 166764 196348
rect 165797 196344 166764 196346
rect 165797 196288 165802 196344
rect 165858 196288 166764 196344
rect 165797 196286 166764 196288
rect 165797 196283 165863 196286
rect 166758 196284 166764 196286
rect 166828 196284 166834 196348
rect 168833 196346 168899 196349
rect 168966 196346 168972 196348
rect 168833 196344 168972 196346
rect 168833 196288 168838 196344
rect 168894 196288 168972 196344
rect 168833 196286 168972 196288
rect 168833 196283 168899 196286
rect 168966 196284 168972 196286
rect 169036 196284 169042 196348
rect 153653 196210 153719 196213
rect 154430 196210 154436 196212
rect 153653 196208 154436 196210
rect 153653 196152 153658 196208
rect 153714 196152 154436 196208
rect 153653 196150 154436 196152
rect 153653 196147 153719 196150
rect 154430 196148 154436 196150
rect 154500 196148 154506 196212
rect 157057 196210 157123 196213
rect 165153 196212 165219 196213
rect 168097 196212 168163 196213
rect 157190 196210 157196 196212
rect 157057 196208 157196 196210
rect 157057 196152 157062 196208
rect 157118 196152 157196 196208
rect 157057 196150 157196 196152
rect 157057 196147 157123 196150
rect 157190 196148 157196 196150
rect 157260 196148 157266 196212
rect 165102 196148 165108 196212
rect 165172 196210 165219 196212
rect 165172 196208 165264 196210
rect 165214 196152 165264 196208
rect 165172 196150 165264 196152
rect 165172 196148 165219 196150
rect 168046 196148 168052 196212
rect 168116 196210 168163 196212
rect 168116 196208 168208 196210
rect 168158 196152 168208 196208
rect 168116 196150 168208 196152
rect 168116 196148 168163 196150
rect 165153 196147 165219 196148
rect 168097 196147 168163 196148
rect 136817 196074 136883 196077
rect 153469 196076 153535 196077
rect 137318 196074 137324 196076
rect 136817 196072 137324 196074
rect -960 195938 480 196028
rect 136817 196016 136822 196072
rect 136878 196016 137324 196072
rect 136817 196014 137324 196016
rect 136817 196011 136883 196014
rect 137318 196012 137324 196014
rect 137388 196012 137394 196076
rect 153469 196074 153516 196076
rect 153424 196072 153516 196074
rect 153424 196016 153474 196072
rect 153424 196014 153516 196016
rect 153469 196012 153516 196014
rect 153580 196012 153586 196076
rect 157006 196012 157012 196076
rect 157076 196074 157082 196076
rect 157333 196074 157399 196077
rect 157076 196072 157399 196074
rect 157076 196016 157338 196072
rect 157394 196016 157399 196072
rect 157076 196014 157399 196016
rect 157076 196012 157082 196014
rect 153469 196011 153535 196012
rect 157333 196011 157399 196014
rect 158662 196012 158668 196076
rect 158732 196074 158738 196076
rect 158989 196074 159055 196077
rect 158732 196072 159055 196074
rect 158732 196016 158994 196072
rect 159050 196016 159055 196072
rect 158732 196014 159055 196016
rect 158732 196012 158738 196014
rect 158989 196011 159055 196014
rect 159541 196074 159607 196077
rect 160318 196074 160324 196076
rect 159541 196072 160324 196074
rect 159541 196016 159546 196072
rect 159602 196016 160324 196072
rect 159541 196014 160324 196016
rect 159541 196011 159607 196014
rect 160318 196012 160324 196014
rect 160388 196012 160394 196076
rect 161105 196074 161171 196077
rect 161238 196074 161244 196076
rect 161105 196072 161244 196074
rect 161105 196016 161110 196072
rect 161166 196016 161244 196072
rect 161105 196014 161244 196016
rect 161105 196011 161171 196014
rect 161238 196012 161244 196014
rect 161308 196012 161314 196076
rect 163129 196074 163195 196077
rect 163998 196074 164004 196076
rect 163129 196072 164004 196074
rect 163129 196016 163134 196072
rect 163190 196016 164004 196072
rect 163129 196014 164004 196016
rect 163129 196011 163195 196014
rect 163998 196012 164004 196014
rect 164068 196012 164074 196076
rect 164325 196074 164391 196077
rect 168966 196074 168972 196076
rect 164325 196072 168972 196074
rect 164325 196016 164330 196072
rect 164386 196016 168972 196072
rect 164325 196014 168972 196016
rect 164325 196011 164391 196014
rect 168966 196012 168972 196014
rect 169036 196012 169042 196076
rect 176653 196074 176719 196077
rect 177062 196074 177068 196076
rect 176653 196072 177068 196074
rect 176653 196016 176658 196072
rect 176714 196016 177068 196072
rect 176653 196014 177068 196016
rect 176653 196011 176719 196014
rect 177062 196012 177068 196014
rect 177132 196012 177138 196076
rect 3417 195938 3483 195941
rect -960 195936 3483 195938
rect -960 195880 3422 195936
rect 3478 195880 3483 195936
rect -960 195878 3483 195880
rect -960 195788 480 195878
rect 3417 195875 3483 195878
rect 91093 195938 91159 195941
rect 122465 195938 122531 195941
rect 91093 195936 122531 195938
rect 91093 195880 91098 195936
rect 91154 195880 122470 195936
rect 122526 195880 122531 195936
rect 91093 195878 122531 195880
rect 91093 195875 91159 195878
rect 122465 195875 122531 195878
rect 122598 195876 122604 195940
rect 122668 195938 122674 195940
rect 122833 195938 122899 195941
rect 133505 195940 133571 195941
rect 122668 195936 122899 195938
rect 122668 195880 122838 195936
rect 122894 195880 122899 195936
rect 122668 195878 122899 195880
rect 122668 195876 122674 195878
rect 122833 195875 122899 195878
rect 133454 195876 133460 195940
rect 133524 195938 133571 195940
rect 136357 195940 136423 195941
rect 136357 195938 136404 195940
rect 133524 195936 133616 195938
rect 133566 195880 133616 195936
rect 133524 195878 133616 195880
rect 136312 195936 136404 195938
rect 136312 195880 136362 195936
rect 136312 195878 136404 195880
rect 133524 195876 133571 195878
rect 133505 195875 133571 195876
rect 136357 195876 136404 195878
rect 136468 195876 136474 195940
rect 138657 195938 138723 195941
rect 139158 195938 139164 195940
rect 138657 195936 139164 195938
rect 138657 195880 138662 195936
rect 138718 195880 139164 195936
rect 138657 195878 139164 195880
rect 136357 195875 136423 195876
rect 138657 195875 138723 195878
rect 139158 195876 139164 195878
rect 139228 195876 139234 195940
rect 147489 195938 147555 195941
rect 574737 195938 574803 195941
rect 147489 195936 574803 195938
rect 147489 195880 147494 195936
rect 147550 195880 574742 195936
rect 574798 195880 574803 195936
rect 147489 195878 574803 195880
rect 147489 195875 147555 195878
rect 574737 195875 574803 195878
rect 104157 195802 104223 195805
rect 170489 195802 170555 195805
rect 104157 195800 170555 195802
rect 104157 195744 104162 195800
rect 104218 195744 170494 195800
rect 170550 195744 170555 195800
rect 104157 195742 170555 195744
rect 104157 195739 104223 195742
rect 170489 195739 170555 195742
rect 182633 195802 182699 195805
rect 215293 195802 215359 195805
rect 182633 195800 215359 195802
rect 182633 195744 182638 195800
rect 182694 195744 215298 195800
rect 215354 195744 215359 195800
rect 182633 195742 215359 195744
rect 182633 195739 182699 195742
rect 215293 195739 215359 195742
rect 140630 195604 140636 195668
rect 140700 195666 140706 195668
rect 141417 195666 141483 195669
rect 140700 195664 141483 195666
rect 140700 195608 141422 195664
rect 141478 195608 141483 195664
rect 140700 195606 141483 195608
rect 140700 195604 140706 195606
rect 141417 195603 141483 195606
rect 166022 195604 166028 195668
rect 166092 195666 166098 195668
rect 200481 195666 200547 195669
rect 214649 195666 214715 195669
rect 376753 195666 376819 195669
rect 166092 195664 200547 195666
rect 166092 195608 200486 195664
rect 200542 195608 200547 195664
rect 166092 195606 200547 195608
rect 166092 195604 166098 195606
rect 200481 195603 200547 195606
rect 209730 195664 376819 195666
rect 209730 195608 214654 195664
rect 214710 195608 376758 195664
rect 376814 195608 376819 195664
rect 209730 195606 376819 195608
rect 122598 195468 122604 195532
rect 122668 195530 122674 195532
rect 145925 195530 145991 195533
rect 147489 195530 147555 195533
rect 122668 195528 147555 195530
rect 122668 195472 145930 195528
rect 145986 195472 147494 195528
rect 147550 195472 147555 195528
rect 122668 195470 147555 195472
rect 122668 195468 122674 195470
rect 145925 195467 145991 195470
rect 147489 195467 147555 195470
rect 155953 195530 156019 195533
rect 170765 195532 170831 195533
rect 162158 195530 162164 195532
rect 155953 195528 162164 195530
rect 155953 195472 155958 195528
rect 156014 195472 162164 195528
rect 155953 195470 162164 195472
rect 155953 195467 156019 195470
rect 162158 195468 162164 195470
rect 162228 195468 162234 195532
rect 170765 195530 170812 195532
rect 170720 195528 170812 195530
rect 170720 195472 170770 195528
rect 170720 195470 170812 195472
rect 170765 195468 170812 195470
rect 170876 195468 170882 195532
rect 209730 195530 209790 195606
rect 214649 195603 214715 195606
rect 376753 195603 376819 195606
rect 172148 195470 209790 195530
rect 215293 195530 215359 195533
rect 215477 195530 215543 195533
rect 577773 195530 577839 195533
rect 215293 195528 577839 195530
rect 215293 195472 215298 195528
rect 215354 195472 215482 195528
rect 215538 195472 577778 195528
rect 577834 195472 577839 195528
rect 215293 195470 577839 195472
rect 170765 195467 170831 195468
rect 113950 195332 113956 195396
rect 114020 195394 114026 195396
rect 146477 195394 146543 195397
rect 168373 195394 168439 195397
rect 114020 195392 168439 195394
rect 114020 195336 146482 195392
rect 146538 195336 168378 195392
rect 168434 195336 168439 195392
rect 114020 195334 168439 195336
rect 114020 195332 114026 195334
rect 146477 195331 146543 195334
rect 168373 195331 168439 195334
rect 170581 195394 170647 195397
rect 172148 195394 172208 195470
rect 215293 195467 215359 195470
rect 215477 195467 215543 195470
rect 577773 195467 577839 195470
rect 170581 195392 172208 195394
rect 170581 195336 170586 195392
rect 170642 195336 172208 195392
rect 170581 195334 172208 195336
rect 170581 195331 170647 195334
rect 172462 195332 172468 195396
rect 172532 195394 172538 195396
rect 214465 195394 214531 195397
rect 577497 195394 577563 195397
rect 172532 195392 577563 195394
rect 172532 195336 214470 195392
rect 214526 195336 577502 195392
rect 577558 195336 577563 195392
rect 172532 195334 577563 195336
rect 172532 195332 172538 195334
rect 214465 195331 214531 195334
rect 577497 195331 577563 195334
rect 105537 195258 105603 195261
rect 117078 195258 117084 195260
rect 105537 195256 117084 195258
rect 105537 195200 105542 195256
rect 105598 195200 117084 195256
rect 105537 195198 117084 195200
rect 105537 195195 105603 195198
rect 117078 195196 117084 195198
rect 117148 195258 117154 195260
rect 150617 195258 150683 195261
rect 117148 195256 150683 195258
rect 117148 195200 150622 195256
rect 150678 195200 150683 195256
rect 117148 195198 150683 195200
rect 117148 195196 117154 195198
rect 150617 195195 150683 195198
rect 169702 195196 169708 195260
rect 169772 195258 169778 195260
rect 211613 195258 211679 195261
rect 580349 195258 580415 195261
rect 169772 195256 580415 195258
rect 169772 195200 211618 195256
rect 211674 195200 580354 195256
rect 580410 195200 580415 195256
rect 169772 195198 580415 195200
rect 169772 195196 169778 195198
rect 211613 195195 211679 195198
rect 580349 195195 580415 195198
rect 163037 195122 163103 195125
rect 197353 195122 197419 195125
rect 163037 195120 197419 195122
rect 163037 195064 163042 195120
rect 163098 195064 197358 195120
rect 197414 195064 197419 195120
rect 163037 195062 197419 195064
rect 163037 195059 163103 195062
rect 197353 195059 197419 195062
rect 176510 194652 176516 194716
rect 176580 194714 176586 194716
rect 177297 194714 177363 194717
rect 176580 194712 177363 194714
rect 176580 194656 177302 194712
rect 177358 194656 177363 194712
rect 176580 194654 177363 194656
rect 176580 194652 176586 194654
rect 177297 194651 177363 194654
rect 84193 194578 84259 194581
rect 84193 194576 157350 194578
rect 84193 194520 84198 194576
rect 84254 194520 157350 194576
rect 84193 194518 157350 194520
rect 84193 194515 84259 194518
rect 126697 194442 126763 194445
rect 137921 194442 137987 194445
rect 126697 194440 137987 194442
rect 126697 194384 126702 194440
rect 126758 194384 137926 194440
rect 137982 194384 137987 194440
rect 126697 194382 137987 194384
rect 126697 194379 126763 194382
rect 137921 194379 137987 194382
rect 123569 194306 123635 194309
rect 133781 194306 133847 194309
rect 123569 194304 133847 194306
rect 123569 194248 123574 194304
rect 123630 194248 133786 194304
rect 133842 194248 133847 194304
rect 123569 194246 133847 194248
rect 123569 194243 123635 194246
rect 133781 194243 133847 194246
rect 121310 194108 121316 194172
rect 121380 194170 121386 194172
rect 141969 194170 142035 194173
rect 121380 194168 142035 194170
rect 121380 194112 141974 194168
rect 142030 194112 142035 194168
rect 121380 194110 142035 194112
rect 157290 194170 157350 194518
rect 196014 194516 196020 194580
rect 196084 194578 196090 194580
rect 196566 194578 196572 194580
rect 196084 194518 196572 194578
rect 196084 194516 196090 194518
rect 196566 194516 196572 194518
rect 196636 194578 196642 194580
rect 571977 194578 572043 194581
rect 196636 194576 572043 194578
rect 196636 194520 571982 194576
rect 572038 194520 572043 194576
rect 196636 194518 572043 194520
rect 196636 194516 196642 194518
rect 571977 194515 572043 194518
rect 167913 194442 167979 194445
rect 181069 194442 181135 194445
rect 167913 194440 181135 194442
rect 167913 194384 167918 194440
rect 167974 194384 181074 194440
rect 181130 194384 181135 194440
rect 167913 194382 181135 194384
rect 167913 194379 167979 194382
rect 181069 194379 181135 194382
rect 182081 194442 182147 194445
rect 391933 194442 391999 194445
rect 182081 194440 391999 194442
rect 182081 194384 182086 194440
rect 182142 194384 391938 194440
rect 391994 194384 391999 194440
rect 182081 194382 391999 194384
rect 182081 194379 182147 194382
rect 391933 194379 391999 194382
rect 172145 194170 172211 194173
rect 205582 194170 205588 194172
rect 157290 194168 205588 194170
rect 157290 194112 172150 194168
rect 172206 194112 205588 194168
rect 157290 194110 205588 194112
rect 121380 194108 121386 194110
rect 141969 194107 142035 194110
rect 172145 194107 172211 194110
rect 205582 194108 205588 194110
rect 205652 194108 205658 194172
rect 121126 193972 121132 194036
rect 121196 194034 121202 194036
rect 128537 194034 128603 194037
rect 135253 194034 135319 194037
rect 175917 194034 175983 194037
rect 121196 194032 128603 194034
rect 121196 193976 128542 194032
rect 128598 193976 128603 194032
rect 121196 193974 128603 193976
rect 121196 193972 121202 193974
rect 128537 193971 128603 193974
rect 133830 194032 175983 194034
rect 133830 193976 135258 194032
rect 135314 193976 175922 194032
rect 175978 193976 175983 194032
rect 133830 193974 175983 193976
rect 97758 193836 97764 193900
rect 97828 193898 97834 193900
rect 133830 193898 133890 193974
rect 135253 193971 135319 193974
rect 175917 193971 175983 193974
rect 97828 193838 133890 193898
rect 97828 193836 97834 193838
rect 134374 193836 134380 193900
rect 134444 193898 134450 193900
rect 134793 193898 134859 193901
rect 134444 193896 134859 193898
rect 134444 193840 134798 193896
rect 134854 193840 134859 193896
rect 134444 193838 134859 193840
rect 134444 193836 134450 193838
rect 134793 193835 134859 193838
rect 161974 193836 161980 193900
rect 162044 193898 162050 193900
rect 217133 193898 217199 193901
rect 581729 193898 581795 193901
rect 162044 193896 581795 193898
rect 162044 193840 217138 193896
rect 217194 193840 581734 193896
rect 581790 193840 581795 193896
rect 162044 193838 581795 193840
rect 162044 193836 162050 193838
rect 217133 193835 217199 193838
rect 581729 193835 581795 193838
rect 170857 193354 170923 193357
rect 187734 193354 187740 193356
rect 170857 193352 187740 193354
rect 170857 193296 170862 193352
rect 170918 193296 187740 193352
rect 170857 193294 187740 193296
rect 170857 193291 170923 193294
rect 187734 193292 187740 193294
rect 187804 193292 187810 193356
rect 117313 193218 117379 193221
rect 162485 193218 162551 193221
rect 117313 193216 162551 193218
rect 117313 193160 117318 193216
rect 117374 193160 162490 193216
rect 162546 193160 162551 193216
rect 117313 193158 162551 193160
rect 117313 193155 117379 193158
rect 162485 193155 162551 193158
rect 579613 193218 579679 193221
rect 583520 193218 584960 193308
rect 579613 193216 584960 193218
rect 579613 193160 579618 193216
rect 579674 193160 584960 193216
rect 579613 193158 584960 193160
rect 579613 193155 579679 193158
rect 135989 193082 136055 193085
rect 556889 193082 556955 193085
rect 135989 193080 556955 193082
rect 135989 193024 135994 193080
rect 136050 193024 556894 193080
rect 556950 193024 556955 193080
rect 583520 193068 584960 193158
rect 135989 193022 556955 193024
rect 135989 193019 136055 193022
rect 556889 193019 556955 193022
rect 89069 192946 89135 192949
rect 169937 192946 170003 192949
rect 89069 192944 170003 192946
rect 89069 192888 89074 192944
rect 89130 192888 169942 192944
rect 169998 192888 170003 192944
rect 89069 192886 170003 192888
rect 89069 192883 89135 192886
rect 169937 192883 170003 192886
rect 136766 192748 136772 192812
rect 136836 192810 136842 192812
rect 136909 192810 136975 192813
rect 136836 192808 136975 192810
rect 136836 192752 136914 192808
rect 136970 192752 136975 192808
rect 136836 192750 136975 192752
rect 136836 192748 136842 192750
rect 136909 192747 136975 192750
rect 175590 192748 175596 192812
rect 175660 192810 175666 192812
rect 215293 192810 215359 192813
rect 342253 192810 342319 192813
rect 175660 192808 342319 192810
rect 175660 192752 215298 192808
rect 215354 192752 342258 192808
rect 342314 192752 342319 192808
rect 175660 192750 342319 192752
rect 175660 192748 175666 192750
rect 215293 192747 215359 192750
rect 342253 192747 342319 192750
rect -960 192538 480 192628
rect 120574 192612 120580 192676
rect 120644 192674 120650 192676
rect 147070 192674 147076 192676
rect 120644 192614 147076 192674
rect 120644 192612 120650 192614
rect 147070 192612 147076 192614
rect 147140 192674 147146 192676
rect 179137 192674 179203 192677
rect 215569 192674 215635 192677
rect 574921 192674 574987 192677
rect 147140 192614 157350 192674
rect 147140 192612 147146 192614
rect 3417 192538 3483 192541
rect -960 192536 3483 192538
rect -960 192480 3422 192536
rect 3478 192480 3483 192536
rect -960 192478 3483 192480
rect -960 192388 480 192478
rect 3417 192475 3483 192478
rect 104341 192538 104407 192541
rect 118049 192538 118115 192541
rect 147990 192538 147996 192540
rect 104341 192536 147996 192538
rect 104341 192480 104346 192536
rect 104402 192480 118054 192536
rect 118110 192480 147996 192536
rect 104341 192478 147996 192480
rect 104341 192475 104407 192478
rect 118049 192475 118115 192478
rect 147990 192476 147996 192478
rect 148060 192476 148066 192540
rect 157290 192402 157350 192614
rect 179137 192672 574987 192674
rect 179137 192616 179142 192672
rect 179198 192616 215574 192672
rect 215630 192616 574926 192672
rect 574982 192616 574987 192672
rect 179137 192614 574987 192616
rect 179137 192611 179203 192614
rect 215569 192611 215635 192614
rect 574921 192611 574987 192614
rect 173801 192538 173867 192541
rect 200982 192538 200988 192540
rect 173801 192536 200988 192538
rect 173801 192480 173806 192536
rect 173862 192480 200988 192536
rect 173801 192478 200988 192480
rect 173801 192475 173867 192478
rect 200982 192476 200988 192478
rect 201052 192538 201058 192540
rect 580533 192538 580599 192541
rect 201052 192536 580599 192538
rect 201052 192480 580538 192536
rect 580594 192480 580599 192536
rect 201052 192478 580599 192480
rect 201052 192476 201058 192478
rect 580533 192475 580599 192478
rect 576209 192402 576275 192405
rect 157290 192400 576275 192402
rect 157290 192344 576214 192400
rect 576270 192344 576275 192400
rect 157290 192342 576275 192344
rect 576209 192339 576275 192342
rect 148317 192130 148383 192133
rect 148910 192130 148916 192132
rect 148317 192128 148916 192130
rect 148317 192072 148322 192128
rect 148378 192072 148916 192128
rect 148317 192070 148916 192072
rect 148317 192067 148383 192070
rect 148910 192068 148916 192070
rect 148980 192130 148986 192132
rect 150341 192130 150407 192133
rect 148980 192128 150407 192130
rect 148980 192072 150346 192128
rect 150402 192072 150407 192128
rect 148980 192070 150407 192072
rect 148980 192068 148986 192070
rect 150341 192067 150407 192070
rect 93117 191722 93183 191725
rect 170765 191722 170831 191725
rect 93117 191720 170831 191722
rect 93117 191664 93122 191720
rect 93178 191664 170770 191720
rect 170826 191664 170831 191720
rect 93117 191662 170831 191664
rect 93117 191659 93183 191662
rect 170765 191659 170831 191662
rect 198774 191660 198780 191724
rect 198844 191722 198850 191724
rect 231853 191722 231919 191725
rect 198844 191720 231919 191722
rect 198844 191664 231858 191720
rect 231914 191664 231919 191720
rect 198844 191662 231919 191664
rect 198844 191660 198850 191662
rect 231853 191659 231919 191662
rect 95734 191524 95740 191588
rect 95804 191586 95810 191588
rect 95804 191526 138030 191586
rect 95804 191524 95810 191526
rect 137970 191450 138030 191526
rect 174302 191524 174308 191588
rect 174372 191586 174378 191588
rect 174372 191526 219450 191586
rect 174372 191524 174378 191526
rect 151854 191450 151860 191452
rect 137970 191390 151860 191450
rect 151854 191388 151860 191390
rect 151924 191450 151930 191452
rect 201534 191450 201540 191452
rect 151924 191390 201540 191450
rect 151924 191388 151930 191390
rect 201534 191388 201540 191390
rect 201604 191388 201610 191452
rect 219390 191450 219450 191526
rect 219617 191450 219683 191453
rect 377397 191450 377463 191453
rect 219390 191448 377463 191450
rect 219390 191392 219622 191448
rect 219678 191392 377402 191448
rect 377458 191392 377463 191448
rect 219390 191390 377463 191392
rect 219617 191387 219683 191390
rect 377397 191387 377463 191390
rect 98637 191314 98703 191317
rect 117262 191314 117268 191316
rect 98637 191312 117268 191314
rect 98637 191256 98642 191312
rect 98698 191256 117268 191312
rect 98637 191254 117268 191256
rect 98637 191251 98703 191254
rect 117262 191252 117268 191254
rect 117332 191252 117338 191316
rect 164182 191252 164188 191316
rect 164252 191314 164258 191316
rect 197486 191314 197492 191316
rect 164252 191254 197492 191314
rect 164252 191252 164258 191254
rect 197486 191252 197492 191254
rect 197556 191314 197562 191316
rect 494053 191314 494119 191317
rect 197556 191312 494119 191314
rect 197556 191256 494058 191312
rect 494114 191256 494119 191312
rect 197556 191254 494119 191256
rect 197556 191252 197562 191254
rect 494053 191251 494119 191254
rect 80789 191178 80855 191181
rect 104566 191178 104572 191180
rect 80789 191176 104572 191178
rect 80789 191120 80794 191176
rect 80850 191120 104572 191176
rect 80789 191118 104572 191120
rect 80789 191115 80855 191118
rect 104566 191116 104572 191118
rect 104636 191178 104642 191180
rect 138841 191178 138907 191181
rect 104636 191176 138907 191178
rect 104636 191120 138846 191176
rect 138902 191120 138907 191176
rect 104636 191118 138907 191120
rect 104636 191116 104642 191118
rect 138841 191115 138907 191118
rect 158662 191116 158668 191180
rect 158732 191178 158738 191180
rect 193254 191178 193260 191180
rect 158732 191118 193260 191178
rect 158732 191116 158738 191118
rect 193254 191116 193260 191118
rect 193324 191178 193330 191180
rect 576301 191178 576367 191181
rect 193324 191176 576367 191178
rect 193324 191120 576306 191176
rect 576362 191120 576367 191176
rect 193324 191118 576367 191120
rect 193324 191116 193330 191118
rect 576301 191115 576367 191118
rect 93301 191042 93367 191045
rect 158621 191042 158687 191045
rect 159541 191042 159607 191045
rect 93301 191040 159607 191042
rect 93301 190984 93306 191040
rect 93362 190984 158626 191040
rect 158682 190984 159546 191040
rect 159602 190984 159607 191040
rect 93301 190982 159607 190984
rect 93301 190979 93367 190982
rect 158621 190979 158687 190982
rect 159541 190979 159607 190982
rect 161381 191042 161447 191045
rect 194542 191042 194548 191044
rect 161381 191040 194548 191042
rect 161381 190984 161386 191040
rect 161442 190984 194548 191040
rect 161381 190982 194548 190984
rect 161381 190979 161447 190982
rect 194542 190980 194548 190982
rect 194612 191042 194618 191044
rect 578877 191042 578943 191045
rect 194612 191040 578943 191042
rect 194612 190984 578882 191040
rect 578938 190984 578943 191040
rect 194612 190982 578943 190984
rect 194612 190980 194618 190982
rect 578877 190979 578943 190982
rect 164233 190906 164299 190909
rect 197077 190906 197143 190909
rect 197353 190908 197419 190909
rect 197302 190906 197308 190908
rect 164233 190904 197143 190906
rect 164233 190848 164238 190904
rect 164294 190848 197082 190904
rect 197138 190848 197143 190904
rect 164233 190846 197143 190848
rect 197262 190846 197308 190906
rect 197372 190904 197419 190908
rect 201769 190906 201835 190909
rect 220813 190906 220879 190909
rect 197414 190848 197419 190904
rect 164233 190843 164299 190846
rect 197077 190843 197143 190846
rect 197302 190844 197308 190846
rect 197372 190844 197419 190848
rect 197353 190843 197419 190844
rect 200070 190904 220879 190906
rect 200070 190848 201774 190904
rect 201830 190848 220818 190904
rect 220874 190848 220879 190904
rect 200070 190846 220879 190848
rect 134517 190772 134583 190773
rect 134517 190770 134564 190772
rect 134472 190768 134564 190770
rect 134472 190712 134522 190768
rect 134472 190710 134564 190712
rect 134517 190708 134564 190710
rect 134628 190708 134634 190772
rect 168230 190708 168236 190772
rect 168300 190770 168306 190772
rect 200070 190770 200130 190846
rect 201769 190843 201835 190846
rect 220813 190843 220879 190846
rect 168300 190710 200130 190770
rect 168300 190708 168306 190710
rect 134517 190707 134583 190708
rect 197077 190634 197143 190637
rect 198774 190634 198780 190636
rect 197077 190632 198780 190634
rect 197077 190576 197082 190632
rect 197138 190576 198780 190632
rect 197077 190574 198780 190576
rect 197077 190571 197143 190574
rect 198774 190572 198780 190574
rect 198844 190572 198850 190636
rect 122465 190498 122531 190501
rect 122782 190498 122788 190500
rect 122465 190496 122788 190498
rect 122465 190440 122470 190496
rect 122526 190440 122788 190496
rect 122465 190438 122788 190440
rect 122465 190435 122531 190438
rect 122782 190436 122788 190438
rect 122852 190436 122858 190500
rect 148225 190498 148291 190501
rect 148358 190498 148364 190500
rect 148225 190496 148364 190498
rect 148225 190440 148230 190496
rect 148286 190440 148364 190496
rect 148225 190438 148364 190440
rect 148225 190435 148291 190438
rect 148358 190436 148364 190438
rect 148428 190436 148434 190500
rect 60733 190362 60799 190365
rect 154614 190362 154620 190364
rect 60733 190360 154620 190362
rect 60733 190304 60738 190360
rect 60794 190304 154620 190360
rect 60733 190302 154620 190304
rect 60733 190299 60799 190302
rect 154614 190300 154620 190302
rect 154684 190362 154690 190364
rect 155401 190362 155467 190365
rect 154684 190360 155467 190362
rect 154684 190304 155406 190360
rect 155462 190304 155467 190360
rect 154684 190302 155467 190304
rect 154684 190300 154690 190302
rect 155401 190299 155467 190302
rect 157190 190300 157196 190364
rect 157260 190362 157266 190364
rect 215661 190362 215727 190365
rect 260097 190362 260163 190365
rect 157260 190360 260163 190362
rect 157260 190304 215666 190360
rect 215722 190304 260102 190360
rect 260158 190304 260163 190360
rect 157260 190302 260163 190304
rect 157260 190300 157266 190302
rect 215661 190299 215727 190302
rect 260097 190299 260163 190302
rect 110413 190226 110479 190229
rect 111558 190226 111564 190228
rect 110413 190224 111564 190226
rect 110413 190168 110418 190224
rect 110474 190168 111564 190224
rect 110413 190166 111564 190168
rect 110413 190163 110479 190166
rect 111558 190164 111564 190166
rect 111628 190226 111634 190228
rect 139485 190226 139551 190229
rect 111628 190224 139551 190226
rect 111628 190168 139490 190224
rect 139546 190168 139551 190224
rect 111628 190166 139551 190168
rect 111628 190164 111634 190166
rect 139485 190163 139551 190166
rect 139894 190164 139900 190228
rect 139964 190226 139970 190228
rect 140129 190226 140195 190229
rect 139964 190224 140195 190226
rect 139964 190168 140134 190224
rect 140190 190168 140195 190224
rect 139964 190166 140195 190168
rect 139964 190164 139970 190166
rect 140129 190163 140195 190166
rect 166206 190164 166212 190228
rect 166276 190226 166282 190228
rect 190494 190226 190500 190228
rect 166276 190166 190500 190226
rect 166276 190164 166282 190166
rect 190494 190164 190500 190166
rect 190564 190226 190570 190228
rect 266353 190226 266419 190229
rect 190564 190224 266419 190226
rect 190564 190168 266358 190224
rect 266414 190168 266419 190224
rect 190564 190166 266419 190168
rect 190564 190164 190570 190166
rect 266353 190163 266419 190166
rect 117262 190028 117268 190092
rect 117332 190090 117338 190092
rect 149605 190090 149671 190093
rect 117332 190088 149671 190090
rect 117332 190032 149610 190088
rect 149666 190032 149671 190088
rect 117332 190030 149671 190032
rect 117332 190028 117338 190030
rect 149605 190027 149671 190030
rect 158294 190028 158300 190092
rect 158364 190090 158370 190092
rect 183277 190090 183343 190093
rect 431217 190090 431283 190093
rect 158364 190088 431283 190090
rect 158364 190032 183282 190088
rect 183338 190032 431222 190088
rect 431278 190032 431283 190088
rect 158364 190030 431283 190032
rect 158364 190028 158370 190030
rect 183277 190027 183343 190030
rect 431217 190027 431283 190030
rect 112437 189954 112503 189957
rect 112989 189954 113055 189957
rect 143574 189954 143580 189956
rect 112437 189952 143580 189954
rect 112437 189896 112442 189952
rect 112498 189896 112994 189952
rect 113050 189896 143580 189952
rect 112437 189894 143580 189896
rect 112437 189891 112503 189894
rect 112989 189891 113055 189894
rect 143574 189892 143580 189894
rect 143644 189892 143650 189956
rect 174854 189892 174860 189956
rect 174924 189954 174930 189956
rect 207606 189954 207612 189956
rect 174924 189894 207612 189954
rect 174924 189892 174930 189894
rect 207606 189892 207612 189894
rect 207676 189954 207682 189956
rect 561673 189954 561739 189957
rect 207676 189952 561739 189954
rect 207676 189896 561678 189952
rect 561734 189896 561739 189952
rect 207676 189894 561739 189896
rect 207676 189892 207682 189894
rect 561673 189891 561739 189894
rect 107326 189756 107332 189820
rect 107396 189818 107402 189820
rect 138565 189818 138631 189821
rect 107396 189816 138631 189818
rect 107396 189760 138570 189816
rect 138626 189760 138631 189816
rect 107396 189758 138631 189760
rect 107396 189756 107402 189758
rect 138565 189755 138631 189758
rect 139485 189818 139551 189821
rect 144453 189818 144519 189821
rect 139485 189816 144519 189818
rect 139485 189760 139490 189816
rect 139546 189760 144458 189816
rect 144514 189760 144519 189816
rect 139485 189758 144519 189760
rect 139485 189755 139551 189758
rect 144453 189755 144519 189758
rect 160737 189818 160803 189821
rect 192150 189818 192156 189820
rect 160737 189816 192156 189818
rect 160737 189760 160742 189816
rect 160798 189760 192156 189816
rect 160737 189758 192156 189760
rect 160737 189755 160803 189758
rect 192150 189756 192156 189758
rect 192220 189756 192226 189820
rect 205766 189756 205772 189820
rect 205836 189818 205842 189820
rect 577865 189818 577931 189821
rect 205836 189816 577931 189818
rect 205836 189760 577870 189816
rect 577926 189760 577931 189816
rect 205836 189758 577931 189760
rect 205836 189756 205842 189758
rect 577865 189755 577931 189758
rect 108614 189620 108620 189684
rect 108684 189682 108690 189684
rect 142613 189682 142679 189685
rect 108684 189680 142679 189682
rect 108684 189624 142618 189680
rect 142674 189624 142679 189680
rect 108684 189622 142679 189624
rect 108684 189620 108690 189622
rect 142613 189619 142679 189622
rect 157006 189620 157012 189684
rect 157076 189682 157082 189684
rect 181989 189682 182055 189685
rect 574829 189682 574895 189685
rect 157076 189680 574895 189682
rect 157076 189624 181994 189680
rect 182050 189624 574834 189680
rect 574890 189624 574895 189680
rect 157076 189622 574895 189624
rect 157076 189620 157082 189622
rect 181989 189619 182055 189622
rect 574829 189619 574895 189622
rect 122741 189546 122807 189549
rect 122966 189546 122972 189548
rect 122696 189544 122972 189546
rect 122696 189488 122746 189544
rect 122802 189488 122972 189544
rect 122696 189486 122972 189488
rect 122741 189483 122807 189486
rect 122966 189484 122972 189486
rect 123036 189484 123042 189548
rect 172278 189484 172284 189548
rect 172348 189546 172354 189548
rect 215385 189546 215451 189549
rect 172348 189544 215451 189546
rect 172348 189488 215390 189544
rect 215446 189488 215451 189544
rect 172348 189486 215451 189488
rect 172348 189484 172354 189486
rect 215385 189483 215451 189486
rect 167453 189140 167519 189141
rect 116894 189076 116900 189140
rect 116964 189138 116970 189140
rect 117262 189138 117268 189140
rect 116964 189078 117268 189138
rect 116964 189076 116970 189078
rect 117262 189076 117268 189078
rect 117332 189076 117338 189140
rect 167453 189136 167500 189140
rect 167564 189138 167570 189140
rect 579981 189138 580047 189141
rect 583520 189138 584960 189228
rect 167453 189080 167458 189136
rect 167453 189076 167500 189080
rect 167564 189078 167610 189138
rect 579981 189136 584960 189138
rect 579981 189080 579986 189136
rect 580042 189080 584960 189136
rect 579981 189078 584960 189080
rect 167564 189076 167570 189078
rect 167453 189075 167519 189076
rect 579981 189075 580047 189078
rect 129089 189002 129155 189005
rect 129641 189002 129707 189005
rect 138933 189004 138999 189005
rect 138933 189002 138980 189004
rect 129089 189000 138030 189002
rect 129089 188944 129094 189000
rect 129150 188944 129646 189000
rect 129702 188944 138030 189000
rect 129089 188942 138030 188944
rect 138888 189000 138980 189002
rect 138888 188944 138938 189000
rect 138888 188942 138980 188944
rect 129089 188939 129155 188942
rect 129641 188939 129707 188942
rect 137970 188866 138030 188942
rect 138933 188940 138980 188942
rect 139044 188940 139050 189004
rect 151721 189002 151787 189005
rect 563789 189002 563855 189005
rect 151721 189000 563855 189002
rect 151721 188944 151726 189000
rect 151782 188944 563794 189000
rect 563850 188944 563855 189000
rect 583520 188988 584960 189078
rect 151721 188942 563855 188944
rect 138933 188939 138999 188940
rect 151721 188939 151787 188942
rect 563789 188939 563855 188942
rect 524413 188866 524479 188869
rect 137970 188864 524479 188866
rect 137970 188808 524418 188864
rect 524474 188808 524479 188864
rect 137970 188806 524479 188808
rect 524413 188803 524479 188806
rect 138933 188730 138999 188733
rect 455413 188730 455479 188733
rect 138933 188728 455479 188730
rect 138933 188672 138938 188728
rect 138994 188672 455418 188728
rect 455474 188672 455479 188728
rect 138933 188670 455479 188672
rect 138933 188667 138999 188670
rect 455413 188667 455479 188670
rect 171685 188594 171751 188597
rect 205766 188594 205772 188596
rect 171685 188592 205772 188594
rect -960 188458 480 188548
rect 171685 188536 171690 188592
rect 171746 188536 205772 188592
rect 171685 188534 205772 188536
rect 171685 188531 171751 188534
rect 205766 188532 205772 188534
rect 205836 188532 205842 188596
rect 3233 188458 3299 188461
rect -960 188456 3299 188458
rect -960 188400 3238 188456
rect 3294 188400 3299 188456
rect -960 188398 3299 188400
rect -960 188308 480 188398
rect 3233 188395 3299 188398
rect 122230 188396 122236 188460
rect 122300 188458 122306 188460
rect 151721 188458 151787 188461
rect 122300 188456 151787 188458
rect 122300 188400 151726 188456
rect 151782 188400 151787 188456
rect 122300 188398 151787 188400
rect 122300 188396 122306 188398
rect 151721 188395 151787 188398
rect 154481 188458 154547 188461
rect 182766 188458 182772 188460
rect 154481 188456 182772 188458
rect 154481 188400 154486 188456
rect 154542 188400 182772 188456
rect 154481 188398 182772 188400
rect 154481 188395 154547 188398
rect 182766 188396 182772 188398
rect 182836 188396 182842 188460
rect 149830 188260 149836 188324
rect 149900 188322 149906 188324
rect 189206 188322 189212 188324
rect 149900 188262 189212 188322
rect 149900 188260 149906 188262
rect 189206 188260 189212 188262
rect 189276 188322 189282 188324
rect 580993 188322 581059 188325
rect 189276 188320 581059 188322
rect 189276 188264 580998 188320
rect 581054 188264 581059 188320
rect 189276 188262 581059 188264
rect 189276 188260 189282 188262
rect 580993 188259 581059 188262
rect 170213 187780 170279 187781
rect 170213 187776 170260 187780
rect 170324 187778 170330 187780
rect 170213 187720 170218 187776
rect 170213 187716 170260 187720
rect 170324 187718 170370 187778
rect 170324 187716 170330 187718
rect 170213 187715 170279 187716
rect 148961 187642 149027 187645
rect 580441 187642 580507 187645
rect 148961 187640 580507 187642
rect 148961 187584 148966 187640
rect 149022 187584 580446 187640
rect 580502 187584 580507 187640
rect 148961 187582 580507 187584
rect 148961 187579 149027 187582
rect 580441 187579 580507 187582
rect 144913 187506 144979 187509
rect 145649 187506 145715 187509
rect 566641 187506 566707 187509
rect 144913 187504 566707 187506
rect 144913 187448 144918 187504
rect 144974 187448 145654 187504
rect 145710 187448 566646 187504
rect 566702 187448 566707 187504
rect 144913 187446 566707 187448
rect 144913 187443 144979 187446
rect 145649 187443 145715 187446
rect 566641 187443 566707 187446
rect 199326 187308 199332 187372
rect 199396 187370 199402 187372
rect 200481 187370 200547 187373
rect 489913 187370 489979 187373
rect 199396 187368 489979 187370
rect 199396 187312 200486 187368
rect 200542 187312 489918 187368
rect 489974 187312 489979 187368
rect 199396 187310 489979 187312
rect 199396 187308 199402 187310
rect 200481 187307 200547 187310
rect 489913 187307 489979 187310
rect 113766 187036 113772 187100
rect 113836 187098 113842 187100
rect 145097 187098 145163 187101
rect 113836 187096 145163 187098
rect 113836 187040 145102 187096
rect 145158 187040 145163 187096
rect 113836 187038 145163 187040
rect 113836 187036 113842 187038
rect 145097 187035 145163 187038
rect 108430 186900 108436 186964
rect 108500 186962 108506 186964
rect 143073 186962 143139 186965
rect 108500 186960 143139 186962
rect 108500 186904 143078 186960
rect 143134 186904 143139 186960
rect 108500 186902 143139 186904
rect 108500 186900 108506 186902
rect 143073 186899 143139 186902
rect 160553 186962 160619 186965
rect 180701 186962 180767 186965
rect 452653 186962 452719 186965
rect 160553 186960 452719 186962
rect 160553 186904 160558 186960
rect 160614 186904 180706 186960
rect 180762 186904 452658 186960
rect 452714 186904 452719 186960
rect 160553 186902 452719 186904
rect 160553 186899 160619 186902
rect 180701 186899 180767 186902
rect 452653 186899 452719 186902
rect 145373 186284 145439 186285
rect 145373 186282 145420 186284
rect 145328 186280 145420 186282
rect 145328 186224 145378 186280
rect 145328 186222 145420 186224
rect 145373 186220 145420 186222
rect 145484 186220 145490 186284
rect 145557 186282 145623 186285
rect 145741 186282 145807 186285
rect 567929 186282 567995 186285
rect 145557 186280 567995 186282
rect 145557 186224 145562 186280
rect 145618 186224 145746 186280
rect 145802 186224 567934 186280
rect 567990 186224 567995 186280
rect 145557 186222 567995 186224
rect 145373 186219 145439 186220
rect 145557 186219 145623 186222
rect 145741 186219 145807 186222
rect 567929 186219 567995 186222
rect 94497 186146 94563 186149
rect 168373 186146 168439 186149
rect 169150 186146 169156 186148
rect 94497 186144 161490 186146
rect 94497 186088 94502 186144
rect 94558 186088 161490 186144
rect 94497 186086 161490 186088
rect 94497 186083 94563 186086
rect 161430 185738 161490 186086
rect 168373 186144 169156 186146
rect 168373 186088 168378 186144
rect 168434 186088 169156 186144
rect 168373 186086 169156 186088
rect 168373 186083 168439 186086
rect 169150 186084 169156 186086
rect 169220 186084 169226 186148
rect 173750 185948 173756 186012
rect 173820 186010 173826 186012
rect 207565 186010 207631 186013
rect 173820 186008 207631 186010
rect 173820 185952 207570 186008
rect 207626 185952 207631 186008
rect 173820 185950 207631 185952
rect 173820 185948 173826 185950
rect 207565 185947 207631 185950
rect 179413 185738 179479 185741
rect 203006 185738 203012 185740
rect 161430 185736 203012 185738
rect 161430 185680 179418 185736
rect 179474 185680 203012 185736
rect 161430 185678 203012 185680
rect 179413 185675 179479 185678
rect 203006 185676 203012 185678
rect 203076 185676 203082 185740
rect 111374 185540 111380 185604
rect 111444 185602 111450 185604
rect 145557 185602 145623 185605
rect 111444 185600 145623 185602
rect 111444 185544 145562 185600
rect 145618 185544 145623 185600
rect 111444 185542 145623 185544
rect 111444 185540 111450 185542
rect 145557 185539 145623 185542
rect 174486 185540 174492 185604
rect 174556 185602 174562 185604
rect 208853 185602 208919 185605
rect 560937 185602 561003 185605
rect 174556 185600 561003 185602
rect 174556 185544 208858 185600
rect 208914 185544 560942 185600
rect 560998 185544 561003 185600
rect 174556 185542 561003 185544
rect 174556 185540 174562 185542
rect 208853 185539 208919 185542
rect 560937 185539 561003 185542
rect 107510 184996 107516 185060
rect 107580 185058 107586 185060
rect 131113 185058 131179 185061
rect 107580 185056 131179 185058
rect 107580 185000 131118 185056
rect 131174 185000 131179 185056
rect 107580 184998 131179 185000
rect 107580 184996 107586 184998
rect 131113 184995 131179 184998
rect 580165 185058 580231 185061
rect 583520 185058 584960 185148
rect 580165 185056 584960 185058
rect 580165 185000 580170 185056
rect 580226 185000 584960 185056
rect 580165 184998 584960 185000
rect 580165 184995 580231 184998
rect 138013 184922 138079 184925
rect 139158 184922 139164 184924
rect 138013 184920 139164 184922
rect 138013 184864 138018 184920
rect 138074 184864 139164 184920
rect 138013 184862 139164 184864
rect 138013 184859 138079 184862
rect 139158 184860 139164 184862
rect 139228 184922 139234 184924
rect 554037 184922 554103 184925
rect 139228 184920 554103 184922
rect 139228 184864 554042 184920
rect 554098 184864 554103 184920
rect 583520 184908 584960 184998
rect 139228 184862 554103 184864
rect 139228 184860 139234 184862
rect 554037 184859 554103 184862
rect 558269 184786 558335 184789
rect 151770 184784 558335 184786
rect 151770 184728 558274 184784
rect 558330 184728 558335 184784
rect 151770 184726 558335 184728
rect -960 184378 480 184468
rect 119838 184452 119844 184516
rect 119908 184514 119914 184516
rect 148041 184514 148107 184517
rect 119908 184512 148107 184514
rect 119908 184456 148046 184512
rect 148102 184456 148107 184512
rect 119908 184454 148107 184456
rect 119908 184452 119914 184454
rect 148041 184451 148107 184454
rect 3141 184378 3207 184381
rect -960 184376 3207 184378
rect -960 184320 3146 184376
rect 3202 184320 3207 184376
rect -960 184318 3207 184320
rect -960 184228 480 184318
rect 3141 184315 3207 184318
rect 112846 184316 112852 184380
rect 112916 184378 112922 184380
rect 146886 184378 146892 184380
rect 112916 184318 146892 184378
rect 112916 184316 112922 184318
rect 146886 184316 146892 184318
rect 146956 184378 146962 184380
rect 151770 184378 151830 184726
rect 558269 184723 558335 184726
rect 163998 184588 164004 184652
rect 164068 184650 164074 184652
rect 186037 184650 186103 184653
rect 436093 184650 436159 184653
rect 164068 184648 436159 184650
rect 164068 184592 186042 184648
rect 186098 184592 436098 184648
rect 436154 184592 436159 184648
rect 164068 184590 436159 184592
rect 164068 184588 164074 184590
rect 186037 184587 186103 184590
rect 436093 184587 436159 184590
rect 166390 184452 166396 184516
rect 166460 184514 166466 184516
rect 218421 184514 218487 184517
rect 511993 184514 512059 184517
rect 166460 184512 512059 184514
rect 166460 184456 218426 184512
rect 218482 184456 511998 184512
rect 512054 184456 512059 184512
rect 166460 184454 512059 184456
rect 166460 184452 166466 184454
rect 218421 184451 218487 184454
rect 511993 184451 512059 184454
rect 146956 184318 151830 184378
rect 146956 184316 146962 184318
rect 170990 184316 170996 184380
rect 171060 184378 171066 184380
rect 204621 184378 204687 184381
rect 548517 184378 548583 184381
rect 171060 184376 548583 184378
rect 171060 184320 204626 184376
rect 204682 184320 548522 184376
rect 548578 184320 548583 184376
rect 171060 184318 548583 184320
rect 171060 184316 171066 184318
rect 204621 184315 204687 184318
rect 548517 184315 548583 184318
rect 108246 184180 108252 184244
rect 108316 184242 108322 184244
rect 147622 184242 147628 184244
rect 108316 184182 147628 184242
rect 108316 184180 108322 184182
rect 147622 184180 147628 184182
rect 147692 184180 147698 184244
rect 168966 184180 168972 184244
rect 169036 184242 169042 184244
rect 198958 184242 198964 184244
rect 169036 184182 198964 184242
rect 169036 184180 169042 184182
rect 198958 184180 198964 184182
rect 199028 184242 199034 184244
rect 561029 184242 561095 184245
rect 199028 184240 561095 184242
rect 199028 184184 561034 184240
rect 561090 184184 561095 184240
rect 199028 184182 561095 184184
rect 199028 184180 199034 184182
rect 561029 184179 561095 184182
rect 158110 183500 158116 183564
rect 158180 183562 158186 183564
rect 219525 183562 219591 183565
rect 220169 183562 220235 183565
rect 158180 183560 220235 183562
rect 158180 183504 219530 183560
rect 219586 183504 220174 183560
rect 220230 183504 220235 183560
rect 158180 183502 220235 183504
rect 158180 183500 158186 183502
rect 219525 183499 219591 183502
rect 220169 183499 220235 183502
rect 189022 183364 189028 183428
rect 189092 183426 189098 183428
rect 189574 183426 189580 183428
rect 189092 183366 189580 183426
rect 189092 183364 189098 183366
rect 189574 183364 189580 183366
rect 189644 183426 189650 183428
rect 485773 183426 485839 183429
rect 189644 183424 485839 183426
rect 189644 183368 485778 183424
rect 485834 183368 485839 183424
rect 189644 183366 485839 183368
rect 189644 183364 189650 183366
rect 485773 183363 485839 183366
rect 152774 183228 152780 183292
rect 152844 183290 152850 183292
rect 219801 183290 219867 183293
rect 543733 183290 543799 183293
rect 152844 183288 543799 183290
rect 152844 183232 219806 183288
rect 219862 183232 543738 183288
rect 543794 183232 543799 183288
rect 152844 183230 543799 183232
rect 152844 183228 152850 183230
rect 219801 183227 219867 183230
rect 543733 183227 543799 183230
rect 154849 183154 154915 183157
rect 189022 183154 189028 183156
rect 154849 183152 189028 183154
rect 154849 183096 154854 183152
rect 154910 183096 189028 183152
rect 154849 183094 189028 183096
rect 154849 183091 154915 183094
rect 189022 183092 189028 183094
rect 189092 183092 189098 183156
rect 573357 183154 573423 183157
rect 216814 183152 573423 183154
rect 216814 183096 573362 183152
rect 573418 183096 573423 183152
rect 216814 183094 573423 183096
rect 216814 183021 216874 183094
rect 573357 183091 573423 183094
rect 154430 182956 154436 183020
rect 154500 183018 154506 183020
rect 216765 183018 216874 183021
rect 154500 183016 216874 183018
rect 154500 182960 216770 183016
rect 216826 182960 216874 183016
rect 154500 182958 216874 182960
rect 220169 183018 220235 183021
rect 576117 183018 576183 183021
rect 220169 183016 576183 183018
rect 220169 182960 220174 183016
rect 220230 182960 576122 183016
rect 576178 182960 576183 183016
rect 220169 182958 576183 182960
rect 154500 182956 154506 182958
rect 216765 182955 216831 182958
rect 220169 182955 220235 182958
rect 576117 182955 576183 182958
rect 159725 182882 159791 182885
rect 188838 182882 188844 182884
rect 159725 182880 188844 182882
rect 159725 182824 159730 182880
rect 159786 182824 188844 182880
rect 159725 182822 188844 182824
rect 159725 182819 159791 182822
rect 188838 182820 188844 182822
rect 188908 182882 188914 182884
rect 552657 182882 552723 182885
rect 188908 182880 552723 182882
rect 188908 182824 552662 182880
rect 552718 182824 552723 182880
rect 188908 182822 552723 182824
rect 188908 182820 188914 182822
rect 552657 182819 552723 182822
rect 152958 181596 152964 181660
rect 153028 181658 153034 181660
rect 219433 181658 219499 181661
rect 535453 181658 535519 181661
rect 153028 181656 535519 181658
rect 153028 181600 219438 181656
rect 219494 181600 535458 181656
rect 535514 181600 535519 181656
rect 153028 181598 535519 181600
rect 153028 181596 153034 181598
rect 219433 181595 219499 181598
rect 535453 181595 535519 181598
rect 122741 181522 122807 181525
rect 122966 181522 122972 181524
rect 122696 181520 122972 181522
rect 122696 181464 122746 181520
rect 122802 181464 122972 181520
rect 122696 181462 122972 181464
rect 122741 181459 122807 181462
rect 122966 181460 122972 181462
rect 123036 181460 123042 181524
rect 151670 181460 151676 181524
rect 151740 181522 151746 181524
rect 220077 181522 220143 181525
rect 570689 181522 570755 181525
rect 151740 181520 570755 181522
rect 151740 181464 220082 181520
rect 220138 181464 570694 181520
rect 570750 181464 570755 181520
rect 151740 181462 570755 181464
rect 151740 181460 151746 181462
rect 220077 181459 220143 181462
rect 570689 181459 570755 181462
rect 107142 181324 107148 181388
rect 107212 181386 107218 181388
rect 138013 181386 138079 181389
rect 107212 181384 138079 181386
rect 107212 181328 138018 181384
rect 138074 181328 138079 181384
rect 107212 181326 138079 181328
rect 107212 181324 107218 181326
rect 138013 181323 138079 181326
rect 150014 181324 150020 181388
rect 150084 181386 150090 181388
rect 219709 181386 219775 181389
rect 578233 181386 578299 181389
rect 150084 181384 578299 181386
rect 150084 181328 219714 181384
rect 219770 181328 578238 181384
rect 578294 181328 578299 181384
rect 150084 181326 578299 181328
rect 150084 181324 150090 181326
rect 219709 181323 219775 181326
rect 578233 181323 578299 181326
rect 106038 181188 106044 181252
rect 106108 181250 106114 181252
rect 127985 181250 128051 181253
rect 106108 181248 128051 181250
rect 106108 181192 127990 181248
rect 128046 181192 128051 181248
rect 106108 181190 128051 181192
rect 106108 181188 106114 181190
rect 127985 181187 128051 181190
rect 103278 181052 103284 181116
rect 103348 181114 103354 181116
rect 128721 181114 128787 181117
rect 103348 181112 128787 181114
rect 103348 181056 128726 181112
rect 128782 181056 128787 181112
rect 103348 181054 128787 181056
rect 103348 181052 103354 181054
rect 128721 181051 128787 181054
rect 101990 180916 101996 180980
rect 102060 180978 102066 180980
rect 129181 180978 129247 180981
rect 102060 180976 129247 180978
rect 102060 180920 129186 180976
rect 129242 180920 129247 180976
rect 102060 180918 129247 180920
rect 102060 180916 102066 180918
rect 129181 180915 129247 180918
rect 580165 180978 580231 180981
rect 583520 180978 584960 181068
rect 580165 180976 584960 180978
rect 580165 180920 580170 180976
rect 580226 180920 584960 180976
rect 580165 180918 584960 180920
rect 580165 180915 580231 180918
rect 100518 180780 100524 180844
rect 100588 180842 100594 180844
rect 128169 180842 128235 180845
rect 100588 180840 128235 180842
rect 100588 180784 128174 180840
rect 128230 180784 128235 180840
rect 583520 180828 584960 180918
rect 100588 180782 128235 180784
rect 100588 180780 100594 180782
rect 128169 180779 128235 180782
rect 122741 180706 122807 180709
rect 122696 180704 122850 180706
rect 122696 180648 122746 180704
rect 122802 180648 122850 180704
rect 122696 180646 122850 180648
rect 122741 180643 122850 180646
rect 122790 180572 122850 180643
rect 122782 180508 122788 180572
rect 122852 180508 122858 180572
rect 169334 180508 169340 180572
rect 169404 180570 169410 180572
rect 203190 180570 203196 180572
rect 169404 180510 203196 180570
rect 169404 180508 169410 180510
rect 203190 180508 203196 180510
rect 203260 180570 203266 180572
rect 204110 180570 204116 180572
rect 203260 180510 204116 180570
rect 203260 180508 203266 180510
rect 204110 180508 204116 180510
rect 204180 180508 204186 180572
rect 305637 180434 305703 180437
rect 180750 180432 305703 180434
rect -960 180298 480 180388
rect 180750 180376 305642 180432
rect 305698 180376 305703 180432
rect 180750 180374 305703 180376
rect 3233 180298 3299 180301
rect -960 180296 3299 180298
rect -960 180240 3238 180296
rect 3294 180240 3299 180296
rect -960 180238 3299 180240
rect -960 180148 480 180238
rect 3233 180235 3299 180238
rect 169201 180298 169267 180301
rect 176469 180298 176535 180301
rect 180750 180298 180810 180374
rect 305637 180371 305703 180374
rect 200614 180298 200620 180300
rect 169201 180296 180810 180298
rect 169201 180240 169206 180296
rect 169262 180240 176474 180296
rect 176530 180240 180810 180296
rect 169201 180238 180810 180240
rect 200070 180238 200620 180298
rect 169201 180235 169267 180238
rect 176469 180235 176535 180238
rect 166574 180100 166580 180164
rect 166644 180162 166650 180164
rect 200070 180162 200130 180238
rect 200614 180236 200620 180238
rect 200684 180298 200690 180300
rect 548609 180298 548675 180301
rect 200684 180296 548675 180298
rect 200684 180240 548614 180296
rect 548670 180240 548675 180296
rect 200684 180238 548675 180240
rect 200684 180236 200690 180238
rect 548609 180235 548675 180238
rect 166644 180102 200130 180162
rect 166644 180100 166650 180102
rect 204110 180100 204116 180164
rect 204180 180162 204186 180164
rect 582833 180162 582899 180165
rect 204180 180160 582899 180162
rect 204180 180104 582838 180160
rect 582894 180104 582899 180160
rect 204180 180102 582899 180104
rect 204180 180100 204186 180102
rect 582833 180099 582899 180102
rect 166758 179964 166764 180028
rect 166828 180026 166834 180028
rect 200798 180026 200804 180028
rect 166828 179966 200804 180026
rect 166828 179964 166834 179966
rect 200798 179964 200804 179966
rect 200868 180026 200874 180028
rect 582741 180026 582807 180029
rect 200868 180024 582807 180026
rect 200868 179968 582746 180024
rect 582802 179968 582807 180024
rect 200868 179966 582807 179968
rect 200868 179964 200874 179966
rect 582741 179963 582807 179966
rect 165286 179284 165292 179348
rect 165356 179346 165362 179348
rect 188337 179346 188403 179349
rect 165356 179344 190470 179346
rect 165356 179288 188342 179344
rect 188398 179288 190470 179344
rect 165356 179286 190470 179288
rect 165356 179284 165362 179286
rect 188337 179283 188403 179286
rect 162485 179210 162551 179213
rect 187182 179210 187188 179212
rect 162485 179208 187188 179210
rect 162485 179152 162490 179208
rect 162546 179152 187188 179208
rect 162485 179150 187188 179152
rect 162485 179147 162551 179150
rect 187182 179148 187188 179150
rect 187252 179148 187258 179212
rect 156045 179074 156111 179077
rect 186078 179074 186084 179076
rect 156045 179072 186084 179074
rect 156045 179016 156050 179072
rect 156106 179016 186084 179072
rect 156045 179014 186084 179016
rect 156045 179011 156111 179014
rect 186078 179012 186084 179014
rect 186148 179012 186154 179076
rect 190410 179074 190470 179286
rect 235993 179074 236059 179077
rect 190410 179072 236059 179074
rect 190410 179016 235998 179072
rect 236054 179016 236059 179072
rect 190410 179014 236059 179016
rect 235993 179011 236059 179014
rect 134374 178876 134380 178940
rect 134444 178938 134450 178940
rect 134517 178938 134583 178941
rect 134444 178936 134583 178938
rect 134444 178880 134522 178936
rect 134578 178880 134583 178936
rect 134444 178878 134583 178880
rect 134444 178876 134450 178878
rect 134517 178875 134583 178878
rect 161238 178876 161244 178940
rect 161308 178938 161314 178940
rect 221181 178938 221247 178941
rect 459553 178938 459619 178941
rect 161308 178936 459619 178938
rect 161308 178880 221186 178936
rect 221242 178880 459558 178936
rect 459614 178880 459619 178936
rect 161308 178878 459619 178880
rect 161308 178876 161314 178878
rect 221181 178875 221247 178878
rect 459553 178875 459619 178878
rect 161054 178740 161060 178804
rect 161124 178802 161130 178804
rect 212901 178802 212967 178805
rect 463693 178802 463759 178805
rect 161124 178800 463759 178802
rect 161124 178744 212906 178800
rect 212962 178744 463698 178800
rect 463754 178744 463759 178800
rect 161124 178742 463759 178744
rect 161124 178740 161130 178742
rect 212901 178739 212967 178742
rect 463693 178739 463759 178742
rect 163037 178666 163103 178669
rect 185158 178666 185164 178668
rect 163037 178664 185164 178666
rect 163037 178608 163042 178664
rect 163098 178608 185164 178664
rect 163037 178606 185164 178608
rect 163037 178603 163103 178606
rect 185158 178604 185164 178606
rect 185228 178666 185234 178668
rect 566825 178666 566891 178669
rect 185228 178664 566891 178666
rect 185228 178608 566830 178664
rect 566886 178608 566891 178664
rect 185228 178606 566891 178608
rect 185228 178604 185234 178606
rect 566825 178603 566891 178606
rect 97574 178060 97580 178124
rect 97644 178122 97650 178124
rect 126605 178122 126671 178125
rect 97644 178120 126671 178122
rect 97644 178064 126610 178120
rect 126666 178064 126671 178120
rect 97644 178062 126671 178064
rect 97644 178060 97650 178062
rect 126605 178059 126671 178062
rect 121126 177924 121132 177988
rect 121196 177986 121202 177988
rect 542997 177986 543063 177989
rect 121196 177984 543063 177986
rect 121196 177928 543002 177984
rect 543058 177928 543063 177984
rect 121196 177926 543063 177928
rect 121196 177924 121202 177926
rect 542997 177923 543063 177926
rect 140630 177850 140636 177852
rect 122790 177790 140636 177850
rect 113030 177380 113036 177444
rect 113100 177442 113106 177444
rect 122790 177442 122850 177790
rect 140630 177788 140636 177790
rect 140700 177850 140706 177852
rect 554129 177850 554195 177853
rect 140700 177848 554195 177850
rect 140700 177792 554134 177848
rect 554190 177792 554195 177848
rect 140700 177790 554195 177792
rect 140700 177788 140706 177790
rect 554129 177787 554195 177790
rect 476757 177714 476823 177717
rect 113100 177382 122850 177442
rect 142110 177712 476823 177714
rect 142110 177656 476762 177712
rect 476818 177656 476823 177712
rect 142110 177654 476823 177656
rect 113100 177380 113106 177382
rect 104382 177244 104388 177308
rect 104452 177306 104458 177308
rect 138606 177306 138612 177308
rect 104452 177246 138612 177306
rect 104452 177244 104458 177246
rect 138606 177244 138612 177246
rect 138676 177306 138682 177308
rect 142110 177306 142170 177654
rect 476757 177651 476823 177654
rect 138676 177246 142170 177306
rect 138676 177244 138682 177246
rect 579797 176898 579863 176901
rect 583520 176898 584960 176988
rect 579797 176896 584960 176898
rect 579797 176840 579802 176896
rect 579858 176840 584960 176896
rect 579797 176838 584960 176840
rect 579797 176835 579863 176838
rect 583520 176748 584960 176838
rect 135846 176564 135852 176628
rect 135916 176626 135922 176628
rect 136541 176626 136607 176629
rect 135916 176624 136607 176626
rect 135916 176568 136546 176624
rect 136602 176568 136607 176624
rect 135916 176566 136607 176568
rect 135916 176564 135922 176566
rect 136541 176563 136607 176566
rect 140773 176628 140839 176629
rect 140773 176624 140820 176628
rect 140884 176626 140890 176628
rect 140773 176568 140778 176624
rect 140773 176564 140820 176568
rect 140884 176566 140930 176626
rect 140884 176564 140890 176566
rect 140773 176563 140839 176564
rect -960 176068 480 176308
rect 140865 175266 140931 175269
rect 140998 175266 141004 175268
rect 140865 175264 141004 175266
rect 140865 175208 140870 175264
rect 140926 175208 141004 175264
rect 140865 175206 141004 175208
rect 140865 175203 140931 175206
rect 140998 175204 141004 175206
rect 141068 175204 141074 175268
rect 137318 175068 137324 175132
rect 137388 175130 137394 175132
rect 559557 175130 559623 175133
rect 137388 175128 559623 175130
rect 137388 175072 559562 175128
rect 559618 175072 559623 175128
rect 137388 175070 559623 175072
rect 137388 175068 137394 175070
rect 559557 175067 559623 175070
rect 137645 174994 137711 174997
rect 381537 174994 381603 174997
rect 137645 174992 381603 174994
rect 137645 174936 137650 174992
rect 137706 174936 381542 174992
rect 381598 174936 381603 174992
rect 137645 174934 381603 174936
rect 137645 174931 137711 174934
rect 381537 174931 381603 174934
rect 122046 174796 122052 174860
rect 122116 174858 122122 174860
rect 556797 174858 556863 174861
rect 122116 174856 556863 174858
rect 122116 174800 556802 174856
rect 556858 174800 556863 174856
rect 122116 174798 556863 174800
rect 122116 174796 122122 174798
rect 556797 174795 556863 174798
rect 102910 174660 102916 174724
rect 102980 174722 102986 174724
rect 137645 174722 137711 174725
rect 102980 174720 137711 174722
rect 102980 174664 137650 174720
rect 137706 174664 137711 174720
rect 102980 174662 137711 174664
rect 102980 174660 102986 174662
rect 137645 174659 137711 174662
rect 103094 174524 103100 174588
rect 103164 174586 103170 174588
rect 137318 174586 137324 174588
rect 103164 174526 137324 174586
rect 103164 174524 103170 174526
rect 137318 174524 137324 174526
rect 137388 174524 137394 174588
rect 580257 172818 580323 172821
rect 583520 172818 584960 172908
rect 580257 172816 584960 172818
rect 580257 172760 580262 172816
rect 580318 172760 584960 172816
rect 580257 172758 584960 172760
rect 580257 172755 580323 172758
rect 583520 172668 584960 172758
rect -960 172138 480 172228
rect 3233 172138 3299 172141
rect -960 172136 3299 172138
rect -960 172080 3238 172136
rect 3294 172080 3299 172136
rect -960 172078 3299 172080
rect -960 171988 480 172078
rect 3233 172075 3299 172078
rect 122741 171188 122807 171189
rect 122741 171186 122788 171188
rect 122696 171184 122788 171186
rect 122852 171186 122858 171188
rect 122696 171128 122746 171184
rect 122696 171126 122788 171128
rect 122741 171124 122788 171126
rect 122852 171126 122934 171186
rect 122852 171124 122858 171126
rect 122741 171123 122807 171124
rect 122741 171052 122807 171053
rect 122741 171050 122788 171052
rect 122696 171048 122788 171050
rect 122852 171050 122858 171052
rect 122696 170992 122746 171048
rect 122696 170990 122788 170992
rect 122741 170988 122788 170990
rect 122852 170990 122934 171050
rect 122852 170988 122858 170990
rect 122741 170987 122807 170988
rect 580349 168738 580415 168741
rect 583520 168738 584960 168828
rect 580349 168736 584960 168738
rect 580349 168680 580354 168736
rect 580410 168680 584960 168736
rect 580349 168678 584960 168680
rect 580349 168675 580415 168678
rect 583520 168588 584960 168678
rect -960 168058 480 168148
rect 3325 168058 3391 168061
rect -960 168056 3391 168058
rect -960 168000 3330 168056
rect 3386 168000 3391 168056
rect -960 167998 3391 168000
rect -960 167908 480 167998
rect 3325 167995 3391 167998
rect 580165 164658 580231 164661
rect 583520 164658 584960 164748
rect 580165 164656 584960 164658
rect 580165 164600 580170 164656
rect 580226 164600 584960 164656
rect 580165 164598 584960 164600
rect 580165 164595 580231 164598
rect 583520 164508 584960 164598
rect -960 163978 480 164068
rect 3049 163978 3115 163981
rect -960 163976 3115 163978
rect -960 163920 3054 163976
rect 3110 163920 3115 163976
rect -960 163918 3115 163920
rect -960 163828 480 163918
rect 3049 163915 3115 163918
rect 122741 161530 122807 161533
rect 122966 161530 122972 161532
rect 122696 161528 122972 161530
rect 122696 161472 122746 161528
rect 122802 161472 122972 161528
rect 122696 161470 122972 161472
rect 122741 161467 122807 161470
rect 122966 161468 122972 161470
rect 123036 161468 123042 161532
rect 122741 161396 122807 161397
rect 122741 161394 122788 161396
rect 122696 161392 122788 161394
rect 122852 161394 122858 161396
rect 122696 161336 122746 161392
rect 122696 161334 122788 161336
rect 122741 161332 122788 161334
rect 122852 161334 122934 161394
rect 122852 161332 122858 161334
rect 122741 161331 122807 161332
rect 583520 160428 584960 160668
rect -960 159898 480 159988
rect 3601 159898 3667 159901
rect -960 159896 3667 159898
rect -960 159840 3606 159896
rect 3662 159840 3667 159896
rect -960 159838 3667 159840
rect -960 159748 480 159838
rect 3601 159835 3667 159838
rect 580165 157178 580231 157181
rect 583520 157178 584960 157268
rect 580165 157176 584960 157178
rect 580165 157120 580170 157176
rect 580226 157120 584960 157176
rect 580165 157118 584960 157120
rect 580165 157115 580231 157118
rect 583520 157028 584960 157118
rect -960 155818 480 155908
rect 3509 155818 3575 155821
rect -960 155816 3575 155818
rect -960 155760 3514 155816
rect 3570 155760 3575 155816
rect -960 155758 3575 155760
rect -960 155668 480 155758
rect 3509 155755 3575 155758
rect 579797 153098 579863 153101
rect 583520 153098 584960 153188
rect 579797 153096 584960 153098
rect 579797 153040 579802 153096
rect 579858 153040 584960 153096
rect 579797 153038 584960 153040
rect 579797 153035 579863 153038
rect 583520 152948 584960 153038
rect -960 152418 480 152508
rect 3601 152418 3667 152421
rect -960 152416 3667 152418
rect -960 152360 3606 152416
rect 3662 152360 3667 152416
rect -960 152358 3667 152360
rect -960 152268 480 152358
rect 3601 152355 3667 152358
rect 122782 151948 122788 152012
rect 122852 151948 122858 152012
rect 122790 151877 122850 151948
rect 122741 151874 122850 151877
rect 122696 151872 122850 151874
rect 122696 151816 122746 151872
rect 122802 151816 122850 151872
rect 122696 151814 122850 151816
rect 122741 151811 122807 151814
rect 122741 151738 122807 151741
rect 122696 151736 122850 151738
rect 122696 151680 122746 151736
rect 122802 151680 122850 151736
rect 122696 151678 122850 151680
rect 122741 151675 122850 151678
rect 122790 151604 122850 151675
rect 122782 151540 122788 151604
rect 122852 151540 122858 151604
rect 583520 148868 584960 149108
rect 111190 148684 111196 148748
rect 111260 148746 111266 148748
rect 129089 148746 129155 148749
rect 111260 148744 129155 148746
rect 111260 148688 129094 148744
rect 129150 148688 129155 148744
rect 111260 148686 129155 148688
rect 111260 148684 111266 148686
rect 129089 148683 129155 148686
rect 100334 148548 100340 148612
rect 100404 148610 100410 148612
rect 125593 148610 125659 148613
rect 100404 148608 125659 148610
rect 100404 148552 125598 148608
rect 125654 148552 125659 148608
rect 100404 148550 125659 148552
rect 100404 148548 100410 148550
rect 125593 148547 125659 148550
rect 99833 148474 99899 148477
rect 125777 148474 125843 148477
rect 99833 148472 125843 148474
rect -960 148188 480 148428
rect 99833 148416 99838 148472
rect 99894 148416 125782 148472
rect 125838 148416 125843 148472
rect 99833 148414 125843 148416
rect 99833 148411 99899 148414
rect 125777 148411 125843 148414
rect 168465 148474 168531 148477
rect 203149 148474 203215 148477
rect 168465 148472 203215 148474
rect 168465 148416 168470 148472
rect 168526 148416 203154 148472
rect 203210 148416 203215 148472
rect 168465 148414 203215 148416
rect 168465 148411 168531 148414
rect 203149 148411 203215 148414
rect 112662 148276 112668 148340
rect 112732 148338 112738 148340
rect 144126 148338 144132 148340
rect 112732 148278 144132 148338
rect 112732 148276 112738 148278
rect 144126 148276 144132 148278
rect 144196 148276 144202 148340
rect 165470 148276 165476 148340
rect 165540 148338 165546 148340
rect 202229 148338 202295 148341
rect 165540 148336 202295 148338
rect 165540 148280 202234 148336
rect 202290 148280 202295 148336
rect 165540 148278 202295 148280
rect 165540 148276 165546 148278
rect 202229 148275 202295 148278
rect 122741 147660 122807 147661
rect 122741 147656 122788 147660
rect 122852 147658 122858 147660
rect 122741 147600 122746 147656
rect 122741 147596 122788 147600
rect 122852 147598 122898 147658
rect 122852 147596 122858 147598
rect 122741 147595 122807 147596
rect 177941 146978 178007 146981
rect 197854 146978 197860 146980
rect 177941 146976 197860 146978
rect 177941 146920 177946 146976
rect 178002 146920 197860 146976
rect 177941 146918 197860 146920
rect 177941 146915 178007 146918
rect 197854 146916 197860 146918
rect 197924 146916 197930 146980
rect 112529 146026 112595 146029
rect 131849 146026 131915 146029
rect 112529 146024 131915 146026
rect 112529 145968 112534 146024
rect 112590 145968 131854 146024
rect 131910 145968 131915 146024
rect 112529 145966 131915 145968
rect 112529 145963 112595 145966
rect 131849 145963 131915 145966
rect 186037 146026 186103 146029
rect 197670 146026 197676 146028
rect 186037 146024 197676 146026
rect 186037 145968 186042 146024
rect 186098 145968 197676 146024
rect 186037 145966 197676 145968
rect 186037 145963 186103 145966
rect 197670 145964 197676 145966
rect 197740 145964 197746 146028
rect 110229 145890 110295 145893
rect 135345 145890 135411 145893
rect 110229 145888 135411 145890
rect 110229 145832 110234 145888
rect 110290 145832 135350 145888
rect 135406 145832 135411 145888
rect 110229 145830 135411 145832
rect 110229 145827 110295 145830
rect 135345 145827 135411 145830
rect 184289 145890 184355 145893
rect 196014 145890 196020 145892
rect 184289 145888 196020 145890
rect 184289 145832 184294 145888
rect 184350 145832 196020 145888
rect 184289 145830 196020 145832
rect 184289 145827 184355 145830
rect 196014 145828 196020 145830
rect 196084 145828 196090 145892
rect 120441 145754 120507 145757
rect 152273 145754 152339 145757
rect 120441 145752 152339 145754
rect 120441 145696 120446 145752
rect 120502 145696 152278 145752
rect 152334 145696 152339 145752
rect 120441 145694 152339 145696
rect 120441 145691 120507 145694
rect 152273 145691 152339 145694
rect 153929 145754 153995 145757
rect 187918 145754 187924 145756
rect 153929 145752 187924 145754
rect 153929 145696 153934 145752
rect 153990 145696 187924 145752
rect 153929 145694 187924 145696
rect 153929 145691 153995 145694
rect 187918 145692 187924 145694
rect 187988 145692 187994 145756
rect 64137 145618 64203 145621
rect 187693 145618 187759 145621
rect 64137 145616 187759 145618
rect 64137 145560 64142 145616
rect 64198 145560 187698 145616
rect 187754 145560 187759 145616
rect 64137 145558 187759 145560
rect 64137 145555 64203 145558
rect 187693 145555 187759 145558
rect 119245 144938 119311 144941
rect 125225 144938 125291 144941
rect 119245 144936 125291 144938
rect 119245 144880 119250 144936
rect 119306 144880 125230 144936
rect 125286 144880 125291 144936
rect 119245 144878 125291 144880
rect 119245 144875 119311 144878
rect 125225 144875 125291 144878
rect 580165 144938 580231 144941
rect 583520 144938 584960 145028
rect 580165 144936 584960 144938
rect 580165 144880 580170 144936
rect 580226 144880 584960 144936
rect 580165 144878 584960 144880
rect 580165 144875 580231 144878
rect 583520 144788 584960 144878
rect 176377 144394 176443 144397
rect 195513 144394 195579 144397
rect 176377 144392 195579 144394
rect -960 144258 480 144348
rect 176377 144336 176382 144392
rect 176438 144336 195518 144392
rect 195574 144336 195579 144392
rect 176377 144334 195579 144336
rect 176377 144331 176443 144334
rect 195513 144331 195579 144334
rect 3141 144258 3207 144261
rect -960 144256 3207 144258
rect -960 144200 3146 144256
rect 3202 144200 3207 144256
rect -960 144198 3207 144200
rect -960 144108 480 144198
rect 3141 144195 3207 144198
rect 111006 144196 111012 144260
rect 111076 144258 111082 144260
rect 137461 144258 137527 144261
rect 111076 144256 137527 144258
rect 111076 144200 137466 144256
rect 137522 144200 137527 144256
rect 111076 144198 137527 144200
rect 111076 144196 111082 144198
rect 137461 144195 137527 144198
rect 177941 144258 178007 144261
rect 198457 144258 198523 144261
rect 177941 144256 198523 144258
rect 177941 144200 177946 144256
rect 178002 144200 198462 144256
rect 198518 144200 198523 144256
rect 177941 144198 198523 144200
rect 177941 144195 178007 144198
rect 198457 144195 198523 144198
rect 115606 144060 115612 144124
rect 115676 144122 115682 144124
rect 149789 144122 149855 144125
rect 115676 144120 149855 144122
rect 115676 144064 149794 144120
rect 149850 144064 149855 144120
rect 115676 144062 149855 144064
rect 115676 144060 115682 144062
rect 149789 144059 149855 144062
rect 170581 144122 170647 144125
rect 199561 144122 199627 144125
rect 170581 144120 199627 144122
rect 170581 144064 170586 144120
rect 170642 144064 199566 144120
rect 199622 144064 199627 144120
rect 170581 144062 199627 144064
rect 170581 144059 170647 144062
rect 199561 144059 199627 144062
rect 186865 143442 186931 143445
rect 186998 143442 187004 143444
rect 186865 143440 187004 143442
rect 186865 143384 186870 143440
rect 186926 143384 187004 143440
rect 186865 143382 187004 143384
rect 186865 143379 186931 143382
rect 186998 143380 187004 143382
rect 187068 143380 187074 143444
rect 115105 143306 115171 143309
rect 124397 143306 124463 143309
rect 115105 143304 124463 143306
rect 115105 143248 115110 143304
rect 115166 143248 124402 143304
rect 124458 143248 124463 143304
rect 115105 143246 124463 143248
rect 115105 143243 115171 143246
rect 124397 143243 124463 143246
rect 185945 143306 186011 143309
rect 194685 143306 194751 143309
rect 185945 143304 194751 143306
rect 185945 143248 185950 143304
rect 186006 143248 194690 143304
rect 194746 143248 194751 143304
rect 185945 143246 194751 143248
rect 185945 143243 186011 143246
rect 194685 143243 194751 143246
rect 118550 143108 118556 143172
rect 118620 143170 118626 143172
rect 131113 143170 131179 143173
rect 118620 143168 131179 143170
rect 118620 143112 131118 143168
rect 131174 143112 131179 143168
rect 118620 143110 131179 143112
rect 118620 143108 118626 143110
rect 131113 143107 131179 143110
rect 173709 143170 173775 143173
rect 191966 143170 191972 143172
rect 173709 143168 191972 143170
rect 173709 143112 173714 143168
rect 173770 143112 191972 143168
rect 173709 143110 191972 143112
rect 173709 143107 173775 143110
rect 191966 143108 191972 143110
rect 192036 143108 192042 143172
rect 117681 143034 117747 143037
rect 145925 143034 145991 143037
rect 117681 143032 145991 143034
rect 117681 142976 117686 143032
rect 117742 142976 145930 143032
rect 145986 142976 145991 143032
rect 117681 142974 145991 142976
rect 117681 142971 117747 142974
rect 145925 142971 145991 142974
rect 171041 143034 171107 143037
rect 191782 143034 191788 143036
rect 171041 143032 191788 143034
rect 171041 142976 171046 143032
rect 171102 142976 191788 143032
rect 171041 142974 191788 142976
rect 171041 142971 171107 142974
rect 191782 142972 191788 142974
rect 191852 142972 191858 143036
rect 119061 142898 119127 142901
rect 153377 142898 153443 142901
rect 119061 142896 153443 142898
rect 119061 142840 119066 142896
rect 119122 142840 153382 142896
rect 153438 142840 153443 142896
rect 119061 142838 153443 142840
rect 119061 142835 119127 142838
rect 153377 142835 153443 142838
rect 163865 142898 163931 142901
rect 193305 142898 193371 142901
rect 163865 142896 193371 142898
rect 163865 142840 163870 142896
rect 163926 142840 193310 142896
rect 193366 142840 193371 142896
rect 163865 142838 193371 142840
rect 163865 142835 163931 142838
rect 193305 142835 193371 142838
rect 115013 142762 115079 142765
rect 149237 142762 149303 142765
rect 115013 142760 149303 142762
rect 115013 142704 115018 142760
rect 115074 142704 149242 142760
rect 149298 142704 149303 142760
rect 115013 142702 149303 142704
rect 115013 142699 115079 142702
rect 149237 142699 149303 142702
rect 156505 142762 156571 142765
rect 190545 142762 190611 142765
rect 156505 142760 190611 142762
rect 156505 142704 156510 142760
rect 156566 142704 190550 142760
rect 190606 142704 190611 142760
rect 156505 142702 190611 142704
rect 156505 142699 156571 142702
rect 190545 142699 190611 142702
rect 185945 142490 186011 142493
rect 186221 142490 186287 142493
rect 185945 142488 186287 142490
rect 185945 142432 185950 142488
rect 186006 142432 186226 142488
rect 186282 142432 186287 142488
rect 185945 142430 186287 142432
rect 185945 142427 186011 142430
rect 186221 142427 186287 142430
rect 113633 142218 113699 142221
rect 136817 142218 136883 142221
rect 113633 142216 136883 142218
rect 113633 142160 113638 142216
rect 113694 142160 136822 142216
rect 136878 142160 136883 142216
rect 113633 142158 136883 142160
rect 113633 142155 113699 142158
rect 136817 142155 136883 142158
rect 117681 141946 117747 141949
rect 131205 141946 131271 141949
rect 117681 141944 131271 141946
rect 117681 141888 117686 141944
rect 117742 141888 131210 141944
rect 131266 141888 131271 141944
rect 117681 141886 131271 141888
rect 117681 141883 117747 141886
rect 131205 141883 131271 141886
rect 186129 141946 186195 141949
rect 194225 141946 194291 141949
rect 186129 141944 194291 141946
rect 186129 141888 186134 141944
rect 186190 141888 194230 141944
rect 194286 141888 194291 141944
rect 186129 141886 194291 141888
rect 186129 141883 186195 141886
rect 194225 141883 194291 141886
rect 118550 141748 118556 141812
rect 118620 141810 118626 141812
rect 149697 141810 149763 141813
rect 118620 141808 149763 141810
rect 118620 141752 149702 141808
rect 149758 141752 149763 141808
rect 118620 141750 149763 141752
rect 118620 141748 118626 141750
rect 149697 141747 149763 141750
rect 183369 141810 183435 141813
rect 193305 141810 193371 141813
rect 183369 141808 193371 141810
rect 183369 141752 183374 141808
rect 183430 141752 193310 141808
rect 193366 141752 193371 141808
rect 183369 141750 193371 141752
rect 183369 141747 183435 141750
rect 193305 141747 193371 141750
rect 115422 141612 115428 141676
rect 115492 141674 115498 141676
rect 148409 141674 148475 141677
rect 115492 141672 148475 141674
rect 115492 141616 148414 141672
rect 148470 141616 148475 141672
rect 115492 141614 148475 141616
rect 115492 141612 115498 141614
rect 148409 141611 148475 141614
rect 180701 141674 180767 141677
rect 194869 141674 194935 141677
rect 180701 141672 194935 141674
rect 180701 141616 180706 141672
rect 180762 141616 194874 141672
rect 194930 141616 194935 141672
rect 180701 141614 194935 141616
rect 180701 141611 180767 141614
rect 194869 141611 194935 141614
rect 118366 141476 118372 141540
rect 118436 141538 118442 141540
rect 152365 141538 152431 141541
rect 118436 141536 152431 141538
rect 118436 141480 152370 141536
rect 152426 141480 152431 141536
rect 118436 141478 152431 141480
rect 118436 141476 118442 141478
rect 152365 141475 152431 141478
rect 155401 141538 155467 141541
rect 191598 141538 191604 141540
rect 155401 141536 191604 141538
rect 155401 141480 155406 141536
rect 155462 141480 191604 141536
rect 155401 141478 191604 141480
rect 155401 141475 155467 141478
rect 191598 141476 191604 141478
rect 191668 141476 191674 141540
rect 119286 141340 119292 141404
rect 119356 141402 119362 141404
rect 180977 141402 181043 141405
rect 119356 141400 181043 141402
rect 119356 141344 180982 141400
rect 181038 141344 181043 141400
rect 119356 141342 181043 141344
rect 119356 141340 119362 141342
rect 180977 141339 181043 141342
rect 184841 141402 184907 141405
rect 195237 141402 195303 141405
rect 184841 141400 195303 141402
rect 184841 141344 184846 141400
rect 184902 141344 195242 141400
rect 195298 141344 195303 141400
rect 184841 141342 195303 141344
rect 184841 141339 184907 141342
rect 195237 141339 195303 141342
rect 580165 140858 580231 140861
rect 583520 140858 584960 140948
rect 580165 140856 584960 140858
rect 580165 140800 580170 140856
rect 580226 140800 584960 140856
rect 580165 140798 584960 140800
rect 580165 140795 580231 140798
rect 186313 140724 186379 140725
rect 186262 140660 186268 140724
rect 186332 140722 186379 140724
rect 186332 140720 186424 140722
rect 186374 140664 186424 140720
rect 583520 140708 584960 140798
rect 186332 140662 186424 140664
rect 186332 140660 186379 140662
rect 186313 140659 186379 140660
rect 115790 140524 115796 140588
rect 115860 140586 115866 140588
rect 137277 140586 137343 140589
rect 115860 140584 137343 140586
rect 115860 140528 137282 140584
rect 137338 140528 137343 140584
rect 115860 140526 137343 140528
rect 115860 140524 115866 140526
rect 137277 140523 137343 140526
rect 173433 140586 173499 140589
rect 185894 140586 185900 140588
rect 173433 140584 185900 140586
rect 173433 140528 173438 140584
rect 173494 140528 185900 140584
rect 173433 140526 185900 140528
rect 173433 140523 173499 140526
rect 185894 140524 185900 140526
rect 185964 140524 185970 140588
rect 186037 140586 186103 140589
rect 195053 140586 195119 140589
rect 186037 140584 195119 140586
rect 186037 140528 186042 140584
rect 186098 140528 195058 140584
rect 195114 140528 195119 140584
rect 186037 140526 195119 140528
rect 186037 140523 186103 140526
rect 195053 140523 195119 140526
rect 116710 140388 116716 140452
rect 116780 140450 116786 140452
rect 146569 140450 146635 140453
rect 116780 140448 146635 140450
rect 116780 140392 146574 140448
rect 146630 140392 146635 140448
rect 116780 140390 146635 140392
rect 116780 140388 116786 140390
rect 146569 140387 146635 140390
rect 178769 140450 178835 140453
rect 191782 140450 191788 140452
rect 178769 140448 191788 140450
rect 178769 140392 178774 140448
rect 178830 140392 191788 140448
rect 178769 140390 191788 140392
rect 178769 140387 178835 140390
rect 191782 140388 191788 140390
rect 191852 140388 191858 140452
rect -960 140178 480 140268
rect 119470 140252 119476 140316
rect 119540 140314 119546 140316
rect 151118 140314 151124 140316
rect 119540 140254 151124 140314
rect 119540 140252 119546 140254
rect 151118 140252 151124 140254
rect 151188 140252 151194 140316
rect 163681 140314 163747 140317
rect 186998 140314 187004 140316
rect 163681 140312 187004 140314
rect 163681 140256 163686 140312
rect 163742 140256 187004 140312
rect 163681 140254 187004 140256
rect 163681 140251 163747 140254
rect 186998 140252 187004 140254
rect 187068 140252 187074 140316
rect 2773 140178 2839 140181
rect -960 140176 2839 140178
rect -960 140120 2778 140176
rect 2834 140120 2839 140176
rect -960 140118 2839 140120
rect -960 140028 480 140118
rect 2773 140115 2839 140118
rect 119654 140116 119660 140180
rect 119724 140178 119730 140180
rect 179597 140178 179663 140181
rect 119724 140176 179663 140178
rect 119724 140120 179602 140176
rect 179658 140120 179663 140176
rect 119724 140118 179663 140120
rect 119724 140116 119730 140118
rect 179597 140115 179663 140118
rect 181989 140178 182055 140181
rect 191281 140178 191347 140181
rect 181989 140176 191347 140178
rect 181989 140120 181994 140176
rect 182050 140120 191286 140176
rect 191342 140120 191347 140176
rect 181989 140118 191347 140120
rect 181989 140115 182055 140118
rect 191281 140115 191347 140118
rect 118182 139980 118188 140044
rect 118252 140042 118258 140044
rect 179505 140042 179571 140045
rect 118252 140040 179571 140042
rect 118252 139984 179510 140040
rect 179566 139984 179571 140040
rect 118252 139982 179571 139984
rect 118252 139980 118258 139982
rect 179505 139979 179571 139982
rect 182081 140042 182147 140045
rect 196382 140042 196388 140044
rect 182081 140040 196388 140042
rect 182081 139984 182086 140040
rect 182142 139984 196388 140040
rect 182081 139982 196388 139984
rect 182081 139979 182147 139982
rect 196382 139980 196388 139982
rect 196452 139980 196458 140044
rect 124213 139636 124279 139637
rect 124213 139632 124260 139636
rect 124324 139634 124330 139636
rect 187325 139634 187391 139637
rect 124213 139576 124218 139632
rect 124213 139572 124260 139576
rect 124324 139574 124370 139634
rect 187325 139632 188354 139634
rect 187325 139576 187330 139632
rect 187386 139576 188354 139632
rect 187325 139574 188354 139576
rect 124324 139572 124330 139574
rect 124213 139571 124279 139572
rect 187325 139571 187391 139574
rect 123158 139438 124322 139498
rect 118601 139362 118667 139365
rect 120901 139362 120967 139365
rect 123158 139362 123218 139438
rect 118601 139360 118710 139362
rect 118601 139304 118606 139360
rect 118662 139304 118710 139360
rect 118601 139299 118710 139304
rect 120901 139360 123218 139362
rect 120901 139304 120906 139360
rect 120962 139304 123218 139360
rect 120901 139302 123218 139304
rect 120901 139299 120967 139302
rect 123334 139300 123340 139364
rect 123404 139362 123410 139364
rect 123569 139362 123635 139365
rect 123404 139360 123635 139362
rect 123404 139304 123574 139360
rect 123630 139304 123635 139360
rect 123404 139302 123635 139304
rect 123404 139300 123410 139302
rect 123569 139299 123635 139302
rect 123886 139300 123892 139364
rect 123956 139362 123962 139364
rect 124121 139362 124187 139365
rect 123956 139360 124187 139362
rect 123956 139304 124126 139360
rect 124182 139304 124187 139360
rect 123956 139302 124187 139304
rect 124262 139362 124322 139438
rect 130694 139436 130700 139500
rect 130764 139498 130770 139500
rect 130837 139498 130903 139501
rect 183185 139500 183251 139501
rect 130764 139496 130903 139498
rect 130764 139440 130842 139496
rect 130898 139440 130903 139496
rect 130764 139438 130903 139440
rect 130764 139436 130770 139438
rect 130837 139435 130903 139438
rect 183134 139436 183140 139500
rect 183204 139498 183251 139500
rect 186497 139498 186563 139501
rect 186630 139498 186636 139500
rect 183204 139496 183296 139498
rect 183246 139440 183296 139496
rect 183204 139438 183296 139440
rect 183878 139438 184306 139498
rect 183204 139436 183251 139438
rect 183185 139435 183251 139436
rect 127617 139362 127683 139365
rect 129181 139362 129247 139365
rect 130837 139362 130903 139365
rect 146661 139362 146727 139365
rect 124262 139360 127683 139362
rect 124262 139304 127622 139360
rect 127678 139304 127683 139360
rect 124262 139302 127683 139304
rect 123956 139300 123962 139302
rect 124121 139299 124187 139302
rect 127617 139299 127683 139302
rect 128310 139360 129247 139362
rect 128310 139304 129186 139360
rect 129242 139304 129247 139360
rect 128310 139302 129247 139304
rect 118650 139090 118710 139299
rect 120942 139164 120948 139228
rect 121012 139226 121018 139228
rect 128310 139226 128370 139302
rect 129181 139299 129247 139302
rect 129414 139360 130903 139362
rect 129414 139304 130842 139360
rect 130898 139304 130903 139360
rect 129414 139302 130903 139304
rect 121012 139166 128370 139226
rect 121012 139164 121018 139166
rect 124254 139090 124260 139092
rect 118650 139030 124260 139090
rect 124254 139028 124260 139030
rect 124324 139028 124330 139092
rect 119337 138954 119403 138957
rect 119337 138952 128370 138954
rect 119337 138896 119342 138952
rect 119398 138896 128370 138952
rect 119337 138894 128370 138896
rect 119337 138891 119403 138894
rect 116526 138756 116532 138820
rect 116596 138818 116602 138820
rect 121729 138818 121795 138821
rect 116596 138816 121795 138818
rect 116596 138760 121734 138816
rect 121790 138760 121795 138816
rect 116596 138758 121795 138760
rect 128310 138818 128370 138894
rect 129414 138818 129474 139302
rect 130837 139299 130903 139302
rect 137970 139360 146727 139362
rect 137970 139304 146666 139360
rect 146722 139304 146727 139360
rect 137970 139302 146727 139304
rect 128310 138758 129474 138818
rect 116596 138756 116602 138758
rect 121729 138755 121795 138758
rect 116761 138682 116827 138685
rect 137970 138682 138030 139302
rect 146661 139299 146727 139302
rect 170673 139362 170739 139365
rect 176469 139364 176535 139365
rect 176469 139362 176516 139364
rect 170673 139360 171150 139362
rect 170673 139304 170678 139360
rect 170734 139304 171150 139360
rect 170673 139302 171150 139304
rect 176424 139360 176516 139362
rect 176424 139304 176474 139360
rect 176424 139302 176516 139304
rect 170673 139299 170739 139302
rect 171090 138818 171150 139302
rect 176469 139300 176516 139302
rect 176580 139300 176586 139364
rect 183093 139362 183159 139365
rect 183878 139362 183938 139438
rect 183093 139360 183938 139362
rect 183093 139304 183098 139360
rect 183154 139304 183938 139360
rect 183093 139302 183938 139304
rect 184013 139362 184079 139365
rect 184013 139360 184122 139362
rect 184013 139304 184018 139360
rect 184074 139304 184122 139360
rect 176469 139299 176535 139300
rect 183093 139299 183159 139302
rect 184013 139299 184122 139304
rect 184062 138954 184122 139299
rect 184246 139090 184306 139438
rect 186497 139496 186636 139498
rect 186497 139440 186502 139496
rect 186558 139440 186636 139496
rect 186497 139438 186636 139440
rect 186497 139435 186563 139438
rect 186630 139436 186636 139438
rect 186700 139436 186706 139500
rect 187969 139498 188035 139501
rect 187742 139496 188035 139498
rect 187742 139440 187974 139496
rect 188030 139440 188035 139496
rect 187742 139438 188035 139440
rect 187742 139226 187802 139438
rect 187969 139435 188035 139438
rect 188294 139362 188354 139574
rect 196198 139362 196204 139364
rect 188294 139302 196204 139362
rect 196198 139300 196204 139302
rect 196268 139300 196274 139364
rect 199142 139226 199148 139228
rect 187742 139166 199148 139226
rect 199142 139164 199148 139166
rect 199212 139164 199218 139228
rect 195329 139090 195395 139093
rect 184246 139088 195395 139090
rect 184246 139032 195334 139088
rect 195390 139032 195395 139088
rect 184246 139030 195395 139032
rect 195329 139027 195395 139030
rect 202321 138954 202387 138957
rect 184062 138952 202387 138954
rect 184062 138896 202326 138952
rect 202382 138896 202387 138952
rect 184062 138894 202387 138896
rect 202321 138891 202387 138894
rect 191097 138818 191163 138821
rect 171090 138816 191163 138818
rect 171090 138760 191102 138816
rect 191158 138760 191163 138816
rect 171090 138758 191163 138760
rect 191097 138755 191163 138758
rect 116761 138680 138030 138682
rect 116761 138624 116766 138680
rect 116822 138624 138030 138680
rect 116761 138622 138030 138624
rect 116761 138619 116827 138622
rect 176510 138620 176516 138684
rect 176580 138682 176586 138684
rect 201718 138682 201724 138684
rect 176580 138622 201724 138682
rect 176580 138620 176586 138622
rect 201718 138620 201724 138622
rect 201788 138620 201794 138684
rect 121729 138546 121795 138549
rect 130694 138546 130700 138548
rect 121729 138544 130700 138546
rect 121729 138488 121734 138544
rect 121790 138488 130700 138544
rect 121729 138486 130700 138488
rect 121729 138483 121795 138486
rect 130694 138484 130700 138486
rect 130764 138484 130770 138548
rect 183134 138484 183140 138548
rect 183204 138546 183210 138548
rect 191966 138546 191972 138548
rect 183204 138486 191972 138546
rect 183204 138484 183210 138486
rect 191966 138484 191972 138486
rect 192036 138484 192042 138548
rect 121729 138138 121795 138141
rect 122782 138138 122788 138140
rect 121729 138136 122788 138138
rect 121729 138080 121734 138136
rect 121790 138080 122788 138136
rect 121729 138078 122788 138080
rect 121729 138075 121795 138078
rect 122782 138076 122788 138078
rect 122852 138076 122858 138140
rect 185158 138076 185164 138140
rect 185228 138138 185234 138140
rect 187366 138138 187372 138140
rect 185228 138078 187372 138138
rect 185228 138076 185234 138078
rect 187366 138076 187372 138078
rect 187436 138076 187442 138140
rect 186630 137940 186636 138004
rect 186700 138002 186706 138004
rect 190637 138002 190703 138005
rect 186700 138000 190703 138002
rect 186700 137944 190642 138000
rect 190698 137944 190703 138000
rect 186700 137942 190703 137944
rect 186700 137940 186706 137942
rect 190637 137939 190703 137942
rect 182766 137804 182772 137868
rect 182836 137866 182842 137868
rect 186814 137866 186820 137868
rect 182836 137806 186820 137866
rect 182836 137804 182842 137806
rect 186814 137804 186820 137806
rect 186884 137804 186890 137868
rect 188838 137532 188844 137596
rect 188908 137594 188914 137596
rect 193438 137594 193444 137596
rect 188908 137534 193444 137594
rect 188908 137532 188914 137534
rect 193438 137532 193444 137534
rect 193508 137532 193514 137596
rect 187182 137396 187188 137460
rect 187252 137458 187258 137460
rect 196341 137458 196407 137461
rect 187252 137456 196407 137458
rect 187252 137400 196346 137456
rect 196402 137400 196407 137456
rect 187252 137398 196407 137400
rect 187252 137396 187258 137398
rect 196341 137395 196407 137398
rect 186262 137260 186268 137324
rect 186332 137322 186338 137324
rect 199101 137322 199167 137325
rect 186332 137320 199167 137322
rect 186332 137264 199106 137320
rect 199162 137264 199167 137320
rect 186332 137262 199167 137264
rect 186332 137260 186338 137262
rect 199101 137259 199167 137262
rect 186262 136580 186268 136644
rect 186332 136642 186338 136644
rect 191005 136642 191071 136645
rect 186332 136640 191071 136642
rect 186332 136584 191010 136640
rect 191066 136584 191071 136640
rect 583520 136628 584960 136868
rect 186332 136582 191071 136584
rect 186332 136580 186338 136582
rect 191005 136579 191071 136582
rect -960 136098 480 136188
rect 3509 136098 3575 136101
rect -960 136096 3575 136098
rect -960 136040 3514 136096
rect 3570 136040 3575 136096
rect -960 136038 3575 136040
rect -960 135948 480 136038
rect 3509 136035 3575 136038
rect 113582 136036 113588 136100
rect 113652 136098 113658 136100
rect 123334 136098 123340 136100
rect 113652 136038 123340 136098
rect 113652 136036 113658 136038
rect 123334 136036 123340 136038
rect 123404 136036 123410 136100
rect 105445 135962 105511 135965
rect 121729 135962 121795 135965
rect 105445 135960 121795 135962
rect 105445 135904 105450 135960
rect 105506 135904 121734 135960
rect 121790 135904 121795 135960
rect 105445 135902 121795 135904
rect 105445 135899 105511 135902
rect 121729 135899 121795 135902
rect 187366 135900 187372 135964
rect 187436 135962 187442 135964
rect 198181 135962 198247 135965
rect 187436 135960 198247 135962
rect 187436 135904 198186 135960
rect 198242 135904 198247 135960
rect 187436 135902 198247 135904
rect 187436 135900 187442 135902
rect 198181 135899 198247 135902
rect 186078 134404 186084 134468
rect 186148 134466 186154 134468
rect 196801 134466 196867 134469
rect 186148 134464 196867 134466
rect 186148 134408 196806 134464
rect 196862 134408 196867 134464
rect 186148 134406 196867 134408
rect 186148 134404 186154 134406
rect 196801 134403 196867 134406
rect 186078 133724 186084 133788
rect 186148 133786 186154 133788
rect 188705 133786 188771 133789
rect 186148 133784 188771 133786
rect 186148 133728 188710 133784
rect 188766 133728 188771 133784
rect 186148 133726 188771 133728
rect 186148 133724 186154 133726
rect 188705 133723 188771 133726
rect 579797 132698 579863 132701
rect 583520 132698 584960 132788
rect 579797 132696 584960 132698
rect 579797 132640 579802 132696
rect 579858 132640 584960 132696
rect 579797 132638 584960 132640
rect 579797 132635 579863 132638
rect 583520 132548 584960 132638
rect -960 132018 480 132108
rect 3325 132018 3391 132021
rect -960 132016 3391 132018
rect -960 131960 3330 132016
rect 3386 131960 3391 132016
rect -960 131958 3391 131960
rect -960 131868 480 131958
rect 3325 131955 3391 131958
rect 580625 128618 580691 128621
rect 583520 128618 584960 128708
rect 580625 128616 584960 128618
rect 580625 128560 580630 128616
rect 580686 128560 584960 128616
rect 580625 128558 584960 128560
rect 580625 128555 580691 128558
rect 583520 128468 584960 128558
rect -960 127938 480 128028
rect 3417 127938 3483 127941
rect -960 127936 3483 127938
rect -960 127880 3422 127936
rect 3478 127880 3483 127936
rect -960 127878 3483 127880
rect -960 127788 480 127878
rect 3417 127875 3483 127878
rect 583520 124388 584960 124628
rect -960 123858 480 123948
rect 3417 123858 3483 123861
rect -960 123856 3483 123858
rect -960 123800 3422 123856
rect 3478 123800 3483 123856
rect -960 123798 3483 123800
rect -960 123708 480 123798
rect 3417 123795 3483 123798
rect 583520 120988 584960 121228
rect -960 119778 480 119868
rect 3325 119778 3391 119781
rect -960 119776 3391 119778
rect -960 119720 3330 119776
rect 3386 119720 3391 119776
rect -960 119718 3391 119720
rect -960 119628 480 119718
rect 3325 119715 3391 119718
rect 580901 117058 580967 117061
rect 583520 117058 584960 117148
rect 580901 117056 584960 117058
rect 580901 117000 580906 117056
rect 580962 117000 584960 117056
rect 580901 116998 584960 117000
rect 580901 116995 580967 116998
rect 583520 116908 584960 116998
rect -960 116378 480 116468
rect 3509 116378 3575 116381
rect -960 116376 3575 116378
rect -960 116320 3514 116376
rect 3570 116320 3575 116376
rect -960 116318 3575 116320
rect -960 116228 480 116318
rect 3509 116315 3575 116318
rect 580809 112978 580875 112981
rect 583520 112978 584960 113068
rect 580809 112976 584960 112978
rect 580809 112920 580814 112976
rect 580870 112920 584960 112976
rect 580809 112918 584960 112920
rect 580809 112915 580875 112918
rect 583520 112828 584960 112918
rect -960 112298 480 112388
rect 3325 112298 3391 112301
rect -960 112296 3391 112298
rect -960 112240 3330 112296
rect 3386 112240 3391 112296
rect -960 112238 3391 112240
rect -960 112148 480 112238
rect 3325 112235 3391 112238
rect 580165 108898 580231 108901
rect 583520 108898 584960 108988
rect 580165 108896 584960 108898
rect 580165 108840 580170 108896
rect 580226 108840 584960 108896
rect 580165 108838 584960 108840
rect 580165 108835 580231 108838
rect 583520 108748 584960 108838
rect -960 108218 480 108308
rect 3049 108218 3115 108221
rect -960 108216 3115 108218
rect -960 108160 3054 108216
rect 3110 108160 3115 108216
rect -960 108158 3115 108160
rect -960 108068 480 108158
rect 3049 108155 3115 108158
rect 580809 104818 580875 104821
rect 583520 104818 584960 104908
rect 580809 104816 584960 104818
rect 580809 104760 580814 104816
rect 580870 104760 584960 104816
rect 580809 104758 584960 104760
rect 580809 104755 580875 104758
rect 583520 104668 584960 104758
rect -960 104138 480 104228
rect 2957 104138 3023 104141
rect -960 104136 3023 104138
rect -960 104080 2962 104136
rect 3018 104080 3023 104136
rect -960 104078 3023 104080
rect -960 103988 480 104078
rect 2957 104075 3023 104078
rect 188889 104138 188955 104141
rect 197854 104138 197860 104140
rect 188889 104136 197860 104138
rect 188889 104080 188894 104136
rect 188950 104080 197860 104136
rect 188889 104078 197860 104080
rect 188889 104075 188955 104078
rect 197854 104076 197860 104078
rect 197924 104076 197930 104140
rect 580901 100738 580967 100741
rect 583520 100738 584960 100828
rect 580901 100736 584960 100738
rect 580901 100680 580906 100736
rect 580962 100680 584960 100736
rect 580901 100678 584960 100680
rect 580901 100675 580967 100678
rect 583520 100588 584960 100678
rect -960 100058 480 100148
rect 2865 100058 2931 100061
rect -960 100056 2931 100058
rect -960 100000 2870 100056
rect 2926 100000 2931 100056
rect -960 99998 2931 100000
rect -960 99908 480 99998
rect 2865 99995 2931 99998
rect 580625 96658 580691 96661
rect 583520 96658 584960 96748
rect 580625 96656 584960 96658
rect 580625 96600 580630 96656
rect 580686 96600 584960 96656
rect 580625 96598 584960 96600
rect 580625 96595 580691 96598
rect 583520 96508 584960 96598
rect -960 95978 480 96068
rect 2957 95978 3023 95981
rect -960 95976 3023 95978
rect -960 95920 2962 95976
rect 3018 95920 3023 95976
rect -960 95918 3023 95920
rect -960 95828 480 95918
rect 2957 95915 3023 95918
rect 119245 95162 119311 95165
rect 120574 95162 120580 95164
rect 119245 95160 120580 95162
rect 119245 95104 119250 95160
rect 119306 95104 120580 95160
rect 119245 95102 120580 95104
rect 119245 95099 119311 95102
rect 120574 95100 120580 95102
rect 120644 95100 120650 95164
rect 580717 92578 580783 92581
rect 583520 92578 584960 92668
rect 580717 92576 584960 92578
rect 580717 92520 580722 92576
rect 580778 92520 584960 92576
rect 580717 92518 584960 92520
rect 580717 92515 580783 92518
rect 583520 92428 584960 92518
rect -960 91898 480 91988
rect 3049 91898 3115 91901
rect -960 91896 3115 91898
rect -960 91840 3054 91896
rect 3110 91840 3115 91896
rect -960 91838 3115 91840
rect -960 91748 480 91838
rect 3049 91835 3115 91838
rect 186998 91836 187004 91900
rect 187068 91898 187074 91900
rect 192661 91898 192727 91901
rect 187068 91896 192727 91898
rect 187068 91840 192666 91896
rect 192722 91840 192727 91896
rect 187068 91838 192727 91840
rect 187068 91836 187074 91838
rect 192661 91835 192727 91838
rect 186078 91156 186084 91220
rect 186148 91218 186154 91220
rect 187182 91218 187188 91220
rect 186148 91158 187188 91218
rect 186148 91156 186154 91158
rect 187182 91156 187188 91158
rect 187252 91156 187258 91220
rect 119429 89858 119495 89861
rect 121729 89858 121795 89861
rect 119429 89856 121795 89858
rect 119429 89800 119434 89856
rect 119490 89800 121734 89856
rect 121790 89800 121795 89856
rect 119429 89798 121795 89800
rect 119429 89795 119495 89798
rect 121729 89795 121795 89798
rect 580717 88498 580783 88501
rect 583520 88498 584960 88588
rect 580717 88496 584960 88498
rect 580717 88440 580722 88496
rect 580778 88440 584960 88496
rect 580717 88438 584960 88440
rect 580717 88435 580783 88438
rect 186814 88300 186820 88364
rect 186884 88362 186890 88364
rect 190085 88362 190151 88365
rect 186884 88360 190151 88362
rect 186884 88304 190090 88360
rect 190146 88304 190151 88360
rect 583520 88348 584960 88438
rect 186884 88302 190151 88304
rect 186884 88300 186890 88302
rect 190085 88299 190151 88302
rect -960 87818 480 87908
rect 3509 87818 3575 87821
rect -960 87816 3575 87818
rect -960 87760 3514 87816
rect 3570 87760 3575 87816
rect -960 87758 3575 87760
rect -960 87668 480 87758
rect 3509 87755 3575 87758
rect 580533 84418 580599 84421
rect 583520 84418 584960 84508
rect 580533 84416 584960 84418
rect 580533 84360 580538 84416
rect 580594 84360 584960 84416
rect 580533 84358 584960 84360
rect 580533 84355 580599 84358
rect 583520 84268 584960 84358
rect -960 83738 480 83828
rect 3509 83738 3575 83741
rect -960 83736 3575 83738
rect -960 83680 3514 83736
rect 3570 83680 3575 83736
rect -960 83678 3575 83680
rect -960 83588 480 83678
rect 3509 83675 3575 83678
rect 186998 83404 187004 83468
rect 187068 83466 187074 83468
rect 196801 83466 196867 83469
rect 187068 83464 196867 83466
rect 187068 83408 196806 83464
rect 196862 83408 196867 83464
rect 187068 83406 196867 83408
rect 187068 83404 187074 83406
rect 196801 83403 196867 83406
rect 189390 82180 189396 82244
rect 189460 82242 189466 82244
rect 217041 82242 217107 82245
rect 189460 82240 217107 82242
rect 189460 82184 217046 82240
rect 217102 82184 217107 82240
rect 189460 82182 217107 82184
rect 189460 82180 189466 82182
rect 217041 82179 217107 82182
rect 186078 82044 186084 82108
rect 186148 82106 186154 82108
rect 217409 82106 217475 82109
rect 186148 82104 217475 82106
rect 186148 82048 217414 82104
rect 217470 82048 217475 82104
rect 186148 82046 217475 82048
rect 186148 82044 186154 82046
rect 217409 82043 217475 82046
rect 96981 81970 97047 81973
rect 133454 81970 133460 81972
rect 96981 81968 133460 81970
rect 96981 81912 96986 81968
rect 97042 81912 133460 81968
rect 96981 81910 133460 81912
rect 96981 81907 97047 81910
rect 133454 81908 133460 81910
rect 133524 81908 133530 81972
rect 172646 81908 172652 81972
rect 172716 81970 172722 81972
rect 204989 81970 205055 81973
rect 172716 81968 205055 81970
rect 172716 81912 204994 81968
rect 205050 81912 205055 81968
rect 172716 81910 205055 81912
rect 172716 81908 172722 81910
rect 204989 81907 205055 81910
rect 101213 81834 101279 81837
rect 132166 81834 132172 81836
rect 101213 81832 132172 81834
rect 101213 81776 101218 81832
rect 101274 81776 132172 81832
rect 101213 81774 132172 81776
rect 101213 81771 101279 81774
rect 132166 81772 132172 81774
rect 132236 81772 132242 81836
rect 175222 81772 175228 81836
rect 175292 81834 175298 81836
rect 199142 81834 199148 81836
rect 175292 81774 199148 81834
rect 175292 81772 175298 81774
rect 199142 81772 199148 81774
rect 199212 81772 199218 81836
rect 116669 81698 116735 81701
rect 129774 81698 129780 81700
rect 116669 81696 129780 81698
rect 116669 81640 116674 81696
rect 116730 81640 129780 81696
rect 116669 81638 129780 81640
rect 116669 81635 116735 81638
rect 129774 81636 129780 81638
rect 129844 81636 129850 81700
rect 185526 81636 185532 81700
rect 185596 81698 185602 81700
rect 206369 81698 206435 81701
rect 185596 81696 206435 81698
rect 185596 81640 206374 81696
rect 206430 81640 206435 81696
rect 185596 81638 206435 81640
rect 185596 81636 185602 81638
rect 206369 81635 206435 81638
rect 122046 81364 122052 81428
rect 122116 81426 122122 81428
rect 135478 81426 135484 81428
rect 122116 81366 135484 81426
rect 122116 81364 122122 81366
rect 135478 81364 135484 81366
rect 135548 81364 135554 81428
rect 189901 81426 189967 81429
rect 191966 81426 191972 81428
rect 189901 81424 191972 81426
rect 189901 81368 189906 81424
rect 189962 81368 191972 81424
rect 189901 81366 191972 81368
rect 189901 81363 189967 81366
rect 191966 81364 191972 81366
rect 192036 81364 192042 81428
rect 107142 81228 107148 81292
rect 107212 81290 107218 81292
rect 138790 81290 138796 81292
rect 107212 81230 138796 81290
rect 107212 81228 107218 81230
rect 138790 81228 138796 81230
rect 138860 81228 138866 81292
rect 171910 81228 171916 81292
rect 171980 81290 171986 81292
rect 202822 81290 202828 81292
rect 171980 81230 202828 81290
rect 171980 81228 171986 81230
rect 202822 81228 202828 81230
rect 202892 81228 202898 81292
rect 119286 81092 119292 81156
rect 119356 81154 119362 81156
rect 151486 81154 151492 81156
rect 119356 81094 151492 81154
rect 119356 81092 119362 81094
rect 151486 81092 151492 81094
rect 151556 81092 151562 81156
rect 158662 81092 158668 81156
rect 158732 81154 158738 81156
rect 191782 81154 191788 81156
rect 158732 81094 191788 81154
rect 158732 81092 158738 81094
rect 191782 81092 191788 81094
rect 191852 81092 191858 81156
rect 101489 81018 101555 81021
rect 134558 81018 134564 81020
rect 101489 81016 134564 81018
rect 101489 80960 101494 81016
rect 101550 80960 134564 81016
rect 101489 80958 134564 80960
rect 101489 80955 101555 80958
rect 134558 80956 134564 80958
rect 134628 80956 134634 81020
rect 157374 80956 157380 81020
rect 157444 81018 157450 81020
rect 191281 81018 191347 81021
rect 157444 81016 191347 81018
rect 157444 80960 191286 81016
rect 191342 80960 191347 81016
rect 157444 80958 191347 80960
rect 157444 80956 157450 80958
rect 191281 80955 191347 80958
rect 580165 81018 580231 81021
rect 583520 81018 584960 81108
rect 580165 81016 584960 81018
rect 580165 80960 580170 81016
rect 580226 80960 584960 81016
rect 580165 80958 584960 80960
rect 580165 80955 580231 80958
rect 105537 80882 105603 80885
rect 139894 80882 139900 80884
rect 105537 80880 139900 80882
rect 105537 80824 105542 80880
rect 105598 80824 139900 80880
rect 105537 80822 139900 80824
rect 105537 80819 105603 80822
rect 139894 80820 139900 80822
rect 139964 80820 139970 80884
rect 164734 80820 164740 80884
rect 164804 80882 164810 80884
rect 175222 80882 175228 80884
rect 164804 80822 175228 80882
rect 164804 80820 164810 80822
rect 175222 80820 175228 80822
rect 175292 80820 175298 80884
rect 191281 80882 191347 80885
rect 212993 80882 213059 80885
rect 191281 80880 213059 80882
rect 191281 80824 191286 80880
rect 191342 80824 212998 80880
rect 213054 80824 213059 80880
rect 583520 80868 584960 80958
rect 191281 80822 213059 80824
rect 191281 80819 191347 80822
rect 212993 80819 213059 80822
rect 100334 80684 100340 80748
rect 100404 80746 100410 80748
rect 131757 80746 131823 80749
rect 132217 80748 132283 80749
rect 100404 80744 131823 80746
rect 100404 80688 131762 80744
rect 131818 80688 131823 80744
rect 100404 80686 131823 80688
rect 100404 80684 100410 80686
rect 131757 80683 131823 80686
rect 132166 80684 132172 80748
rect 132236 80746 132283 80748
rect 133822 80746 133828 80748
rect 132236 80744 133828 80746
rect 132278 80688 133828 80744
rect 132236 80686 133828 80688
rect 132236 80684 132283 80686
rect 133822 80684 133828 80686
rect 133892 80684 133898 80748
rect 152222 80684 152228 80748
rect 152292 80746 152298 80748
rect 220077 80746 220143 80749
rect 152292 80744 220143 80746
rect 152292 80688 220082 80744
rect 220138 80688 220143 80744
rect 152292 80686 220143 80688
rect 152292 80684 152298 80686
rect 132217 80683 132283 80684
rect 220077 80683 220143 80686
rect 120942 80548 120948 80612
rect 121012 80610 121018 80612
rect 123477 80610 123543 80613
rect 121012 80608 123543 80610
rect 121012 80552 123482 80608
rect 123538 80552 123543 80608
rect 121012 80550 123543 80552
rect 121012 80548 121018 80550
rect 123477 80547 123543 80550
rect 124070 80548 124076 80612
rect 124140 80610 124146 80612
rect 136582 80610 136588 80612
rect 124140 80550 136588 80610
rect 124140 80548 124146 80550
rect 136582 80548 136588 80550
rect 136652 80548 136658 80612
rect 177757 80610 177823 80613
rect 191281 80610 191347 80613
rect 177757 80608 191347 80610
rect 177757 80552 177762 80608
rect 177818 80552 191286 80608
rect 191342 80552 191347 80608
rect 177757 80550 191347 80552
rect 177757 80547 177823 80550
rect 191281 80547 191347 80550
rect 171726 80412 171732 80476
rect 171796 80474 171802 80476
rect 178585 80474 178651 80477
rect 171796 80472 178651 80474
rect 171796 80416 178590 80472
rect 178646 80416 178651 80472
rect 171796 80414 178651 80416
rect 171796 80412 171802 80414
rect 178585 80411 178651 80414
rect 187049 80474 187115 80477
rect 192150 80474 192156 80476
rect 187049 80472 192156 80474
rect 187049 80416 187054 80472
rect 187110 80416 192156 80472
rect 187049 80414 192156 80416
rect 187049 80411 187115 80414
rect 192150 80412 192156 80414
rect 192220 80412 192226 80476
rect 115422 80276 115428 80340
rect 115492 80338 115498 80340
rect 122373 80338 122439 80341
rect 115492 80336 122439 80338
rect 115492 80280 122378 80336
rect 122434 80280 122439 80336
rect 115492 80278 122439 80280
rect 115492 80276 115498 80278
rect 122373 80275 122439 80278
rect 131941 80338 132007 80341
rect 134926 80338 134932 80340
rect 131941 80336 134932 80338
rect 131941 80280 131946 80336
rect 132002 80280 134932 80336
rect 131941 80278 134932 80280
rect 131941 80275 132007 80278
rect 134926 80276 134932 80278
rect 134996 80276 135002 80340
rect 115606 80140 115612 80204
rect 115676 80202 115682 80204
rect 120717 80202 120783 80205
rect 137134 80202 137140 80204
rect 115676 80200 120783 80202
rect 115676 80144 120722 80200
rect 120778 80144 120783 80200
rect 115676 80142 120783 80144
rect 115676 80140 115682 80142
rect 120717 80139 120783 80142
rect 125550 80142 137140 80202
rect 112662 80004 112668 80068
rect 112732 80066 112738 80068
rect 112732 80006 122850 80066
rect 112732 80004 112738 80006
rect -960 79658 480 79748
rect 3509 79658 3575 79661
rect -960 79656 3575 79658
rect -960 79600 3514 79656
rect 3570 79600 3575 79656
rect -960 79598 3575 79600
rect 122790 79658 122850 80006
rect 125550 79658 125610 80142
rect 137134 80140 137140 80142
rect 137204 80140 137210 80204
rect 137502 80140 137508 80204
rect 137572 80202 137578 80204
rect 155534 80202 155540 80204
rect 137572 80142 144562 80202
rect 137572 80140 137578 80142
rect 131849 80066 131915 80069
rect 131849 80064 134304 80066
rect 131849 80008 131854 80064
rect 131910 80008 134304 80064
rect 131849 80006 134304 80008
rect 131849 80003 131915 80006
rect 126329 79930 126395 79933
rect 133091 79932 133157 79933
rect 133086 79930 133092 79932
rect 126329 79928 131130 79930
rect 126329 79872 126334 79928
rect 126390 79872 131130 79928
rect 126329 79870 131130 79872
rect 133000 79870 133092 79930
rect 126329 79867 126395 79870
rect 131070 79794 131130 79870
rect 133086 79868 133092 79870
rect 133156 79868 133162 79932
rect 133459 79928 133525 79933
rect 133643 79932 133709 79933
rect 134011 79932 134077 79933
rect 133459 79872 133464 79928
rect 133520 79872 133525 79928
rect 133091 79867 133157 79868
rect 133459 79867 133525 79872
rect 133638 79868 133644 79932
rect 133708 79930 133714 79932
rect 134006 79930 134012 79932
rect 133708 79870 133800 79930
rect 133920 79870 134012 79930
rect 133708 79868 133714 79870
rect 134006 79868 134012 79870
rect 134076 79868 134082 79932
rect 134244 79930 134304 80006
rect 140262 80004 140268 80068
rect 140332 80066 140338 80068
rect 140332 80006 142584 80066
rect 140332 80004 140338 80006
rect 134379 79962 134445 79967
rect 134379 79930 134384 79962
rect 134244 79906 134384 79930
rect 134440 79906 134445 79962
rect 134244 79901 134445 79906
rect 134747 79962 134813 79967
rect 135575 79964 135641 79967
rect 134747 79906 134752 79962
rect 134808 79906 134813 79962
rect 135532 79962 135641 79964
rect 135532 79932 135580 79962
rect 134747 79901 134813 79906
rect 134244 79870 134442 79901
rect 133643 79867 133709 79868
rect 134011 79867 134077 79868
rect 133462 79797 133522 79867
rect 132125 79794 132191 79797
rect 131070 79792 132191 79794
rect 131070 79736 132130 79792
rect 132186 79736 132191 79792
rect 131070 79734 132191 79736
rect 132125 79731 132191 79734
rect 133413 79792 133522 79797
rect 133413 79736 133418 79792
rect 133474 79736 133522 79792
rect 133413 79734 133522 79736
rect 133413 79731 133479 79734
rect 133822 79732 133828 79796
rect 133892 79794 133898 79796
rect 133965 79794 134031 79797
rect 134609 79796 134675 79797
rect 134558 79794 134564 79796
rect 133892 79792 134031 79794
rect 133892 79736 133970 79792
rect 134026 79736 134031 79792
rect 133892 79734 134031 79736
rect 134518 79734 134564 79794
rect 134628 79792 134675 79796
rect 134670 79736 134675 79792
rect 133892 79732 133898 79734
rect 133965 79731 134031 79734
rect 134558 79732 134564 79734
rect 134628 79732 134675 79736
rect 134609 79731 134675 79732
rect 122790 79598 125610 79658
rect 133137 79658 133203 79661
rect 134057 79660 134123 79661
rect 133454 79658 133460 79660
rect 133137 79656 133460 79658
rect 133137 79600 133142 79656
rect 133198 79600 133460 79656
rect 133137 79598 133460 79600
rect -960 79508 480 79598
rect 3509 79595 3575 79598
rect 133137 79595 133203 79598
rect 133454 79596 133460 79598
rect 133524 79596 133530 79660
rect 134006 79658 134012 79660
rect 133966 79598 134012 79658
rect 134076 79656 134123 79660
rect 134118 79600 134123 79656
rect 134006 79596 134012 79598
rect 134076 79596 134123 79600
rect 134057 79595 134123 79596
rect 134609 79658 134675 79661
rect 134750 79658 134810 79901
rect 135478 79868 135484 79932
rect 135548 79906 135580 79932
rect 135636 79906 135641 79962
rect 135548 79901 135641 79906
rect 135851 79962 135917 79967
rect 135851 79906 135856 79962
rect 135912 79906 135917 79962
rect 136771 79962 136837 79967
rect 135851 79901 135917 79906
rect 136127 79930 136193 79933
rect 136771 79932 136776 79962
rect 136832 79932 136837 79962
rect 137323 79962 137389 79967
rect 136398 79930 136404 79932
rect 136127 79928 136404 79930
rect 135548 79870 135592 79901
rect 135548 79868 135554 79870
rect 135854 79794 135914 79901
rect 136127 79872 136132 79928
rect 136188 79872 136404 79928
rect 136127 79870 136404 79872
rect 136127 79867 136193 79870
rect 136398 79868 136404 79870
rect 136468 79868 136474 79932
rect 136766 79868 136772 79932
rect 136836 79930 136842 79932
rect 136836 79870 136894 79930
rect 137139 79928 137205 79933
rect 137139 79872 137144 79928
rect 137200 79872 137205 79928
rect 137323 79906 137328 79962
rect 137384 79906 137389 79962
rect 137323 79901 137389 79906
rect 138059 79962 138125 79967
rect 138887 79964 138953 79967
rect 138059 79906 138064 79962
rect 138120 79906 138125 79962
rect 138844 79962 138953 79964
rect 138427 79932 138493 79933
rect 138844 79932 138892 79962
rect 138422 79930 138428 79932
rect 138059 79901 138125 79906
rect 136836 79868 136842 79870
rect 137139 79867 137205 79872
rect 137142 79797 137202 79867
rect 136817 79794 136883 79797
rect 135854 79792 136883 79794
rect 135854 79736 136822 79792
rect 136878 79736 136883 79792
rect 135854 79734 136883 79736
rect 137142 79792 137251 79797
rect 137142 79736 137190 79792
rect 137246 79736 137251 79792
rect 137142 79734 137251 79736
rect 136817 79731 136883 79734
rect 137185 79731 137251 79734
rect 134609 79656 134810 79658
rect 134609 79600 134614 79656
rect 134670 79600 134810 79656
rect 134609 79598 134810 79600
rect 134609 79595 134675 79598
rect 134926 79596 134932 79660
rect 134996 79658 135002 79660
rect 136173 79658 136239 79661
rect 134996 79656 136239 79658
rect 134996 79600 136178 79656
rect 136234 79600 136239 79656
rect 134996 79598 136239 79600
rect 134996 79596 135002 79598
rect 136173 79595 136239 79598
rect 136582 79596 136588 79660
rect 136652 79658 136658 79660
rect 136817 79658 136883 79661
rect 136652 79656 136883 79658
rect 136652 79600 136822 79656
rect 136878 79600 136883 79656
rect 136652 79598 136883 79600
rect 137326 79658 137386 79901
rect 138062 79794 138122 79901
rect 138336 79870 138428 79930
rect 138422 79868 138428 79870
rect 138492 79868 138498 79932
rect 138790 79868 138796 79932
rect 138860 79906 138892 79932
rect 138948 79906 138953 79962
rect 139531 79932 139597 79933
rect 139526 79930 139532 79932
rect 138860 79901 138953 79906
rect 138860 79870 138904 79901
rect 139440 79870 139532 79930
rect 138860 79868 138866 79870
rect 139526 79868 139532 79870
rect 139596 79868 139602 79932
rect 139715 79928 139781 79933
rect 140543 79930 140609 79933
rect 139715 79872 139720 79928
rect 139776 79872 139781 79928
rect 138427 79867 138493 79868
rect 139531 79867 139597 79868
rect 139715 79867 139781 79872
rect 140500 79928 140609 79930
rect 140500 79872 140548 79928
rect 140604 79872 140609 79928
rect 140500 79867 140609 79872
rect 140819 79928 140885 79933
rect 141095 79930 141161 79933
rect 141279 79930 141345 79933
rect 140819 79872 140824 79928
rect 140880 79872 140885 79928
rect 140819 79867 140885 79872
rect 140960 79928 141161 79930
rect 140960 79872 141100 79928
rect 141156 79872 141161 79928
rect 140960 79870 141161 79872
rect 138238 79794 138244 79796
rect 138062 79734 138244 79794
rect 138238 79732 138244 79734
rect 138308 79732 138314 79796
rect 139342 79732 139348 79796
rect 139412 79794 139418 79796
rect 139718 79794 139778 79867
rect 139412 79734 139778 79794
rect 139853 79796 139919 79797
rect 139853 79792 139900 79796
rect 139964 79794 139970 79796
rect 139853 79736 139858 79792
rect 139412 79732 139418 79734
rect 139853 79732 139900 79736
rect 139964 79734 140010 79794
rect 139964 79732 139970 79734
rect 139853 79731 139919 79732
rect 140500 79661 140560 79867
rect 137461 79658 137527 79661
rect 137326 79656 137527 79658
rect 137326 79600 137466 79656
rect 137522 79600 137527 79656
rect 137326 79598 137527 79600
rect 136652 79596 136658 79598
rect 136817 79595 136883 79598
rect 137461 79595 137527 79598
rect 140497 79656 140563 79661
rect 140497 79600 140502 79656
rect 140558 79600 140563 79656
rect 140497 79595 140563 79600
rect 105629 79522 105695 79525
rect 138289 79522 138355 79525
rect 105629 79520 138355 79522
rect 105629 79464 105634 79520
rect 105690 79464 138294 79520
rect 138350 79464 138355 79520
rect 105629 79462 138355 79464
rect 105629 79459 105695 79462
rect 138289 79459 138355 79462
rect 140822 79389 140882 79867
rect 140960 79797 141020 79870
rect 141095 79867 141161 79870
rect 141236 79928 141345 79930
rect 141236 79872 141284 79928
rect 141340 79872 141345 79928
rect 141236 79867 141345 79872
rect 141550 79868 141556 79932
rect 141620 79930 141626 79932
rect 141923 79930 141989 79933
rect 141620 79928 141989 79930
rect 141620 79872 141928 79928
rect 141984 79872 141989 79928
rect 141620 79870 141989 79872
rect 141620 79868 141626 79870
rect 141923 79867 141989 79870
rect 142102 79868 142108 79932
rect 142172 79930 142178 79932
rect 142291 79930 142357 79933
rect 142172 79928 142357 79930
rect 142172 79872 142296 79928
rect 142352 79872 142357 79928
rect 142172 79870 142357 79872
rect 142524 79930 142584 80006
rect 144502 79967 144562 80142
rect 154898 80142 155540 80202
rect 145046 80004 145052 80068
rect 145116 80066 145122 80068
rect 145116 80006 145620 80066
rect 145116 80004 145122 80006
rect 142751 79962 142817 79967
rect 142751 79930 142756 79962
rect 142524 79906 142756 79930
rect 142812 79906 142817 79962
rect 142524 79901 142817 79906
rect 143027 79962 143093 79967
rect 143027 79906 143032 79962
rect 143088 79906 143093 79962
rect 144499 79962 144565 79967
rect 143027 79901 143093 79906
rect 142524 79870 142814 79901
rect 142172 79868 142178 79870
rect 142291 79867 142357 79870
rect 140957 79792 141023 79797
rect 140957 79736 140962 79792
rect 141018 79736 141023 79792
rect 140957 79731 141023 79736
rect 141236 79661 141296 79867
rect 141233 79656 141299 79661
rect 141693 79658 141759 79661
rect 141233 79600 141238 79656
rect 141294 79600 141299 79656
rect 141233 79595 141299 79600
rect 141512 79656 141759 79658
rect 141512 79600 141698 79656
rect 141754 79600 141759 79656
rect 141512 79598 141759 79600
rect 141512 79525 141572 79598
rect 141693 79595 141759 79598
rect 142102 79596 142108 79660
rect 142172 79658 142178 79660
rect 143030 79658 143090 79901
rect 143942 79868 143948 79932
rect 144012 79930 144018 79932
rect 144223 79930 144289 79933
rect 144012 79928 144289 79930
rect 144012 79872 144228 79928
rect 144284 79872 144289 79928
rect 144499 79906 144504 79962
rect 144560 79906 144565 79962
rect 144867 79962 144933 79967
rect 144867 79932 144872 79962
rect 144928 79932 144933 79962
rect 144499 79901 144565 79906
rect 144012 79870 144289 79872
rect 144012 79868 144018 79870
rect 144223 79867 144289 79870
rect 144862 79868 144868 79932
rect 144932 79930 144938 79932
rect 144932 79870 144990 79930
rect 145327 79928 145393 79933
rect 145327 79872 145332 79928
rect 145388 79872 145393 79928
rect 144932 79868 144938 79870
rect 145327 79867 145393 79872
rect 145560 79930 145620 80006
rect 154898 79967 154958 80142
rect 155534 80140 155540 80142
rect 155604 80140 155610 80204
rect 184933 80202 184999 80205
rect 157014 80200 184999 80202
rect 157014 80144 184938 80200
rect 184994 80144 184999 80200
rect 157014 80142 184999 80144
rect 145971 79962 146037 79967
rect 146247 79964 146313 79967
rect 145971 79930 145976 79962
rect 145560 79906 145976 79930
rect 146032 79906 146037 79962
rect 146204 79962 146313 79964
rect 146204 79932 146252 79962
rect 145560 79901 146037 79906
rect 145560 79870 146034 79901
rect 146150 79868 146156 79932
rect 146220 79906 146252 79932
rect 146308 79906 146313 79962
rect 146523 79962 146589 79967
rect 146523 79932 146528 79962
rect 146584 79932 146589 79962
rect 148179 79962 148245 79967
rect 147075 79932 147141 79933
rect 146220 79901 146313 79906
rect 146220 79870 146264 79901
rect 146220 79868 146226 79870
rect 146518 79868 146524 79932
rect 146588 79930 146594 79932
rect 147070 79930 147076 79932
rect 146588 79870 146646 79930
rect 146707 79894 146773 79899
rect 146588 79868 146594 79870
rect 143574 79732 143580 79796
rect 143644 79794 143650 79796
rect 144729 79794 144795 79797
rect 145330 79794 145390 79867
rect 146707 79838 146712 79894
rect 146768 79838 146773 79894
rect 146984 79870 147076 79930
rect 147070 79868 147076 79870
rect 147140 79868 147146 79932
rect 147719 79930 147785 79933
rect 148179 79932 148184 79962
rect 148240 79932 148245 79962
rect 148363 79962 148429 79967
rect 147676 79928 147785 79930
rect 147676 79872 147724 79928
rect 147780 79872 147785 79928
rect 147075 79867 147141 79868
rect 147676 79867 147785 79872
rect 147995 79894 148061 79899
rect 146707 79833 146773 79838
rect 143644 79792 144795 79794
rect 143644 79736 144734 79792
rect 144790 79736 144795 79792
rect 143644 79734 144795 79736
rect 143644 79732 143650 79734
rect 144729 79731 144795 79734
rect 145054 79734 145390 79794
rect 143809 79658 143875 79661
rect 142172 79598 143090 79658
rect 143214 79656 143875 79658
rect 143214 79600 143814 79656
rect 143870 79600 143875 79656
rect 143214 79598 143875 79600
rect 142172 79596 142178 79598
rect 141509 79520 141575 79525
rect 141509 79464 141514 79520
rect 141570 79464 141575 79520
rect 141509 79459 141575 79464
rect 141693 79522 141759 79525
rect 143214 79522 143274 79598
rect 143809 79595 143875 79598
rect 144177 79658 144243 79661
rect 145054 79658 145114 79734
rect 144177 79656 145114 79658
rect 144177 79600 144182 79656
rect 144238 79600 145114 79656
rect 144177 79598 145114 79600
rect 146569 79658 146635 79661
rect 146710 79658 146770 79833
rect 147676 79794 147736 79867
rect 147995 79838 148000 79894
rect 148056 79838 148061 79894
rect 148174 79868 148180 79932
rect 148244 79930 148250 79932
rect 148244 79870 148302 79930
rect 148363 79906 148368 79962
rect 148424 79906 148429 79962
rect 150571 79962 150637 79967
rect 148731 79932 148797 79933
rect 148726 79930 148732 79932
rect 148363 79901 148429 79906
rect 148244 79868 148250 79870
rect 147995 79833 148061 79838
rect 147806 79794 147812 79796
rect 147676 79734 147812 79794
rect 147806 79732 147812 79734
rect 147876 79732 147882 79796
rect 146569 79656 146770 79658
rect 146569 79600 146574 79656
rect 146630 79600 146770 79656
rect 146569 79598 146770 79600
rect 147998 79658 148058 79833
rect 148366 79661 148426 79901
rect 148640 79870 148732 79930
rect 148726 79868 148732 79870
rect 148796 79868 148802 79932
rect 150571 79906 150576 79962
rect 150632 79906 150637 79962
rect 150571 79901 150637 79906
rect 150939 79962 151005 79967
rect 150939 79906 150944 79962
rect 151000 79906 151005 79962
rect 151491 79964 151557 79967
rect 151491 79962 151614 79964
rect 151491 79932 151496 79962
rect 151552 79932 151614 79962
rect 153147 79962 153213 79967
rect 153975 79964 154041 79967
rect 150939 79901 151005 79906
rect 148731 79867 148797 79868
rect 149283 79826 149349 79831
rect 149283 79770 149288 79826
rect 149344 79770 149349 79826
rect 149283 79765 149349 79770
rect 148225 79658 148291 79661
rect 147998 79656 148291 79658
rect 147998 79600 148230 79656
rect 148286 79600 148291 79656
rect 147998 79598 148291 79600
rect 148366 79656 148475 79661
rect 148366 79600 148414 79656
rect 148470 79600 148475 79656
rect 148366 79598 148475 79600
rect 144177 79595 144243 79598
rect 146569 79595 146635 79598
rect 148225 79595 148291 79598
rect 148409 79595 148475 79598
rect 141693 79520 143274 79522
rect 141693 79464 141698 79520
rect 141754 79464 143274 79520
rect 141693 79462 143274 79464
rect 149286 79525 149346 79765
rect 149421 79660 149487 79661
rect 149421 79656 149468 79660
rect 149532 79658 149538 79660
rect 149421 79600 149426 79656
rect 149421 79596 149468 79600
rect 149532 79598 149578 79658
rect 149532 79596 149538 79598
rect 149421 79595 149487 79596
rect 150574 79525 150634 79901
rect 150942 79661 151002 79901
rect 151486 79868 151492 79932
rect 151556 79904 151614 79932
rect 151556 79868 151562 79904
rect 152038 79868 152044 79932
rect 152108 79930 152114 79932
rect 152319 79930 152385 79933
rect 152108 79928 152385 79930
rect 152108 79872 152324 79928
rect 152380 79872 152385 79928
rect 152108 79870 152385 79872
rect 152108 79868 152114 79870
rect 152319 79867 152385 79870
rect 152503 79930 152569 79933
rect 152958 79930 152964 79932
rect 152503 79928 152964 79930
rect 152503 79872 152508 79928
rect 152564 79872 152964 79928
rect 152503 79870 152964 79872
rect 152503 79867 152569 79870
rect 152958 79868 152964 79870
rect 153028 79868 153034 79932
rect 153147 79906 153152 79962
rect 153208 79906 153213 79962
rect 153147 79901 153213 79906
rect 153932 79962 154041 79964
rect 153932 79906 153980 79962
rect 154036 79906 154041 79962
rect 154711 79962 154777 79967
rect 153932 79901 154041 79906
rect 154159 79930 154225 79933
rect 154430 79930 154436 79932
rect 154159 79928 154436 79930
rect 150893 79656 151002 79661
rect 150893 79600 150898 79656
rect 150954 79600 151002 79656
rect 150893 79598 151002 79600
rect 151445 79658 151511 79661
rect 153150 79658 153210 79901
rect 153791 79794 153857 79797
rect 151445 79656 153210 79658
rect 151445 79600 151450 79656
rect 151506 79600 153210 79656
rect 151445 79598 153210 79600
rect 153518 79792 153857 79794
rect 153518 79736 153796 79792
rect 153852 79736 153857 79792
rect 153518 79734 153857 79736
rect 153518 79658 153578 79734
rect 153791 79731 153857 79734
rect 153932 79661 153992 79901
rect 154159 79872 154164 79928
rect 154220 79872 154436 79928
rect 154159 79870 154436 79872
rect 154159 79867 154225 79870
rect 154430 79868 154436 79870
rect 154500 79868 154506 79932
rect 154711 79906 154716 79962
rect 154772 79906 154777 79962
rect 154711 79901 154777 79906
rect 154895 79962 154961 79967
rect 154895 79906 154900 79962
rect 154956 79906 154961 79962
rect 156091 79962 156157 79967
rect 154895 79901 154961 79906
rect 155079 79930 155145 79933
rect 155079 79928 155280 79930
rect 154714 79794 154774 79901
rect 155079 79872 155084 79928
rect 155140 79872 155280 79928
rect 155079 79870 155280 79872
rect 155079 79867 155145 79870
rect 155220 79797 155280 79870
rect 155355 79928 155421 79933
rect 155355 79872 155360 79928
rect 155416 79872 155421 79928
rect 156091 79906 156096 79962
rect 156152 79906 156157 79962
rect 156091 79901 156157 79906
rect 156275 79928 156341 79933
rect 155355 79867 155421 79872
rect 155723 79894 155789 79899
rect 154982 79794 154988 79796
rect 154714 79734 154988 79794
rect 154982 79732 154988 79734
rect 155052 79732 155058 79796
rect 155217 79792 155283 79797
rect 155217 79736 155222 79792
rect 155278 79736 155283 79792
rect 155217 79731 155283 79736
rect 153745 79658 153811 79661
rect 153518 79656 153811 79658
rect 153518 79600 153750 79656
rect 153806 79600 153811 79656
rect 153518 79598 153811 79600
rect 150893 79595 150959 79598
rect 151445 79595 151511 79598
rect 153745 79595 153811 79598
rect 153929 79656 153995 79661
rect 154665 79660 154731 79661
rect 154614 79658 154620 79660
rect 153929 79600 153934 79656
rect 153990 79600 153995 79656
rect 153929 79595 153995 79600
rect 154574 79598 154620 79658
rect 154684 79656 154731 79660
rect 154726 79600 154731 79656
rect 154614 79596 154620 79598
rect 154684 79596 154731 79600
rect 154665 79595 154731 79596
rect 149286 79520 149395 79525
rect 149286 79464 149334 79520
rect 149390 79464 149395 79520
rect 149286 79462 149395 79464
rect 150574 79520 150683 79525
rect 152181 79524 152247 79525
rect 152181 79522 152228 79524
rect 150574 79464 150622 79520
rect 150678 79464 150683 79520
rect 150574 79462 150683 79464
rect 152136 79520 152228 79522
rect 152136 79464 152186 79520
rect 152136 79462 152228 79464
rect 141693 79459 141759 79462
rect 149329 79459 149395 79462
rect 150617 79459 150683 79462
rect 152181 79460 152228 79462
rect 152292 79460 152298 79524
rect 152181 79459 152247 79460
rect 111006 79324 111012 79388
rect 111076 79386 111082 79388
rect 137553 79386 137619 79389
rect 111076 79384 137619 79386
rect 111076 79328 137558 79384
rect 137614 79328 137619 79384
rect 111076 79326 137619 79328
rect 140822 79384 140931 79389
rect 140822 79328 140870 79384
rect 140926 79328 140931 79384
rect 140822 79326 140931 79328
rect 111076 79324 111082 79326
rect 137553 79323 137619 79326
rect 140865 79323 140931 79326
rect 152549 79386 152615 79389
rect 155358 79386 155418 79867
rect 155723 79838 155728 79894
rect 155784 79838 155789 79894
rect 155723 79833 155789 79838
rect 155726 79661 155786 79833
rect 156094 79661 156154 79901
rect 156275 79872 156280 79928
rect 156336 79872 156341 79928
rect 156275 79867 156341 79872
rect 155677 79656 155786 79661
rect 155677 79600 155682 79656
rect 155738 79600 155786 79656
rect 155677 79598 155786 79600
rect 156045 79656 156154 79661
rect 156045 79600 156050 79656
rect 156106 79600 156154 79656
rect 156045 79598 156154 79600
rect 156278 79658 156338 79867
rect 157014 79831 157074 80142
rect 184933 80139 184999 80142
rect 172278 80066 172284 80068
rect 171688 80006 172284 80066
rect 171688 79967 171748 80006
rect 172278 80004 172284 80006
rect 172348 80004 172354 80068
rect 177941 80066 178007 80069
rect 177254 80064 178007 80066
rect 177254 80008 177946 80064
rect 178002 80008 178007 80064
rect 177254 80006 178007 80008
rect 157287 79964 157353 79967
rect 157287 79962 157396 79964
rect 157287 79906 157292 79962
rect 157348 79932 157396 79962
rect 157931 79962 157997 79967
rect 157348 79906 157380 79932
rect 157287 79901 157380 79906
rect 157336 79870 157380 79901
rect 157374 79868 157380 79870
rect 157444 79868 157450 79932
rect 157747 79928 157813 79933
rect 157747 79872 157752 79928
rect 157808 79872 157813 79928
rect 157931 79906 157936 79962
rect 157992 79930 157997 79962
rect 159587 79962 159653 79967
rect 158667 79932 158733 79933
rect 158478 79930 158484 79932
rect 157992 79906 158484 79930
rect 157931 79901 158484 79906
rect 157747 79867 157813 79872
rect 157934 79870 158484 79901
rect 158478 79868 158484 79870
rect 158548 79868 158554 79932
rect 158662 79868 158668 79932
rect 158732 79930 158738 79932
rect 158732 79870 158824 79930
rect 159587 79906 159592 79962
rect 159648 79906 159653 79962
rect 159587 79901 159653 79906
rect 159771 79962 159837 79967
rect 159771 79906 159776 79962
rect 159832 79906 159837 79962
rect 159771 79901 159837 79906
rect 160139 79962 160205 79967
rect 160139 79906 160144 79962
rect 160200 79906 160205 79962
rect 160783 79964 160849 79967
rect 161059 79964 161125 79967
rect 161335 79964 161401 79967
rect 160783 79962 160892 79964
rect 160139 79901 160205 79906
rect 160323 79928 160389 79933
rect 158732 79868 158738 79870
rect 158667 79867 158733 79868
rect 157011 79826 157077 79831
rect 157011 79770 157016 79826
rect 157072 79770 157077 79826
rect 157011 79765 157077 79770
rect 157750 79794 157810 79867
rect 158110 79794 158116 79796
rect 157750 79734 158116 79794
rect 158110 79732 158116 79734
rect 158180 79732 158186 79796
rect 157977 79658 158043 79661
rect 156278 79656 158043 79658
rect 156278 79600 157982 79656
rect 158038 79600 158043 79656
rect 156278 79598 158043 79600
rect 155677 79595 155743 79598
rect 156045 79595 156111 79598
rect 157977 79595 158043 79598
rect 158989 79658 159055 79661
rect 159590 79658 159650 79901
rect 158989 79656 159650 79658
rect 158989 79600 158994 79656
rect 159050 79600 159650 79656
rect 158989 79598 159650 79600
rect 159774 79658 159834 79901
rect 160142 79661 160202 79901
rect 160323 79872 160328 79928
rect 160384 79872 160389 79928
rect 160323 79867 160389 79872
rect 160599 79928 160665 79933
rect 160599 79872 160604 79928
rect 160660 79872 160665 79928
rect 160783 79906 160788 79962
rect 160844 79932 160892 79962
rect 161059 79962 161182 79964
rect 161059 79932 161064 79962
rect 161120 79932 161182 79962
rect 160844 79906 160876 79932
rect 160783 79901 160876 79906
rect 160599 79867 160665 79872
rect 160832 79870 160876 79901
rect 160870 79868 160876 79870
rect 160940 79868 160946 79932
rect 161054 79868 161060 79932
rect 161124 79904 161182 79932
rect 161335 79962 161444 79964
rect 161335 79906 161340 79962
rect 161396 79930 161444 79962
rect 161795 79962 161861 79967
rect 161606 79930 161612 79932
rect 161396 79906 161612 79930
rect 161124 79868 161130 79904
rect 161335 79901 161612 79906
rect 161384 79870 161612 79901
rect 161606 79868 161612 79870
rect 161676 79868 161682 79932
rect 161795 79906 161800 79962
rect 161856 79906 161861 79962
rect 161795 79901 161861 79906
rect 161979 79962 162045 79967
rect 161979 79906 161984 79962
rect 162040 79906 162045 79962
rect 162531 79964 162597 79967
rect 162531 79962 162654 79964
rect 162531 79932 162536 79962
rect 162592 79932 162654 79962
rect 161979 79901 162045 79906
rect 159909 79658 159975 79661
rect 159774 79656 159975 79658
rect 159774 79600 159914 79656
rect 159970 79600 159975 79656
rect 159774 79598 159975 79600
rect 160142 79656 160251 79661
rect 160142 79600 160190 79656
rect 160246 79600 160251 79656
rect 160142 79598 160251 79600
rect 160326 79658 160386 79867
rect 160602 79794 160662 79867
rect 161798 79797 161858 79901
rect 161013 79794 161079 79797
rect 160602 79792 161079 79794
rect 160602 79736 161018 79792
rect 161074 79736 161079 79792
rect 160602 79734 161079 79736
rect 161798 79792 161907 79797
rect 161798 79736 161846 79792
rect 161902 79736 161907 79792
rect 161798 79734 161907 79736
rect 161982 79794 162042 79901
rect 162526 79868 162532 79932
rect 162596 79904 162654 79932
rect 162715 79962 162781 79967
rect 162715 79906 162720 79962
rect 162776 79906 162781 79962
rect 164003 79962 164069 79967
rect 162596 79868 162602 79904
rect 162715 79901 162781 79906
rect 162899 79930 162965 79933
rect 163267 79932 163333 79933
rect 163078 79930 163084 79932
rect 162899 79928 163084 79930
rect 162117 79794 162183 79797
rect 162718 79796 162778 79901
rect 162899 79872 162904 79928
rect 162960 79872 163084 79928
rect 162899 79870 163084 79872
rect 162899 79867 162965 79870
rect 163078 79868 163084 79870
rect 163148 79868 163154 79932
rect 163262 79868 163268 79932
rect 163332 79930 163338 79932
rect 163332 79870 163424 79930
rect 164003 79906 164008 79962
rect 164064 79906 164069 79962
rect 164003 79901 164069 79906
rect 164187 79962 164253 79967
rect 164187 79906 164192 79962
rect 164248 79930 164253 79962
rect 164647 79964 164713 79967
rect 164923 79964 164989 79967
rect 164647 79962 164756 79964
rect 164366 79930 164372 79932
rect 164248 79906 164372 79930
rect 164187 79901 164372 79906
rect 163332 79868 163338 79870
rect 163267 79867 163333 79868
rect 161982 79792 162183 79794
rect 161982 79736 162122 79792
rect 162178 79736 162183 79792
rect 161982 79734 162183 79736
rect 161013 79731 161079 79734
rect 161841 79731 161907 79734
rect 162117 79731 162183 79734
rect 162710 79732 162716 79796
rect 162780 79732 162786 79796
rect 163083 79792 163149 79797
rect 163083 79736 163088 79792
rect 163144 79736 163149 79792
rect 163083 79731 163149 79736
rect 163497 79794 163563 79797
rect 163727 79794 163793 79797
rect 163497 79792 163793 79794
rect 163497 79736 163502 79792
rect 163558 79736 163732 79792
rect 163788 79736 163793 79792
rect 163497 79734 163793 79736
rect 163497 79731 163563 79734
rect 163727 79731 163793 79734
rect 161289 79658 161355 79661
rect 160326 79656 161355 79658
rect 160326 79600 161294 79656
rect 161350 79600 161355 79656
rect 160326 79598 161355 79600
rect 158989 79595 159055 79598
rect 159909 79595 159975 79598
rect 160185 79595 160251 79598
rect 161289 79595 161355 79598
rect 161933 79658 161999 79661
rect 162761 79658 162827 79661
rect 161933 79656 162827 79658
rect 161933 79600 161938 79656
rect 161994 79600 162766 79656
rect 162822 79600 162827 79656
rect 161933 79598 162827 79600
rect 163086 79658 163146 79731
rect 163313 79658 163379 79661
rect 163086 79656 163379 79658
rect 163086 79600 163318 79656
rect 163374 79600 163379 79656
rect 163086 79598 163379 79600
rect 164006 79658 164066 79901
rect 164190 79870 164372 79901
rect 164366 79868 164372 79870
rect 164436 79868 164442 79932
rect 164647 79906 164652 79962
rect 164708 79932 164756 79962
rect 164923 79962 165046 79964
rect 164923 79932 164928 79962
rect 164984 79932 165046 79962
rect 164708 79906 164740 79932
rect 164647 79901 164740 79906
rect 164696 79870 164740 79901
rect 164734 79868 164740 79870
rect 164804 79868 164810 79932
rect 164918 79868 164924 79932
rect 164988 79904 165046 79932
rect 165475 79962 165541 79967
rect 165475 79906 165480 79962
rect 165536 79906 165541 79962
rect 164988 79868 164994 79904
rect 165475 79901 165541 79906
rect 165659 79962 165725 79967
rect 165659 79906 165664 79962
rect 165720 79930 165725 79962
rect 166211 79962 166277 79967
rect 165720 79906 166090 79930
rect 165659 79901 166090 79906
rect 166211 79906 166216 79962
rect 166272 79906 166277 79962
rect 166211 79901 166277 79906
rect 166579 79962 166645 79967
rect 166579 79906 166584 79962
rect 166640 79906 166645 79962
rect 166579 79901 166645 79906
rect 167131 79962 167197 79967
rect 167131 79906 167136 79962
rect 167192 79906 167197 79962
rect 168051 79962 168117 79967
rect 167131 79901 167197 79906
rect 164279 79794 164345 79797
rect 165102 79794 165108 79796
rect 164279 79792 165108 79794
rect 164279 79736 164284 79792
rect 164340 79736 165108 79792
rect 164279 79734 165108 79736
rect 164279 79731 164345 79734
rect 165102 79732 165108 79734
rect 165172 79732 165178 79796
rect 164601 79658 164667 79661
rect 164006 79656 164667 79658
rect 164006 79600 164606 79656
rect 164662 79600 164667 79656
rect 164006 79598 164667 79600
rect 161933 79595 161999 79598
rect 162761 79595 162827 79598
rect 163313 79595 163379 79598
rect 164601 79595 164667 79598
rect 164233 79522 164299 79525
rect 164918 79522 164924 79524
rect 164233 79520 164924 79522
rect 164233 79464 164238 79520
rect 164294 79464 164924 79520
rect 164233 79462 164924 79464
rect 164233 79459 164299 79462
rect 164918 79460 164924 79462
rect 164988 79460 164994 79524
rect 152549 79384 155418 79386
rect 152549 79328 152554 79384
rect 152610 79328 155418 79384
rect 152549 79326 155418 79328
rect 155493 79386 155559 79389
rect 160686 79386 160692 79388
rect 155493 79384 160692 79386
rect 155493 79328 155498 79384
rect 155554 79328 160692 79384
rect 155493 79326 160692 79328
rect 152549 79323 152615 79326
rect 155493 79323 155559 79326
rect 160686 79324 160692 79326
rect 160756 79324 160762 79388
rect 163037 79386 163103 79389
rect 163262 79386 163268 79388
rect 163037 79384 163268 79386
rect 163037 79328 163042 79384
rect 163098 79328 163268 79384
rect 163037 79326 163268 79328
rect 163037 79323 163103 79326
rect 163262 79324 163268 79326
rect 163332 79324 163338 79388
rect 165478 79386 165538 79901
rect 165662 79870 166090 79901
rect 166030 79522 166090 79870
rect 166214 79797 166274 79901
rect 166165 79792 166274 79797
rect 166165 79736 166170 79792
rect 166226 79736 166274 79792
rect 166165 79734 166274 79736
rect 166165 79731 166231 79734
rect 166582 79658 166642 79901
rect 166855 79828 166921 79831
rect 166812 79826 166921 79828
rect 166812 79796 166860 79826
rect 166758 79732 166764 79796
rect 166828 79770 166860 79796
rect 166916 79770 166921 79826
rect 166828 79765 166921 79770
rect 167134 79794 167194 79901
rect 167678 79868 167684 79932
rect 167748 79930 167754 79932
rect 168051 79930 168056 79962
rect 167748 79906 168056 79930
rect 168112 79906 168117 79962
rect 169523 79962 169589 79967
rect 169523 79930 169528 79962
rect 167748 79901 168117 79906
rect 168376 79906 169528 79930
rect 169584 79906 169589 79962
rect 170811 79962 170877 79967
rect 168376 79901 169589 79906
rect 169891 79928 169957 79933
rect 167748 79870 168114 79901
rect 168235 79894 168301 79899
rect 167748 79868 167754 79870
rect 168235 79838 168240 79894
rect 168296 79838 168301 79894
rect 168235 79833 168301 79838
rect 168376 79870 169586 79901
rect 169891 79872 169896 79928
rect 169952 79872 169957 79928
rect 167862 79794 167868 79796
rect 166828 79734 166872 79765
rect 167134 79734 167868 79794
rect 166828 79732 166834 79734
rect 167862 79732 167868 79734
rect 167932 79732 167938 79796
rect 168238 79661 168298 79833
rect 168376 79661 168436 79870
rect 169891 79867 169957 79872
rect 170167 79930 170233 79933
rect 170438 79930 170444 79932
rect 170167 79928 170444 79930
rect 170167 79872 170172 79928
rect 170228 79872 170444 79928
rect 170167 79870 170444 79872
rect 170167 79867 170233 79870
rect 170438 79868 170444 79870
rect 170508 79868 170514 79932
rect 170811 79906 170816 79962
rect 170872 79930 170877 79962
rect 171639 79962 171748 79967
rect 170872 79906 171426 79930
rect 170811 79901 171426 79906
rect 171639 79906 171644 79962
rect 171700 79906 171748 79962
rect 172467 79962 172533 79967
rect 172467 79932 172472 79962
rect 172528 79932 172533 79962
rect 173755 79962 173821 79967
rect 171639 79904 171748 79906
rect 171639 79901 171705 79904
rect 170814 79870 171426 79901
rect 168603 79792 168669 79797
rect 168603 79736 168608 79792
rect 168664 79736 168669 79792
rect 168603 79731 168669 79736
rect 167545 79658 167611 79661
rect 166582 79656 167611 79658
rect 166582 79600 167550 79656
rect 167606 79600 167611 79656
rect 166582 79598 167611 79600
rect 167545 79595 167611 79598
rect 168189 79656 168298 79661
rect 168189 79600 168194 79656
rect 168250 79600 168298 79656
rect 168189 79598 168298 79600
rect 168373 79656 168439 79661
rect 168373 79600 168378 79656
rect 168434 79600 168439 79656
rect 168189 79595 168255 79598
rect 168373 79595 168439 79600
rect 166717 79522 166783 79525
rect 166030 79520 166783 79522
rect 166030 79464 166722 79520
rect 166778 79464 166783 79520
rect 166030 79462 166783 79464
rect 168606 79522 168666 79731
rect 169894 79658 169954 79867
rect 170806 79732 170812 79796
rect 170876 79794 170882 79796
rect 170995 79794 171061 79797
rect 170876 79792 171061 79794
rect 170876 79736 171000 79792
rect 171056 79736 171061 79792
rect 170876 79734 171061 79736
rect 170876 79732 170882 79734
rect 170995 79731 171061 79734
rect 170990 79658 170996 79660
rect 169894 79598 170996 79658
rect 170990 79596 170996 79598
rect 171060 79596 171066 79660
rect 171366 79658 171426 79870
rect 172462 79868 172468 79932
rect 172532 79930 172538 79932
rect 172651 79930 172717 79933
rect 172830 79930 172836 79932
rect 172532 79870 172590 79930
rect 172651 79928 172836 79930
rect 172651 79872 172656 79928
rect 172712 79872 172836 79928
rect 172651 79870 172836 79872
rect 172532 79868 172538 79870
rect 172651 79867 172717 79870
rect 172830 79868 172836 79870
rect 172900 79868 172906 79932
rect 173111 79930 173177 79933
rect 173755 79932 173760 79962
rect 173816 79932 173821 79962
rect 173939 79962 174005 79967
rect 173566 79930 173572 79932
rect 173111 79928 173572 79930
rect 173111 79872 173116 79928
rect 173172 79872 173572 79928
rect 173111 79870 173572 79872
rect 173111 79867 173177 79870
rect 173566 79868 173572 79870
rect 173636 79868 173642 79932
rect 173750 79868 173756 79932
rect 173820 79930 173826 79932
rect 173820 79870 173878 79930
rect 173939 79906 173944 79962
rect 174000 79930 174005 79962
rect 175227 79962 175293 79967
rect 174675 79930 174741 79933
rect 174000 79906 174554 79930
rect 173939 79901 174554 79906
rect 173942 79870 174554 79901
rect 173820 79868 173826 79870
rect 171726 79732 171732 79796
rect 171796 79794 171802 79796
rect 172007 79794 172073 79797
rect 172605 79796 172671 79797
rect 172605 79794 172652 79796
rect 171796 79792 172073 79794
rect 171796 79736 172012 79792
rect 172068 79736 172073 79792
rect 171796 79734 172073 79736
rect 172560 79792 172652 79794
rect 172560 79736 172610 79792
rect 172560 79734 172652 79736
rect 171796 79732 171802 79734
rect 172007 79731 172073 79734
rect 172605 79732 172652 79734
rect 172716 79732 172722 79796
rect 174031 79792 174097 79797
rect 174031 79736 174036 79792
rect 174092 79736 174097 79792
rect 172605 79731 172671 79732
rect 174031 79731 174097 79736
rect 174494 79794 174554 79870
rect 174675 79928 175060 79930
rect 174675 79872 174680 79928
rect 174736 79872 175060 79928
rect 175227 79906 175232 79962
rect 175288 79906 175293 79962
rect 176607 79962 176673 79967
rect 175963 79932 176029 79933
rect 175958 79930 175964 79932
rect 175227 79901 175293 79906
rect 174675 79870 175060 79872
rect 174675 79867 174741 79870
rect 174854 79794 174860 79796
rect 174494 79734 174860 79794
rect 174854 79732 174860 79734
rect 174924 79732 174930 79796
rect 171593 79658 171659 79661
rect 171366 79656 171659 79658
rect 171366 79600 171598 79656
rect 171654 79600 171659 79656
rect 171366 79598 171659 79600
rect 171593 79595 171659 79598
rect 173157 79658 173223 79661
rect 173801 79658 173867 79661
rect 173157 79656 173867 79658
rect 173157 79600 173162 79656
rect 173218 79600 173806 79656
rect 173862 79600 173867 79656
rect 173157 79598 173867 79600
rect 174034 79658 174094 79731
rect 175000 79661 175060 79870
rect 175230 79794 175290 79901
rect 175872 79870 175964 79930
rect 175958 79868 175964 79870
rect 176028 79868 176034 79932
rect 176326 79868 176332 79932
rect 176396 79930 176402 79932
rect 176607 79930 176612 79962
rect 176396 79906 176612 79930
rect 176668 79906 176673 79962
rect 176396 79901 176673 79906
rect 176883 79962 176949 79967
rect 176883 79906 176888 79962
rect 176944 79930 176949 79962
rect 177254 79930 177314 80006
rect 177941 80003 178007 80006
rect 176944 79906 177314 79930
rect 176883 79901 177314 79906
rect 176396 79870 176670 79901
rect 176886 79870 177314 79901
rect 177435 79930 177501 79933
rect 181621 79930 181687 79933
rect 177435 79928 181687 79930
rect 177435 79872 177440 79928
rect 177496 79872 181626 79928
rect 181682 79872 181687 79928
rect 177435 79870 181687 79872
rect 176396 79868 176402 79870
rect 175963 79867 176029 79868
rect 177435 79867 177501 79870
rect 181621 79867 181687 79870
rect 181529 79794 181595 79797
rect 175230 79792 181595 79794
rect 175230 79736 181534 79792
rect 181590 79736 181595 79792
rect 175230 79734 181595 79736
rect 181529 79731 181595 79734
rect 174670 79658 174676 79660
rect 174034 79598 174676 79658
rect 173157 79595 173223 79598
rect 173801 79595 173867 79598
rect 174670 79596 174676 79598
rect 174740 79596 174746 79660
rect 174997 79656 175063 79661
rect 174997 79600 175002 79656
rect 175058 79600 175063 79656
rect 174997 79595 175063 79600
rect 189390 79522 189396 79524
rect 168606 79462 189396 79522
rect 166717 79459 166783 79462
rect 189390 79460 189396 79462
rect 189460 79460 189466 79524
rect 185526 79386 185532 79388
rect 165478 79326 185532 79386
rect 185526 79324 185532 79326
rect 185596 79324 185602 79388
rect 186957 79386 187023 79389
rect 189206 79386 189212 79388
rect 186957 79384 189212 79386
rect 186957 79328 186962 79384
rect 187018 79328 189212 79384
rect 186957 79326 189212 79328
rect 186957 79323 187023 79326
rect 189206 79324 189212 79326
rect 189276 79324 189282 79388
rect 107326 79188 107332 79252
rect 107396 79250 107402 79252
rect 137369 79250 137435 79253
rect 107396 79248 137435 79250
rect 107396 79192 137374 79248
rect 137430 79192 137435 79248
rect 107396 79190 137435 79192
rect 107396 79188 107402 79190
rect 137369 79187 137435 79190
rect 154430 79188 154436 79252
rect 154500 79250 154506 79252
rect 186078 79250 186084 79252
rect 154500 79190 186084 79250
rect 154500 79188 154506 79190
rect 186078 79188 186084 79190
rect 186148 79188 186154 79252
rect 116526 79052 116532 79116
rect 116596 79114 116602 79116
rect 148317 79114 148383 79117
rect 163129 79116 163195 79117
rect 163078 79114 163084 79116
rect 116596 79112 148383 79114
rect 116596 79056 148322 79112
rect 148378 79056 148383 79112
rect 116596 79054 148383 79056
rect 163038 79054 163084 79114
rect 163148 79112 163195 79116
rect 163190 79056 163195 79112
rect 116596 79052 116602 79054
rect 148317 79051 148383 79054
rect 163078 79052 163084 79054
rect 163148 79052 163195 79056
rect 163129 79051 163195 79052
rect 169753 79114 169819 79117
rect 211613 79114 211679 79117
rect 169753 79112 211679 79114
rect 169753 79056 169758 79112
rect 169814 79056 211618 79112
rect 211674 79056 211679 79112
rect 169753 79054 211679 79056
rect 169753 79051 169819 79054
rect 211613 79051 211679 79054
rect 122414 78916 122420 78980
rect 122484 78978 122490 78980
rect 159449 78978 159515 78981
rect 122484 78976 159515 78978
rect 122484 78920 159454 78976
rect 159510 78920 159515 78976
rect 122484 78918 159515 78920
rect 122484 78916 122490 78918
rect 159449 78915 159515 78918
rect 165797 78978 165863 78981
rect 168005 78980 168071 78981
rect 171869 78980 171935 78981
rect 166758 78978 166764 78980
rect 165797 78976 166764 78978
rect 165797 78920 165802 78976
rect 165858 78920 166764 78976
rect 165797 78918 166764 78920
rect 165797 78915 165863 78918
rect 166758 78916 166764 78918
rect 166828 78916 166834 78980
rect 168005 78976 168052 78980
rect 168116 78978 168122 78980
rect 171869 78978 171916 78980
rect 168005 78920 168010 78976
rect 168005 78916 168052 78920
rect 168116 78918 168162 78978
rect 171824 78976 171916 78978
rect 171824 78920 171874 78976
rect 171824 78918 171916 78920
rect 168116 78916 168122 78918
rect 171869 78916 171916 78918
rect 171980 78916 171986 78980
rect 175273 78978 175339 78981
rect 218237 78978 218303 78981
rect 175273 78976 218303 78978
rect 175273 78920 175278 78976
rect 175334 78920 218242 78976
rect 218298 78920 218303 78976
rect 175273 78918 218303 78920
rect 168005 78915 168071 78916
rect 171869 78915 171935 78916
rect 175273 78915 175339 78918
rect 218237 78915 218303 78918
rect 108246 78780 108252 78844
rect 108316 78842 108322 78844
rect 146150 78842 146156 78844
rect 108316 78782 146156 78842
rect 108316 78780 108322 78782
rect 146150 78780 146156 78782
rect 146220 78780 146226 78844
rect 166809 78842 166875 78845
rect 218421 78842 218487 78845
rect 166809 78840 218487 78842
rect 166809 78784 166814 78840
rect 166870 78784 218426 78840
rect 218482 78784 218487 78840
rect 166809 78782 218487 78784
rect 166809 78779 166875 78782
rect 218421 78779 218487 78782
rect 133137 78708 133203 78709
rect 133086 78644 133092 78708
rect 133156 78706 133203 78708
rect 133156 78704 133248 78706
rect 133198 78648 133248 78704
rect 133156 78646 133248 78648
rect 133156 78644 133203 78646
rect 138606 78644 138612 78708
rect 138676 78706 138682 78708
rect 142153 78706 142219 78709
rect 138676 78704 142219 78706
rect 138676 78648 142158 78704
rect 142214 78648 142219 78704
rect 138676 78646 142219 78648
rect 138676 78644 138682 78646
rect 133137 78643 133203 78644
rect 142153 78643 142219 78646
rect 142286 78644 142292 78708
rect 142356 78706 142362 78708
rect 142889 78706 142955 78709
rect 142356 78704 142955 78706
rect 142356 78648 142894 78704
rect 142950 78648 142955 78704
rect 142356 78646 142955 78648
rect 142356 78644 142362 78646
rect 142889 78643 142955 78646
rect 143533 78706 143599 78709
rect 143758 78706 143764 78708
rect 143533 78704 143764 78706
rect 143533 78648 143538 78704
rect 143594 78648 143764 78704
rect 143533 78646 143764 78648
rect 143533 78643 143599 78646
rect 143758 78644 143764 78646
rect 143828 78644 143834 78708
rect 580901 78706 580967 78709
rect 144870 78704 580967 78706
rect 144870 78648 580906 78704
rect 580962 78648 580967 78704
rect 144870 78646 580967 78648
rect 119470 78508 119476 78572
rect 119540 78570 119546 78572
rect 119797 78570 119863 78573
rect 119540 78568 119863 78570
rect 119540 78512 119802 78568
rect 119858 78512 119863 78568
rect 119540 78510 119863 78512
rect 119540 78508 119546 78510
rect 119797 78507 119863 78510
rect 121126 78508 121132 78572
rect 121196 78570 121202 78572
rect 133045 78570 133111 78573
rect 121196 78568 133111 78570
rect 121196 78512 133050 78568
rect 133106 78512 133111 78568
rect 121196 78510 133111 78512
rect 121196 78508 121202 78510
rect 133045 78507 133111 78510
rect 134977 78570 135043 78573
rect 139117 78570 139183 78573
rect 139577 78572 139643 78573
rect 134977 78568 139183 78570
rect 134977 78512 134982 78568
rect 135038 78512 139122 78568
rect 139178 78512 139183 78568
rect 134977 78510 139183 78512
rect 134977 78507 135043 78510
rect 139117 78507 139183 78510
rect 139526 78508 139532 78572
rect 139596 78570 139643 78572
rect 139596 78568 139688 78570
rect 139638 78512 139688 78568
rect 139596 78510 139688 78512
rect 139596 78508 139643 78510
rect 141550 78508 141556 78572
rect 141620 78570 141626 78572
rect 141877 78570 141943 78573
rect 141620 78568 141943 78570
rect 141620 78512 141882 78568
rect 141938 78512 141943 78568
rect 141620 78510 141943 78512
rect 141620 78508 141626 78510
rect 139577 78507 139643 78508
rect 141877 78507 141943 78510
rect 142797 78570 142863 78573
rect 144870 78570 144930 78646
rect 580901 78643 580967 78646
rect 142797 78568 144930 78570
rect 142797 78512 142802 78568
rect 142858 78512 144930 78568
rect 142797 78510 144930 78512
rect 154573 78572 154639 78573
rect 154573 78568 154620 78572
rect 154684 78570 154690 78572
rect 154849 78570 154915 78573
rect 154982 78570 154988 78572
rect 154573 78512 154578 78568
rect 142797 78507 142863 78510
rect 154573 78508 154620 78512
rect 154684 78510 154730 78570
rect 154849 78568 154988 78570
rect 154849 78512 154854 78568
rect 154910 78512 154988 78568
rect 154849 78510 154988 78512
rect 154684 78508 154690 78510
rect 154573 78507 154639 78508
rect 154849 78507 154915 78510
rect 154982 78508 154988 78510
rect 155052 78508 155058 78572
rect 161749 78570 161815 78573
rect 172421 78572 172487 78573
rect 162710 78570 162716 78572
rect 161749 78568 162716 78570
rect 161749 78512 161754 78568
rect 161810 78512 162716 78568
rect 161749 78510 162716 78512
rect 161749 78507 161815 78510
rect 162710 78508 162716 78510
rect 162780 78508 162786 78572
rect 172421 78570 172468 78572
rect 172376 78568 172468 78570
rect 172376 78512 172426 78568
rect 172376 78510 172468 78512
rect 172421 78508 172468 78510
rect 172532 78508 172538 78572
rect 172605 78570 172671 78573
rect 175917 78572 175983 78573
rect 172830 78570 172836 78572
rect 172605 78568 172836 78570
rect 172605 78512 172610 78568
rect 172666 78512 172836 78568
rect 172605 78510 172836 78512
rect 172421 78507 172487 78508
rect 172605 78507 172671 78510
rect 172830 78508 172836 78510
rect 172900 78508 172906 78572
rect 175917 78570 175964 78572
rect 175872 78568 175964 78570
rect 175872 78512 175922 78568
rect 175872 78510 175964 78512
rect 175917 78508 175964 78510
rect 176028 78508 176034 78572
rect 176326 78508 176332 78572
rect 176396 78570 176402 78572
rect 176469 78570 176535 78573
rect 176396 78568 176535 78570
rect 176396 78512 176474 78568
rect 176530 78512 176535 78568
rect 176396 78510 176535 78512
rect 176396 78508 176402 78510
rect 175917 78507 175983 78508
rect 176469 78507 176535 78510
rect 101990 78372 101996 78436
rect 102060 78434 102066 78436
rect 132861 78434 132927 78437
rect 102060 78432 132927 78434
rect 102060 78376 132866 78432
rect 132922 78376 132927 78432
rect 102060 78374 132927 78376
rect 102060 78372 102066 78374
rect 132861 78371 132927 78374
rect 133086 78372 133092 78436
rect 133156 78434 133162 78436
rect 141417 78434 141483 78437
rect 133156 78432 141483 78434
rect 133156 78376 141422 78432
rect 141478 78376 141483 78432
rect 133156 78374 141483 78376
rect 133156 78372 133162 78374
rect 141417 78371 141483 78374
rect 166073 78434 166139 78437
rect 169150 78434 169156 78436
rect 166073 78432 169156 78434
rect 166073 78376 166078 78432
rect 166134 78376 169156 78432
rect 166073 78374 169156 78376
rect 166073 78371 166139 78374
rect 169150 78372 169156 78374
rect 169220 78372 169226 78436
rect 170673 78434 170739 78437
rect 171726 78434 171732 78436
rect 170673 78432 171732 78434
rect 170673 78376 170678 78432
rect 170734 78376 171732 78432
rect 170673 78374 171732 78376
rect 170673 78371 170739 78374
rect 171726 78372 171732 78374
rect 171796 78372 171802 78436
rect 173249 78434 173315 78437
rect 207197 78434 207263 78437
rect 173249 78432 207263 78434
rect 173249 78376 173254 78432
rect 173310 78376 207202 78432
rect 207258 78376 207263 78432
rect 173249 78374 207263 78376
rect 173249 78371 173315 78374
rect 207197 78371 207263 78374
rect 103278 78236 103284 78300
rect 103348 78298 103354 78300
rect 129181 78298 129247 78301
rect 103348 78296 129247 78298
rect 103348 78240 129186 78296
rect 129242 78240 129247 78296
rect 103348 78238 129247 78240
rect 103348 78236 103354 78238
rect 129181 78235 129247 78238
rect 135110 78236 135116 78300
rect 135180 78298 135186 78300
rect 136766 78298 136772 78300
rect 135180 78238 136772 78298
rect 135180 78236 135186 78238
rect 136766 78236 136772 78238
rect 136836 78236 136842 78300
rect 139117 78298 139183 78301
rect 141918 78298 141924 78300
rect 139117 78296 141924 78298
rect 139117 78240 139122 78296
rect 139178 78240 141924 78296
rect 139117 78238 141924 78240
rect 139117 78235 139183 78238
rect 141918 78236 141924 78238
rect 141988 78236 141994 78300
rect 170857 78298 170923 78301
rect 181621 78298 181687 78301
rect 211102 78298 211108 78300
rect 170857 78296 176670 78298
rect 170857 78240 170862 78296
rect 170918 78240 176670 78296
rect 170857 78238 176670 78240
rect 170857 78235 170923 78238
rect 123886 78100 123892 78164
rect 123956 78162 123962 78164
rect 135713 78162 135779 78165
rect 123956 78160 135779 78162
rect 123956 78104 135718 78160
rect 135774 78104 135779 78160
rect 123956 78102 135779 78104
rect 123956 78100 123962 78102
rect 135713 78099 135779 78102
rect 136582 78100 136588 78164
rect 136652 78162 136658 78164
rect 145833 78162 145899 78165
rect 136652 78160 145899 78162
rect 136652 78104 145838 78160
rect 145894 78104 145899 78160
rect 136652 78102 145899 78104
rect 176610 78162 176670 78238
rect 181621 78296 211108 78298
rect 181621 78240 181626 78296
rect 181682 78240 211108 78296
rect 181621 78238 211108 78240
rect 181621 78235 181687 78238
rect 211102 78236 211108 78238
rect 211172 78236 211178 78300
rect 187734 78162 187740 78164
rect 176610 78102 187740 78162
rect 136652 78100 136658 78102
rect 145833 78099 145899 78102
rect 187734 78100 187740 78102
rect 187804 78100 187810 78164
rect 126329 78026 126395 78029
rect 122790 78024 126395 78026
rect 122790 77968 126334 78024
rect 126390 77968 126395 78024
rect 122790 77966 126395 77968
rect 104750 77828 104756 77892
rect 104820 77890 104826 77892
rect 122790 77890 122850 77966
rect 126329 77963 126395 77966
rect 134977 78026 135043 78029
rect 138105 78028 138171 78029
rect 136398 78026 136404 78028
rect 134977 78024 136404 78026
rect 134977 77968 134982 78024
rect 135038 77968 136404 78024
rect 134977 77966 136404 77968
rect 134977 77963 135043 77966
rect 136398 77964 136404 77966
rect 136468 77964 136474 78028
rect 138054 78026 138060 78028
rect 138014 77966 138060 78026
rect 138124 78024 138171 78028
rect 138166 77968 138171 78024
rect 138054 77964 138060 77966
rect 138124 77964 138171 77968
rect 140630 77964 140636 78028
rect 140700 78026 140706 78028
rect 149605 78026 149671 78029
rect 140700 78024 149671 78026
rect 140700 77968 149610 78024
rect 149666 77968 149671 78024
rect 140700 77966 149671 77968
rect 140700 77964 140706 77966
rect 138105 77963 138171 77964
rect 149605 77963 149671 77966
rect 152825 78026 152891 78029
rect 161422 78026 161428 78028
rect 152825 78024 161428 78026
rect 152825 77968 152830 78024
rect 152886 77968 161428 78024
rect 152825 77966 161428 77968
rect 152825 77963 152891 77966
rect 161422 77964 161428 77966
rect 161492 77964 161498 78028
rect 170949 78026 171015 78029
rect 180701 78026 180767 78029
rect 195329 78026 195395 78029
rect 170949 78024 179430 78026
rect 170949 77968 170954 78024
rect 171010 77968 179430 78024
rect 170949 77966 179430 77968
rect 170949 77963 171015 77966
rect 135253 77890 135319 77893
rect 104820 77830 122850 77890
rect 128310 77888 135319 77890
rect 128310 77832 135258 77888
rect 135314 77832 135319 77888
rect 128310 77830 135319 77832
rect 104820 77828 104826 77830
rect 97758 77556 97764 77620
rect 97828 77618 97834 77620
rect 128310 77618 128370 77830
rect 135253 77827 135319 77830
rect 142654 77828 142660 77892
rect 142724 77890 142730 77892
rect 151537 77890 151603 77893
rect 142724 77888 151603 77890
rect 142724 77832 151542 77888
rect 151598 77832 151603 77888
rect 142724 77830 151603 77832
rect 142724 77828 142730 77830
rect 151537 77827 151603 77830
rect 152958 77828 152964 77892
rect 153028 77890 153034 77892
rect 155493 77890 155559 77893
rect 173709 77892 173775 77893
rect 153028 77888 155559 77890
rect 153028 77832 155498 77888
rect 155554 77832 155559 77888
rect 153028 77830 155559 77832
rect 153028 77828 153034 77830
rect 155493 77827 155559 77830
rect 158478 77828 158484 77892
rect 158548 77890 158554 77892
rect 173709 77890 173756 77892
rect 158548 77830 159098 77890
rect 173664 77888 173756 77890
rect 173664 77832 173714 77888
rect 173664 77830 173756 77832
rect 158548 77828 158554 77830
rect 141325 77754 141391 77757
rect 97828 77558 128370 77618
rect 133094 77752 141391 77754
rect 133094 77696 141330 77752
rect 141386 77696 141391 77752
rect 133094 77694 141391 77696
rect 97828 77556 97834 77558
rect 121310 77420 121316 77484
rect 121380 77482 121386 77484
rect 133094 77482 133154 77694
rect 141325 77691 141391 77694
rect 142061 77754 142127 77757
rect 148174 77754 148180 77756
rect 142061 77752 148180 77754
rect 142061 77696 142066 77752
rect 142122 77696 148180 77752
rect 142061 77694 148180 77696
rect 142061 77691 142127 77694
rect 148174 77692 148180 77694
rect 148244 77692 148250 77756
rect 149973 77754 150039 77757
rect 158621 77754 158687 77757
rect 149973 77752 158687 77754
rect 149973 77696 149978 77752
rect 150034 77696 158626 77752
rect 158682 77696 158687 77752
rect 149973 77694 158687 77696
rect 159038 77754 159098 77830
rect 173709 77828 173756 77830
rect 173820 77828 173826 77892
rect 175549 77890 175615 77893
rect 176510 77890 176516 77892
rect 175549 77888 176516 77890
rect 175549 77832 175554 77888
rect 175610 77832 176516 77888
rect 175549 77830 176516 77832
rect 173709 77827 173775 77828
rect 175549 77827 175615 77830
rect 176510 77828 176516 77830
rect 176580 77828 176586 77892
rect 172462 77754 172468 77756
rect 159038 77694 172468 77754
rect 149973 77691 150039 77694
rect 158621 77691 158687 77694
rect 172462 77692 172468 77694
rect 172532 77692 172538 77756
rect 179370 77754 179430 77966
rect 180701 78024 195395 78026
rect 180701 77968 180706 78024
rect 180762 77968 195334 78024
rect 195390 77968 195395 78024
rect 180701 77966 195395 77968
rect 180701 77963 180767 77966
rect 195329 77963 195395 77966
rect 182909 77890 182975 77893
rect 209957 77890 210023 77893
rect 182909 77888 210023 77890
rect 182909 77832 182914 77888
rect 182970 77832 209962 77888
rect 210018 77832 210023 77888
rect 182909 77830 210023 77832
rect 182909 77827 182975 77830
rect 209957 77827 210023 77830
rect 188981 77754 189047 77757
rect 179370 77752 189047 77754
rect 179370 77696 188986 77752
rect 189042 77696 189047 77752
rect 179370 77694 189047 77696
rect 188981 77691 189047 77694
rect 150157 77618 150223 77621
rect 140638 77616 150223 77618
rect 140638 77560 150162 77616
rect 150218 77560 150223 77616
rect 140638 77558 150223 77560
rect 121380 77422 133154 77482
rect 121380 77420 121386 77422
rect 140446 77420 140452 77484
rect 140516 77482 140522 77484
rect 140638 77482 140698 77558
rect 150157 77555 150223 77558
rect 140516 77422 140698 77482
rect 140516 77420 140522 77422
rect 160870 77420 160876 77484
rect 160940 77482 160946 77484
rect 160940 77422 176670 77482
rect 160940 77420 160946 77422
rect 135846 77284 135852 77348
rect 135916 77346 135922 77348
rect 137185 77346 137251 77349
rect 135916 77344 137251 77346
rect 135916 77288 137190 77344
rect 137246 77288 137251 77344
rect 135916 77286 137251 77288
rect 176610 77346 176670 77422
rect 214741 77346 214807 77349
rect 176610 77344 214807 77346
rect 176610 77288 214746 77344
rect 214802 77288 214807 77344
rect 176610 77286 214807 77288
rect 135916 77284 135922 77286
rect 137185 77283 137251 77286
rect 214741 77283 214807 77286
rect 104382 77148 104388 77212
rect 104452 77210 104458 77212
rect 104525 77210 104591 77213
rect 104452 77208 104591 77210
rect 104452 77152 104530 77208
rect 104586 77152 104591 77208
rect 104452 77150 104591 77152
rect 104452 77148 104458 77150
rect 104525 77147 104591 77150
rect 135294 77148 135300 77212
rect 135364 77210 135370 77212
rect 140497 77210 140563 77213
rect 135364 77208 140563 77210
rect 135364 77152 140502 77208
rect 140558 77152 140563 77208
rect 135364 77150 140563 77152
rect 135364 77148 135370 77150
rect 140497 77147 140563 77150
rect 160645 77210 160711 77213
rect 180701 77210 180767 77213
rect 160645 77208 180767 77210
rect 160645 77152 160650 77208
rect 160706 77152 180706 77208
rect 180762 77152 180767 77208
rect 160645 77150 180767 77152
rect 160645 77147 160711 77150
rect 180701 77147 180767 77150
rect 181437 77210 181503 77213
rect 193581 77210 193647 77213
rect 194501 77210 194567 77213
rect 181437 77208 194567 77210
rect 181437 77152 181442 77208
rect 181498 77152 193586 77208
rect 193642 77152 194506 77208
rect 194562 77152 194567 77208
rect 181437 77150 194567 77152
rect 181437 77147 181503 77150
rect 193581 77147 193647 77150
rect 194501 77147 194567 77150
rect 104566 77012 104572 77076
rect 104636 77074 104642 77076
rect 138657 77074 138723 77077
rect 104636 77072 138723 77074
rect 104636 77016 138662 77072
rect 138718 77016 138723 77072
rect 104636 77014 138723 77016
rect 104636 77012 104642 77014
rect 138657 77011 138723 77014
rect 164734 77012 164740 77076
rect 164804 77074 164810 77076
rect 170622 77074 170628 77076
rect 164804 77014 170628 77074
rect 164804 77012 164810 77014
rect 170622 77012 170628 77014
rect 170692 77012 170698 77076
rect 180609 77074 180675 77077
rect 220905 77074 220971 77077
rect 180609 77072 220971 77074
rect 180609 77016 180614 77072
rect 180670 77016 220910 77072
rect 220966 77016 220971 77072
rect 180609 77014 220971 77016
rect 180609 77011 180675 77014
rect 220905 77011 220971 77014
rect 108798 76876 108804 76940
rect 108868 76938 108874 76940
rect 136633 76938 136699 76941
rect 108868 76936 136699 76938
rect 108868 76880 136638 76936
rect 136694 76880 136699 76936
rect 108868 76878 136699 76880
rect 108868 76876 108874 76878
rect 136633 76875 136699 76878
rect 167913 76938 167979 76941
rect 180333 76938 180399 76941
rect 167913 76936 180399 76938
rect 167913 76880 167918 76936
rect 167974 76880 180338 76936
rect 180394 76880 180399 76936
rect 167913 76878 180399 76880
rect 167913 76875 167979 76878
rect 180333 76875 180399 76878
rect 580441 76938 580507 76941
rect 583520 76938 584960 77028
rect 580441 76936 584960 76938
rect 580441 76880 580446 76936
rect 580502 76880 584960 76936
rect 580441 76878 584960 76880
rect 580441 76875 580507 76878
rect 113766 76740 113772 76804
rect 113836 76802 113842 76804
rect 137001 76802 137067 76805
rect 113836 76800 137067 76802
rect 113836 76744 137006 76800
rect 137062 76744 137067 76800
rect 113836 76742 137067 76744
rect 113836 76740 113842 76742
rect 137001 76739 137067 76742
rect 161013 76802 161079 76805
rect 169017 76802 169083 76805
rect 161013 76800 169083 76802
rect 161013 76744 161018 76800
rect 161074 76744 169022 76800
rect 169078 76744 169083 76800
rect 161013 76742 169083 76744
rect 161013 76739 161079 76742
rect 169017 76739 169083 76742
rect 169385 76802 169451 76805
rect 203190 76802 203196 76804
rect 169385 76800 203196 76802
rect 169385 76744 169390 76800
rect 169446 76744 203196 76800
rect 169385 76742 203196 76744
rect 169385 76739 169451 76742
rect 203190 76740 203196 76742
rect 203260 76740 203266 76804
rect 583520 76788 584960 76878
rect 116894 76604 116900 76668
rect 116964 76666 116970 76668
rect 140630 76666 140636 76668
rect 116964 76606 140636 76666
rect 116964 76604 116970 76606
rect 140630 76604 140636 76606
rect 140700 76604 140706 76668
rect 140814 76604 140820 76668
rect 140884 76666 140890 76668
rect 141141 76666 141207 76669
rect 140884 76664 141207 76666
rect 140884 76608 141146 76664
rect 141202 76608 141207 76664
rect 140884 76606 141207 76608
rect 140884 76604 140890 76606
rect 141141 76603 141207 76606
rect 141417 76666 141483 76669
rect 144821 76668 144887 76669
rect 143942 76666 143948 76668
rect 141417 76664 143948 76666
rect 141417 76608 141422 76664
rect 141478 76608 143948 76664
rect 141417 76606 143948 76608
rect 141417 76603 141483 76606
rect 143942 76604 143948 76606
rect 144012 76604 144018 76668
rect 144821 76666 144868 76668
rect 144776 76664 144868 76666
rect 144776 76608 144826 76664
rect 144776 76606 144868 76608
rect 144821 76604 144868 76606
rect 144932 76604 144938 76668
rect 146477 76666 146543 76669
rect 146702 76666 146708 76668
rect 146477 76664 146708 76666
rect 146477 76608 146482 76664
rect 146538 76608 146708 76664
rect 146477 76606 146708 76608
rect 144821 76603 144887 76604
rect 146477 76603 146543 76606
rect 146702 76604 146708 76606
rect 146772 76604 146778 76668
rect 156137 76666 156203 76669
rect 156454 76666 156460 76668
rect 156137 76664 156460 76666
rect 156137 76608 156142 76664
rect 156198 76608 156460 76664
rect 156137 76606 156460 76608
rect 156137 76603 156203 76606
rect 156454 76604 156460 76606
rect 156524 76604 156530 76668
rect 162526 76604 162532 76668
rect 162596 76666 162602 76668
rect 170254 76666 170260 76668
rect 162596 76606 170260 76666
rect 162596 76604 162602 76606
rect 170254 76604 170260 76606
rect 170324 76604 170330 76668
rect 173985 76666 174051 76669
rect 200982 76666 200988 76668
rect 173985 76664 200988 76666
rect 173985 76608 173990 76664
rect 174046 76608 200988 76664
rect 173985 76606 200988 76608
rect 173985 76603 174051 76606
rect 200982 76604 200988 76606
rect 201052 76604 201058 76668
rect 95141 76530 95207 76533
rect 135069 76530 135135 76533
rect 95141 76528 135135 76530
rect 95141 76472 95146 76528
rect 95202 76472 135074 76528
rect 135130 76472 135135 76528
rect 95141 76470 135135 76472
rect 95141 76467 95207 76470
rect 135069 76467 135135 76470
rect 138381 76532 138447 76533
rect 138381 76528 138428 76532
rect 138492 76530 138498 76532
rect 172421 76530 172487 76533
rect 214465 76530 214531 76533
rect 138381 76472 138386 76528
rect 138381 76468 138428 76472
rect 138492 76470 138538 76530
rect 172421 76528 214531 76530
rect 172421 76472 172426 76528
rect 172482 76472 214470 76528
rect 214526 76472 214531 76528
rect 172421 76470 214531 76472
rect 138492 76468 138498 76470
rect 138381 76467 138447 76468
rect 172421 76467 172487 76470
rect 214465 76467 214531 76470
rect -960 76258 480 76348
rect 129774 76332 129780 76396
rect 129844 76394 129850 76396
rect 151077 76394 151143 76397
rect 129844 76392 151143 76394
rect 129844 76336 151082 76392
rect 151138 76336 151143 76392
rect 129844 76334 151143 76336
rect 129844 76332 129850 76334
rect 151077 76331 151143 76334
rect 156229 76394 156295 76397
rect 190494 76394 190500 76396
rect 156229 76392 190500 76394
rect 156229 76336 156234 76392
rect 156290 76336 190500 76392
rect 156229 76334 190500 76336
rect 156229 76331 156295 76334
rect 190494 76332 190500 76334
rect 190564 76332 190570 76396
rect 2865 76258 2931 76261
rect -960 76256 2931 76258
rect -960 76200 2870 76256
rect 2926 76200 2931 76256
rect -960 76198 2931 76200
rect -960 76108 480 76198
rect 2865 76195 2931 76198
rect 134006 76196 134012 76260
rect 134076 76258 134082 76260
rect 135529 76258 135595 76261
rect 134076 76256 135595 76258
rect 134076 76200 135534 76256
rect 135590 76200 135595 76256
rect 134076 76198 135595 76200
rect 134076 76196 134082 76198
rect 135529 76195 135595 76198
rect 176009 76258 176075 76261
rect 215569 76258 215635 76261
rect 176009 76256 215635 76258
rect 176009 76200 176014 76256
rect 176070 76200 215574 76256
rect 215630 76200 215635 76256
rect 176009 76198 215635 76200
rect 176009 76195 176075 76198
rect 215569 76195 215635 76198
rect 152457 75986 152523 75989
rect 152958 75986 152964 75988
rect 152457 75984 152964 75986
rect 152457 75928 152462 75984
rect 152518 75928 152964 75984
rect 152457 75926 152964 75928
rect 152457 75923 152523 75926
rect 152958 75924 152964 75926
rect 153028 75924 153034 75988
rect 154246 75924 154252 75988
rect 154316 75986 154322 75988
rect 154665 75986 154731 75989
rect 154316 75984 154731 75986
rect 154316 75928 154670 75984
rect 154726 75928 154731 75984
rect 154316 75926 154731 75928
rect 154316 75924 154322 75926
rect 154665 75923 154731 75926
rect 155309 75986 155375 75989
rect 157926 75986 157932 75988
rect 155309 75984 157932 75986
rect 155309 75928 155314 75984
rect 155370 75928 157932 75984
rect 155309 75926 157932 75928
rect 155309 75923 155375 75926
rect 157926 75924 157932 75926
rect 157996 75924 158002 75988
rect 169753 75986 169819 75989
rect 170438 75986 170444 75988
rect 169753 75984 170444 75986
rect 169753 75928 169758 75984
rect 169814 75928 170444 75984
rect 169753 75926 170444 75928
rect 169753 75923 169819 75926
rect 170438 75924 170444 75926
rect 170508 75924 170514 75988
rect 104709 75850 104775 75853
rect 145281 75850 145347 75853
rect 104709 75848 145347 75850
rect 104709 75792 104714 75848
rect 104770 75792 145286 75848
rect 145342 75792 145347 75848
rect 104709 75790 145347 75792
rect 104709 75787 104775 75790
rect 145281 75787 145347 75790
rect 153837 75850 153903 75853
rect 154430 75850 154436 75852
rect 153837 75848 154436 75850
rect 153837 75792 153842 75848
rect 153898 75792 154436 75848
rect 153837 75790 154436 75792
rect 153837 75787 153903 75790
rect 154430 75788 154436 75790
rect 154500 75788 154506 75852
rect 169661 75850 169727 75853
rect 192150 75850 192156 75852
rect 169661 75848 192156 75850
rect 169661 75792 169666 75848
rect 169722 75792 192156 75848
rect 169661 75790 192156 75792
rect 169661 75787 169727 75790
rect 192150 75788 192156 75790
rect 192220 75788 192226 75852
rect 113950 75652 113956 75716
rect 114020 75714 114026 75716
rect 146518 75714 146524 75716
rect 114020 75654 146524 75714
rect 114020 75652 114026 75654
rect 146518 75652 146524 75654
rect 146588 75652 146594 75716
rect 161422 75652 161428 75716
rect 161492 75714 161498 75716
rect 219801 75714 219867 75717
rect 161492 75712 219867 75714
rect 161492 75656 219806 75712
rect 219862 75656 219867 75712
rect 161492 75654 219867 75656
rect 161492 75652 161498 75654
rect 219801 75651 219867 75654
rect 114134 75516 114140 75580
rect 114204 75578 114210 75580
rect 147397 75578 147463 75581
rect 114204 75576 147463 75578
rect 114204 75520 147402 75576
rect 147458 75520 147463 75576
rect 114204 75518 147463 75520
rect 114204 75516 114210 75518
rect 147397 75515 147463 75518
rect 161606 75516 161612 75580
rect 161676 75578 161682 75580
rect 212901 75578 212967 75581
rect 161676 75576 212967 75578
rect 161676 75520 212906 75576
rect 212962 75520 212967 75576
rect 161676 75518 212967 75520
rect 161676 75516 161682 75518
rect 212901 75515 212967 75518
rect 109861 75442 109927 75445
rect 143165 75442 143231 75445
rect 109861 75440 143231 75442
rect 109861 75384 109866 75440
rect 109922 75384 143170 75440
rect 143226 75384 143231 75440
rect 109861 75382 143231 75384
rect 109861 75379 109927 75382
rect 143165 75379 143231 75382
rect 151997 75442 152063 75445
rect 201534 75442 201540 75444
rect 151997 75440 201540 75442
rect 151997 75384 152002 75440
rect 152058 75384 201540 75440
rect 151997 75382 201540 75384
rect 151997 75379 152063 75382
rect 201534 75380 201540 75382
rect 201604 75380 201610 75444
rect 102910 75244 102916 75308
rect 102980 75306 102986 75308
rect 137093 75306 137159 75309
rect 102980 75304 137159 75306
rect 102980 75248 137098 75304
rect 137154 75248 137159 75304
rect 102980 75246 137159 75248
rect 102980 75244 102986 75246
rect 137093 75243 137159 75246
rect 162761 75306 162827 75309
rect 186998 75306 187004 75308
rect 162761 75304 187004 75306
rect 162761 75248 162766 75304
rect 162822 75248 187004 75304
rect 162761 75246 187004 75248
rect 162761 75243 162827 75246
rect 186998 75244 187004 75246
rect 187068 75244 187074 75308
rect 133321 75170 133387 75173
rect 133638 75170 133644 75172
rect 133321 75168 133644 75170
rect 133321 75112 133326 75168
rect 133382 75112 133644 75168
rect 133321 75110 133644 75112
rect 133321 75107 133387 75110
rect 133638 75108 133644 75110
rect 133708 75108 133714 75172
rect 145281 75170 145347 75173
rect 534073 75170 534139 75173
rect 145281 75168 534139 75170
rect 145281 75112 145286 75168
rect 145342 75112 534078 75168
rect 534134 75112 534139 75168
rect 145281 75110 534139 75112
rect 145281 75107 145347 75110
rect 534073 75107 534139 75110
rect 118182 74972 118188 75036
rect 118252 75034 118258 75036
rect 149789 75034 149855 75037
rect 118252 75032 149855 75034
rect 118252 74976 149794 75032
rect 149850 74976 149855 75032
rect 118252 74974 149855 74976
rect 118252 74972 118258 74974
rect 149789 74971 149855 74974
rect 159817 75034 159883 75037
rect 166206 75034 166212 75036
rect 159817 75032 166212 75034
rect 159817 74976 159822 75032
rect 159878 74976 166212 75032
rect 159817 74974 166212 74976
rect 159817 74971 159883 74974
rect 166206 74972 166212 74974
rect 166276 74972 166282 75036
rect 176326 74972 176332 75036
rect 176396 75034 176402 75036
rect 176561 75034 176627 75037
rect 176396 75032 176627 75034
rect 176396 74976 176566 75032
rect 176622 74976 176627 75032
rect 176396 74974 176627 74976
rect 176396 74972 176402 74974
rect 176561 74971 176627 74974
rect 119245 74898 119311 74901
rect 147070 74898 147076 74900
rect 119245 74896 147076 74898
rect 119245 74840 119250 74896
rect 119306 74840 147076 74896
rect 119245 74838 147076 74840
rect 119245 74835 119311 74838
rect 147070 74836 147076 74838
rect 147140 74836 147146 74900
rect 148726 74836 148732 74900
rect 148796 74898 148802 74900
rect 216673 74898 216739 74901
rect 148796 74896 216739 74898
rect 148796 74840 216678 74896
rect 216734 74840 216739 74896
rect 148796 74838 216739 74840
rect 148796 74836 148802 74838
rect 216673 74835 216739 74838
rect 122373 74490 122439 74493
rect 147673 74490 147739 74493
rect 122373 74488 147739 74490
rect 122373 74432 122378 74488
rect 122434 74432 147678 74488
rect 147734 74432 147739 74488
rect 122373 74430 147739 74432
rect 122373 74427 122439 74430
rect 147673 74427 147739 74430
rect 170622 74428 170628 74492
rect 170692 74490 170698 74492
rect 197486 74490 197492 74492
rect 170692 74430 197492 74490
rect 170692 74428 170698 74430
rect 197486 74428 197492 74430
rect 197556 74428 197562 74492
rect 111374 74292 111380 74356
rect 111444 74354 111450 74356
rect 144177 74354 144243 74357
rect 111444 74352 144243 74354
rect 111444 74296 144182 74352
rect 144238 74296 144243 74352
rect 111444 74294 144243 74296
rect 111444 74292 111450 74294
rect 144177 74291 144243 74294
rect 161473 74354 161539 74357
rect 194542 74354 194548 74356
rect 161473 74352 194548 74354
rect 161473 74296 161478 74352
rect 161534 74296 194548 74352
rect 161473 74294 194548 74296
rect 161473 74291 161539 74294
rect 194542 74292 194548 74294
rect 194612 74292 194618 74356
rect 119654 74156 119660 74220
rect 119724 74218 119730 74220
rect 153653 74218 153719 74221
rect 119724 74216 153719 74218
rect 119724 74160 153658 74216
rect 153714 74160 153719 74216
rect 119724 74158 153719 74160
rect 119724 74156 119730 74158
rect 153653 74155 153719 74158
rect 178309 74218 178375 74221
rect 208853 74218 208919 74221
rect 178309 74216 208919 74218
rect 178309 74160 178314 74216
rect 178370 74160 208858 74216
rect 208914 74160 208919 74216
rect 178309 74158 208919 74160
rect 178309 74155 178375 74158
rect 208853 74155 208919 74158
rect 103094 74020 103100 74084
rect 103164 74082 103170 74084
rect 135110 74082 135116 74084
rect 103164 74022 135116 74082
rect 103164 74020 103170 74022
rect 135110 74020 135116 74022
rect 135180 74020 135186 74084
rect 166165 74082 166231 74085
rect 200113 74082 200179 74085
rect 166165 74080 200179 74082
rect 166165 74024 166170 74080
rect 166226 74024 200118 74080
rect 200174 74024 200179 74080
rect 166165 74022 200179 74024
rect 166165 74019 166231 74022
rect 200113 74019 200179 74022
rect 207013 74082 207079 74085
rect 207606 74082 207612 74084
rect 207013 74080 207612 74082
rect 207013 74024 207018 74080
rect 207074 74024 207612 74080
rect 207013 74022 207612 74024
rect 207013 74019 207079 74022
rect 207606 74020 207612 74022
rect 207676 74020 207682 74084
rect 116710 73884 116716 73948
rect 116780 73946 116786 73948
rect 146937 73946 147003 73949
rect 153929 73946 153995 73949
rect 116780 73944 153995 73946
rect 116780 73888 146942 73944
rect 146998 73888 153934 73944
rect 153990 73888 153995 73944
rect 116780 73886 153995 73888
rect 116780 73884 116786 73886
rect 146937 73883 147003 73886
rect 153929 73883 153995 73886
rect 164141 73946 164207 73949
rect 193673 73946 193739 73949
rect 164141 73944 193739 73946
rect 164141 73888 164146 73944
rect 164202 73888 193678 73944
rect 193734 73888 193739 73944
rect 164141 73886 193739 73888
rect 164141 73883 164207 73886
rect 193673 73883 193739 73886
rect 117078 73748 117084 73812
rect 117148 73810 117154 73812
rect 140037 73810 140103 73813
rect 117148 73808 140103 73810
rect 117148 73752 140042 73808
rect 140098 73752 140103 73808
rect 117148 73750 140103 73752
rect 117148 73748 117154 73750
rect 140037 73747 140103 73750
rect 166165 73810 166231 73813
rect 166574 73810 166580 73812
rect 166165 73808 166580 73810
rect 166165 73752 166170 73808
rect 166226 73752 166580 73808
rect 166165 73750 166580 73752
rect 166165 73747 166231 73750
rect 166574 73748 166580 73750
rect 166644 73748 166650 73812
rect 170254 73748 170260 73812
rect 170324 73810 170330 73812
rect 196566 73810 196572 73812
rect 170324 73750 196572 73810
rect 170324 73748 170330 73750
rect 196566 73748 196572 73750
rect 196636 73748 196642 73812
rect 118366 73612 118372 73676
rect 118436 73674 118442 73676
rect 151445 73674 151511 73677
rect 118436 73672 151511 73674
rect 118436 73616 151450 73672
rect 151506 73616 151511 73672
rect 118436 73614 151511 73616
rect 118436 73612 118442 73614
rect 151445 73611 151511 73614
rect 160461 73674 160527 73677
rect 193254 73674 193260 73676
rect 160461 73672 193260 73674
rect 160461 73616 160466 73672
rect 160522 73616 193260 73672
rect 160461 73614 193260 73616
rect 160461 73611 160527 73614
rect 193254 73612 193260 73614
rect 193324 73612 193330 73676
rect 118550 73068 118556 73132
rect 118620 73130 118626 73132
rect 140446 73130 140452 73132
rect 118620 73070 140452 73130
rect 118620 73068 118626 73070
rect 140446 73068 140452 73070
rect 140516 73068 140522 73132
rect 172462 73068 172468 73132
rect 172532 73130 172538 73132
rect 187049 73130 187115 73133
rect 172532 73128 187115 73130
rect 172532 73072 187054 73128
rect 187110 73072 187115 73128
rect 172532 73070 187115 73072
rect 172532 73068 172538 73070
rect 187049 73067 187115 73070
rect 112846 72932 112852 72996
rect 112916 72994 112922 72996
rect 146702 72994 146708 72996
rect 112916 72934 146708 72994
rect 112916 72932 112922 72934
rect 146702 72932 146708 72934
rect 146772 72932 146778 72996
rect 162761 72994 162827 72997
rect 196382 72994 196388 72996
rect 162761 72992 196388 72994
rect 162761 72936 162766 72992
rect 162822 72936 196388 72992
rect 162761 72934 196388 72936
rect 162761 72931 162827 72934
rect 196382 72932 196388 72934
rect 196452 72932 196458 72996
rect 119797 72858 119863 72861
rect 152038 72858 152044 72860
rect 119797 72856 152044 72858
rect 119797 72800 119802 72856
rect 119858 72800 152044 72856
rect 119797 72798 152044 72800
rect 119797 72795 119863 72798
rect 152038 72796 152044 72798
rect 152108 72796 152114 72860
rect 163865 72858 163931 72861
rect 197302 72858 197308 72860
rect 163865 72856 197308 72858
rect 163865 72800 163870 72856
rect 163926 72800 197308 72856
rect 163865 72798 197308 72800
rect 163865 72795 163931 72798
rect 197302 72796 197308 72798
rect 197372 72796 197378 72860
rect 580165 72858 580231 72861
rect 583520 72858 584960 72948
rect 580165 72856 584960 72858
rect 580165 72800 580170 72856
rect 580226 72800 584960 72856
rect 580165 72798 584960 72800
rect 580165 72795 580231 72798
rect 115790 72660 115796 72724
rect 115860 72722 115866 72724
rect 143993 72722 144059 72725
rect 115860 72720 144059 72722
rect 115860 72664 143998 72720
rect 144054 72664 144059 72720
rect 115860 72662 144059 72664
rect 115860 72660 115866 72662
rect 143993 72659 144059 72662
rect 164877 72722 164943 72725
rect 198774 72722 198780 72724
rect 164877 72720 198780 72722
rect 164877 72664 164882 72720
rect 164938 72664 198780 72720
rect 164877 72662 198780 72664
rect 164877 72659 164943 72662
rect 198774 72660 198780 72662
rect 198844 72660 198850 72724
rect 583520 72708 584960 72798
rect 112437 72586 112503 72589
rect 136582 72586 136588 72588
rect 112437 72584 136588 72586
rect 112437 72528 112442 72584
rect 112498 72528 136588 72584
rect 112437 72526 136588 72528
rect 112437 72523 112503 72526
rect 136582 72524 136588 72526
rect 136652 72524 136658 72588
rect 170857 72586 170923 72589
rect 196065 72586 196131 72589
rect 170857 72584 196131 72586
rect 170857 72528 170862 72584
rect 170918 72528 196070 72584
rect 196126 72528 196131 72584
rect 170857 72526 196131 72528
rect 170857 72523 170923 72526
rect 196065 72523 196131 72526
rect 112713 72450 112779 72453
rect 147990 72450 147996 72452
rect 112713 72448 147996 72450
rect 112713 72392 112718 72448
rect 112774 72392 147996 72448
rect 112713 72390 147996 72392
rect 112713 72387 112779 72390
rect 147990 72388 147996 72390
rect 148060 72388 148066 72452
rect 165337 72450 165403 72453
rect 199326 72450 199332 72452
rect 165337 72448 199332 72450
rect 165337 72392 165342 72448
rect 165398 72392 199332 72448
rect 165337 72390 199332 72392
rect 165337 72387 165403 72390
rect 199326 72388 199332 72390
rect 199396 72388 199402 72452
rect -960 72178 480 72268
rect 3141 72178 3207 72181
rect -960 72176 3207 72178
rect -960 72120 3146 72176
rect 3202 72120 3207 72176
rect -960 72118 3207 72120
rect -960 72028 480 72118
rect 3141 72115 3207 72118
rect 97073 71770 97139 71773
rect 146293 71770 146359 71773
rect 97073 71768 146359 71770
rect 97073 71712 97078 71768
rect 97134 71712 146298 71768
rect 146354 71712 146359 71768
rect 97073 71710 146359 71712
rect 97073 71707 97139 71710
rect 146293 71707 146359 71710
rect 155534 71708 155540 71772
rect 155604 71770 155610 71772
rect 218329 71770 218395 71773
rect 155604 71768 218395 71770
rect 155604 71712 218334 71768
rect 218390 71712 218395 71768
rect 155604 71710 218395 71712
rect 155604 71708 155610 71710
rect 218329 71707 218395 71710
rect 107510 71572 107516 71636
rect 107580 71634 107586 71636
rect 145005 71634 145071 71637
rect 107580 71632 145071 71634
rect 107580 71576 145010 71632
rect 145066 71576 145071 71632
rect 107580 71574 145071 71576
rect 107580 71572 107586 71574
rect 145005 71571 145071 71574
rect 158110 71572 158116 71636
rect 158180 71634 158186 71636
rect 219525 71634 219591 71637
rect 158180 71632 219591 71634
rect 158180 71576 219530 71632
rect 219586 71576 219591 71632
rect 158180 71574 219591 71576
rect 158180 71572 158186 71574
rect 219525 71571 219591 71574
rect 108430 71436 108436 71500
rect 108500 71498 108506 71500
rect 142286 71498 142292 71500
rect 108500 71438 142292 71498
rect 108500 71436 108506 71438
rect 142286 71436 142292 71438
rect 142356 71436 142362 71500
rect 167678 71436 167684 71500
rect 167748 71498 167754 71500
rect 216949 71498 217015 71501
rect 167748 71496 217015 71498
rect 167748 71440 216954 71496
rect 217010 71440 217015 71496
rect 167748 71438 217015 71440
rect 167748 71436 167754 71438
rect 216949 71435 217015 71438
rect 108614 71300 108620 71364
rect 108684 71362 108690 71364
rect 140262 71362 140268 71364
rect 108684 71302 140268 71362
rect 108684 71300 108690 71302
rect 140262 71300 140268 71302
rect 140332 71300 140338 71364
rect 173566 71300 173572 71364
rect 173636 71362 173642 71364
rect 207105 71362 207171 71365
rect 173636 71360 207171 71362
rect 173636 71304 207110 71360
rect 207166 71304 207171 71360
rect 173636 71302 207171 71304
rect 173636 71300 173642 71302
rect 207105 71299 207171 71302
rect 112989 71226 113055 71229
rect 144453 71226 144519 71229
rect 112989 71224 144519 71226
rect 112989 71168 112994 71224
rect 113050 71168 144458 71224
rect 144514 71168 144519 71224
rect 112989 71166 144519 71168
rect 112989 71163 113055 71166
rect 144453 71163 144519 71166
rect 171961 71226 172027 71229
rect 205766 71226 205772 71228
rect 171961 71224 205772 71226
rect 171961 71168 171966 71224
rect 172022 71168 205772 71224
rect 171961 71166 205772 71168
rect 171961 71163 172027 71166
rect 205766 71164 205772 71166
rect 205836 71164 205842 71228
rect 105813 71090 105879 71093
rect 135294 71090 135300 71092
rect 105813 71088 135300 71090
rect 105813 71032 105818 71088
rect 105874 71032 135300 71088
rect 105813 71030 135300 71032
rect 105813 71027 105879 71030
rect 135294 71028 135300 71030
rect 135364 71028 135370 71092
rect 156454 71028 156460 71092
rect 156524 71090 156530 71092
rect 191598 71090 191604 71092
rect 156524 71030 191604 71090
rect 156524 71028 156530 71030
rect 191598 71028 191604 71030
rect 191668 71028 191674 71092
rect 149462 70892 149468 70956
rect 149532 70954 149538 70956
rect 189022 70954 189028 70956
rect 149532 70894 189028 70954
rect 149532 70892 149538 70894
rect 189022 70892 189028 70894
rect 189092 70892 189098 70956
rect 141969 70410 142035 70413
rect 142102 70410 142108 70412
rect 141969 70408 142108 70410
rect 141969 70352 141974 70408
rect 142030 70352 142108 70408
rect 141969 70350 142108 70352
rect 141969 70347 142035 70350
rect 142102 70348 142108 70350
rect 142172 70348 142178 70412
rect 106917 70274 106983 70277
rect 133086 70274 133092 70276
rect 106917 70272 133092 70274
rect 106917 70216 106922 70272
rect 106978 70216 133092 70272
rect 106917 70214 133092 70216
rect 106917 70211 106983 70214
rect 133086 70212 133092 70214
rect 133156 70212 133162 70276
rect 170213 70274 170279 70277
rect 204805 70274 204871 70277
rect 170213 70272 204871 70274
rect 170213 70216 170218 70272
rect 170274 70216 204810 70272
rect 204866 70216 204871 70272
rect 170213 70214 204871 70216
rect 170213 70211 170279 70214
rect 204805 70211 204871 70214
rect 122230 70076 122236 70140
rect 122300 70138 122306 70140
rect 142654 70138 142660 70140
rect 122300 70078 142660 70138
rect 122300 70076 122306 70078
rect 142654 70076 142660 70078
rect 142724 70076 142730 70140
rect 173617 70138 173683 70141
rect 205582 70138 205588 70140
rect 173617 70136 205588 70138
rect 173617 70080 173622 70136
rect 173678 70080 205588 70136
rect 173617 70078 205588 70080
rect 173617 70075 173683 70078
rect 205582 70076 205588 70078
rect 205652 70076 205658 70140
rect 109534 69940 109540 70004
rect 109604 70002 109610 70004
rect 143574 70002 143580 70004
rect 109604 69942 143580 70002
rect 109604 69940 109610 69942
rect 143574 69940 143580 69942
rect 143644 69940 143650 70004
rect 171409 70002 171475 70005
rect 204345 70002 204411 70005
rect 171409 70000 204411 70002
rect 171409 69944 171414 70000
rect 171470 69944 204350 70000
rect 204406 69944 204411 70000
rect 171409 69942 204411 69944
rect 171409 69939 171475 69942
rect 204345 69939 204411 69942
rect 111558 69804 111564 69868
rect 111628 69866 111634 69868
rect 143901 69866 143967 69869
rect 111628 69864 143967 69866
rect 111628 69808 143906 69864
rect 143962 69808 143967 69864
rect 111628 69806 143967 69808
rect 111628 69804 111634 69806
rect 143901 69803 143967 69806
rect 174854 69804 174860 69868
rect 174924 69866 174930 69868
rect 207054 69866 207060 69868
rect 174924 69806 207060 69866
rect 174924 69804 174930 69806
rect 207054 69804 207060 69806
rect 207124 69804 207130 69868
rect 111190 69668 111196 69732
rect 111260 69730 111266 69732
rect 141969 69730 142035 69733
rect 111260 69728 142035 69730
rect 111260 69672 141974 69728
rect 142030 69672 142035 69728
rect 111260 69670 142035 69672
rect 111260 69668 111266 69670
rect 141969 69667 142035 69670
rect 171726 69668 171732 69732
rect 171796 69730 171802 69732
rect 202965 69730 203031 69733
rect 171796 69728 203031 69730
rect 171796 69672 202970 69728
rect 203026 69672 203031 69728
rect 171796 69670 203031 69672
rect 171796 69668 171802 69670
rect 202965 69667 203031 69670
rect 99833 69594 99899 69597
rect 138238 69594 138244 69596
rect 99833 69592 138244 69594
rect 99833 69536 99838 69592
rect 99894 69536 138244 69592
rect 99833 69534 138244 69536
rect 99833 69531 99899 69534
rect 138238 69532 138244 69534
rect 138308 69532 138314 69596
rect 155125 69594 155191 69597
rect 189349 69594 189415 69597
rect 579613 69594 579679 69597
rect 155125 69592 579679 69594
rect 155125 69536 155130 69592
rect 155186 69536 189354 69592
rect 189410 69536 579618 69592
rect 579674 69536 579679 69592
rect 155125 69534 579679 69536
rect 155125 69531 155191 69534
rect 189349 69531 189415 69534
rect 579613 69531 579679 69534
rect 107101 69458 107167 69461
rect 143758 69458 143764 69460
rect 107101 69456 143764 69458
rect 107101 69400 107106 69456
rect 107162 69400 143764 69456
rect 107101 69398 143764 69400
rect 107101 69395 107167 69398
rect 143758 69396 143764 69398
rect 143828 69396 143834 69460
rect 122598 68852 122604 68916
rect 122668 68914 122674 68916
rect 145046 68914 145052 68916
rect 122668 68854 145052 68914
rect 122668 68852 122674 68854
rect 145046 68852 145052 68854
rect 145116 68852 145122 68916
rect 170806 68852 170812 68916
rect 170876 68914 170882 68916
rect 218145 68914 218211 68917
rect 170876 68912 218211 68914
rect 170876 68856 218150 68912
rect 218206 68856 218211 68912
rect 170876 68854 218211 68856
rect 170876 68852 170882 68854
rect 218145 68851 218211 68854
rect 100518 68716 100524 68780
rect 100588 68778 100594 68780
rect 140814 68778 140820 68780
rect 100588 68718 140820 68778
rect 100588 68716 100594 68718
rect 140814 68716 140820 68718
rect 140884 68716 140890 68780
rect 166206 68716 166212 68780
rect 166276 68778 166282 68780
rect 203006 68778 203012 68780
rect 166276 68718 203012 68778
rect 166276 68716 166282 68718
rect 203006 68716 203012 68718
rect 203076 68716 203082 68780
rect 580349 68778 580415 68781
rect 583520 68778 584960 68868
rect 580349 68776 584960 68778
rect 580349 68720 580354 68776
rect 580410 68720 584960 68776
rect 580349 68718 584960 68720
rect 580349 68715 580415 68718
rect 103145 68642 103211 68645
rect 138054 68642 138060 68644
rect 103145 68640 138060 68642
rect 103145 68584 103150 68640
rect 103206 68584 138060 68640
rect 103145 68582 138060 68584
rect 103145 68579 103211 68582
rect 138054 68580 138060 68582
rect 138124 68580 138130 68644
rect 163221 68642 163287 68645
rect 197670 68642 197676 68644
rect 163221 68640 197676 68642
rect 163221 68584 163226 68640
rect 163282 68584 197676 68640
rect 163221 68582 197676 68584
rect 163221 68579 163287 68582
rect 197670 68580 197676 68582
rect 197740 68580 197746 68644
rect 583520 68628 584960 68718
rect 106038 68444 106044 68508
rect 106108 68506 106114 68508
rect 135846 68506 135852 68508
rect 106108 68446 135852 68506
rect 106108 68444 106114 68446
rect 135846 68444 135852 68446
rect 135916 68444 135922 68508
rect 161933 68506 161999 68509
rect 196014 68506 196020 68508
rect 161933 68504 196020 68506
rect 161933 68448 161938 68504
rect 161994 68448 196020 68504
rect 161933 68446 196020 68448
rect 161933 68443 161999 68446
rect 196014 68444 196020 68446
rect 196084 68444 196090 68508
rect 97574 68308 97580 68372
rect 97644 68370 97650 68372
rect 139342 68370 139348 68372
rect 97644 68310 139348 68370
rect 97644 68308 97650 68310
rect 139342 68308 139348 68310
rect 139412 68308 139418 68372
rect 165102 68308 165108 68372
rect 165172 68370 165178 68372
rect 198958 68370 198964 68372
rect 165172 68310 198964 68370
rect 165172 68308 165178 68310
rect 198958 68308 198964 68310
rect 199028 68308 199034 68372
rect -960 68098 480 68188
rect 3509 68098 3575 68101
rect -960 68096 3575 68098
rect -960 68040 3514 68096
rect 3570 68040 3575 68096
rect -960 68038 3575 68040
rect -960 67948 480 68038
rect 3509 68035 3575 68038
rect 103329 67554 103395 67557
rect 145741 67554 145807 67557
rect 103329 67552 145807 67554
rect 103329 67496 103334 67552
rect 103390 67496 145746 67552
rect 145802 67496 145807 67552
rect 103329 67494 145807 67496
rect 103329 67491 103395 67494
rect 145741 67491 145807 67494
rect 146753 67554 146819 67557
rect 147121 67554 147187 67557
rect 146753 67552 147187 67554
rect 146753 67496 146758 67552
rect 146814 67496 147126 67552
rect 147182 67496 147187 67552
rect 146753 67494 147187 67496
rect 146753 67491 146819 67494
rect 147121 67491 147187 67494
rect 152958 67492 152964 67556
rect 153028 67554 153034 67556
rect 219433 67554 219499 67557
rect 153028 67552 219499 67554
rect 153028 67496 219438 67552
rect 219494 67496 219499 67552
rect 153028 67494 219499 67496
rect 153028 67492 153034 67494
rect 219433 67491 219499 67494
rect 97717 67418 97783 67421
rect 138606 67418 138612 67420
rect 97717 67416 138612 67418
rect 97717 67360 97722 67416
rect 97778 67360 138612 67416
rect 97717 67358 138612 67360
rect 97717 67355 97783 67358
rect 138606 67356 138612 67358
rect 138676 67356 138682 67420
rect 159081 67418 159147 67421
rect 193438 67418 193444 67420
rect 159081 67416 193444 67418
rect 159081 67360 159086 67416
rect 159142 67360 193444 67416
rect 159081 67358 193444 67360
rect 159081 67355 159147 67358
rect 193438 67356 193444 67358
rect 193508 67356 193514 67420
rect 104801 67282 104867 67285
rect 138289 67282 138355 67285
rect 104801 67280 138355 67282
rect 104801 67224 104806 67280
rect 104862 67224 138294 67280
rect 138350 67224 138355 67280
rect 104801 67222 138355 67224
rect 104801 67219 104867 67222
rect 138289 67219 138355 67222
rect 174670 67220 174676 67284
rect 174740 67282 174746 67284
rect 208669 67282 208735 67285
rect 174740 67280 208735 67282
rect 174740 67224 208674 67280
rect 208730 67224 208735 67280
rect 174740 67222 208735 67224
rect 174740 67220 174746 67222
rect 208669 67219 208735 67222
rect 99281 67146 99347 67149
rect 132769 67146 132835 67149
rect 99281 67144 132835 67146
rect 99281 67088 99286 67144
rect 99342 67088 132774 67144
rect 132830 67088 132835 67144
rect 99281 67086 132835 67088
rect 99281 67083 99347 67086
rect 132769 67083 132835 67086
rect 176326 67084 176332 67148
rect 176396 67146 176402 67148
rect 208485 67146 208551 67149
rect 176396 67144 208551 67146
rect 176396 67088 208490 67144
rect 208546 67088 208551 67144
rect 176396 67086 208551 67088
rect 176396 67084 176402 67086
rect 208485 67083 208551 67086
rect 115473 67010 115539 67013
rect 147121 67010 147187 67013
rect 115473 67008 147187 67010
rect 115473 66952 115478 67008
rect 115534 66952 147126 67008
rect 147182 66952 147187 67008
rect 115473 66950 147187 66952
rect 115473 66947 115539 66950
rect 147121 66947 147187 66950
rect 157926 66948 157932 67012
rect 157996 67010 158002 67012
rect 186957 67010 187023 67013
rect 157996 67008 187023 67010
rect 157996 66952 186962 67008
rect 187018 66952 187023 67008
rect 157996 66950 187023 66952
rect 157996 66948 158002 66950
rect 186957 66947 187023 66950
rect 119838 66132 119844 66196
rect 119908 66194 119914 66196
rect 149881 66194 149947 66197
rect 119908 66192 149947 66194
rect 119908 66136 149886 66192
rect 149942 66136 149947 66192
rect 119908 66134 149947 66136
rect 119908 66132 119914 66134
rect 149881 66131 149947 66134
rect 154246 66132 154252 66196
rect 154316 66194 154322 66196
rect 218237 66194 218303 66197
rect 154316 66192 218303 66194
rect 154316 66136 218242 66192
rect 218298 66136 218303 66192
rect 154316 66134 218303 66136
rect 154316 66132 154322 66134
rect 218237 66131 218303 66134
rect 113030 65996 113036 66060
rect 113100 66058 113106 66060
rect 141233 66058 141299 66061
rect 113100 66056 141299 66058
rect 113100 66000 141238 66056
rect 141294 66000 141299 66056
rect 113100 65998 141299 66000
rect 113100 65996 113106 65998
rect 141233 65995 141299 65998
rect 154430 65996 154436 66060
rect 154500 66058 154506 66060
rect 216765 66058 216831 66061
rect 154500 66056 216831 66058
rect 154500 66000 216770 66056
rect 216826 66000 216831 66056
rect 154500 65998 216831 66000
rect 154500 65996 154506 65998
rect 216765 65995 216831 65998
rect 160686 65860 160692 65924
rect 160756 65922 160762 65924
rect 221089 65922 221155 65925
rect 160756 65920 221155 65922
rect 160756 65864 221094 65920
rect 221150 65864 221155 65920
rect 160756 65862 221155 65864
rect 160756 65860 160762 65862
rect 221089 65859 221155 65862
rect 154941 65786 155007 65789
rect 161289 65786 161355 65789
rect 154941 65784 161355 65786
rect 154941 65728 154946 65784
rect 155002 65728 161294 65784
rect 161350 65728 161355 65784
rect 154941 65726 161355 65728
rect 154941 65723 155007 65726
rect 161289 65723 161355 65726
rect 170990 65724 170996 65788
rect 171060 65786 171066 65788
rect 204621 65786 204687 65789
rect 171060 65784 204687 65786
rect 171060 65728 204626 65784
rect 204682 65728 204687 65784
rect 171060 65726 204687 65728
rect 171060 65724 171066 65726
rect 204621 65723 204687 65726
rect 161289 65514 161355 65517
rect 187182 65514 187188 65516
rect 161289 65512 187188 65514
rect 161289 65456 161294 65512
rect 161350 65456 187188 65512
rect 161289 65454 187188 65456
rect 161289 65451 161355 65454
rect 187182 65452 187188 65454
rect 187252 65452 187258 65516
rect 102041 64834 102107 64837
rect 133822 64834 133828 64836
rect 102041 64832 133828 64834
rect 102041 64776 102046 64832
rect 102102 64776 133828 64832
rect 102041 64774 133828 64776
rect 102041 64771 102107 64774
rect 133822 64772 133828 64774
rect 133892 64772 133898 64836
rect 172094 64772 172100 64836
rect 172164 64834 172170 64836
rect 214005 64834 214071 64837
rect 172164 64832 214071 64834
rect 172164 64776 214010 64832
rect 214066 64776 214071 64832
rect 172164 64774 214071 64776
rect 172164 64772 172170 64774
rect 214005 64771 214071 64774
rect 113582 64636 113588 64700
rect 113652 64698 113658 64700
rect 141601 64698 141667 64701
rect 113652 64696 141667 64698
rect 113652 64640 141606 64696
rect 141662 64640 141667 64696
rect 113652 64638 141667 64640
rect 113652 64636 113658 64638
rect 141601 64635 141667 64638
rect 176510 64636 176516 64700
rect 176580 64698 176586 64700
rect 215293 64698 215359 64701
rect 176580 64696 215359 64698
rect 176580 64640 215298 64696
rect 215354 64640 215359 64696
rect 176580 64638 215359 64640
rect 176580 64636 176586 64638
rect 215293 64635 215359 64638
rect 161657 64562 161723 64565
rect 196198 64562 196204 64564
rect 161657 64560 196204 64562
rect 161657 64504 161662 64560
rect 161718 64504 196204 64560
rect 161657 64502 196204 64504
rect 161657 64499 161723 64502
rect 196198 64500 196204 64502
rect 196268 64500 196274 64564
rect 583520 64548 584960 64788
rect 166758 64364 166764 64428
rect 166828 64426 166834 64428
rect 200798 64426 200804 64428
rect 166828 64366 200804 64426
rect 166828 64364 166834 64366
rect 200798 64364 200804 64366
rect 200868 64364 200874 64428
rect 167862 64228 167868 64292
rect 167932 64290 167938 64292
rect 201585 64290 201651 64293
rect 167932 64288 201651 64290
rect 167932 64232 201590 64288
rect 201646 64232 201651 64288
rect 167932 64230 201651 64232
rect 167932 64228 167938 64230
rect 201585 64227 201651 64230
rect -960 63868 480 64108
rect 168046 64092 168052 64156
rect 168116 64154 168122 64156
rect 201718 64154 201724 64156
rect 168116 64094 201724 64154
rect 168116 64092 168122 64094
rect 201718 64092 201724 64094
rect 201788 64092 201794 64156
rect 169150 63956 169156 64020
rect 169220 64018 169226 64020
rect 200614 64018 200620 64020
rect 169220 63958 200620 64018
rect 169220 63956 169226 63958
rect 200614 63956 200620 63958
rect 200684 63956 200690 64020
rect 133822 63412 133828 63476
rect 133892 63474 133898 63476
rect 580625 63474 580691 63477
rect 133892 63472 580691 63474
rect 133892 63416 580630 63472
rect 580686 63416 580691 63472
rect 133892 63414 580691 63416
rect 133892 63412 133898 63414
rect 580625 63411 580691 63414
rect 161054 63276 161060 63340
rect 161124 63338 161130 63340
rect 221181 63338 221247 63341
rect 161124 63336 221247 63338
rect 161124 63280 221186 63336
rect 221242 63280 221247 63336
rect 161124 63278 221247 63280
rect 161124 63276 161130 63278
rect 221181 63275 221247 63278
rect 580257 60618 580323 60621
rect 583520 60618 584960 60708
rect 580257 60616 584960 60618
rect 580257 60560 580262 60616
rect 580318 60560 584960 60616
rect 580257 60558 584960 60560
rect 580257 60555 580323 60558
rect 583520 60468 584960 60558
rect -960 59938 480 60028
rect 3509 59938 3575 59941
rect -960 59936 3575 59938
rect -960 59880 3514 59936
rect 3570 59880 3575 59936
rect -960 59878 3575 59880
rect -960 59788 480 59878
rect 3509 59875 3575 59878
rect 579889 56538 579955 56541
rect 583520 56538 584960 56628
rect 579889 56536 584960 56538
rect 579889 56480 579894 56536
rect 579950 56480 584960 56536
rect 579889 56478 584960 56480
rect 579889 56475 579955 56478
rect 583520 56388 584960 56478
rect -960 55708 480 55948
rect 579889 52458 579955 52461
rect 583520 52458 584960 52548
rect 579889 52456 584960 52458
rect 579889 52400 579894 52456
rect 579950 52400 584960 52456
rect 579889 52398 584960 52400
rect 579889 52395 579955 52398
rect 583520 52308 584960 52398
rect -960 51778 480 51868
rect 3509 51778 3575 51781
rect -960 51776 3575 51778
rect -960 51720 3514 51776
rect 3570 51720 3575 51776
rect -960 51718 3575 51720
rect -960 51628 480 51718
rect 3509 51715 3575 51718
rect 580165 48378 580231 48381
rect 583520 48378 584960 48468
rect 580165 48376 584960 48378
rect 580165 48320 580170 48376
rect 580226 48320 584960 48376
rect 580165 48318 584960 48320
rect 580165 48315 580231 48318
rect 583520 48228 584960 48318
rect -960 47698 480 47788
rect 3509 47698 3575 47701
rect -960 47696 3575 47698
rect -960 47640 3514 47696
rect 3570 47640 3575 47696
rect -960 47638 3575 47640
rect -960 47548 480 47638
rect 3509 47635 3575 47638
rect 579981 44298 580047 44301
rect 583520 44298 584960 44388
rect 579981 44296 584960 44298
rect 579981 44240 579986 44296
rect 580042 44240 584960 44296
rect 579981 44238 584960 44240
rect 579981 44235 580047 44238
rect 583520 44148 584960 44238
rect -960 43618 480 43708
rect 3509 43618 3575 43621
rect -960 43616 3575 43618
rect -960 43560 3514 43616
rect 3570 43560 3575 43616
rect -960 43558 3575 43560
rect -960 43468 480 43558
rect 3509 43555 3575 43558
rect 580165 40898 580231 40901
rect 583520 40898 584960 40988
rect 580165 40896 584960 40898
rect 580165 40840 580170 40896
rect 580226 40840 584960 40896
rect 580165 40838 584960 40840
rect 580165 40835 580231 40838
rect 583520 40748 584960 40838
rect -960 39538 480 39628
rect 3509 39538 3575 39541
rect -960 39536 3575 39538
rect -960 39480 3514 39536
rect 3570 39480 3575 39536
rect -960 39478 3575 39480
rect -960 39388 480 39478
rect 3509 39475 3575 39478
rect 580165 36818 580231 36821
rect 583520 36818 584960 36908
rect 580165 36816 584960 36818
rect 580165 36760 580170 36816
rect 580226 36760 584960 36816
rect 580165 36758 584960 36760
rect 580165 36755 580231 36758
rect 583520 36668 584960 36758
rect -960 36138 480 36228
rect 3141 36138 3207 36141
rect -960 36136 3207 36138
rect -960 36080 3146 36136
rect 3202 36080 3207 36136
rect -960 36078 3207 36080
rect -960 35988 480 36078
rect 3141 36075 3207 36078
rect 191782 34444 191788 34508
rect 191852 34506 191858 34508
rect 191925 34506 191991 34509
rect 191852 34504 191991 34506
rect 191852 34448 191930 34504
rect 191986 34448 191991 34504
rect 191852 34446 191991 34448
rect 191852 34444 191858 34446
rect 191925 34443 191991 34446
rect 580165 32738 580231 32741
rect 583520 32738 584960 32828
rect 580165 32736 584960 32738
rect 580165 32680 580170 32736
rect 580226 32680 584960 32736
rect 580165 32678 584960 32680
rect 580165 32675 580231 32678
rect 583520 32588 584960 32678
rect -960 31908 480 32148
rect 580165 28658 580231 28661
rect 583520 28658 584960 28748
rect 580165 28656 584960 28658
rect 580165 28600 580170 28656
rect 580226 28600 584960 28656
rect 580165 28598 584960 28600
rect 580165 28595 580231 28598
rect 583520 28508 584960 28598
rect -960 27978 480 28068
rect 3141 27978 3207 27981
rect -960 27976 3207 27978
rect -960 27920 3146 27976
rect 3202 27920 3207 27976
rect -960 27918 3207 27920
rect -960 27828 480 27918
rect 3141 27915 3207 27918
rect 580165 24578 580231 24581
rect 583520 24578 584960 24668
rect 580165 24576 584960 24578
rect 580165 24520 580170 24576
rect 580226 24520 584960 24576
rect 580165 24518 584960 24520
rect 580165 24515 580231 24518
rect 583520 24428 584960 24518
rect -960 23898 480 23988
rect 3417 23898 3483 23901
rect -960 23896 3483 23898
rect -960 23840 3422 23896
rect 3478 23840 3483 23896
rect -960 23838 3483 23840
rect -960 23748 480 23838
rect 3417 23835 3483 23838
rect 580165 20498 580231 20501
rect 583520 20498 584960 20588
rect 580165 20496 584960 20498
rect 580165 20440 580170 20496
rect 580226 20440 584960 20496
rect 580165 20438 584960 20440
rect 580165 20435 580231 20438
rect 583520 20348 584960 20438
rect -960 19818 480 19908
rect 3141 19818 3207 19821
rect -960 19816 3207 19818
rect -960 19760 3146 19816
rect 3202 19760 3207 19816
rect -960 19758 3207 19760
rect -960 19668 480 19758
rect 3141 19755 3207 19758
rect 580165 16418 580231 16421
rect 583520 16418 584960 16508
rect 580165 16416 584960 16418
rect 580165 16360 580170 16416
rect 580226 16360 584960 16416
rect 580165 16358 584960 16360
rect 580165 16355 580231 16358
rect 583520 16268 584960 16358
rect -960 15738 480 15828
rect 3325 15738 3391 15741
rect -960 15736 3391 15738
rect -960 15680 3330 15736
rect 3386 15680 3391 15736
rect -960 15678 3391 15680
rect -960 15588 480 15678
rect 3325 15675 3391 15678
rect 580165 12338 580231 12341
rect 583520 12338 584960 12428
rect 580165 12336 584960 12338
rect 580165 12280 580170 12336
rect 580226 12280 584960 12336
rect 580165 12278 584960 12280
rect 580165 12275 580231 12278
rect 583520 12188 584960 12278
rect -960 11658 480 11748
rect 3049 11658 3115 11661
rect -960 11656 3115 11658
rect -960 11600 3054 11656
rect 3110 11600 3115 11656
rect -960 11598 3115 11600
rect -960 11508 480 11598
rect 3049 11595 3115 11598
rect 580165 8258 580231 8261
rect 583520 8258 584960 8348
rect 580165 8256 584960 8258
rect 580165 8200 580170 8256
rect 580226 8200 584960 8256
rect 580165 8198 584960 8200
rect 580165 8195 580231 8198
rect 583520 8108 584960 8198
rect -960 7578 480 7668
rect 2957 7578 3023 7581
rect -960 7576 3023 7578
rect -960 7520 2962 7576
rect 3018 7520 3023 7576
rect -960 7518 3023 7520
rect -960 7428 480 7518
rect 2957 7515 3023 7518
rect 580165 4858 580231 4861
rect 583520 4858 584960 4948
rect 580165 4856 584960 4858
rect 580165 4800 580170 4856
rect 580226 4800 584960 4856
rect 580165 4798 584960 4800
rect 580165 4795 580231 4798
rect 583520 4708 584960 4798
rect -960 3498 480 3588
rect 2773 3498 2839 3501
rect -960 3496 2839 3498
rect -960 3440 2778 3496
rect 2834 3440 2839 3496
rect -960 3438 2839 3440
rect -960 3348 480 3438
rect 2773 3435 2839 3438
rect 578877 778 578943 781
rect 583520 778 584960 868
rect 578877 776 584960 778
rect 578877 720 578882 776
rect 578938 720 584960 776
rect 578877 718 584960 720
rect 578877 715 578943 718
rect 583520 628 584960 718
<< via3 >>
rect 95740 656916 95804 656980
rect 191972 263740 192036 263804
rect 118556 263604 118620 263668
rect 191788 263604 191852 263668
rect 187004 259932 187068 259996
rect 187924 259660 187988 259724
rect 122604 259584 122668 259588
rect 122604 259528 122618 259584
rect 122618 259528 122668 259584
rect 122604 259524 122668 259528
rect 187188 259584 187252 259588
rect 187188 259528 187202 259584
rect 187202 259528 187252 259584
rect 187188 259524 187252 259528
rect 188292 233276 188356 233340
rect 122052 227700 122116 227764
rect 186820 220900 186884 220964
rect 122236 211108 122300 211172
rect 186268 208388 186332 208452
rect 121868 207028 121932 207092
rect 176332 201452 176396 201516
rect 122052 200908 122116 200972
rect 121500 200772 121564 200836
rect 156828 200772 156892 200836
rect 168236 200772 168300 200836
rect 186820 200772 186884 200836
rect 203012 200772 203076 200836
rect 138612 200636 138676 200700
rect 152412 200636 152476 200700
rect 186084 200636 186148 200700
rect 187188 200636 187252 200700
rect 207060 200636 207124 200700
rect 138244 200500 138308 200564
rect 173020 200500 173084 200564
rect 145604 200364 145668 200428
rect 176148 200364 176212 200428
rect 139348 200228 139412 200292
rect 121500 200092 121564 200156
rect 122420 200092 122484 200156
rect 147996 200092 148060 200156
rect 149468 200092 149532 200156
rect 153332 200092 153396 200156
rect 154436 200092 154500 200156
rect 133092 199880 133156 199884
rect 133092 199824 133096 199880
rect 133096 199824 133152 199880
rect 133152 199824 133156 199880
rect 133092 199820 133156 199824
rect 133276 199820 133340 199884
rect 133828 199820 133892 199884
rect 134380 199880 134444 199884
rect 134380 199824 134384 199880
rect 134384 199824 134440 199880
rect 134440 199824 134444 199880
rect 134380 199820 134444 199824
rect 138060 199956 138124 200020
rect 136036 199820 136100 199884
rect 137324 199858 137328 199884
rect 137328 199858 137384 199884
rect 137384 199858 137388 199884
rect 137324 199820 137388 199858
rect 138060 199820 138124 199884
rect 160324 200228 160388 200292
rect 161612 200228 161676 200292
rect 160508 200092 160572 200156
rect 161428 200092 161492 200156
rect 203012 200228 203076 200292
rect 138980 199820 139044 199884
rect 139164 199820 139228 199884
rect 139532 199858 139536 199884
rect 139536 199858 139592 199884
rect 139592 199858 139596 199884
rect 139532 199820 139596 199858
rect 139900 199858 139904 199884
rect 139904 199858 139960 199884
rect 139960 199858 139964 199884
rect 139900 199820 139964 199858
rect 140268 199858 140272 199884
rect 140272 199858 140328 199884
rect 140328 199858 140332 199884
rect 140268 199820 140332 199858
rect 140636 199858 140640 199884
rect 140640 199858 140696 199884
rect 140696 199858 140700 199884
rect 140636 199820 140700 199858
rect 141188 199820 141252 199884
rect 142476 199858 142480 199884
rect 142480 199858 142536 199884
rect 142536 199858 142540 199884
rect 142476 199820 142540 199858
rect 143028 199820 143092 199884
rect 144316 199858 144320 199884
rect 144320 199858 144376 199884
rect 144376 199858 144380 199884
rect 144316 199820 144380 199858
rect 144868 199820 144932 199884
rect 145420 199820 145484 199884
rect 145604 199858 145608 199884
rect 145608 199858 145664 199884
rect 145664 199858 145668 199884
rect 145604 199820 145668 199858
rect 146156 199858 146160 199884
rect 146160 199858 146216 199884
rect 146216 199858 146220 199884
rect 146156 199820 146220 199858
rect 146524 199820 146588 199884
rect 147812 199858 147816 199884
rect 147816 199858 147872 199884
rect 147872 199858 147876 199884
rect 147812 199820 147876 199858
rect 148364 199820 148428 199884
rect 148548 199858 148552 199884
rect 148552 199858 148608 199884
rect 148608 199858 148612 199884
rect 148548 199820 148612 199858
rect 148916 199858 148920 199884
rect 148920 199858 148976 199884
rect 148976 199858 148980 199884
rect 148916 199820 148980 199858
rect 149284 199820 149348 199884
rect 149652 199858 149656 199884
rect 149656 199858 149712 199884
rect 149712 199858 149716 199884
rect 149652 199820 149716 199858
rect 150204 199858 150208 199884
rect 150208 199858 150264 199884
rect 150264 199858 150268 199884
rect 150204 199820 150268 199858
rect 150572 199820 150636 199884
rect 151492 199820 151556 199884
rect 152044 199858 152048 199884
rect 152048 199858 152104 199884
rect 152104 199858 152108 199884
rect 152044 199820 152108 199858
rect 152412 199858 152416 199884
rect 152416 199858 152472 199884
rect 152472 199858 152476 199884
rect 152412 199820 152476 199858
rect 153148 199858 153152 199884
rect 153152 199858 153208 199884
rect 153208 199858 153212 199884
rect 153148 199820 153212 199858
rect 153516 199858 153520 199884
rect 153520 199858 153576 199884
rect 153576 199858 153580 199884
rect 153516 199820 153580 199858
rect 154252 199858 154256 199884
rect 154256 199858 154312 199884
rect 154312 199858 154316 199884
rect 154252 199820 154316 199858
rect 154804 199858 154808 199884
rect 154808 199858 154864 199884
rect 154864 199858 154868 199884
rect 154804 199820 154868 199858
rect 156828 199858 156832 199884
rect 156832 199858 156888 199884
rect 156888 199858 156892 199884
rect 156828 199820 156892 199858
rect 158300 199820 158364 199884
rect 158852 199858 158856 199884
rect 158856 199858 158912 199884
rect 158912 199858 158916 199884
rect 158852 199820 158916 199858
rect 159220 199820 159284 199884
rect 160876 199820 160940 199884
rect 161244 199858 161248 199884
rect 161248 199858 161304 199884
rect 161304 199858 161308 199884
rect 161244 199820 161308 199858
rect 161980 199820 162044 199884
rect 162532 199820 162596 199884
rect 162900 199858 162904 199884
rect 162904 199858 162960 199884
rect 162960 199858 162964 199884
rect 162900 199820 162964 199858
rect 163820 199820 163884 199884
rect 164188 199858 164192 199884
rect 164192 199858 164248 199884
rect 164248 199858 164252 199884
rect 164188 199820 164252 199858
rect 165108 199880 165172 199884
rect 165108 199824 165112 199880
rect 165112 199824 165168 199880
rect 165168 199824 165172 199880
rect 165108 199820 165172 199824
rect 166028 199820 166092 199884
rect 168052 199820 168116 199884
rect 168236 199880 168300 199884
rect 168236 199824 168240 199880
rect 168240 199824 168296 199880
rect 168296 199824 168300 199880
rect 168236 199820 168300 199824
rect 160692 199684 160756 199748
rect 122236 199548 122300 199612
rect 161060 199548 161124 199612
rect 161428 199548 161492 199612
rect 162164 199548 162228 199612
rect 166396 199684 166460 199748
rect 121868 199412 121932 199476
rect 133092 199336 133156 199340
rect 133092 199280 133142 199336
rect 133142 199280 133156 199336
rect 133092 199276 133156 199280
rect 133460 199336 133524 199340
rect 133460 199280 133510 199336
rect 133510 199280 133524 199336
rect 133460 199276 133524 199280
rect 133828 199276 133892 199340
rect 134564 199276 134628 199340
rect 135852 199276 135916 199340
rect 136404 199276 136468 199340
rect 136956 199276 137020 199340
rect 137324 199336 137388 199340
rect 137324 199280 137374 199336
rect 137374 199280 137388 199336
rect 137324 199276 137388 199280
rect 138244 199276 138308 199340
rect 153148 199276 153212 199340
rect 160876 199276 160940 199340
rect 161244 199336 161308 199340
rect 161244 199280 161294 199336
rect 161294 199280 161308 199336
rect 161244 199276 161308 199280
rect 161612 199276 161676 199340
rect 162532 199336 162596 199340
rect 162532 199280 162546 199336
rect 162546 199280 162596 199336
rect 162532 199276 162596 199280
rect 162900 199336 162964 199340
rect 162900 199280 162950 199336
rect 162950 199280 162964 199336
rect 162900 199276 162964 199280
rect 133276 199140 133340 199204
rect 134380 199140 134444 199204
rect 136772 199140 136836 199204
rect 138060 199140 138124 199204
rect 139348 199140 139412 199204
rect 141188 199140 141252 199204
rect 143948 199140 144012 199204
rect 146892 199140 146956 199204
rect 147076 199140 147140 199204
rect 149468 199140 149532 199204
rect 158116 199140 158180 199204
rect 158300 199140 158364 199204
rect 167500 199412 167564 199476
rect 168972 199820 169036 199884
rect 169708 199880 169772 199884
rect 169708 199824 169712 199880
rect 169712 199824 169768 199880
rect 169768 199824 169772 199880
rect 169708 199820 169772 199824
rect 170444 199858 170448 199884
rect 170448 199858 170504 199884
rect 170504 199858 170508 199884
rect 170444 199820 170508 199858
rect 172284 199820 172348 199884
rect 173020 199820 173084 199884
rect 173204 199858 173208 199884
rect 173208 199858 173264 199884
rect 173264 199858 173268 199884
rect 173204 199820 173268 199858
rect 169156 199684 169220 199748
rect 173572 199744 173636 199748
rect 173572 199688 173622 199744
rect 173622 199688 173636 199744
rect 173572 199684 173636 199688
rect 170996 199548 171060 199612
rect 173756 199548 173820 199612
rect 174124 199858 174128 199884
rect 174128 199858 174184 199884
rect 174184 199858 174188 199884
rect 174124 199820 174188 199858
rect 177068 200092 177132 200156
rect 176792 199880 176856 199884
rect 176792 199824 176796 199880
rect 176796 199824 176852 199880
rect 176852 199824 176856 199880
rect 176792 199820 176856 199824
rect 177252 199820 177316 199884
rect 174860 199684 174924 199748
rect 207060 200092 207124 200156
rect 176148 199608 176212 199612
rect 176148 199552 176162 199608
rect 176162 199552 176212 199608
rect 176148 199548 176212 199552
rect 176332 199548 176396 199612
rect 177068 199548 177132 199612
rect 169340 199140 169404 199204
rect 170812 199140 170876 199204
rect 211108 199276 211172 199340
rect 114140 199004 114204 199068
rect 150204 199064 150268 199068
rect 150204 199008 150218 199064
rect 150218 199008 150268 199064
rect 150204 199004 150268 199008
rect 151676 199064 151740 199068
rect 151676 199008 151726 199064
rect 151726 199008 151740 199064
rect 151676 199004 151740 199008
rect 109540 198868 109604 198932
rect 149284 198868 149348 198932
rect 188292 198868 188356 198932
rect 138612 198732 138676 198796
rect 140820 198732 140884 198796
rect 144316 198792 144380 198796
rect 144316 198736 144366 198792
rect 144366 198736 144380 198792
rect 144316 198732 144380 198736
rect 149836 198732 149900 198796
rect 150020 198792 150084 198796
rect 150020 198736 150034 198792
rect 150034 198736 150084 198792
rect 150020 198732 150084 198736
rect 151124 198732 151188 198796
rect 153332 198732 153396 198796
rect 154252 198732 154316 198796
rect 154436 198732 154500 198796
rect 158852 198792 158916 198796
rect 158852 198736 158902 198792
rect 158902 198736 158916 198792
rect 158852 198732 158916 198736
rect 159220 198732 159284 198796
rect 160692 198732 160756 198796
rect 165476 198732 165540 198796
rect 124076 198460 124140 198524
rect 136220 198520 136284 198524
rect 136220 198464 136234 198520
rect 136234 198464 136284 198520
rect 122052 198324 122116 198388
rect 136220 198460 136284 198464
rect 136956 198520 137020 198524
rect 136956 198464 137006 198520
rect 137006 198464 137020 198520
rect 136956 198460 137020 198464
rect 138796 198596 138860 198660
rect 141004 198596 141068 198660
rect 144316 198656 144380 198660
rect 144316 198600 144330 198656
rect 144330 198600 144380 198656
rect 144316 198596 144380 198600
rect 138612 198460 138676 198524
rect 146156 198460 146220 198524
rect 150572 198324 150636 198388
rect 151492 198324 151556 198388
rect 154804 198324 154868 198388
rect 166580 198460 166644 198524
rect 172468 198656 172532 198660
rect 172468 198600 172482 198656
rect 172482 198600 172532 198656
rect 172468 198596 172532 198600
rect 174124 198656 174188 198660
rect 174124 198600 174138 198656
rect 174138 198600 174188 198656
rect 174124 198596 174188 198600
rect 175596 198656 175660 198660
rect 175596 198600 175610 198656
rect 175610 198600 175660 198656
rect 175596 198596 175660 198600
rect 173204 198324 173268 198388
rect 139164 198188 139228 198252
rect 139900 198188 139964 198252
rect 104756 197916 104820 197980
rect 138612 198052 138676 198116
rect 138980 198052 139044 198116
rect 139900 198052 139964 198116
rect 143028 198052 143092 198116
rect 144868 198052 144932 198116
rect 148548 198052 148612 198116
rect 152412 198052 152476 198116
rect 154620 198052 154684 198116
rect 165292 198052 165356 198116
rect 166212 198052 166276 198116
rect 168236 198112 168300 198116
rect 168236 198056 168250 198112
rect 168250 198056 168300 198112
rect 149652 197916 149716 197980
rect 138612 197780 138676 197844
rect 146524 197780 146588 197844
rect 168236 198052 168300 198056
rect 174492 198052 174556 198116
rect 139532 197644 139596 197708
rect 140636 197508 140700 197572
rect 140268 197372 140332 197436
rect 147812 197432 147876 197436
rect 147812 197376 147862 197432
rect 147862 197376 147876 197432
rect 147812 197372 147876 197376
rect 142476 197100 142540 197164
rect 173572 196888 173636 196892
rect 173572 196832 173622 196888
rect 173622 196832 173636 196888
rect 173572 196828 173636 196832
rect 174308 196888 174372 196892
rect 174308 196832 174322 196888
rect 174322 196832 174372 196888
rect 174308 196828 174372 196832
rect 108804 196556 108868 196620
rect 142476 196556 142540 196620
rect 147812 196556 147876 196620
rect 152780 196480 152844 196484
rect 152780 196424 152794 196480
rect 152794 196424 152844 196480
rect 152780 196420 152844 196424
rect 158300 196420 158364 196484
rect 160508 196420 160572 196484
rect 196020 196420 196084 196484
rect 138428 196344 138492 196348
rect 138428 196288 138478 196344
rect 138478 196288 138492 196344
rect 138428 196284 138492 196288
rect 152964 196284 153028 196348
rect 163820 196284 163884 196348
rect 166764 196284 166828 196348
rect 168972 196284 169036 196348
rect 154436 196148 154500 196212
rect 157196 196148 157260 196212
rect 165108 196208 165172 196212
rect 165108 196152 165158 196208
rect 165158 196152 165172 196208
rect 165108 196148 165172 196152
rect 168052 196208 168116 196212
rect 168052 196152 168102 196208
rect 168102 196152 168116 196208
rect 168052 196148 168116 196152
rect 137324 196012 137388 196076
rect 153516 196072 153580 196076
rect 153516 196016 153530 196072
rect 153530 196016 153580 196072
rect 153516 196012 153580 196016
rect 157012 196012 157076 196076
rect 158668 196012 158732 196076
rect 160324 196012 160388 196076
rect 161244 196012 161308 196076
rect 164004 196012 164068 196076
rect 168972 196012 169036 196076
rect 177068 196012 177132 196076
rect 122604 195876 122668 195940
rect 133460 195936 133524 195940
rect 133460 195880 133510 195936
rect 133510 195880 133524 195936
rect 133460 195876 133524 195880
rect 136404 195936 136468 195940
rect 136404 195880 136418 195936
rect 136418 195880 136468 195936
rect 136404 195876 136468 195880
rect 139164 195876 139228 195940
rect 140636 195604 140700 195668
rect 166028 195604 166092 195668
rect 122604 195468 122668 195532
rect 162164 195468 162228 195532
rect 170812 195528 170876 195532
rect 170812 195472 170826 195528
rect 170826 195472 170876 195528
rect 170812 195468 170876 195472
rect 113956 195332 114020 195396
rect 172468 195332 172532 195396
rect 117084 195196 117148 195260
rect 169708 195196 169772 195260
rect 176516 194652 176580 194716
rect 121316 194108 121380 194172
rect 196020 194516 196084 194580
rect 196572 194516 196636 194580
rect 205588 194108 205652 194172
rect 121132 193972 121196 194036
rect 97764 193836 97828 193900
rect 134380 193836 134444 193900
rect 161980 193836 162044 193900
rect 187740 193292 187804 193356
rect 136772 192748 136836 192812
rect 175596 192748 175660 192812
rect 120580 192612 120644 192676
rect 147076 192612 147140 192676
rect 147996 192476 148060 192540
rect 200988 192476 201052 192540
rect 148916 192068 148980 192132
rect 198780 191660 198844 191724
rect 95740 191524 95804 191588
rect 174308 191524 174372 191588
rect 151860 191388 151924 191452
rect 201540 191388 201604 191452
rect 117268 191252 117332 191316
rect 164188 191252 164252 191316
rect 197492 191252 197556 191316
rect 104572 191116 104636 191180
rect 158668 191116 158732 191180
rect 193260 191116 193324 191180
rect 194548 190980 194612 191044
rect 197308 190904 197372 190908
rect 197308 190848 197358 190904
rect 197358 190848 197372 190904
rect 197308 190844 197372 190848
rect 134564 190768 134628 190772
rect 134564 190712 134578 190768
rect 134578 190712 134628 190768
rect 134564 190708 134628 190712
rect 168236 190708 168300 190772
rect 198780 190572 198844 190636
rect 122788 190436 122852 190500
rect 148364 190436 148428 190500
rect 154620 190300 154684 190364
rect 157196 190300 157260 190364
rect 111564 190164 111628 190228
rect 139900 190164 139964 190228
rect 166212 190164 166276 190228
rect 190500 190164 190564 190228
rect 117268 190028 117332 190092
rect 158300 190028 158364 190092
rect 143580 189892 143644 189956
rect 174860 189892 174924 189956
rect 207612 189892 207676 189956
rect 107332 189756 107396 189820
rect 192156 189756 192220 189820
rect 205772 189756 205836 189820
rect 108620 189620 108684 189684
rect 157012 189620 157076 189684
rect 122972 189484 123036 189548
rect 172284 189484 172348 189548
rect 116900 189076 116964 189140
rect 117268 189076 117332 189140
rect 167500 189136 167564 189140
rect 167500 189080 167514 189136
rect 167514 189080 167564 189136
rect 167500 189076 167564 189080
rect 138980 189000 139044 189004
rect 138980 188944 138994 189000
rect 138994 188944 139044 189000
rect 138980 188940 139044 188944
rect 205772 188532 205836 188596
rect 122236 188396 122300 188460
rect 182772 188396 182836 188460
rect 149836 188260 149900 188324
rect 189212 188260 189276 188324
rect 170260 187776 170324 187780
rect 170260 187720 170274 187776
rect 170274 187720 170324 187776
rect 170260 187716 170324 187720
rect 199332 187308 199396 187372
rect 113772 187036 113836 187100
rect 108436 186900 108500 186964
rect 145420 186280 145484 186284
rect 145420 186224 145434 186280
rect 145434 186224 145484 186280
rect 145420 186220 145484 186224
rect 169156 186084 169220 186148
rect 173756 185948 173820 186012
rect 203012 185676 203076 185740
rect 111380 185540 111444 185604
rect 174492 185540 174556 185604
rect 107516 184996 107580 185060
rect 139164 184860 139228 184924
rect 119844 184452 119908 184516
rect 112852 184316 112916 184380
rect 146892 184316 146956 184380
rect 164004 184588 164068 184652
rect 166396 184452 166460 184516
rect 170996 184316 171060 184380
rect 108252 184180 108316 184244
rect 147628 184180 147692 184244
rect 168972 184180 169036 184244
rect 198964 184180 199028 184244
rect 158116 183500 158180 183564
rect 189028 183364 189092 183428
rect 189580 183364 189644 183428
rect 152780 183228 152844 183292
rect 189028 183092 189092 183156
rect 154436 182956 154500 183020
rect 188844 182820 188908 182884
rect 152964 181596 153028 181660
rect 122972 181460 123036 181524
rect 151676 181460 151740 181524
rect 107148 181324 107212 181388
rect 150020 181324 150084 181388
rect 106044 181188 106108 181252
rect 103284 181052 103348 181116
rect 101996 180916 102060 180980
rect 100524 180780 100588 180844
rect 122788 180508 122852 180572
rect 169340 180508 169404 180572
rect 203196 180508 203260 180572
rect 204116 180508 204180 180572
rect 166580 180100 166644 180164
rect 200620 180236 200684 180300
rect 204116 180100 204180 180164
rect 166764 179964 166828 180028
rect 200804 179964 200868 180028
rect 165292 179284 165356 179348
rect 187188 179148 187252 179212
rect 186084 179012 186148 179076
rect 134380 178876 134444 178940
rect 161244 178876 161308 178940
rect 161060 178740 161124 178804
rect 185164 178604 185228 178668
rect 97580 178060 97644 178124
rect 121132 177924 121196 177988
rect 113036 177380 113100 177444
rect 140636 177788 140700 177852
rect 104388 177244 104452 177308
rect 138612 177244 138676 177308
rect 135852 176564 135916 176628
rect 140820 176624 140884 176628
rect 140820 176568 140834 176624
rect 140834 176568 140884 176624
rect 140820 176564 140884 176568
rect 141004 175204 141068 175268
rect 137324 175068 137388 175132
rect 122052 174796 122116 174860
rect 102916 174660 102980 174724
rect 103100 174524 103164 174588
rect 137324 174524 137388 174588
rect 122788 171184 122852 171188
rect 122788 171128 122802 171184
rect 122802 171128 122852 171184
rect 122788 171124 122852 171128
rect 122788 171048 122852 171052
rect 122788 170992 122802 171048
rect 122802 170992 122852 171048
rect 122788 170988 122852 170992
rect 122972 161468 123036 161532
rect 122788 161392 122852 161396
rect 122788 161336 122802 161392
rect 122802 161336 122852 161392
rect 122788 161332 122852 161336
rect 122788 151948 122852 152012
rect 122788 151540 122852 151604
rect 111196 148684 111260 148748
rect 100340 148548 100404 148612
rect 112668 148276 112732 148340
rect 144132 148276 144196 148340
rect 165476 148276 165540 148340
rect 122788 147656 122852 147660
rect 122788 147600 122802 147656
rect 122802 147600 122852 147656
rect 122788 147596 122852 147600
rect 197860 146916 197924 146980
rect 197676 145964 197740 146028
rect 196020 145828 196084 145892
rect 187924 145692 187988 145756
rect 111012 144196 111076 144260
rect 115612 144060 115676 144124
rect 187004 143380 187068 143444
rect 118556 143108 118620 143172
rect 191972 143108 192036 143172
rect 191788 142972 191852 143036
rect 118556 141748 118620 141812
rect 115428 141612 115492 141676
rect 118372 141476 118436 141540
rect 191604 141476 191668 141540
rect 119292 141340 119356 141404
rect 186268 140720 186332 140724
rect 186268 140664 186318 140720
rect 186318 140664 186332 140720
rect 186268 140660 186332 140664
rect 115796 140524 115860 140588
rect 185900 140524 185964 140588
rect 116716 140388 116780 140452
rect 191788 140388 191852 140452
rect 119476 140252 119540 140316
rect 151124 140252 151188 140316
rect 187004 140252 187068 140316
rect 119660 140116 119724 140180
rect 118188 139980 118252 140044
rect 196388 139980 196452 140044
rect 124260 139632 124324 139636
rect 124260 139576 124274 139632
rect 124274 139576 124324 139632
rect 124260 139572 124324 139576
rect 123340 139300 123404 139364
rect 123892 139300 123956 139364
rect 130700 139436 130764 139500
rect 183140 139496 183204 139500
rect 183140 139440 183190 139496
rect 183190 139440 183204 139496
rect 183140 139436 183204 139440
rect 120948 139164 121012 139228
rect 124260 139028 124324 139092
rect 116532 138756 116596 138820
rect 176516 139360 176580 139364
rect 176516 139304 176530 139360
rect 176530 139304 176580 139360
rect 176516 139300 176580 139304
rect 186636 139436 186700 139500
rect 196204 139300 196268 139364
rect 199148 139164 199212 139228
rect 176516 138620 176580 138684
rect 201724 138620 201788 138684
rect 130700 138484 130764 138548
rect 183140 138484 183204 138548
rect 191972 138484 192036 138548
rect 122788 138076 122852 138140
rect 185164 138076 185228 138140
rect 187372 138076 187436 138140
rect 186636 137940 186700 138004
rect 182772 137804 182836 137868
rect 186820 137804 186884 137868
rect 188844 137532 188908 137596
rect 193444 137532 193508 137596
rect 187188 137396 187252 137460
rect 186268 137260 186332 137324
rect 186268 136580 186332 136644
rect 113588 136036 113652 136100
rect 123340 136036 123404 136100
rect 187372 135900 187436 135964
rect 186084 134404 186148 134468
rect 186084 133724 186148 133788
rect 197860 104076 197924 104140
rect 120580 95100 120644 95164
rect 187004 91836 187068 91900
rect 186084 91156 186148 91220
rect 187188 91156 187252 91220
rect 186820 88300 186884 88364
rect 187004 83404 187068 83468
rect 189396 82180 189460 82244
rect 186084 82044 186148 82108
rect 133460 81908 133524 81972
rect 172652 81908 172716 81972
rect 132172 81772 132236 81836
rect 175228 81772 175292 81836
rect 199148 81772 199212 81836
rect 129780 81636 129844 81700
rect 185532 81636 185596 81700
rect 122052 81364 122116 81428
rect 135484 81364 135548 81428
rect 191972 81364 192036 81428
rect 107148 81228 107212 81292
rect 138796 81228 138860 81292
rect 171916 81228 171980 81292
rect 202828 81228 202892 81292
rect 119292 81092 119356 81156
rect 151492 81092 151556 81156
rect 158668 81092 158732 81156
rect 191788 81092 191852 81156
rect 134564 80956 134628 81020
rect 157380 80956 157444 81020
rect 139900 80820 139964 80884
rect 164740 80820 164804 80884
rect 175228 80820 175292 80884
rect 100340 80684 100404 80748
rect 132172 80744 132236 80748
rect 132172 80688 132222 80744
rect 132222 80688 132236 80744
rect 132172 80684 132236 80688
rect 133828 80684 133892 80748
rect 152228 80684 152292 80748
rect 120948 80548 121012 80612
rect 124076 80548 124140 80612
rect 136588 80548 136652 80612
rect 171732 80412 171796 80476
rect 192156 80412 192220 80476
rect 115428 80276 115492 80340
rect 134932 80276 134996 80340
rect 115612 80140 115676 80204
rect 112668 80004 112732 80068
rect 137140 80140 137204 80204
rect 137508 80140 137572 80204
rect 133092 79928 133156 79932
rect 133092 79872 133096 79928
rect 133096 79872 133152 79928
rect 133152 79872 133156 79928
rect 133092 79868 133156 79872
rect 133644 79928 133708 79932
rect 133644 79872 133648 79928
rect 133648 79872 133704 79928
rect 133704 79872 133708 79928
rect 133644 79868 133708 79872
rect 134012 79928 134076 79932
rect 134012 79872 134016 79928
rect 134016 79872 134072 79928
rect 134072 79872 134076 79928
rect 134012 79868 134076 79872
rect 140268 80004 140332 80068
rect 133828 79732 133892 79796
rect 134564 79792 134628 79796
rect 134564 79736 134614 79792
rect 134614 79736 134628 79792
rect 134564 79732 134628 79736
rect 133460 79596 133524 79660
rect 134012 79656 134076 79660
rect 134012 79600 134062 79656
rect 134062 79600 134076 79656
rect 134012 79596 134076 79600
rect 135484 79868 135548 79932
rect 136404 79868 136468 79932
rect 136772 79906 136776 79932
rect 136776 79906 136832 79932
rect 136832 79906 136836 79932
rect 136772 79868 136836 79906
rect 134932 79596 134996 79660
rect 136588 79596 136652 79660
rect 138428 79928 138492 79932
rect 138428 79872 138432 79928
rect 138432 79872 138488 79928
rect 138488 79872 138492 79928
rect 138428 79868 138492 79872
rect 138796 79868 138860 79932
rect 139532 79928 139596 79932
rect 139532 79872 139536 79928
rect 139536 79872 139592 79928
rect 139592 79872 139596 79928
rect 139532 79868 139596 79872
rect 138244 79732 138308 79796
rect 139348 79732 139412 79796
rect 139900 79792 139964 79796
rect 139900 79736 139914 79792
rect 139914 79736 139964 79792
rect 139900 79732 139964 79736
rect 141556 79868 141620 79932
rect 142108 79868 142172 79932
rect 145052 80004 145116 80068
rect 142108 79596 142172 79660
rect 143948 79868 144012 79932
rect 144868 79906 144872 79932
rect 144872 79906 144928 79932
rect 144928 79906 144932 79932
rect 144868 79868 144932 79906
rect 155540 80140 155604 80204
rect 146156 79868 146220 79932
rect 146524 79906 146528 79932
rect 146528 79906 146584 79932
rect 146584 79906 146588 79932
rect 146524 79868 146588 79906
rect 143580 79732 143644 79796
rect 147076 79928 147140 79932
rect 147076 79872 147080 79928
rect 147080 79872 147136 79928
rect 147136 79872 147140 79928
rect 147076 79868 147140 79872
rect 148180 79906 148184 79932
rect 148184 79906 148240 79932
rect 148240 79906 148244 79932
rect 148180 79868 148244 79906
rect 147812 79732 147876 79796
rect 148732 79928 148796 79932
rect 148732 79872 148736 79928
rect 148736 79872 148792 79928
rect 148792 79872 148796 79928
rect 148732 79868 148796 79872
rect 149468 79656 149532 79660
rect 149468 79600 149482 79656
rect 149482 79600 149532 79656
rect 149468 79596 149532 79600
rect 151492 79906 151496 79932
rect 151496 79906 151552 79932
rect 151552 79906 151556 79932
rect 151492 79868 151556 79906
rect 152044 79868 152108 79932
rect 152964 79868 153028 79932
rect 154436 79868 154500 79932
rect 154988 79732 155052 79796
rect 154620 79656 154684 79660
rect 154620 79600 154670 79656
rect 154670 79600 154684 79656
rect 154620 79596 154684 79600
rect 152228 79520 152292 79524
rect 152228 79464 152242 79520
rect 152242 79464 152292 79520
rect 152228 79460 152292 79464
rect 111012 79324 111076 79388
rect 172284 80004 172348 80068
rect 157380 79868 157444 79932
rect 158484 79868 158548 79932
rect 158668 79928 158732 79932
rect 158668 79872 158672 79928
rect 158672 79872 158728 79928
rect 158728 79872 158732 79928
rect 158668 79868 158732 79872
rect 158116 79732 158180 79796
rect 160876 79868 160940 79932
rect 161060 79906 161064 79932
rect 161064 79906 161120 79932
rect 161120 79906 161124 79932
rect 161060 79868 161124 79906
rect 161612 79868 161676 79932
rect 162532 79906 162536 79932
rect 162536 79906 162592 79932
rect 162592 79906 162596 79932
rect 162532 79868 162596 79906
rect 163084 79868 163148 79932
rect 163268 79928 163332 79932
rect 163268 79872 163272 79928
rect 163272 79872 163328 79928
rect 163328 79872 163332 79928
rect 163268 79868 163332 79872
rect 162716 79732 162780 79796
rect 164372 79868 164436 79932
rect 164740 79868 164804 79932
rect 164924 79906 164928 79932
rect 164928 79906 164984 79932
rect 164984 79906 164988 79932
rect 164924 79868 164988 79906
rect 165108 79732 165172 79796
rect 164924 79460 164988 79524
rect 160692 79324 160756 79388
rect 163268 79324 163332 79388
rect 166764 79732 166828 79796
rect 167684 79868 167748 79932
rect 167868 79732 167932 79796
rect 170444 79868 170508 79932
rect 170812 79732 170876 79796
rect 170996 79596 171060 79660
rect 172468 79906 172472 79932
rect 172472 79906 172528 79932
rect 172528 79906 172532 79932
rect 172468 79868 172532 79906
rect 172836 79868 172900 79932
rect 173572 79868 173636 79932
rect 173756 79906 173760 79932
rect 173760 79906 173816 79932
rect 173816 79906 173820 79932
rect 173756 79868 173820 79906
rect 171732 79732 171796 79796
rect 172652 79792 172716 79796
rect 172652 79736 172666 79792
rect 172666 79736 172716 79792
rect 172652 79732 172716 79736
rect 174860 79732 174924 79796
rect 175964 79928 176028 79932
rect 175964 79872 175968 79928
rect 175968 79872 176024 79928
rect 176024 79872 176028 79928
rect 175964 79868 176028 79872
rect 176332 79868 176396 79932
rect 174676 79596 174740 79660
rect 189396 79460 189460 79524
rect 185532 79324 185596 79388
rect 189212 79324 189276 79388
rect 107332 79188 107396 79252
rect 154436 79188 154500 79252
rect 186084 79188 186148 79252
rect 116532 79052 116596 79116
rect 163084 79112 163148 79116
rect 163084 79056 163134 79112
rect 163134 79056 163148 79112
rect 163084 79052 163148 79056
rect 122420 78916 122484 78980
rect 166764 78916 166828 78980
rect 168052 78976 168116 78980
rect 168052 78920 168066 78976
rect 168066 78920 168116 78976
rect 168052 78916 168116 78920
rect 171916 78976 171980 78980
rect 171916 78920 171930 78976
rect 171930 78920 171980 78976
rect 171916 78916 171980 78920
rect 108252 78780 108316 78844
rect 146156 78780 146220 78844
rect 133092 78704 133156 78708
rect 133092 78648 133142 78704
rect 133142 78648 133156 78704
rect 133092 78644 133156 78648
rect 138612 78644 138676 78708
rect 142292 78644 142356 78708
rect 143764 78644 143828 78708
rect 119476 78508 119540 78572
rect 121132 78508 121196 78572
rect 139532 78568 139596 78572
rect 139532 78512 139582 78568
rect 139582 78512 139596 78568
rect 139532 78508 139596 78512
rect 141556 78508 141620 78572
rect 154620 78568 154684 78572
rect 154620 78512 154634 78568
rect 154634 78512 154684 78568
rect 154620 78508 154684 78512
rect 154988 78508 155052 78572
rect 162716 78508 162780 78572
rect 172468 78568 172532 78572
rect 172468 78512 172482 78568
rect 172482 78512 172532 78568
rect 172468 78508 172532 78512
rect 172836 78508 172900 78572
rect 175964 78568 176028 78572
rect 175964 78512 175978 78568
rect 175978 78512 176028 78568
rect 175964 78508 176028 78512
rect 176332 78508 176396 78572
rect 101996 78372 102060 78436
rect 133092 78372 133156 78436
rect 169156 78372 169220 78436
rect 171732 78372 171796 78436
rect 103284 78236 103348 78300
rect 135116 78236 135180 78300
rect 136772 78236 136836 78300
rect 141924 78236 141988 78300
rect 123892 78100 123956 78164
rect 136588 78100 136652 78164
rect 211108 78236 211172 78300
rect 187740 78100 187804 78164
rect 104756 77828 104820 77892
rect 136404 77964 136468 78028
rect 138060 78024 138124 78028
rect 138060 77968 138110 78024
rect 138110 77968 138124 78024
rect 138060 77964 138124 77968
rect 140636 77964 140700 78028
rect 161428 77964 161492 78028
rect 97764 77556 97828 77620
rect 142660 77828 142724 77892
rect 152964 77828 153028 77892
rect 158484 77828 158548 77892
rect 173756 77888 173820 77892
rect 173756 77832 173770 77888
rect 173770 77832 173820 77888
rect 121316 77420 121380 77484
rect 148180 77692 148244 77756
rect 173756 77828 173820 77832
rect 176516 77828 176580 77892
rect 172468 77692 172532 77756
rect 140452 77420 140516 77484
rect 160876 77420 160940 77484
rect 135852 77284 135916 77348
rect 104388 77148 104452 77212
rect 135300 77148 135364 77212
rect 104572 77012 104636 77076
rect 164740 77012 164804 77076
rect 170628 77012 170692 77076
rect 108804 76876 108868 76940
rect 113772 76740 113836 76804
rect 203196 76740 203260 76804
rect 116900 76604 116964 76668
rect 140636 76604 140700 76668
rect 140820 76604 140884 76668
rect 143948 76604 144012 76668
rect 144868 76664 144932 76668
rect 144868 76608 144882 76664
rect 144882 76608 144932 76664
rect 144868 76604 144932 76608
rect 146708 76604 146772 76668
rect 156460 76604 156524 76668
rect 162532 76604 162596 76668
rect 170260 76604 170324 76668
rect 200988 76604 201052 76668
rect 138428 76528 138492 76532
rect 138428 76472 138442 76528
rect 138442 76472 138492 76528
rect 138428 76468 138492 76472
rect 129780 76332 129844 76396
rect 190500 76332 190564 76396
rect 134012 76196 134076 76260
rect 152964 75924 153028 75988
rect 154252 75924 154316 75988
rect 157932 75924 157996 75988
rect 170444 75924 170508 75988
rect 154436 75788 154500 75852
rect 192156 75788 192220 75852
rect 113956 75652 114020 75716
rect 146524 75652 146588 75716
rect 161428 75652 161492 75716
rect 114140 75516 114204 75580
rect 161612 75516 161676 75580
rect 201540 75380 201604 75444
rect 102916 75244 102980 75308
rect 187004 75244 187068 75308
rect 133644 75108 133708 75172
rect 118188 74972 118252 75036
rect 166212 74972 166276 75036
rect 176332 74972 176396 75036
rect 147076 74836 147140 74900
rect 148732 74836 148796 74900
rect 170628 74428 170692 74492
rect 197492 74428 197556 74492
rect 111380 74292 111444 74356
rect 194548 74292 194612 74356
rect 119660 74156 119724 74220
rect 103100 74020 103164 74084
rect 135116 74020 135180 74084
rect 207612 74020 207676 74084
rect 116716 73884 116780 73948
rect 117084 73748 117148 73812
rect 166580 73748 166644 73812
rect 170260 73748 170324 73812
rect 196572 73748 196636 73812
rect 118372 73612 118436 73676
rect 193260 73612 193324 73676
rect 118556 73068 118620 73132
rect 140452 73068 140516 73132
rect 172468 73068 172532 73132
rect 112852 72932 112916 72996
rect 146708 72932 146772 72996
rect 196388 72932 196452 72996
rect 152044 72796 152108 72860
rect 197308 72796 197372 72860
rect 115796 72660 115860 72724
rect 198780 72660 198844 72724
rect 136588 72524 136652 72588
rect 147996 72388 148060 72452
rect 199332 72388 199396 72452
rect 155540 71708 155604 71772
rect 107516 71572 107580 71636
rect 158116 71572 158180 71636
rect 108436 71436 108500 71500
rect 142292 71436 142356 71500
rect 167684 71436 167748 71500
rect 108620 71300 108684 71364
rect 140268 71300 140332 71364
rect 173572 71300 173636 71364
rect 205772 71164 205836 71228
rect 135300 71028 135364 71092
rect 156460 71028 156524 71092
rect 191604 71028 191668 71092
rect 149468 70892 149532 70956
rect 189028 70892 189092 70956
rect 142108 70348 142172 70412
rect 133092 70212 133156 70276
rect 122236 70076 122300 70140
rect 142660 70076 142724 70140
rect 205588 70076 205652 70140
rect 109540 69940 109604 70004
rect 143580 69940 143644 70004
rect 111564 69804 111628 69868
rect 174860 69804 174924 69868
rect 207060 69804 207124 69868
rect 111196 69668 111260 69732
rect 171732 69668 171796 69732
rect 138244 69532 138308 69596
rect 143764 69396 143828 69460
rect 122604 68852 122668 68916
rect 145052 68852 145116 68916
rect 170812 68852 170876 68916
rect 100524 68716 100588 68780
rect 140820 68716 140884 68780
rect 166212 68716 166276 68780
rect 203012 68716 203076 68780
rect 138060 68580 138124 68644
rect 197676 68580 197740 68644
rect 106044 68444 106108 68508
rect 135852 68444 135916 68508
rect 196020 68444 196084 68508
rect 97580 68308 97644 68372
rect 139348 68308 139412 68372
rect 165108 68308 165172 68372
rect 198964 68308 199028 68372
rect 152964 67492 153028 67556
rect 138612 67356 138676 67420
rect 193444 67356 193508 67420
rect 174676 67220 174740 67284
rect 176332 67084 176396 67148
rect 157932 66948 157996 67012
rect 119844 66132 119908 66196
rect 154252 66132 154316 66196
rect 113036 65996 113100 66060
rect 154436 65996 154500 66060
rect 160692 65860 160756 65924
rect 170996 65724 171060 65788
rect 187188 65452 187252 65516
rect 133828 64772 133892 64836
rect 172100 64772 172164 64836
rect 113588 64636 113652 64700
rect 176516 64636 176580 64700
rect 196204 64500 196268 64564
rect 166764 64364 166828 64428
rect 200804 64364 200868 64428
rect 167868 64228 167932 64292
rect 168052 64092 168116 64156
rect 201724 64092 201788 64156
rect 169156 63956 169220 64020
rect 200620 63956 200684 64020
rect 133828 63412 133892 63476
rect 161060 63276 161124 63340
rect 191788 34444 191852 34508
<< metal4 >>
rect -8726 711558 -8106 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 -8106 711558
rect -8726 711238 -8106 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 -8106 711238
rect -8726 682954 -8106 711002
rect -8726 682718 -8694 682954
rect -8458 682718 -8374 682954
rect -8138 682718 -8106 682954
rect -8726 682634 -8106 682718
rect -8726 682398 -8694 682634
rect -8458 682398 -8374 682634
rect -8138 682398 -8106 682634
rect -8726 646954 -8106 682398
rect -8726 646718 -8694 646954
rect -8458 646718 -8374 646954
rect -8138 646718 -8106 646954
rect -8726 646634 -8106 646718
rect -8726 646398 -8694 646634
rect -8458 646398 -8374 646634
rect -8138 646398 -8106 646634
rect -8726 610954 -8106 646398
rect -8726 610718 -8694 610954
rect -8458 610718 -8374 610954
rect -8138 610718 -8106 610954
rect -8726 610634 -8106 610718
rect -8726 610398 -8694 610634
rect -8458 610398 -8374 610634
rect -8138 610398 -8106 610634
rect -8726 574954 -8106 610398
rect -8726 574718 -8694 574954
rect -8458 574718 -8374 574954
rect -8138 574718 -8106 574954
rect -8726 574634 -8106 574718
rect -8726 574398 -8694 574634
rect -8458 574398 -8374 574634
rect -8138 574398 -8106 574634
rect -8726 538954 -8106 574398
rect -8726 538718 -8694 538954
rect -8458 538718 -8374 538954
rect -8138 538718 -8106 538954
rect -8726 538634 -8106 538718
rect -8726 538398 -8694 538634
rect -8458 538398 -8374 538634
rect -8138 538398 -8106 538634
rect -8726 502954 -8106 538398
rect -8726 502718 -8694 502954
rect -8458 502718 -8374 502954
rect -8138 502718 -8106 502954
rect -8726 502634 -8106 502718
rect -8726 502398 -8694 502634
rect -8458 502398 -8374 502634
rect -8138 502398 -8106 502634
rect -8726 466954 -8106 502398
rect -8726 466718 -8694 466954
rect -8458 466718 -8374 466954
rect -8138 466718 -8106 466954
rect -8726 466634 -8106 466718
rect -8726 466398 -8694 466634
rect -8458 466398 -8374 466634
rect -8138 466398 -8106 466634
rect -8726 430954 -8106 466398
rect -8726 430718 -8694 430954
rect -8458 430718 -8374 430954
rect -8138 430718 -8106 430954
rect -8726 430634 -8106 430718
rect -8726 430398 -8694 430634
rect -8458 430398 -8374 430634
rect -8138 430398 -8106 430634
rect -8726 394954 -8106 430398
rect -8726 394718 -8694 394954
rect -8458 394718 -8374 394954
rect -8138 394718 -8106 394954
rect -8726 394634 -8106 394718
rect -8726 394398 -8694 394634
rect -8458 394398 -8374 394634
rect -8138 394398 -8106 394634
rect -8726 358954 -8106 394398
rect -8726 358718 -8694 358954
rect -8458 358718 -8374 358954
rect -8138 358718 -8106 358954
rect -8726 358634 -8106 358718
rect -8726 358398 -8694 358634
rect -8458 358398 -8374 358634
rect -8138 358398 -8106 358634
rect -8726 322954 -8106 358398
rect -8726 322718 -8694 322954
rect -8458 322718 -8374 322954
rect -8138 322718 -8106 322954
rect -8726 322634 -8106 322718
rect -8726 322398 -8694 322634
rect -8458 322398 -8374 322634
rect -8138 322398 -8106 322634
rect -8726 286954 -8106 322398
rect -8726 286718 -8694 286954
rect -8458 286718 -8374 286954
rect -8138 286718 -8106 286954
rect -8726 286634 -8106 286718
rect -8726 286398 -8694 286634
rect -8458 286398 -8374 286634
rect -8138 286398 -8106 286634
rect -8726 250954 -8106 286398
rect -8726 250718 -8694 250954
rect -8458 250718 -8374 250954
rect -8138 250718 -8106 250954
rect -8726 250634 -8106 250718
rect -8726 250398 -8694 250634
rect -8458 250398 -8374 250634
rect -8138 250398 -8106 250634
rect -8726 214954 -8106 250398
rect -8726 214718 -8694 214954
rect -8458 214718 -8374 214954
rect -8138 214718 -8106 214954
rect -8726 214634 -8106 214718
rect -8726 214398 -8694 214634
rect -8458 214398 -8374 214634
rect -8138 214398 -8106 214634
rect -8726 178954 -8106 214398
rect -8726 178718 -8694 178954
rect -8458 178718 -8374 178954
rect -8138 178718 -8106 178954
rect -8726 178634 -8106 178718
rect -8726 178398 -8694 178634
rect -8458 178398 -8374 178634
rect -8138 178398 -8106 178634
rect -8726 142954 -8106 178398
rect -8726 142718 -8694 142954
rect -8458 142718 -8374 142954
rect -8138 142718 -8106 142954
rect -8726 142634 -8106 142718
rect -8726 142398 -8694 142634
rect -8458 142398 -8374 142634
rect -8138 142398 -8106 142634
rect -8726 106954 -8106 142398
rect -8726 106718 -8694 106954
rect -8458 106718 -8374 106954
rect -8138 106718 -8106 106954
rect -8726 106634 -8106 106718
rect -8726 106398 -8694 106634
rect -8458 106398 -8374 106634
rect -8138 106398 -8106 106634
rect -8726 70954 -8106 106398
rect -8726 70718 -8694 70954
rect -8458 70718 -8374 70954
rect -8138 70718 -8106 70954
rect -8726 70634 -8106 70718
rect -8726 70398 -8694 70634
rect -8458 70398 -8374 70634
rect -8138 70398 -8106 70634
rect -8726 34954 -8106 70398
rect -8726 34718 -8694 34954
rect -8458 34718 -8374 34954
rect -8138 34718 -8106 34954
rect -8726 34634 -8106 34718
rect -8726 34398 -8694 34634
rect -8458 34398 -8374 34634
rect -8138 34398 -8106 34634
rect -8726 -7066 -8106 34398
rect -7766 710598 -7146 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 -7146 710598
rect -7766 710278 -7146 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 -7146 710278
rect -7766 678454 -7146 710042
rect -7766 678218 -7734 678454
rect -7498 678218 -7414 678454
rect -7178 678218 -7146 678454
rect -7766 678134 -7146 678218
rect -7766 677898 -7734 678134
rect -7498 677898 -7414 678134
rect -7178 677898 -7146 678134
rect -7766 642454 -7146 677898
rect -7766 642218 -7734 642454
rect -7498 642218 -7414 642454
rect -7178 642218 -7146 642454
rect -7766 642134 -7146 642218
rect -7766 641898 -7734 642134
rect -7498 641898 -7414 642134
rect -7178 641898 -7146 642134
rect -7766 606454 -7146 641898
rect -7766 606218 -7734 606454
rect -7498 606218 -7414 606454
rect -7178 606218 -7146 606454
rect -7766 606134 -7146 606218
rect -7766 605898 -7734 606134
rect -7498 605898 -7414 606134
rect -7178 605898 -7146 606134
rect -7766 570454 -7146 605898
rect -7766 570218 -7734 570454
rect -7498 570218 -7414 570454
rect -7178 570218 -7146 570454
rect -7766 570134 -7146 570218
rect -7766 569898 -7734 570134
rect -7498 569898 -7414 570134
rect -7178 569898 -7146 570134
rect -7766 534454 -7146 569898
rect -7766 534218 -7734 534454
rect -7498 534218 -7414 534454
rect -7178 534218 -7146 534454
rect -7766 534134 -7146 534218
rect -7766 533898 -7734 534134
rect -7498 533898 -7414 534134
rect -7178 533898 -7146 534134
rect -7766 498454 -7146 533898
rect -7766 498218 -7734 498454
rect -7498 498218 -7414 498454
rect -7178 498218 -7146 498454
rect -7766 498134 -7146 498218
rect -7766 497898 -7734 498134
rect -7498 497898 -7414 498134
rect -7178 497898 -7146 498134
rect -7766 462454 -7146 497898
rect -7766 462218 -7734 462454
rect -7498 462218 -7414 462454
rect -7178 462218 -7146 462454
rect -7766 462134 -7146 462218
rect -7766 461898 -7734 462134
rect -7498 461898 -7414 462134
rect -7178 461898 -7146 462134
rect -7766 426454 -7146 461898
rect -7766 426218 -7734 426454
rect -7498 426218 -7414 426454
rect -7178 426218 -7146 426454
rect -7766 426134 -7146 426218
rect -7766 425898 -7734 426134
rect -7498 425898 -7414 426134
rect -7178 425898 -7146 426134
rect -7766 390454 -7146 425898
rect -7766 390218 -7734 390454
rect -7498 390218 -7414 390454
rect -7178 390218 -7146 390454
rect -7766 390134 -7146 390218
rect -7766 389898 -7734 390134
rect -7498 389898 -7414 390134
rect -7178 389898 -7146 390134
rect -7766 354454 -7146 389898
rect -7766 354218 -7734 354454
rect -7498 354218 -7414 354454
rect -7178 354218 -7146 354454
rect -7766 354134 -7146 354218
rect -7766 353898 -7734 354134
rect -7498 353898 -7414 354134
rect -7178 353898 -7146 354134
rect -7766 318454 -7146 353898
rect -7766 318218 -7734 318454
rect -7498 318218 -7414 318454
rect -7178 318218 -7146 318454
rect -7766 318134 -7146 318218
rect -7766 317898 -7734 318134
rect -7498 317898 -7414 318134
rect -7178 317898 -7146 318134
rect -7766 282454 -7146 317898
rect -7766 282218 -7734 282454
rect -7498 282218 -7414 282454
rect -7178 282218 -7146 282454
rect -7766 282134 -7146 282218
rect -7766 281898 -7734 282134
rect -7498 281898 -7414 282134
rect -7178 281898 -7146 282134
rect -7766 246454 -7146 281898
rect -7766 246218 -7734 246454
rect -7498 246218 -7414 246454
rect -7178 246218 -7146 246454
rect -7766 246134 -7146 246218
rect -7766 245898 -7734 246134
rect -7498 245898 -7414 246134
rect -7178 245898 -7146 246134
rect -7766 210454 -7146 245898
rect -7766 210218 -7734 210454
rect -7498 210218 -7414 210454
rect -7178 210218 -7146 210454
rect -7766 210134 -7146 210218
rect -7766 209898 -7734 210134
rect -7498 209898 -7414 210134
rect -7178 209898 -7146 210134
rect -7766 174454 -7146 209898
rect -7766 174218 -7734 174454
rect -7498 174218 -7414 174454
rect -7178 174218 -7146 174454
rect -7766 174134 -7146 174218
rect -7766 173898 -7734 174134
rect -7498 173898 -7414 174134
rect -7178 173898 -7146 174134
rect -7766 138454 -7146 173898
rect -7766 138218 -7734 138454
rect -7498 138218 -7414 138454
rect -7178 138218 -7146 138454
rect -7766 138134 -7146 138218
rect -7766 137898 -7734 138134
rect -7498 137898 -7414 138134
rect -7178 137898 -7146 138134
rect -7766 102454 -7146 137898
rect -7766 102218 -7734 102454
rect -7498 102218 -7414 102454
rect -7178 102218 -7146 102454
rect -7766 102134 -7146 102218
rect -7766 101898 -7734 102134
rect -7498 101898 -7414 102134
rect -7178 101898 -7146 102134
rect -7766 66454 -7146 101898
rect -7766 66218 -7734 66454
rect -7498 66218 -7414 66454
rect -7178 66218 -7146 66454
rect -7766 66134 -7146 66218
rect -7766 65898 -7734 66134
rect -7498 65898 -7414 66134
rect -7178 65898 -7146 66134
rect -7766 30454 -7146 65898
rect -7766 30218 -7734 30454
rect -7498 30218 -7414 30454
rect -7178 30218 -7146 30454
rect -7766 30134 -7146 30218
rect -7766 29898 -7734 30134
rect -7498 29898 -7414 30134
rect -7178 29898 -7146 30134
rect -7766 -6106 -7146 29898
rect -6806 709638 -6186 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 -6186 709638
rect -6806 709318 -6186 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 -6186 709318
rect -6806 673954 -6186 709082
rect -6806 673718 -6774 673954
rect -6538 673718 -6454 673954
rect -6218 673718 -6186 673954
rect -6806 673634 -6186 673718
rect -6806 673398 -6774 673634
rect -6538 673398 -6454 673634
rect -6218 673398 -6186 673634
rect -6806 637954 -6186 673398
rect -6806 637718 -6774 637954
rect -6538 637718 -6454 637954
rect -6218 637718 -6186 637954
rect -6806 637634 -6186 637718
rect -6806 637398 -6774 637634
rect -6538 637398 -6454 637634
rect -6218 637398 -6186 637634
rect -6806 601954 -6186 637398
rect -6806 601718 -6774 601954
rect -6538 601718 -6454 601954
rect -6218 601718 -6186 601954
rect -6806 601634 -6186 601718
rect -6806 601398 -6774 601634
rect -6538 601398 -6454 601634
rect -6218 601398 -6186 601634
rect -6806 565954 -6186 601398
rect -6806 565718 -6774 565954
rect -6538 565718 -6454 565954
rect -6218 565718 -6186 565954
rect -6806 565634 -6186 565718
rect -6806 565398 -6774 565634
rect -6538 565398 -6454 565634
rect -6218 565398 -6186 565634
rect -6806 529954 -6186 565398
rect -6806 529718 -6774 529954
rect -6538 529718 -6454 529954
rect -6218 529718 -6186 529954
rect -6806 529634 -6186 529718
rect -6806 529398 -6774 529634
rect -6538 529398 -6454 529634
rect -6218 529398 -6186 529634
rect -6806 493954 -6186 529398
rect -6806 493718 -6774 493954
rect -6538 493718 -6454 493954
rect -6218 493718 -6186 493954
rect -6806 493634 -6186 493718
rect -6806 493398 -6774 493634
rect -6538 493398 -6454 493634
rect -6218 493398 -6186 493634
rect -6806 457954 -6186 493398
rect -6806 457718 -6774 457954
rect -6538 457718 -6454 457954
rect -6218 457718 -6186 457954
rect -6806 457634 -6186 457718
rect -6806 457398 -6774 457634
rect -6538 457398 -6454 457634
rect -6218 457398 -6186 457634
rect -6806 421954 -6186 457398
rect -6806 421718 -6774 421954
rect -6538 421718 -6454 421954
rect -6218 421718 -6186 421954
rect -6806 421634 -6186 421718
rect -6806 421398 -6774 421634
rect -6538 421398 -6454 421634
rect -6218 421398 -6186 421634
rect -6806 385954 -6186 421398
rect -6806 385718 -6774 385954
rect -6538 385718 -6454 385954
rect -6218 385718 -6186 385954
rect -6806 385634 -6186 385718
rect -6806 385398 -6774 385634
rect -6538 385398 -6454 385634
rect -6218 385398 -6186 385634
rect -6806 349954 -6186 385398
rect -6806 349718 -6774 349954
rect -6538 349718 -6454 349954
rect -6218 349718 -6186 349954
rect -6806 349634 -6186 349718
rect -6806 349398 -6774 349634
rect -6538 349398 -6454 349634
rect -6218 349398 -6186 349634
rect -6806 313954 -6186 349398
rect -6806 313718 -6774 313954
rect -6538 313718 -6454 313954
rect -6218 313718 -6186 313954
rect -6806 313634 -6186 313718
rect -6806 313398 -6774 313634
rect -6538 313398 -6454 313634
rect -6218 313398 -6186 313634
rect -6806 277954 -6186 313398
rect -6806 277718 -6774 277954
rect -6538 277718 -6454 277954
rect -6218 277718 -6186 277954
rect -6806 277634 -6186 277718
rect -6806 277398 -6774 277634
rect -6538 277398 -6454 277634
rect -6218 277398 -6186 277634
rect -6806 241954 -6186 277398
rect -6806 241718 -6774 241954
rect -6538 241718 -6454 241954
rect -6218 241718 -6186 241954
rect -6806 241634 -6186 241718
rect -6806 241398 -6774 241634
rect -6538 241398 -6454 241634
rect -6218 241398 -6186 241634
rect -6806 205954 -6186 241398
rect -6806 205718 -6774 205954
rect -6538 205718 -6454 205954
rect -6218 205718 -6186 205954
rect -6806 205634 -6186 205718
rect -6806 205398 -6774 205634
rect -6538 205398 -6454 205634
rect -6218 205398 -6186 205634
rect -6806 169954 -6186 205398
rect -6806 169718 -6774 169954
rect -6538 169718 -6454 169954
rect -6218 169718 -6186 169954
rect -6806 169634 -6186 169718
rect -6806 169398 -6774 169634
rect -6538 169398 -6454 169634
rect -6218 169398 -6186 169634
rect -6806 133954 -6186 169398
rect -6806 133718 -6774 133954
rect -6538 133718 -6454 133954
rect -6218 133718 -6186 133954
rect -6806 133634 -6186 133718
rect -6806 133398 -6774 133634
rect -6538 133398 -6454 133634
rect -6218 133398 -6186 133634
rect -6806 97954 -6186 133398
rect -6806 97718 -6774 97954
rect -6538 97718 -6454 97954
rect -6218 97718 -6186 97954
rect -6806 97634 -6186 97718
rect -6806 97398 -6774 97634
rect -6538 97398 -6454 97634
rect -6218 97398 -6186 97634
rect -6806 61954 -6186 97398
rect -6806 61718 -6774 61954
rect -6538 61718 -6454 61954
rect -6218 61718 -6186 61954
rect -6806 61634 -6186 61718
rect -6806 61398 -6774 61634
rect -6538 61398 -6454 61634
rect -6218 61398 -6186 61634
rect -6806 25954 -6186 61398
rect -6806 25718 -6774 25954
rect -6538 25718 -6454 25954
rect -6218 25718 -6186 25954
rect -6806 25634 -6186 25718
rect -6806 25398 -6774 25634
rect -6538 25398 -6454 25634
rect -6218 25398 -6186 25634
rect -6806 -5146 -6186 25398
rect -5846 708678 -5226 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 -5226 708678
rect -5846 708358 -5226 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 -5226 708358
rect -5846 669454 -5226 708122
rect -5846 669218 -5814 669454
rect -5578 669218 -5494 669454
rect -5258 669218 -5226 669454
rect -5846 669134 -5226 669218
rect -5846 668898 -5814 669134
rect -5578 668898 -5494 669134
rect -5258 668898 -5226 669134
rect -5846 633454 -5226 668898
rect -5846 633218 -5814 633454
rect -5578 633218 -5494 633454
rect -5258 633218 -5226 633454
rect -5846 633134 -5226 633218
rect -5846 632898 -5814 633134
rect -5578 632898 -5494 633134
rect -5258 632898 -5226 633134
rect -5846 597454 -5226 632898
rect -5846 597218 -5814 597454
rect -5578 597218 -5494 597454
rect -5258 597218 -5226 597454
rect -5846 597134 -5226 597218
rect -5846 596898 -5814 597134
rect -5578 596898 -5494 597134
rect -5258 596898 -5226 597134
rect -5846 561454 -5226 596898
rect -5846 561218 -5814 561454
rect -5578 561218 -5494 561454
rect -5258 561218 -5226 561454
rect -5846 561134 -5226 561218
rect -5846 560898 -5814 561134
rect -5578 560898 -5494 561134
rect -5258 560898 -5226 561134
rect -5846 525454 -5226 560898
rect -5846 525218 -5814 525454
rect -5578 525218 -5494 525454
rect -5258 525218 -5226 525454
rect -5846 525134 -5226 525218
rect -5846 524898 -5814 525134
rect -5578 524898 -5494 525134
rect -5258 524898 -5226 525134
rect -5846 489454 -5226 524898
rect -5846 489218 -5814 489454
rect -5578 489218 -5494 489454
rect -5258 489218 -5226 489454
rect -5846 489134 -5226 489218
rect -5846 488898 -5814 489134
rect -5578 488898 -5494 489134
rect -5258 488898 -5226 489134
rect -5846 453454 -5226 488898
rect -5846 453218 -5814 453454
rect -5578 453218 -5494 453454
rect -5258 453218 -5226 453454
rect -5846 453134 -5226 453218
rect -5846 452898 -5814 453134
rect -5578 452898 -5494 453134
rect -5258 452898 -5226 453134
rect -5846 417454 -5226 452898
rect -5846 417218 -5814 417454
rect -5578 417218 -5494 417454
rect -5258 417218 -5226 417454
rect -5846 417134 -5226 417218
rect -5846 416898 -5814 417134
rect -5578 416898 -5494 417134
rect -5258 416898 -5226 417134
rect -5846 381454 -5226 416898
rect -5846 381218 -5814 381454
rect -5578 381218 -5494 381454
rect -5258 381218 -5226 381454
rect -5846 381134 -5226 381218
rect -5846 380898 -5814 381134
rect -5578 380898 -5494 381134
rect -5258 380898 -5226 381134
rect -5846 345454 -5226 380898
rect -5846 345218 -5814 345454
rect -5578 345218 -5494 345454
rect -5258 345218 -5226 345454
rect -5846 345134 -5226 345218
rect -5846 344898 -5814 345134
rect -5578 344898 -5494 345134
rect -5258 344898 -5226 345134
rect -5846 309454 -5226 344898
rect -5846 309218 -5814 309454
rect -5578 309218 -5494 309454
rect -5258 309218 -5226 309454
rect -5846 309134 -5226 309218
rect -5846 308898 -5814 309134
rect -5578 308898 -5494 309134
rect -5258 308898 -5226 309134
rect -5846 273454 -5226 308898
rect -5846 273218 -5814 273454
rect -5578 273218 -5494 273454
rect -5258 273218 -5226 273454
rect -5846 273134 -5226 273218
rect -5846 272898 -5814 273134
rect -5578 272898 -5494 273134
rect -5258 272898 -5226 273134
rect -5846 237454 -5226 272898
rect -5846 237218 -5814 237454
rect -5578 237218 -5494 237454
rect -5258 237218 -5226 237454
rect -5846 237134 -5226 237218
rect -5846 236898 -5814 237134
rect -5578 236898 -5494 237134
rect -5258 236898 -5226 237134
rect -5846 201454 -5226 236898
rect -5846 201218 -5814 201454
rect -5578 201218 -5494 201454
rect -5258 201218 -5226 201454
rect -5846 201134 -5226 201218
rect -5846 200898 -5814 201134
rect -5578 200898 -5494 201134
rect -5258 200898 -5226 201134
rect -5846 165454 -5226 200898
rect -5846 165218 -5814 165454
rect -5578 165218 -5494 165454
rect -5258 165218 -5226 165454
rect -5846 165134 -5226 165218
rect -5846 164898 -5814 165134
rect -5578 164898 -5494 165134
rect -5258 164898 -5226 165134
rect -5846 129454 -5226 164898
rect -5846 129218 -5814 129454
rect -5578 129218 -5494 129454
rect -5258 129218 -5226 129454
rect -5846 129134 -5226 129218
rect -5846 128898 -5814 129134
rect -5578 128898 -5494 129134
rect -5258 128898 -5226 129134
rect -5846 93454 -5226 128898
rect -5846 93218 -5814 93454
rect -5578 93218 -5494 93454
rect -5258 93218 -5226 93454
rect -5846 93134 -5226 93218
rect -5846 92898 -5814 93134
rect -5578 92898 -5494 93134
rect -5258 92898 -5226 93134
rect -5846 57454 -5226 92898
rect -5846 57218 -5814 57454
rect -5578 57218 -5494 57454
rect -5258 57218 -5226 57454
rect -5846 57134 -5226 57218
rect -5846 56898 -5814 57134
rect -5578 56898 -5494 57134
rect -5258 56898 -5226 57134
rect -5846 21454 -5226 56898
rect -5846 21218 -5814 21454
rect -5578 21218 -5494 21454
rect -5258 21218 -5226 21454
rect -5846 21134 -5226 21218
rect -5846 20898 -5814 21134
rect -5578 20898 -5494 21134
rect -5258 20898 -5226 21134
rect -5846 -4186 -5226 20898
rect -4886 707718 -4266 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 -4266 707718
rect -4886 707398 -4266 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 -4266 707398
rect -4886 700954 -4266 707162
rect -4886 700718 -4854 700954
rect -4618 700718 -4534 700954
rect -4298 700718 -4266 700954
rect -4886 700634 -4266 700718
rect -4886 700398 -4854 700634
rect -4618 700398 -4534 700634
rect -4298 700398 -4266 700634
rect -4886 664954 -4266 700398
rect -4886 664718 -4854 664954
rect -4618 664718 -4534 664954
rect -4298 664718 -4266 664954
rect -4886 664634 -4266 664718
rect -4886 664398 -4854 664634
rect -4618 664398 -4534 664634
rect -4298 664398 -4266 664634
rect -4886 628954 -4266 664398
rect -4886 628718 -4854 628954
rect -4618 628718 -4534 628954
rect -4298 628718 -4266 628954
rect -4886 628634 -4266 628718
rect -4886 628398 -4854 628634
rect -4618 628398 -4534 628634
rect -4298 628398 -4266 628634
rect -4886 592954 -4266 628398
rect -4886 592718 -4854 592954
rect -4618 592718 -4534 592954
rect -4298 592718 -4266 592954
rect -4886 592634 -4266 592718
rect -4886 592398 -4854 592634
rect -4618 592398 -4534 592634
rect -4298 592398 -4266 592634
rect -4886 556954 -4266 592398
rect -4886 556718 -4854 556954
rect -4618 556718 -4534 556954
rect -4298 556718 -4266 556954
rect -4886 556634 -4266 556718
rect -4886 556398 -4854 556634
rect -4618 556398 -4534 556634
rect -4298 556398 -4266 556634
rect -4886 520954 -4266 556398
rect -4886 520718 -4854 520954
rect -4618 520718 -4534 520954
rect -4298 520718 -4266 520954
rect -4886 520634 -4266 520718
rect -4886 520398 -4854 520634
rect -4618 520398 -4534 520634
rect -4298 520398 -4266 520634
rect -4886 484954 -4266 520398
rect -4886 484718 -4854 484954
rect -4618 484718 -4534 484954
rect -4298 484718 -4266 484954
rect -4886 484634 -4266 484718
rect -4886 484398 -4854 484634
rect -4618 484398 -4534 484634
rect -4298 484398 -4266 484634
rect -4886 448954 -4266 484398
rect -4886 448718 -4854 448954
rect -4618 448718 -4534 448954
rect -4298 448718 -4266 448954
rect -4886 448634 -4266 448718
rect -4886 448398 -4854 448634
rect -4618 448398 -4534 448634
rect -4298 448398 -4266 448634
rect -4886 412954 -4266 448398
rect -4886 412718 -4854 412954
rect -4618 412718 -4534 412954
rect -4298 412718 -4266 412954
rect -4886 412634 -4266 412718
rect -4886 412398 -4854 412634
rect -4618 412398 -4534 412634
rect -4298 412398 -4266 412634
rect -4886 376954 -4266 412398
rect -4886 376718 -4854 376954
rect -4618 376718 -4534 376954
rect -4298 376718 -4266 376954
rect -4886 376634 -4266 376718
rect -4886 376398 -4854 376634
rect -4618 376398 -4534 376634
rect -4298 376398 -4266 376634
rect -4886 340954 -4266 376398
rect -4886 340718 -4854 340954
rect -4618 340718 -4534 340954
rect -4298 340718 -4266 340954
rect -4886 340634 -4266 340718
rect -4886 340398 -4854 340634
rect -4618 340398 -4534 340634
rect -4298 340398 -4266 340634
rect -4886 304954 -4266 340398
rect -4886 304718 -4854 304954
rect -4618 304718 -4534 304954
rect -4298 304718 -4266 304954
rect -4886 304634 -4266 304718
rect -4886 304398 -4854 304634
rect -4618 304398 -4534 304634
rect -4298 304398 -4266 304634
rect -4886 268954 -4266 304398
rect -4886 268718 -4854 268954
rect -4618 268718 -4534 268954
rect -4298 268718 -4266 268954
rect -4886 268634 -4266 268718
rect -4886 268398 -4854 268634
rect -4618 268398 -4534 268634
rect -4298 268398 -4266 268634
rect -4886 232954 -4266 268398
rect -4886 232718 -4854 232954
rect -4618 232718 -4534 232954
rect -4298 232718 -4266 232954
rect -4886 232634 -4266 232718
rect -4886 232398 -4854 232634
rect -4618 232398 -4534 232634
rect -4298 232398 -4266 232634
rect -4886 196954 -4266 232398
rect -4886 196718 -4854 196954
rect -4618 196718 -4534 196954
rect -4298 196718 -4266 196954
rect -4886 196634 -4266 196718
rect -4886 196398 -4854 196634
rect -4618 196398 -4534 196634
rect -4298 196398 -4266 196634
rect -4886 160954 -4266 196398
rect -4886 160718 -4854 160954
rect -4618 160718 -4534 160954
rect -4298 160718 -4266 160954
rect -4886 160634 -4266 160718
rect -4886 160398 -4854 160634
rect -4618 160398 -4534 160634
rect -4298 160398 -4266 160634
rect -4886 124954 -4266 160398
rect -4886 124718 -4854 124954
rect -4618 124718 -4534 124954
rect -4298 124718 -4266 124954
rect -4886 124634 -4266 124718
rect -4886 124398 -4854 124634
rect -4618 124398 -4534 124634
rect -4298 124398 -4266 124634
rect -4886 88954 -4266 124398
rect -4886 88718 -4854 88954
rect -4618 88718 -4534 88954
rect -4298 88718 -4266 88954
rect -4886 88634 -4266 88718
rect -4886 88398 -4854 88634
rect -4618 88398 -4534 88634
rect -4298 88398 -4266 88634
rect -4886 52954 -4266 88398
rect -4886 52718 -4854 52954
rect -4618 52718 -4534 52954
rect -4298 52718 -4266 52954
rect -4886 52634 -4266 52718
rect -4886 52398 -4854 52634
rect -4618 52398 -4534 52634
rect -4298 52398 -4266 52634
rect -4886 16954 -4266 52398
rect -4886 16718 -4854 16954
rect -4618 16718 -4534 16954
rect -4298 16718 -4266 16954
rect -4886 16634 -4266 16718
rect -4886 16398 -4854 16634
rect -4618 16398 -4534 16634
rect -4298 16398 -4266 16634
rect -4886 -3226 -4266 16398
rect -3926 706758 -3306 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 -3306 706758
rect -3926 706438 -3306 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 -3306 706438
rect -3926 696454 -3306 706202
rect -3926 696218 -3894 696454
rect -3658 696218 -3574 696454
rect -3338 696218 -3306 696454
rect -3926 696134 -3306 696218
rect -3926 695898 -3894 696134
rect -3658 695898 -3574 696134
rect -3338 695898 -3306 696134
rect -3926 660454 -3306 695898
rect -3926 660218 -3894 660454
rect -3658 660218 -3574 660454
rect -3338 660218 -3306 660454
rect -3926 660134 -3306 660218
rect -3926 659898 -3894 660134
rect -3658 659898 -3574 660134
rect -3338 659898 -3306 660134
rect -3926 624454 -3306 659898
rect -3926 624218 -3894 624454
rect -3658 624218 -3574 624454
rect -3338 624218 -3306 624454
rect -3926 624134 -3306 624218
rect -3926 623898 -3894 624134
rect -3658 623898 -3574 624134
rect -3338 623898 -3306 624134
rect -3926 588454 -3306 623898
rect -3926 588218 -3894 588454
rect -3658 588218 -3574 588454
rect -3338 588218 -3306 588454
rect -3926 588134 -3306 588218
rect -3926 587898 -3894 588134
rect -3658 587898 -3574 588134
rect -3338 587898 -3306 588134
rect -3926 552454 -3306 587898
rect -3926 552218 -3894 552454
rect -3658 552218 -3574 552454
rect -3338 552218 -3306 552454
rect -3926 552134 -3306 552218
rect -3926 551898 -3894 552134
rect -3658 551898 -3574 552134
rect -3338 551898 -3306 552134
rect -3926 516454 -3306 551898
rect -3926 516218 -3894 516454
rect -3658 516218 -3574 516454
rect -3338 516218 -3306 516454
rect -3926 516134 -3306 516218
rect -3926 515898 -3894 516134
rect -3658 515898 -3574 516134
rect -3338 515898 -3306 516134
rect -3926 480454 -3306 515898
rect -3926 480218 -3894 480454
rect -3658 480218 -3574 480454
rect -3338 480218 -3306 480454
rect -3926 480134 -3306 480218
rect -3926 479898 -3894 480134
rect -3658 479898 -3574 480134
rect -3338 479898 -3306 480134
rect -3926 444454 -3306 479898
rect -3926 444218 -3894 444454
rect -3658 444218 -3574 444454
rect -3338 444218 -3306 444454
rect -3926 444134 -3306 444218
rect -3926 443898 -3894 444134
rect -3658 443898 -3574 444134
rect -3338 443898 -3306 444134
rect -3926 408454 -3306 443898
rect -3926 408218 -3894 408454
rect -3658 408218 -3574 408454
rect -3338 408218 -3306 408454
rect -3926 408134 -3306 408218
rect -3926 407898 -3894 408134
rect -3658 407898 -3574 408134
rect -3338 407898 -3306 408134
rect -3926 372454 -3306 407898
rect -3926 372218 -3894 372454
rect -3658 372218 -3574 372454
rect -3338 372218 -3306 372454
rect -3926 372134 -3306 372218
rect -3926 371898 -3894 372134
rect -3658 371898 -3574 372134
rect -3338 371898 -3306 372134
rect -3926 336454 -3306 371898
rect -3926 336218 -3894 336454
rect -3658 336218 -3574 336454
rect -3338 336218 -3306 336454
rect -3926 336134 -3306 336218
rect -3926 335898 -3894 336134
rect -3658 335898 -3574 336134
rect -3338 335898 -3306 336134
rect -3926 300454 -3306 335898
rect -3926 300218 -3894 300454
rect -3658 300218 -3574 300454
rect -3338 300218 -3306 300454
rect -3926 300134 -3306 300218
rect -3926 299898 -3894 300134
rect -3658 299898 -3574 300134
rect -3338 299898 -3306 300134
rect -3926 264454 -3306 299898
rect -3926 264218 -3894 264454
rect -3658 264218 -3574 264454
rect -3338 264218 -3306 264454
rect -3926 264134 -3306 264218
rect -3926 263898 -3894 264134
rect -3658 263898 -3574 264134
rect -3338 263898 -3306 264134
rect -3926 228454 -3306 263898
rect -3926 228218 -3894 228454
rect -3658 228218 -3574 228454
rect -3338 228218 -3306 228454
rect -3926 228134 -3306 228218
rect -3926 227898 -3894 228134
rect -3658 227898 -3574 228134
rect -3338 227898 -3306 228134
rect -3926 192454 -3306 227898
rect -3926 192218 -3894 192454
rect -3658 192218 -3574 192454
rect -3338 192218 -3306 192454
rect -3926 192134 -3306 192218
rect -3926 191898 -3894 192134
rect -3658 191898 -3574 192134
rect -3338 191898 -3306 192134
rect -3926 156454 -3306 191898
rect -3926 156218 -3894 156454
rect -3658 156218 -3574 156454
rect -3338 156218 -3306 156454
rect -3926 156134 -3306 156218
rect -3926 155898 -3894 156134
rect -3658 155898 -3574 156134
rect -3338 155898 -3306 156134
rect -3926 120454 -3306 155898
rect -3926 120218 -3894 120454
rect -3658 120218 -3574 120454
rect -3338 120218 -3306 120454
rect -3926 120134 -3306 120218
rect -3926 119898 -3894 120134
rect -3658 119898 -3574 120134
rect -3338 119898 -3306 120134
rect -3926 84454 -3306 119898
rect -3926 84218 -3894 84454
rect -3658 84218 -3574 84454
rect -3338 84218 -3306 84454
rect -3926 84134 -3306 84218
rect -3926 83898 -3894 84134
rect -3658 83898 -3574 84134
rect -3338 83898 -3306 84134
rect -3926 48454 -3306 83898
rect -3926 48218 -3894 48454
rect -3658 48218 -3574 48454
rect -3338 48218 -3306 48454
rect -3926 48134 -3306 48218
rect -3926 47898 -3894 48134
rect -3658 47898 -3574 48134
rect -3338 47898 -3306 48134
rect -3926 12454 -3306 47898
rect -3926 12218 -3894 12454
rect -3658 12218 -3574 12454
rect -3338 12218 -3306 12454
rect -3926 12134 -3306 12218
rect -3926 11898 -3894 12134
rect -3658 11898 -3574 12134
rect -3338 11898 -3306 12134
rect -3926 -2266 -3306 11898
rect -2966 705798 -2346 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 -2346 705798
rect -2966 705478 -2346 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 -2346 705478
rect -2966 691954 -2346 705242
rect -2966 691718 -2934 691954
rect -2698 691718 -2614 691954
rect -2378 691718 -2346 691954
rect -2966 691634 -2346 691718
rect -2966 691398 -2934 691634
rect -2698 691398 -2614 691634
rect -2378 691398 -2346 691634
rect -2966 655954 -2346 691398
rect -2966 655718 -2934 655954
rect -2698 655718 -2614 655954
rect -2378 655718 -2346 655954
rect -2966 655634 -2346 655718
rect -2966 655398 -2934 655634
rect -2698 655398 -2614 655634
rect -2378 655398 -2346 655634
rect -2966 619954 -2346 655398
rect -2966 619718 -2934 619954
rect -2698 619718 -2614 619954
rect -2378 619718 -2346 619954
rect -2966 619634 -2346 619718
rect -2966 619398 -2934 619634
rect -2698 619398 -2614 619634
rect -2378 619398 -2346 619634
rect -2966 583954 -2346 619398
rect -2966 583718 -2934 583954
rect -2698 583718 -2614 583954
rect -2378 583718 -2346 583954
rect -2966 583634 -2346 583718
rect -2966 583398 -2934 583634
rect -2698 583398 -2614 583634
rect -2378 583398 -2346 583634
rect -2966 547954 -2346 583398
rect -2966 547718 -2934 547954
rect -2698 547718 -2614 547954
rect -2378 547718 -2346 547954
rect -2966 547634 -2346 547718
rect -2966 547398 -2934 547634
rect -2698 547398 -2614 547634
rect -2378 547398 -2346 547634
rect -2966 511954 -2346 547398
rect -2966 511718 -2934 511954
rect -2698 511718 -2614 511954
rect -2378 511718 -2346 511954
rect -2966 511634 -2346 511718
rect -2966 511398 -2934 511634
rect -2698 511398 -2614 511634
rect -2378 511398 -2346 511634
rect -2966 475954 -2346 511398
rect -2966 475718 -2934 475954
rect -2698 475718 -2614 475954
rect -2378 475718 -2346 475954
rect -2966 475634 -2346 475718
rect -2966 475398 -2934 475634
rect -2698 475398 -2614 475634
rect -2378 475398 -2346 475634
rect -2966 439954 -2346 475398
rect -2966 439718 -2934 439954
rect -2698 439718 -2614 439954
rect -2378 439718 -2346 439954
rect -2966 439634 -2346 439718
rect -2966 439398 -2934 439634
rect -2698 439398 -2614 439634
rect -2378 439398 -2346 439634
rect -2966 403954 -2346 439398
rect -2966 403718 -2934 403954
rect -2698 403718 -2614 403954
rect -2378 403718 -2346 403954
rect -2966 403634 -2346 403718
rect -2966 403398 -2934 403634
rect -2698 403398 -2614 403634
rect -2378 403398 -2346 403634
rect -2966 367954 -2346 403398
rect -2966 367718 -2934 367954
rect -2698 367718 -2614 367954
rect -2378 367718 -2346 367954
rect -2966 367634 -2346 367718
rect -2966 367398 -2934 367634
rect -2698 367398 -2614 367634
rect -2378 367398 -2346 367634
rect -2966 331954 -2346 367398
rect -2966 331718 -2934 331954
rect -2698 331718 -2614 331954
rect -2378 331718 -2346 331954
rect -2966 331634 -2346 331718
rect -2966 331398 -2934 331634
rect -2698 331398 -2614 331634
rect -2378 331398 -2346 331634
rect -2966 295954 -2346 331398
rect -2966 295718 -2934 295954
rect -2698 295718 -2614 295954
rect -2378 295718 -2346 295954
rect -2966 295634 -2346 295718
rect -2966 295398 -2934 295634
rect -2698 295398 -2614 295634
rect -2378 295398 -2346 295634
rect -2966 259954 -2346 295398
rect -2966 259718 -2934 259954
rect -2698 259718 -2614 259954
rect -2378 259718 -2346 259954
rect -2966 259634 -2346 259718
rect -2966 259398 -2934 259634
rect -2698 259398 -2614 259634
rect -2378 259398 -2346 259634
rect -2966 223954 -2346 259398
rect -2966 223718 -2934 223954
rect -2698 223718 -2614 223954
rect -2378 223718 -2346 223954
rect -2966 223634 -2346 223718
rect -2966 223398 -2934 223634
rect -2698 223398 -2614 223634
rect -2378 223398 -2346 223634
rect -2966 187954 -2346 223398
rect -2966 187718 -2934 187954
rect -2698 187718 -2614 187954
rect -2378 187718 -2346 187954
rect -2966 187634 -2346 187718
rect -2966 187398 -2934 187634
rect -2698 187398 -2614 187634
rect -2378 187398 -2346 187634
rect -2966 151954 -2346 187398
rect -2966 151718 -2934 151954
rect -2698 151718 -2614 151954
rect -2378 151718 -2346 151954
rect -2966 151634 -2346 151718
rect -2966 151398 -2934 151634
rect -2698 151398 -2614 151634
rect -2378 151398 -2346 151634
rect -2966 115954 -2346 151398
rect -2966 115718 -2934 115954
rect -2698 115718 -2614 115954
rect -2378 115718 -2346 115954
rect -2966 115634 -2346 115718
rect -2966 115398 -2934 115634
rect -2698 115398 -2614 115634
rect -2378 115398 -2346 115634
rect -2966 79954 -2346 115398
rect -2966 79718 -2934 79954
rect -2698 79718 -2614 79954
rect -2378 79718 -2346 79954
rect -2966 79634 -2346 79718
rect -2966 79398 -2934 79634
rect -2698 79398 -2614 79634
rect -2378 79398 -2346 79634
rect -2966 43954 -2346 79398
rect -2966 43718 -2934 43954
rect -2698 43718 -2614 43954
rect -2378 43718 -2346 43954
rect -2966 43634 -2346 43718
rect -2966 43398 -2934 43634
rect -2698 43398 -2614 43634
rect -2378 43398 -2346 43634
rect -2966 7954 -2346 43398
rect -2966 7718 -2934 7954
rect -2698 7718 -2614 7954
rect -2378 7718 -2346 7954
rect -2966 7634 -2346 7718
rect -2966 7398 -2934 7634
rect -2698 7398 -2614 7634
rect -2378 7398 -2346 7634
rect -2966 -1306 -2346 7398
rect -2006 704838 -1386 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 -1386 704838
rect -2006 704518 -1386 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 -1386 704518
rect -2006 687454 -1386 704282
rect -2006 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 -1386 687454
rect -2006 687134 -1386 687218
rect -2006 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 -1386 687134
rect -2006 651454 -1386 686898
rect -2006 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 -1386 651454
rect -2006 651134 -1386 651218
rect -2006 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 -1386 651134
rect -2006 615454 -1386 650898
rect -2006 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 -1386 615454
rect -2006 615134 -1386 615218
rect -2006 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 -1386 615134
rect -2006 579454 -1386 614898
rect -2006 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 -1386 579454
rect -2006 579134 -1386 579218
rect -2006 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 -1386 579134
rect -2006 543454 -1386 578898
rect -2006 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 -1386 543454
rect -2006 543134 -1386 543218
rect -2006 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 -1386 543134
rect -2006 507454 -1386 542898
rect -2006 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 -1386 507454
rect -2006 507134 -1386 507218
rect -2006 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 -1386 507134
rect -2006 471454 -1386 506898
rect -2006 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 -1386 471454
rect -2006 471134 -1386 471218
rect -2006 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 -1386 471134
rect -2006 435454 -1386 470898
rect -2006 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 -1386 435454
rect -2006 435134 -1386 435218
rect -2006 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 -1386 435134
rect -2006 399454 -1386 434898
rect -2006 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 -1386 399454
rect -2006 399134 -1386 399218
rect -2006 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 -1386 399134
rect -2006 363454 -1386 398898
rect -2006 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 -1386 363454
rect -2006 363134 -1386 363218
rect -2006 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 -1386 363134
rect -2006 327454 -1386 362898
rect -2006 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 -1386 327454
rect -2006 327134 -1386 327218
rect -2006 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 -1386 327134
rect -2006 291454 -1386 326898
rect -2006 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 -1386 291454
rect -2006 291134 -1386 291218
rect -2006 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 -1386 291134
rect -2006 255454 -1386 290898
rect -2006 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 -1386 255454
rect -2006 255134 -1386 255218
rect -2006 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 -1386 255134
rect -2006 219454 -1386 254898
rect -2006 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 -1386 219454
rect -2006 219134 -1386 219218
rect -2006 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 -1386 219134
rect -2006 183454 -1386 218898
rect -2006 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 -1386 183454
rect -2006 183134 -1386 183218
rect -2006 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 -1386 183134
rect -2006 147454 -1386 182898
rect -2006 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 -1386 147454
rect -2006 147134 -1386 147218
rect -2006 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 -1386 147134
rect -2006 111454 -1386 146898
rect -2006 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 -1386 111454
rect -2006 111134 -1386 111218
rect -2006 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 -1386 111134
rect -2006 75454 -1386 110898
rect -2006 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 -1386 75454
rect -2006 75134 -1386 75218
rect -2006 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 -1386 75134
rect -2006 39454 -1386 74898
rect -2006 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 -1386 39454
rect -2006 39134 -1386 39218
rect -2006 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 -1386 39134
rect -2006 3454 -1386 38898
rect -2006 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 -1386 3454
rect -2006 3134 -1386 3218
rect -2006 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 -1386 3134
rect -2006 -346 -1386 2898
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 -1386 -346
rect -2006 -666 -1386 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 -1386 -666
rect -2006 -934 -1386 -902
rect 1794 704838 2414 711590
rect 1794 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 2414 704838
rect 1794 704518 2414 704602
rect 1794 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 2414 704518
rect 1794 687454 2414 704282
rect 1794 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 2414 687454
rect 1794 687134 2414 687218
rect 1794 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 2414 687134
rect 1794 651454 2414 686898
rect 1794 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 2414 651454
rect 1794 651134 2414 651218
rect 1794 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 2414 651134
rect 1794 615454 2414 650898
rect 1794 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 2414 615454
rect 1794 615134 2414 615218
rect 1794 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 2414 615134
rect 1794 579454 2414 614898
rect 1794 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 2414 579454
rect 1794 579134 2414 579218
rect 1794 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 2414 579134
rect 1794 543454 2414 578898
rect 1794 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 2414 543454
rect 1794 543134 2414 543218
rect 1794 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 2414 543134
rect 1794 507454 2414 542898
rect 1794 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 2414 507454
rect 1794 507134 2414 507218
rect 1794 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 2414 507134
rect 1794 471454 2414 506898
rect 1794 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 2414 471454
rect 1794 471134 2414 471218
rect 1794 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 2414 471134
rect 1794 435454 2414 470898
rect 1794 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 2414 435454
rect 1794 435134 2414 435218
rect 1794 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 2414 435134
rect 1794 399454 2414 434898
rect 1794 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 2414 399454
rect 1794 399134 2414 399218
rect 1794 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 2414 399134
rect 1794 363454 2414 398898
rect 1794 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 2414 363454
rect 1794 363134 2414 363218
rect 1794 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 2414 363134
rect 1794 327454 2414 362898
rect 1794 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 2414 327454
rect 1794 327134 2414 327218
rect 1794 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 2414 327134
rect 1794 291454 2414 326898
rect 1794 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 2414 291454
rect 1794 291134 2414 291218
rect 1794 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 2414 291134
rect 1794 255454 2414 290898
rect 1794 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 2414 255454
rect 1794 255134 2414 255218
rect 1794 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 2414 255134
rect 1794 219454 2414 254898
rect 1794 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 2414 219454
rect 1794 219134 2414 219218
rect 1794 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 2414 219134
rect 1794 183454 2414 218898
rect 1794 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 2414 183454
rect 1794 183134 2414 183218
rect 1794 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 2414 183134
rect 1794 147454 2414 182898
rect 1794 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 2414 147454
rect 1794 147134 2414 147218
rect 1794 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 2414 147134
rect 1794 111454 2414 146898
rect 1794 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 2414 111454
rect 1794 111134 2414 111218
rect 1794 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 2414 111134
rect 1794 75454 2414 110898
rect 1794 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 2414 75454
rect 1794 75134 2414 75218
rect 1794 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 2414 75134
rect 1794 39454 2414 74898
rect 1794 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 2414 39454
rect 1794 39134 2414 39218
rect 1794 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 2414 39134
rect 1794 3454 2414 38898
rect 1794 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 2414 3454
rect 1794 3134 2414 3218
rect 1794 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 2414 3134
rect 1794 -346 2414 2898
rect 1794 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 2414 -346
rect 1794 -666 2414 -582
rect 1794 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 2414 -666
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 -2346 -1306
rect -2966 -1626 -2346 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 -2346 -1626
rect -2966 -1894 -2346 -1862
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 -3306 -2266
rect -3926 -2586 -3306 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 -3306 -2586
rect -3926 -2854 -3306 -2822
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 -4266 -3226
rect -4886 -3546 -4266 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 -4266 -3546
rect -4886 -3814 -4266 -3782
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 -5226 -4186
rect -5846 -4506 -5226 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 -5226 -4506
rect -5846 -4774 -5226 -4742
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 -6186 -5146
rect -6806 -5466 -6186 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 -6186 -5466
rect -6806 -5734 -6186 -5702
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 -7146 -6106
rect -7766 -6426 -7146 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 -7146 -6426
rect -7766 -6694 -7146 -6662
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 -8106 -7066
rect -8726 -7386 -8106 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 -8106 -7386
rect -8726 -7654 -8106 -7622
rect 1794 -7654 2414 -902
rect 6294 705798 6914 711590
rect 6294 705562 6326 705798
rect 6562 705562 6646 705798
rect 6882 705562 6914 705798
rect 6294 705478 6914 705562
rect 6294 705242 6326 705478
rect 6562 705242 6646 705478
rect 6882 705242 6914 705478
rect 6294 691954 6914 705242
rect 6294 691718 6326 691954
rect 6562 691718 6646 691954
rect 6882 691718 6914 691954
rect 6294 691634 6914 691718
rect 6294 691398 6326 691634
rect 6562 691398 6646 691634
rect 6882 691398 6914 691634
rect 6294 655954 6914 691398
rect 6294 655718 6326 655954
rect 6562 655718 6646 655954
rect 6882 655718 6914 655954
rect 6294 655634 6914 655718
rect 6294 655398 6326 655634
rect 6562 655398 6646 655634
rect 6882 655398 6914 655634
rect 6294 619954 6914 655398
rect 6294 619718 6326 619954
rect 6562 619718 6646 619954
rect 6882 619718 6914 619954
rect 6294 619634 6914 619718
rect 6294 619398 6326 619634
rect 6562 619398 6646 619634
rect 6882 619398 6914 619634
rect 6294 583954 6914 619398
rect 6294 583718 6326 583954
rect 6562 583718 6646 583954
rect 6882 583718 6914 583954
rect 6294 583634 6914 583718
rect 6294 583398 6326 583634
rect 6562 583398 6646 583634
rect 6882 583398 6914 583634
rect 6294 547954 6914 583398
rect 6294 547718 6326 547954
rect 6562 547718 6646 547954
rect 6882 547718 6914 547954
rect 6294 547634 6914 547718
rect 6294 547398 6326 547634
rect 6562 547398 6646 547634
rect 6882 547398 6914 547634
rect 6294 511954 6914 547398
rect 6294 511718 6326 511954
rect 6562 511718 6646 511954
rect 6882 511718 6914 511954
rect 6294 511634 6914 511718
rect 6294 511398 6326 511634
rect 6562 511398 6646 511634
rect 6882 511398 6914 511634
rect 6294 475954 6914 511398
rect 6294 475718 6326 475954
rect 6562 475718 6646 475954
rect 6882 475718 6914 475954
rect 6294 475634 6914 475718
rect 6294 475398 6326 475634
rect 6562 475398 6646 475634
rect 6882 475398 6914 475634
rect 6294 439954 6914 475398
rect 6294 439718 6326 439954
rect 6562 439718 6646 439954
rect 6882 439718 6914 439954
rect 6294 439634 6914 439718
rect 6294 439398 6326 439634
rect 6562 439398 6646 439634
rect 6882 439398 6914 439634
rect 6294 403954 6914 439398
rect 6294 403718 6326 403954
rect 6562 403718 6646 403954
rect 6882 403718 6914 403954
rect 6294 403634 6914 403718
rect 6294 403398 6326 403634
rect 6562 403398 6646 403634
rect 6882 403398 6914 403634
rect 6294 367954 6914 403398
rect 6294 367718 6326 367954
rect 6562 367718 6646 367954
rect 6882 367718 6914 367954
rect 6294 367634 6914 367718
rect 6294 367398 6326 367634
rect 6562 367398 6646 367634
rect 6882 367398 6914 367634
rect 6294 331954 6914 367398
rect 6294 331718 6326 331954
rect 6562 331718 6646 331954
rect 6882 331718 6914 331954
rect 6294 331634 6914 331718
rect 6294 331398 6326 331634
rect 6562 331398 6646 331634
rect 6882 331398 6914 331634
rect 6294 295954 6914 331398
rect 6294 295718 6326 295954
rect 6562 295718 6646 295954
rect 6882 295718 6914 295954
rect 6294 295634 6914 295718
rect 6294 295398 6326 295634
rect 6562 295398 6646 295634
rect 6882 295398 6914 295634
rect 6294 259954 6914 295398
rect 6294 259718 6326 259954
rect 6562 259718 6646 259954
rect 6882 259718 6914 259954
rect 6294 259634 6914 259718
rect 6294 259398 6326 259634
rect 6562 259398 6646 259634
rect 6882 259398 6914 259634
rect 6294 223954 6914 259398
rect 6294 223718 6326 223954
rect 6562 223718 6646 223954
rect 6882 223718 6914 223954
rect 6294 223634 6914 223718
rect 6294 223398 6326 223634
rect 6562 223398 6646 223634
rect 6882 223398 6914 223634
rect 6294 187954 6914 223398
rect 6294 187718 6326 187954
rect 6562 187718 6646 187954
rect 6882 187718 6914 187954
rect 6294 187634 6914 187718
rect 6294 187398 6326 187634
rect 6562 187398 6646 187634
rect 6882 187398 6914 187634
rect 6294 151954 6914 187398
rect 6294 151718 6326 151954
rect 6562 151718 6646 151954
rect 6882 151718 6914 151954
rect 6294 151634 6914 151718
rect 6294 151398 6326 151634
rect 6562 151398 6646 151634
rect 6882 151398 6914 151634
rect 6294 115954 6914 151398
rect 6294 115718 6326 115954
rect 6562 115718 6646 115954
rect 6882 115718 6914 115954
rect 6294 115634 6914 115718
rect 6294 115398 6326 115634
rect 6562 115398 6646 115634
rect 6882 115398 6914 115634
rect 6294 79954 6914 115398
rect 6294 79718 6326 79954
rect 6562 79718 6646 79954
rect 6882 79718 6914 79954
rect 6294 79634 6914 79718
rect 6294 79398 6326 79634
rect 6562 79398 6646 79634
rect 6882 79398 6914 79634
rect 6294 43954 6914 79398
rect 6294 43718 6326 43954
rect 6562 43718 6646 43954
rect 6882 43718 6914 43954
rect 6294 43634 6914 43718
rect 6294 43398 6326 43634
rect 6562 43398 6646 43634
rect 6882 43398 6914 43634
rect 6294 7954 6914 43398
rect 6294 7718 6326 7954
rect 6562 7718 6646 7954
rect 6882 7718 6914 7954
rect 6294 7634 6914 7718
rect 6294 7398 6326 7634
rect 6562 7398 6646 7634
rect 6882 7398 6914 7634
rect 6294 -1306 6914 7398
rect 6294 -1542 6326 -1306
rect 6562 -1542 6646 -1306
rect 6882 -1542 6914 -1306
rect 6294 -1626 6914 -1542
rect 6294 -1862 6326 -1626
rect 6562 -1862 6646 -1626
rect 6882 -1862 6914 -1626
rect 6294 -7654 6914 -1862
rect 10794 706758 11414 711590
rect 10794 706522 10826 706758
rect 11062 706522 11146 706758
rect 11382 706522 11414 706758
rect 10794 706438 11414 706522
rect 10794 706202 10826 706438
rect 11062 706202 11146 706438
rect 11382 706202 11414 706438
rect 10794 696454 11414 706202
rect 10794 696218 10826 696454
rect 11062 696218 11146 696454
rect 11382 696218 11414 696454
rect 10794 696134 11414 696218
rect 10794 695898 10826 696134
rect 11062 695898 11146 696134
rect 11382 695898 11414 696134
rect 10794 660454 11414 695898
rect 10794 660218 10826 660454
rect 11062 660218 11146 660454
rect 11382 660218 11414 660454
rect 10794 660134 11414 660218
rect 10794 659898 10826 660134
rect 11062 659898 11146 660134
rect 11382 659898 11414 660134
rect 10794 624454 11414 659898
rect 10794 624218 10826 624454
rect 11062 624218 11146 624454
rect 11382 624218 11414 624454
rect 10794 624134 11414 624218
rect 10794 623898 10826 624134
rect 11062 623898 11146 624134
rect 11382 623898 11414 624134
rect 10794 588454 11414 623898
rect 10794 588218 10826 588454
rect 11062 588218 11146 588454
rect 11382 588218 11414 588454
rect 10794 588134 11414 588218
rect 10794 587898 10826 588134
rect 11062 587898 11146 588134
rect 11382 587898 11414 588134
rect 10794 552454 11414 587898
rect 10794 552218 10826 552454
rect 11062 552218 11146 552454
rect 11382 552218 11414 552454
rect 10794 552134 11414 552218
rect 10794 551898 10826 552134
rect 11062 551898 11146 552134
rect 11382 551898 11414 552134
rect 10794 516454 11414 551898
rect 10794 516218 10826 516454
rect 11062 516218 11146 516454
rect 11382 516218 11414 516454
rect 10794 516134 11414 516218
rect 10794 515898 10826 516134
rect 11062 515898 11146 516134
rect 11382 515898 11414 516134
rect 10794 480454 11414 515898
rect 10794 480218 10826 480454
rect 11062 480218 11146 480454
rect 11382 480218 11414 480454
rect 10794 480134 11414 480218
rect 10794 479898 10826 480134
rect 11062 479898 11146 480134
rect 11382 479898 11414 480134
rect 10794 444454 11414 479898
rect 10794 444218 10826 444454
rect 11062 444218 11146 444454
rect 11382 444218 11414 444454
rect 10794 444134 11414 444218
rect 10794 443898 10826 444134
rect 11062 443898 11146 444134
rect 11382 443898 11414 444134
rect 10794 408454 11414 443898
rect 10794 408218 10826 408454
rect 11062 408218 11146 408454
rect 11382 408218 11414 408454
rect 10794 408134 11414 408218
rect 10794 407898 10826 408134
rect 11062 407898 11146 408134
rect 11382 407898 11414 408134
rect 10794 372454 11414 407898
rect 10794 372218 10826 372454
rect 11062 372218 11146 372454
rect 11382 372218 11414 372454
rect 10794 372134 11414 372218
rect 10794 371898 10826 372134
rect 11062 371898 11146 372134
rect 11382 371898 11414 372134
rect 10794 336454 11414 371898
rect 10794 336218 10826 336454
rect 11062 336218 11146 336454
rect 11382 336218 11414 336454
rect 10794 336134 11414 336218
rect 10794 335898 10826 336134
rect 11062 335898 11146 336134
rect 11382 335898 11414 336134
rect 10794 300454 11414 335898
rect 10794 300218 10826 300454
rect 11062 300218 11146 300454
rect 11382 300218 11414 300454
rect 10794 300134 11414 300218
rect 10794 299898 10826 300134
rect 11062 299898 11146 300134
rect 11382 299898 11414 300134
rect 10794 264454 11414 299898
rect 10794 264218 10826 264454
rect 11062 264218 11146 264454
rect 11382 264218 11414 264454
rect 10794 264134 11414 264218
rect 10794 263898 10826 264134
rect 11062 263898 11146 264134
rect 11382 263898 11414 264134
rect 10794 228454 11414 263898
rect 10794 228218 10826 228454
rect 11062 228218 11146 228454
rect 11382 228218 11414 228454
rect 10794 228134 11414 228218
rect 10794 227898 10826 228134
rect 11062 227898 11146 228134
rect 11382 227898 11414 228134
rect 10794 192454 11414 227898
rect 10794 192218 10826 192454
rect 11062 192218 11146 192454
rect 11382 192218 11414 192454
rect 10794 192134 11414 192218
rect 10794 191898 10826 192134
rect 11062 191898 11146 192134
rect 11382 191898 11414 192134
rect 10794 156454 11414 191898
rect 10794 156218 10826 156454
rect 11062 156218 11146 156454
rect 11382 156218 11414 156454
rect 10794 156134 11414 156218
rect 10794 155898 10826 156134
rect 11062 155898 11146 156134
rect 11382 155898 11414 156134
rect 10794 120454 11414 155898
rect 10794 120218 10826 120454
rect 11062 120218 11146 120454
rect 11382 120218 11414 120454
rect 10794 120134 11414 120218
rect 10794 119898 10826 120134
rect 11062 119898 11146 120134
rect 11382 119898 11414 120134
rect 10794 84454 11414 119898
rect 10794 84218 10826 84454
rect 11062 84218 11146 84454
rect 11382 84218 11414 84454
rect 10794 84134 11414 84218
rect 10794 83898 10826 84134
rect 11062 83898 11146 84134
rect 11382 83898 11414 84134
rect 10794 48454 11414 83898
rect 10794 48218 10826 48454
rect 11062 48218 11146 48454
rect 11382 48218 11414 48454
rect 10794 48134 11414 48218
rect 10794 47898 10826 48134
rect 11062 47898 11146 48134
rect 11382 47898 11414 48134
rect 10794 12454 11414 47898
rect 10794 12218 10826 12454
rect 11062 12218 11146 12454
rect 11382 12218 11414 12454
rect 10794 12134 11414 12218
rect 10794 11898 10826 12134
rect 11062 11898 11146 12134
rect 11382 11898 11414 12134
rect 10794 -2266 11414 11898
rect 10794 -2502 10826 -2266
rect 11062 -2502 11146 -2266
rect 11382 -2502 11414 -2266
rect 10794 -2586 11414 -2502
rect 10794 -2822 10826 -2586
rect 11062 -2822 11146 -2586
rect 11382 -2822 11414 -2586
rect 10794 -7654 11414 -2822
rect 15294 707718 15914 711590
rect 15294 707482 15326 707718
rect 15562 707482 15646 707718
rect 15882 707482 15914 707718
rect 15294 707398 15914 707482
rect 15294 707162 15326 707398
rect 15562 707162 15646 707398
rect 15882 707162 15914 707398
rect 15294 700954 15914 707162
rect 15294 700718 15326 700954
rect 15562 700718 15646 700954
rect 15882 700718 15914 700954
rect 15294 700634 15914 700718
rect 15294 700398 15326 700634
rect 15562 700398 15646 700634
rect 15882 700398 15914 700634
rect 15294 664954 15914 700398
rect 15294 664718 15326 664954
rect 15562 664718 15646 664954
rect 15882 664718 15914 664954
rect 15294 664634 15914 664718
rect 15294 664398 15326 664634
rect 15562 664398 15646 664634
rect 15882 664398 15914 664634
rect 15294 628954 15914 664398
rect 15294 628718 15326 628954
rect 15562 628718 15646 628954
rect 15882 628718 15914 628954
rect 15294 628634 15914 628718
rect 15294 628398 15326 628634
rect 15562 628398 15646 628634
rect 15882 628398 15914 628634
rect 15294 592954 15914 628398
rect 15294 592718 15326 592954
rect 15562 592718 15646 592954
rect 15882 592718 15914 592954
rect 15294 592634 15914 592718
rect 15294 592398 15326 592634
rect 15562 592398 15646 592634
rect 15882 592398 15914 592634
rect 15294 556954 15914 592398
rect 15294 556718 15326 556954
rect 15562 556718 15646 556954
rect 15882 556718 15914 556954
rect 15294 556634 15914 556718
rect 15294 556398 15326 556634
rect 15562 556398 15646 556634
rect 15882 556398 15914 556634
rect 15294 520954 15914 556398
rect 15294 520718 15326 520954
rect 15562 520718 15646 520954
rect 15882 520718 15914 520954
rect 15294 520634 15914 520718
rect 15294 520398 15326 520634
rect 15562 520398 15646 520634
rect 15882 520398 15914 520634
rect 15294 484954 15914 520398
rect 15294 484718 15326 484954
rect 15562 484718 15646 484954
rect 15882 484718 15914 484954
rect 15294 484634 15914 484718
rect 15294 484398 15326 484634
rect 15562 484398 15646 484634
rect 15882 484398 15914 484634
rect 15294 448954 15914 484398
rect 15294 448718 15326 448954
rect 15562 448718 15646 448954
rect 15882 448718 15914 448954
rect 15294 448634 15914 448718
rect 15294 448398 15326 448634
rect 15562 448398 15646 448634
rect 15882 448398 15914 448634
rect 15294 412954 15914 448398
rect 15294 412718 15326 412954
rect 15562 412718 15646 412954
rect 15882 412718 15914 412954
rect 15294 412634 15914 412718
rect 15294 412398 15326 412634
rect 15562 412398 15646 412634
rect 15882 412398 15914 412634
rect 15294 376954 15914 412398
rect 15294 376718 15326 376954
rect 15562 376718 15646 376954
rect 15882 376718 15914 376954
rect 15294 376634 15914 376718
rect 15294 376398 15326 376634
rect 15562 376398 15646 376634
rect 15882 376398 15914 376634
rect 15294 340954 15914 376398
rect 15294 340718 15326 340954
rect 15562 340718 15646 340954
rect 15882 340718 15914 340954
rect 15294 340634 15914 340718
rect 15294 340398 15326 340634
rect 15562 340398 15646 340634
rect 15882 340398 15914 340634
rect 15294 304954 15914 340398
rect 15294 304718 15326 304954
rect 15562 304718 15646 304954
rect 15882 304718 15914 304954
rect 15294 304634 15914 304718
rect 15294 304398 15326 304634
rect 15562 304398 15646 304634
rect 15882 304398 15914 304634
rect 15294 268954 15914 304398
rect 15294 268718 15326 268954
rect 15562 268718 15646 268954
rect 15882 268718 15914 268954
rect 15294 268634 15914 268718
rect 15294 268398 15326 268634
rect 15562 268398 15646 268634
rect 15882 268398 15914 268634
rect 15294 232954 15914 268398
rect 15294 232718 15326 232954
rect 15562 232718 15646 232954
rect 15882 232718 15914 232954
rect 15294 232634 15914 232718
rect 15294 232398 15326 232634
rect 15562 232398 15646 232634
rect 15882 232398 15914 232634
rect 15294 196954 15914 232398
rect 15294 196718 15326 196954
rect 15562 196718 15646 196954
rect 15882 196718 15914 196954
rect 15294 196634 15914 196718
rect 15294 196398 15326 196634
rect 15562 196398 15646 196634
rect 15882 196398 15914 196634
rect 15294 160954 15914 196398
rect 15294 160718 15326 160954
rect 15562 160718 15646 160954
rect 15882 160718 15914 160954
rect 15294 160634 15914 160718
rect 15294 160398 15326 160634
rect 15562 160398 15646 160634
rect 15882 160398 15914 160634
rect 15294 124954 15914 160398
rect 15294 124718 15326 124954
rect 15562 124718 15646 124954
rect 15882 124718 15914 124954
rect 15294 124634 15914 124718
rect 15294 124398 15326 124634
rect 15562 124398 15646 124634
rect 15882 124398 15914 124634
rect 15294 88954 15914 124398
rect 15294 88718 15326 88954
rect 15562 88718 15646 88954
rect 15882 88718 15914 88954
rect 15294 88634 15914 88718
rect 15294 88398 15326 88634
rect 15562 88398 15646 88634
rect 15882 88398 15914 88634
rect 15294 52954 15914 88398
rect 15294 52718 15326 52954
rect 15562 52718 15646 52954
rect 15882 52718 15914 52954
rect 15294 52634 15914 52718
rect 15294 52398 15326 52634
rect 15562 52398 15646 52634
rect 15882 52398 15914 52634
rect 15294 16954 15914 52398
rect 15294 16718 15326 16954
rect 15562 16718 15646 16954
rect 15882 16718 15914 16954
rect 15294 16634 15914 16718
rect 15294 16398 15326 16634
rect 15562 16398 15646 16634
rect 15882 16398 15914 16634
rect 15294 -3226 15914 16398
rect 15294 -3462 15326 -3226
rect 15562 -3462 15646 -3226
rect 15882 -3462 15914 -3226
rect 15294 -3546 15914 -3462
rect 15294 -3782 15326 -3546
rect 15562 -3782 15646 -3546
rect 15882 -3782 15914 -3546
rect 15294 -7654 15914 -3782
rect 19794 708678 20414 711590
rect 19794 708442 19826 708678
rect 20062 708442 20146 708678
rect 20382 708442 20414 708678
rect 19794 708358 20414 708442
rect 19794 708122 19826 708358
rect 20062 708122 20146 708358
rect 20382 708122 20414 708358
rect 19794 669454 20414 708122
rect 19794 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 20414 669454
rect 19794 669134 20414 669218
rect 19794 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 20414 669134
rect 19794 633454 20414 668898
rect 19794 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 20414 633454
rect 19794 633134 20414 633218
rect 19794 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 20414 633134
rect 19794 597454 20414 632898
rect 19794 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 20414 597454
rect 19794 597134 20414 597218
rect 19794 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 20414 597134
rect 19794 561454 20414 596898
rect 19794 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 20414 561454
rect 19794 561134 20414 561218
rect 19794 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 20414 561134
rect 19794 525454 20414 560898
rect 19794 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 20414 525454
rect 19794 525134 20414 525218
rect 19794 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 20414 525134
rect 19794 489454 20414 524898
rect 19794 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 20414 489454
rect 19794 489134 20414 489218
rect 19794 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 20414 489134
rect 19794 453454 20414 488898
rect 19794 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 20414 453454
rect 19794 453134 20414 453218
rect 19794 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 20414 453134
rect 19794 417454 20414 452898
rect 19794 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 20414 417454
rect 19794 417134 20414 417218
rect 19794 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 20414 417134
rect 19794 381454 20414 416898
rect 19794 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 20414 381454
rect 19794 381134 20414 381218
rect 19794 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 20414 381134
rect 19794 345454 20414 380898
rect 19794 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 20414 345454
rect 19794 345134 20414 345218
rect 19794 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 20414 345134
rect 19794 309454 20414 344898
rect 19794 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 20414 309454
rect 19794 309134 20414 309218
rect 19794 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 20414 309134
rect 19794 273454 20414 308898
rect 19794 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 20414 273454
rect 19794 273134 20414 273218
rect 19794 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 20414 273134
rect 19794 237454 20414 272898
rect 19794 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 20414 237454
rect 19794 237134 20414 237218
rect 19794 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 20414 237134
rect 19794 201454 20414 236898
rect 19794 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 20414 201454
rect 19794 201134 20414 201218
rect 19794 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 20414 201134
rect 19794 165454 20414 200898
rect 19794 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 20414 165454
rect 19794 165134 20414 165218
rect 19794 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 20414 165134
rect 19794 129454 20414 164898
rect 19794 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 20414 129454
rect 19794 129134 20414 129218
rect 19794 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 20414 129134
rect 19794 93454 20414 128898
rect 19794 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 20414 93454
rect 19794 93134 20414 93218
rect 19794 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 20414 93134
rect 19794 57454 20414 92898
rect 19794 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 20414 57454
rect 19794 57134 20414 57218
rect 19794 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 20414 57134
rect 19794 21454 20414 56898
rect 19794 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 20414 21454
rect 19794 21134 20414 21218
rect 19794 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 20414 21134
rect 19794 -4186 20414 20898
rect 19794 -4422 19826 -4186
rect 20062 -4422 20146 -4186
rect 20382 -4422 20414 -4186
rect 19794 -4506 20414 -4422
rect 19794 -4742 19826 -4506
rect 20062 -4742 20146 -4506
rect 20382 -4742 20414 -4506
rect 19794 -7654 20414 -4742
rect 24294 709638 24914 711590
rect 24294 709402 24326 709638
rect 24562 709402 24646 709638
rect 24882 709402 24914 709638
rect 24294 709318 24914 709402
rect 24294 709082 24326 709318
rect 24562 709082 24646 709318
rect 24882 709082 24914 709318
rect 24294 673954 24914 709082
rect 24294 673718 24326 673954
rect 24562 673718 24646 673954
rect 24882 673718 24914 673954
rect 24294 673634 24914 673718
rect 24294 673398 24326 673634
rect 24562 673398 24646 673634
rect 24882 673398 24914 673634
rect 24294 637954 24914 673398
rect 24294 637718 24326 637954
rect 24562 637718 24646 637954
rect 24882 637718 24914 637954
rect 24294 637634 24914 637718
rect 24294 637398 24326 637634
rect 24562 637398 24646 637634
rect 24882 637398 24914 637634
rect 24294 601954 24914 637398
rect 24294 601718 24326 601954
rect 24562 601718 24646 601954
rect 24882 601718 24914 601954
rect 24294 601634 24914 601718
rect 24294 601398 24326 601634
rect 24562 601398 24646 601634
rect 24882 601398 24914 601634
rect 24294 565954 24914 601398
rect 24294 565718 24326 565954
rect 24562 565718 24646 565954
rect 24882 565718 24914 565954
rect 24294 565634 24914 565718
rect 24294 565398 24326 565634
rect 24562 565398 24646 565634
rect 24882 565398 24914 565634
rect 24294 529954 24914 565398
rect 24294 529718 24326 529954
rect 24562 529718 24646 529954
rect 24882 529718 24914 529954
rect 24294 529634 24914 529718
rect 24294 529398 24326 529634
rect 24562 529398 24646 529634
rect 24882 529398 24914 529634
rect 24294 493954 24914 529398
rect 24294 493718 24326 493954
rect 24562 493718 24646 493954
rect 24882 493718 24914 493954
rect 24294 493634 24914 493718
rect 24294 493398 24326 493634
rect 24562 493398 24646 493634
rect 24882 493398 24914 493634
rect 24294 457954 24914 493398
rect 24294 457718 24326 457954
rect 24562 457718 24646 457954
rect 24882 457718 24914 457954
rect 24294 457634 24914 457718
rect 24294 457398 24326 457634
rect 24562 457398 24646 457634
rect 24882 457398 24914 457634
rect 24294 421954 24914 457398
rect 24294 421718 24326 421954
rect 24562 421718 24646 421954
rect 24882 421718 24914 421954
rect 24294 421634 24914 421718
rect 24294 421398 24326 421634
rect 24562 421398 24646 421634
rect 24882 421398 24914 421634
rect 24294 385954 24914 421398
rect 24294 385718 24326 385954
rect 24562 385718 24646 385954
rect 24882 385718 24914 385954
rect 24294 385634 24914 385718
rect 24294 385398 24326 385634
rect 24562 385398 24646 385634
rect 24882 385398 24914 385634
rect 24294 349954 24914 385398
rect 24294 349718 24326 349954
rect 24562 349718 24646 349954
rect 24882 349718 24914 349954
rect 24294 349634 24914 349718
rect 24294 349398 24326 349634
rect 24562 349398 24646 349634
rect 24882 349398 24914 349634
rect 24294 313954 24914 349398
rect 24294 313718 24326 313954
rect 24562 313718 24646 313954
rect 24882 313718 24914 313954
rect 24294 313634 24914 313718
rect 24294 313398 24326 313634
rect 24562 313398 24646 313634
rect 24882 313398 24914 313634
rect 24294 277954 24914 313398
rect 24294 277718 24326 277954
rect 24562 277718 24646 277954
rect 24882 277718 24914 277954
rect 24294 277634 24914 277718
rect 24294 277398 24326 277634
rect 24562 277398 24646 277634
rect 24882 277398 24914 277634
rect 24294 241954 24914 277398
rect 24294 241718 24326 241954
rect 24562 241718 24646 241954
rect 24882 241718 24914 241954
rect 24294 241634 24914 241718
rect 24294 241398 24326 241634
rect 24562 241398 24646 241634
rect 24882 241398 24914 241634
rect 24294 205954 24914 241398
rect 24294 205718 24326 205954
rect 24562 205718 24646 205954
rect 24882 205718 24914 205954
rect 24294 205634 24914 205718
rect 24294 205398 24326 205634
rect 24562 205398 24646 205634
rect 24882 205398 24914 205634
rect 24294 169954 24914 205398
rect 24294 169718 24326 169954
rect 24562 169718 24646 169954
rect 24882 169718 24914 169954
rect 24294 169634 24914 169718
rect 24294 169398 24326 169634
rect 24562 169398 24646 169634
rect 24882 169398 24914 169634
rect 24294 133954 24914 169398
rect 24294 133718 24326 133954
rect 24562 133718 24646 133954
rect 24882 133718 24914 133954
rect 24294 133634 24914 133718
rect 24294 133398 24326 133634
rect 24562 133398 24646 133634
rect 24882 133398 24914 133634
rect 24294 97954 24914 133398
rect 24294 97718 24326 97954
rect 24562 97718 24646 97954
rect 24882 97718 24914 97954
rect 24294 97634 24914 97718
rect 24294 97398 24326 97634
rect 24562 97398 24646 97634
rect 24882 97398 24914 97634
rect 24294 61954 24914 97398
rect 24294 61718 24326 61954
rect 24562 61718 24646 61954
rect 24882 61718 24914 61954
rect 24294 61634 24914 61718
rect 24294 61398 24326 61634
rect 24562 61398 24646 61634
rect 24882 61398 24914 61634
rect 24294 25954 24914 61398
rect 24294 25718 24326 25954
rect 24562 25718 24646 25954
rect 24882 25718 24914 25954
rect 24294 25634 24914 25718
rect 24294 25398 24326 25634
rect 24562 25398 24646 25634
rect 24882 25398 24914 25634
rect 24294 -5146 24914 25398
rect 24294 -5382 24326 -5146
rect 24562 -5382 24646 -5146
rect 24882 -5382 24914 -5146
rect 24294 -5466 24914 -5382
rect 24294 -5702 24326 -5466
rect 24562 -5702 24646 -5466
rect 24882 -5702 24914 -5466
rect 24294 -7654 24914 -5702
rect 28794 710598 29414 711590
rect 28794 710362 28826 710598
rect 29062 710362 29146 710598
rect 29382 710362 29414 710598
rect 28794 710278 29414 710362
rect 28794 710042 28826 710278
rect 29062 710042 29146 710278
rect 29382 710042 29414 710278
rect 28794 678454 29414 710042
rect 28794 678218 28826 678454
rect 29062 678218 29146 678454
rect 29382 678218 29414 678454
rect 28794 678134 29414 678218
rect 28794 677898 28826 678134
rect 29062 677898 29146 678134
rect 29382 677898 29414 678134
rect 28794 642454 29414 677898
rect 28794 642218 28826 642454
rect 29062 642218 29146 642454
rect 29382 642218 29414 642454
rect 28794 642134 29414 642218
rect 28794 641898 28826 642134
rect 29062 641898 29146 642134
rect 29382 641898 29414 642134
rect 28794 606454 29414 641898
rect 28794 606218 28826 606454
rect 29062 606218 29146 606454
rect 29382 606218 29414 606454
rect 28794 606134 29414 606218
rect 28794 605898 28826 606134
rect 29062 605898 29146 606134
rect 29382 605898 29414 606134
rect 28794 570454 29414 605898
rect 28794 570218 28826 570454
rect 29062 570218 29146 570454
rect 29382 570218 29414 570454
rect 28794 570134 29414 570218
rect 28794 569898 28826 570134
rect 29062 569898 29146 570134
rect 29382 569898 29414 570134
rect 28794 534454 29414 569898
rect 28794 534218 28826 534454
rect 29062 534218 29146 534454
rect 29382 534218 29414 534454
rect 28794 534134 29414 534218
rect 28794 533898 28826 534134
rect 29062 533898 29146 534134
rect 29382 533898 29414 534134
rect 28794 498454 29414 533898
rect 28794 498218 28826 498454
rect 29062 498218 29146 498454
rect 29382 498218 29414 498454
rect 28794 498134 29414 498218
rect 28794 497898 28826 498134
rect 29062 497898 29146 498134
rect 29382 497898 29414 498134
rect 28794 462454 29414 497898
rect 28794 462218 28826 462454
rect 29062 462218 29146 462454
rect 29382 462218 29414 462454
rect 28794 462134 29414 462218
rect 28794 461898 28826 462134
rect 29062 461898 29146 462134
rect 29382 461898 29414 462134
rect 28794 426454 29414 461898
rect 28794 426218 28826 426454
rect 29062 426218 29146 426454
rect 29382 426218 29414 426454
rect 28794 426134 29414 426218
rect 28794 425898 28826 426134
rect 29062 425898 29146 426134
rect 29382 425898 29414 426134
rect 28794 390454 29414 425898
rect 28794 390218 28826 390454
rect 29062 390218 29146 390454
rect 29382 390218 29414 390454
rect 28794 390134 29414 390218
rect 28794 389898 28826 390134
rect 29062 389898 29146 390134
rect 29382 389898 29414 390134
rect 28794 354454 29414 389898
rect 28794 354218 28826 354454
rect 29062 354218 29146 354454
rect 29382 354218 29414 354454
rect 28794 354134 29414 354218
rect 28794 353898 28826 354134
rect 29062 353898 29146 354134
rect 29382 353898 29414 354134
rect 28794 318454 29414 353898
rect 28794 318218 28826 318454
rect 29062 318218 29146 318454
rect 29382 318218 29414 318454
rect 28794 318134 29414 318218
rect 28794 317898 28826 318134
rect 29062 317898 29146 318134
rect 29382 317898 29414 318134
rect 28794 282454 29414 317898
rect 28794 282218 28826 282454
rect 29062 282218 29146 282454
rect 29382 282218 29414 282454
rect 28794 282134 29414 282218
rect 28794 281898 28826 282134
rect 29062 281898 29146 282134
rect 29382 281898 29414 282134
rect 28794 246454 29414 281898
rect 28794 246218 28826 246454
rect 29062 246218 29146 246454
rect 29382 246218 29414 246454
rect 28794 246134 29414 246218
rect 28794 245898 28826 246134
rect 29062 245898 29146 246134
rect 29382 245898 29414 246134
rect 28794 210454 29414 245898
rect 28794 210218 28826 210454
rect 29062 210218 29146 210454
rect 29382 210218 29414 210454
rect 28794 210134 29414 210218
rect 28794 209898 28826 210134
rect 29062 209898 29146 210134
rect 29382 209898 29414 210134
rect 28794 174454 29414 209898
rect 28794 174218 28826 174454
rect 29062 174218 29146 174454
rect 29382 174218 29414 174454
rect 28794 174134 29414 174218
rect 28794 173898 28826 174134
rect 29062 173898 29146 174134
rect 29382 173898 29414 174134
rect 28794 138454 29414 173898
rect 28794 138218 28826 138454
rect 29062 138218 29146 138454
rect 29382 138218 29414 138454
rect 28794 138134 29414 138218
rect 28794 137898 28826 138134
rect 29062 137898 29146 138134
rect 29382 137898 29414 138134
rect 28794 102454 29414 137898
rect 28794 102218 28826 102454
rect 29062 102218 29146 102454
rect 29382 102218 29414 102454
rect 28794 102134 29414 102218
rect 28794 101898 28826 102134
rect 29062 101898 29146 102134
rect 29382 101898 29414 102134
rect 28794 66454 29414 101898
rect 28794 66218 28826 66454
rect 29062 66218 29146 66454
rect 29382 66218 29414 66454
rect 28794 66134 29414 66218
rect 28794 65898 28826 66134
rect 29062 65898 29146 66134
rect 29382 65898 29414 66134
rect 28794 30454 29414 65898
rect 28794 30218 28826 30454
rect 29062 30218 29146 30454
rect 29382 30218 29414 30454
rect 28794 30134 29414 30218
rect 28794 29898 28826 30134
rect 29062 29898 29146 30134
rect 29382 29898 29414 30134
rect 28794 -6106 29414 29898
rect 28794 -6342 28826 -6106
rect 29062 -6342 29146 -6106
rect 29382 -6342 29414 -6106
rect 28794 -6426 29414 -6342
rect 28794 -6662 28826 -6426
rect 29062 -6662 29146 -6426
rect 29382 -6662 29414 -6426
rect 28794 -7654 29414 -6662
rect 33294 711558 33914 711590
rect 33294 711322 33326 711558
rect 33562 711322 33646 711558
rect 33882 711322 33914 711558
rect 33294 711238 33914 711322
rect 33294 711002 33326 711238
rect 33562 711002 33646 711238
rect 33882 711002 33914 711238
rect 33294 682954 33914 711002
rect 33294 682718 33326 682954
rect 33562 682718 33646 682954
rect 33882 682718 33914 682954
rect 33294 682634 33914 682718
rect 33294 682398 33326 682634
rect 33562 682398 33646 682634
rect 33882 682398 33914 682634
rect 33294 646954 33914 682398
rect 33294 646718 33326 646954
rect 33562 646718 33646 646954
rect 33882 646718 33914 646954
rect 33294 646634 33914 646718
rect 33294 646398 33326 646634
rect 33562 646398 33646 646634
rect 33882 646398 33914 646634
rect 33294 610954 33914 646398
rect 33294 610718 33326 610954
rect 33562 610718 33646 610954
rect 33882 610718 33914 610954
rect 33294 610634 33914 610718
rect 33294 610398 33326 610634
rect 33562 610398 33646 610634
rect 33882 610398 33914 610634
rect 33294 574954 33914 610398
rect 33294 574718 33326 574954
rect 33562 574718 33646 574954
rect 33882 574718 33914 574954
rect 33294 574634 33914 574718
rect 33294 574398 33326 574634
rect 33562 574398 33646 574634
rect 33882 574398 33914 574634
rect 33294 538954 33914 574398
rect 33294 538718 33326 538954
rect 33562 538718 33646 538954
rect 33882 538718 33914 538954
rect 33294 538634 33914 538718
rect 33294 538398 33326 538634
rect 33562 538398 33646 538634
rect 33882 538398 33914 538634
rect 33294 502954 33914 538398
rect 33294 502718 33326 502954
rect 33562 502718 33646 502954
rect 33882 502718 33914 502954
rect 33294 502634 33914 502718
rect 33294 502398 33326 502634
rect 33562 502398 33646 502634
rect 33882 502398 33914 502634
rect 33294 466954 33914 502398
rect 33294 466718 33326 466954
rect 33562 466718 33646 466954
rect 33882 466718 33914 466954
rect 33294 466634 33914 466718
rect 33294 466398 33326 466634
rect 33562 466398 33646 466634
rect 33882 466398 33914 466634
rect 33294 430954 33914 466398
rect 33294 430718 33326 430954
rect 33562 430718 33646 430954
rect 33882 430718 33914 430954
rect 33294 430634 33914 430718
rect 33294 430398 33326 430634
rect 33562 430398 33646 430634
rect 33882 430398 33914 430634
rect 33294 394954 33914 430398
rect 33294 394718 33326 394954
rect 33562 394718 33646 394954
rect 33882 394718 33914 394954
rect 33294 394634 33914 394718
rect 33294 394398 33326 394634
rect 33562 394398 33646 394634
rect 33882 394398 33914 394634
rect 33294 358954 33914 394398
rect 33294 358718 33326 358954
rect 33562 358718 33646 358954
rect 33882 358718 33914 358954
rect 33294 358634 33914 358718
rect 33294 358398 33326 358634
rect 33562 358398 33646 358634
rect 33882 358398 33914 358634
rect 33294 322954 33914 358398
rect 33294 322718 33326 322954
rect 33562 322718 33646 322954
rect 33882 322718 33914 322954
rect 33294 322634 33914 322718
rect 33294 322398 33326 322634
rect 33562 322398 33646 322634
rect 33882 322398 33914 322634
rect 33294 286954 33914 322398
rect 33294 286718 33326 286954
rect 33562 286718 33646 286954
rect 33882 286718 33914 286954
rect 33294 286634 33914 286718
rect 33294 286398 33326 286634
rect 33562 286398 33646 286634
rect 33882 286398 33914 286634
rect 33294 250954 33914 286398
rect 33294 250718 33326 250954
rect 33562 250718 33646 250954
rect 33882 250718 33914 250954
rect 33294 250634 33914 250718
rect 33294 250398 33326 250634
rect 33562 250398 33646 250634
rect 33882 250398 33914 250634
rect 33294 214954 33914 250398
rect 33294 214718 33326 214954
rect 33562 214718 33646 214954
rect 33882 214718 33914 214954
rect 33294 214634 33914 214718
rect 33294 214398 33326 214634
rect 33562 214398 33646 214634
rect 33882 214398 33914 214634
rect 33294 178954 33914 214398
rect 33294 178718 33326 178954
rect 33562 178718 33646 178954
rect 33882 178718 33914 178954
rect 33294 178634 33914 178718
rect 33294 178398 33326 178634
rect 33562 178398 33646 178634
rect 33882 178398 33914 178634
rect 33294 142954 33914 178398
rect 33294 142718 33326 142954
rect 33562 142718 33646 142954
rect 33882 142718 33914 142954
rect 33294 142634 33914 142718
rect 33294 142398 33326 142634
rect 33562 142398 33646 142634
rect 33882 142398 33914 142634
rect 33294 106954 33914 142398
rect 33294 106718 33326 106954
rect 33562 106718 33646 106954
rect 33882 106718 33914 106954
rect 33294 106634 33914 106718
rect 33294 106398 33326 106634
rect 33562 106398 33646 106634
rect 33882 106398 33914 106634
rect 33294 70954 33914 106398
rect 33294 70718 33326 70954
rect 33562 70718 33646 70954
rect 33882 70718 33914 70954
rect 33294 70634 33914 70718
rect 33294 70398 33326 70634
rect 33562 70398 33646 70634
rect 33882 70398 33914 70634
rect 33294 34954 33914 70398
rect 33294 34718 33326 34954
rect 33562 34718 33646 34954
rect 33882 34718 33914 34954
rect 33294 34634 33914 34718
rect 33294 34398 33326 34634
rect 33562 34398 33646 34634
rect 33882 34398 33914 34634
rect 33294 -7066 33914 34398
rect 33294 -7302 33326 -7066
rect 33562 -7302 33646 -7066
rect 33882 -7302 33914 -7066
rect 33294 -7386 33914 -7302
rect 33294 -7622 33326 -7386
rect 33562 -7622 33646 -7386
rect 33882 -7622 33914 -7386
rect 33294 -7654 33914 -7622
rect 37794 704838 38414 711590
rect 37794 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 38414 704838
rect 37794 704518 38414 704602
rect 37794 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 38414 704518
rect 37794 687454 38414 704282
rect 37794 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 38414 687454
rect 37794 687134 38414 687218
rect 37794 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 38414 687134
rect 37794 651454 38414 686898
rect 37794 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 38414 651454
rect 37794 651134 38414 651218
rect 37794 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 38414 651134
rect 37794 615454 38414 650898
rect 37794 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 38414 615454
rect 37794 615134 38414 615218
rect 37794 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 38414 615134
rect 37794 579454 38414 614898
rect 37794 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 38414 579454
rect 37794 579134 38414 579218
rect 37794 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 38414 579134
rect 37794 543454 38414 578898
rect 37794 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 38414 543454
rect 37794 543134 38414 543218
rect 37794 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 38414 543134
rect 37794 507454 38414 542898
rect 37794 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 38414 507454
rect 37794 507134 38414 507218
rect 37794 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 38414 507134
rect 37794 471454 38414 506898
rect 37794 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 38414 471454
rect 37794 471134 38414 471218
rect 37794 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 38414 471134
rect 37794 435454 38414 470898
rect 37794 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 38414 435454
rect 37794 435134 38414 435218
rect 37794 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 38414 435134
rect 37794 399454 38414 434898
rect 37794 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 38414 399454
rect 37794 399134 38414 399218
rect 37794 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 38414 399134
rect 37794 363454 38414 398898
rect 37794 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 38414 363454
rect 37794 363134 38414 363218
rect 37794 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 38414 363134
rect 37794 327454 38414 362898
rect 37794 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 38414 327454
rect 37794 327134 38414 327218
rect 37794 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 38414 327134
rect 37794 291454 38414 326898
rect 37794 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 38414 291454
rect 37794 291134 38414 291218
rect 37794 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 38414 291134
rect 37794 255454 38414 290898
rect 37794 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 38414 255454
rect 37794 255134 38414 255218
rect 37794 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 38414 255134
rect 37794 219454 38414 254898
rect 37794 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 38414 219454
rect 37794 219134 38414 219218
rect 37794 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 38414 219134
rect 37794 183454 38414 218898
rect 37794 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 38414 183454
rect 37794 183134 38414 183218
rect 37794 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 38414 183134
rect 37794 147454 38414 182898
rect 37794 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 38414 147454
rect 37794 147134 38414 147218
rect 37794 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 38414 147134
rect 37794 111454 38414 146898
rect 37794 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 38414 111454
rect 37794 111134 38414 111218
rect 37794 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 38414 111134
rect 37794 75454 38414 110898
rect 37794 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 38414 75454
rect 37794 75134 38414 75218
rect 37794 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 38414 75134
rect 37794 39454 38414 74898
rect 37794 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 38414 39454
rect 37794 39134 38414 39218
rect 37794 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 38414 39134
rect 37794 3454 38414 38898
rect 37794 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 38414 3454
rect 37794 3134 38414 3218
rect 37794 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 38414 3134
rect 37794 -346 38414 2898
rect 37794 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 38414 -346
rect 37794 -666 38414 -582
rect 37794 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 38414 -666
rect 37794 -7654 38414 -902
rect 42294 705798 42914 711590
rect 42294 705562 42326 705798
rect 42562 705562 42646 705798
rect 42882 705562 42914 705798
rect 42294 705478 42914 705562
rect 42294 705242 42326 705478
rect 42562 705242 42646 705478
rect 42882 705242 42914 705478
rect 42294 691954 42914 705242
rect 42294 691718 42326 691954
rect 42562 691718 42646 691954
rect 42882 691718 42914 691954
rect 42294 691634 42914 691718
rect 42294 691398 42326 691634
rect 42562 691398 42646 691634
rect 42882 691398 42914 691634
rect 42294 655954 42914 691398
rect 42294 655718 42326 655954
rect 42562 655718 42646 655954
rect 42882 655718 42914 655954
rect 42294 655634 42914 655718
rect 42294 655398 42326 655634
rect 42562 655398 42646 655634
rect 42882 655398 42914 655634
rect 42294 619954 42914 655398
rect 42294 619718 42326 619954
rect 42562 619718 42646 619954
rect 42882 619718 42914 619954
rect 42294 619634 42914 619718
rect 42294 619398 42326 619634
rect 42562 619398 42646 619634
rect 42882 619398 42914 619634
rect 42294 583954 42914 619398
rect 42294 583718 42326 583954
rect 42562 583718 42646 583954
rect 42882 583718 42914 583954
rect 42294 583634 42914 583718
rect 42294 583398 42326 583634
rect 42562 583398 42646 583634
rect 42882 583398 42914 583634
rect 42294 547954 42914 583398
rect 42294 547718 42326 547954
rect 42562 547718 42646 547954
rect 42882 547718 42914 547954
rect 42294 547634 42914 547718
rect 42294 547398 42326 547634
rect 42562 547398 42646 547634
rect 42882 547398 42914 547634
rect 42294 511954 42914 547398
rect 42294 511718 42326 511954
rect 42562 511718 42646 511954
rect 42882 511718 42914 511954
rect 42294 511634 42914 511718
rect 42294 511398 42326 511634
rect 42562 511398 42646 511634
rect 42882 511398 42914 511634
rect 42294 475954 42914 511398
rect 42294 475718 42326 475954
rect 42562 475718 42646 475954
rect 42882 475718 42914 475954
rect 42294 475634 42914 475718
rect 42294 475398 42326 475634
rect 42562 475398 42646 475634
rect 42882 475398 42914 475634
rect 42294 439954 42914 475398
rect 42294 439718 42326 439954
rect 42562 439718 42646 439954
rect 42882 439718 42914 439954
rect 42294 439634 42914 439718
rect 42294 439398 42326 439634
rect 42562 439398 42646 439634
rect 42882 439398 42914 439634
rect 42294 403954 42914 439398
rect 42294 403718 42326 403954
rect 42562 403718 42646 403954
rect 42882 403718 42914 403954
rect 42294 403634 42914 403718
rect 42294 403398 42326 403634
rect 42562 403398 42646 403634
rect 42882 403398 42914 403634
rect 42294 367954 42914 403398
rect 42294 367718 42326 367954
rect 42562 367718 42646 367954
rect 42882 367718 42914 367954
rect 42294 367634 42914 367718
rect 42294 367398 42326 367634
rect 42562 367398 42646 367634
rect 42882 367398 42914 367634
rect 42294 331954 42914 367398
rect 42294 331718 42326 331954
rect 42562 331718 42646 331954
rect 42882 331718 42914 331954
rect 42294 331634 42914 331718
rect 42294 331398 42326 331634
rect 42562 331398 42646 331634
rect 42882 331398 42914 331634
rect 42294 295954 42914 331398
rect 42294 295718 42326 295954
rect 42562 295718 42646 295954
rect 42882 295718 42914 295954
rect 42294 295634 42914 295718
rect 42294 295398 42326 295634
rect 42562 295398 42646 295634
rect 42882 295398 42914 295634
rect 42294 259954 42914 295398
rect 42294 259718 42326 259954
rect 42562 259718 42646 259954
rect 42882 259718 42914 259954
rect 42294 259634 42914 259718
rect 42294 259398 42326 259634
rect 42562 259398 42646 259634
rect 42882 259398 42914 259634
rect 42294 223954 42914 259398
rect 42294 223718 42326 223954
rect 42562 223718 42646 223954
rect 42882 223718 42914 223954
rect 42294 223634 42914 223718
rect 42294 223398 42326 223634
rect 42562 223398 42646 223634
rect 42882 223398 42914 223634
rect 42294 187954 42914 223398
rect 42294 187718 42326 187954
rect 42562 187718 42646 187954
rect 42882 187718 42914 187954
rect 42294 187634 42914 187718
rect 42294 187398 42326 187634
rect 42562 187398 42646 187634
rect 42882 187398 42914 187634
rect 42294 151954 42914 187398
rect 42294 151718 42326 151954
rect 42562 151718 42646 151954
rect 42882 151718 42914 151954
rect 42294 151634 42914 151718
rect 42294 151398 42326 151634
rect 42562 151398 42646 151634
rect 42882 151398 42914 151634
rect 42294 115954 42914 151398
rect 42294 115718 42326 115954
rect 42562 115718 42646 115954
rect 42882 115718 42914 115954
rect 42294 115634 42914 115718
rect 42294 115398 42326 115634
rect 42562 115398 42646 115634
rect 42882 115398 42914 115634
rect 42294 79954 42914 115398
rect 42294 79718 42326 79954
rect 42562 79718 42646 79954
rect 42882 79718 42914 79954
rect 42294 79634 42914 79718
rect 42294 79398 42326 79634
rect 42562 79398 42646 79634
rect 42882 79398 42914 79634
rect 42294 43954 42914 79398
rect 42294 43718 42326 43954
rect 42562 43718 42646 43954
rect 42882 43718 42914 43954
rect 42294 43634 42914 43718
rect 42294 43398 42326 43634
rect 42562 43398 42646 43634
rect 42882 43398 42914 43634
rect 42294 7954 42914 43398
rect 42294 7718 42326 7954
rect 42562 7718 42646 7954
rect 42882 7718 42914 7954
rect 42294 7634 42914 7718
rect 42294 7398 42326 7634
rect 42562 7398 42646 7634
rect 42882 7398 42914 7634
rect 42294 -1306 42914 7398
rect 42294 -1542 42326 -1306
rect 42562 -1542 42646 -1306
rect 42882 -1542 42914 -1306
rect 42294 -1626 42914 -1542
rect 42294 -1862 42326 -1626
rect 42562 -1862 42646 -1626
rect 42882 -1862 42914 -1626
rect 42294 -7654 42914 -1862
rect 46794 706758 47414 711590
rect 46794 706522 46826 706758
rect 47062 706522 47146 706758
rect 47382 706522 47414 706758
rect 46794 706438 47414 706522
rect 46794 706202 46826 706438
rect 47062 706202 47146 706438
rect 47382 706202 47414 706438
rect 46794 696454 47414 706202
rect 46794 696218 46826 696454
rect 47062 696218 47146 696454
rect 47382 696218 47414 696454
rect 46794 696134 47414 696218
rect 46794 695898 46826 696134
rect 47062 695898 47146 696134
rect 47382 695898 47414 696134
rect 46794 660454 47414 695898
rect 46794 660218 46826 660454
rect 47062 660218 47146 660454
rect 47382 660218 47414 660454
rect 46794 660134 47414 660218
rect 46794 659898 46826 660134
rect 47062 659898 47146 660134
rect 47382 659898 47414 660134
rect 46794 624454 47414 659898
rect 46794 624218 46826 624454
rect 47062 624218 47146 624454
rect 47382 624218 47414 624454
rect 46794 624134 47414 624218
rect 46794 623898 46826 624134
rect 47062 623898 47146 624134
rect 47382 623898 47414 624134
rect 46794 588454 47414 623898
rect 46794 588218 46826 588454
rect 47062 588218 47146 588454
rect 47382 588218 47414 588454
rect 46794 588134 47414 588218
rect 46794 587898 46826 588134
rect 47062 587898 47146 588134
rect 47382 587898 47414 588134
rect 46794 552454 47414 587898
rect 46794 552218 46826 552454
rect 47062 552218 47146 552454
rect 47382 552218 47414 552454
rect 46794 552134 47414 552218
rect 46794 551898 46826 552134
rect 47062 551898 47146 552134
rect 47382 551898 47414 552134
rect 46794 516454 47414 551898
rect 46794 516218 46826 516454
rect 47062 516218 47146 516454
rect 47382 516218 47414 516454
rect 46794 516134 47414 516218
rect 46794 515898 46826 516134
rect 47062 515898 47146 516134
rect 47382 515898 47414 516134
rect 46794 480454 47414 515898
rect 46794 480218 46826 480454
rect 47062 480218 47146 480454
rect 47382 480218 47414 480454
rect 46794 480134 47414 480218
rect 46794 479898 46826 480134
rect 47062 479898 47146 480134
rect 47382 479898 47414 480134
rect 46794 444454 47414 479898
rect 46794 444218 46826 444454
rect 47062 444218 47146 444454
rect 47382 444218 47414 444454
rect 46794 444134 47414 444218
rect 46794 443898 46826 444134
rect 47062 443898 47146 444134
rect 47382 443898 47414 444134
rect 46794 408454 47414 443898
rect 46794 408218 46826 408454
rect 47062 408218 47146 408454
rect 47382 408218 47414 408454
rect 46794 408134 47414 408218
rect 46794 407898 46826 408134
rect 47062 407898 47146 408134
rect 47382 407898 47414 408134
rect 46794 372454 47414 407898
rect 46794 372218 46826 372454
rect 47062 372218 47146 372454
rect 47382 372218 47414 372454
rect 46794 372134 47414 372218
rect 46794 371898 46826 372134
rect 47062 371898 47146 372134
rect 47382 371898 47414 372134
rect 46794 336454 47414 371898
rect 46794 336218 46826 336454
rect 47062 336218 47146 336454
rect 47382 336218 47414 336454
rect 46794 336134 47414 336218
rect 46794 335898 46826 336134
rect 47062 335898 47146 336134
rect 47382 335898 47414 336134
rect 46794 300454 47414 335898
rect 46794 300218 46826 300454
rect 47062 300218 47146 300454
rect 47382 300218 47414 300454
rect 46794 300134 47414 300218
rect 46794 299898 46826 300134
rect 47062 299898 47146 300134
rect 47382 299898 47414 300134
rect 46794 264454 47414 299898
rect 46794 264218 46826 264454
rect 47062 264218 47146 264454
rect 47382 264218 47414 264454
rect 46794 264134 47414 264218
rect 46794 263898 46826 264134
rect 47062 263898 47146 264134
rect 47382 263898 47414 264134
rect 46794 228454 47414 263898
rect 46794 228218 46826 228454
rect 47062 228218 47146 228454
rect 47382 228218 47414 228454
rect 46794 228134 47414 228218
rect 46794 227898 46826 228134
rect 47062 227898 47146 228134
rect 47382 227898 47414 228134
rect 46794 192454 47414 227898
rect 46794 192218 46826 192454
rect 47062 192218 47146 192454
rect 47382 192218 47414 192454
rect 46794 192134 47414 192218
rect 46794 191898 46826 192134
rect 47062 191898 47146 192134
rect 47382 191898 47414 192134
rect 46794 156454 47414 191898
rect 46794 156218 46826 156454
rect 47062 156218 47146 156454
rect 47382 156218 47414 156454
rect 46794 156134 47414 156218
rect 46794 155898 46826 156134
rect 47062 155898 47146 156134
rect 47382 155898 47414 156134
rect 46794 120454 47414 155898
rect 46794 120218 46826 120454
rect 47062 120218 47146 120454
rect 47382 120218 47414 120454
rect 46794 120134 47414 120218
rect 46794 119898 46826 120134
rect 47062 119898 47146 120134
rect 47382 119898 47414 120134
rect 46794 84454 47414 119898
rect 46794 84218 46826 84454
rect 47062 84218 47146 84454
rect 47382 84218 47414 84454
rect 46794 84134 47414 84218
rect 46794 83898 46826 84134
rect 47062 83898 47146 84134
rect 47382 83898 47414 84134
rect 46794 48454 47414 83898
rect 46794 48218 46826 48454
rect 47062 48218 47146 48454
rect 47382 48218 47414 48454
rect 46794 48134 47414 48218
rect 46794 47898 46826 48134
rect 47062 47898 47146 48134
rect 47382 47898 47414 48134
rect 46794 12454 47414 47898
rect 46794 12218 46826 12454
rect 47062 12218 47146 12454
rect 47382 12218 47414 12454
rect 46794 12134 47414 12218
rect 46794 11898 46826 12134
rect 47062 11898 47146 12134
rect 47382 11898 47414 12134
rect 46794 -2266 47414 11898
rect 46794 -2502 46826 -2266
rect 47062 -2502 47146 -2266
rect 47382 -2502 47414 -2266
rect 46794 -2586 47414 -2502
rect 46794 -2822 46826 -2586
rect 47062 -2822 47146 -2586
rect 47382 -2822 47414 -2586
rect 46794 -7654 47414 -2822
rect 51294 707718 51914 711590
rect 51294 707482 51326 707718
rect 51562 707482 51646 707718
rect 51882 707482 51914 707718
rect 51294 707398 51914 707482
rect 51294 707162 51326 707398
rect 51562 707162 51646 707398
rect 51882 707162 51914 707398
rect 51294 700954 51914 707162
rect 51294 700718 51326 700954
rect 51562 700718 51646 700954
rect 51882 700718 51914 700954
rect 51294 700634 51914 700718
rect 51294 700398 51326 700634
rect 51562 700398 51646 700634
rect 51882 700398 51914 700634
rect 51294 664954 51914 700398
rect 51294 664718 51326 664954
rect 51562 664718 51646 664954
rect 51882 664718 51914 664954
rect 51294 664634 51914 664718
rect 51294 664398 51326 664634
rect 51562 664398 51646 664634
rect 51882 664398 51914 664634
rect 51294 628954 51914 664398
rect 51294 628718 51326 628954
rect 51562 628718 51646 628954
rect 51882 628718 51914 628954
rect 51294 628634 51914 628718
rect 51294 628398 51326 628634
rect 51562 628398 51646 628634
rect 51882 628398 51914 628634
rect 51294 592954 51914 628398
rect 51294 592718 51326 592954
rect 51562 592718 51646 592954
rect 51882 592718 51914 592954
rect 51294 592634 51914 592718
rect 51294 592398 51326 592634
rect 51562 592398 51646 592634
rect 51882 592398 51914 592634
rect 51294 556954 51914 592398
rect 51294 556718 51326 556954
rect 51562 556718 51646 556954
rect 51882 556718 51914 556954
rect 51294 556634 51914 556718
rect 51294 556398 51326 556634
rect 51562 556398 51646 556634
rect 51882 556398 51914 556634
rect 51294 520954 51914 556398
rect 51294 520718 51326 520954
rect 51562 520718 51646 520954
rect 51882 520718 51914 520954
rect 51294 520634 51914 520718
rect 51294 520398 51326 520634
rect 51562 520398 51646 520634
rect 51882 520398 51914 520634
rect 51294 484954 51914 520398
rect 51294 484718 51326 484954
rect 51562 484718 51646 484954
rect 51882 484718 51914 484954
rect 51294 484634 51914 484718
rect 51294 484398 51326 484634
rect 51562 484398 51646 484634
rect 51882 484398 51914 484634
rect 51294 448954 51914 484398
rect 51294 448718 51326 448954
rect 51562 448718 51646 448954
rect 51882 448718 51914 448954
rect 51294 448634 51914 448718
rect 51294 448398 51326 448634
rect 51562 448398 51646 448634
rect 51882 448398 51914 448634
rect 51294 412954 51914 448398
rect 51294 412718 51326 412954
rect 51562 412718 51646 412954
rect 51882 412718 51914 412954
rect 51294 412634 51914 412718
rect 51294 412398 51326 412634
rect 51562 412398 51646 412634
rect 51882 412398 51914 412634
rect 51294 376954 51914 412398
rect 51294 376718 51326 376954
rect 51562 376718 51646 376954
rect 51882 376718 51914 376954
rect 51294 376634 51914 376718
rect 51294 376398 51326 376634
rect 51562 376398 51646 376634
rect 51882 376398 51914 376634
rect 51294 340954 51914 376398
rect 51294 340718 51326 340954
rect 51562 340718 51646 340954
rect 51882 340718 51914 340954
rect 51294 340634 51914 340718
rect 51294 340398 51326 340634
rect 51562 340398 51646 340634
rect 51882 340398 51914 340634
rect 51294 304954 51914 340398
rect 51294 304718 51326 304954
rect 51562 304718 51646 304954
rect 51882 304718 51914 304954
rect 51294 304634 51914 304718
rect 51294 304398 51326 304634
rect 51562 304398 51646 304634
rect 51882 304398 51914 304634
rect 51294 268954 51914 304398
rect 51294 268718 51326 268954
rect 51562 268718 51646 268954
rect 51882 268718 51914 268954
rect 51294 268634 51914 268718
rect 51294 268398 51326 268634
rect 51562 268398 51646 268634
rect 51882 268398 51914 268634
rect 51294 232954 51914 268398
rect 51294 232718 51326 232954
rect 51562 232718 51646 232954
rect 51882 232718 51914 232954
rect 51294 232634 51914 232718
rect 51294 232398 51326 232634
rect 51562 232398 51646 232634
rect 51882 232398 51914 232634
rect 51294 196954 51914 232398
rect 51294 196718 51326 196954
rect 51562 196718 51646 196954
rect 51882 196718 51914 196954
rect 51294 196634 51914 196718
rect 51294 196398 51326 196634
rect 51562 196398 51646 196634
rect 51882 196398 51914 196634
rect 51294 160954 51914 196398
rect 51294 160718 51326 160954
rect 51562 160718 51646 160954
rect 51882 160718 51914 160954
rect 51294 160634 51914 160718
rect 51294 160398 51326 160634
rect 51562 160398 51646 160634
rect 51882 160398 51914 160634
rect 51294 124954 51914 160398
rect 51294 124718 51326 124954
rect 51562 124718 51646 124954
rect 51882 124718 51914 124954
rect 51294 124634 51914 124718
rect 51294 124398 51326 124634
rect 51562 124398 51646 124634
rect 51882 124398 51914 124634
rect 51294 88954 51914 124398
rect 51294 88718 51326 88954
rect 51562 88718 51646 88954
rect 51882 88718 51914 88954
rect 51294 88634 51914 88718
rect 51294 88398 51326 88634
rect 51562 88398 51646 88634
rect 51882 88398 51914 88634
rect 51294 52954 51914 88398
rect 51294 52718 51326 52954
rect 51562 52718 51646 52954
rect 51882 52718 51914 52954
rect 51294 52634 51914 52718
rect 51294 52398 51326 52634
rect 51562 52398 51646 52634
rect 51882 52398 51914 52634
rect 51294 16954 51914 52398
rect 51294 16718 51326 16954
rect 51562 16718 51646 16954
rect 51882 16718 51914 16954
rect 51294 16634 51914 16718
rect 51294 16398 51326 16634
rect 51562 16398 51646 16634
rect 51882 16398 51914 16634
rect 51294 -3226 51914 16398
rect 51294 -3462 51326 -3226
rect 51562 -3462 51646 -3226
rect 51882 -3462 51914 -3226
rect 51294 -3546 51914 -3462
rect 51294 -3782 51326 -3546
rect 51562 -3782 51646 -3546
rect 51882 -3782 51914 -3546
rect 51294 -7654 51914 -3782
rect 55794 708678 56414 711590
rect 55794 708442 55826 708678
rect 56062 708442 56146 708678
rect 56382 708442 56414 708678
rect 55794 708358 56414 708442
rect 55794 708122 55826 708358
rect 56062 708122 56146 708358
rect 56382 708122 56414 708358
rect 55794 669454 56414 708122
rect 55794 669218 55826 669454
rect 56062 669218 56146 669454
rect 56382 669218 56414 669454
rect 55794 669134 56414 669218
rect 55794 668898 55826 669134
rect 56062 668898 56146 669134
rect 56382 668898 56414 669134
rect 55794 633454 56414 668898
rect 55794 633218 55826 633454
rect 56062 633218 56146 633454
rect 56382 633218 56414 633454
rect 55794 633134 56414 633218
rect 55794 632898 55826 633134
rect 56062 632898 56146 633134
rect 56382 632898 56414 633134
rect 55794 597454 56414 632898
rect 55794 597218 55826 597454
rect 56062 597218 56146 597454
rect 56382 597218 56414 597454
rect 55794 597134 56414 597218
rect 55794 596898 55826 597134
rect 56062 596898 56146 597134
rect 56382 596898 56414 597134
rect 55794 561454 56414 596898
rect 55794 561218 55826 561454
rect 56062 561218 56146 561454
rect 56382 561218 56414 561454
rect 55794 561134 56414 561218
rect 55794 560898 55826 561134
rect 56062 560898 56146 561134
rect 56382 560898 56414 561134
rect 55794 525454 56414 560898
rect 55794 525218 55826 525454
rect 56062 525218 56146 525454
rect 56382 525218 56414 525454
rect 55794 525134 56414 525218
rect 55794 524898 55826 525134
rect 56062 524898 56146 525134
rect 56382 524898 56414 525134
rect 55794 489454 56414 524898
rect 55794 489218 55826 489454
rect 56062 489218 56146 489454
rect 56382 489218 56414 489454
rect 55794 489134 56414 489218
rect 55794 488898 55826 489134
rect 56062 488898 56146 489134
rect 56382 488898 56414 489134
rect 55794 453454 56414 488898
rect 55794 453218 55826 453454
rect 56062 453218 56146 453454
rect 56382 453218 56414 453454
rect 55794 453134 56414 453218
rect 55794 452898 55826 453134
rect 56062 452898 56146 453134
rect 56382 452898 56414 453134
rect 55794 417454 56414 452898
rect 55794 417218 55826 417454
rect 56062 417218 56146 417454
rect 56382 417218 56414 417454
rect 55794 417134 56414 417218
rect 55794 416898 55826 417134
rect 56062 416898 56146 417134
rect 56382 416898 56414 417134
rect 55794 381454 56414 416898
rect 55794 381218 55826 381454
rect 56062 381218 56146 381454
rect 56382 381218 56414 381454
rect 55794 381134 56414 381218
rect 55794 380898 55826 381134
rect 56062 380898 56146 381134
rect 56382 380898 56414 381134
rect 55794 345454 56414 380898
rect 55794 345218 55826 345454
rect 56062 345218 56146 345454
rect 56382 345218 56414 345454
rect 55794 345134 56414 345218
rect 55794 344898 55826 345134
rect 56062 344898 56146 345134
rect 56382 344898 56414 345134
rect 55794 309454 56414 344898
rect 55794 309218 55826 309454
rect 56062 309218 56146 309454
rect 56382 309218 56414 309454
rect 55794 309134 56414 309218
rect 55794 308898 55826 309134
rect 56062 308898 56146 309134
rect 56382 308898 56414 309134
rect 55794 273454 56414 308898
rect 55794 273218 55826 273454
rect 56062 273218 56146 273454
rect 56382 273218 56414 273454
rect 55794 273134 56414 273218
rect 55794 272898 55826 273134
rect 56062 272898 56146 273134
rect 56382 272898 56414 273134
rect 55794 237454 56414 272898
rect 55794 237218 55826 237454
rect 56062 237218 56146 237454
rect 56382 237218 56414 237454
rect 55794 237134 56414 237218
rect 55794 236898 55826 237134
rect 56062 236898 56146 237134
rect 56382 236898 56414 237134
rect 55794 201454 56414 236898
rect 55794 201218 55826 201454
rect 56062 201218 56146 201454
rect 56382 201218 56414 201454
rect 55794 201134 56414 201218
rect 55794 200898 55826 201134
rect 56062 200898 56146 201134
rect 56382 200898 56414 201134
rect 55794 165454 56414 200898
rect 55794 165218 55826 165454
rect 56062 165218 56146 165454
rect 56382 165218 56414 165454
rect 55794 165134 56414 165218
rect 55794 164898 55826 165134
rect 56062 164898 56146 165134
rect 56382 164898 56414 165134
rect 55794 129454 56414 164898
rect 55794 129218 55826 129454
rect 56062 129218 56146 129454
rect 56382 129218 56414 129454
rect 55794 129134 56414 129218
rect 55794 128898 55826 129134
rect 56062 128898 56146 129134
rect 56382 128898 56414 129134
rect 55794 93454 56414 128898
rect 55794 93218 55826 93454
rect 56062 93218 56146 93454
rect 56382 93218 56414 93454
rect 55794 93134 56414 93218
rect 55794 92898 55826 93134
rect 56062 92898 56146 93134
rect 56382 92898 56414 93134
rect 55794 57454 56414 92898
rect 55794 57218 55826 57454
rect 56062 57218 56146 57454
rect 56382 57218 56414 57454
rect 55794 57134 56414 57218
rect 55794 56898 55826 57134
rect 56062 56898 56146 57134
rect 56382 56898 56414 57134
rect 55794 21454 56414 56898
rect 55794 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 56414 21454
rect 55794 21134 56414 21218
rect 55794 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 56414 21134
rect 55794 -4186 56414 20898
rect 55794 -4422 55826 -4186
rect 56062 -4422 56146 -4186
rect 56382 -4422 56414 -4186
rect 55794 -4506 56414 -4422
rect 55794 -4742 55826 -4506
rect 56062 -4742 56146 -4506
rect 56382 -4742 56414 -4506
rect 55794 -7654 56414 -4742
rect 60294 709638 60914 711590
rect 60294 709402 60326 709638
rect 60562 709402 60646 709638
rect 60882 709402 60914 709638
rect 60294 709318 60914 709402
rect 60294 709082 60326 709318
rect 60562 709082 60646 709318
rect 60882 709082 60914 709318
rect 60294 673954 60914 709082
rect 60294 673718 60326 673954
rect 60562 673718 60646 673954
rect 60882 673718 60914 673954
rect 60294 673634 60914 673718
rect 60294 673398 60326 673634
rect 60562 673398 60646 673634
rect 60882 673398 60914 673634
rect 60294 637954 60914 673398
rect 60294 637718 60326 637954
rect 60562 637718 60646 637954
rect 60882 637718 60914 637954
rect 60294 637634 60914 637718
rect 60294 637398 60326 637634
rect 60562 637398 60646 637634
rect 60882 637398 60914 637634
rect 60294 601954 60914 637398
rect 60294 601718 60326 601954
rect 60562 601718 60646 601954
rect 60882 601718 60914 601954
rect 60294 601634 60914 601718
rect 60294 601398 60326 601634
rect 60562 601398 60646 601634
rect 60882 601398 60914 601634
rect 60294 565954 60914 601398
rect 60294 565718 60326 565954
rect 60562 565718 60646 565954
rect 60882 565718 60914 565954
rect 60294 565634 60914 565718
rect 60294 565398 60326 565634
rect 60562 565398 60646 565634
rect 60882 565398 60914 565634
rect 60294 529954 60914 565398
rect 60294 529718 60326 529954
rect 60562 529718 60646 529954
rect 60882 529718 60914 529954
rect 60294 529634 60914 529718
rect 60294 529398 60326 529634
rect 60562 529398 60646 529634
rect 60882 529398 60914 529634
rect 60294 493954 60914 529398
rect 60294 493718 60326 493954
rect 60562 493718 60646 493954
rect 60882 493718 60914 493954
rect 60294 493634 60914 493718
rect 60294 493398 60326 493634
rect 60562 493398 60646 493634
rect 60882 493398 60914 493634
rect 60294 457954 60914 493398
rect 60294 457718 60326 457954
rect 60562 457718 60646 457954
rect 60882 457718 60914 457954
rect 60294 457634 60914 457718
rect 60294 457398 60326 457634
rect 60562 457398 60646 457634
rect 60882 457398 60914 457634
rect 60294 421954 60914 457398
rect 60294 421718 60326 421954
rect 60562 421718 60646 421954
rect 60882 421718 60914 421954
rect 60294 421634 60914 421718
rect 60294 421398 60326 421634
rect 60562 421398 60646 421634
rect 60882 421398 60914 421634
rect 60294 385954 60914 421398
rect 60294 385718 60326 385954
rect 60562 385718 60646 385954
rect 60882 385718 60914 385954
rect 60294 385634 60914 385718
rect 60294 385398 60326 385634
rect 60562 385398 60646 385634
rect 60882 385398 60914 385634
rect 60294 349954 60914 385398
rect 60294 349718 60326 349954
rect 60562 349718 60646 349954
rect 60882 349718 60914 349954
rect 60294 349634 60914 349718
rect 60294 349398 60326 349634
rect 60562 349398 60646 349634
rect 60882 349398 60914 349634
rect 60294 313954 60914 349398
rect 60294 313718 60326 313954
rect 60562 313718 60646 313954
rect 60882 313718 60914 313954
rect 60294 313634 60914 313718
rect 60294 313398 60326 313634
rect 60562 313398 60646 313634
rect 60882 313398 60914 313634
rect 60294 277954 60914 313398
rect 60294 277718 60326 277954
rect 60562 277718 60646 277954
rect 60882 277718 60914 277954
rect 60294 277634 60914 277718
rect 60294 277398 60326 277634
rect 60562 277398 60646 277634
rect 60882 277398 60914 277634
rect 60294 241954 60914 277398
rect 60294 241718 60326 241954
rect 60562 241718 60646 241954
rect 60882 241718 60914 241954
rect 60294 241634 60914 241718
rect 60294 241398 60326 241634
rect 60562 241398 60646 241634
rect 60882 241398 60914 241634
rect 60294 205954 60914 241398
rect 60294 205718 60326 205954
rect 60562 205718 60646 205954
rect 60882 205718 60914 205954
rect 60294 205634 60914 205718
rect 60294 205398 60326 205634
rect 60562 205398 60646 205634
rect 60882 205398 60914 205634
rect 60294 169954 60914 205398
rect 60294 169718 60326 169954
rect 60562 169718 60646 169954
rect 60882 169718 60914 169954
rect 60294 169634 60914 169718
rect 60294 169398 60326 169634
rect 60562 169398 60646 169634
rect 60882 169398 60914 169634
rect 60294 133954 60914 169398
rect 60294 133718 60326 133954
rect 60562 133718 60646 133954
rect 60882 133718 60914 133954
rect 60294 133634 60914 133718
rect 60294 133398 60326 133634
rect 60562 133398 60646 133634
rect 60882 133398 60914 133634
rect 60294 97954 60914 133398
rect 60294 97718 60326 97954
rect 60562 97718 60646 97954
rect 60882 97718 60914 97954
rect 60294 97634 60914 97718
rect 60294 97398 60326 97634
rect 60562 97398 60646 97634
rect 60882 97398 60914 97634
rect 60294 61954 60914 97398
rect 60294 61718 60326 61954
rect 60562 61718 60646 61954
rect 60882 61718 60914 61954
rect 60294 61634 60914 61718
rect 60294 61398 60326 61634
rect 60562 61398 60646 61634
rect 60882 61398 60914 61634
rect 60294 25954 60914 61398
rect 60294 25718 60326 25954
rect 60562 25718 60646 25954
rect 60882 25718 60914 25954
rect 60294 25634 60914 25718
rect 60294 25398 60326 25634
rect 60562 25398 60646 25634
rect 60882 25398 60914 25634
rect 60294 -5146 60914 25398
rect 60294 -5382 60326 -5146
rect 60562 -5382 60646 -5146
rect 60882 -5382 60914 -5146
rect 60294 -5466 60914 -5382
rect 60294 -5702 60326 -5466
rect 60562 -5702 60646 -5466
rect 60882 -5702 60914 -5466
rect 60294 -7654 60914 -5702
rect 64794 710598 65414 711590
rect 64794 710362 64826 710598
rect 65062 710362 65146 710598
rect 65382 710362 65414 710598
rect 64794 710278 65414 710362
rect 64794 710042 64826 710278
rect 65062 710042 65146 710278
rect 65382 710042 65414 710278
rect 64794 678454 65414 710042
rect 64794 678218 64826 678454
rect 65062 678218 65146 678454
rect 65382 678218 65414 678454
rect 64794 678134 65414 678218
rect 64794 677898 64826 678134
rect 65062 677898 65146 678134
rect 65382 677898 65414 678134
rect 64794 642454 65414 677898
rect 64794 642218 64826 642454
rect 65062 642218 65146 642454
rect 65382 642218 65414 642454
rect 64794 642134 65414 642218
rect 64794 641898 64826 642134
rect 65062 641898 65146 642134
rect 65382 641898 65414 642134
rect 64794 606454 65414 641898
rect 64794 606218 64826 606454
rect 65062 606218 65146 606454
rect 65382 606218 65414 606454
rect 64794 606134 65414 606218
rect 64794 605898 64826 606134
rect 65062 605898 65146 606134
rect 65382 605898 65414 606134
rect 64794 570454 65414 605898
rect 64794 570218 64826 570454
rect 65062 570218 65146 570454
rect 65382 570218 65414 570454
rect 64794 570134 65414 570218
rect 64794 569898 64826 570134
rect 65062 569898 65146 570134
rect 65382 569898 65414 570134
rect 64794 534454 65414 569898
rect 64794 534218 64826 534454
rect 65062 534218 65146 534454
rect 65382 534218 65414 534454
rect 64794 534134 65414 534218
rect 64794 533898 64826 534134
rect 65062 533898 65146 534134
rect 65382 533898 65414 534134
rect 64794 498454 65414 533898
rect 64794 498218 64826 498454
rect 65062 498218 65146 498454
rect 65382 498218 65414 498454
rect 64794 498134 65414 498218
rect 64794 497898 64826 498134
rect 65062 497898 65146 498134
rect 65382 497898 65414 498134
rect 64794 462454 65414 497898
rect 64794 462218 64826 462454
rect 65062 462218 65146 462454
rect 65382 462218 65414 462454
rect 64794 462134 65414 462218
rect 64794 461898 64826 462134
rect 65062 461898 65146 462134
rect 65382 461898 65414 462134
rect 64794 426454 65414 461898
rect 64794 426218 64826 426454
rect 65062 426218 65146 426454
rect 65382 426218 65414 426454
rect 64794 426134 65414 426218
rect 64794 425898 64826 426134
rect 65062 425898 65146 426134
rect 65382 425898 65414 426134
rect 64794 390454 65414 425898
rect 64794 390218 64826 390454
rect 65062 390218 65146 390454
rect 65382 390218 65414 390454
rect 64794 390134 65414 390218
rect 64794 389898 64826 390134
rect 65062 389898 65146 390134
rect 65382 389898 65414 390134
rect 64794 354454 65414 389898
rect 64794 354218 64826 354454
rect 65062 354218 65146 354454
rect 65382 354218 65414 354454
rect 64794 354134 65414 354218
rect 64794 353898 64826 354134
rect 65062 353898 65146 354134
rect 65382 353898 65414 354134
rect 64794 318454 65414 353898
rect 64794 318218 64826 318454
rect 65062 318218 65146 318454
rect 65382 318218 65414 318454
rect 64794 318134 65414 318218
rect 64794 317898 64826 318134
rect 65062 317898 65146 318134
rect 65382 317898 65414 318134
rect 64794 282454 65414 317898
rect 64794 282218 64826 282454
rect 65062 282218 65146 282454
rect 65382 282218 65414 282454
rect 64794 282134 65414 282218
rect 64794 281898 64826 282134
rect 65062 281898 65146 282134
rect 65382 281898 65414 282134
rect 64794 246454 65414 281898
rect 64794 246218 64826 246454
rect 65062 246218 65146 246454
rect 65382 246218 65414 246454
rect 64794 246134 65414 246218
rect 64794 245898 64826 246134
rect 65062 245898 65146 246134
rect 65382 245898 65414 246134
rect 64794 210454 65414 245898
rect 64794 210218 64826 210454
rect 65062 210218 65146 210454
rect 65382 210218 65414 210454
rect 64794 210134 65414 210218
rect 64794 209898 64826 210134
rect 65062 209898 65146 210134
rect 65382 209898 65414 210134
rect 64794 174454 65414 209898
rect 64794 174218 64826 174454
rect 65062 174218 65146 174454
rect 65382 174218 65414 174454
rect 64794 174134 65414 174218
rect 64794 173898 64826 174134
rect 65062 173898 65146 174134
rect 65382 173898 65414 174134
rect 64794 138454 65414 173898
rect 64794 138218 64826 138454
rect 65062 138218 65146 138454
rect 65382 138218 65414 138454
rect 64794 138134 65414 138218
rect 64794 137898 64826 138134
rect 65062 137898 65146 138134
rect 65382 137898 65414 138134
rect 64794 102454 65414 137898
rect 64794 102218 64826 102454
rect 65062 102218 65146 102454
rect 65382 102218 65414 102454
rect 64794 102134 65414 102218
rect 64794 101898 64826 102134
rect 65062 101898 65146 102134
rect 65382 101898 65414 102134
rect 64794 66454 65414 101898
rect 64794 66218 64826 66454
rect 65062 66218 65146 66454
rect 65382 66218 65414 66454
rect 64794 66134 65414 66218
rect 64794 65898 64826 66134
rect 65062 65898 65146 66134
rect 65382 65898 65414 66134
rect 64794 30454 65414 65898
rect 64794 30218 64826 30454
rect 65062 30218 65146 30454
rect 65382 30218 65414 30454
rect 64794 30134 65414 30218
rect 64794 29898 64826 30134
rect 65062 29898 65146 30134
rect 65382 29898 65414 30134
rect 64794 -6106 65414 29898
rect 64794 -6342 64826 -6106
rect 65062 -6342 65146 -6106
rect 65382 -6342 65414 -6106
rect 64794 -6426 65414 -6342
rect 64794 -6662 64826 -6426
rect 65062 -6662 65146 -6426
rect 65382 -6662 65414 -6426
rect 64794 -7654 65414 -6662
rect 69294 711558 69914 711590
rect 69294 711322 69326 711558
rect 69562 711322 69646 711558
rect 69882 711322 69914 711558
rect 69294 711238 69914 711322
rect 69294 711002 69326 711238
rect 69562 711002 69646 711238
rect 69882 711002 69914 711238
rect 69294 682954 69914 711002
rect 69294 682718 69326 682954
rect 69562 682718 69646 682954
rect 69882 682718 69914 682954
rect 69294 682634 69914 682718
rect 69294 682398 69326 682634
rect 69562 682398 69646 682634
rect 69882 682398 69914 682634
rect 69294 646954 69914 682398
rect 69294 646718 69326 646954
rect 69562 646718 69646 646954
rect 69882 646718 69914 646954
rect 69294 646634 69914 646718
rect 69294 646398 69326 646634
rect 69562 646398 69646 646634
rect 69882 646398 69914 646634
rect 69294 610954 69914 646398
rect 69294 610718 69326 610954
rect 69562 610718 69646 610954
rect 69882 610718 69914 610954
rect 69294 610634 69914 610718
rect 69294 610398 69326 610634
rect 69562 610398 69646 610634
rect 69882 610398 69914 610634
rect 69294 574954 69914 610398
rect 69294 574718 69326 574954
rect 69562 574718 69646 574954
rect 69882 574718 69914 574954
rect 69294 574634 69914 574718
rect 69294 574398 69326 574634
rect 69562 574398 69646 574634
rect 69882 574398 69914 574634
rect 69294 538954 69914 574398
rect 69294 538718 69326 538954
rect 69562 538718 69646 538954
rect 69882 538718 69914 538954
rect 69294 538634 69914 538718
rect 69294 538398 69326 538634
rect 69562 538398 69646 538634
rect 69882 538398 69914 538634
rect 69294 502954 69914 538398
rect 69294 502718 69326 502954
rect 69562 502718 69646 502954
rect 69882 502718 69914 502954
rect 69294 502634 69914 502718
rect 69294 502398 69326 502634
rect 69562 502398 69646 502634
rect 69882 502398 69914 502634
rect 69294 466954 69914 502398
rect 69294 466718 69326 466954
rect 69562 466718 69646 466954
rect 69882 466718 69914 466954
rect 69294 466634 69914 466718
rect 69294 466398 69326 466634
rect 69562 466398 69646 466634
rect 69882 466398 69914 466634
rect 69294 430954 69914 466398
rect 69294 430718 69326 430954
rect 69562 430718 69646 430954
rect 69882 430718 69914 430954
rect 69294 430634 69914 430718
rect 69294 430398 69326 430634
rect 69562 430398 69646 430634
rect 69882 430398 69914 430634
rect 69294 394954 69914 430398
rect 69294 394718 69326 394954
rect 69562 394718 69646 394954
rect 69882 394718 69914 394954
rect 69294 394634 69914 394718
rect 69294 394398 69326 394634
rect 69562 394398 69646 394634
rect 69882 394398 69914 394634
rect 69294 358954 69914 394398
rect 69294 358718 69326 358954
rect 69562 358718 69646 358954
rect 69882 358718 69914 358954
rect 69294 358634 69914 358718
rect 69294 358398 69326 358634
rect 69562 358398 69646 358634
rect 69882 358398 69914 358634
rect 69294 322954 69914 358398
rect 69294 322718 69326 322954
rect 69562 322718 69646 322954
rect 69882 322718 69914 322954
rect 69294 322634 69914 322718
rect 69294 322398 69326 322634
rect 69562 322398 69646 322634
rect 69882 322398 69914 322634
rect 69294 286954 69914 322398
rect 69294 286718 69326 286954
rect 69562 286718 69646 286954
rect 69882 286718 69914 286954
rect 69294 286634 69914 286718
rect 69294 286398 69326 286634
rect 69562 286398 69646 286634
rect 69882 286398 69914 286634
rect 69294 250954 69914 286398
rect 69294 250718 69326 250954
rect 69562 250718 69646 250954
rect 69882 250718 69914 250954
rect 69294 250634 69914 250718
rect 69294 250398 69326 250634
rect 69562 250398 69646 250634
rect 69882 250398 69914 250634
rect 69294 214954 69914 250398
rect 69294 214718 69326 214954
rect 69562 214718 69646 214954
rect 69882 214718 69914 214954
rect 69294 214634 69914 214718
rect 69294 214398 69326 214634
rect 69562 214398 69646 214634
rect 69882 214398 69914 214634
rect 69294 178954 69914 214398
rect 69294 178718 69326 178954
rect 69562 178718 69646 178954
rect 69882 178718 69914 178954
rect 69294 178634 69914 178718
rect 69294 178398 69326 178634
rect 69562 178398 69646 178634
rect 69882 178398 69914 178634
rect 69294 142954 69914 178398
rect 69294 142718 69326 142954
rect 69562 142718 69646 142954
rect 69882 142718 69914 142954
rect 69294 142634 69914 142718
rect 69294 142398 69326 142634
rect 69562 142398 69646 142634
rect 69882 142398 69914 142634
rect 69294 106954 69914 142398
rect 69294 106718 69326 106954
rect 69562 106718 69646 106954
rect 69882 106718 69914 106954
rect 69294 106634 69914 106718
rect 69294 106398 69326 106634
rect 69562 106398 69646 106634
rect 69882 106398 69914 106634
rect 69294 70954 69914 106398
rect 69294 70718 69326 70954
rect 69562 70718 69646 70954
rect 69882 70718 69914 70954
rect 69294 70634 69914 70718
rect 69294 70398 69326 70634
rect 69562 70398 69646 70634
rect 69882 70398 69914 70634
rect 69294 34954 69914 70398
rect 69294 34718 69326 34954
rect 69562 34718 69646 34954
rect 69882 34718 69914 34954
rect 69294 34634 69914 34718
rect 69294 34398 69326 34634
rect 69562 34398 69646 34634
rect 69882 34398 69914 34634
rect 69294 -7066 69914 34398
rect 69294 -7302 69326 -7066
rect 69562 -7302 69646 -7066
rect 69882 -7302 69914 -7066
rect 69294 -7386 69914 -7302
rect 69294 -7622 69326 -7386
rect 69562 -7622 69646 -7386
rect 69882 -7622 69914 -7386
rect 69294 -7654 69914 -7622
rect 73794 704838 74414 711590
rect 73794 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 74414 704838
rect 73794 704518 74414 704602
rect 73794 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 74414 704518
rect 73794 687454 74414 704282
rect 73794 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 74414 687454
rect 73794 687134 74414 687218
rect 73794 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 74414 687134
rect 73794 651454 74414 686898
rect 73794 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 74414 651454
rect 73794 651134 74414 651218
rect 73794 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 74414 651134
rect 73794 615454 74414 650898
rect 73794 615218 73826 615454
rect 74062 615218 74146 615454
rect 74382 615218 74414 615454
rect 73794 615134 74414 615218
rect 73794 614898 73826 615134
rect 74062 614898 74146 615134
rect 74382 614898 74414 615134
rect 73794 579454 74414 614898
rect 73794 579218 73826 579454
rect 74062 579218 74146 579454
rect 74382 579218 74414 579454
rect 73794 579134 74414 579218
rect 73794 578898 73826 579134
rect 74062 578898 74146 579134
rect 74382 578898 74414 579134
rect 73794 543454 74414 578898
rect 73794 543218 73826 543454
rect 74062 543218 74146 543454
rect 74382 543218 74414 543454
rect 73794 543134 74414 543218
rect 73794 542898 73826 543134
rect 74062 542898 74146 543134
rect 74382 542898 74414 543134
rect 73794 507454 74414 542898
rect 73794 507218 73826 507454
rect 74062 507218 74146 507454
rect 74382 507218 74414 507454
rect 73794 507134 74414 507218
rect 73794 506898 73826 507134
rect 74062 506898 74146 507134
rect 74382 506898 74414 507134
rect 73794 471454 74414 506898
rect 73794 471218 73826 471454
rect 74062 471218 74146 471454
rect 74382 471218 74414 471454
rect 73794 471134 74414 471218
rect 73794 470898 73826 471134
rect 74062 470898 74146 471134
rect 74382 470898 74414 471134
rect 73794 435454 74414 470898
rect 73794 435218 73826 435454
rect 74062 435218 74146 435454
rect 74382 435218 74414 435454
rect 73794 435134 74414 435218
rect 73794 434898 73826 435134
rect 74062 434898 74146 435134
rect 74382 434898 74414 435134
rect 73794 399454 74414 434898
rect 73794 399218 73826 399454
rect 74062 399218 74146 399454
rect 74382 399218 74414 399454
rect 73794 399134 74414 399218
rect 73794 398898 73826 399134
rect 74062 398898 74146 399134
rect 74382 398898 74414 399134
rect 73794 363454 74414 398898
rect 73794 363218 73826 363454
rect 74062 363218 74146 363454
rect 74382 363218 74414 363454
rect 73794 363134 74414 363218
rect 73794 362898 73826 363134
rect 74062 362898 74146 363134
rect 74382 362898 74414 363134
rect 73794 327454 74414 362898
rect 73794 327218 73826 327454
rect 74062 327218 74146 327454
rect 74382 327218 74414 327454
rect 73794 327134 74414 327218
rect 73794 326898 73826 327134
rect 74062 326898 74146 327134
rect 74382 326898 74414 327134
rect 73794 291454 74414 326898
rect 73794 291218 73826 291454
rect 74062 291218 74146 291454
rect 74382 291218 74414 291454
rect 73794 291134 74414 291218
rect 73794 290898 73826 291134
rect 74062 290898 74146 291134
rect 74382 290898 74414 291134
rect 73794 255454 74414 290898
rect 73794 255218 73826 255454
rect 74062 255218 74146 255454
rect 74382 255218 74414 255454
rect 73794 255134 74414 255218
rect 73794 254898 73826 255134
rect 74062 254898 74146 255134
rect 74382 254898 74414 255134
rect 73794 219454 74414 254898
rect 73794 219218 73826 219454
rect 74062 219218 74146 219454
rect 74382 219218 74414 219454
rect 73794 219134 74414 219218
rect 73794 218898 73826 219134
rect 74062 218898 74146 219134
rect 74382 218898 74414 219134
rect 73794 183454 74414 218898
rect 73794 183218 73826 183454
rect 74062 183218 74146 183454
rect 74382 183218 74414 183454
rect 73794 183134 74414 183218
rect 73794 182898 73826 183134
rect 74062 182898 74146 183134
rect 74382 182898 74414 183134
rect 73794 147454 74414 182898
rect 73794 147218 73826 147454
rect 74062 147218 74146 147454
rect 74382 147218 74414 147454
rect 73794 147134 74414 147218
rect 73794 146898 73826 147134
rect 74062 146898 74146 147134
rect 74382 146898 74414 147134
rect 73794 111454 74414 146898
rect 73794 111218 73826 111454
rect 74062 111218 74146 111454
rect 74382 111218 74414 111454
rect 73794 111134 74414 111218
rect 73794 110898 73826 111134
rect 74062 110898 74146 111134
rect 74382 110898 74414 111134
rect 73794 75454 74414 110898
rect 73794 75218 73826 75454
rect 74062 75218 74146 75454
rect 74382 75218 74414 75454
rect 73794 75134 74414 75218
rect 73794 74898 73826 75134
rect 74062 74898 74146 75134
rect 74382 74898 74414 75134
rect 73794 39454 74414 74898
rect 73794 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 74414 39454
rect 73794 39134 74414 39218
rect 73794 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 74414 39134
rect 73794 3454 74414 38898
rect 73794 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 74414 3454
rect 73794 3134 74414 3218
rect 73794 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 74414 3134
rect 73794 -346 74414 2898
rect 73794 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 74414 -346
rect 73794 -666 74414 -582
rect 73794 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 74414 -666
rect 73794 -7654 74414 -902
rect 78294 705798 78914 711590
rect 78294 705562 78326 705798
rect 78562 705562 78646 705798
rect 78882 705562 78914 705798
rect 78294 705478 78914 705562
rect 78294 705242 78326 705478
rect 78562 705242 78646 705478
rect 78882 705242 78914 705478
rect 78294 691954 78914 705242
rect 78294 691718 78326 691954
rect 78562 691718 78646 691954
rect 78882 691718 78914 691954
rect 78294 691634 78914 691718
rect 78294 691398 78326 691634
rect 78562 691398 78646 691634
rect 78882 691398 78914 691634
rect 78294 655954 78914 691398
rect 78294 655718 78326 655954
rect 78562 655718 78646 655954
rect 78882 655718 78914 655954
rect 78294 655634 78914 655718
rect 78294 655398 78326 655634
rect 78562 655398 78646 655634
rect 78882 655398 78914 655634
rect 78294 619954 78914 655398
rect 78294 619718 78326 619954
rect 78562 619718 78646 619954
rect 78882 619718 78914 619954
rect 78294 619634 78914 619718
rect 78294 619398 78326 619634
rect 78562 619398 78646 619634
rect 78882 619398 78914 619634
rect 78294 583954 78914 619398
rect 78294 583718 78326 583954
rect 78562 583718 78646 583954
rect 78882 583718 78914 583954
rect 78294 583634 78914 583718
rect 78294 583398 78326 583634
rect 78562 583398 78646 583634
rect 78882 583398 78914 583634
rect 78294 547954 78914 583398
rect 78294 547718 78326 547954
rect 78562 547718 78646 547954
rect 78882 547718 78914 547954
rect 78294 547634 78914 547718
rect 78294 547398 78326 547634
rect 78562 547398 78646 547634
rect 78882 547398 78914 547634
rect 78294 511954 78914 547398
rect 78294 511718 78326 511954
rect 78562 511718 78646 511954
rect 78882 511718 78914 511954
rect 78294 511634 78914 511718
rect 78294 511398 78326 511634
rect 78562 511398 78646 511634
rect 78882 511398 78914 511634
rect 78294 475954 78914 511398
rect 78294 475718 78326 475954
rect 78562 475718 78646 475954
rect 78882 475718 78914 475954
rect 78294 475634 78914 475718
rect 78294 475398 78326 475634
rect 78562 475398 78646 475634
rect 78882 475398 78914 475634
rect 78294 439954 78914 475398
rect 78294 439718 78326 439954
rect 78562 439718 78646 439954
rect 78882 439718 78914 439954
rect 78294 439634 78914 439718
rect 78294 439398 78326 439634
rect 78562 439398 78646 439634
rect 78882 439398 78914 439634
rect 78294 403954 78914 439398
rect 78294 403718 78326 403954
rect 78562 403718 78646 403954
rect 78882 403718 78914 403954
rect 78294 403634 78914 403718
rect 78294 403398 78326 403634
rect 78562 403398 78646 403634
rect 78882 403398 78914 403634
rect 78294 367954 78914 403398
rect 78294 367718 78326 367954
rect 78562 367718 78646 367954
rect 78882 367718 78914 367954
rect 78294 367634 78914 367718
rect 78294 367398 78326 367634
rect 78562 367398 78646 367634
rect 78882 367398 78914 367634
rect 78294 331954 78914 367398
rect 78294 331718 78326 331954
rect 78562 331718 78646 331954
rect 78882 331718 78914 331954
rect 78294 331634 78914 331718
rect 78294 331398 78326 331634
rect 78562 331398 78646 331634
rect 78882 331398 78914 331634
rect 78294 295954 78914 331398
rect 78294 295718 78326 295954
rect 78562 295718 78646 295954
rect 78882 295718 78914 295954
rect 78294 295634 78914 295718
rect 78294 295398 78326 295634
rect 78562 295398 78646 295634
rect 78882 295398 78914 295634
rect 78294 259954 78914 295398
rect 78294 259718 78326 259954
rect 78562 259718 78646 259954
rect 78882 259718 78914 259954
rect 78294 259634 78914 259718
rect 78294 259398 78326 259634
rect 78562 259398 78646 259634
rect 78882 259398 78914 259634
rect 78294 223954 78914 259398
rect 78294 223718 78326 223954
rect 78562 223718 78646 223954
rect 78882 223718 78914 223954
rect 78294 223634 78914 223718
rect 78294 223398 78326 223634
rect 78562 223398 78646 223634
rect 78882 223398 78914 223634
rect 78294 187954 78914 223398
rect 78294 187718 78326 187954
rect 78562 187718 78646 187954
rect 78882 187718 78914 187954
rect 78294 187634 78914 187718
rect 78294 187398 78326 187634
rect 78562 187398 78646 187634
rect 78882 187398 78914 187634
rect 78294 151954 78914 187398
rect 78294 151718 78326 151954
rect 78562 151718 78646 151954
rect 78882 151718 78914 151954
rect 78294 151634 78914 151718
rect 78294 151398 78326 151634
rect 78562 151398 78646 151634
rect 78882 151398 78914 151634
rect 78294 115954 78914 151398
rect 78294 115718 78326 115954
rect 78562 115718 78646 115954
rect 78882 115718 78914 115954
rect 78294 115634 78914 115718
rect 78294 115398 78326 115634
rect 78562 115398 78646 115634
rect 78882 115398 78914 115634
rect 78294 79954 78914 115398
rect 78294 79718 78326 79954
rect 78562 79718 78646 79954
rect 78882 79718 78914 79954
rect 78294 79634 78914 79718
rect 78294 79398 78326 79634
rect 78562 79398 78646 79634
rect 78882 79398 78914 79634
rect 78294 43954 78914 79398
rect 78294 43718 78326 43954
rect 78562 43718 78646 43954
rect 78882 43718 78914 43954
rect 78294 43634 78914 43718
rect 78294 43398 78326 43634
rect 78562 43398 78646 43634
rect 78882 43398 78914 43634
rect 78294 7954 78914 43398
rect 78294 7718 78326 7954
rect 78562 7718 78646 7954
rect 78882 7718 78914 7954
rect 78294 7634 78914 7718
rect 78294 7398 78326 7634
rect 78562 7398 78646 7634
rect 78882 7398 78914 7634
rect 78294 -1306 78914 7398
rect 78294 -1542 78326 -1306
rect 78562 -1542 78646 -1306
rect 78882 -1542 78914 -1306
rect 78294 -1626 78914 -1542
rect 78294 -1862 78326 -1626
rect 78562 -1862 78646 -1626
rect 78882 -1862 78914 -1626
rect 78294 -7654 78914 -1862
rect 82794 706758 83414 711590
rect 82794 706522 82826 706758
rect 83062 706522 83146 706758
rect 83382 706522 83414 706758
rect 82794 706438 83414 706522
rect 82794 706202 82826 706438
rect 83062 706202 83146 706438
rect 83382 706202 83414 706438
rect 82794 696454 83414 706202
rect 82794 696218 82826 696454
rect 83062 696218 83146 696454
rect 83382 696218 83414 696454
rect 82794 696134 83414 696218
rect 82794 695898 82826 696134
rect 83062 695898 83146 696134
rect 83382 695898 83414 696134
rect 82794 660454 83414 695898
rect 82794 660218 82826 660454
rect 83062 660218 83146 660454
rect 83382 660218 83414 660454
rect 82794 660134 83414 660218
rect 82794 659898 82826 660134
rect 83062 659898 83146 660134
rect 83382 659898 83414 660134
rect 82794 624454 83414 659898
rect 82794 624218 82826 624454
rect 83062 624218 83146 624454
rect 83382 624218 83414 624454
rect 82794 624134 83414 624218
rect 82794 623898 82826 624134
rect 83062 623898 83146 624134
rect 83382 623898 83414 624134
rect 82794 588454 83414 623898
rect 82794 588218 82826 588454
rect 83062 588218 83146 588454
rect 83382 588218 83414 588454
rect 82794 588134 83414 588218
rect 82794 587898 82826 588134
rect 83062 587898 83146 588134
rect 83382 587898 83414 588134
rect 82794 552454 83414 587898
rect 82794 552218 82826 552454
rect 83062 552218 83146 552454
rect 83382 552218 83414 552454
rect 82794 552134 83414 552218
rect 82794 551898 82826 552134
rect 83062 551898 83146 552134
rect 83382 551898 83414 552134
rect 82794 516454 83414 551898
rect 82794 516218 82826 516454
rect 83062 516218 83146 516454
rect 83382 516218 83414 516454
rect 82794 516134 83414 516218
rect 82794 515898 82826 516134
rect 83062 515898 83146 516134
rect 83382 515898 83414 516134
rect 82794 480454 83414 515898
rect 82794 480218 82826 480454
rect 83062 480218 83146 480454
rect 83382 480218 83414 480454
rect 82794 480134 83414 480218
rect 82794 479898 82826 480134
rect 83062 479898 83146 480134
rect 83382 479898 83414 480134
rect 82794 444454 83414 479898
rect 82794 444218 82826 444454
rect 83062 444218 83146 444454
rect 83382 444218 83414 444454
rect 82794 444134 83414 444218
rect 82794 443898 82826 444134
rect 83062 443898 83146 444134
rect 83382 443898 83414 444134
rect 82794 408454 83414 443898
rect 82794 408218 82826 408454
rect 83062 408218 83146 408454
rect 83382 408218 83414 408454
rect 82794 408134 83414 408218
rect 82794 407898 82826 408134
rect 83062 407898 83146 408134
rect 83382 407898 83414 408134
rect 82794 372454 83414 407898
rect 82794 372218 82826 372454
rect 83062 372218 83146 372454
rect 83382 372218 83414 372454
rect 82794 372134 83414 372218
rect 82794 371898 82826 372134
rect 83062 371898 83146 372134
rect 83382 371898 83414 372134
rect 82794 336454 83414 371898
rect 82794 336218 82826 336454
rect 83062 336218 83146 336454
rect 83382 336218 83414 336454
rect 82794 336134 83414 336218
rect 82794 335898 82826 336134
rect 83062 335898 83146 336134
rect 83382 335898 83414 336134
rect 82794 300454 83414 335898
rect 82794 300218 82826 300454
rect 83062 300218 83146 300454
rect 83382 300218 83414 300454
rect 82794 300134 83414 300218
rect 82794 299898 82826 300134
rect 83062 299898 83146 300134
rect 83382 299898 83414 300134
rect 82794 264454 83414 299898
rect 82794 264218 82826 264454
rect 83062 264218 83146 264454
rect 83382 264218 83414 264454
rect 82794 264134 83414 264218
rect 82794 263898 82826 264134
rect 83062 263898 83146 264134
rect 83382 263898 83414 264134
rect 82794 228454 83414 263898
rect 82794 228218 82826 228454
rect 83062 228218 83146 228454
rect 83382 228218 83414 228454
rect 82794 228134 83414 228218
rect 82794 227898 82826 228134
rect 83062 227898 83146 228134
rect 83382 227898 83414 228134
rect 82794 192454 83414 227898
rect 82794 192218 82826 192454
rect 83062 192218 83146 192454
rect 83382 192218 83414 192454
rect 82794 192134 83414 192218
rect 82794 191898 82826 192134
rect 83062 191898 83146 192134
rect 83382 191898 83414 192134
rect 82794 156454 83414 191898
rect 82794 156218 82826 156454
rect 83062 156218 83146 156454
rect 83382 156218 83414 156454
rect 82794 156134 83414 156218
rect 82794 155898 82826 156134
rect 83062 155898 83146 156134
rect 83382 155898 83414 156134
rect 82794 120454 83414 155898
rect 82794 120218 82826 120454
rect 83062 120218 83146 120454
rect 83382 120218 83414 120454
rect 82794 120134 83414 120218
rect 82794 119898 82826 120134
rect 83062 119898 83146 120134
rect 83382 119898 83414 120134
rect 82794 84454 83414 119898
rect 82794 84218 82826 84454
rect 83062 84218 83146 84454
rect 83382 84218 83414 84454
rect 82794 84134 83414 84218
rect 82794 83898 82826 84134
rect 83062 83898 83146 84134
rect 83382 83898 83414 84134
rect 82794 48454 83414 83898
rect 82794 48218 82826 48454
rect 83062 48218 83146 48454
rect 83382 48218 83414 48454
rect 82794 48134 83414 48218
rect 82794 47898 82826 48134
rect 83062 47898 83146 48134
rect 83382 47898 83414 48134
rect 82794 12454 83414 47898
rect 82794 12218 82826 12454
rect 83062 12218 83146 12454
rect 83382 12218 83414 12454
rect 82794 12134 83414 12218
rect 82794 11898 82826 12134
rect 83062 11898 83146 12134
rect 83382 11898 83414 12134
rect 82794 -2266 83414 11898
rect 82794 -2502 82826 -2266
rect 83062 -2502 83146 -2266
rect 83382 -2502 83414 -2266
rect 82794 -2586 83414 -2502
rect 82794 -2822 82826 -2586
rect 83062 -2822 83146 -2586
rect 83382 -2822 83414 -2586
rect 82794 -7654 83414 -2822
rect 87294 707718 87914 711590
rect 87294 707482 87326 707718
rect 87562 707482 87646 707718
rect 87882 707482 87914 707718
rect 87294 707398 87914 707482
rect 87294 707162 87326 707398
rect 87562 707162 87646 707398
rect 87882 707162 87914 707398
rect 87294 700954 87914 707162
rect 87294 700718 87326 700954
rect 87562 700718 87646 700954
rect 87882 700718 87914 700954
rect 87294 700634 87914 700718
rect 87294 700398 87326 700634
rect 87562 700398 87646 700634
rect 87882 700398 87914 700634
rect 87294 664954 87914 700398
rect 87294 664718 87326 664954
rect 87562 664718 87646 664954
rect 87882 664718 87914 664954
rect 87294 664634 87914 664718
rect 87294 664398 87326 664634
rect 87562 664398 87646 664634
rect 87882 664398 87914 664634
rect 87294 628954 87914 664398
rect 87294 628718 87326 628954
rect 87562 628718 87646 628954
rect 87882 628718 87914 628954
rect 87294 628634 87914 628718
rect 87294 628398 87326 628634
rect 87562 628398 87646 628634
rect 87882 628398 87914 628634
rect 87294 592954 87914 628398
rect 87294 592718 87326 592954
rect 87562 592718 87646 592954
rect 87882 592718 87914 592954
rect 87294 592634 87914 592718
rect 87294 592398 87326 592634
rect 87562 592398 87646 592634
rect 87882 592398 87914 592634
rect 87294 556954 87914 592398
rect 87294 556718 87326 556954
rect 87562 556718 87646 556954
rect 87882 556718 87914 556954
rect 87294 556634 87914 556718
rect 87294 556398 87326 556634
rect 87562 556398 87646 556634
rect 87882 556398 87914 556634
rect 87294 520954 87914 556398
rect 87294 520718 87326 520954
rect 87562 520718 87646 520954
rect 87882 520718 87914 520954
rect 87294 520634 87914 520718
rect 87294 520398 87326 520634
rect 87562 520398 87646 520634
rect 87882 520398 87914 520634
rect 87294 484954 87914 520398
rect 87294 484718 87326 484954
rect 87562 484718 87646 484954
rect 87882 484718 87914 484954
rect 87294 484634 87914 484718
rect 87294 484398 87326 484634
rect 87562 484398 87646 484634
rect 87882 484398 87914 484634
rect 87294 448954 87914 484398
rect 87294 448718 87326 448954
rect 87562 448718 87646 448954
rect 87882 448718 87914 448954
rect 87294 448634 87914 448718
rect 87294 448398 87326 448634
rect 87562 448398 87646 448634
rect 87882 448398 87914 448634
rect 87294 412954 87914 448398
rect 87294 412718 87326 412954
rect 87562 412718 87646 412954
rect 87882 412718 87914 412954
rect 87294 412634 87914 412718
rect 87294 412398 87326 412634
rect 87562 412398 87646 412634
rect 87882 412398 87914 412634
rect 87294 376954 87914 412398
rect 87294 376718 87326 376954
rect 87562 376718 87646 376954
rect 87882 376718 87914 376954
rect 87294 376634 87914 376718
rect 87294 376398 87326 376634
rect 87562 376398 87646 376634
rect 87882 376398 87914 376634
rect 87294 340954 87914 376398
rect 87294 340718 87326 340954
rect 87562 340718 87646 340954
rect 87882 340718 87914 340954
rect 87294 340634 87914 340718
rect 87294 340398 87326 340634
rect 87562 340398 87646 340634
rect 87882 340398 87914 340634
rect 87294 304954 87914 340398
rect 87294 304718 87326 304954
rect 87562 304718 87646 304954
rect 87882 304718 87914 304954
rect 87294 304634 87914 304718
rect 87294 304398 87326 304634
rect 87562 304398 87646 304634
rect 87882 304398 87914 304634
rect 87294 268954 87914 304398
rect 87294 268718 87326 268954
rect 87562 268718 87646 268954
rect 87882 268718 87914 268954
rect 87294 268634 87914 268718
rect 87294 268398 87326 268634
rect 87562 268398 87646 268634
rect 87882 268398 87914 268634
rect 87294 232954 87914 268398
rect 87294 232718 87326 232954
rect 87562 232718 87646 232954
rect 87882 232718 87914 232954
rect 87294 232634 87914 232718
rect 87294 232398 87326 232634
rect 87562 232398 87646 232634
rect 87882 232398 87914 232634
rect 87294 196954 87914 232398
rect 87294 196718 87326 196954
rect 87562 196718 87646 196954
rect 87882 196718 87914 196954
rect 87294 196634 87914 196718
rect 87294 196398 87326 196634
rect 87562 196398 87646 196634
rect 87882 196398 87914 196634
rect 87294 160954 87914 196398
rect 87294 160718 87326 160954
rect 87562 160718 87646 160954
rect 87882 160718 87914 160954
rect 87294 160634 87914 160718
rect 87294 160398 87326 160634
rect 87562 160398 87646 160634
rect 87882 160398 87914 160634
rect 87294 124954 87914 160398
rect 87294 124718 87326 124954
rect 87562 124718 87646 124954
rect 87882 124718 87914 124954
rect 87294 124634 87914 124718
rect 87294 124398 87326 124634
rect 87562 124398 87646 124634
rect 87882 124398 87914 124634
rect 87294 88954 87914 124398
rect 87294 88718 87326 88954
rect 87562 88718 87646 88954
rect 87882 88718 87914 88954
rect 87294 88634 87914 88718
rect 87294 88398 87326 88634
rect 87562 88398 87646 88634
rect 87882 88398 87914 88634
rect 87294 52954 87914 88398
rect 87294 52718 87326 52954
rect 87562 52718 87646 52954
rect 87882 52718 87914 52954
rect 87294 52634 87914 52718
rect 87294 52398 87326 52634
rect 87562 52398 87646 52634
rect 87882 52398 87914 52634
rect 87294 16954 87914 52398
rect 87294 16718 87326 16954
rect 87562 16718 87646 16954
rect 87882 16718 87914 16954
rect 87294 16634 87914 16718
rect 87294 16398 87326 16634
rect 87562 16398 87646 16634
rect 87882 16398 87914 16634
rect 87294 -3226 87914 16398
rect 87294 -3462 87326 -3226
rect 87562 -3462 87646 -3226
rect 87882 -3462 87914 -3226
rect 87294 -3546 87914 -3462
rect 87294 -3782 87326 -3546
rect 87562 -3782 87646 -3546
rect 87882 -3782 87914 -3546
rect 87294 -7654 87914 -3782
rect 91794 708678 92414 711590
rect 91794 708442 91826 708678
rect 92062 708442 92146 708678
rect 92382 708442 92414 708678
rect 91794 708358 92414 708442
rect 91794 708122 91826 708358
rect 92062 708122 92146 708358
rect 92382 708122 92414 708358
rect 91794 669454 92414 708122
rect 91794 669218 91826 669454
rect 92062 669218 92146 669454
rect 92382 669218 92414 669454
rect 91794 669134 92414 669218
rect 91794 668898 91826 669134
rect 92062 668898 92146 669134
rect 92382 668898 92414 669134
rect 91794 633454 92414 668898
rect 96294 709638 96914 711590
rect 96294 709402 96326 709638
rect 96562 709402 96646 709638
rect 96882 709402 96914 709638
rect 96294 709318 96914 709402
rect 96294 709082 96326 709318
rect 96562 709082 96646 709318
rect 96882 709082 96914 709318
rect 96294 673954 96914 709082
rect 96294 673718 96326 673954
rect 96562 673718 96646 673954
rect 96882 673718 96914 673954
rect 96294 673634 96914 673718
rect 96294 673398 96326 673634
rect 96562 673398 96646 673634
rect 96882 673398 96914 673634
rect 95739 656980 95805 656981
rect 95739 656916 95740 656980
rect 95804 656916 95805 656980
rect 95739 656915 95805 656916
rect 91794 633218 91826 633454
rect 92062 633218 92146 633454
rect 92382 633218 92414 633454
rect 91794 633134 92414 633218
rect 91794 632898 91826 633134
rect 92062 632898 92146 633134
rect 92382 632898 92414 633134
rect 91794 597454 92414 632898
rect 91794 597218 91826 597454
rect 92062 597218 92146 597454
rect 92382 597218 92414 597454
rect 91794 597134 92414 597218
rect 91794 596898 91826 597134
rect 92062 596898 92146 597134
rect 92382 596898 92414 597134
rect 91794 561454 92414 596898
rect 91794 561218 91826 561454
rect 92062 561218 92146 561454
rect 92382 561218 92414 561454
rect 91794 561134 92414 561218
rect 91794 560898 91826 561134
rect 92062 560898 92146 561134
rect 92382 560898 92414 561134
rect 91794 525454 92414 560898
rect 91794 525218 91826 525454
rect 92062 525218 92146 525454
rect 92382 525218 92414 525454
rect 91794 525134 92414 525218
rect 91794 524898 91826 525134
rect 92062 524898 92146 525134
rect 92382 524898 92414 525134
rect 91794 489454 92414 524898
rect 91794 489218 91826 489454
rect 92062 489218 92146 489454
rect 92382 489218 92414 489454
rect 91794 489134 92414 489218
rect 91794 488898 91826 489134
rect 92062 488898 92146 489134
rect 92382 488898 92414 489134
rect 91794 453454 92414 488898
rect 91794 453218 91826 453454
rect 92062 453218 92146 453454
rect 92382 453218 92414 453454
rect 91794 453134 92414 453218
rect 91794 452898 91826 453134
rect 92062 452898 92146 453134
rect 92382 452898 92414 453134
rect 91794 417454 92414 452898
rect 91794 417218 91826 417454
rect 92062 417218 92146 417454
rect 92382 417218 92414 417454
rect 91794 417134 92414 417218
rect 91794 416898 91826 417134
rect 92062 416898 92146 417134
rect 92382 416898 92414 417134
rect 91794 381454 92414 416898
rect 91794 381218 91826 381454
rect 92062 381218 92146 381454
rect 92382 381218 92414 381454
rect 91794 381134 92414 381218
rect 91794 380898 91826 381134
rect 92062 380898 92146 381134
rect 92382 380898 92414 381134
rect 91794 345454 92414 380898
rect 91794 345218 91826 345454
rect 92062 345218 92146 345454
rect 92382 345218 92414 345454
rect 91794 345134 92414 345218
rect 91794 344898 91826 345134
rect 92062 344898 92146 345134
rect 92382 344898 92414 345134
rect 91794 309454 92414 344898
rect 91794 309218 91826 309454
rect 92062 309218 92146 309454
rect 92382 309218 92414 309454
rect 91794 309134 92414 309218
rect 91794 308898 91826 309134
rect 92062 308898 92146 309134
rect 92382 308898 92414 309134
rect 91794 273454 92414 308898
rect 91794 273218 91826 273454
rect 92062 273218 92146 273454
rect 92382 273218 92414 273454
rect 91794 273134 92414 273218
rect 91794 272898 91826 273134
rect 92062 272898 92146 273134
rect 92382 272898 92414 273134
rect 91794 237454 92414 272898
rect 91794 237218 91826 237454
rect 92062 237218 92146 237454
rect 92382 237218 92414 237454
rect 91794 237134 92414 237218
rect 91794 236898 91826 237134
rect 92062 236898 92146 237134
rect 92382 236898 92414 237134
rect 91794 201454 92414 236898
rect 91794 201218 91826 201454
rect 92062 201218 92146 201454
rect 92382 201218 92414 201454
rect 91794 201134 92414 201218
rect 91794 200898 91826 201134
rect 92062 200898 92146 201134
rect 92382 200898 92414 201134
rect 91794 165454 92414 200898
rect 95742 191589 95802 656915
rect 96294 637954 96914 673398
rect 96294 637718 96326 637954
rect 96562 637718 96646 637954
rect 96882 637718 96914 637954
rect 96294 637634 96914 637718
rect 96294 637398 96326 637634
rect 96562 637398 96646 637634
rect 96882 637398 96914 637634
rect 96294 601954 96914 637398
rect 96294 601718 96326 601954
rect 96562 601718 96646 601954
rect 96882 601718 96914 601954
rect 96294 601634 96914 601718
rect 96294 601398 96326 601634
rect 96562 601398 96646 601634
rect 96882 601398 96914 601634
rect 96294 565954 96914 601398
rect 96294 565718 96326 565954
rect 96562 565718 96646 565954
rect 96882 565718 96914 565954
rect 96294 565634 96914 565718
rect 96294 565398 96326 565634
rect 96562 565398 96646 565634
rect 96882 565398 96914 565634
rect 96294 529954 96914 565398
rect 96294 529718 96326 529954
rect 96562 529718 96646 529954
rect 96882 529718 96914 529954
rect 96294 529634 96914 529718
rect 96294 529398 96326 529634
rect 96562 529398 96646 529634
rect 96882 529398 96914 529634
rect 96294 493954 96914 529398
rect 96294 493718 96326 493954
rect 96562 493718 96646 493954
rect 96882 493718 96914 493954
rect 96294 493634 96914 493718
rect 96294 493398 96326 493634
rect 96562 493398 96646 493634
rect 96882 493398 96914 493634
rect 96294 457954 96914 493398
rect 96294 457718 96326 457954
rect 96562 457718 96646 457954
rect 96882 457718 96914 457954
rect 96294 457634 96914 457718
rect 96294 457398 96326 457634
rect 96562 457398 96646 457634
rect 96882 457398 96914 457634
rect 96294 421954 96914 457398
rect 96294 421718 96326 421954
rect 96562 421718 96646 421954
rect 96882 421718 96914 421954
rect 96294 421634 96914 421718
rect 96294 421398 96326 421634
rect 96562 421398 96646 421634
rect 96882 421398 96914 421634
rect 96294 385954 96914 421398
rect 96294 385718 96326 385954
rect 96562 385718 96646 385954
rect 96882 385718 96914 385954
rect 96294 385634 96914 385718
rect 96294 385398 96326 385634
rect 96562 385398 96646 385634
rect 96882 385398 96914 385634
rect 96294 349954 96914 385398
rect 96294 349718 96326 349954
rect 96562 349718 96646 349954
rect 96882 349718 96914 349954
rect 96294 349634 96914 349718
rect 96294 349398 96326 349634
rect 96562 349398 96646 349634
rect 96882 349398 96914 349634
rect 96294 313954 96914 349398
rect 96294 313718 96326 313954
rect 96562 313718 96646 313954
rect 96882 313718 96914 313954
rect 96294 313634 96914 313718
rect 96294 313398 96326 313634
rect 96562 313398 96646 313634
rect 96882 313398 96914 313634
rect 96294 277954 96914 313398
rect 96294 277718 96326 277954
rect 96562 277718 96646 277954
rect 96882 277718 96914 277954
rect 96294 277634 96914 277718
rect 96294 277398 96326 277634
rect 96562 277398 96646 277634
rect 96882 277398 96914 277634
rect 96294 241954 96914 277398
rect 96294 241718 96326 241954
rect 96562 241718 96646 241954
rect 96882 241718 96914 241954
rect 96294 241634 96914 241718
rect 96294 241398 96326 241634
rect 96562 241398 96646 241634
rect 96882 241398 96914 241634
rect 96294 205954 96914 241398
rect 96294 205718 96326 205954
rect 96562 205718 96646 205954
rect 96882 205718 96914 205954
rect 96294 205634 96914 205718
rect 96294 205398 96326 205634
rect 96562 205398 96646 205634
rect 96882 205398 96914 205634
rect 95739 191588 95805 191589
rect 95739 191524 95740 191588
rect 95804 191524 95805 191588
rect 95739 191523 95805 191524
rect 91794 165218 91826 165454
rect 92062 165218 92146 165454
rect 92382 165218 92414 165454
rect 91794 165134 92414 165218
rect 91794 164898 91826 165134
rect 92062 164898 92146 165134
rect 92382 164898 92414 165134
rect 91794 129454 92414 164898
rect 91794 129218 91826 129454
rect 92062 129218 92146 129454
rect 92382 129218 92414 129454
rect 91794 129134 92414 129218
rect 91794 128898 91826 129134
rect 92062 128898 92146 129134
rect 92382 128898 92414 129134
rect 91794 93454 92414 128898
rect 91794 93218 91826 93454
rect 92062 93218 92146 93454
rect 92382 93218 92414 93454
rect 91794 93134 92414 93218
rect 91794 92898 91826 93134
rect 92062 92898 92146 93134
rect 92382 92898 92414 93134
rect 91794 57454 92414 92898
rect 91794 57218 91826 57454
rect 92062 57218 92146 57454
rect 92382 57218 92414 57454
rect 91794 57134 92414 57218
rect 91794 56898 91826 57134
rect 92062 56898 92146 57134
rect 92382 56898 92414 57134
rect 91794 21454 92414 56898
rect 91794 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 92414 21454
rect 91794 21134 92414 21218
rect 91794 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 92414 21134
rect 91794 -4186 92414 20898
rect 91794 -4422 91826 -4186
rect 92062 -4422 92146 -4186
rect 92382 -4422 92414 -4186
rect 91794 -4506 92414 -4422
rect 91794 -4742 91826 -4506
rect 92062 -4742 92146 -4506
rect 92382 -4742 92414 -4506
rect 91794 -7654 92414 -4742
rect 96294 169954 96914 205398
rect 100794 710598 101414 711590
rect 100794 710362 100826 710598
rect 101062 710362 101146 710598
rect 101382 710362 101414 710598
rect 100794 710278 101414 710362
rect 100794 710042 100826 710278
rect 101062 710042 101146 710278
rect 101382 710042 101414 710278
rect 100794 678454 101414 710042
rect 100794 678218 100826 678454
rect 101062 678218 101146 678454
rect 101382 678218 101414 678454
rect 100794 678134 101414 678218
rect 100794 677898 100826 678134
rect 101062 677898 101146 678134
rect 101382 677898 101414 678134
rect 100794 642454 101414 677898
rect 100794 642218 100826 642454
rect 101062 642218 101146 642454
rect 101382 642218 101414 642454
rect 100794 642134 101414 642218
rect 100794 641898 100826 642134
rect 101062 641898 101146 642134
rect 101382 641898 101414 642134
rect 100794 606454 101414 641898
rect 100794 606218 100826 606454
rect 101062 606218 101146 606454
rect 101382 606218 101414 606454
rect 100794 606134 101414 606218
rect 100794 605898 100826 606134
rect 101062 605898 101146 606134
rect 101382 605898 101414 606134
rect 100794 570454 101414 605898
rect 100794 570218 100826 570454
rect 101062 570218 101146 570454
rect 101382 570218 101414 570454
rect 100794 570134 101414 570218
rect 100794 569898 100826 570134
rect 101062 569898 101146 570134
rect 101382 569898 101414 570134
rect 100794 534454 101414 569898
rect 100794 534218 100826 534454
rect 101062 534218 101146 534454
rect 101382 534218 101414 534454
rect 100794 534134 101414 534218
rect 100794 533898 100826 534134
rect 101062 533898 101146 534134
rect 101382 533898 101414 534134
rect 100794 498454 101414 533898
rect 100794 498218 100826 498454
rect 101062 498218 101146 498454
rect 101382 498218 101414 498454
rect 100794 498134 101414 498218
rect 100794 497898 100826 498134
rect 101062 497898 101146 498134
rect 101382 497898 101414 498134
rect 100794 462454 101414 497898
rect 100794 462218 100826 462454
rect 101062 462218 101146 462454
rect 101382 462218 101414 462454
rect 100794 462134 101414 462218
rect 100794 461898 100826 462134
rect 101062 461898 101146 462134
rect 101382 461898 101414 462134
rect 100794 426454 101414 461898
rect 100794 426218 100826 426454
rect 101062 426218 101146 426454
rect 101382 426218 101414 426454
rect 100794 426134 101414 426218
rect 100794 425898 100826 426134
rect 101062 425898 101146 426134
rect 101382 425898 101414 426134
rect 100794 390454 101414 425898
rect 100794 390218 100826 390454
rect 101062 390218 101146 390454
rect 101382 390218 101414 390454
rect 100794 390134 101414 390218
rect 100794 389898 100826 390134
rect 101062 389898 101146 390134
rect 101382 389898 101414 390134
rect 100794 354454 101414 389898
rect 100794 354218 100826 354454
rect 101062 354218 101146 354454
rect 101382 354218 101414 354454
rect 100794 354134 101414 354218
rect 100794 353898 100826 354134
rect 101062 353898 101146 354134
rect 101382 353898 101414 354134
rect 100794 318454 101414 353898
rect 100794 318218 100826 318454
rect 101062 318218 101146 318454
rect 101382 318218 101414 318454
rect 100794 318134 101414 318218
rect 100794 317898 100826 318134
rect 101062 317898 101146 318134
rect 101382 317898 101414 318134
rect 100794 282454 101414 317898
rect 100794 282218 100826 282454
rect 101062 282218 101146 282454
rect 101382 282218 101414 282454
rect 100794 282134 101414 282218
rect 100794 281898 100826 282134
rect 101062 281898 101146 282134
rect 101382 281898 101414 282134
rect 100794 246454 101414 281898
rect 100794 246218 100826 246454
rect 101062 246218 101146 246454
rect 101382 246218 101414 246454
rect 100794 246134 101414 246218
rect 100794 245898 100826 246134
rect 101062 245898 101146 246134
rect 101382 245898 101414 246134
rect 100794 210454 101414 245898
rect 100794 210218 100826 210454
rect 101062 210218 101146 210454
rect 101382 210218 101414 210454
rect 100794 210134 101414 210218
rect 100794 209898 100826 210134
rect 101062 209898 101146 210134
rect 101382 209898 101414 210134
rect 97763 193900 97829 193901
rect 97763 193836 97764 193900
rect 97828 193836 97829 193900
rect 97763 193835 97829 193836
rect 97579 178124 97645 178125
rect 97579 178060 97580 178124
rect 97644 178060 97645 178124
rect 97579 178059 97645 178060
rect 96294 169718 96326 169954
rect 96562 169718 96646 169954
rect 96882 169718 96914 169954
rect 96294 169634 96914 169718
rect 96294 169398 96326 169634
rect 96562 169398 96646 169634
rect 96882 169398 96914 169634
rect 96294 133954 96914 169398
rect 96294 133718 96326 133954
rect 96562 133718 96646 133954
rect 96882 133718 96914 133954
rect 96294 133634 96914 133718
rect 96294 133398 96326 133634
rect 96562 133398 96646 133634
rect 96882 133398 96914 133634
rect 96294 97954 96914 133398
rect 96294 97718 96326 97954
rect 96562 97718 96646 97954
rect 96882 97718 96914 97954
rect 96294 97634 96914 97718
rect 96294 97398 96326 97634
rect 96562 97398 96646 97634
rect 96882 97398 96914 97634
rect 96294 61954 96914 97398
rect 97582 68373 97642 178059
rect 97766 77621 97826 193835
rect 100523 180844 100589 180845
rect 100523 180780 100524 180844
rect 100588 180780 100589 180844
rect 100523 180779 100589 180780
rect 100339 148612 100405 148613
rect 100339 148548 100340 148612
rect 100404 148548 100405 148612
rect 100339 148547 100405 148548
rect 100342 80749 100402 148547
rect 100339 80748 100405 80749
rect 100339 80684 100340 80748
rect 100404 80684 100405 80748
rect 100339 80683 100405 80684
rect 97763 77620 97829 77621
rect 97763 77556 97764 77620
rect 97828 77556 97829 77620
rect 97763 77555 97829 77556
rect 100526 68781 100586 180779
rect 100794 174454 101414 209898
rect 105294 711558 105914 711590
rect 105294 711322 105326 711558
rect 105562 711322 105646 711558
rect 105882 711322 105914 711558
rect 105294 711238 105914 711322
rect 105294 711002 105326 711238
rect 105562 711002 105646 711238
rect 105882 711002 105914 711238
rect 105294 682954 105914 711002
rect 105294 682718 105326 682954
rect 105562 682718 105646 682954
rect 105882 682718 105914 682954
rect 105294 682634 105914 682718
rect 105294 682398 105326 682634
rect 105562 682398 105646 682634
rect 105882 682398 105914 682634
rect 105294 646954 105914 682398
rect 105294 646718 105326 646954
rect 105562 646718 105646 646954
rect 105882 646718 105914 646954
rect 105294 646634 105914 646718
rect 105294 646398 105326 646634
rect 105562 646398 105646 646634
rect 105882 646398 105914 646634
rect 105294 610954 105914 646398
rect 105294 610718 105326 610954
rect 105562 610718 105646 610954
rect 105882 610718 105914 610954
rect 105294 610634 105914 610718
rect 105294 610398 105326 610634
rect 105562 610398 105646 610634
rect 105882 610398 105914 610634
rect 105294 574954 105914 610398
rect 105294 574718 105326 574954
rect 105562 574718 105646 574954
rect 105882 574718 105914 574954
rect 105294 574634 105914 574718
rect 105294 574398 105326 574634
rect 105562 574398 105646 574634
rect 105882 574398 105914 574634
rect 105294 538954 105914 574398
rect 105294 538718 105326 538954
rect 105562 538718 105646 538954
rect 105882 538718 105914 538954
rect 105294 538634 105914 538718
rect 105294 538398 105326 538634
rect 105562 538398 105646 538634
rect 105882 538398 105914 538634
rect 105294 502954 105914 538398
rect 105294 502718 105326 502954
rect 105562 502718 105646 502954
rect 105882 502718 105914 502954
rect 105294 502634 105914 502718
rect 105294 502398 105326 502634
rect 105562 502398 105646 502634
rect 105882 502398 105914 502634
rect 105294 466954 105914 502398
rect 105294 466718 105326 466954
rect 105562 466718 105646 466954
rect 105882 466718 105914 466954
rect 105294 466634 105914 466718
rect 105294 466398 105326 466634
rect 105562 466398 105646 466634
rect 105882 466398 105914 466634
rect 105294 430954 105914 466398
rect 105294 430718 105326 430954
rect 105562 430718 105646 430954
rect 105882 430718 105914 430954
rect 105294 430634 105914 430718
rect 105294 430398 105326 430634
rect 105562 430398 105646 430634
rect 105882 430398 105914 430634
rect 105294 394954 105914 430398
rect 105294 394718 105326 394954
rect 105562 394718 105646 394954
rect 105882 394718 105914 394954
rect 105294 394634 105914 394718
rect 105294 394398 105326 394634
rect 105562 394398 105646 394634
rect 105882 394398 105914 394634
rect 105294 358954 105914 394398
rect 105294 358718 105326 358954
rect 105562 358718 105646 358954
rect 105882 358718 105914 358954
rect 105294 358634 105914 358718
rect 105294 358398 105326 358634
rect 105562 358398 105646 358634
rect 105882 358398 105914 358634
rect 105294 322954 105914 358398
rect 105294 322718 105326 322954
rect 105562 322718 105646 322954
rect 105882 322718 105914 322954
rect 105294 322634 105914 322718
rect 105294 322398 105326 322634
rect 105562 322398 105646 322634
rect 105882 322398 105914 322634
rect 105294 286954 105914 322398
rect 105294 286718 105326 286954
rect 105562 286718 105646 286954
rect 105882 286718 105914 286954
rect 105294 286634 105914 286718
rect 105294 286398 105326 286634
rect 105562 286398 105646 286634
rect 105882 286398 105914 286634
rect 105294 250954 105914 286398
rect 105294 250718 105326 250954
rect 105562 250718 105646 250954
rect 105882 250718 105914 250954
rect 105294 250634 105914 250718
rect 105294 250398 105326 250634
rect 105562 250398 105646 250634
rect 105882 250398 105914 250634
rect 105294 214954 105914 250398
rect 105294 214718 105326 214954
rect 105562 214718 105646 214954
rect 105882 214718 105914 214954
rect 105294 214634 105914 214718
rect 105294 214398 105326 214634
rect 105562 214398 105646 214634
rect 105882 214398 105914 214634
rect 104755 197980 104821 197981
rect 104755 197916 104756 197980
rect 104820 197916 104821 197980
rect 104755 197915 104821 197916
rect 104571 191180 104637 191181
rect 104571 191116 104572 191180
rect 104636 191116 104637 191180
rect 104571 191115 104637 191116
rect 103283 181116 103349 181117
rect 103283 181052 103284 181116
rect 103348 181052 103349 181116
rect 103283 181051 103349 181052
rect 101995 180980 102061 180981
rect 101995 180916 101996 180980
rect 102060 180916 102061 180980
rect 101995 180915 102061 180916
rect 100794 174218 100826 174454
rect 101062 174218 101146 174454
rect 101382 174218 101414 174454
rect 100794 174134 101414 174218
rect 100794 173898 100826 174134
rect 101062 173898 101146 174134
rect 101382 173898 101414 174134
rect 100794 138454 101414 173898
rect 100794 138218 100826 138454
rect 101062 138218 101146 138454
rect 101382 138218 101414 138454
rect 100794 138134 101414 138218
rect 100794 137898 100826 138134
rect 101062 137898 101146 138134
rect 101382 137898 101414 138134
rect 100794 102454 101414 137898
rect 100794 102218 100826 102454
rect 101062 102218 101146 102454
rect 101382 102218 101414 102454
rect 100794 102134 101414 102218
rect 100794 101898 100826 102134
rect 101062 101898 101146 102134
rect 101382 101898 101414 102134
rect 100523 68780 100589 68781
rect 100523 68716 100524 68780
rect 100588 68716 100589 68780
rect 100523 68715 100589 68716
rect 97579 68372 97645 68373
rect 97579 68308 97580 68372
rect 97644 68308 97645 68372
rect 97579 68307 97645 68308
rect 96294 61718 96326 61954
rect 96562 61718 96646 61954
rect 96882 61718 96914 61954
rect 96294 61634 96914 61718
rect 96294 61398 96326 61634
rect 96562 61398 96646 61634
rect 96882 61398 96914 61634
rect 96294 25954 96914 61398
rect 96294 25718 96326 25954
rect 96562 25718 96646 25954
rect 96882 25718 96914 25954
rect 96294 25634 96914 25718
rect 96294 25398 96326 25634
rect 96562 25398 96646 25634
rect 96882 25398 96914 25634
rect 96294 -5146 96914 25398
rect 96294 -5382 96326 -5146
rect 96562 -5382 96646 -5146
rect 96882 -5382 96914 -5146
rect 96294 -5466 96914 -5382
rect 96294 -5702 96326 -5466
rect 96562 -5702 96646 -5466
rect 96882 -5702 96914 -5466
rect 96294 -7654 96914 -5702
rect 100794 66454 101414 101898
rect 101998 78437 102058 180915
rect 102915 174724 102981 174725
rect 102915 174660 102916 174724
rect 102980 174660 102981 174724
rect 102915 174659 102981 174660
rect 101995 78436 102061 78437
rect 101995 78372 101996 78436
rect 102060 78372 102061 78436
rect 101995 78371 102061 78372
rect 102918 75309 102978 174659
rect 103099 174588 103165 174589
rect 103099 174524 103100 174588
rect 103164 174524 103165 174588
rect 103099 174523 103165 174524
rect 102915 75308 102981 75309
rect 102915 75244 102916 75308
rect 102980 75244 102981 75308
rect 102915 75243 102981 75244
rect 103102 74085 103162 174523
rect 103286 78301 103346 181051
rect 104387 177308 104453 177309
rect 104387 177244 104388 177308
rect 104452 177244 104453 177308
rect 104387 177243 104453 177244
rect 103283 78300 103349 78301
rect 103283 78236 103284 78300
rect 103348 78236 103349 78300
rect 103283 78235 103349 78236
rect 104390 77213 104450 177243
rect 104387 77212 104453 77213
rect 104387 77148 104388 77212
rect 104452 77148 104453 77212
rect 104387 77147 104453 77148
rect 104574 77077 104634 191115
rect 104758 77893 104818 197915
rect 105294 178954 105914 214398
rect 109794 704838 110414 711590
rect 109794 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 110414 704838
rect 109794 704518 110414 704602
rect 109794 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 110414 704518
rect 109794 687454 110414 704282
rect 109794 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 110414 687454
rect 109794 687134 110414 687218
rect 109794 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 110414 687134
rect 109794 651454 110414 686898
rect 109794 651218 109826 651454
rect 110062 651218 110146 651454
rect 110382 651218 110414 651454
rect 109794 651134 110414 651218
rect 109794 650898 109826 651134
rect 110062 650898 110146 651134
rect 110382 650898 110414 651134
rect 109794 615454 110414 650898
rect 109794 615218 109826 615454
rect 110062 615218 110146 615454
rect 110382 615218 110414 615454
rect 109794 615134 110414 615218
rect 109794 614898 109826 615134
rect 110062 614898 110146 615134
rect 110382 614898 110414 615134
rect 109794 579454 110414 614898
rect 109794 579218 109826 579454
rect 110062 579218 110146 579454
rect 110382 579218 110414 579454
rect 109794 579134 110414 579218
rect 109794 578898 109826 579134
rect 110062 578898 110146 579134
rect 110382 578898 110414 579134
rect 109794 543454 110414 578898
rect 109794 543218 109826 543454
rect 110062 543218 110146 543454
rect 110382 543218 110414 543454
rect 109794 543134 110414 543218
rect 109794 542898 109826 543134
rect 110062 542898 110146 543134
rect 110382 542898 110414 543134
rect 109794 507454 110414 542898
rect 109794 507218 109826 507454
rect 110062 507218 110146 507454
rect 110382 507218 110414 507454
rect 109794 507134 110414 507218
rect 109794 506898 109826 507134
rect 110062 506898 110146 507134
rect 110382 506898 110414 507134
rect 109794 471454 110414 506898
rect 109794 471218 109826 471454
rect 110062 471218 110146 471454
rect 110382 471218 110414 471454
rect 109794 471134 110414 471218
rect 109794 470898 109826 471134
rect 110062 470898 110146 471134
rect 110382 470898 110414 471134
rect 109794 435454 110414 470898
rect 109794 435218 109826 435454
rect 110062 435218 110146 435454
rect 110382 435218 110414 435454
rect 109794 435134 110414 435218
rect 109794 434898 109826 435134
rect 110062 434898 110146 435134
rect 110382 434898 110414 435134
rect 109794 399454 110414 434898
rect 109794 399218 109826 399454
rect 110062 399218 110146 399454
rect 110382 399218 110414 399454
rect 109794 399134 110414 399218
rect 109794 398898 109826 399134
rect 110062 398898 110146 399134
rect 110382 398898 110414 399134
rect 109794 363454 110414 398898
rect 109794 363218 109826 363454
rect 110062 363218 110146 363454
rect 110382 363218 110414 363454
rect 109794 363134 110414 363218
rect 109794 362898 109826 363134
rect 110062 362898 110146 363134
rect 110382 362898 110414 363134
rect 109794 327454 110414 362898
rect 109794 327218 109826 327454
rect 110062 327218 110146 327454
rect 110382 327218 110414 327454
rect 109794 327134 110414 327218
rect 109794 326898 109826 327134
rect 110062 326898 110146 327134
rect 110382 326898 110414 327134
rect 109794 291454 110414 326898
rect 109794 291218 109826 291454
rect 110062 291218 110146 291454
rect 110382 291218 110414 291454
rect 109794 291134 110414 291218
rect 109794 290898 109826 291134
rect 110062 290898 110146 291134
rect 110382 290898 110414 291134
rect 109794 255454 110414 290898
rect 109794 255218 109826 255454
rect 110062 255218 110146 255454
rect 110382 255218 110414 255454
rect 109794 255134 110414 255218
rect 109794 254898 109826 255134
rect 110062 254898 110146 255134
rect 110382 254898 110414 255134
rect 109794 219454 110414 254898
rect 109794 219218 109826 219454
rect 110062 219218 110146 219454
rect 110382 219218 110414 219454
rect 109794 219134 110414 219218
rect 109794 218898 109826 219134
rect 110062 218898 110146 219134
rect 110382 218898 110414 219134
rect 109539 198932 109605 198933
rect 109539 198868 109540 198932
rect 109604 198868 109605 198932
rect 109539 198867 109605 198868
rect 108803 196620 108869 196621
rect 108803 196556 108804 196620
rect 108868 196556 108869 196620
rect 108803 196555 108869 196556
rect 107331 189820 107397 189821
rect 107331 189756 107332 189820
rect 107396 189756 107397 189820
rect 107331 189755 107397 189756
rect 107147 181388 107213 181389
rect 107147 181324 107148 181388
rect 107212 181324 107213 181388
rect 107147 181323 107213 181324
rect 106043 181252 106109 181253
rect 106043 181188 106044 181252
rect 106108 181188 106109 181252
rect 106043 181187 106109 181188
rect 105294 178718 105326 178954
rect 105562 178718 105646 178954
rect 105882 178718 105914 178954
rect 105294 178634 105914 178718
rect 105294 178398 105326 178634
rect 105562 178398 105646 178634
rect 105882 178398 105914 178634
rect 105294 142954 105914 178398
rect 105294 142718 105326 142954
rect 105562 142718 105646 142954
rect 105882 142718 105914 142954
rect 105294 142634 105914 142718
rect 105294 142398 105326 142634
rect 105562 142398 105646 142634
rect 105882 142398 105914 142634
rect 105294 106954 105914 142398
rect 105294 106718 105326 106954
rect 105562 106718 105646 106954
rect 105882 106718 105914 106954
rect 105294 106634 105914 106718
rect 105294 106398 105326 106634
rect 105562 106398 105646 106634
rect 105882 106398 105914 106634
rect 104755 77892 104821 77893
rect 104755 77828 104756 77892
rect 104820 77828 104821 77892
rect 104755 77827 104821 77828
rect 104571 77076 104637 77077
rect 104571 77012 104572 77076
rect 104636 77012 104637 77076
rect 104571 77011 104637 77012
rect 103099 74084 103165 74085
rect 103099 74020 103100 74084
rect 103164 74020 103165 74084
rect 103099 74019 103165 74020
rect 100794 66218 100826 66454
rect 101062 66218 101146 66454
rect 101382 66218 101414 66454
rect 100794 66134 101414 66218
rect 100794 65898 100826 66134
rect 101062 65898 101146 66134
rect 101382 65898 101414 66134
rect 100794 30454 101414 65898
rect 100794 30218 100826 30454
rect 101062 30218 101146 30454
rect 101382 30218 101414 30454
rect 100794 30134 101414 30218
rect 100794 29898 100826 30134
rect 101062 29898 101146 30134
rect 101382 29898 101414 30134
rect 100794 -6106 101414 29898
rect 100794 -6342 100826 -6106
rect 101062 -6342 101146 -6106
rect 101382 -6342 101414 -6106
rect 100794 -6426 101414 -6342
rect 100794 -6662 100826 -6426
rect 101062 -6662 101146 -6426
rect 101382 -6662 101414 -6426
rect 100794 -7654 101414 -6662
rect 105294 70954 105914 106398
rect 105294 70718 105326 70954
rect 105562 70718 105646 70954
rect 105882 70718 105914 70954
rect 105294 70634 105914 70718
rect 105294 70398 105326 70634
rect 105562 70398 105646 70634
rect 105882 70398 105914 70634
rect 105294 34954 105914 70398
rect 106046 68509 106106 181187
rect 107150 81293 107210 181323
rect 107147 81292 107213 81293
rect 107147 81228 107148 81292
rect 107212 81228 107213 81292
rect 107147 81227 107213 81228
rect 107334 79253 107394 189755
rect 108619 189684 108685 189685
rect 108619 189620 108620 189684
rect 108684 189620 108685 189684
rect 108619 189619 108685 189620
rect 108435 186964 108501 186965
rect 108435 186900 108436 186964
rect 108500 186900 108501 186964
rect 108435 186899 108501 186900
rect 107515 185060 107581 185061
rect 107515 184996 107516 185060
rect 107580 184996 107581 185060
rect 107515 184995 107581 184996
rect 107331 79252 107397 79253
rect 107331 79188 107332 79252
rect 107396 79188 107397 79252
rect 107331 79187 107397 79188
rect 107518 71637 107578 184995
rect 108251 184244 108317 184245
rect 108251 184180 108252 184244
rect 108316 184180 108317 184244
rect 108251 184179 108317 184180
rect 108254 78845 108314 184179
rect 108251 78844 108317 78845
rect 108251 78780 108252 78844
rect 108316 78780 108317 78844
rect 108251 78779 108317 78780
rect 107515 71636 107581 71637
rect 107515 71572 107516 71636
rect 107580 71572 107581 71636
rect 107515 71571 107581 71572
rect 108438 71501 108498 186899
rect 108435 71500 108501 71501
rect 108435 71436 108436 71500
rect 108500 71436 108501 71500
rect 108435 71435 108501 71436
rect 108622 71365 108682 189619
rect 108806 76941 108866 196555
rect 108803 76940 108869 76941
rect 108803 76876 108804 76940
rect 108868 76876 108869 76940
rect 108803 76875 108869 76876
rect 108619 71364 108685 71365
rect 108619 71300 108620 71364
rect 108684 71300 108685 71364
rect 108619 71299 108685 71300
rect 109542 70005 109602 198867
rect 109794 183454 110414 218898
rect 114294 705798 114914 711590
rect 114294 705562 114326 705798
rect 114562 705562 114646 705798
rect 114882 705562 114914 705798
rect 114294 705478 114914 705562
rect 114294 705242 114326 705478
rect 114562 705242 114646 705478
rect 114882 705242 114914 705478
rect 114294 691954 114914 705242
rect 114294 691718 114326 691954
rect 114562 691718 114646 691954
rect 114882 691718 114914 691954
rect 114294 691634 114914 691718
rect 114294 691398 114326 691634
rect 114562 691398 114646 691634
rect 114882 691398 114914 691634
rect 114294 655954 114914 691398
rect 114294 655718 114326 655954
rect 114562 655718 114646 655954
rect 114882 655718 114914 655954
rect 114294 655634 114914 655718
rect 114294 655398 114326 655634
rect 114562 655398 114646 655634
rect 114882 655398 114914 655634
rect 114294 619954 114914 655398
rect 114294 619718 114326 619954
rect 114562 619718 114646 619954
rect 114882 619718 114914 619954
rect 114294 619634 114914 619718
rect 114294 619398 114326 619634
rect 114562 619398 114646 619634
rect 114882 619398 114914 619634
rect 114294 583954 114914 619398
rect 114294 583718 114326 583954
rect 114562 583718 114646 583954
rect 114882 583718 114914 583954
rect 114294 583634 114914 583718
rect 114294 583398 114326 583634
rect 114562 583398 114646 583634
rect 114882 583398 114914 583634
rect 114294 547954 114914 583398
rect 114294 547718 114326 547954
rect 114562 547718 114646 547954
rect 114882 547718 114914 547954
rect 114294 547634 114914 547718
rect 114294 547398 114326 547634
rect 114562 547398 114646 547634
rect 114882 547398 114914 547634
rect 114294 511954 114914 547398
rect 114294 511718 114326 511954
rect 114562 511718 114646 511954
rect 114882 511718 114914 511954
rect 114294 511634 114914 511718
rect 114294 511398 114326 511634
rect 114562 511398 114646 511634
rect 114882 511398 114914 511634
rect 114294 475954 114914 511398
rect 114294 475718 114326 475954
rect 114562 475718 114646 475954
rect 114882 475718 114914 475954
rect 114294 475634 114914 475718
rect 114294 475398 114326 475634
rect 114562 475398 114646 475634
rect 114882 475398 114914 475634
rect 114294 439954 114914 475398
rect 114294 439718 114326 439954
rect 114562 439718 114646 439954
rect 114882 439718 114914 439954
rect 114294 439634 114914 439718
rect 114294 439398 114326 439634
rect 114562 439398 114646 439634
rect 114882 439398 114914 439634
rect 114294 403954 114914 439398
rect 114294 403718 114326 403954
rect 114562 403718 114646 403954
rect 114882 403718 114914 403954
rect 114294 403634 114914 403718
rect 114294 403398 114326 403634
rect 114562 403398 114646 403634
rect 114882 403398 114914 403634
rect 114294 367954 114914 403398
rect 114294 367718 114326 367954
rect 114562 367718 114646 367954
rect 114882 367718 114914 367954
rect 114294 367634 114914 367718
rect 114294 367398 114326 367634
rect 114562 367398 114646 367634
rect 114882 367398 114914 367634
rect 114294 331954 114914 367398
rect 114294 331718 114326 331954
rect 114562 331718 114646 331954
rect 114882 331718 114914 331954
rect 114294 331634 114914 331718
rect 114294 331398 114326 331634
rect 114562 331398 114646 331634
rect 114882 331398 114914 331634
rect 114294 295954 114914 331398
rect 114294 295718 114326 295954
rect 114562 295718 114646 295954
rect 114882 295718 114914 295954
rect 114294 295634 114914 295718
rect 114294 295398 114326 295634
rect 114562 295398 114646 295634
rect 114882 295398 114914 295634
rect 114294 259954 114914 295398
rect 118794 706758 119414 711590
rect 118794 706522 118826 706758
rect 119062 706522 119146 706758
rect 119382 706522 119414 706758
rect 118794 706438 119414 706522
rect 118794 706202 118826 706438
rect 119062 706202 119146 706438
rect 119382 706202 119414 706438
rect 118794 696454 119414 706202
rect 118794 696218 118826 696454
rect 119062 696218 119146 696454
rect 119382 696218 119414 696454
rect 118794 696134 119414 696218
rect 118794 695898 118826 696134
rect 119062 695898 119146 696134
rect 119382 695898 119414 696134
rect 118794 660454 119414 695898
rect 118794 660218 118826 660454
rect 119062 660218 119146 660454
rect 119382 660218 119414 660454
rect 118794 660134 119414 660218
rect 118794 659898 118826 660134
rect 119062 659898 119146 660134
rect 119382 659898 119414 660134
rect 118794 624454 119414 659898
rect 118794 624218 118826 624454
rect 119062 624218 119146 624454
rect 119382 624218 119414 624454
rect 118794 624134 119414 624218
rect 118794 623898 118826 624134
rect 119062 623898 119146 624134
rect 119382 623898 119414 624134
rect 118794 588454 119414 623898
rect 118794 588218 118826 588454
rect 119062 588218 119146 588454
rect 119382 588218 119414 588454
rect 118794 588134 119414 588218
rect 118794 587898 118826 588134
rect 119062 587898 119146 588134
rect 119382 587898 119414 588134
rect 118794 552454 119414 587898
rect 118794 552218 118826 552454
rect 119062 552218 119146 552454
rect 119382 552218 119414 552454
rect 118794 552134 119414 552218
rect 118794 551898 118826 552134
rect 119062 551898 119146 552134
rect 119382 551898 119414 552134
rect 118794 516454 119414 551898
rect 118794 516218 118826 516454
rect 119062 516218 119146 516454
rect 119382 516218 119414 516454
rect 118794 516134 119414 516218
rect 118794 515898 118826 516134
rect 119062 515898 119146 516134
rect 119382 515898 119414 516134
rect 118794 480454 119414 515898
rect 118794 480218 118826 480454
rect 119062 480218 119146 480454
rect 119382 480218 119414 480454
rect 118794 480134 119414 480218
rect 118794 479898 118826 480134
rect 119062 479898 119146 480134
rect 119382 479898 119414 480134
rect 118794 444454 119414 479898
rect 118794 444218 118826 444454
rect 119062 444218 119146 444454
rect 119382 444218 119414 444454
rect 118794 444134 119414 444218
rect 118794 443898 118826 444134
rect 119062 443898 119146 444134
rect 119382 443898 119414 444134
rect 118794 408454 119414 443898
rect 118794 408218 118826 408454
rect 119062 408218 119146 408454
rect 119382 408218 119414 408454
rect 118794 408134 119414 408218
rect 118794 407898 118826 408134
rect 119062 407898 119146 408134
rect 119382 407898 119414 408134
rect 118794 372454 119414 407898
rect 118794 372218 118826 372454
rect 119062 372218 119146 372454
rect 119382 372218 119414 372454
rect 118794 372134 119414 372218
rect 118794 371898 118826 372134
rect 119062 371898 119146 372134
rect 119382 371898 119414 372134
rect 118794 336454 119414 371898
rect 118794 336218 118826 336454
rect 119062 336218 119146 336454
rect 119382 336218 119414 336454
rect 118794 336134 119414 336218
rect 118794 335898 118826 336134
rect 119062 335898 119146 336134
rect 119382 335898 119414 336134
rect 118794 300454 119414 335898
rect 118794 300218 118826 300454
rect 119062 300218 119146 300454
rect 119382 300218 119414 300454
rect 118794 300134 119414 300218
rect 118794 299898 118826 300134
rect 119062 299898 119146 300134
rect 119382 299898 119414 300134
rect 118794 264454 119414 299898
rect 118794 264218 118826 264454
rect 119062 264218 119146 264454
rect 119382 264218 119414 264454
rect 118794 264134 119414 264218
rect 118794 263898 118826 264134
rect 119062 263898 119146 264134
rect 119382 263898 119414 264134
rect 118555 263668 118621 263669
rect 118555 263604 118556 263668
rect 118620 263604 118621 263668
rect 118555 263603 118621 263604
rect 114294 259718 114326 259954
rect 114562 259718 114646 259954
rect 114882 259718 114914 259954
rect 114294 259634 114914 259718
rect 114294 259398 114326 259634
rect 114562 259398 114646 259634
rect 114882 259398 114914 259634
rect 114294 223954 114914 259398
rect 114294 223718 114326 223954
rect 114562 223718 114646 223954
rect 114882 223718 114914 223954
rect 114294 223634 114914 223718
rect 114294 223398 114326 223634
rect 114562 223398 114646 223634
rect 114882 223398 114914 223634
rect 114139 199068 114205 199069
rect 114139 199004 114140 199068
rect 114204 199004 114205 199068
rect 114139 199003 114205 199004
rect 113955 195396 114021 195397
rect 113955 195332 113956 195396
rect 114020 195332 114021 195396
rect 113955 195331 114021 195332
rect 111563 190228 111629 190229
rect 111563 190164 111564 190228
rect 111628 190164 111629 190228
rect 111563 190163 111629 190164
rect 111379 185604 111445 185605
rect 111379 185540 111380 185604
rect 111444 185540 111445 185604
rect 111379 185539 111445 185540
rect 109794 183218 109826 183454
rect 110062 183218 110146 183454
rect 110382 183218 110414 183454
rect 109794 183134 110414 183218
rect 109794 182898 109826 183134
rect 110062 182898 110146 183134
rect 110382 182898 110414 183134
rect 109794 147454 110414 182898
rect 111195 148748 111261 148749
rect 111195 148684 111196 148748
rect 111260 148684 111261 148748
rect 111195 148683 111261 148684
rect 109794 147218 109826 147454
rect 110062 147218 110146 147454
rect 110382 147218 110414 147454
rect 109794 147134 110414 147218
rect 109794 146898 109826 147134
rect 110062 146898 110146 147134
rect 110382 146898 110414 147134
rect 109794 111454 110414 146898
rect 111011 144260 111077 144261
rect 111011 144196 111012 144260
rect 111076 144196 111077 144260
rect 111011 144195 111077 144196
rect 109794 111218 109826 111454
rect 110062 111218 110146 111454
rect 110382 111218 110414 111454
rect 109794 111134 110414 111218
rect 109794 110898 109826 111134
rect 110062 110898 110146 111134
rect 110382 110898 110414 111134
rect 109794 75454 110414 110898
rect 111014 79389 111074 144195
rect 111011 79388 111077 79389
rect 111011 79324 111012 79388
rect 111076 79324 111077 79388
rect 111011 79323 111077 79324
rect 109794 75218 109826 75454
rect 110062 75218 110146 75454
rect 110382 75218 110414 75454
rect 109794 75134 110414 75218
rect 109794 74898 109826 75134
rect 110062 74898 110146 75134
rect 110382 74898 110414 75134
rect 109539 70004 109605 70005
rect 109539 69940 109540 70004
rect 109604 69940 109605 70004
rect 109539 69939 109605 69940
rect 106043 68508 106109 68509
rect 106043 68444 106044 68508
rect 106108 68444 106109 68508
rect 106043 68443 106109 68444
rect 105294 34718 105326 34954
rect 105562 34718 105646 34954
rect 105882 34718 105914 34954
rect 105294 34634 105914 34718
rect 105294 34398 105326 34634
rect 105562 34398 105646 34634
rect 105882 34398 105914 34634
rect 105294 -7066 105914 34398
rect 105294 -7302 105326 -7066
rect 105562 -7302 105646 -7066
rect 105882 -7302 105914 -7066
rect 105294 -7386 105914 -7302
rect 105294 -7622 105326 -7386
rect 105562 -7622 105646 -7386
rect 105882 -7622 105914 -7386
rect 105294 -7654 105914 -7622
rect 109794 39454 110414 74898
rect 111198 69733 111258 148683
rect 111382 74357 111442 185539
rect 111379 74356 111445 74357
rect 111379 74292 111380 74356
rect 111444 74292 111445 74356
rect 111379 74291 111445 74292
rect 111566 69869 111626 190163
rect 113771 187100 113837 187101
rect 113771 187036 113772 187100
rect 113836 187036 113837 187100
rect 113771 187035 113837 187036
rect 112851 184380 112917 184381
rect 112851 184316 112852 184380
rect 112916 184316 112917 184380
rect 112851 184315 112917 184316
rect 112667 148340 112733 148341
rect 112667 148276 112668 148340
rect 112732 148276 112733 148340
rect 112667 148275 112733 148276
rect 112670 80069 112730 148275
rect 112667 80068 112733 80069
rect 112667 80004 112668 80068
rect 112732 80004 112733 80068
rect 112667 80003 112733 80004
rect 112854 72997 112914 184315
rect 113035 177444 113101 177445
rect 113035 177380 113036 177444
rect 113100 177380 113101 177444
rect 113035 177379 113101 177380
rect 112851 72996 112917 72997
rect 112851 72932 112852 72996
rect 112916 72932 112917 72996
rect 112851 72931 112917 72932
rect 111563 69868 111629 69869
rect 111563 69804 111564 69868
rect 111628 69804 111629 69868
rect 111563 69803 111629 69804
rect 111195 69732 111261 69733
rect 111195 69668 111196 69732
rect 111260 69668 111261 69732
rect 111195 69667 111261 69668
rect 113038 66061 113098 177379
rect 113587 136100 113653 136101
rect 113587 136036 113588 136100
rect 113652 136036 113653 136100
rect 113587 136035 113653 136036
rect 113035 66060 113101 66061
rect 113035 65996 113036 66060
rect 113100 65996 113101 66060
rect 113035 65995 113101 65996
rect 113590 64701 113650 136035
rect 113774 76805 113834 187035
rect 113771 76804 113837 76805
rect 113771 76740 113772 76804
rect 113836 76740 113837 76804
rect 113771 76739 113837 76740
rect 113958 75717 114018 195331
rect 113955 75716 114021 75717
rect 113955 75652 113956 75716
rect 114020 75652 114021 75716
rect 113955 75651 114021 75652
rect 114142 75581 114202 199003
rect 114294 187954 114914 223398
rect 117083 195260 117149 195261
rect 117083 195196 117084 195260
rect 117148 195196 117149 195260
rect 117083 195195 117149 195196
rect 116899 189140 116965 189141
rect 116899 189076 116900 189140
rect 116964 189076 116965 189140
rect 116899 189075 116965 189076
rect 114294 187718 114326 187954
rect 114562 187718 114646 187954
rect 114882 187718 114914 187954
rect 114294 187634 114914 187718
rect 114294 187398 114326 187634
rect 114562 187398 114646 187634
rect 114882 187398 114914 187634
rect 114294 151954 114914 187398
rect 114294 151718 114326 151954
rect 114562 151718 114646 151954
rect 114882 151718 114914 151954
rect 114294 151634 114914 151718
rect 114294 151398 114326 151634
rect 114562 151398 114646 151634
rect 114882 151398 114914 151634
rect 114294 115954 114914 151398
rect 115611 144124 115677 144125
rect 115611 144060 115612 144124
rect 115676 144060 115677 144124
rect 115611 144059 115677 144060
rect 115427 141676 115493 141677
rect 115427 141612 115428 141676
rect 115492 141612 115493 141676
rect 115427 141611 115493 141612
rect 114294 115718 114326 115954
rect 114562 115718 114646 115954
rect 114882 115718 114914 115954
rect 114294 115634 114914 115718
rect 114294 115398 114326 115634
rect 114562 115398 114646 115634
rect 114882 115398 114914 115634
rect 114294 79954 114914 115398
rect 115430 80341 115490 141611
rect 115427 80340 115493 80341
rect 115427 80276 115428 80340
rect 115492 80276 115493 80340
rect 115427 80275 115493 80276
rect 115614 80205 115674 144059
rect 115795 140588 115861 140589
rect 115795 140524 115796 140588
rect 115860 140524 115861 140588
rect 115795 140523 115861 140524
rect 115611 80204 115677 80205
rect 115611 80140 115612 80204
rect 115676 80140 115677 80204
rect 115611 80139 115677 80140
rect 114294 79718 114326 79954
rect 114562 79718 114646 79954
rect 114882 79718 114914 79954
rect 114294 79634 114914 79718
rect 114294 79398 114326 79634
rect 114562 79398 114646 79634
rect 114882 79398 114914 79634
rect 114139 75580 114205 75581
rect 114139 75516 114140 75580
rect 114204 75516 114205 75580
rect 114139 75515 114205 75516
rect 113587 64700 113653 64701
rect 113587 64636 113588 64700
rect 113652 64636 113653 64700
rect 113587 64635 113653 64636
rect 109794 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 110414 39454
rect 109794 39134 110414 39218
rect 109794 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 110414 39134
rect 109794 3454 110414 38898
rect 109794 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 110414 3454
rect 109794 3134 110414 3218
rect 109794 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 110414 3134
rect 109794 -346 110414 2898
rect 109794 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 110414 -346
rect 109794 -666 110414 -582
rect 109794 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 110414 -666
rect 109794 -7654 110414 -902
rect 114294 43954 114914 79398
rect 115798 72725 115858 140523
rect 116715 140452 116781 140453
rect 116715 140388 116716 140452
rect 116780 140388 116781 140452
rect 116715 140387 116781 140388
rect 116531 138820 116597 138821
rect 116531 138756 116532 138820
rect 116596 138756 116597 138820
rect 116531 138755 116597 138756
rect 116534 79117 116594 138755
rect 116531 79116 116597 79117
rect 116531 79052 116532 79116
rect 116596 79052 116597 79116
rect 116531 79051 116597 79052
rect 116718 73949 116778 140387
rect 116902 76669 116962 189075
rect 116899 76668 116965 76669
rect 116899 76604 116900 76668
rect 116964 76604 116965 76668
rect 116899 76603 116965 76604
rect 116715 73948 116781 73949
rect 116715 73884 116716 73948
rect 116780 73884 116781 73948
rect 116715 73883 116781 73884
rect 117086 73813 117146 195195
rect 117267 191316 117333 191317
rect 117267 191252 117268 191316
rect 117332 191252 117333 191316
rect 117267 191251 117333 191252
rect 117270 190093 117330 191251
rect 117267 190092 117333 190093
rect 117267 190028 117268 190092
rect 117332 190028 117333 190092
rect 117267 190027 117333 190028
rect 117270 189141 117330 190027
rect 117267 189140 117333 189141
rect 117267 189076 117268 189140
rect 117332 189076 117333 189140
rect 117267 189075 117333 189076
rect 118558 143173 118618 263603
rect 118794 262000 119414 263898
rect 123294 707718 123914 711590
rect 123294 707482 123326 707718
rect 123562 707482 123646 707718
rect 123882 707482 123914 707718
rect 123294 707398 123914 707482
rect 123294 707162 123326 707398
rect 123562 707162 123646 707398
rect 123882 707162 123914 707398
rect 123294 700954 123914 707162
rect 123294 700718 123326 700954
rect 123562 700718 123646 700954
rect 123882 700718 123914 700954
rect 123294 700634 123914 700718
rect 123294 700398 123326 700634
rect 123562 700398 123646 700634
rect 123882 700398 123914 700634
rect 123294 664954 123914 700398
rect 123294 664718 123326 664954
rect 123562 664718 123646 664954
rect 123882 664718 123914 664954
rect 123294 664634 123914 664718
rect 123294 664398 123326 664634
rect 123562 664398 123646 664634
rect 123882 664398 123914 664634
rect 123294 628954 123914 664398
rect 123294 628718 123326 628954
rect 123562 628718 123646 628954
rect 123882 628718 123914 628954
rect 123294 628634 123914 628718
rect 123294 628398 123326 628634
rect 123562 628398 123646 628634
rect 123882 628398 123914 628634
rect 123294 592954 123914 628398
rect 123294 592718 123326 592954
rect 123562 592718 123646 592954
rect 123882 592718 123914 592954
rect 123294 592634 123914 592718
rect 123294 592398 123326 592634
rect 123562 592398 123646 592634
rect 123882 592398 123914 592634
rect 123294 556954 123914 592398
rect 123294 556718 123326 556954
rect 123562 556718 123646 556954
rect 123882 556718 123914 556954
rect 123294 556634 123914 556718
rect 123294 556398 123326 556634
rect 123562 556398 123646 556634
rect 123882 556398 123914 556634
rect 123294 520954 123914 556398
rect 123294 520718 123326 520954
rect 123562 520718 123646 520954
rect 123882 520718 123914 520954
rect 123294 520634 123914 520718
rect 123294 520398 123326 520634
rect 123562 520398 123646 520634
rect 123882 520398 123914 520634
rect 123294 484954 123914 520398
rect 123294 484718 123326 484954
rect 123562 484718 123646 484954
rect 123882 484718 123914 484954
rect 123294 484634 123914 484718
rect 123294 484398 123326 484634
rect 123562 484398 123646 484634
rect 123882 484398 123914 484634
rect 123294 448954 123914 484398
rect 123294 448718 123326 448954
rect 123562 448718 123646 448954
rect 123882 448718 123914 448954
rect 123294 448634 123914 448718
rect 123294 448398 123326 448634
rect 123562 448398 123646 448634
rect 123882 448398 123914 448634
rect 123294 412954 123914 448398
rect 123294 412718 123326 412954
rect 123562 412718 123646 412954
rect 123882 412718 123914 412954
rect 123294 412634 123914 412718
rect 123294 412398 123326 412634
rect 123562 412398 123646 412634
rect 123882 412398 123914 412634
rect 123294 376954 123914 412398
rect 123294 376718 123326 376954
rect 123562 376718 123646 376954
rect 123882 376718 123914 376954
rect 123294 376634 123914 376718
rect 123294 376398 123326 376634
rect 123562 376398 123646 376634
rect 123882 376398 123914 376634
rect 123294 340954 123914 376398
rect 123294 340718 123326 340954
rect 123562 340718 123646 340954
rect 123882 340718 123914 340954
rect 123294 340634 123914 340718
rect 123294 340398 123326 340634
rect 123562 340398 123646 340634
rect 123882 340398 123914 340634
rect 123294 304954 123914 340398
rect 123294 304718 123326 304954
rect 123562 304718 123646 304954
rect 123882 304718 123914 304954
rect 123294 304634 123914 304718
rect 123294 304398 123326 304634
rect 123562 304398 123646 304634
rect 123882 304398 123914 304634
rect 123294 268954 123914 304398
rect 123294 268718 123326 268954
rect 123562 268718 123646 268954
rect 123882 268718 123914 268954
rect 123294 268634 123914 268718
rect 123294 268398 123326 268634
rect 123562 268398 123646 268634
rect 123882 268398 123914 268634
rect 123294 262000 123914 268398
rect 127794 708678 128414 711590
rect 127794 708442 127826 708678
rect 128062 708442 128146 708678
rect 128382 708442 128414 708678
rect 127794 708358 128414 708442
rect 127794 708122 127826 708358
rect 128062 708122 128146 708358
rect 128382 708122 128414 708358
rect 127794 669454 128414 708122
rect 127794 669218 127826 669454
rect 128062 669218 128146 669454
rect 128382 669218 128414 669454
rect 127794 669134 128414 669218
rect 127794 668898 127826 669134
rect 128062 668898 128146 669134
rect 128382 668898 128414 669134
rect 127794 633454 128414 668898
rect 127794 633218 127826 633454
rect 128062 633218 128146 633454
rect 128382 633218 128414 633454
rect 127794 633134 128414 633218
rect 127794 632898 127826 633134
rect 128062 632898 128146 633134
rect 128382 632898 128414 633134
rect 127794 597454 128414 632898
rect 127794 597218 127826 597454
rect 128062 597218 128146 597454
rect 128382 597218 128414 597454
rect 127794 597134 128414 597218
rect 127794 596898 127826 597134
rect 128062 596898 128146 597134
rect 128382 596898 128414 597134
rect 127794 561454 128414 596898
rect 127794 561218 127826 561454
rect 128062 561218 128146 561454
rect 128382 561218 128414 561454
rect 127794 561134 128414 561218
rect 127794 560898 127826 561134
rect 128062 560898 128146 561134
rect 128382 560898 128414 561134
rect 127794 525454 128414 560898
rect 127794 525218 127826 525454
rect 128062 525218 128146 525454
rect 128382 525218 128414 525454
rect 127794 525134 128414 525218
rect 127794 524898 127826 525134
rect 128062 524898 128146 525134
rect 128382 524898 128414 525134
rect 127794 489454 128414 524898
rect 127794 489218 127826 489454
rect 128062 489218 128146 489454
rect 128382 489218 128414 489454
rect 127794 489134 128414 489218
rect 127794 488898 127826 489134
rect 128062 488898 128146 489134
rect 128382 488898 128414 489134
rect 127794 453454 128414 488898
rect 127794 453218 127826 453454
rect 128062 453218 128146 453454
rect 128382 453218 128414 453454
rect 127794 453134 128414 453218
rect 127794 452898 127826 453134
rect 128062 452898 128146 453134
rect 128382 452898 128414 453134
rect 127794 417454 128414 452898
rect 127794 417218 127826 417454
rect 128062 417218 128146 417454
rect 128382 417218 128414 417454
rect 127794 417134 128414 417218
rect 127794 416898 127826 417134
rect 128062 416898 128146 417134
rect 128382 416898 128414 417134
rect 127794 381454 128414 416898
rect 127794 381218 127826 381454
rect 128062 381218 128146 381454
rect 128382 381218 128414 381454
rect 127794 381134 128414 381218
rect 127794 380898 127826 381134
rect 128062 380898 128146 381134
rect 128382 380898 128414 381134
rect 127794 345454 128414 380898
rect 127794 345218 127826 345454
rect 128062 345218 128146 345454
rect 128382 345218 128414 345454
rect 127794 345134 128414 345218
rect 127794 344898 127826 345134
rect 128062 344898 128146 345134
rect 128382 344898 128414 345134
rect 127794 309454 128414 344898
rect 127794 309218 127826 309454
rect 128062 309218 128146 309454
rect 128382 309218 128414 309454
rect 127794 309134 128414 309218
rect 127794 308898 127826 309134
rect 128062 308898 128146 309134
rect 128382 308898 128414 309134
rect 127794 273454 128414 308898
rect 127794 273218 127826 273454
rect 128062 273218 128146 273454
rect 128382 273218 128414 273454
rect 127794 273134 128414 273218
rect 127794 272898 127826 273134
rect 128062 272898 128146 273134
rect 128382 272898 128414 273134
rect 127794 262000 128414 272898
rect 132294 709638 132914 711590
rect 132294 709402 132326 709638
rect 132562 709402 132646 709638
rect 132882 709402 132914 709638
rect 132294 709318 132914 709402
rect 132294 709082 132326 709318
rect 132562 709082 132646 709318
rect 132882 709082 132914 709318
rect 132294 673954 132914 709082
rect 132294 673718 132326 673954
rect 132562 673718 132646 673954
rect 132882 673718 132914 673954
rect 132294 673634 132914 673718
rect 132294 673398 132326 673634
rect 132562 673398 132646 673634
rect 132882 673398 132914 673634
rect 132294 637954 132914 673398
rect 132294 637718 132326 637954
rect 132562 637718 132646 637954
rect 132882 637718 132914 637954
rect 132294 637634 132914 637718
rect 132294 637398 132326 637634
rect 132562 637398 132646 637634
rect 132882 637398 132914 637634
rect 132294 601954 132914 637398
rect 132294 601718 132326 601954
rect 132562 601718 132646 601954
rect 132882 601718 132914 601954
rect 132294 601634 132914 601718
rect 132294 601398 132326 601634
rect 132562 601398 132646 601634
rect 132882 601398 132914 601634
rect 132294 565954 132914 601398
rect 132294 565718 132326 565954
rect 132562 565718 132646 565954
rect 132882 565718 132914 565954
rect 132294 565634 132914 565718
rect 132294 565398 132326 565634
rect 132562 565398 132646 565634
rect 132882 565398 132914 565634
rect 132294 529954 132914 565398
rect 132294 529718 132326 529954
rect 132562 529718 132646 529954
rect 132882 529718 132914 529954
rect 132294 529634 132914 529718
rect 132294 529398 132326 529634
rect 132562 529398 132646 529634
rect 132882 529398 132914 529634
rect 132294 493954 132914 529398
rect 132294 493718 132326 493954
rect 132562 493718 132646 493954
rect 132882 493718 132914 493954
rect 132294 493634 132914 493718
rect 132294 493398 132326 493634
rect 132562 493398 132646 493634
rect 132882 493398 132914 493634
rect 132294 457954 132914 493398
rect 132294 457718 132326 457954
rect 132562 457718 132646 457954
rect 132882 457718 132914 457954
rect 132294 457634 132914 457718
rect 132294 457398 132326 457634
rect 132562 457398 132646 457634
rect 132882 457398 132914 457634
rect 132294 421954 132914 457398
rect 132294 421718 132326 421954
rect 132562 421718 132646 421954
rect 132882 421718 132914 421954
rect 132294 421634 132914 421718
rect 132294 421398 132326 421634
rect 132562 421398 132646 421634
rect 132882 421398 132914 421634
rect 132294 385954 132914 421398
rect 132294 385718 132326 385954
rect 132562 385718 132646 385954
rect 132882 385718 132914 385954
rect 132294 385634 132914 385718
rect 132294 385398 132326 385634
rect 132562 385398 132646 385634
rect 132882 385398 132914 385634
rect 132294 349954 132914 385398
rect 132294 349718 132326 349954
rect 132562 349718 132646 349954
rect 132882 349718 132914 349954
rect 132294 349634 132914 349718
rect 132294 349398 132326 349634
rect 132562 349398 132646 349634
rect 132882 349398 132914 349634
rect 132294 313954 132914 349398
rect 132294 313718 132326 313954
rect 132562 313718 132646 313954
rect 132882 313718 132914 313954
rect 132294 313634 132914 313718
rect 132294 313398 132326 313634
rect 132562 313398 132646 313634
rect 132882 313398 132914 313634
rect 132294 277954 132914 313398
rect 132294 277718 132326 277954
rect 132562 277718 132646 277954
rect 132882 277718 132914 277954
rect 132294 277634 132914 277718
rect 132294 277398 132326 277634
rect 132562 277398 132646 277634
rect 132882 277398 132914 277634
rect 132294 262000 132914 277398
rect 136794 710598 137414 711590
rect 136794 710362 136826 710598
rect 137062 710362 137146 710598
rect 137382 710362 137414 710598
rect 136794 710278 137414 710362
rect 136794 710042 136826 710278
rect 137062 710042 137146 710278
rect 137382 710042 137414 710278
rect 136794 678454 137414 710042
rect 136794 678218 136826 678454
rect 137062 678218 137146 678454
rect 137382 678218 137414 678454
rect 136794 678134 137414 678218
rect 136794 677898 136826 678134
rect 137062 677898 137146 678134
rect 137382 677898 137414 678134
rect 136794 642454 137414 677898
rect 136794 642218 136826 642454
rect 137062 642218 137146 642454
rect 137382 642218 137414 642454
rect 136794 642134 137414 642218
rect 136794 641898 136826 642134
rect 137062 641898 137146 642134
rect 137382 641898 137414 642134
rect 136794 606454 137414 641898
rect 136794 606218 136826 606454
rect 137062 606218 137146 606454
rect 137382 606218 137414 606454
rect 136794 606134 137414 606218
rect 136794 605898 136826 606134
rect 137062 605898 137146 606134
rect 137382 605898 137414 606134
rect 136794 570454 137414 605898
rect 136794 570218 136826 570454
rect 137062 570218 137146 570454
rect 137382 570218 137414 570454
rect 136794 570134 137414 570218
rect 136794 569898 136826 570134
rect 137062 569898 137146 570134
rect 137382 569898 137414 570134
rect 136794 534454 137414 569898
rect 136794 534218 136826 534454
rect 137062 534218 137146 534454
rect 137382 534218 137414 534454
rect 136794 534134 137414 534218
rect 136794 533898 136826 534134
rect 137062 533898 137146 534134
rect 137382 533898 137414 534134
rect 136794 498454 137414 533898
rect 136794 498218 136826 498454
rect 137062 498218 137146 498454
rect 137382 498218 137414 498454
rect 136794 498134 137414 498218
rect 136794 497898 136826 498134
rect 137062 497898 137146 498134
rect 137382 497898 137414 498134
rect 136794 462454 137414 497898
rect 136794 462218 136826 462454
rect 137062 462218 137146 462454
rect 137382 462218 137414 462454
rect 136794 462134 137414 462218
rect 136794 461898 136826 462134
rect 137062 461898 137146 462134
rect 137382 461898 137414 462134
rect 136794 426454 137414 461898
rect 136794 426218 136826 426454
rect 137062 426218 137146 426454
rect 137382 426218 137414 426454
rect 136794 426134 137414 426218
rect 136794 425898 136826 426134
rect 137062 425898 137146 426134
rect 137382 425898 137414 426134
rect 136794 390454 137414 425898
rect 136794 390218 136826 390454
rect 137062 390218 137146 390454
rect 137382 390218 137414 390454
rect 136794 390134 137414 390218
rect 136794 389898 136826 390134
rect 137062 389898 137146 390134
rect 137382 389898 137414 390134
rect 136794 354454 137414 389898
rect 136794 354218 136826 354454
rect 137062 354218 137146 354454
rect 137382 354218 137414 354454
rect 136794 354134 137414 354218
rect 136794 353898 136826 354134
rect 137062 353898 137146 354134
rect 137382 353898 137414 354134
rect 136794 318454 137414 353898
rect 136794 318218 136826 318454
rect 137062 318218 137146 318454
rect 137382 318218 137414 318454
rect 136794 318134 137414 318218
rect 136794 317898 136826 318134
rect 137062 317898 137146 318134
rect 137382 317898 137414 318134
rect 136794 282454 137414 317898
rect 136794 282218 136826 282454
rect 137062 282218 137146 282454
rect 137382 282218 137414 282454
rect 136794 282134 137414 282218
rect 136794 281898 136826 282134
rect 137062 281898 137146 282134
rect 137382 281898 137414 282134
rect 136794 262000 137414 281898
rect 141294 711558 141914 711590
rect 141294 711322 141326 711558
rect 141562 711322 141646 711558
rect 141882 711322 141914 711558
rect 141294 711238 141914 711322
rect 141294 711002 141326 711238
rect 141562 711002 141646 711238
rect 141882 711002 141914 711238
rect 141294 682954 141914 711002
rect 141294 682718 141326 682954
rect 141562 682718 141646 682954
rect 141882 682718 141914 682954
rect 141294 682634 141914 682718
rect 141294 682398 141326 682634
rect 141562 682398 141646 682634
rect 141882 682398 141914 682634
rect 141294 646954 141914 682398
rect 141294 646718 141326 646954
rect 141562 646718 141646 646954
rect 141882 646718 141914 646954
rect 141294 646634 141914 646718
rect 141294 646398 141326 646634
rect 141562 646398 141646 646634
rect 141882 646398 141914 646634
rect 141294 610954 141914 646398
rect 141294 610718 141326 610954
rect 141562 610718 141646 610954
rect 141882 610718 141914 610954
rect 141294 610634 141914 610718
rect 141294 610398 141326 610634
rect 141562 610398 141646 610634
rect 141882 610398 141914 610634
rect 141294 574954 141914 610398
rect 141294 574718 141326 574954
rect 141562 574718 141646 574954
rect 141882 574718 141914 574954
rect 141294 574634 141914 574718
rect 141294 574398 141326 574634
rect 141562 574398 141646 574634
rect 141882 574398 141914 574634
rect 141294 538954 141914 574398
rect 141294 538718 141326 538954
rect 141562 538718 141646 538954
rect 141882 538718 141914 538954
rect 141294 538634 141914 538718
rect 141294 538398 141326 538634
rect 141562 538398 141646 538634
rect 141882 538398 141914 538634
rect 141294 502954 141914 538398
rect 141294 502718 141326 502954
rect 141562 502718 141646 502954
rect 141882 502718 141914 502954
rect 141294 502634 141914 502718
rect 141294 502398 141326 502634
rect 141562 502398 141646 502634
rect 141882 502398 141914 502634
rect 141294 466954 141914 502398
rect 141294 466718 141326 466954
rect 141562 466718 141646 466954
rect 141882 466718 141914 466954
rect 141294 466634 141914 466718
rect 141294 466398 141326 466634
rect 141562 466398 141646 466634
rect 141882 466398 141914 466634
rect 141294 430954 141914 466398
rect 141294 430718 141326 430954
rect 141562 430718 141646 430954
rect 141882 430718 141914 430954
rect 141294 430634 141914 430718
rect 141294 430398 141326 430634
rect 141562 430398 141646 430634
rect 141882 430398 141914 430634
rect 141294 394954 141914 430398
rect 141294 394718 141326 394954
rect 141562 394718 141646 394954
rect 141882 394718 141914 394954
rect 141294 394634 141914 394718
rect 141294 394398 141326 394634
rect 141562 394398 141646 394634
rect 141882 394398 141914 394634
rect 141294 358954 141914 394398
rect 141294 358718 141326 358954
rect 141562 358718 141646 358954
rect 141882 358718 141914 358954
rect 141294 358634 141914 358718
rect 141294 358398 141326 358634
rect 141562 358398 141646 358634
rect 141882 358398 141914 358634
rect 141294 322954 141914 358398
rect 141294 322718 141326 322954
rect 141562 322718 141646 322954
rect 141882 322718 141914 322954
rect 141294 322634 141914 322718
rect 141294 322398 141326 322634
rect 141562 322398 141646 322634
rect 141882 322398 141914 322634
rect 141294 286954 141914 322398
rect 141294 286718 141326 286954
rect 141562 286718 141646 286954
rect 141882 286718 141914 286954
rect 141294 286634 141914 286718
rect 141294 286398 141326 286634
rect 141562 286398 141646 286634
rect 141882 286398 141914 286634
rect 141294 262000 141914 286398
rect 145794 704838 146414 711590
rect 145794 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 146414 704838
rect 145794 704518 146414 704602
rect 145794 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 146414 704518
rect 145794 687454 146414 704282
rect 145794 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 146414 687454
rect 145794 687134 146414 687218
rect 145794 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 146414 687134
rect 145794 651454 146414 686898
rect 145794 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 146414 651454
rect 145794 651134 146414 651218
rect 145794 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 146414 651134
rect 145794 615454 146414 650898
rect 145794 615218 145826 615454
rect 146062 615218 146146 615454
rect 146382 615218 146414 615454
rect 145794 615134 146414 615218
rect 145794 614898 145826 615134
rect 146062 614898 146146 615134
rect 146382 614898 146414 615134
rect 145794 579454 146414 614898
rect 145794 579218 145826 579454
rect 146062 579218 146146 579454
rect 146382 579218 146414 579454
rect 145794 579134 146414 579218
rect 145794 578898 145826 579134
rect 146062 578898 146146 579134
rect 146382 578898 146414 579134
rect 145794 543454 146414 578898
rect 145794 543218 145826 543454
rect 146062 543218 146146 543454
rect 146382 543218 146414 543454
rect 145794 543134 146414 543218
rect 145794 542898 145826 543134
rect 146062 542898 146146 543134
rect 146382 542898 146414 543134
rect 145794 507454 146414 542898
rect 145794 507218 145826 507454
rect 146062 507218 146146 507454
rect 146382 507218 146414 507454
rect 145794 507134 146414 507218
rect 145794 506898 145826 507134
rect 146062 506898 146146 507134
rect 146382 506898 146414 507134
rect 145794 471454 146414 506898
rect 145794 471218 145826 471454
rect 146062 471218 146146 471454
rect 146382 471218 146414 471454
rect 145794 471134 146414 471218
rect 145794 470898 145826 471134
rect 146062 470898 146146 471134
rect 146382 470898 146414 471134
rect 145794 435454 146414 470898
rect 145794 435218 145826 435454
rect 146062 435218 146146 435454
rect 146382 435218 146414 435454
rect 145794 435134 146414 435218
rect 145794 434898 145826 435134
rect 146062 434898 146146 435134
rect 146382 434898 146414 435134
rect 145794 399454 146414 434898
rect 145794 399218 145826 399454
rect 146062 399218 146146 399454
rect 146382 399218 146414 399454
rect 145794 399134 146414 399218
rect 145794 398898 145826 399134
rect 146062 398898 146146 399134
rect 146382 398898 146414 399134
rect 145794 363454 146414 398898
rect 145794 363218 145826 363454
rect 146062 363218 146146 363454
rect 146382 363218 146414 363454
rect 145794 363134 146414 363218
rect 145794 362898 145826 363134
rect 146062 362898 146146 363134
rect 146382 362898 146414 363134
rect 145794 327454 146414 362898
rect 145794 327218 145826 327454
rect 146062 327218 146146 327454
rect 146382 327218 146414 327454
rect 145794 327134 146414 327218
rect 145794 326898 145826 327134
rect 146062 326898 146146 327134
rect 146382 326898 146414 327134
rect 145794 291454 146414 326898
rect 145794 291218 145826 291454
rect 146062 291218 146146 291454
rect 146382 291218 146414 291454
rect 145794 291134 146414 291218
rect 145794 290898 145826 291134
rect 146062 290898 146146 291134
rect 146382 290898 146414 291134
rect 145794 262000 146414 290898
rect 150294 705798 150914 711590
rect 150294 705562 150326 705798
rect 150562 705562 150646 705798
rect 150882 705562 150914 705798
rect 150294 705478 150914 705562
rect 150294 705242 150326 705478
rect 150562 705242 150646 705478
rect 150882 705242 150914 705478
rect 150294 691954 150914 705242
rect 150294 691718 150326 691954
rect 150562 691718 150646 691954
rect 150882 691718 150914 691954
rect 150294 691634 150914 691718
rect 150294 691398 150326 691634
rect 150562 691398 150646 691634
rect 150882 691398 150914 691634
rect 150294 655954 150914 691398
rect 150294 655718 150326 655954
rect 150562 655718 150646 655954
rect 150882 655718 150914 655954
rect 150294 655634 150914 655718
rect 150294 655398 150326 655634
rect 150562 655398 150646 655634
rect 150882 655398 150914 655634
rect 150294 619954 150914 655398
rect 150294 619718 150326 619954
rect 150562 619718 150646 619954
rect 150882 619718 150914 619954
rect 150294 619634 150914 619718
rect 150294 619398 150326 619634
rect 150562 619398 150646 619634
rect 150882 619398 150914 619634
rect 150294 583954 150914 619398
rect 150294 583718 150326 583954
rect 150562 583718 150646 583954
rect 150882 583718 150914 583954
rect 150294 583634 150914 583718
rect 150294 583398 150326 583634
rect 150562 583398 150646 583634
rect 150882 583398 150914 583634
rect 150294 547954 150914 583398
rect 150294 547718 150326 547954
rect 150562 547718 150646 547954
rect 150882 547718 150914 547954
rect 150294 547634 150914 547718
rect 150294 547398 150326 547634
rect 150562 547398 150646 547634
rect 150882 547398 150914 547634
rect 150294 511954 150914 547398
rect 150294 511718 150326 511954
rect 150562 511718 150646 511954
rect 150882 511718 150914 511954
rect 150294 511634 150914 511718
rect 150294 511398 150326 511634
rect 150562 511398 150646 511634
rect 150882 511398 150914 511634
rect 150294 475954 150914 511398
rect 150294 475718 150326 475954
rect 150562 475718 150646 475954
rect 150882 475718 150914 475954
rect 150294 475634 150914 475718
rect 150294 475398 150326 475634
rect 150562 475398 150646 475634
rect 150882 475398 150914 475634
rect 150294 439954 150914 475398
rect 150294 439718 150326 439954
rect 150562 439718 150646 439954
rect 150882 439718 150914 439954
rect 150294 439634 150914 439718
rect 150294 439398 150326 439634
rect 150562 439398 150646 439634
rect 150882 439398 150914 439634
rect 150294 403954 150914 439398
rect 150294 403718 150326 403954
rect 150562 403718 150646 403954
rect 150882 403718 150914 403954
rect 150294 403634 150914 403718
rect 150294 403398 150326 403634
rect 150562 403398 150646 403634
rect 150882 403398 150914 403634
rect 150294 367954 150914 403398
rect 150294 367718 150326 367954
rect 150562 367718 150646 367954
rect 150882 367718 150914 367954
rect 150294 367634 150914 367718
rect 150294 367398 150326 367634
rect 150562 367398 150646 367634
rect 150882 367398 150914 367634
rect 150294 331954 150914 367398
rect 150294 331718 150326 331954
rect 150562 331718 150646 331954
rect 150882 331718 150914 331954
rect 150294 331634 150914 331718
rect 150294 331398 150326 331634
rect 150562 331398 150646 331634
rect 150882 331398 150914 331634
rect 150294 295954 150914 331398
rect 150294 295718 150326 295954
rect 150562 295718 150646 295954
rect 150882 295718 150914 295954
rect 150294 295634 150914 295718
rect 150294 295398 150326 295634
rect 150562 295398 150646 295634
rect 150882 295398 150914 295634
rect 150294 262000 150914 295398
rect 154794 706758 155414 711590
rect 154794 706522 154826 706758
rect 155062 706522 155146 706758
rect 155382 706522 155414 706758
rect 154794 706438 155414 706522
rect 154794 706202 154826 706438
rect 155062 706202 155146 706438
rect 155382 706202 155414 706438
rect 154794 696454 155414 706202
rect 154794 696218 154826 696454
rect 155062 696218 155146 696454
rect 155382 696218 155414 696454
rect 154794 696134 155414 696218
rect 154794 695898 154826 696134
rect 155062 695898 155146 696134
rect 155382 695898 155414 696134
rect 154794 660454 155414 695898
rect 154794 660218 154826 660454
rect 155062 660218 155146 660454
rect 155382 660218 155414 660454
rect 154794 660134 155414 660218
rect 154794 659898 154826 660134
rect 155062 659898 155146 660134
rect 155382 659898 155414 660134
rect 154794 624454 155414 659898
rect 154794 624218 154826 624454
rect 155062 624218 155146 624454
rect 155382 624218 155414 624454
rect 154794 624134 155414 624218
rect 154794 623898 154826 624134
rect 155062 623898 155146 624134
rect 155382 623898 155414 624134
rect 154794 588454 155414 623898
rect 154794 588218 154826 588454
rect 155062 588218 155146 588454
rect 155382 588218 155414 588454
rect 154794 588134 155414 588218
rect 154794 587898 154826 588134
rect 155062 587898 155146 588134
rect 155382 587898 155414 588134
rect 154794 552454 155414 587898
rect 154794 552218 154826 552454
rect 155062 552218 155146 552454
rect 155382 552218 155414 552454
rect 154794 552134 155414 552218
rect 154794 551898 154826 552134
rect 155062 551898 155146 552134
rect 155382 551898 155414 552134
rect 154794 516454 155414 551898
rect 154794 516218 154826 516454
rect 155062 516218 155146 516454
rect 155382 516218 155414 516454
rect 154794 516134 155414 516218
rect 154794 515898 154826 516134
rect 155062 515898 155146 516134
rect 155382 515898 155414 516134
rect 154794 480454 155414 515898
rect 154794 480218 154826 480454
rect 155062 480218 155146 480454
rect 155382 480218 155414 480454
rect 154794 480134 155414 480218
rect 154794 479898 154826 480134
rect 155062 479898 155146 480134
rect 155382 479898 155414 480134
rect 154794 444454 155414 479898
rect 154794 444218 154826 444454
rect 155062 444218 155146 444454
rect 155382 444218 155414 444454
rect 154794 444134 155414 444218
rect 154794 443898 154826 444134
rect 155062 443898 155146 444134
rect 155382 443898 155414 444134
rect 154794 408454 155414 443898
rect 154794 408218 154826 408454
rect 155062 408218 155146 408454
rect 155382 408218 155414 408454
rect 154794 408134 155414 408218
rect 154794 407898 154826 408134
rect 155062 407898 155146 408134
rect 155382 407898 155414 408134
rect 154794 372454 155414 407898
rect 154794 372218 154826 372454
rect 155062 372218 155146 372454
rect 155382 372218 155414 372454
rect 154794 372134 155414 372218
rect 154794 371898 154826 372134
rect 155062 371898 155146 372134
rect 155382 371898 155414 372134
rect 154794 336454 155414 371898
rect 154794 336218 154826 336454
rect 155062 336218 155146 336454
rect 155382 336218 155414 336454
rect 154794 336134 155414 336218
rect 154794 335898 154826 336134
rect 155062 335898 155146 336134
rect 155382 335898 155414 336134
rect 154794 300454 155414 335898
rect 154794 300218 154826 300454
rect 155062 300218 155146 300454
rect 155382 300218 155414 300454
rect 154794 300134 155414 300218
rect 154794 299898 154826 300134
rect 155062 299898 155146 300134
rect 155382 299898 155414 300134
rect 154794 264454 155414 299898
rect 154794 264218 154826 264454
rect 155062 264218 155146 264454
rect 155382 264218 155414 264454
rect 154794 264134 155414 264218
rect 154794 263898 154826 264134
rect 155062 263898 155146 264134
rect 155382 263898 155414 264134
rect 154794 262000 155414 263898
rect 159294 707718 159914 711590
rect 159294 707482 159326 707718
rect 159562 707482 159646 707718
rect 159882 707482 159914 707718
rect 159294 707398 159914 707482
rect 159294 707162 159326 707398
rect 159562 707162 159646 707398
rect 159882 707162 159914 707398
rect 159294 700954 159914 707162
rect 159294 700718 159326 700954
rect 159562 700718 159646 700954
rect 159882 700718 159914 700954
rect 159294 700634 159914 700718
rect 159294 700398 159326 700634
rect 159562 700398 159646 700634
rect 159882 700398 159914 700634
rect 159294 664954 159914 700398
rect 159294 664718 159326 664954
rect 159562 664718 159646 664954
rect 159882 664718 159914 664954
rect 159294 664634 159914 664718
rect 159294 664398 159326 664634
rect 159562 664398 159646 664634
rect 159882 664398 159914 664634
rect 159294 628954 159914 664398
rect 159294 628718 159326 628954
rect 159562 628718 159646 628954
rect 159882 628718 159914 628954
rect 159294 628634 159914 628718
rect 159294 628398 159326 628634
rect 159562 628398 159646 628634
rect 159882 628398 159914 628634
rect 159294 592954 159914 628398
rect 159294 592718 159326 592954
rect 159562 592718 159646 592954
rect 159882 592718 159914 592954
rect 159294 592634 159914 592718
rect 159294 592398 159326 592634
rect 159562 592398 159646 592634
rect 159882 592398 159914 592634
rect 159294 556954 159914 592398
rect 159294 556718 159326 556954
rect 159562 556718 159646 556954
rect 159882 556718 159914 556954
rect 159294 556634 159914 556718
rect 159294 556398 159326 556634
rect 159562 556398 159646 556634
rect 159882 556398 159914 556634
rect 159294 520954 159914 556398
rect 159294 520718 159326 520954
rect 159562 520718 159646 520954
rect 159882 520718 159914 520954
rect 159294 520634 159914 520718
rect 159294 520398 159326 520634
rect 159562 520398 159646 520634
rect 159882 520398 159914 520634
rect 159294 484954 159914 520398
rect 159294 484718 159326 484954
rect 159562 484718 159646 484954
rect 159882 484718 159914 484954
rect 159294 484634 159914 484718
rect 159294 484398 159326 484634
rect 159562 484398 159646 484634
rect 159882 484398 159914 484634
rect 159294 448954 159914 484398
rect 159294 448718 159326 448954
rect 159562 448718 159646 448954
rect 159882 448718 159914 448954
rect 159294 448634 159914 448718
rect 159294 448398 159326 448634
rect 159562 448398 159646 448634
rect 159882 448398 159914 448634
rect 159294 412954 159914 448398
rect 159294 412718 159326 412954
rect 159562 412718 159646 412954
rect 159882 412718 159914 412954
rect 159294 412634 159914 412718
rect 159294 412398 159326 412634
rect 159562 412398 159646 412634
rect 159882 412398 159914 412634
rect 159294 376954 159914 412398
rect 159294 376718 159326 376954
rect 159562 376718 159646 376954
rect 159882 376718 159914 376954
rect 159294 376634 159914 376718
rect 159294 376398 159326 376634
rect 159562 376398 159646 376634
rect 159882 376398 159914 376634
rect 159294 340954 159914 376398
rect 159294 340718 159326 340954
rect 159562 340718 159646 340954
rect 159882 340718 159914 340954
rect 159294 340634 159914 340718
rect 159294 340398 159326 340634
rect 159562 340398 159646 340634
rect 159882 340398 159914 340634
rect 159294 304954 159914 340398
rect 159294 304718 159326 304954
rect 159562 304718 159646 304954
rect 159882 304718 159914 304954
rect 159294 304634 159914 304718
rect 159294 304398 159326 304634
rect 159562 304398 159646 304634
rect 159882 304398 159914 304634
rect 159294 268954 159914 304398
rect 159294 268718 159326 268954
rect 159562 268718 159646 268954
rect 159882 268718 159914 268954
rect 159294 268634 159914 268718
rect 159294 268398 159326 268634
rect 159562 268398 159646 268634
rect 159882 268398 159914 268634
rect 159294 262000 159914 268398
rect 163794 708678 164414 711590
rect 163794 708442 163826 708678
rect 164062 708442 164146 708678
rect 164382 708442 164414 708678
rect 163794 708358 164414 708442
rect 163794 708122 163826 708358
rect 164062 708122 164146 708358
rect 164382 708122 164414 708358
rect 163794 669454 164414 708122
rect 163794 669218 163826 669454
rect 164062 669218 164146 669454
rect 164382 669218 164414 669454
rect 163794 669134 164414 669218
rect 163794 668898 163826 669134
rect 164062 668898 164146 669134
rect 164382 668898 164414 669134
rect 163794 633454 164414 668898
rect 163794 633218 163826 633454
rect 164062 633218 164146 633454
rect 164382 633218 164414 633454
rect 163794 633134 164414 633218
rect 163794 632898 163826 633134
rect 164062 632898 164146 633134
rect 164382 632898 164414 633134
rect 163794 597454 164414 632898
rect 163794 597218 163826 597454
rect 164062 597218 164146 597454
rect 164382 597218 164414 597454
rect 163794 597134 164414 597218
rect 163794 596898 163826 597134
rect 164062 596898 164146 597134
rect 164382 596898 164414 597134
rect 163794 561454 164414 596898
rect 163794 561218 163826 561454
rect 164062 561218 164146 561454
rect 164382 561218 164414 561454
rect 163794 561134 164414 561218
rect 163794 560898 163826 561134
rect 164062 560898 164146 561134
rect 164382 560898 164414 561134
rect 163794 525454 164414 560898
rect 163794 525218 163826 525454
rect 164062 525218 164146 525454
rect 164382 525218 164414 525454
rect 163794 525134 164414 525218
rect 163794 524898 163826 525134
rect 164062 524898 164146 525134
rect 164382 524898 164414 525134
rect 163794 489454 164414 524898
rect 163794 489218 163826 489454
rect 164062 489218 164146 489454
rect 164382 489218 164414 489454
rect 163794 489134 164414 489218
rect 163794 488898 163826 489134
rect 164062 488898 164146 489134
rect 164382 488898 164414 489134
rect 163794 453454 164414 488898
rect 163794 453218 163826 453454
rect 164062 453218 164146 453454
rect 164382 453218 164414 453454
rect 163794 453134 164414 453218
rect 163794 452898 163826 453134
rect 164062 452898 164146 453134
rect 164382 452898 164414 453134
rect 163794 417454 164414 452898
rect 163794 417218 163826 417454
rect 164062 417218 164146 417454
rect 164382 417218 164414 417454
rect 163794 417134 164414 417218
rect 163794 416898 163826 417134
rect 164062 416898 164146 417134
rect 164382 416898 164414 417134
rect 163794 381454 164414 416898
rect 163794 381218 163826 381454
rect 164062 381218 164146 381454
rect 164382 381218 164414 381454
rect 163794 381134 164414 381218
rect 163794 380898 163826 381134
rect 164062 380898 164146 381134
rect 164382 380898 164414 381134
rect 163794 345454 164414 380898
rect 163794 345218 163826 345454
rect 164062 345218 164146 345454
rect 164382 345218 164414 345454
rect 163794 345134 164414 345218
rect 163794 344898 163826 345134
rect 164062 344898 164146 345134
rect 164382 344898 164414 345134
rect 163794 309454 164414 344898
rect 163794 309218 163826 309454
rect 164062 309218 164146 309454
rect 164382 309218 164414 309454
rect 163794 309134 164414 309218
rect 163794 308898 163826 309134
rect 164062 308898 164146 309134
rect 164382 308898 164414 309134
rect 163794 273454 164414 308898
rect 163794 273218 163826 273454
rect 164062 273218 164146 273454
rect 164382 273218 164414 273454
rect 163794 273134 164414 273218
rect 163794 272898 163826 273134
rect 164062 272898 164146 273134
rect 164382 272898 164414 273134
rect 163794 262000 164414 272898
rect 168294 709638 168914 711590
rect 168294 709402 168326 709638
rect 168562 709402 168646 709638
rect 168882 709402 168914 709638
rect 168294 709318 168914 709402
rect 168294 709082 168326 709318
rect 168562 709082 168646 709318
rect 168882 709082 168914 709318
rect 168294 673954 168914 709082
rect 168294 673718 168326 673954
rect 168562 673718 168646 673954
rect 168882 673718 168914 673954
rect 168294 673634 168914 673718
rect 168294 673398 168326 673634
rect 168562 673398 168646 673634
rect 168882 673398 168914 673634
rect 168294 637954 168914 673398
rect 168294 637718 168326 637954
rect 168562 637718 168646 637954
rect 168882 637718 168914 637954
rect 168294 637634 168914 637718
rect 168294 637398 168326 637634
rect 168562 637398 168646 637634
rect 168882 637398 168914 637634
rect 168294 601954 168914 637398
rect 168294 601718 168326 601954
rect 168562 601718 168646 601954
rect 168882 601718 168914 601954
rect 168294 601634 168914 601718
rect 168294 601398 168326 601634
rect 168562 601398 168646 601634
rect 168882 601398 168914 601634
rect 168294 565954 168914 601398
rect 168294 565718 168326 565954
rect 168562 565718 168646 565954
rect 168882 565718 168914 565954
rect 168294 565634 168914 565718
rect 168294 565398 168326 565634
rect 168562 565398 168646 565634
rect 168882 565398 168914 565634
rect 168294 529954 168914 565398
rect 168294 529718 168326 529954
rect 168562 529718 168646 529954
rect 168882 529718 168914 529954
rect 168294 529634 168914 529718
rect 168294 529398 168326 529634
rect 168562 529398 168646 529634
rect 168882 529398 168914 529634
rect 168294 493954 168914 529398
rect 168294 493718 168326 493954
rect 168562 493718 168646 493954
rect 168882 493718 168914 493954
rect 168294 493634 168914 493718
rect 168294 493398 168326 493634
rect 168562 493398 168646 493634
rect 168882 493398 168914 493634
rect 168294 457954 168914 493398
rect 168294 457718 168326 457954
rect 168562 457718 168646 457954
rect 168882 457718 168914 457954
rect 168294 457634 168914 457718
rect 168294 457398 168326 457634
rect 168562 457398 168646 457634
rect 168882 457398 168914 457634
rect 168294 421954 168914 457398
rect 168294 421718 168326 421954
rect 168562 421718 168646 421954
rect 168882 421718 168914 421954
rect 168294 421634 168914 421718
rect 168294 421398 168326 421634
rect 168562 421398 168646 421634
rect 168882 421398 168914 421634
rect 168294 385954 168914 421398
rect 168294 385718 168326 385954
rect 168562 385718 168646 385954
rect 168882 385718 168914 385954
rect 168294 385634 168914 385718
rect 168294 385398 168326 385634
rect 168562 385398 168646 385634
rect 168882 385398 168914 385634
rect 168294 349954 168914 385398
rect 168294 349718 168326 349954
rect 168562 349718 168646 349954
rect 168882 349718 168914 349954
rect 168294 349634 168914 349718
rect 168294 349398 168326 349634
rect 168562 349398 168646 349634
rect 168882 349398 168914 349634
rect 168294 313954 168914 349398
rect 168294 313718 168326 313954
rect 168562 313718 168646 313954
rect 168882 313718 168914 313954
rect 168294 313634 168914 313718
rect 168294 313398 168326 313634
rect 168562 313398 168646 313634
rect 168882 313398 168914 313634
rect 168294 277954 168914 313398
rect 168294 277718 168326 277954
rect 168562 277718 168646 277954
rect 168882 277718 168914 277954
rect 168294 277634 168914 277718
rect 168294 277398 168326 277634
rect 168562 277398 168646 277634
rect 168882 277398 168914 277634
rect 168294 262000 168914 277398
rect 172794 710598 173414 711590
rect 172794 710362 172826 710598
rect 173062 710362 173146 710598
rect 173382 710362 173414 710598
rect 172794 710278 173414 710362
rect 172794 710042 172826 710278
rect 173062 710042 173146 710278
rect 173382 710042 173414 710278
rect 172794 678454 173414 710042
rect 172794 678218 172826 678454
rect 173062 678218 173146 678454
rect 173382 678218 173414 678454
rect 172794 678134 173414 678218
rect 172794 677898 172826 678134
rect 173062 677898 173146 678134
rect 173382 677898 173414 678134
rect 172794 642454 173414 677898
rect 172794 642218 172826 642454
rect 173062 642218 173146 642454
rect 173382 642218 173414 642454
rect 172794 642134 173414 642218
rect 172794 641898 172826 642134
rect 173062 641898 173146 642134
rect 173382 641898 173414 642134
rect 172794 606454 173414 641898
rect 172794 606218 172826 606454
rect 173062 606218 173146 606454
rect 173382 606218 173414 606454
rect 172794 606134 173414 606218
rect 172794 605898 172826 606134
rect 173062 605898 173146 606134
rect 173382 605898 173414 606134
rect 172794 570454 173414 605898
rect 172794 570218 172826 570454
rect 173062 570218 173146 570454
rect 173382 570218 173414 570454
rect 172794 570134 173414 570218
rect 172794 569898 172826 570134
rect 173062 569898 173146 570134
rect 173382 569898 173414 570134
rect 172794 534454 173414 569898
rect 172794 534218 172826 534454
rect 173062 534218 173146 534454
rect 173382 534218 173414 534454
rect 172794 534134 173414 534218
rect 172794 533898 172826 534134
rect 173062 533898 173146 534134
rect 173382 533898 173414 534134
rect 172794 498454 173414 533898
rect 172794 498218 172826 498454
rect 173062 498218 173146 498454
rect 173382 498218 173414 498454
rect 172794 498134 173414 498218
rect 172794 497898 172826 498134
rect 173062 497898 173146 498134
rect 173382 497898 173414 498134
rect 172794 462454 173414 497898
rect 172794 462218 172826 462454
rect 173062 462218 173146 462454
rect 173382 462218 173414 462454
rect 172794 462134 173414 462218
rect 172794 461898 172826 462134
rect 173062 461898 173146 462134
rect 173382 461898 173414 462134
rect 172794 426454 173414 461898
rect 172794 426218 172826 426454
rect 173062 426218 173146 426454
rect 173382 426218 173414 426454
rect 172794 426134 173414 426218
rect 172794 425898 172826 426134
rect 173062 425898 173146 426134
rect 173382 425898 173414 426134
rect 172794 390454 173414 425898
rect 172794 390218 172826 390454
rect 173062 390218 173146 390454
rect 173382 390218 173414 390454
rect 172794 390134 173414 390218
rect 172794 389898 172826 390134
rect 173062 389898 173146 390134
rect 173382 389898 173414 390134
rect 172794 354454 173414 389898
rect 172794 354218 172826 354454
rect 173062 354218 173146 354454
rect 173382 354218 173414 354454
rect 172794 354134 173414 354218
rect 172794 353898 172826 354134
rect 173062 353898 173146 354134
rect 173382 353898 173414 354134
rect 172794 318454 173414 353898
rect 172794 318218 172826 318454
rect 173062 318218 173146 318454
rect 173382 318218 173414 318454
rect 172794 318134 173414 318218
rect 172794 317898 172826 318134
rect 173062 317898 173146 318134
rect 173382 317898 173414 318134
rect 172794 282454 173414 317898
rect 172794 282218 172826 282454
rect 173062 282218 173146 282454
rect 173382 282218 173414 282454
rect 172794 282134 173414 282218
rect 172794 281898 172826 282134
rect 173062 281898 173146 282134
rect 173382 281898 173414 282134
rect 172794 262000 173414 281898
rect 177294 711558 177914 711590
rect 177294 711322 177326 711558
rect 177562 711322 177646 711558
rect 177882 711322 177914 711558
rect 177294 711238 177914 711322
rect 177294 711002 177326 711238
rect 177562 711002 177646 711238
rect 177882 711002 177914 711238
rect 177294 682954 177914 711002
rect 177294 682718 177326 682954
rect 177562 682718 177646 682954
rect 177882 682718 177914 682954
rect 177294 682634 177914 682718
rect 177294 682398 177326 682634
rect 177562 682398 177646 682634
rect 177882 682398 177914 682634
rect 177294 646954 177914 682398
rect 177294 646718 177326 646954
rect 177562 646718 177646 646954
rect 177882 646718 177914 646954
rect 177294 646634 177914 646718
rect 177294 646398 177326 646634
rect 177562 646398 177646 646634
rect 177882 646398 177914 646634
rect 177294 610954 177914 646398
rect 177294 610718 177326 610954
rect 177562 610718 177646 610954
rect 177882 610718 177914 610954
rect 177294 610634 177914 610718
rect 177294 610398 177326 610634
rect 177562 610398 177646 610634
rect 177882 610398 177914 610634
rect 177294 574954 177914 610398
rect 177294 574718 177326 574954
rect 177562 574718 177646 574954
rect 177882 574718 177914 574954
rect 177294 574634 177914 574718
rect 177294 574398 177326 574634
rect 177562 574398 177646 574634
rect 177882 574398 177914 574634
rect 177294 538954 177914 574398
rect 177294 538718 177326 538954
rect 177562 538718 177646 538954
rect 177882 538718 177914 538954
rect 177294 538634 177914 538718
rect 177294 538398 177326 538634
rect 177562 538398 177646 538634
rect 177882 538398 177914 538634
rect 177294 502954 177914 538398
rect 177294 502718 177326 502954
rect 177562 502718 177646 502954
rect 177882 502718 177914 502954
rect 177294 502634 177914 502718
rect 177294 502398 177326 502634
rect 177562 502398 177646 502634
rect 177882 502398 177914 502634
rect 177294 466954 177914 502398
rect 177294 466718 177326 466954
rect 177562 466718 177646 466954
rect 177882 466718 177914 466954
rect 177294 466634 177914 466718
rect 177294 466398 177326 466634
rect 177562 466398 177646 466634
rect 177882 466398 177914 466634
rect 177294 430954 177914 466398
rect 177294 430718 177326 430954
rect 177562 430718 177646 430954
rect 177882 430718 177914 430954
rect 177294 430634 177914 430718
rect 177294 430398 177326 430634
rect 177562 430398 177646 430634
rect 177882 430398 177914 430634
rect 177294 394954 177914 430398
rect 177294 394718 177326 394954
rect 177562 394718 177646 394954
rect 177882 394718 177914 394954
rect 177294 394634 177914 394718
rect 177294 394398 177326 394634
rect 177562 394398 177646 394634
rect 177882 394398 177914 394634
rect 177294 358954 177914 394398
rect 177294 358718 177326 358954
rect 177562 358718 177646 358954
rect 177882 358718 177914 358954
rect 177294 358634 177914 358718
rect 177294 358398 177326 358634
rect 177562 358398 177646 358634
rect 177882 358398 177914 358634
rect 177294 322954 177914 358398
rect 177294 322718 177326 322954
rect 177562 322718 177646 322954
rect 177882 322718 177914 322954
rect 177294 322634 177914 322718
rect 177294 322398 177326 322634
rect 177562 322398 177646 322634
rect 177882 322398 177914 322634
rect 177294 286954 177914 322398
rect 177294 286718 177326 286954
rect 177562 286718 177646 286954
rect 177882 286718 177914 286954
rect 177294 286634 177914 286718
rect 177294 286398 177326 286634
rect 177562 286398 177646 286634
rect 177882 286398 177914 286634
rect 177294 262000 177914 286398
rect 181794 704838 182414 711590
rect 181794 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 182414 704838
rect 181794 704518 182414 704602
rect 181794 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 182414 704518
rect 181794 687454 182414 704282
rect 181794 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 182414 687454
rect 181794 687134 182414 687218
rect 181794 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 182414 687134
rect 181794 651454 182414 686898
rect 181794 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 182414 651454
rect 181794 651134 182414 651218
rect 181794 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 182414 651134
rect 181794 615454 182414 650898
rect 181794 615218 181826 615454
rect 182062 615218 182146 615454
rect 182382 615218 182414 615454
rect 181794 615134 182414 615218
rect 181794 614898 181826 615134
rect 182062 614898 182146 615134
rect 182382 614898 182414 615134
rect 181794 579454 182414 614898
rect 181794 579218 181826 579454
rect 182062 579218 182146 579454
rect 182382 579218 182414 579454
rect 181794 579134 182414 579218
rect 181794 578898 181826 579134
rect 182062 578898 182146 579134
rect 182382 578898 182414 579134
rect 181794 543454 182414 578898
rect 181794 543218 181826 543454
rect 182062 543218 182146 543454
rect 182382 543218 182414 543454
rect 181794 543134 182414 543218
rect 181794 542898 181826 543134
rect 182062 542898 182146 543134
rect 182382 542898 182414 543134
rect 181794 507454 182414 542898
rect 181794 507218 181826 507454
rect 182062 507218 182146 507454
rect 182382 507218 182414 507454
rect 181794 507134 182414 507218
rect 181794 506898 181826 507134
rect 182062 506898 182146 507134
rect 182382 506898 182414 507134
rect 181794 471454 182414 506898
rect 181794 471218 181826 471454
rect 182062 471218 182146 471454
rect 182382 471218 182414 471454
rect 181794 471134 182414 471218
rect 181794 470898 181826 471134
rect 182062 470898 182146 471134
rect 182382 470898 182414 471134
rect 181794 435454 182414 470898
rect 181794 435218 181826 435454
rect 182062 435218 182146 435454
rect 182382 435218 182414 435454
rect 181794 435134 182414 435218
rect 181794 434898 181826 435134
rect 182062 434898 182146 435134
rect 182382 434898 182414 435134
rect 181794 399454 182414 434898
rect 181794 399218 181826 399454
rect 182062 399218 182146 399454
rect 182382 399218 182414 399454
rect 181794 399134 182414 399218
rect 181794 398898 181826 399134
rect 182062 398898 182146 399134
rect 182382 398898 182414 399134
rect 181794 363454 182414 398898
rect 181794 363218 181826 363454
rect 182062 363218 182146 363454
rect 182382 363218 182414 363454
rect 181794 363134 182414 363218
rect 181794 362898 181826 363134
rect 182062 362898 182146 363134
rect 182382 362898 182414 363134
rect 181794 327454 182414 362898
rect 181794 327218 181826 327454
rect 182062 327218 182146 327454
rect 182382 327218 182414 327454
rect 181794 327134 182414 327218
rect 181794 326898 181826 327134
rect 182062 326898 182146 327134
rect 182382 326898 182414 327134
rect 181794 291454 182414 326898
rect 181794 291218 181826 291454
rect 182062 291218 182146 291454
rect 182382 291218 182414 291454
rect 181794 291134 182414 291218
rect 181794 290898 181826 291134
rect 182062 290898 182146 291134
rect 182382 290898 182414 291134
rect 181794 262000 182414 290898
rect 186294 705798 186914 711590
rect 186294 705562 186326 705798
rect 186562 705562 186646 705798
rect 186882 705562 186914 705798
rect 186294 705478 186914 705562
rect 186294 705242 186326 705478
rect 186562 705242 186646 705478
rect 186882 705242 186914 705478
rect 186294 691954 186914 705242
rect 186294 691718 186326 691954
rect 186562 691718 186646 691954
rect 186882 691718 186914 691954
rect 186294 691634 186914 691718
rect 186294 691398 186326 691634
rect 186562 691398 186646 691634
rect 186882 691398 186914 691634
rect 186294 655954 186914 691398
rect 186294 655718 186326 655954
rect 186562 655718 186646 655954
rect 186882 655718 186914 655954
rect 186294 655634 186914 655718
rect 186294 655398 186326 655634
rect 186562 655398 186646 655634
rect 186882 655398 186914 655634
rect 186294 619954 186914 655398
rect 186294 619718 186326 619954
rect 186562 619718 186646 619954
rect 186882 619718 186914 619954
rect 186294 619634 186914 619718
rect 186294 619398 186326 619634
rect 186562 619398 186646 619634
rect 186882 619398 186914 619634
rect 186294 583954 186914 619398
rect 186294 583718 186326 583954
rect 186562 583718 186646 583954
rect 186882 583718 186914 583954
rect 186294 583634 186914 583718
rect 186294 583398 186326 583634
rect 186562 583398 186646 583634
rect 186882 583398 186914 583634
rect 186294 547954 186914 583398
rect 186294 547718 186326 547954
rect 186562 547718 186646 547954
rect 186882 547718 186914 547954
rect 186294 547634 186914 547718
rect 186294 547398 186326 547634
rect 186562 547398 186646 547634
rect 186882 547398 186914 547634
rect 186294 511954 186914 547398
rect 186294 511718 186326 511954
rect 186562 511718 186646 511954
rect 186882 511718 186914 511954
rect 186294 511634 186914 511718
rect 186294 511398 186326 511634
rect 186562 511398 186646 511634
rect 186882 511398 186914 511634
rect 186294 475954 186914 511398
rect 186294 475718 186326 475954
rect 186562 475718 186646 475954
rect 186882 475718 186914 475954
rect 186294 475634 186914 475718
rect 186294 475398 186326 475634
rect 186562 475398 186646 475634
rect 186882 475398 186914 475634
rect 186294 439954 186914 475398
rect 186294 439718 186326 439954
rect 186562 439718 186646 439954
rect 186882 439718 186914 439954
rect 186294 439634 186914 439718
rect 186294 439398 186326 439634
rect 186562 439398 186646 439634
rect 186882 439398 186914 439634
rect 186294 403954 186914 439398
rect 186294 403718 186326 403954
rect 186562 403718 186646 403954
rect 186882 403718 186914 403954
rect 186294 403634 186914 403718
rect 186294 403398 186326 403634
rect 186562 403398 186646 403634
rect 186882 403398 186914 403634
rect 186294 367954 186914 403398
rect 186294 367718 186326 367954
rect 186562 367718 186646 367954
rect 186882 367718 186914 367954
rect 186294 367634 186914 367718
rect 186294 367398 186326 367634
rect 186562 367398 186646 367634
rect 186882 367398 186914 367634
rect 186294 331954 186914 367398
rect 186294 331718 186326 331954
rect 186562 331718 186646 331954
rect 186882 331718 186914 331954
rect 186294 331634 186914 331718
rect 186294 331398 186326 331634
rect 186562 331398 186646 331634
rect 186882 331398 186914 331634
rect 186294 295954 186914 331398
rect 186294 295718 186326 295954
rect 186562 295718 186646 295954
rect 186882 295718 186914 295954
rect 186294 295634 186914 295718
rect 186294 295398 186326 295634
rect 186562 295398 186646 295634
rect 186882 295398 186914 295634
rect 186294 262000 186914 295398
rect 190794 706758 191414 711590
rect 190794 706522 190826 706758
rect 191062 706522 191146 706758
rect 191382 706522 191414 706758
rect 190794 706438 191414 706522
rect 190794 706202 190826 706438
rect 191062 706202 191146 706438
rect 191382 706202 191414 706438
rect 190794 696454 191414 706202
rect 190794 696218 190826 696454
rect 191062 696218 191146 696454
rect 191382 696218 191414 696454
rect 190794 696134 191414 696218
rect 190794 695898 190826 696134
rect 191062 695898 191146 696134
rect 191382 695898 191414 696134
rect 190794 660454 191414 695898
rect 190794 660218 190826 660454
rect 191062 660218 191146 660454
rect 191382 660218 191414 660454
rect 190794 660134 191414 660218
rect 190794 659898 190826 660134
rect 191062 659898 191146 660134
rect 191382 659898 191414 660134
rect 190794 624454 191414 659898
rect 190794 624218 190826 624454
rect 191062 624218 191146 624454
rect 191382 624218 191414 624454
rect 190794 624134 191414 624218
rect 190794 623898 190826 624134
rect 191062 623898 191146 624134
rect 191382 623898 191414 624134
rect 190794 588454 191414 623898
rect 190794 588218 190826 588454
rect 191062 588218 191146 588454
rect 191382 588218 191414 588454
rect 190794 588134 191414 588218
rect 190794 587898 190826 588134
rect 191062 587898 191146 588134
rect 191382 587898 191414 588134
rect 190794 552454 191414 587898
rect 190794 552218 190826 552454
rect 191062 552218 191146 552454
rect 191382 552218 191414 552454
rect 190794 552134 191414 552218
rect 190794 551898 190826 552134
rect 191062 551898 191146 552134
rect 191382 551898 191414 552134
rect 190794 516454 191414 551898
rect 190794 516218 190826 516454
rect 191062 516218 191146 516454
rect 191382 516218 191414 516454
rect 190794 516134 191414 516218
rect 190794 515898 190826 516134
rect 191062 515898 191146 516134
rect 191382 515898 191414 516134
rect 190794 480454 191414 515898
rect 190794 480218 190826 480454
rect 191062 480218 191146 480454
rect 191382 480218 191414 480454
rect 190794 480134 191414 480218
rect 190794 479898 190826 480134
rect 191062 479898 191146 480134
rect 191382 479898 191414 480134
rect 190794 444454 191414 479898
rect 190794 444218 190826 444454
rect 191062 444218 191146 444454
rect 191382 444218 191414 444454
rect 190794 444134 191414 444218
rect 190794 443898 190826 444134
rect 191062 443898 191146 444134
rect 191382 443898 191414 444134
rect 190794 408454 191414 443898
rect 190794 408218 190826 408454
rect 191062 408218 191146 408454
rect 191382 408218 191414 408454
rect 190794 408134 191414 408218
rect 190794 407898 190826 408134
rect 191062 407898 191146 408134
rect 191382 407898 191414 408134
rect 190794 372454 191414 407898
rect 190794 372218 190826 372454
rect 191062 372218 191146 372454
rect 191382 372218 191414 372454
rect 190794 372134 191414 372218
rect 190794 371898 190826 372134
rect 191062 371898 191146 372134
rect 191382 371898 191414 372134
rect 190794 336454 191414 371898
rect 190794 336218 190826 336454
rect 191062 336218 191146 336454
rect 191382 336218 191414 336454
rect 190794 336134 191414 336218
rect 190794 335898 190826 336134
rect 191062 335898 191146 336134
rect 191382 335898 191414 336134
rect 190794 300454 191414 335898
rect 190794 300218 190826 300454
rect 191062 300218 191146 300454
rect 191382 300218 191414 300454
rect 190794 300134 191414 300218
rect 190794 299898 190826 300134
rect 191062 299898 191146 300134
rect 191382 299898 191414 300134
rect 190794 264454 191414 299898
rect 190794 264218 190826 264454
rect 191062 264218 191146 264454
rect 191382 264218 191414 264454
rect 190794 264134 191414 264218
rect 190794 263898 190826 264134
rect 191062 263898 191146 264134
rect 191382 263898 191414 264134
rect 190794 262000 191414 263898
rect 195294 707718 195914 711590
rect 195294 707482 195326 707718
rect 195562 707482 195646 707718
rect 195882 707482 195914 707718
rect 195294 707398 195914 707482
rect 195294 707162 195326 707398
rect 195562 707162 195646 707398
rect 195882 707162 195914 707398
rect 195294 700954 195914 707162
rect 195294 700718 195326 700954
rect 195562 700718 195646 700954
rect 195882 700718 195914 700954
rect 195294 700634 195914 700718
rect 195294 700398 195326 700634
rect 195562 700398 195646 700634
rect 195882 700398 195914 700634
rect 195294 664954 195914 700398
rect 195294 664718 195326 664954
rect 195562 664718 195646 664954
rect 195882 664718 195914 664954
rect 195294 664634 195914 664718
rect 195294 664398 195326 664634
rect 195562 664398 195646 664634
rect 195882 664398 195914 664634
rect 195294 628954 195914 664398
rect 195294 628718 195326 628954
rect 195562 628718 195646 628954
rect 195882 628718 195914 628954
rect 195294 628634 195914 628718
rect 195294 628398 195326 628634
rect 195562 628398 195646 628634
rect 195882 628398 195914 628634
rect 195294 592954 195914 628398
rect 195294 592718 195326 592954
rect 195562 592718 195646 592954
rect 195882 592718 195914 592954
rect 195294 592634 195914 592718
rect 195294 592398 195326 592634
rect 195562 592398 195646 592634
rect 195882 592398 195914 592634
rect 195294 556954 195914 592398
rect 195294 556718 195326 556954
rect 195562 556718 195646 556954
rect 195882 556718 195914 556954
rect 195294 556634 195914 556718
rect 195294 556398 195326 556634
rect 195562 556398 195646 556634
rect 195882 556398 195914 556634
rect 195294 520954 195914 556398
rect 195294 520718 195326 520954
rect 195562 520718 195646 520954
rect 195882 520718 195914 520954
rect 195294 520634 195914 520718
rect 195294 520398 195326 520634
rect 195562 520398 195646 520634
rect 195882 520398 195914 520634
rect 195294 484954 195914 520398
rect 195294 484718 195326 484954
rect 195562 484718 195646 484954
rect 195882 484718 195914 484954
rect 195294 484634 195914 484718
rect 195294 484398 195326 484634
rect 195562 484398 195646 484634
rect 195882 484398 195914 484634
rect 195294 448954 195914 484398
rect 195294 448718 195326 448954
rect 195562 448718 195646 448954
rect 195882 448718 195914 448954
rect 195294 448634 195914 448718
rect 195294 448398 195326 448634
rect 195562 448398 195646 448634
rect 195882 448398 195914 448634
rect 195294 412954 195914 448398
rect 195294 412718 195326 412954
rect 195562 412718 195646 412954
rect 195882 412718 195914 412954
rect 195294 412634 195914 412718
rect 195294 412398 195326 412634
rect 195562 412398 195646 412634
rect 195882 412398 195914 412634
rect 195294 376954 195914 412398
rect 195294 376718 195326 376954
rect 195562 376718 195646 376954
rect 195882 376718 195914 376954
rect 195294 376634 195914 376718
rect 195294 376398 195326 376634
rect 195562 376398 195646 376634
rect 195882 376398 195914 376634
rect 195294 340954 195914 376398
rect 195294 340718 195326 340954
rect 195562 340718 195646 340954
rect 195882 340718 195914 340954
rect 195294 340634 195914 340718
rect 195294 340398 195326 340634
rect 195562 340398 195646 340634
rect 195882 340398 195914 340634
rect 195294 304954 195914 340398
rect 195294 304718 195326 304954
rect 195562 304718 195646 304954
rect 195882 304718 195914 304954
rect 195294 304634 195914 304718
rect 195294 304398 195326 304634
rect 195562 304398 195646 304634
rect 195882 304398 195914 304634
rect 195294 268954 195914 304398
rect 195294 268718 195326 268954
rect 195562 268718 195646 268954
rect 195882 268718 195914 268954
rect 195294 268634 195914 268718
rect 195294 268398 195326 268634
rect 195562 268398 195646 268634
rect 195882 268398 195914 268634
rect 191971 263804 192037 263805
rect 191971 263740 191972 263804
rect 192036 263740 192037 263804
rect 191971 263739 192037 263740
rect 191787 263668 191853 263669
rect 191787 263604 191788 263668
rect 191852 263604 191853 263668
rect 191787 263603 191853 263604
rect 187003 259996 187069 259997
rect 187003 259932 187004 259996
rect 187068 259932 187069 259996
rect 187003 259931 187069 259932
rect 122603 259588 122669 259589
rect 122603 259524 122604 259588
rect 122668 259524 122669 259588
rect 122603 259523 122669 259524
rect 122051 227764 122117 227765
rect 122051 227700 122052 227764
rect 122116 227700 122117 227764
rect 122051 227699 122117 227700
rect 121867 207092 121933 207093
rect 121867 207028 121868 207092
rect 121932 207028 121933 207092
rect 121867 207027 121933 207028
rect 121499 200836 121565 200837
rect 121499 200772 121500 200836
rect 121564 200772 121565 200836
rect 121499 200771 121565 200772
rect 121502 200157 121562 200771
rect 121499 200156 121565 200157
rect 121499 200092 121500 200156
rect 121564 200092 121565 200156
rect 121499 200091 121565 200092
rect 121870 199477 121930 207027
rect 122054 200973 122114 227699
rect 122235 211172 122301 211173
rect 122235 211108 122236 211172
rect 122300 211108 122301 211172
rect 122235 211107 122301 211108
rect 122051 200972 122117 200973
rect 122051 200908 122052 200972
rect 122116 200908 122117 200972
rect 122051 200907 122117 200908
rect 122238 199613 122298 211107
rect 122419 200156 122485 200157
rect 122419 200092 122420 200156
rect 122484 200092 122485 200156
rect 122419 200091 122485 200092
rect 122235 199612 122301 199613
rect 122235 199548 122236 199612
rect 122300 199548 122301 199612
rect 122235 199547 122301 199548
rect 121867 199476 121933 199477
rect 121867 199412 121868 199476
rect 121932 199412 121933 199476
rect 121867 199411 121933 199412
rect 122051 198388 122117 198389
rect 122051 198324 122052 198388
rect 122116 198324 122117 198388
rect 122051 198323 122117 198324
rect 118794 192454 119414 198000
rect 121315 194172 121381 194173
rect 121315 194108 121316 194172
rect 121380 194108 121381 194172
rect 121315 194107 121381 194108
rect 121131 194036 121197 194037
rect 121131 193972 121132 194036
rect 121196 193972 121197 194036
rect 121131 193971 121197 193972
rect 120579 192676 120645 192677
rect 120579 192612 120580 192676
rect 120644 192612 120645 192676
rect 120579 192611 120645 192612
rect 118794 192218 118826 192454
rect 119062 192218 119146 192454
rect 119382 192218 119414 192454
rect 118794 192134 119414 192218
rect 118794 191898 118826 192134
rect 119062 191898 119146 192134
rect 119382 191898 119414 192134
rect 118794 156454 119414 191898
rect 119843 184516 119909 184517
rect 119843 184452 119844 184516
rect 119908 184452 119909 184516
rect 119843 184451 119909 184452
rect 118794 156218 118826 156454
rect 119062 156218 119146 156454
rect 119382 156218 119414 156454
rect 118794 156134 119414 156218
rect 118794 155898 118826 156134
rect 119062 155898 119146 156134
rect 119382 155898 119414 156134
rect 118555 143172 118621 143173
rect 118555 143108 118556 143172
rect 118620 143108 118621 143172
rect 118555 143107 118621 143108
rect 118794 142000 119414 155898
rect 118555 141812 118621 141813
rect 118555 141748 118556 141812
rect 118620 141748 118621 141812
rect 118555 141747 118621 141748
rect 118371 141540 118437 141541
rect 118371 141476 118372 141540
rect 118436 141476 118437 141540
rect 118371 141475 118437 141476
rect 118187 140044 118253 140045
rect 118187 139980 118188 140044
rect 118252 139980 118253 140044
rect 118187 139979 118253 139980
rect 118190 75037 118250 139979
rect 118187 75036 118253 75037
rect 118187 74972 118188 75036
rect 118252 74972 118253 75036
rect 118187 74971 118253 74972
rect 117083 73812 117149 73813
rect 117083 73748 117084 73812
rect 117148 73748 117149 73812
rect 117083 73747 117149 73748
rect 118374 73677 118434 141475
rect 118371 73676 118437 73677
rect 118371 73612 118372 73676
rect 118436 73612 118437 73676
rect 118371 73611 118437 73612
rect 118558 73133 118618 141747
rect 119291 141404 119357 141405
rect 119291 141340 119292 141404
rect 119356 141340 119357 141404
rect 119291 141339 119357 141340
rect 119294 81157 119354 141339
rect 119475 140316 119541 140317
rect 119475 140252 119476 140316
rect 119540 140252 119541 140316
rect 119475 140251 119541 140252
rect 119291 81156 119357 81157
rect 119291 81092 119292 81156
rect 119356 81092 119357 81156
rect 119291 81091 119357 81092
rect 119478 78573 119538 140251
rect 119659 140180 119725 140181
rect 119659 140116 119660 140180
rect 119724 140116 119725 140180
rect 119659 140115 119725 140116
rect 119475 78572 119541 78573
rect 119475 78508 119476 78572
rect 119540 78508 119541 78572
rect 119475 78507 119541 78508
rect 118555 73132 118621 73133
rect 118555 73068 118556 73132
rect 118620 73068 118621 73132
rect 118555 73067 118621 73068
rect 115795 72724 115861 72725
rect 115795 72660 115796 72724
rect 115860 72660 115861 72724
rect 115795 72659 115861 72660
rect 114294 43718 114326 43954
rect 114562 43718 114646 43954
rect 114882 43718 114914 43954
rect 114294 43634 114914 43718
rect 114294 43398 114326 43634
rect 114562 43398 114646 43634
rect 114882 43398 114914 43634
rect 114294 7954 114914 43398
rect 114294 7718 114326 7954
rect 114562 7718 114646 7954
rect 114882 7718 114914 7954
rect 114294 7634 114914 7718
rect 114294 7398 114326 7634
rect 114562 7398 114646 7634
rect 114882 7398 114914 7634
rect 114294 -1306 114914 7398
rect 114294 -1542 114326 -1306
rect 114562 -1542 114646 -1306
rect 114882 -1542 114914 -1306
rect 114294 -1626 114914 -1542
rect 114294 -1862 114326 -1626
rect 114562 -1862 114646 -1626
rect 114882 -1862 114914 -1626
rect 114294 -7654 114914 -1862
rect 118794 48454 119414 78000
rect 119662 74221 119722 140115
rect 119659 74220 119725 74221
rect 119659 74156 119660 74220
rect 119724 74156 119725 74220
rect 119659 74155 119725 74156
rect 119846 66197 119906 184451
rect 120582 95165 120642 192611
rect 121134 177989 121194 193971
rect 121131 177988 121197 177989
rect 121131 177924 121132 177988
rect 121196 177924 121197 177988
rect 121131 177923 121197 177924
rect 120947 139228 121013 139229
rect 120947 139164 120948 139228
rect 121012 139164 121013 139228
rect 120947 139163 121013 139164
rect 120579 95164 120645 95165
rect 120579 95100 120580 95164
rect 120644 95100 120645 95164
rect 120579 95099 120645 95100
rect 120950 80613 121010 139163
rect 120947 80612 121013 80613
rect 120947 80548 120948 80612
rect 121012 80548 121013 80612
rect 120947 80547 121013 80548
rect 121134 78573 121194 177923
rect 121131 78572 121197 78573
rect 121131 78508 121132 78572
rect 121196 78508 121197 78572
rect 121131 78507 121197 78508
rect 121318 77485 121378 194107
rect 122054 174861 122114 198323
rect 122235 188460 122301 188461
rect 122235 188396 122236 188460
rect 122300 188396 122301 188460
rect 122235 188395 122301 188396
rect 122051 174860 122117 174861
rect 122051 174796 122052 174860
rect 122116 174796 122117 174860
rect 122051 174795 122117 174796
rect 122054 81429 122114 174795
rect 122051 81428 122117 81429
rect 122051 81364 122052 81428
rect 122116 81364 122117 81428
rect 122051 81363 122117 81364
rect 121315 77484 121381 77485
rect 121315 77420 121316 77484
rect 121380 77420 121381 77484
rect 121315 77419 121381 77420
rect 122238 70141 122298 188395
rect 122422 78981 122482 200091
rect 122606 195941 122666 259523
rect 124208 255454 124528 255486
rect 124208 255218 124250 255454
rect 124486 255218 124528 255454
rect 124208 255134 124528 255218
rect 124208 254898 124250 255134
rect 124486 254898 124528 255134
rect 124208 254866 124528 254898
rect 154928 255454 155248 255486
rect 154928 255218 154970 255454
rect 155206 255218 155248 255454
rect 154928 255134 155248 255218
rect 154928 254898 154970 255134
rect 155206 254898 155248 255134
rect 154928 254866 155248 254898
rect 185648 255454 185968 255486
rect 185648 255218 185690 255454
rect 185926 255218 185968 255454
rect 185648 255134 185968 255218
rect 185648 254898 185690 255134
rect 185926 254898 185968 255134
rect 185648 254866 185968 254898
rect 139568 223954 139888 223986
rect 139568 223718 139610 223954
rect 139846 223718 139888 223954
rect 139568 223634 139888 223718
rect 139568 223398 139610 223634
rect 139846 223398 139888 223634
rect 139568 223366 139888 223398
rect 170288 223954 170608 223986
rect 170288 223718 170330 223954
rect 170566 223718 170608 223954
rect 170288 223634 170608 223718
rect 170288 223398 170330 223634
rect 170566 223398 170608 223634
rect 170288 223366 170608 223398
rect 186819 220964 186885 220965
rect 186819 220900 186820 220964
rect 186884 220900 186885 220964
rect 186819 220899 186885 220900
rect 124208 219454 124528 219486
rect 124208 219218 124250 219454
rect 124486 219218 124528 219454
rect 124208 219134 124528 219218
rect 124208 218898 124250 219134
rect 124486 218898 124528 219134
rect 124208 218866 124528 218898
rect 154928 219454 155248 219486
rect 154928 219218 154970 219454
rect 155206 219218 155248 219454
rect 154928 219134 155248 219218
rect 154928 218898 154970 219134
rect 155206 218898 155248 219134
rect 154928 218866 155248 218898
rect 185648 219454 185968 219486
rect 185648 219218 185690 219454
rect 185926 219218 185968 219454
rect 185648 219134 185968 219218
rect 185648 218898 185690 219134
rect 185926 218898 185968 219134
rect 185648 218866 185968 218898
rect 186267 208452 186333 208453
rect 186267 208388 186268 208452
rect 186332 208388 186333 208452
rect 186267 208387 186333 208388
rect 186270 205650 186330 208387
rect 186086 205590 186330 205650
rect 176331 201516 176397 201517
rect 176331 201452 176332 201516
rect 176396 201452 176397 201516
rect 176331 201451 176397 201452
rect 156827 200836 156893 200837
rect 156827 200772 156828 200836
rect 156892 200772 156893 200836
rect 156827 200771 156893 200772
rect 168235 200836 168301 200837
rect 168235 200772 168236 200836
rect 168300 200772 168301 200836
rect 168235 200771 168301 200772
rect 138611 200700 138677 200701
rect 138062 200638 138490 200698
rect 138062 200021 138122 200638
rect 138243 200564 138309 200565
rect 138243 200500 138244 200564
rect 138308 200500 138309 200564
rect 138243 200499 138309 200500
rect 138059 200020 138125 200021
rect 138059 199956 138060 200020
rect 138124 199956 138125 200020
rect 138059 199955 138125 199956
rect 133091 199884 133157 199885
rect 133091 199820 133092 199884
rect 133156 199820 133157 199884
rect 133091 199819 133157 199820
rect 133275 199884 133341 199885
rect 133275 199820 133276 199884
rect 133340 199820 133341 199884
rect 133275 199819 133341 199820
rect 133827 199884 133893 199885
rect 133827 199820 133828 199884
rect 133892 199820 133893 199884
rect 133827 199819 133893 199820
rect 134379 199884 134445 199885
rect 134379 199820 134380 199884
rect 134444 199820 134445 199884
rect 134379 199819 134445 199820
rect 136035 199884 136101 199885
rect 136035 199820 136036 199884
rect 136100 199820 136101 199884
rect 136035 199819 136101 199820
rect 137323 199884 137389 199885
rect 137323 199820 137324 199884
rect 137388 199820 137389 199884
rect 137323 199819 137389 199820
rect 138059 199884 138125 199885
rect 138059 199820 138060 199884
rect 138124 199820 138125 199884
rect 138059 199819 138125 199820
rect 133094 199341 133154 199819
rect 133091 199340 133157 199341
rect 133091 199276 133092 199340
rect 133156 199276 133157 199340
rect 133091 199275 133157 199276
rect 133278 199205 133338 199819
rect 133830 199341 133890 199819
rect 133459 199340 133525 199341
rect 133459 199276 133460 199340
rect 133524 199276 133525 199340
rect 133459 199275 133525 199276
rect 133827 199340 133893 199341
rect 133827 199276 133828 199340
rect 133892 199276 133893 199340
rect 133827 199275 133893 199276
rect 133275 199204 133341 199205
rect 133275 199140 133276 199204
rect 133340 199140 133341 199204
rect 133275 199139 133341 199140
rect 124075 198524 124141 198525
rect 124075 198460 124076 198524
rect 124140 198460 124141 198524
rect 124075 198459 124141 198460
rect 123294 196954 123914 198000
rect 123294 196718 123326 196954
rect 123562 196718 123646 196954
rect 123882 196718 123914 196954
rect 123294 196634 123914 196718
rect 123294 196398 123326 196634
rect 123562 196398 123646 196634
rect 123882 196398 123914 196634
rect 122603 195940 122669 195941
rect 122603 195876 122604 195940
rect 122668 195876 122669 195940
rect 122603 195875 122669 195876
rect 122603 195532 122669 195533
rect 122603 195468 122604 195532
rect 122668 195468 122669 195532
rect 122603 195467 122669 195468
rect 122419 78980 122485 78981
rect 122419 78916 122420 78980
rect 122484 78916 122485 78980
rect 122419 78915 122485 78916
rect 122235 70140 122301 70141
rect 122235 70076 122236 70140
rect 122300 70076 122301 70140
rect 122235 70075 122301 70076
rect 122606 68917 122666 195467
rect 122787 190500 122853 190501
rect 122787 190436 122788 190500
rect 122852 190470 122853 190500
rect 122852 190436 123034 190470
rect 122787 190435 123034 190436
rect 122790 190410 123034 190435
rect 122974 189549 123034 190410
rect 122971 189548 123037 189549
rect 122971 189484 122972 189548
rect 123036 189484 123037 189548
rect 122971 189483 123037 189484
rect 122971 181524 123037 181525
rect 122971 181460 122972 181524
rect 123036 181460 123037 181524
rect 122971 181459 123037 181460
rect 122974 180810 123034 181459
rect 122790 180750 123034 180810
rect 122790 180573 122850 180750
rect 122787 180572 122853 180573
rect 122787 180508 122788 180572
rect 122852 180508 122853 180572
rect 122787 180507 122853 180508
rect 122787 171188 122853 171189
rect 122787 171124 122788 171188
rect 122852 171124 122853 171188
rect 122787 171123 122853 171124
rect 122790 171053 122850 171123
rect 122787 171052 122853 171053
rect 122787 170988 122788 171052
rect 122852 170988 122853 171052
rect 122787 170987 122853 170988
rect 122971 161532 123037 161533
rect 122971 161530 122972 161532
rect 122790 161470 122972 161530
rect 122790 161397 122850 161470
rect 122971 161468 122972 161470
rect 123036 161468 123037 161532
rect 122971 161467 123037 161468
rect 122787 161396 122853 161397
rect 122787 161332 122788 161396
rect 122852 161332 122853 161396
rect 122787 161331 122853 161332
rect 123294 160954 123914 196398
rect 123294 160718 123326 160954
rect 123562 160718 123646 160954
rect 123882 160718 123914 160954
rect 123294 160634 123914 160718
rect 123294 160398 123326 160634
rect 123562 160398 123646 160634
rect 123882 160398 123914 160634
rect 122787 152012 122853 152013
rect 122787 151948 122788 152012
rect 122852 151948 122853 152012
rect 122787 151947 122853 151948
rect 122790 151605 122850 151947
rect 122787 151604 122853 151605
rect 122787 151540 122788 151604
rect 122852 151540 122853 151604
rect 122787 151539 122853 151540
rect 122787 147660 122853 147661
rect 122787 147596 122788 147660
rect 122852 147596 122853 147660
rect 122787 147595 122853 147596
rect 122790 138141 122850 147595
rect 123294 142000 123914 160398
rect 123339 139364 123405 139365
rect 123339 139300 123340 139364
rect 123404 139300 123405 139364
rect 123339 139299 123405 139300
rect 123891 139364 123957 139365
rect 123891 139300 123892 139364
rect 123956 139300 123957 139364
rect 123891 139299 123957 139300
rect 122787 138140 122853 138141
rect 122787 138076 122788 138140
rect 122852 138076 122853 138140
rect 122787 138075 122853 138076
rect 123342 136101 123402 139299
rect 123339 136100 123405 136101
rect 123339 136036 123340 136100
rect 123404 136036 123405 136100
rect 123339 136035 123405 136036
rect 123894 78165 123954 139299
rect 124078 80613 124138 198459
rect 133462 195941 133522 199275
rect 134382 199205 134442 199819
rect 134563 199340 134629 199341
rect 134563 199276 134564 199340
rect 134628 199276 134629 199340
rect 134563 199275 134629 199276
rect 135851 199340 135917 199341
rect 135851 199276 135852 199340
rect 135916 199276 135917 199340
rect 135851 199275 135917 199276
rect 134379 199204 134445 199205
rect 134379 199140 134380 199204
rect 134444 199140 134445 199204
rect 134379 199139 134445 199140
rect 133459 195940 133525 195941
rect 133459 195876 133460 195940
rect 133524 195876 133525 195940
rect 133459 195875 133525 195876
rect 134379 193900 134445 193901
rect 134379 193836 134380 193900
rect 134444 193836 134445 193900
rect 134379 193835 134445 193836
rect 134382 178941 134442 193835
rect 134566 190773 134626 199275
rect 134563 190772 134629 190773
rect 134563 190708 134564 190772
rect 134628 190708 134629 190772
rect 134563 190707 134629 190708
rect 134379 178940 134445 178941
rect 134379 178876 134380 178940
rect 134444 178876 134445 178940
rect 134379 178875 134445 178876
rect 135854 176629 135914 199275
rect 136038 198750 136098 199819
rect 137326 199341 137386 199819
rect 136403 199340 136469 199341
rect 136403 199276 136404 199340
rect 136468 199276 136469 199340
rect 136403 199275 136469 199276
rect 136955 199340 137021 199341
rect 136955 199276 136956 199340
rect 137020 199276 137021 199340
rect 136955 199275 137021 199276
rect 137323 199340 137389 199341
rect 137323 199276 137324 199340
rect 137388 199276 137389 199340
rect 137323 199275 137389 199276
rect 136038 198690 136282 198750
rect 136222 198525 136282 198690
rect 136219 198524 136285 198525
rect 136219 198460 136220 198524
rect 136284 198460 136285 198524
rect 136219 198459 136285 198460
rect 136406 195941 136466 199275
rect 136771 199204 136837 199205
rect 136771 199140 136772 199204
rect 136836 199140 136837 199204
rect 136771 199139 136837 199140
rect 136403 195940 136469 195941
rect 136403 195876 136404 195940
rect 136468 195876 136469 195940
rect 136403 195875 136469 195876
rect 136774 192813 136834 199139
rect 136958 198525 137018 199275
rect 138062 199205 138122 199819
rect 138246 199341 138306 200499
rect 138243 199340 138309 199341
rect 138243 199276 138244 199340
rect 138308 199276 138309 199340
rect 138243 199275 138309 199276
rect 138059 199204 138125 199205
rect 138059 199140 138060 199204
rect 138124 199140 138125 199204
rect 138059 199139 138125 199140
rect 136955 198524 137021 198525
rect 136955 198460 136956 198524
rect 137020 198460 137021 198524
rect 136955 198459 137021 198460
rect 138430 196349 138490 200638
rect 138611 200636 138612 200700
rect 138676 200636 138677 200700
rect 138611 200635 138677 200636
rect 152411 200700 152477 200701
rect 152411 200636 152412 200700
rect 152476 200636 152477 200700
rect 152411 200635 152477 200636
rect 138614 198797 138674 200635
rect 145603 200428 145669 200429
rect 145603 200364 145604 200428
rect 145668 200364 145669 200428
rect 145603 200363 145669 200364
rect 139347 200292 139413 200293
rect 139347 200228 139348 200292
rect 139412 200228 139413 200292
rect 139347 200227 139413 200228
rect 138979 199884 139045 199885
rect 138979 199820 138980 199884
rect 139044 199820 139045 199884
rect 138979 199819 139045 199820
rect 139163 199884 139229 199885
rect 139163 199820 139164 199884
rect 139228 199820 139229 199884
rect 139163 199819 139229 199820
rect 138611 198796 138677 198797
rect 138611 198732 138612 198796
rect 138676 198732 138677 198796
rect 138611 198731 138677 198732
rect 138795 198660 138861 198661
rect 138795 198596 138796 198660
rect 138860 198596 138861 198660
rect 138795 198595 138861 198596
rect 138611 198524 138677 198525
rect 138611 198460 138612 198524
rect 138676 198460 138677 198524
rect 138611 198459 138677 198460
rect 138614 198117 138674 198459
rect 138611 198116 138677 198117
rect 138611 198052 138612 198116
rect 138676 198052 138677 198116
rect 138611 198051 138677 198052
rect 138611 197844 138677 197845
rect 138611 197780 138612 197844
rect 138676 197780 138677 197844
rect 138611 197779 138677 197780
rect 138427 196348 138493 196349
rect 138427 196284 138428 196348
rect 138492 196284 138493 196348
rect 138427 196283 138493 196284
rect 137323 196076 137389 196077
rect 137323 196012 137324 196076
rect 137388 196012 137389 196076
rect 137323 196011 137389 196012
rect 136771 192812 136837 192813
rect 136771 192748 136772 192812
rect 136836 192748 136837 192812
rect 136771 192747 136837 192748
rect 135851 176628 135917 176629
rect 135851 176564 135852 176628
rect 135916 176564 135917 176628
rect 135851 176563 135917 176564
rect 137326 175133 137386 196011
rect 138614 177309 138674 197779
rect 138798 191850 138858 198595
rect 138982 198117 139042 199819
rect 139166 198253 139226 199819
rect 139350 199205 139410 200227
rect 145606 199885 145666 200363
rect 147995 200156 148061 200157
rect 147995 200092 147996 200156
rect 148060 200092 148061 200156
rect 147995 200091 148061 200092
rect 149467 200156 149533 200157
rect 149467 200092 149468 200156
rect 149532 200092 149533 200156
rect 149467 200091 149533 200092
rect 139531 199884 139597 199885
rect 139531 199820 139532 199884
rect 139596 199820 139597 199884
rect 139531 199819 139597 199820
rect 139899 199884 139965 199885
rect 139899 199820 139900 199884
rect 139964 199820 139965 199884
rect 139899 199819 139965 199820
rect 140267 199884 140333 199885
rect 140267 199820 140268 199884
rect 140332 199820 140333 199884
rect 140267 199819 140333 199820
rect 140635 199884 140701 199885
rect 140635 199820 140636 199884
rect 140700 199820 140701 199884
rect 140635 199819 140701 199820
rect 141187 199884 141253 199885
rect 141187 199820 141188 199884
rect 141252 199820 141253 199884
rect 141187 199819 141253 199820
rect 142475 199884 142541 199885
rect 142475 199820 142476 199884
rect 142540 199820 142541 199884
rect 142475 199819 142541 199820
rect 143027 199884 143093 199885
rect 143027 199820 143028 199884
rect 143092 199820 143093 199884
rect 143027 199819 143093 199820
rect 144315 199884 144381 199885
rect 144315 199820 144316 199884
rect 144380 199820 144381 199884
rect 144315 199819 144381 199820
rect 144867 199884 144933 199885
rect 144867 199820 144868 199884
rect 144932 199820 144933 199884
rect 144867 199819 144933 199820
rect 145419 199884 145485 199885
rect 145419 199820 145420 199884
rect 145484 199820 145485 199884
rect 145419 199819 145485 199820
rect 145603 199884 145669 199885
rect 145603 199820 145604 199884
rect 145668 199820 145669 199884
rect 145603 199819 145669 199820
rect 146155 199884 146221 199885
rect 146155 199820 146156 199884
rect 146220 199820 146221 199884
rect 146155 199819 146221 199820
rect 146523 199884 146589 199885
rect 146523 199820 146524 199884
rect 146588 199820 146589 199884
rect 146523 199819 146589 199820
rect 147811 199884 147877 199885
rect 147811 199820 147812 199884
rect 147876 199820 147877 199884
rect 147811 199819 147877 199820
rect 139347 199204 139413 199205
rect 139347 199140 139348 199204
rect 139412 199140 139413 199204
rect 139347 199139 139413 199140
rect 139163 198252 139229 198253
rect 139163 198188 139164 198252
rect 139228 198188 139229 198252
rect 139163 198187 139229 198188
rect 138979 198116 139045 198117
rect 138979 198052 138980 198116
rect 139044 198052 139045 198116
rect 138979 198051 139045 198052
rect 139534 197709 139594 199819
rect 139902 198253 139962 199819
rect 139899 198252 139965 198253
rect 139899 198188 139900 198252
rect 139964 198188 139965 198252
rect 139899 198187 139965 198188
rect 139899 198116 139965 198117
rect 139899 198052 139900 198116
rect 139964 198052 139965 198116
rect 139899 198051 139965 198052
rect 139531 197708 139597 197709
rect 139531 197644 139532 197708
rect 139596 197644 139597 197708
rect 139531 197643 139597 197644
rect 139163 195940 139229 195941
rect 139163 195876 139164 195940
rect 139228 195876 139229 195940
rect 139163 195875 139229 195876
rect 138798 191790 139042 191850
rect 138982 189005 139042 191790
rect 138979 189004 139045 189005
rect 138979 188940 138980 189004
rect 139044 188940 139045 189004
rect 138979 188939 139045 188940
rect 139166 184925 139226 195875
rect 139902 190229 139962 198051
rect 140270 197437 140330 199819
rect 140638 197573 140698 199819
rect 141190 199205 141250 199819
rect 141187 199204 141253 199205
rect 141187 199140 141188 199204
rect 141252 199140 141253 199204
rect 141187 199139 141253 199140
rect 140819 198796 140885 198797
rect 140819 198732 140820 198796
rect 140884 198732 140885 198796
rect 140819 198731 140885 198732
rect 140635 197572 140701 197573
rect 140635 197508 140636 197572
rect 140700 197508 140701 197572
rect 140635 197507 140701 197508
rect 140267 197436 140333 197437
rect 140267 197372 140268 197436
rect 140332 197372 140333 197436
rect 140267 197371 140333 197372
rect 140635 195668 140701 195669
rect 140635 195604 140636 195668
rect 140700 195604 140701 195668
rect 140635 195603 140701 195604
rect 139899 190228 139965 190229
rect 139899 190164 139900 190228
rect 139964 190164 139965 190228
rect 139899 190163 139965 190164
rect 139163 184924 139229 184925
rect 139163 184860 139164 184924
rect 139228 184860 139229 184924
rect 139163 184859 139229 184860
rect 140638 177853 140698 195603
rect 140635 177852 140701 177853
rect 140635 177788 140636 177852
rect 140700 177788 140701 177852
rect 140635 177787 140701 177788
rect 138611 177308 138677 177309
rect 138611 177244 138612 177308
rect 138676 177244 138677 177308
rect 138611 177243 138677 177244
rect 140822 176629 140882 198731
rect 141003 198660 141069 198661
rect 141003 198596 141004 198660
rect 141068 198596 141069 198660
rect 141003 198595 141069 198596
rect 140819 176628 140885 176629
rect 140819 176564 140820 176628
rect 140884 176564 140885 176628
rect 140819 176563 140885 176564
rect 141006 175269 141066 198595
rect 141294 178954 141914 198000
rect 142478 197165 142538 199819
rect 143030 198117 143090 199819
rect 143947 199204 144013 199205
rect 143947 199140 143948 199204
rect 144012 199140 144013 199204
rect 143947 199139 144013 199140
rect 143027 198116 143093 198117
rect 143027 198052 143028 198116
rect 143092 198052 143093 198116
rect 143027 198051 143093 198052
rect 142475 197164 142541 197165
rect 142475 197100 142476 197164
rect 142540 197100 142541 197164
rect 142475 197099 142541 197100
rect 142478 196621 142538 197099
rect 142475 196620 142541 196621
rect 142475 196556 142476 196620
rect 142540 196556 142541 196620
rect 142475 196555 142541 196556
rect 143950 193230 144010 199139
rect 144318 198797 144378 199819
rect 144315 198796 144381 198797
rect 144315 198732 144316 198796
rect 144380 198732 144381 198796
rect 144315 198731 144381 198732
rect 144315 198660 144381 198661
rect 144315 198596 144316 198660
rect 144380 198596 144381 198660
rect 144315 198595 144381 198596
rect 143582 193170 144010 193230
rect 143582 189957 143642 193170
rect 144318 191850 144378 198595
rect 144870 198117 144930 199819
rect 144867 198116 144933 198117
rect 144867 198052 144868 198116
rect 144932 198052 144933 198116
rect 144867 198051 144933 198052
rect 144134 191790 144378 191850
rect 143579 189956 143645 189957
rect 143579 189892 143580 189956
rect 143644 189892 143645 189956
rect 143579 189891 143645 189892
rect 141294 178718 141326 178954
rect 141562 178718 141646 178954
rect 141882 178718 141914 178954
rect 141294 178634 141914 178718
rect 141294 178398 141326 178634
rect 141562 178398 141646 178634
rect 141882 178398 141914 178634
rect 141003 175268 141069 175269
rect 141003 175204 141004 175268
rect 141068 175204 141069 175268
rect 141003 175203 141069 175204
rect 137323 175132 137389 175133
rect 137323 175068 137324 175132
rect 137388 175068 137389 175132
rect 137323 175067 137389 175068
rect 137326 174589 137386 175067
rect 137323 174588 137389 174589
rect 137323 174524 137324 174588
rect 137388 174524 137389 174588
rect 137323 174523 137389 174524
rect 141294 142954 141914 178398
rect 144134 148341 144194 191790
rect 145422 186285 145482 199819
rect 146158 198525 146218 199819
rect 146155 198524 146221 198525
rect 146155 198460 146156 198524
rect 146220 198460 146221 198524
rect 146155 198459 146221 198460
rect 145419 186284 145485 186285
rect 145419 186220 145420 186284
rect 145484 186220 145485 186284
rect 145419 186219 145485 186220
rect 145794 183454 146414 198000
rect 146526 197845 146586 199819
rect 146891 199204 146957 199205
rect 146891 199140 146892 199204
rect 146956 199140 146957 199204
rect 146891 199139 146957 199140
rect 147075 199204 147141 199205
rect 147075 199140 147076 199204
rect 147140 199140 147141 199204
rect 147075 199139 147141 199140
rect 146523 197844 146589 197845
rect 146523 197780 146524 197844
rect 146588 197780 146589 197844
rect 146523 197779 146589 197780
rect 146894 184381 146954 199139
rect 147078 192677 147138 199139
rect 147814 197437 147874 199819
rect 147811 197436 147877 197437
rect 147811 197372 147812 197436
rect 147876 197372 147877 197436
rect 147811 197371 147877 197372
rect 147811 196620 147877 196621
rect 147811 196556 147812 196620
rect 147876 196556 147877 196620
rect 147811 196555 147877 196556
rect 147075 192676 147141 192677
rect 147075 192612 147076 192676
rect 147140 192612 147141 192676
rect 147075 192611 147141 192612
rect 147814 186330 147874 196555
rect 147998 192541 148058 200091
rect 148363 199884 148429 199885
rect 148363 199820 148364 199884
rect 148428 199820 148429 199884
rect 148363 199819 148429 199820
rect 148547 199884 148613 199885
rect 148547 199820 148548 199884
rect 148612 199820 148613 199884
rect 148547 199819 148613 199820
rect 148915 199884 148981 199885
rect 148915 199820 148916 199884
rect 148980 199820 148981 199884
rect 148915 199819 148981 199820
rect 149283 199884 149349 199885
rect 149283 199820 149284 199884
rect 149348 199820 149349 199884
rect 149283 199819 149349 199820
rect 147995 192540 148061 192541
rect 147995 192476 147996 192540
rect 148060 192476 148061 192540
rect 147995 192475 148061 192476
rect 148366 190501 148426 199819
rect 148550 198117 148610 199819
rect 148547 198116 148613 198117
rect 148547 198052 148548 198116
rect 148612 198052 148613 198116
rect 148547 198051 148613 198052
rect 148918 192133 148978 199819
rect 149286 198933 149346 199819
rect 149470 199205 149530 200091
rect 152414 199885 152474 200635
rect 153331 200156 153397 200157
rect 153331 200092 153332 200156
rect 153396 200092 153397 200156
rect 153331 200091 153397 200092
rect 154435 200156 154501 200157
rect 154435 200092 154436 200156
rect 154500 200092 154501 200156
rect 154435 200091 154501 200092
rect 149651 199884 149717 199885
rect 149651 199820 149652 199884
rect 149716 199820 149717 199884
rect 149651 199819 149717 199820
rect 150203 199884 150269 199885
rect 150203 199820 150204 199884
rect 150268 199820 150269 199884
rect 150203 199819 150269 199820
rect 150571 199884 150637 199885
rect 150571 199820 150572 199884
rect 150636 199820 150637 199884
rect 150571 199819 150637 199820
rect 151491 199884 151557 199885
rect 151491 199820 151492 199884
rect 151556 199820 151557 199884
rect 151491 199819 151557 199820
rect 152043 199884 152109 199885
rect 152043 199820 152044 199884
rect 152108 199820 152109 199884
rect 152043 199819 152109 199820
rect 152411 199884 152477 199885
rect 152411 199820 152412 199884
rect 152476 199820 152477 199884
rect 152411 199819 152477 199820
rect 153147 199884 153213 199885
rect 153147 199820 153148 199884
rect 153212 199820 153213 199884
rect 153147 199819 153213 199820
rect 149467 199204 149533 199205
rect 149467 199140 149468 199204
rect 149532 199140 149533 199204
rect 149467 199139 149533 199140
rect 149283 198932 149349 198933
rect 149283 198868 149284 198932
rect 149348 198868 149349 198932
rect 149283 198867 149349 198868
rect 149654 197981 149714 199819
rect 150206 199069 150266 199819
rect 150203 199068 150269 199069
rect 150203 199004 150204 199068
rect 150268 199004 150269 199068
rect 150203 199003 150269 199004
rect 149835 198796 149901 198797
rect 149835 198732 149836 198796
rect 149900 198732 149901 198796
rect 149835 198731 149901 198732
rect 150019 198796 150085 198797
rect 150019 198732 150020 198796
rect 150084 198732 150085 198796
rect 150019 198731 150085 198732
rect 149651 197980 149717 197981
rect 149651 197916 149652 197980
rect 149716 197916 149717 197980
rect 149651 197915 149717 197916
rect 148915 192132 148981 192133
rect 148915 192068 148916 192132
rect 148980 192068 148981 192132
rect 148915 192067 148981 192068
rect 148363 190500 148429 190501
rect 148363 190436 148364 190500
rect 148428 190436 148429 190500
rect 148363 190435 148429 190436
rect 149838 188325 149898 198731
rect 149835 188324 149901 188325
rect 149835 188260 149836 188324
rect 149900 188260 149901 188324
rect 149835 188259 149901 188260
rect 147630 186270 147874 186330
rect 146891 184380 146957 184381
rect 146891 184316 146892 184380
rect 146956 184316 146957 184380
rect 146891 184315 146957 184316
rect 147630 184245 147690 186270
rect 147627 184244 147693 184245
rect 147627 184180 147628 184244
rect 147692 184180 147693 184244
rect 147627 184179 147693 184180
rect 145794 183218 145826 183454
rect 146062 183218 146146 183454
rect 146382 183218 146414 183454
rect 145794 183134 146414 183218
rect 145794 182898 145826 183134
rect 146062 182898 146146 183134
rect 146382 182898 146414 183134
rect 144131 148340 144197 148341
rect 144131 148276 144132 148340
rect 144196 148276 144197 148340
rect 144131 148275 144197 148276
rect 141294 142718 141326 142954
rect 141562 142718 141646 142954
rect 141882 142718 141914 142954
rect 141294 142634 141914 142718
rect 141294 142398 141326 142634
rect 141562 142398 141646 142634
rect 141882 142398 141914 142634
rect 141294 142000 141914 142398
rect 145794 147454 146414 182898
rect 150022 181389 150082 198731
rect 150574 198389 150634 199819
rect 151123 198796 151189 198797
rect 151123 198732 151124 198796
rect 151188 198732 151189 198796
rect 151123 198731 151189 198732
rect 150571 198388 150637 198389
rect 150571 198324 150572 198388
rect 150636 198324 150637 198388
rect 150571 198323 150637 198324
rect 150294 187954 150914 198000
rect 150294 187718 150326 187954
rect 150562 187718 150646 187954
rect 150882 187718 150914 187954
rect 150294 187634 150914 187718
rect 150294 187398 150326 187634
rect 150562 187398 150646 187634
rect 150882 187398 150914 187634
rect 150019 181388 150085 181389
rect 150019 181324 150020 181388
rect 150084 181324 150085 181388
rect 150019 181323 150085 181324
rect 145794 147218 145826 147454
rect 146062 147218 146146 147454
rect 146382 147218 146414 147454
rect 145794 147134 146414 147218
rect 145794 146898 145826 147134
rect 146062 146898 146146 147134
rect 146382 146898 146414 147134
rect 145794 142000 146414 146898
rect 150294 151954 150914 187398
rect 150294 151718 150326 151954
rect 150562 151718 150646 151954
rect 150882 151718 150914 151954
rect 150294 151634 150914 151718
rect 150294 151398 150326 151634
rect 150562 151398 150646 151634
rect 150882 151398 150914 151634
rect 150294 142000 150914 151398
rect 151126 140317 151186 198731
rect 151494 198389 151554 199819
rect 151675 199068 151741 199069
rect 151675 199004 151676 199068
rect 151740 199004 151741 199068
rect 151675 199003 151741 199004
rect 151491 198388 151557 198389
rect 151491 198324 151492 198388
rect 151556 198324 151557 198388
rect 151491 198323 151557 198324
rect 151678 181525 151738 199003
rect 152046 193230 152106 199819
rect 152414 198117 152474 199819
rect 153150 199341 153210 199819
rect 153147 199340 153213 199341
rect 153147 199276 153148 199340
rect 153212 199276 153213 199340
rect 153147 199275 153213 199276
rect 153334 198797 153394 200091
rect 153515 199884 153581 199885
rect 153515 199820 153516 199884
rect 153580 199820 153581 199884
rect 153515 199819 153581 199820
rect 154251 199884 154317 199885
rect 154251 199820 154252 199884
rect 154316 199820 154317 199884
rect 154251 199819 154317 199820
rect 153331 198796 153397 198797
rect 153331 198732 153332 198796
rect 153396 198732 153397 198796
rect 153331 198731 153397 198732
rect 152411 198116 152477 198117
rect 152411 198052 152412 198116
rect 152476 198052 152477 198116
rect 152411 198051 152477 198052
rect 152779 196484 152845 196485
rect 152779 196420 152780 196484
rect 152844 196420 152845 196484
rect 152779 196419 152845 196420
rect 151862 193170 152106 193230
rect 151862 191453 151922 193170
rect 151859 191452 151925 191453
rect 151859 191388 151860 191452
rect 151924 191388 151925 191452
rect 151859 191387 151925 191388
rect 152782 183293 152842 196419
rect 152963 196348 153029 196349
rect 152963 196284 152964 196348
rect 153028 196284 153029 196348
rect 152963 196283 153029 196284
rect 152779 183292 152845 183293
rect 152779 183228 152780 183292
rect 152844 183228 152845 183292
rect 152779 183227 152845 183228
rect 152966 181661 153026 196283
rect 153518 196077 153578 199819
rect 154254 198797 154314 199819
rect 154438 198797 154498 200091
rect 156830 199885 156890 200771
rect 160323 200292 160389 200293
rect 160323 200228 160324 200292
rect 160388 200228 160389 200292
rect 160323 200227 160389 200228
rect 161611 200292 161677 200293
rect 161611 200228 161612 200292
rect 161676 200228 161677 200292
rect 161611 200227 161677 200228
rect 154803 199884 154869 199885
rect 154803 199820 154804 199884
rect 154868 199820 154869 199884
rect 154803 199819 154869 199820
rect 156827 199884 156893 199885
rect 156827 199820 156828 199884
rect 156892 199820 156893 199884
rect 156827 199819 156893 199820
rect 158299 199884 158365 199885
rect 158299 199820 158300 199884
rect 158364 199820 158365 199884
rect 158299 199819 158365 199820
rect 158851 199884 158917 199885
rect 158851 199820 158852 199884
rect 158916 199820 158917 199884
rect 158851 199819 158917 199820
rect 159219 199884 159285 199885
rect 159219 199820 159220 199884
rect 159284 199820 159285 199884
rect 159219 199819 159285 199820
rect 154251 198796 154317 198797
rect 154251 198732 154252 198796
rect 154316 198732 154317 198796
rect 154251 198731 154317 198732
rect 154435 198796 154501 198797
rect 154435 198732 154436 198796
rect 154500 198732 154501 198796
rect 154435 198731 154501 198732
rect 154806 198389 154866 199819
rect 158302 199205 158362 199819
rect 158115 199204 158181 199205
rect 158115 199140 158116 199204
rect 158180 199140 158181 199204
rect 158115 199139 158181 199140
rect 158299 199204 158365 199205
rect 158299 199140 158300 199204
rect 158364 199140 158365 199204
rect 158299 199139 158365 199140
rect 154803 198388 154869 198389
rect 154803 198324 154804 198388
rect 154868 198324 154869 198388
rect 154803 198323 154869 198324
rect 154619 198116 154685 198117
rect 154619 198052 154620 198116
rect 154684 198052 154685 198116
rect 154619 198051 154685 198052
rect 154435 196212 154501 196213
rect 154435 196148 154436 196212
rect 154500 196148 154501 196212
rect 154435 196147 154501 196148
rect 153515 196076 153581 196077
rect 153515 196012 153516 196076
rect 153580 196012 153581 196076
rect 153515 196011 153581 196012
rect 154438 183021 154498 196147
rect 154622 190365 154682 198051
rect 154794 192454 155414 198000
rect 157195 196212 157261 196213
rect 157195 196148 157196 196212
rect 157260 196148 157261 196212
rect 157195 196147 157261 196148
rect 157011 196076 157077 196077
rect 157011 196012 157012 196076
rect 157076 196012 157077 196076
rect 157011 196011 157077 196012
rect 154794 192218 154826 192454
rect 155062 192218 155146 192454
rect 155382 192218 155414 192454
rect 154794 192134 155414 192218
rect 154794 191898 154826 192134
rect 155062 191898 155146 192134
rect 155382 191898 155414 192134
rect 154619 190364 154685 190365
rect 154619 190300 154620 190364
rect 154684 190300 154685 190364
rect 154619 190299 154685 190300
rect 154435 183020 154501 183021
rect 154435 182956 154436 183020
rect 154500 182956 154501 183020
rect 154435 182955 154501 182956
rect 152963 181660 153029 181661
rect 152963 181596 152964 181660
rect 153028 181596 153029 181660
rect 152963 181595 153029 181596
rect 151675 181524 151741 181525
rect 151675 181460 151676 181524
rect 151740 181460 151741 181524
rect 151675 181459 151741 181460
rect 154794 156454 155414 191898
rect 157014 189685 157074 196011
rect 157198 190365 157258 196147
rect 157195 190364 157261 190365
rect 157195 190300 157196 190364
rect 157260 190300 157261 190364
rect 157195 190299 157261 190300
rect 157011 189684 157077 189685
rect 157011 189620 157012 189684
rect 157076 189620 157077 189684
rect 157011 189619 157077 189620
rect 158118 183565 158178 199139
rect 158854 198797 158914 199819
rect 159222 198797 159282 199819
rect 158851 198796 158917 198797
rect 158851 198732 158852 198796
rect 158916 198732 158917 198796
rect 158851 198731 158917 198732
rect 159219 198796 159285 198797
rect 159219 198732 159220 198796
rect 159284 198732 159285 198796
rect 159219 198731 159285 198732
rect 159294 196954 159914 198000
rect 159294 196718 159326 196954
rect 159562 196718 159646 196954
rect 159882 196718 159914 196954
rect 159294 196634 159914 196718
rect 158299 196484 158365 196485
rect 158299 196420 158300 196484
rect 158364 196420 158365 196484
rect 158299 196419 158365 196420
rect 158302 190093 158362 196419
rect 159294 196398 159326 196634
rect 159562 196398 159646 196634
rect 159882 196398 159914 196634
rect 158667 196076 158733 196077
rect 158667 196012 158668 196076
rect 158732 196012 158733 196076
rect 158667 196011 158733 196012
rect 158670 191181 158730 196011
rect 158667 191180 158733 191181
rect 158667 191116 158668 191180
rect 158732 191116 158733 191180
rect 158667 191115 158733 191116
rect 158299 190092 158365 190093
rect 158299 190028 158300 190092
rect 158364 190028 158365 190092
rect 158299 190027 158365 190028
rect 158115 183564 158181 183565
rect 158115 183500 158116 183564
rect 158180 183500 158181 183564
rect 158115 183499 158181 183500
rect 154794 156218 154826 156454
rect 155062 156218 155146 156454
rect 155382 156218 155414 156454
rect 154794 156134 155414 156218
rect 154794 155898 154826 156134
rect 155062 155898 155146 156134
rect 155382 155898 155414 156134
rect 154794 142000 155414 155898
rect 159294 160954 159914 196398
rect 160326 196077 160386 200227
rect 160507 200156 160573 200157
rect 160507 200092 160508 200156
rect 160572 200092 160573 200156
rect 160507 200091 160573 200092
rect 161427 200156 161493 200157
rect 161427 200092 161428 200156
rect 161492 200092 161493 200156
rect 161427 200091 161493 200092
rect 160510 196485 160570 200091
rect 160875 199884 160941 199885
rect 160875 199820 160876 199884
rect 160940 199820 160941 199884
rect 160875 199819 160941 199820
rect 161243 199884 161309 199885
rect 161243 199820 161244 199884
rect 161308 199820 161309 199884
rect 161243 199819 161309 199820
rect 160691 199748 160757 199749
rect 160691 199684 160692 199748
rect 160756 199684 160757 199748
rect 160691 199683 160757 199684
rect 160694 198797 160754 199683
rect 160878 199341 160938 199819
rect 161059 199612 161125 199613
rect 161059 199548 161060 199612
rect 161124 199548 161125 199612
rect 161059 199547 161125 199548
rect 160875 199340 160941 199341
rect 160875 199276 160876 199340
rect 160940 199276 160941 199340
rect 160875 199275 160941 199276
rect 160691 198796 160757 198797
rect 160691 198732 160692 198796
rect 160756 198732 160757 198796
rect 160691 198731 160757 198732
rect 160507 196484 160573 196485
rect 160507 196420 160508 196484
rect 160572 196420 160573 196484
rect 160507 196419 160573 196420
rect 160323 196076 160389 196077
rect 160323 196012 160324 196076
rect 160388 196012 160389 196076
rect 160323 196011 160389 196012
rect 161062 178805 161122 199547
rect 161246 199341 161306 199819
rect 161430 199613 161490 200091
rect 161427 199612 161493 199613
rect 161427 199548 161428 199612
rect 161492 199548 161493 199612
rect 161427 199547 161493 199548
rect 161614 199341 161674 200227
rect 168238 199885 168298 200771
rect 173019 200564 173085 200565
rect 173019 200500 173020 200564
rect 173084 200500 173085 200564
rect 173019 200499 173085 200500
rect 173022 199885 173082 200499
rect 176147 200428 176213 200429
rect 176147 200364 176148 200428
rect 176212 200364 176213 200428
rect 176147 200363 176213 200364
rect 161979 199884 162045 199885
rect 161979 199820 161980 199884
rect 162044 199820 162045 199884
rect 161979 199819 162045 199820
rect 162531 199884 162597 199885
rect 162531 199820 162532 199884
rect 162596 199820 162597 199884
rect 162531 199819 162597 199820
rect 162899 199884 162965 199885
rect 162899 199820 162900 199884
rect 162964 199820 162965 199884
rect 162899 199819 162965 199820
rect 163819 199884 163885 199885
rect 163819 199820 163820 199884
rect 163884 199820 163885 199884
rect 163819 199819 163885 199820
rect 164187 199884 164253 199885
rect 164187 199820 164188 199884
rect 164252 199820 164253 199884
rect 164187 199819 164253 199820
rect 165107 199884 165173 199885
rect 165107 199820 165108 199884
rect 165172 199820 165173 199884
rect 165107 199819 165173 199820
rect 166027 199884 166093 199885
rect 166027 199820 166028 199884
rect 166092 199820 166093 199884
rect 166027 199819 166093 199820
rect 168051 199884 168117 199885
rect 168051 199820 168052 199884
rect 168116 199820 168117 199884
rect 168051 199819 168117 199820
rect 168235 199884 168301 199885
rect 168235 199820 168236 199884
rect 168300 199820 168301 199884
rect 168235 199819 168301 199820
rect 168971 199884 169037 199885
rect 168971 199820 168972 199884
rect 169036 199820 169037 199884
rect 168971 199819 169037 199820
rect 169707 199884 169773 199885
rect 169707 199820 169708 199884
rect 169772 199820 169773 199884
rect 169707 199819 169773 199820
rect 170443 199884 170509 199885
rect 170443 199820 170444 199884
rect 170508 199820 170509 199884
rect 170443 199819 170509 199820
rect 172283 199884 172349 199885
rect 172283 199820 172284 199884
rect 172348 199820 172349 199884
rect 172283 199819 172349 199820
rect 173019 199884 173085 199885
rect 173019 199820 173020 199884
rect 173084 199820 173085 199884
rect 173019 199819 173085 199820
rect 173203 199884 173269 199885
rect 173203 199820 173204 199884
rect 173268 199820 173269 199884
rect 173203 199819 173269 199820
rect 174123 199884 174189 199885
rect 174123 199820 174124 199884
rect 174188 199820 174189 199884
rect 174123 199819 174189 199820
rect 161243 199340 161309 199341
rect 161243 199276 161244 199340
rect 161308 199276 161309 199340
rect 161243 199275 161309 199276
rect 161611 199340 161677 199341
rect 161611 199276 161612 199340
rect 161676 199276 161677 199340
rect 161611 199275 161677 199276
rect 161243 196076 161309 196077
rect 161243 196012 161244 196076
rect 161308 196012 161309 196076
rect 161243 196011 161309 196012
rect 161246 178941 161306 196011
rect 161982 193901 162042 199819
rect 162163 199612 162229 199613
rect 162163 199548 162164 199612
rect 162228 199548 162229 199612
rect 162163 199547 162229 199548
rect 162166 195533 162226 199547
rect 162534 199341 162594 199819
rect 162902 199341 162962 199819
rect 162531 199340 162597 199341
rect 162531 199276 162532 199340
rect 162596 199276 162597 199340
rect 162531 199275 162597 199276
rect 162899 199340 162965 199341
rect 162899 199276 162900 199340
rect 162964 199276 162965 199340
rect 162899 199275 162965 199276
rect 163822 196349 163882 199819
rect 163819 196348 163885 196349
rect 163819 196284 163820 196348
rect 163884 196284 163885 196348
rect 163819 196283 163885 196284
rect 164003 196076 164069 196077
rect 164003 196012 164004 196076
rect 164068 196012 164069 196076
rect 164003 196011 164069 196012
rect 162163 195532 162229 195533
rect 162163 195468 162164 195532
rect 162228 195468 162229 195532
rect 162163 195467 162229 195468
rect 161979 193900 162045 193901
rect 161979 193836 161980 193900
rect 162044 193836 162045 193900
rect 161979 193835 162045 193836
rect 164006 184653 164066 196011
rect 164190 191317 164250 199819
rect 165110 196213 165170 199819
rect 165475 198796 165541 198797
rect 165475 198732 165476 198796
rect 165540 198732 165541 198796
rect 165475 198731 165541 198732
rect 165291 198116 165357 198117
rect 165291 198052 165292 198116
rect 165356 198052 165357 198116
rect 165291 198051 165357 198052
rect 165107 196212 165173 196213
rect 165107 196148 165108 196212
rect 165172 196148 165173 196212
rect 165107 196147 165173 196148
rect 164187 191316 164253 191317
rect 164187 191252 164188 191316
rect 164252 191252 164253 191316
rect 164187 191251 164253 191252
rect 164003 184652 164069 184653
rect 164003 184588 164004 184652
rect 164068 184588 164069 184652
rect 164003 184587 164069 184588
rect 165294 179349 165354 198051
rect 165291 179348 165357 179349
rect 165291 179284 165292 179348
rect 165356 179284 165357 179348
rect 165291 179283 165357 179284
rect 161243 178940 161309 178941
rect 161243 178876 161244 178940
rect 161308 178876 161309 178940
rect 161243 178875 161309 178876
rect 161059 178804 161125 178805
rect 161059 178740 161060 178804
rect 161124 178740 161125 178804
rect 161059 178739 161125 178740
rect 159294 160718 159326 160954
rect 159562 160718 159646 160954
rect 159882 160718 159914 160954
rect 159294 160634 159914 160718
rect 159294 160398 159326 160634
rect 159562 160398 159646 160634
rect 159882 160398 159914 160634
rect 159294 142000 159914 160398
rect 165478 148341 165538 198731
rect 166030 195669 166090 199819
rect 166395 199748 166461 199749
rect 166395 199684 166396 199748
rect 166460 199684 166461 199748
rect 166395 199683 166461 199684
rect 166211 198116 166277 198117
rect 166211 198052 166212 198116
rect 166276 198052 166277 198116
rect 166211 198051 166277 198052
rect 166027 195668 166093 195669
rect 166027 195604 166028 195668
rect 166092 195604 166093 195668
rect 166027 195603 166093 195604
rect 166214 190229 166274 198051
rect 166211 190228 166277 190229
rect 166211 190164 166212 190228
rect 166276 190164 166277 190228
rect 166211 190163 166277 190164
rect 166398 184517 166458 199683
rect 167499 199476 167565 199477
rect 167499 199412 167500 199476
rect 167564 199412 167565 199476
rect 167499 199411 167565 199412
rect 166579 198524 166645 198525
rect 166579 198460 166580 198524
rect 166644 198460 166645 198524
rect 166579 198459 166645 198460
rect 166395 184516 166461 184517
rect 166395 184452 166396 184516
rect 166460 184452 166461 184516
rect 166395 184451 166461 184452
rect 166582 180165 166642 198459
rect 166763 196348 166829 196349
rect 166763 196284 166764 196348
rect 166828 196284 166829 196348
rect 166763 196283 166829 196284
rect 166579 180164 166645 180165
rect 166579 180100 166580 180164
rect 166644 180100 166645 180164
rect 166579 180099 166645 180100
rect 166766 180029 166826 196283
rect 167502 189141 167562 199411
rect 168054 196213 168114 199819
rect 168235 198116 168301 198117
rect 168235 198052 168236 198116
rect 168300 198052 168301 198116
rect 168235 198051 168301 198052
rect 168051 196212 168117 196213
rect 168051 196148 168052 196212
rect 168116 196148 168117 196212
rect 168051 196147 168117 196148
rect 168238 190773 168298 198051
rect 168974 196349 169034 199819
rect 169155 199748 169221 199749
rect 169155 199684 169156 199748
rect 169220 199684 169221 199748
rect 169155 199683 169221 199684
rect 168971 196348 169037 196349
rect 168971 196284 168972 196348
rect 169036 196284 169037 196348
rect 168971 196283 169037 196284
rect 168971 196076 169037 196077
rect 168971 196012 168972 196076
rect 169036 196012 169037 196076
rect 168971 196011 169037 196012
rect 168235 190772 168301 190773
rect 168235 190708 168236 190772
rect 168300 190708 168301 190772
rect 168235 190707 168301 190708
rect 167499 189140 167565 189141
rect 167499 189076 167500 189140
rect 167564 189076 167565 189140
rect 167499 189075 167565 189076
rect 168974 184245 169034 196011
rect 169158 186149 169218 199683
rect 169339 199204 169405 199205
rect 169339 199140 169340 199204
rect 169404 199140 169405 199204
rect 169339 199139 169405 199140
rect 169155 186148 169221 186149
rect 169155 186084 169156 186148
rect 169220 186084 169221 186148
rect 169155 186083 169221 186084
rect 168971 184244 169037 184245
rect 168971 184180 168972 184244
rect 169036 184180 169037 184244
rect 168971 184179 169037 184180
rect 169342 180573 169402 199139
rect 169710 195261 169770 199819
rect 170446 197370 170506 199819
rect 170995 199612 171061 199613
rect 170995 199548 170996 199612
rect 171060 199548 171061 199612
rect 170995 199547 171061 199548
rect 170811 199204 170877 199205
rect 170811 199140 170812 199204
rect 170876 199140 170877 199204
rect 170811 199139 170877 199140
rect 170262 197310 170506 197370
rect 169707 195260 169773 195261
rect 169707 195196 169708 195260
rect 169772 195196 169773 195260
rect 169707 195195 169773 195196
rect 170262 187781 170322 197310
rect 170814 195533 170874 199139
rect 170811 195532 170877 195533
rect 170811 195468 170812 195532
rect 170876 195468 170877 195532
rect 170811 195467 170877 195468
rect 170259 187780 170325 187781
rect 170259 187716 170260 187780
rect 170324 187716 170325 187780
rect 170259 187715 170325 187716
rect 170998 184381 171058 199547
rect 172286 189549 172346 199819
rect 172467 198660 172533 198661
rect 172467 198596 172468 198660
rect 172532 198596 172533 198660
rect 172467 198595 172533 198596
rect 172470 195397 172530 198595
rect 173206 198389 173266 199819
rect 173571 199748 173637 199749
rect 173571 199684 173572 199748
rect 173636 199684 173637 199748
rect 173571 199683 173637 199684
rect 173203 198388 173269 198389
rect 173203 198324 173204 198388
rect 173268 198324 173269 198388
rect 173203 198323 173269 198324
rect 173574 196893 173634 199683
rect 173755 199612 173821 199613
rect 173755 199548 173756 199612
rect 173820 199548 173821 199612
rect 173755 199547 173821 199548
rect 173571 196892 173637 196893
rect 173571 196828 173572 196892
rect 173636 196828 173637 196892
rect 173571 196827 173637 196828
rect 172467 195396 172533 195397
rect 172467 195332 172468 195396
rect 172532 195332 172533 195396
rect 172467 195331 172533 195332
rect 172283 189548 172349 189549
rect 172283 189484 172284 189548
rect 172348 189484 172349 189548
rect 172283 189483 172349 189484
rect 173758 186013 173818 199547
rect 174126 198661 174186 199819
rect 174859 199748 174925 199749
rect 174859 199684 174860 199748
rect 174924 199684 174925 199748
rect 174859 199683 174925 199684
rect 174123 198660 174189 198661
rect 174123 198596 174124 198660
rect 174188 198596 174189 198660
rect 174123 198595 174189 198596
rect 174491 198116 174557 198117
rect 174491 198052 174492 198116
rect 174556 198052 174557 198116
rect 174491 198051 174557 198052
rect 174307 196892 174373 196893
rect 174307 196828 174308 196892
rect 174372 196828 174373 196892
rect 174307 196827 174373 196828
rect 174310 191589 174370 196827
rect 174307 191588 174373 191589
rect 174307 191524 174308 191588
rect 174372 191524 174373 191588
rect 174307 191523 174373 191524
rect 173755 186012 173821 186013
rect 173755 185948 173756 186012
rect 173820 185948 173821 186012
rect 173755 185947 173821 185948
rect 174494 185605 174554 198051
rect 174862 189957 174922 199683
rect 176150 199613 176210 200363
rect 176334 199613 176394 201451
rect 186086 200701 186146 205590
rect 186822 200837 186882 220899
rect 186819 200836 186885 200837
rect 186819 200772 186820 200836
rect 186884 200772 186885 200836
rect 186819 200771 186885 200772
rect 186083 200700 186149 200701
rect 186083 200636 186084 200700
rect 186148 200636 186149 200700
rect 186083 200635 186149 200636
rect 177067 200156 177133 200157
rect 177067 200092 177068 200156
rect 177132 200092 177133 200156
rect 177067 200091 177133 200092
rect 176791 199884 176857 199885
rect 176791 199882 176792 199884
rect 176518 199822 176792 199882
rect 176147 199612 176213 199613
rect 176147 199548 176148 199612
rect 176212 199548 176213 199612
rect 176147 199547 176213 199548
rect 176331 199612 176397 199613
rect 176331 199548 176332 199612
rect 176396 199548 176397 199612
rect 176331 199547 176397 199548
rect 175595 198660 175661 198661
rect 175595 198596 175596 198660
rect 175660 198596 175661 198660
rect 175595 198595 175661 198596
rect 175598 192813 175658 198595
rect 176518 194717 176578 199822
rect 176791 199820 176792 199822
rect 176856 199820 176857 199884
rect 176791 199819 176857 199820
rect 177070 199613 177130 200091
rect 177251 199884 177317 199885
rect 177251 199820 177252 199884
rect 177316 199820 177317 199884
rect 177251 199819 177317 199820
rect 177067 199612 177133 199613
rect 177067 199548 177068 199612
rect 177132 199548 177133 199612
rect 177067 199547 177133 199548
rect 177254 198658 177314 199819
rect 177070 198598 177314 198658
rect 177070 196077 177130 198598
rect 177067 196076 177133 196077
rect 177067 196012 177068 196076
rect 177132 196012 177133 196076
rect 177067 196011 177133 196012
rect 176515 194716 176581 194717
rect 176515 194652 176516 194716
rect 176580 194652 176581 194716
rect 176515 194651 176581 194652
rect 175595 192812 175661 192813
rect 175595 192748 175596 192812
rect 175660 192748 175661 192812
rect 175595 192747 175661 192748
rect 174859 189956 174925 189957
rect 174859 189892 174860 189956
rect 174924 189892 174925 189956
rect 174859 189891 174925 189892
rect 174491 185604 174557 185605
rect 174491 185540 174492 185604
rect 174556 185540 174557 185604
rect 174491 185539 174557 185540
rect 170995 184380 171061 184381
rect 170995 184316 170996 184380
rect 171060 184316 171061 184380
rect 170995 184315 171061 184316
rect 169339 180572 169405 180573
rect 169339 180508 169340 180572
rect 169404 180508 169405 180572
rect 169339 180507 169405 180508
rect 166763 180028 166829 180029
rect 166763 179964 166764 180028
rect 166828 179964 166829 180028
rect 166763 179963 166829 179964
rect 177294 178954 177914 198000
rect 177294 178718 177326 178954
rect 177562 178718 177646 178954
rect 177882 178718 177914 178954
rect 177294 178634 177914 178718
rect 177294 178398 177326 178634
rect 177562 178398 177646 178634
rect 177882 178398 177914 178634
rect 165475 148340 165541 148341
rect 165475 148276 165476 148340
rect 165540 148276 165541 148340
rect 165475 148275 165541 148276
rect 177294 142954 177914 178398
rect 177294 142718 177326 142954
rect 177562 142718 177646 142954
rect 177882 142718 177914 142954
rect 177294 142634 177914 142718
rect 177294 142398 177326 142634
rect 177562 142398 177646 142634
rect 177882 142398 177914 142634
rect 177294 142000 177914 142398
rect 181794 183454 182414 198000
rect 182771 188460 182837 188461
rect 182771 188396 182772 188460
rect 182836 188396 182837 188460
rect 182771 188395 182837 188396
rect 181794 183218 181826 183454
rect 182062 183218 182146 183454
rect 182382 183218 182414 183454
rect 181794 183134 182414 183218
rect 181794 182898 181826 183134
rect 182062 182898 182146 183134
rect 182382 182898 182414 183134
rect 181794 147454 182414 182898
rect 181794 147218 181826 147454
rect 182062 147218 182146 147454
rect 182382 147218 182414 147454
rect 181794 147134 182414 147218
rect 181794 146898 181826 147134
rect 182062 146898 182146 147134
rect 182382 146898 182414 147134
rect 181794 142000 182414 146898
rect 151123 140316 151189 140317
rect 151123 140252 151124 140316
rect 151188 140252 151189 140316
rect 151123 140251 151189 140252
rect 124259 139636 124325 139637
rect 124259 139572 124260 139636
rect 124324 139572 124325 139636
rect 124259 139571 124325 139572
rect 124262 139093 124322 139571
rect 130699 139500 130765 139501
rect 130699 139436 130700 139500
rect 130764 139436 130765 139500
rect 130699 139435 130765 139436
rect 124259 139092 124325 139093
rect 124259 139028 124260 139092
rect 124324 139028 124325 139092
rect 124259 139027 124325 139028
rect 130702 138549 130762 139435
rect 176515 139364 176581 139365
rect 176515 139300 176516 139364
rect 176580 139300 176581 139364
rect 176515 139299 176581 139300
rect 176518 138685 176578 139299
rect 176515 138684 176581 138685
rect 176515 138620 176516 138684
rect 176580 138620 176581 138684
rect 176515 138619 176581 138620
rect 130699 138548 130765 138549
rect 130699 138484 130700 138548
rect 130764 138484 130765 138548
rect 130699 138483 130765 138484
rect 182774 137869 182834 188395
rect 186294 187954 186914 198000
rect 186294 187718 186326 187954
rect 186562 187718 186646 187954
rect 186882 187718 186914 187954
rect 186294 187634 186914 187718
rect 186294 187398 186326 187634
rect 186562 187398 186646 187634
rect 186882 187398 186914 187634
rect 186083 179076 186149 179077
rect 186083 179012 186084 179076
rect 186148 179012 186149 179076
rect 186083 179011 186149 179012
rect 185163 178668 185229 178669
rect 185163 178604 185164 178668
rect 185228 178604 185229 178668
rect 185163 178603 185229 178604
rect 183139 139500 183205 139501
rect 183139 139436 183140 139500
rect 183204 139436 183205 139500
rect 183139 139435 183205 139436
rect 183142 138549 183202 139435
rect 183139 138548 183205 138549
rect 183139 138484 183140 138548
rect 183204 138484 183205 138548
rect 183139 138483 183205 138484
rect 185166 138141 185226 178603
rect 186086 141130 186146 179011
rect 186294 151954 186914 187398
rect 186294 151718 186326 151954
rect 186562 151718 186646 151954
rect 186882 151718 186914 151954
rect 186294 151634 186914 151718
rect 186294 151398 186326 151634
rect 186562 151398 186646 151634
rect 186882 151398 186914 151634
rect 186294 142000 186914 151398
rect 187006 143445 187066 259931
rect 187923 259724 187989 259725
rect 187923 259660 187924 259724
rect 187988 259660 187989 259724
rect 187923 259659 187989 259660
rect 187187 259588 187253 259589
rect 187187 259524 187188 259588
rect 187252 259524 187253 259588
rect 187187 259523 187253 259524
rect 187190 200701 187250 259523
rect 187187 200700 187253 200701
rect 187187 200636 187188 200700
rect 187252 200636 187253 200700
rect 187187 200635 187253 200636
rect 187739 193356 187805 193357
rect 187739 193292 187740 193356
rect 187804 193292 187805 193356
rect 187739 193291 187805 193292
rect 187187 179212 187253 179213
rect 187187 179148 187188 179212
rect 187252 179148 187253 179212
rect 187187 179147 187253 179148
rect 187003 143444 187069 143445
rect 187003 143380 187004 143444
rect 187068 143380 187069 143444
rect 187003 143379 187069 143380
rect 186086 141070 186514 141130
rect 186267 140724 186333 140725
rect 186267 140660 186268 140724
rect 186332 140660 186333 140724
rect 186267 140659 186333 140660
rect 185899 140588 185965 140589
rect 185899 140524 185900 140588
rect 185964 140524 185965 140588
rect 185899 140523 185965 140524
rect 185902 140450 185962 140523
rect 185902 140390 186146 140450
rect 185163 138140 185229 138141
rect 185163 138076 185164 138140
rect 185228 138076 185229 138140
rect 185163 138075 185229 138076
rect 182771 137868 182837 137869
rect 182771 137804 182772 137868
rect 182836 137804 182837 137868
rect 182771 137803 182837 137804
rect 186086 134469 186146 140390
rect 186270 137325 186330 140659
rect 186267 137324 186333 137325
rect 186267 137260 186268 137324
rect 186332 137260 186333 137324
rect 186267 137259 186333 137260
rect 186454 137050 186514 141070
rect 187003 140316 187069 140317
rect 187003 140252 187004 140316
rect 187068 140252 187069 140316
rect 187003 140251 187069 140252
rect 186635 139500 186701 139501
rect 186635 139436 186636 139500
rect 186700 139436 186701 139500
rect 186635 139435 186701 139436
rect 186638 138005 186698 139435
rect 186635 138004 186701 138005
rect 186635 137940 186636 138004
rect 186700 137940 186701 138004
rect 186635 137939 186701 137940
rect 186819 137868 186885 137869
rect 186819 137804 186820 137868
rect 186884 137804 186885 137868
rect 186819 137803 186885 137804
rect 186270 136990 186514 137050
rect 186270 136645 186330 136990
rect 186267 136644 186333 136645
rect 186267 136580 186268 136644
rect 186332 136580 186333 136644
rect 186267 136579 186333 136580
rect 186083 134468 186149 134469
rect 186083 134404 186084 134468
rect 186148 134404 186149 134468
rect 186083 134403 186149 134404
rect 186083 133788 186149 133789
rect 186083 133724 186084 133788
rect 186148 133724 186149 133788
rect 186083 133723 186149 133724
rect 139568 115954 139888 115986
rect 139568 115718 139610 115954
rect 139846 115718 139888 115954
rect 139568 115634 139888 115718
rect 139568 115398 139610 115634
rect 139846 115398 139888 115634
rect 139568 115366 139888 115398
rect 170288 115954 170608 115986
rect 170288 115718 170330 115954
rect 170566 115718 170608 115954
rect 170288 115634 170608 115718
rect 170288 115398 170330 115634
rect 170566 115398 170608 115634
rect 170288 115366 170608 115398
rect 124208 111454 124528 111486
rect 124208 111218 124250 111454
rect 124486 111218 124528 111454
rect 124208 111134 124528 111218
rect 124208 110898 124250 111134
rect 124486 110898 124528 111134
rect 124208 110866 124528 110898
rect 154928 111454 155248 111486
rect 154928 111218 154970 111454
rect 155206 111218 155248 111454
rect 154928 111134 155248 111218
rect 154928 110898 154970 111134
rect 155206 110898 155248 111134
rect 154928 110866 155248 110898
rect 185648 111454 185968 111486
rect 185648 111218 185690 111454
rect 185926 111218 185968 111454
rect 185648 111134 185968 111218
rect 185648 110898 185690 111134
rect 185926 110898 185968 111134
rect 185648 110866 185968 110898
rect 186086 91221 186146 133723
rect 186083 91220 186149 91221
rect 186083 91156 186084 91220
rect 186148 91156 186149 91220
rect 186083 91155 186149 91156
rect 186822 88365 186882 137803
rect 187006 91901 187066 140251
rect 187190 137461 187250 179147
rect 187371 138140 187437 138141
rect 187371 138076 187372 138140
rect 187436 138076 187437 138140
rect 187371 138075 187437 138076
rect 187187 137460 187253 137461
rect 187187 137396 187188 137460
rect 187252 137396 187253 137460
rect 187187 137395 187253 137396
rect 187374 135965 187434 138075
rect 187371 135964 187437 135965
rect 187371 135900 187372 135964
rect 187436 135900 187437 135964
rect 187371 135899 187437 135900
rect 187003 91900 187069 91901
rect 187003 91836 187004 91900
rect 187068 91836 187069 91900
rect 187003 91835 187069 91836
rect 187187 91220 187253 91221
rect 187187 91156 187188 91220
rect 187252 91156 187253 91220
rect 187187 91155 187253 91156
rect 186819 88364 186885 88365
rect 186819 88300 186820 88364
rect 186884 88300 186885 88364
rect 186819 88299 186885 88300
rect 187003 83468 187069 83469
rect 187003 83404 187004 83468
rect 187068 83404 187069 83468
rect 187003 83403 187069 83404
rect 186083 82108 186149 82109
rect 186083 82044 186084 82108
rect 186148 82044 186149 82108
rect 186083 82043 186149 82044
rect 133459 81972 133525 81973
rect 133459 81908 133460 81972
rect 133524 81908 133525 81972
rect 133459 81907 133525 81908
rect 172651 81972 172717 81973
rect 172651 81908 172652 81972
rect 172716 81908 172717 81972
rect 172651 81907 172717 81908
rect 132171 81836 132237 81837
rect 132171 81772 132172 81836
rect 132236 81772 132237 81836
rect 132171 81771 132237 81772
rect 129779 81700 129845 81701
rect 129779 81636 129780 81700
rect 129844 81636 129845 81700
rect 129779 81635 129845 81636
rect 124075 80612 124141 80613
rect 124075 80548 124076 80612
rect 124140 80548 124141 80612
rect 124075 80547 124141 80548
rect 123891 78164 123957 78165
rect 123891 78100 123892 78164
rect 123956 78100 123957 78164
rect 123891 78099 123957 78100
rect 122603 68916 122669 68917
rect 122603 68852 122604 68916
rect 122668 68852 122669 68916
rect 122603 68851 122669 68852
rect 119843 66196 119909 66197
rect 119843 66132 119844 66196
rect 119908 66132 119909 66196
rect 119843 66131 119909 66132
rect 118794 48218 118826 48454
rect 119062 48218 119146 48454
rect 119382 48218 119414 48454
rect 118794 48134 119414 48218
rect 118794 47898 118826 48134
rect 119062 47898 119146 48134
rect 119382 47898 119414 48134
rect 118794 12454 119414 47898
rect 118794 12218 118826 12454
rect 119062 12218 119146 12454
rect 119382 12218 119414 12454
rect 118794 12134 119414 12218
rect 118794 11898 118826 12134
rect 119062 11898 119146 12134
rect 119382 11898 119414 12134
rect 118794 -2266 119414 11898
rect 118794 -2502 118826 -2266
rect 119062 -2502 119146 -2266
rect 119382 -2502 119414 -2266
rect 118794 -2586 119414 -2502
rect 118794 -2822 118826 -2586
rect 119062 -2822 119146 -2586
rect 119382 -2822 119414 -2586
rect 118794 -7654 119414 -2822
rect 123294 52954 123914 78000
rect 123294 52718 123326 52954
rect 123562 52718 123646 52954
rect 123882 52718 123914 52954
rect 123294 52634 123914 52718
rect 123294 52398 123326 52634
rect 123562 52398 123646 52634
rect 123882 52398 123914 52634
rect 123294 16954 123914 52398
rect 123294 16718 123326 16954
rect 123562 16718 123646 16954
rect 123882 16718 123914 16954
rect 123294 16634 123914 16718
rect 123294 16398 123326 16634
rect 123562 16398 123646 16634
rect 123882 16398 123914 16634
rect 123294 -3226 123914 16398
rect 123294 -3462 123326 -3226
rect 123562 -3462 123646 -3226
rect 123882 -3462 123914 -3226
rect 123294 -3546 123914 -3462
rect 123294 -3782 123326 -3546
rect 123562 -3782 123646 -3546
rect 123882 -3782 123914 -3546
rect 123294 -7654 123914 -3782
rect 127794 57454 128414 78000
rect 129782 76397 129842 81635
rect 132174 80749 132234 81771
rect 132171 80748 132237 80749
rect 132171 80684 132172 80748
rect 132236 80684 132237 80748
rect 132171 80683 132237 80684
rect 133091 79932 133157 79933
rect 133091 79868 133092 79932
rect 133156 79868 133157 79932
rect 133091 79867 133157 79868
rect 133094 78709 133154 79867
rect 133462 79661 133522 81907
rect 135483 81428 135549 81429
rect 135483 81364 135484 81428
rect 135548 81364 135549 81428
rect 135483 81363 135549 81364
rect 134563 81020 134629 81021
rect 134563 80956 134564 81020
rect 134628 80956 134629 81020
rect 134563 80955 134629 80956
rect 133827 80748 133893 80749
rect 133827 80684 133828 80748
rect 133892 80684 133893 80748
rect 133827 80683 133893 80684
rect 133643 79932 133709 79933
rect 133643 79868 133644 79932
rect 133708 79868 133709 79932
rect 133643 79867 133709 79868
rect 133459 79660 133525 79661
rect 133459 79596 133460 79660
rect 133524 79596 133525 79660
rect 133459 79595 133525 79596
rect 133091 78708 133157 78709
rect 133091 78644 133092 78708
rect 133156 78644 133157 78708
rect 133091 78643 133157 78644
rect 133091 78436 133157 78437
rect 133091 78372 133092 78436
rect 133156 78372 133157 78436
rect 133091 78371 133157 78372
rect 129779 76396 129845 76397
rect 129779 76332 129780 76396
rect 129844 76332 129845 76396
rect 129779 76331 129845 76332
rect 127794 57218 127826 57454
rect 128062 57218 128146 57454
rect 128382 57218 128414 57454
rect 127794 57134 128414 57218
rect 127794 56898 127826 57134
rect 128062 56898 128146 57134
rect 128382 56898 128414 57134
rect 127794 21454 128414 56898
rect 127794 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 128414 21454
rect 127794 21134 128414 21218
rect 127794 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 128414 21134
rect 127794 -4186 128414 20898
rect 127794 -4422 127826 -4186
rect 128062 -4422 128146 -4186
rect 128382 -4422 128414 -4186
rect 127794 -4506 128414 -4422
rect 127794 -4742 127826 -4506
rect 128062 -4742 128146 -4506
rect 128382 -4742 128414 -4506
rect 127794 -7654 128414 -4742
rect 132294 61954 132914 78000
rect 133094 70277 133154 78371
rect 133646 75173 133706 79867
rect 133830 79797 133890 80683
rect 134011 79932 134077 79933
rect 134011 79868 134012 79932
rect 134076 79868 134077 79932
rect 134011 79867 134077 79868
rect 133827 79796 133893 79797
rect 133827 79732 133828 79796
rect 133892 79732 133893 79796
rect 133827 79731 133893 79732
rect 134014 79661 134074 79867
rect 134566 79797 134626 80955
rect 134931 80340 134997 80341
rect 134931 80276 134932 80340
rect 134996 80276 134997 80340
rect 134931 80275 134997 80276
rect 134563 79796 134629 79797
rect 134563 79732 134564 79796
rect 134628 79732 134629 79796
rect 134563 79731 134629 79732
rect 134934 79661 134994 80275
rect 135486 79933 135546 81363
rect 138795 81292 138861 81293
rect 138795 81228 138796 81292
rect 138860 81228 138861 81292
rect 138795 81227 138861 81228
rect 171915 81292 171981 81293
rect 171915 81228 171916 81292
rect 171980 81228 171981 81292
rect 171915 81227 171981 81228
rect 136587 80612 136653 80613
rect 136587 80548 136588 80612
rect 136652 80548 136653 80612
rect 136587 80547 136653 80548
rect 135483 79932 135549 79933
rect 135483 79868 135484 79932
rect 135548 79868 135549 79932
rect 135483 79867 135549 79868
rect 136403 79932 136469 79933
rect 136403 79868 136404 79932
rect 136468 79868 136469 79932
rect 136403 79867 136469 79868
rect 134011 79660 134077 79661
rect 134011 79596 134012 79660
rect 134076 79596 134077 79660
rect 134011 79595 134077 79596
rect 134931 79660 134997 79661
rect 134931 79596 134932 79660
rect 134996 79596 134997 79660
rect 134931 79595 134997 79596
rect 135115 78300 135181 78301
rect 135115 78236 135116 78300
rect 135180 78236 135181 78300
rect 135115 78235 135181 78236
rect 134011 76260 134077 76261
rect 134011 76196 134012 76260
rect 134076 76196 134077 76260
rect 134011 76195 134077 76196
rect 133643 75172 133709 75173
rect 133643 75108 133644 75172
rect 133708 75108 133709 75172
rect 133643 75107 133709 75108
rect 133091 70276 133157 70277
rect 133091 70212 133092 70276
rect 133156 70212 133157 70276
rect 133091 70211 133157 70212
rect 134014 64890 134074 76195
rect 135118 74085 135178 78235
rect 136406 78029 136466 79867
rect 136590 79661 136650 80547
rect 137139 80204 137205 80205
rect 137139 80140 137140 80204
rect 137204 80202 137205 80204
rect 137507 80204 137573 80205
rect 137507 80202 137508 80204
rect 137204 80142 137508 80202
rect 137204 80140 137205 80142
rect 137139 80139 137205 80140
rect 137507 80140 137508 80142
rect 137572 80140 137573 80204
rect 137507 80139 137573 80140
rect 138798 79933 138858 81227
rect 151491 81156 151557 81157
rect 151491 81092 151492 81156
rect 151556 81092 151557 81156
rect 151491 81091 151557 81092
rect 158667 81156 158733 81157
rect 158667 81092 158668 81156
rect 158732 81092 158733 81156
rect 158667 81091 158733 81092
rect 139899 80884 139965 80885
rect 139899 80820 139900 80884
rect 139964 80820 139965 80884
rect 139899 80819 139965 80820
rect 136771 79932 136837 79933
rect 136771 79868 136772 79932
rect 136836 79868 136837 79932
rect 136771 79867 136837 79868
rect 138427 79932 138493 79933
rect 138427 79868 138428 79932
rect 138492 79868 138493 79932
rect 138427 79867 138493 79868
rect 138795 79932 138861 79933
rect 138795 79868 138796 79932
rect 138860 79868 138861 79932
rect 138795 79867 138861 79868
rect 139531 79932 139597 79933
rect 139531 79868 139532 79932
rect 139596 79868 139597 79932
rect 139531 79867 139597 79868
rect 136587 79660 136653 79661
rect 136587 79596 136588 79660
rect 136652 79596 136653 79660
rect 136587 79595 136653 79596
rect 136774 78301 136834 79867
rect 138243 79796 138309 79797
rect 138243 79732 138244 79796
rect 138308 79732 138309 79796
rect 138243 79731 138309 79732
rect 136771 78300 136837 78301
rect 136771 78236 136772 78300
rect 136836 78236 136837 78300
rect 136771 78235 136837 78236
rect 136587 78164 136653 78165
rect 136587 78100 136588 78164
rect 136652 78100 136653 78164
rect 136587 78099 136653 78100
rect 136403 78028 136469 78029
rect 136403 77964 136404 78028
rect 136468 77964 136469 78028
rect 136403 77963 136469 77964
rect 135851 77348 135917 77349
rect 135851 77284 135852 77348
rect 135916 77284 135917 77348
rect 135851 77283 135917 77284
rect 135299 77212 135365 77213
rect 135299 77148 135300 77212
rect 135364 77148 135365 77212
rect 135299 77147 135365 77148
rect 135115 74084 135181 74085
rect 135115 74020 135116 74084
rect 135180 74020 135181 74084
rect 135115 74019 135181 74020
rect 135302 71093 135362 77147
rect 135299 71092 135365 71093
rect 135299 71028 135300 71092
rect 135364 71028 135365 71092
rect 135299 71027 135365 71028
rect 135854 68509 135914 77283
rect 136590 72589 136650 78099
rect 138059 78028 138125 78029
rect 136587 72588 136653 72589
rect 136587 72524 136588 72588
rect 136652 72524 136653 72588
rect 136587 72523 136653 72524
rect 135851 68508 135917 68509
rect 135851 68444 135852 68508
rect 135916 68444 135917 68508
rect 135851 68443 135917 68444
rect 133830 64837 134074 64890
rect 133827 64836 134074 64837
rect 133827 64772 133828 64836
rect 133892 64830 134074 64836
rect 136794 66454 137414 78000
rect 138059 77964 138060 78028
rect 138124 77964 138125 78028
rect 138059 77963 138125 77964
rect 138062 68645 138122 77963
rect 138246 69597 138306 79731
rect 138430 76533 138490 79867
rect 139347 79796 139413 79797
rect 139347 79732 139348 79796
rect 139412 79732 139413 79796
rect 139347 79731 139413 79732
rect 138611 78708 138677 78709
rect 138611 78644 138612 78708
rect 138676 78644 138677 78708
rect 138611 78643 138677 78644
rect 138427 76532 138493 76533
rect 138427 76468 138428 76532
rect 138492 76468 138493 76532
rect 138427 76467 138493 76468
rect 138243 69596 138309 69597
rect 138243 69532 138244 69596
rect 138308 69532 138309 69596
rect 138243 69531 138309 69532
rect 138059 68644 138125 68645
rect 138059 68580 138060 68644
rect 138124 68580 138125 68644
rect 138059 68579 138125 68580
rect 138614 67421 138674 78643
rect 139350 68373 139410 79731
rect 139534 78573 139594 79867
rect 139902 79797 139962 80819
rect 140267 80068 140333 80069
rect 140267 80004 140268 80068
rect 140332 80004 140333 80068
rect 140267 80003 140333 80004
rect 145051 80068 145117 80069
rect 145051 80004 145052 80068
rect 145116 80004 145117 80068
rect 145051 80003 145117 80004
rect 139899 79796 139965 79797
rect 139899 79732 139900 79796
rect 139964 79732 139965 79796
rect 139899 79731 139965 79732
rect 139531 78572 139597 78573
rect 139531 78508 139532 78572
rect 139596 78508 139597 78572
rect 139531 78507 139597 78508
rect 140270 71365 140330 80003
rect 141555 79932 141621 79933
rect 141555 79868 141556 79932
rect 141620 79868 141621 79932
rect 142107 79932 142173 79933
rect 142107 79930 142108 79932
rect 141555 79867 141621 79868
rect 141926 79870 142108 79930
rect 141558 78573 141618 79867
rect 141555 78572 141621 78573
rect 141555 78508 141556 78572
rect 141620 78508 141621 78572
rect 141555 78507 141621 78508
rect 141926 78301 141986 79870
rect 142107 79868 142108 79870
rect 142172 79868 142173 79932
rect 142107 79867 142173 79868
rect 143947 79932 144013 79933
rect 143947 79868 143948 79932
rect 144012 79868 144013 79932
rect 143947 79867 144013 79868
rect 144867 79932 144933 79933
rect 144867 79868 144868 79932
rect 144932 79868 144933 79932
rect 144867 79867 144933 79868
rect 143579 79796 143645 79797
rect 143579 79732 143580 79796
rect 143644 79732 143645 79796
rect 143579 79731 143645 79732
rect 142107 79660 142173 79661
rect 142107 79596 142108 79660
rect 142172 79596 142173 79660
rect 142107 79595 142173 79596
rect 141923 78300 141989 78301
rect 141923 78236 141924 78300
rect 141988 78236 141989 78300
rect 141923 78235 141989 78236
rect 140635 78028 140701 78029
rect 140635 77964 140636 78028
rect 140700 77964 140701 78028
rect 140635 77963 140701 77964
rect 140451 77484 140517 77485
rect 140451 77420 140452 77484
rect 140516 77420 140517 77484
rect 140451 77419 140517 77420
rect 140454 73133 140514 77419
rect 140638 76669 140698 77963
rect 140635 76668 140701 76669
rect 140635 76604 140636 76668
rect 140700 76604 140701 76668
rect 140635 76603 140701 76604
rect 140819 76668 140885 76669
rect 140819 76604 140820 76668
rect 140884 76604 140885 76668
rect 140819 76603 140885 76604
rect 140451 73132 140517 73133
rect 140451 73068 140452 73132
rect 140516 73068 140517 73132
rect 140451 73067 140517 73068
rect 140267 71364 140333 71365
rect 140267 71300 140268 71364
rect 140332 71300 140333 71364
rect 140267 71299 140333 71300
rect 140822 68781 140882 76603
rect 141294 70954 141914 78000
rect 141294 70718 141326 70954
rect 141562 70718 141646 70954
rect 141882 70718 141914 70954
rect 141294 70634 141914 70718
rect 141294 70398 141326 70634
rect 141562 70398 141646 70634
rect 141882 70398 141914 70634
rect 142110 70413 142170 79595
rect 142291 78708 142357 78709
rect 142291 78644 142292 78708
rect 142356 78644 142357 78708
rect 142291 78643 142357 78644
rect 142294 71501 142354 78643
rect 142659 77892 142725 77893
rect 142659 77828 142660 77892
rect 142724 77828 142725 77892
rect 142659 77827 142725 77828
rect 142291 71500 142357 71501
rect 142291 71436 142292 71500
rect 142356 71436 142357 71500
rect 142291 71435 142357 71436
rect 140819 68780 140885 68781
rect 140819 68716 140820 68780
rect 140884 68716 140885 68780
rect 140819 68715 140885 68716
rect 139347 68372 139413 68373
rect 139347 68308 139348 68372
rect 139412 68308 139413 68372
rect 139347 68307 139413 68308
rect 138611 67420 138677 67421
rect 138611 67356 138612 67420
rect 138676 67356 138677 67420
rect 138611 67355 138677 67356
rect 136794 66218 136826 66454
rect 137062 66218 137146 66454
rect 137382 66218 137414 66454
rect 136794 66134 137414 66218
rect 136794 65898 136826 66134
rect 137062 65898 137146 66134
rect 137382 65898 137414 66134
rect 133892 64772 133893 64830
rect 133827 64771 133893 64772
rect 133830 63477 133890 64771
rect 133827 63476 133893 63477
rect 133827 63412 133828 63476
rect 133892 63412 133893 63476
rect 133827 63411 133893 63412
rect 132294 61718 132326 61954
rect 132562 61718 132646 61954
rect 132882 61718 132914 61954
rect 132294 61634 132914 61718
rect 132294 61398 132326 61634
rect 132562 61398 132646 61634
rect 132882 61398 132914 61634
rect 132294 25954 132914 61398
rect 132294 25718 132326 25954
rect 132562 25718 132646 25954
rect 132882 25718 132914 25954
rect 132294 25634 132914 25718
rect 132294 25398 132326 25634
rect 132562 25398 132646 25634
rect 132882 25398 132914 25634
rect 132294 -5146 132914 25398
rect 132294 -5382 132326 -5146
rect 132562 -5382 132646 -5146
rect 132882 -5382 132914 -5146
rect 132294 -5466 132914 -5382
rect 132294 -5702 132326 -5466
rect 132562 -5702 132646 -5466
rect 132882 -5702 132914 -5466
rect 132294 -7654 132914 -5702
rect 136794 30454 137414 65898
rect 136794 30218 136826 30454
rect 137062 30218 137146 30454
rect 137382 30218 137414 30454
rect 136794 30134 137414 30218
rect 136794 29898 136826 30134
rect 137062 29898 137146 30134
rect 137382 29898 137414 30134
rect 136794 -6106 137414 29898
rect 136794 -6342 136826 -6106
rect 137062 -6342 137146 -6106
rect 137382 -6342 137414 -6106
rect 136794 -6426 137414 -6342
rect 136794 -6662 136826 -6426
rect 137062 -6662 137146 -6426
rect 137382 -6662 137414 -6426
rect 136794 -7654 137414 -6662
rect 141294 34954 141914 70398
rect 142107 70412 142173 70413
rect 142107 70348 142108 70412
rect 142172 70348 142173 70412
rect 142107 70347 142173 70348
rect 142662 70141 142722 77827
rect 142659 70140 142725 70141
rect 142659 70076 142660 70140
rect 142724 70076 142725 70140
rect 142659 70075 142725 70076
rect 143582 70005 143642 79731
rect 143763 78708 143829 78709
rect 143763 78644 143764 78708
rect 143828 78644 143829 78708
rect 143763 78643 143829 78644
rect 143579 70004 143645 70005
rect 143579 69940 143580 70004
rect 143644 69940 143645 70004
rect 143579 69939 143645 69940
rect 143766 69461 143826 78643
rect 143950 76669 144010 79867
rect 144870 76669 144930 79867
rect 143947 76668 144013 76669
rect 143947 76604 143948 76668
rect 144012 76604 144013 76668
rect 143947 76603 144013 76604
rect 144867 76668 144933 76669
rect 144867 76604 144868 76668
rect 144932 76604 144933 76668
rect 144867 76603 144933 76604
rect 143763 69460 143829 69461
rect 143763 69396 143764 69460
rect 143828 69396 143829 69460
rect 143763 69395 143829 69396
rect 145054 68917 145114 80003
rect 151494 79933 151554 81091
rect 157379 81020 157445 81021
rect 157379 80956 157380 81020
rect 157444 80956 157445 81020
rect 157379 80955 157445 80956
rect 152227 80748 152293 80749
rect 152227 80684 152228 80748
rect 152292 80684 152293 80748
rect 152227 80683 152293 80684
rect 146155 79932 146221 79933
rect 146155 79868 146156 79932
rect 146220 79868 146221 79932
rect 146155 79867 146221 79868
rect 146523 79932 146589 79933
rect 146523 79868 146524 79932
rect 146588 79868 146589 79932
rect 146523 79867 146589 79868
rect 147075 79932 147141 79933
rect 147075 79868 147076 79932
rect 147140 79868 147141 79932
rect 147075 79867 147141 79868
rect 148179 79932 148245 79933
rect 148179 79868 148180 79932
rect 148244 79868 148245 79932
rect 148179 79867 148245 79868
rect 148731 79932 148797 79933
rect 148731 79868 148732 79932
rect 148796 79868 148797 79932
rect 148731 79867 148797 79868
rect 151491 79932 151557 79933
rect 151491 79868 151492 79932
rect 151556 79868 151557 79932
rect 151491 79867 151557 79868
rect 152043 79932 152109 79933
rect 152043 79868 152044 79932
rect 152108 79868 152109 79932
rect 152043 79867 152109 79868
rect 146158 78845 146218 79867
rect 146155 78844 146221 78845
rect 146155 78780 146156 78844
rect 146220 78780 146221 78844
rect 146155 78779 146221 78780
rect 145794 75454 146414 78000
rect 146526 75717 146586 79867
rect 146707 76668 146773 76669
rect 146707 76604 146708 76668
rect 146772 76604 146773 76668
rect 146707 76603 146773 76604
rect 146523 75716 146589 75717
rect 146523 75652 146524 75716
rect 146588 75652 146589 75716
rect 146523 75651 146589 75652
rect 145794 75218 145826 75454
rect 146062 75218 146146 75454
rect 146382 75218 146414 75454
rect 145794 75134 146414 75218
rect 145794 74898 145826 75134
rect 146062 74898 146146 75134
rect 146382 74898 146414 75134
rect 145051 68916 145117 68917
rect 145051 68852 145052 68916
rect 145116 68852 145117 68916
rect 145051 68851 145117 68852
rect 141294 34718 141326 34954
rect 141562 34718 141646 34954
rect 141882 34718 141914 34954
rect 141294 34634 141914 34718
rect 141294 34398 141326 34634
rect 141562 34398 141646 34634
rect 141882 34398 141914 34634
rect 141294 -7066 141914 34398
rect 141294 -7302 141326 -7066
rect 141562 -7302 141646 -7066
rect 141882 -7302 141914 -7066
rect 141294 -7386 141914 -7302
rect 141294 -7622 141326 -7386
rect 141562 -7622 141646 -7386
rect 141882 -7622 141914 -7386
rect 141294 -7654 141914 -7622
rect 145794 39454 146414 74898
rect 146710 72997 146770 76603
rect 147078 74901 147138 79867
rect 147811 79796 147877 79797
rect 147811 79732 147812 79796
rect 147876 79794 147877 79796
rect 147876 79734 148058 79794
rect 147876 79732 147877 79734
rect 147811 79731 147877 79732
rect 147075 74900 147141 74901
rect 147075 74836 147076 74900
rect 147140 74836 147141 74900
rect 147075 74835 147141 74836
rect 146707 72996 146773 72997
rect 146707 72932 146708 72996
rect 146772 72932 146773 72996
rect 146707 72931 146773 72932
rect 147998 72453 148058 79734
rect 148182 77757 148242 79867
rect 148179 77756 148245 77757
rect 148179 77692 148180 77756
rect 148244 77692 148245 77756
rect 148179 77691 148245 77692
rect 148734 74901 148794 79867
rect 149467 79660 149533 79661
rect 149467 79596 149468 79660
rect 149532 79596 149533 79660
rect 149467 79595 149533 79596
rect 148731 74900 148797 74901
rect 148731 74836 148732 74900
rect 148796 74836 148797 74900
rect 148731 74835 148797 74836
rect 147995 72452 148061 72453
rect 147995 72388 147996 72452
rect 148060 72388 148061 72452
rect 147995 72387 148061 72388
rect 149470 70957 149530 79595
rect 149467 70956 149533 70957
rect 149467 70892 149468 70956
rect 149532 70892 149533 70956
rect 149467 70891 149533 70892
rect 145794 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 146414 39454
rect 145794 39134 146414 39218
rect 145794 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 146414 39134
rect 145794 3454 146414 38898
rect 145794 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 146414 3454
rect 145794 3134 146414 3218
rect 145794 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 146414 3134
rect 145794 -346 146414 2898
rect 145794 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 146414 -346
rect 145794 -666 146414 -582
rect 145794 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 146414 -666
rect 145794 -7654 146414 -902
rect 150294 43954 150914 78000
rect 152046 72861 152106 79867
rect 152230 79525 152290 80683
rect 155539 80204 155605 80205
rect 155539 80140 155540 80204
rect 155604 80140 155605 80204
rect 155539 80139 155605 80140
rect 152963 79932 153029 79933
rect 152963 79868 152964 79932
rect 153028 79868 153029 79932
rect 152963 79867 153029 79868
rect 154435 79932 154501 79933
rect 154435 79868 154436 79932
rect 154500 79868 154501 79932
rect 154435 79867 154501 79868
rect 152227 79524 152293 79525
rect 152227 79460 152228 79524
rect 152292 79460 152293 79524
rect 152227 79459 152293 79460
rect 152966 77893 153026 79867
rect 154438 79253 154498 79867
rect 154987 79796 155053 79797
rect 154987 79732 154988 79796
rect 155052 79732 155053 79796
rect 154987 79731 155053 79732
rect 154619 79660 154685 79661
rect 154619 79596 154620 79660
rect 154684 79596 154685 79660
rect 154619 79595 154685 79596
rect 154435 79252 154501 79253
rect 154435 79188 154436 79252
rect 154500 79188 154501 79252
rect 154435 79187 154501 79188
rect 154622 78573 154682 79595
rect 154990 78573 155050 79731
rect 154619 78572 154685 78573
rect 154619 78508 154620 78572
rect 154684 78508 154685 78572
rect 154619 78507 154685 78508
rect 154987 78572 155053 78573
rect 154987 78508 154988 78572
rect 155052 78508 155053 78572
rect 154987 78507 155053 78508
rect 152963 77892 153029 77893
rect 152963 77828 152964 77892
rect 153028 77828 153029 77892
rect 152963 77827 153029 77828
rect 152963 75988 153029 75989
rect 152963 75924 152964 75988
rect 153028 75924 153029 75988
rect 152963 75923 153029 75924
rect 154251 75988 154317 75989
rect 154251 75924 154252 75988
rect 154316 75924 154317 75988
rect 154251 75923 154317 75924
rect 152043 72860 152109 72861
rect 152043 72796 152044 72860
rect 152108 72796 152109 72860
rect 152043 72795 152109 72796
rect 152966 67557 153026 75923
rect 152963 67556 153029 67557
rect 152963 67492 152964 67556
rect 153028 67492 153029 67556
rect 152963 67491 153029 67492
rect 154254 66197 154314 75923
rect 154435 75852 154501 75853
rect 154435 75788 154436 75852
rect 154500 75788 154501 75852
rect 154435 75787 154501 75788
rect 154251 66196 154317 66197
rect 154251 66132 154252 66196
rect 154316 66132 154317 66196
rect 154251 66131 154317 66132
rect 154438 66061 154498 75787
rect 154435 66060 154501 66061
rect 154435 65996 154436 66060
rect 154500 65996 154501 66060
rect 154435 65995 154501 65996
rect 150294 43718 150326 43954
rect 150562 43718 150646 43954
rect 150882 43718 150914 43954
rect 150294 43634 150914 43718
rect 150294 43398 150326 43634
rect 150562 43398 150646 43634
rect 150882 43398 150914 43634
rect 150294 7954 150914 43398
rect 150294 7718 150326 7954
rect 150562 7718 150646 7954
rect 150882 7718 150914 7954
rect 150294 7634 150914 7718
rect 150294 7398 150326 7634
rect 150562 7398 150646 7634
rect 150882 7398 150914 7634
rect 150294 -1306 150914 7398
rect 150294 -1542 150326 -1306
rect 150562 -1542 150646 -1306
rect 150882 -1542 150914 -1306
rect 150294 -1626 150914 -1542
rect 150294 -1862 150326 -1626
rect 150562 -1862 150646 -1626
rect 150882 -1862 150914 -1626
rect 150294 -7654 150914 -1862
rect 154794 48454 155414 78000
rect 155542 71773 155602 80139
rect 157382 79933 157442 80955
rect 158670 79933 158730 81091
rect 164739 80884 164805 80885
rect 164739 80820 164740 80884
rect 164804 80820 164805 80884
rect 164739 80819 164805 80820
rect 164742 79933 164802 80819
rect 171731 80476 171797 80477
rect 171731 80412 171732 80476
rect 171796 80412 171797 80476
rect 171731 80411 171797 80412
rect 157379 79932 157445 79933
rect 157379 79868 157380 79932
rect 157444 79868 157445 79932
rect 157379 79867 157445 79868
rect 158483 79932 158549 79933
rect 158483 79868 158484 79932
rect 158548 79868 158549 79932
rect 158483 79867 158549 79868
rect 158667 79932 158733 79933
rect 158667 79868 158668 79932
rect 158732 79868 158733 79932
rect 158667 79867 158733 79868
rect 160875 79932 160941 79933
rect 160875 79868 160876 79932
rect 160940 79868 160941 79932
rect 160875 79867 160941 79868
rect 161059 79932 161125 79933
rect 161059 79868 161060 79932
rect 161124 79868 161125 79932
rect 161059 79867 161125 79868
rect 161611 79932 161677 79933
rect 161611 79868 161612 79932
rect 161676 79868 161677 79932
rect 161611 79867 161677 79868
rect 162531 79932 162597 79933
rect 162531 79868 162532 79932
rect 162596 79868 162597 79932
rect 162531 79867 162597 79868
rect 163083 79932 163149 79933
rect 163083 79868 163084 79932
rect 163148 79868 163149 79932
rect 163083 79867 163149 79868
rect 163267 79932 163333 79933
rect 163267 79868 163268 79932
rect 163332 79868 163333 79932
rect 163267 79867 163333 79868
rect 164371 79932 164437 79933
rect 164371 79868 164372 79932
rect 164436 79868 164437 79932
rect 164371 79867 164437 79868
rect 164739 79932 164805 79933
rect 164739 79868 164740 79932
rect 164804 79868 164805 79932
rect 164739 79867 164805 79868
rect 164923 79932 164989 79933
rect 164923 79868 164924 79932
rect 164988 79868 164989 79932
rect 164923 79867 164989 79868
rect 167683 79932 167749 79933
rect 167683 79868 167684 79932
rect 167748 79868 167749 79932
rect 167683 79867 167749 79868
rect 170443 79932 170509 79933
rect 170443 79868 170444 79932
rect 170508 79868 170509 79932
rect 170443 79867 170509 79868
rect 158115 79796 158181 79797
rect 158115 79732 158116 79796
rect 158180 79732 158181 79796
rect 158115 79731 158181 79732
rect 156459 76668 156525 76669
rect 156459 76604 156460 76668
rect 156524 76604 156525 76668
rect 156459 76603 156525 76604
rect 155539 71772 155605 71773
rect 155539 71708 155540 71772
rect 155604 71708 155605 71772
rect 155539 71707 155605 71708
rect 156462 71093 156522 76603
rect 157931 75988 157997 75989
rect 157931 75924 157932 75988
rect 157996 75924 157997 75988
rect 157931 75923 157997 75924
rect 156459 71092 156525 71093
rect 156459 71028 156460 71092
rect 156524 71028 156525 71092
rect 156459 71027 156525 71028
rect 157934 67013 157994 75923
rect 158118 71637 158178 79731
rect 158486 77893 158546 79867
rect 160691 79388 160757 79389
rect 160691 79324 160692 79388
rect 160756 79324 160757 79388
rect 160691 79323 160757 79324
rect 158483 77892 158549 77893
rect 158483 77828 158484 77892
rect 158548 77828 158549 77892
rect 158483 77827 158549 77828
rect 158115 71636 158181 71637
rect 158115 71572 158116 71636
rect 158180 71572 158181 71636
rect 158115 71571 158181 71572
rect 157931 67012 157997 67013
rect 157931 66948 157932 67012
rect 157996 66948 157997 67012
rect 157931 66947 157997 66948
rect 154794 48218 154826 48454
rect 155062 48218 155146 48454
rect 155382 48218 155414 48454
rect 154794 48134 155414 48218
rect 154794 47898 154826 48134
rect 155062 47898 155146 48134
rect 155382 47898 155414 48134
rect 154794 12454 155414 47898
rect 154794 12218 154826 12454
rect 155062 12218 155146 12454
rect 155382 12218 155414 12454
rect 154794 12134 155414 12218
rect 154794 11898 154826 12134
rect 155062 11898 155146 12134
rect 155382 11898 155414 12134
rect 154794 -2266 155414 11898
rect 154794 -2502 154826 -2266
rect 155062 -2502 155146 -2266
rect 155382 -2502 155414 -2266
rect 154794 -2586 155414 -2502
rect 154794 -2822 154826 -2586
rect 155062 -2822 155146 -2586
rect 155382 -2822 155414 -2586
rect 154794 -7654 155414 -2822
rect 159294 52954 159914 78000
rect 160694 65925 160754 79323
rect 160878 77485 160938 79867
rect 160875 77484 160941 77485
rect 160875 77420 160876 77484
rect 160940 77420 160941 77484
rect 160875 77419 160941 77420
rect 160691 65924 160757 65925
rect 160691 65860 160692 65924
rect 160756 65860 160757 65924
rect 160691 65859 160757 65860
rect 161062 63341 161122 79867
rect 161427 78028 161493 78029
rect 161427 77964 161428 78028
rect 161492 77964 161493 78028
rect 161427 77963 161493 77964
rect 161430 75717 161490 77963
rect 161427 75716 161493 75717
rect 161427 75652 161428 75716
rect 161492 75652 161493 75716
rect 161427 75651 161493 75652
rect 161614 75581 161674 79867
rect 162534 76669 162594 79867
rect 162715 79796 162781 79797
rect 162715 79732 162716 79796
rect 162780 79732 162781 79796
rect 162715 79731 162781 79732
rect 162718 78573 162778 79731
rect 163086 79117 163146 79867
rect 163270 79389 163330 79867
rect 164374 79794 164434 79867
rect 164374 79734 164802 79794
rect 163267 79388 163333 79389
rect 163267 79324 163268 79388
rect 163332 79324 163333 79388
rect 163267 79323 163333 79324
rect 163083 79116 163149 79117
rect 163083 79052 163084 79116
rect 163148 79052 163149 79116
rect 163083 79051 163149 79052
rect 162715 78572 162781 78573
rect 162715 78508 162716 78572
rect 162780 78508 162781 78572
rect 162715 78507 162781 78508
rect 162531 76668 162597 76669
rect 162531 76604 162532 76668
rect 162596 76604 162597 76668
rect 162531 76603 162597 76604
rect 161611 75580 161677 75581
rect 161611 75516 161612 75580
rect 161676 75516 161677 75580
rect 161611 75515 161677 75516
rect 161059 63340 161125 63341
rect 161059 63276 161060 63340
rect 161124 63276 161125 63340
rect 161059 63275 161125 63276
rect 159294 52718 159326 52954
rect 159562 52718 159646 52954
rect 159882 52718 159914 52954
rect 159294 52634 159914 52718
rect 159294 52398 159326 52634
rect 159562 52398 159646 52634
rect 159882 52398 159914 52634
rect 159294 16954 159914 52398
rect 159294 16718 159326 16954
rect 159562 16718 159646 16954
rect 159882 16718 159914 16954
rect 159294 16634 159914 16718
rect 159294 16398 159326 16634
rect 159562 16398 159646 16634
rect 159882 16398 159914 16634
rect 159294 -3226 159914 16398
rect 159294 -3462 159326 -3226
rect 159562 -3462 159646 -3226
rect 159882 -3462 159914 -3226
rect 159294 -3546 159914 -3462
rect 159294 -3782 159326 -3546
rect 159562 -3782 159646 -3546
rect 159882 -3782 159914 -3546
rect 159294 -7654 159914 -3782
rect 163794 57454 164414 78000
rect 164742 77077 164802 79734
rect 164926 79525 164986 79867
rect 165107 79796 165173 79797
rect 165107 79732 165108 79796
rect 165172 79732 165173 79796
rect 166763 79796 166829 79797
rect 166763 79794 166764 79796
rect 165107 79731 165173 79732
rect 166582 79734 166764 79794
rect 164923 79524 164989 79525
rect 164923 79460 164924 79524
rect 164988 79460 164989 79524
rect 164923 79459 164989 79460
rect 164739 77076 164805 77077
rect 164739 77012 164740 77076
rect 164804 77012 164805 77076
rect 164739 77011 164805 77012
rect 165110 68373 165170 79731
rect 166211 75036 166277 75037
rect 166211 74972 166212 75036
rect 166276 74972 166277 75036
rect 166211 74971 166277 74972
rect 166214 68781 166274 74971
rect 166582 73813 166642 79734
rect 166763 79732 166764 79734
rect 166828 79732 166829 79796
rect 166763 79731 166829 79732
rect 166763 78980 166829 78981
rect 166763 78916 166764 78980
rect 166828 78916 166829 78980
rect 166763 78915 166829 78916
rect 166579 73812 166645 73813
rect 166579 73748 166580 73812
rect 166644 73748 166645 73812
rect 166579 73747 166645 73748
rect 166211 68780 166277 68781
rect 166211 68716 166212 68780
rect 166276 68716 166277 68780
rect 166211 68715 166277 68716
rect 165107 68372 165173 68373
rect 165107 68308 165108 68372
rect 165172 68308 165173 68372
rect 165107 68307 165173 68308
rect 166766 64429 166826 78915
rect 167686 71501 167746 79867
rect 167867 79796 167933 79797
rect 167867 79732 167868 79796
rect 167932 79732 167933 79796
rect 167867 79731 167933 79732
rect 167683 71500 167749 71501
rect 167683 71436 167684 71500
rect 167748 71436 167749 71500
rect 167683 71435 167749 71436
rect 166763 64428 166829 64429
rect 166763 64364 166764 64428
rect 166828 64364 166829 64428
rect 166763 64363 166829 64364
rect 167870 64293 167930 79731
rect 168051 78980 168117 78981
rect 168051 78916 168052 78980
rect 168116 78916 168117 78980
rect 168051 78915 168117 78916
rect 167867 64292 167933 64293
rect 167867 64228 167868 64292
rect 167932 64228 167933 64292
rect 167867 64227 167933 64228
rect 168054 64157 168114 78915
rect 169155 78436 169221 78437
rect 169155 78372 169156 78436
rect 169220 78372 169221 78436
rect 169155 78371 169221 78372
rect 168051 64156 168117 64157
rect 168051 64092 168052 64156
rect 168116 64092 168117 64156
rect 168051 64091 168117 64092
rect 163794 57218 163826 57454
rect 164062 57218 164146 57454
rect 164382 57218 164414 57454
rect 163794 57134 164414 57218
rect 163794 56898 163826 57134
rect 164062 56898 164146 57134
rect 164382 56898 164414 57134
rect 163794 21454 164414 56898
rect 163794 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 164414 21454
rect 163794 21134 164414 21218
rect 163794 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 164414 21134
rect 163794 -4186 164414 20898
rect 163794 -4422 163826 -4186
rect 164062 -4422 164146 -4186
rect 164382 -4422 164414 -4186
rect 163794 -4506 164414 -4422
rect 163794 -4742 163826 -4506
rect 164062 -4742 164146 -4506
rect 164382 -4742 164414 -4506
rect 163794 -7654 164414 -4742
rect 168294 61954 168914 78000
rect 169158 64021 169218 78371
rect 170259 76668 170325 76669
rect 170259 76604 170260 76668
rect 170324 76604 170325 76668
rect 170259 76603 170325 76604
rect 170262 73813 170322 76603
rect 170446 75989 170506 79867
rect 171734 79797 171794 80411
rect 170811 79796 170877 79797
rect 170811 79732 170812 79796
rect 170876 79732 170877 79796
rect 170811 79731 170877 79732
rect 171731 79796 171797 79797
rect 171731 79732 171732 79796
rect 171796 79732 171797 79796
rect 171731 79731 171797 79732
rect 170627 77076 170693 77077
rect 170627 77012 170628 77076
rect 170692 77012 170693 77076
rect 170627 77011 170693 77012
rect 170443 75988 170509 75989
rect 170443 75924 170444 75988
rect 170508 75924 170509 75988
rect 170443 75923 170509 75924
rect 170630 74493 170690 77011
rect 170627 74492 170693 74493
rect 170627 74428 170628 74492
rect 170692 74428 170693 74492
rect 170627 74427 170693 74428
rect 170259 73812 170325 73813
rect 170259 73748 170260 73812
rect 170324 73748 170325 73812
rect 170259 73747 170325 73748
rect 170814 68917 170874 79731
rect 170995 79660 171061 79661
rect 170995 79596 170996 79660
rect 171060 79596 171061 79660
rect 170995 79595 171061 79596
rect 170811 68916 170877 68917
rect 170811 68852 170812 68916
rect 170876 68852 170877 68916
rect 170811 68851 170877 68852
rect 170998 65789 171058 79595
rect 171918 78981 171978 81227
rect 172283 80068 172349 80069
rect 172283 80004 172284 80068
rect 172348 80004 172349 80068
rect 172283 80003 172349 80004
rect 171915 78980 171981 78981
rect 171915 78916 171916 78980
rect 171980 78916 171981 78980
rect 171915 78915 171981 78916
rect 171731 78436 171797 78437
rect 171731 78372 171732 78436
rect 171796 78372 171797 78436
rect 171731 78371 171797 78372
rect 171734 69733 171794 78371
rect 172286 73170 172346 80003
rect 172467 79932 172533 79933
rect 172467 79868 172468 79932
rect 172532 79868 172533 79932
rect 172467 79867 172533 79868
rect 172470 78573 172530 79867
rect 172654 79797 172714 81907
rect 175227 81836 175293 81837
rect 175227 81772 175228 81836
rect 175292 81772 175293 81836
rect 175227 81771 175293 81772
rect 175230 80885 175290 81771
rect 185531 81700 185597 81701
rect 185531 81636 185532 81700
rect 185596 81636 185597 81700
rect 185531 81635 185597 81636
rect 175227 80884 175293 80885
rect 175227 80820 175228 80884
rect 175292 80820 175293 80884
rect 175227 80819 175293 80820
rect 172835 79932 172901 79933
rect 172835 79868 172836 79932
rect 172900 79868 172901 79932
rect 172835 79867 172901 79868
rect 173571 79932 173637 79933
rect 173571 79868 173572 79932
rect 173636 79868 173637 79932
rect 173571 79867 173637 79868
rect 173755 79932 173821 79933
rect 173755 79868 173756 79932
rect 173820 79868 173821 79932
rect 173755 79867 173821 79868
rect 175963 79932 176029 79933
rect 175963 79868 175964 79932
rect 176028 79868 176029 79932
rect 175963 79867 176029 79868
rect 176331 79932 176397 79933
rect 176331 79868 176332 79932
rect 176396 79868 176397 79932
rect 176331 79867 176397 79868
rect 172651 79796 172717 79797
rect 172651 79732 172652 79796
rect 172716 79732 172717 79796
rect 172651 79731 172717 79732
rect 172838 78573 172898 79867
rect 172467 78572 172533 78573
rect 172467 78508 172468 78572
rect 172532 78508 172533 78572
rect 172467 78507 172533 78508
rect 172835 78572 172901 78573
rect 172835 78508 172836 78572
rect 172900 78508 172901 78572
rect 172835 78507 172901 78508
rect 172467 77756 172533 77757
rect 172467 77692 172468 77756
rect 172532 77692 172533 77756
rect 172467 77691 172533 77692
rect 172102 73110 172346 73170
rect 172470 73133 172530 77691
rect 172467 73132 172533 73133
rect 171731 69732 171797 69733
rect 171731 69668 171732 69732
rect 171796 69668 171797 69732
rect 171731 69667 171797 69668
rect 170995 65788 171061 65789
rect 170995 65724 170996 65788
rect 171060 65724 171061 65788
rect 170995 65723 171061 65724
rect 172102 64837 172162 73110
rect 172467 73068 172468 73132
rect 172532 73068 172533 73132
rect 172467 73067 172533 73068
rect 172794 66454 173414 78000
rect 173574 71365 173634 79867
rect 173758 77893 173818 79867
rect 174859 79796 174925 79797
rect 174859 79732 174860 79796
rect 174924 79732 174925 79796
rect 174859 79731 174925 79732
rect 174675 79660 174741 79661
rect 174675 79596 174676 79660
rect 174740 79596 174741 79660
rect 174675 79595 174741 79596
rect 173755 77892 173821 77893
rect 173755 77828 173756 77892
rect 173820 77828 173821 77892
rect 173755 77827 173821 77828
rect 173571 71364 173637 71365
rect 173571 71300 173572 71364
rect 173636 71300 173637 71364
rect 173571 71299 173637 71300
rect 174678 67285 174738 79595
rect 174862 69869 174922 79731
rect 175966 78573 176026 79867
rect 176334 78573 176394 79867
rect 185534 79389 185594 81635
rect 185531 79388 185597 79389
rect 185531 79324 185532 79388
rect 185596 79324 185597 79388
rect 185531 79323 185597 79324
rect 186086 79253 186146 82043
rect 186083 79252 186149 79253
rect 186083 79188 186084 79252
rect 186148 79188 186149 79252
rect 186083 79187 186149 79188
rect 175963 78572 176029 78573
rect 175963 78508 175964 78572
rect 176028 78508 176029 78572
rect 175963 78507 176029 78508
rect 176331 78572 176397 78573
rect 176331 78508 176332 78572
rect 176396 78508 176397 78572
rect 176331 78507 176397 78508
rect 176515 77892 176581 77893
rect 176515 77828 176516 77892
rect 176580 77828 176581 77892
rect 176515 77827 176581 77828
rect 176331 75036 176397 75037
rect 176331 74972 176332 75036
rect 176396 74972 176397 75036
rect 176331 74971 176397 74972
rect 174859 69868 174925 69869
rect 174859 69804 174860 69868
rect 174924 69804 174925 69868
rect 174859 69803 174925 69804
rect 174675 67284 174741 67285
rect 174675 67220 174676 67284
rect 174740 67220 174741 67284
rect 174675 67219 174741 67220
rect 176334 67149 176394 74971
rect 176331 67148 176397 67149
rect 176331 67084 176332 67148
rect 176396 67084 176397 67148
rect 176331 67083 176397 67084
rect 172794 66218 172826 66454
rect 173062 66218 173146 66454
rect 173382 66218 173414 66454
rect 172794 66134 173414 66218
rect 172794 65898 172826 66134
rect 173062 65898 173146 66134
rect 173382 65898 173414 66134
rect 172099 64836 172165 64837
rect 172099 64772 172100 64836
rect 172164 64772 172165 64836
rect 172099 64771 172165 64772
rect 169155 64020 169221 64021
rect 169155 63956 169156 64020
rect 169220 63956 169221 64020
rect 169155 63955 169221 63956
rect 168294 61718 168326 61954
rect 168562 61718 168646 61954
rect 168882 61718 168914 61954
rect 168294 61634 168914 61718
rect 168294 61398 168326 61634
rect 168562 61398 168646 61634
rect 168882 61398 168914 61634
rect 168294 25954 168914 61398
rect 168294 25718 168326 25954
rect 168562 25718 168646 25954
rect 168882 25718 168914 25954
rect 168294 25634 168914 25718
rect 168294 25398 168326 25634
rect 168562 25398 168646 25634
rect 168882 25398 168914 25634
rect 168294 -5146 168914 25398
rect 168294 -5382 168326 -5146
rect 168562 -5382 168646 -5146
rect 168882 -5382 168914 -5146
rect 168294 -5466 168914 -5382
rect 168294 -5702 168326 -5466
rect 168562 -5702 168646 -5466
rect 168882 -5702 168914 -5466
rect 168294 -7654 168914 -5702
rect 172794 30454 173414 65898
rect 176518 64701 176578 77827
rect 177294 70954 177914 78000
rect 177294 70718 177326 70954
rect 177562 70718 177646 70954
rect 177882 70718 177914 70954
rect 177294 70634 177914 70718
rect 177294 70398 177326 70634
rect 177562 70398 177646 70634
rect 177882 70398 177914 70634
rect 176515 64700 176581 64701
rect 176515 64636 176516 64700
rect 176580 64636 176581 64700
rect 176515 64635 176581 64636
rect 172794 30218 172826 30454
rect 173062 30218 173146 30454
rect 173382 30218 173414 30454
rect 172794 30134 173414 30218
rect 172794 29898 172826 30134
rect 173062 29898 173146 30134
rect 173382 29898 173414 30134
rect 172794 -6106 173414 29898
rect 172794 -6342 172826 -6106
rect 173062 -6342 173146 -6106
rect 173382 -6342 173414 -6106
rect 172794 -6426 173414 -6342
rect 172794 -6662 172826 -6426
rect 173062 -6662 173146 -6426
rect 173382 -6662 173414 -6426
rect 172794 -7654 173414 -6662
rect 177294 34954 177914 70398
rect 177294 34718 177326 34954
rect 177562 34718 177646 34954
rect 177882 34718 177914 34954
rect 177294 34634 177914 34718
rect 177294 34398 177326 34634
rect 177562 34398 177646 34634
rect 177882 34398 177914 34634
rect 177294 -7066 177914 34398
rect 177294 -7302 177326 -7066
rect 177562 -7302 177646 -7066
rect 177882 -7302 177914 -7066
rect 177294 -7386 177914 -7302
rect 177294 -7622 177326 -7386
rect 177562 -7622 177646 -7386
rect 177882 -7622 177914 -7386
rect 177294 -7654 177914 -7622
rect 181794 75454 182414 78000
rect 181794 75218 181826 75454
rect 182062 75218 182146 75454
rect 182382 75218 182414 75454
rect 181794 75134 182414 75218
rect 181794 74898 181826 75134
rect 182062 74898 182146 75134
rect 182382 74898 182414 75134
rect 181794 39454 182414 74898
rect 181794 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 182414 39454
rect 181794 39134 182414 39218
rect 181794 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 182414 39134
rect 181794 3454 182414 38898
rect 181794 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 182414 3454
rect 181794 3134 182414 3218
rect 181794 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 182414 3134
rect 181794 -346 182414 2898
rect 181794 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 182414 -346
rect 181794 -666 182414 -582
rect 181794 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 182414 -666
rect 181794 -7654 182414 -902
rect 186294 43954 186914 78000
rect 187006 75309 187066 83403
rect 187003 75308 187069 75309
rect 187003 75244 187004 75308
rect 187068 75244 187069 75308
rect 187003 75243 187069 75244
rect 187190 65517 187250 91155
rect 187742 78165 187802 193291
rect 187926 145757 187986 259659
rect 188291 233340 188357 233341
rect 188291 233276 188292 233340
rect 188356 233276 188357 233340
rect 188291 233275 188357 233276
rect 188294 198933 188354 233275
rect 188291 198932 188357 198933
rect 188291 198868 188292 198932
rect 188356 198868 188357 198932
rect 188291 198867 188357 198868
rect 190794 192454 191414 198000
rect 190794 192218 190826 192454
rect 191062 192218 191146 192454
rect 191382 192218 191414 192454
rect 190794 192134 191414 192218
rect 190794 191898 190826 192134
rect 191062 191898 191146 192134
rect 191382 191898 191414 192134
rect 190499 190228 190565 190229
rect 190499 190164 190500 190228
rect 190564 190164 190565 190228
rect 190499 190163 190565 190164
rect 189211 188324 189277 188325
rect 189211 188260 189212 188324
rect 189276 188260 189277 188324
rect 189211 188259 189277 188260
rect 189027 183428 189093 183429
rect 189027 183364 189028 183428
rect 189092 183364 189093 183428
rect 189027 183363 189093 183364
rect 189030 183157 189090 183363
rect 189027 183156 189093 183157
rect 189027 183092 189028 183156
rect 189092 183092 189093 183156
rect 189027 183091 189093 183092
rect 188843 182884 188909 182885
rect 188843 182820 188844 182884
rect 188908 182820 188909 182884
rect 188843 182819 188909 182820
rect 187923 145756 187989 145757
rect 187923 145692 187924 145756
rect 187988 145692 187989 145756
rect 187923 145691 187989 145692
rect 188846 137597 188906 182819
rect 189214 182610 189274 188259
rect 189579 183428 189645 183429
rect 189579 183364 189580 183428
rect 189644 183364 189645 183428
rect 189579 183363 189645 183364
rect 189030 182550 189274 182610
rect 188843 137596 188909 137597
rect 188843 137532 188844 137596
rect 188908 137532 188909 137596
rect 188843 137531 188909 137532
rect 187739 78164 187805 78165
rect 187739 78100 187740 78164
rect 187804 78100 187805 78164
rect 187739 78099 187805 78100
rect 189030 70957 189090 182550
rect 189582 181250 189642 183363
rect 189214 181190 189642 181250
rect 189214 79389 189274 181190
rect 189395 82244 189461 82245
rect 189395 82180 189396 82244
rect 189460 82180 189461 82244
rect 189395 82179 189461 82180
rect 189398 79525 189458 82179
rect 189395 79524 189461 79525
rect 189395 79460 189396 79524
rect 189460 79460 189461 79524
rect 189395 79459 189461 79460
rect 189211 79388 189277 79389
rect 189211 79324 189212 79388
rect 189276 79324 189277 79388
rect 189211 79323 189277 79324
rect 190502 76397 190562 190163
rect 190794 156454 191414 191898
rect 190794 156218 190826 156454
rect 191062 156218 191146 156454
rect 191382 156218 191414 156454
rect 190794 156134 191414 156218
rect 190794 155898 190826 156134
rect 191062 155898 191146 156134
rect 191382 155898 191414 156134
rect 190794 142000 191414 155898
rect 191790 143037 191850 263603
rect 191974 143173 192034 263739
rect 195294 232954 195914 268398
rect 195294 232718 195326 232954
rect 195562 232718 195646 232954
rect 195882 232718 195914 232954
rect 195294 232634 195914 232718
rect 195294 232398 195326 232634
rect 195562 232398 195646 232634
rect 195882 232398 195914 232634
rect 195294 196954 195914 232398
rect 195294 196718 195326 196954
rect 195562 196718 195646 196954
rect 195882 196718 195914 196954
rect 195294 196634 195914 196718
rect 195294 196398 195326 196634
rect 195562 196398 195646 196634
rect 195882 196398 195914 196634
rect 199794 708678 200414 711590
rect 199794 708442 199826 708678
rect 200062 708442 200146 708678
rect 200382 708442 200414 708678
rect 199794 708358 200414 708442
rect 199794 708122 199826 708358
rect 200062 708122 200146 708358
rect 200382 708122 200414 708358
rect 199794 669454 200414 708122
rect 199794 669218 199826 669454
rect 200062 669218 200146 669454
rect 200382 669218 200414 669454
rect 199794 669134 200414 669218
rect 199794 668898 199826 669134
rect 200062 668898 200146 669134
rect 200382 668898 200414 669134
rect 199794 633454 200414 668898
rect 199794 633218 199826 633454
rect 200062 633218 200146 633454
rect 200382 633218 200414 633454
rect 199794 633134 200414 633218
rect 199794 632898 199826 633134
rect 200062 632898 200146 633134
rect 200382 632898 200414 633134
rect 199794 597454 200414 632898
rect 199794 597218 199826 597454
rect 200062 597218 200146 597454
rect 200382 597218 200414 597454
rect 199794 597134 200414 597218
rect 199794 596898 199826 597134
rect 200062 596898 200146 597134
rect 200382 596898 200414 597134
rect 199794 561454 200414 596898
rect 199794 561218 199826 561454
rect 200062 561218 200146 561454
rect 200382 561218 200414 561454
rect 199794 561134 200414 561218
rect 199794 560898 199826 561134
rect 200062 560898 200146 561134
rect 200382 560898 200414 561134
rect 199794 525454 200414 560898
rect 199794 525218 199826 525454
rect 200062 525218 200146 525454
rect 200382 525218 200414 525454
rect 199794 525134 200414 525218
rect 199794 524898 199826 525134
rect 200062 524898 200146 525134
rect 200382 524898 200414 525134
rect 199794 489454 200414 524898
rect 199794 489218 199826 489454
rect 200062 489218 200146 489454
rect 200382 489218 200414 489454
rect 199794 489134 200414 489218
rect 199794 488898 199826 489134
rect 200062 488898 200146 489134
rect 200382 488898 200414 489134
rect 199794 453454 200414 488898
rect 199794 453218 199826 453454
rect 200062 453218 200146 453454
rect 200382 453218 200414 453454
rect 199794 453134 200414 453218
rect 199794 452898 199826 453134
rect 200062 452898 200146 453134
rect 200382 452898 200414 453134
rect 199794 417454 200414 452898
rect 199794 417218 199826 417454
rect 200062 417218 200146 417454
rect 200382 417218 200414 417454
rect 199794 417134 200414 417218
rect 199794 416898 199826 417134
rect 200062 416898 200146 417134
rect 200382 416898 200414 417134
rect 199794 381454 200414 416898
rect 199794 381218 199826 381454
rect 200062 381218 200146 381454
rect 200382 381218 200414 381454
rect 199794 381134 200414 381218
rect 199794 380898 199826 381134
rect 200062 380898 200146 381134
rect 200382 380898 200414 381134
rect 199794 345454 200414 380898
rect 199794 345218 199826 345454
rect 200062 345218 200146 345454
rect 200382 345218 200414 345454
rect 199794 345134 200414 345218
rect 199794 344898 199826 345134
rect 200062 344898 200146 345134
rect 200382 344898 200414 345134
rect 199794 309454 200414 344898
rect 199794 309218 199826 309454
rect 200062 309218 200146 309454
rect 200382 309218 200414 309454
rect 199794 309134 200414 309218
rect 199794 308898 199826 309134
rect 200062 308898 200146 309134
rect 200382 308898 200414 309134
rect 199794 273454 200414 308898
rect 199794 273218 199826 273454
rect 200062 273218 200146 273454
rect 200382 273218 200414 273454
rect 199794 273134 200414 273218
rect 199794 272898 199826 273134
rect 200062 272898 200146 273134
rect 200382 272898 200414 273134
rect 199794 237454 200414 272898
rect 199794 237218 199826 237454
rect 200062 237218 200146 237454
rect 200382 237218 200414 237454
rect 199794 237134 200414 237218
rect 199794 236898 199826 237134
rect 200062 236898 200146 237134
rect 200382 236898 200414 237134
rect 199794 201454 200414 236898
rect 199794 201218 199826 201454
rect 200062 201218 200146 201454
rect 200382 201218 200414 201454
rect 199794 201134 200414 201218
rect 199794 200898 199826 201134
rect 200062 200898 200146 201134
rect 200382 200898 200414 201134
rect 196019 196484 196085 196485
rect 196019 196420 196020 196484
rect 196084 196420 196085 196484
rect 196019 196419 196085 196420
rect 193259 191180 193325 191181
rect 193259 191116 193260 191180
rect 193324 191116 193325 191180
rect 193259 191115 193325 191116
rect 192155 189820 192221 189821
rect 192155 189756 192156 189820
rect 192220 189756 192221 189820
rect 192155 189755 192221 189756
rect 191971 143172 192037 143173
rect 191971 143108 191972 143172
rect 192036 143108 192037 143172
rect 191971 143107 192037 143108
rect 191787 143036 191853 143037
rect 191787 142972 191788 143036
rect 191852 142972 191853 143036
rect 191787 142971 191853 142972
rect 191603 141540 191669 141541
rect 191603 141476 191604 141540
rect 191668 141476 191669 141540
rect 191603 141475 191669 141476
rect 190499 76396 190565 76397
rect 190499 76332 190500 76396
rect 190564 76332 190565 76396
rect 190499 76331 190565 76332
rect 189027 70956 189093 70957
rect 189027 70892 189028 70956
rect 189092 70892 189093 70956
rect 189027 70891 189093 70892
rect 187187 65516 187253 65517
rect 187187 65452 187188 65516
rect 187252 65452 187253 65516
rect 187187 65451 187253 65452
rect 186294 43718 186326 43954
rect 186562 43718 186646 43954
rect 186882 43718 186914 43954
rect 186294 43634 186914 43718
rect 186294 43398 186326 43634
rect 186562 43398 186646 43634
rect 186882 43398 186914 43634
rect 186294 7954 186914 43398
rect 186294 7718 186326 7954
rect 186562 7718 186646 7954
rect 186882 7718 186914 7954
rect 186294 7634 186914 7718
rect 186294 7398 186326 7634
rect 186562 7398 186646 7634
rect 186882 7398 186914 7634
rect 186294 -1306 186914 7398
rect 186294 -1542 186326 -1306
rect 186562 -1542 186646 -1306
rect 186882 -1542 186914 -1306
rect 186294 -1626 186914 -1542
rect 186294 -1862 186326 -1626
rect 186562 -1862 186646 -1626
rect 186882 -1862 186914 -1626
rect 186294 -7654 186914 -1862
rect 190794 48454 191414 78000
rect 191606 71093 191666 141475
rect 191787 140452 191853 140453
rect 191787 140388 191788 140452
rect 191852 140388 191853 140452
rect 191787 140387 191853 140388
rect 191790 81157 191850 140387
rect 191971 138548 192037 138549
rect 191971 138484 191972 138548
rect 192036 138484 192037 138548
rect 191971 138483 192037 138484
rect 191974 81970 192034 138483
rect 192158 82106 192218 189755
rect 192158 82046 192586 82106
rect 191974 81910 192218 81970
rect 191971 81428 192037 81429
rect 191971 81364 191972 81428
rect 192036 81364 192037 81428
rect 191971 81363 192037 81364
rect 191787 81156 191853 81157
rect 191787 81092 191788 81156
rect 191852 81092 191853 81156
rect 191787 81091 191853 81092
rect 191603 71092 191669 71093
rect 191603 71028 191604 71092
rect 191668 71028 191669 71092
rect 191603 71027 191669 71028
rect 191974 64890 192034 81363
rect 192158 80477 192218 81910
rect 192155 80476 192221 80477
rect 192155 80412 192156 80476
rect 192220 80412 192221 80476
rect 192155 80411 192221 80412
rect 192526 80070 192586 82046
rect 192158 80010 192586 80070
rect 192158 75853 192218 80010
rect 192155 75852 192221 75853
rect 192155 75788 192156 75852
rect 192220 75788 192221 75852
rect 192155 75787 192221 75788
rect 193262 73677 193322 191115
rect 194547 191044 194613 191045
rect 194547 190980 194548 191044
rect 194612 190980 194613 191044
rect 194547 190979 194613 190980
rect 193443 137596 193509 137597
rect 193443 137532 193444 137596
rect 193508 137532 193509 137596
rect 193443 137531 193509 137532
rect 193259 73676 193325 73677
rect 193259 73612 193260 73676
rect 193324 73612 193325 73676
rect 193259 73611 193325 73612
rect 193446 67421 193506 137531
rect 194550 74357 194610 190979
rect 195294 160954 195914 196398
rect 196022 194581 196082 196419
rect 196019 194580 196085 194581
rect 196019 194516 196020 194580
rect 196084 194516 196085 194580
rect 196019 194515 196085 194516
rect 196571 194580 196637 194581
rect 196571 194516 196572 194580
rect 196636 194516 196637 194580
rect 196571 194515 196637 194516
rect 195294 160718 195326 160954
rect 195562 160718 195646 160954
rect 195882 160718 195914 160954
rect 195294 160634 195914 160718
rect 195294 160398 195326 160634
rect 195562 160398 195646 160634
rect 195882 160398 195914 160634
rect 195294 124954 195914 160398
rect 196019 145892 196085 145893
rect 196019 145828 196020 145892
rect 196084 145828 196085 145892
rect 196019 145827 196085 145828
rect 195294 124718 195326 124954
rect 195562 124718 195646 124954
rect 195882 124718 195914 124954
rect 195294 124634 195914 124718
rect 195294 124398 195326 124634
rect 195562 124398 195646 124634
rect 195882 124398 195914 124634
rect 195294 88954 195914 124398
rect 195294 88718 195326 88954
rect 195562 88718 195646 88954
rect 195882 88718 195914 88954
rect 195294 88634 195914 88718
rect 195294 88398 195326 88634
rect 195562 88398 195646 88634
rect 195882 88398 195914 88634
rect 194547 74356 194613 74357
rect 194547 74292 194548 74356
rect 194612 74292 194613 74356
rect 194547 74291 194613 74292
rect 193443 67420 193509 67421
rect 193443 67356 193444 67420
rect 193508 67356 193509 67420
rect 193443 67355 193509 67356
rect 190794 48218 190826 48454
rect 191062 48218 191146 48454
rect 191382 48218 191414 48454
rect 190794 48134 191414 48218
rect 190794 47898 190826 48134
rect 191062 47898 191146 48134
rect 191382 47898 191414 48134
rect 190794 12454 191414 47898
rect 191790 64830 192034 64890
rect 191790 34509 191850 64830
rect 195294 52954 195914 88398
rect 196022 68509 196082 145827
rect 196387 140044 196453 140045
rect 196387 139980 196388 140044
rect 196452 139980 196453 140044
rect 196387 139979 196453 139980
rect 196203 139364 196269 139365
rect 196203 139300 196204 139364
rect 196268 139300 196269 139364
rect 196203 139299 196269 139300
rect 196019 68508 196085 68509
rect 196019 68444 196020 68508
rect 196084 68444 196085 68508
rect 196019 68443 196085 68444
rect 196206 64565 196266 139299
rect 196390 72997 196450 139979
rect 196574 73813 196634 194515
rect 198779 191724 198845 191725
rect 198779 191660 198780 191724
rect 198844 191660 198845 191724
rect 198779 191659 198845 191660
rect 197491 191316 197557 191317
rect 197491 191252 197492 191316
rect 197556 191252 197557 191316
rect 197491 191251 197557 191252
rect 197307 190908 197373 190909
rect 197307 190844 197308 190908
rect 197372 190844 197373 190908
rect 197307 190843 197373 190844
rect 196571 73812 196637 73813
rect 196571 73748 196572 73812
rect 196636 73748 196637 73812
rect 196571 73747 196637 73748
rect 196387 72996 196453 72997
rect 196387 72932 196388 72996
rect 196452 72932 196453 72996
rect 196387 72931 196453 72932
rect 197310 72861 197370 190843
rect 197494 74493 197554 191251
rect 198782 190637 198842 191659
rect 198779 190636 198845 190637
rect 198779 190572 198780 190636
rect 198844 190572 198845 190636
rect 198779 190571 198845 190572
rect 197859 146980 197925 146981
rect 197859 146916 197860 146980
rect 197924 146916 197925 146980
rect 197859 146915 197925 146916
rect 197675 146028 197741 146029
rect 197675 145964 197676 146028
rect 197740 145964 197741 146028
rect 197675 145963 197741 145964
rect 197491 74492 197557 74493
rect 197491 74428 197492 74492
rect 197556 74428 197557 74492
rect 197491 74427 197557 74428
rect 197307 72860 197373 72861
rect 197307 72796 197308 72860
rect 197372 72796 197373 72860
rect 197307 72795 197373 72796
rect 197678 68645 197738 145963
rect 197862 104141 197922 146915
rect 197859 104140 197925 104141
rect 197859 104076 197860 104140
rect 197924 104076 197925 104140
rect 197859 104075 197925 104076
rect 198782 72725 198842 190571
rect 199331 187372 199397 187373
rect 199331 187308 199332 187372
rect 199396 187308 199397 187372
rect 199331 187307 199397 187308
rect 198963 184244 199029 184245
rect 198963 184180 198964 184244
rect 199028 184180 199029 184244
rect 198963 184179 199029 184180
rect 198779 72724 198845 72725
rect 198779 72660 198780 72724
rect 198844 72660 198845 72724
rect 198779 72659 198845 72660
rect 197675 68644 197741 68645
rect 197675 68580 197676 68644
rect 197740 68580 197741 68644
rect 197675 68579 197741 68580
rect 198966 68373 199026 184179
rect 199147 139228 199213 139229
rect 199147 139164 199148 139228
rect 199212 139164 199213 139228
rect 199147 139163 199213 139164
rect 199150 81837 199210 139163
rect 199147 81836 199213 81837
rect 199147 81772 199148 81836
rect 199212 81772 199213 81836
rect 199147 81771 199213 81772
rect 199334 72453 199394 187307
rect 199794 165454 200414 200898
rect 204294 709638 204914 711590
rect 204294 709402 204326 709638
rect 204562 709402 204646 709638
rect 204882 709402 204914 709638
rect 204294 709318 204914 709402
rect 204294 709082 204326 709318
rect 204562 709082 204646 709318
rect 204882 709082 204914 709318
rect 204294 673954 204914 709082
rect 204294 673718 204326 673954
rect 204562 673718 204646 673954
rect 204882 673718 204914 673954
rect 204294 673634 204914 673718
rect 204294 673398 204326 673634
rect 204562 673398 204646 673634
rect 204882 673398 204914 673634
rect 204294 637954 204914 673398
rect 204294 637718 204326 637954
rect 204562 637718 204646 637954
rect 204882 637718 204914 637954
rect 204294 637634 204914 637718
rect 204294 637398 204326 637634
rect 204562 637398 204646 637634
rect 204882 637398 204914 637634
rect 204294 601954 204914 637398
rect 204294 601718 204326 601954
rect 204562 601718 204646 601954
rect 204882 601718 204914 601954
rect 204294 601634 204914 601718
rect 204294 601398 204326 601634
rect 204562 601398 204646 601634
rect 204882 601398 204914 601634
rect 204294 565954 204914 601398
rect 204294 565718 204326 565954
rect 204562 565718 204646 565954
rect 204882 565718 204914 565954
rect 204294 565634 204914 565718
rect 204294 565398 204326 565634
rect 204562 565398 204646 565634
rect 204882 565398 204914 565634
rect 204294 529954 204914 565398
rect 204294 529718 204326 529954
rect 204562 529718 204646 529954
rect 204882 529718 204914 529954
rect 204294 529634 204914 529718
rect 204294 529398 204326 529634
rect 204562 529398 204646 529634
rect 204882 529398 204914 529634
rect 204294 493954 204914 529398
rect 204294 493718 204326 493954
rect 204562 493718 204646 493954
rect 204882 493718 204914 493954
rect 204294 493634 204914 493718
rect 204294 493398 204326 493634
rect 204562 493398 204646 493634
rect 204882 493398 204914 493634
rect 204294 457954 204914 493398
rect 204294 457718 204326 457954
rect 204562 457718 204646 457954
rect 204882 457718 204914 457954
rect 204294 457634 204914 457718
rect 204294 457398 204326 457634
rect 204562 457398 204646 457634
rect 204882 457398 204914 457634
rect 204294 421954 204914 457398
rect 204294 421718 204326 421954
rect 204562 421718 204646 421954
rect 204882 421718 204914 421954
rect 204294 421634 204914 421718
rect 204294 421398 204326 421634
rect 204562 421398 204646 421634
rect 204882 421398 204914 421634
rect 204294 385954 204914 421398
rect 204294 385718 204326 385954
rect 204562 385718 204646 385954
rect 204882 385718 204914 385954
rect 204294 385634 204914 385718
rect 204294 385398 204326 385634
rect 204562 385398 204646 385634
rect 204882 385398 204914 385634
rect 204294 349954 204914 385398
rect 204294 349718 204326 349954
rect 204562 349718 204646 349954
rect 204882 349718 204914 349954
rect 204294 349634 204914 349718
rect 204294 349398 204326 349634
rect 204562 349398 204646 349634
rect 204882 349398 204914 349634
rect 204294 313954 204914 349398
rect 204294 313718 204326 313954
rect 204562 313718 204646 313954
rect 204882 313718 204914 313954
rect 204294 313634 204914 313718
rect 204294 313398 204326 313634
rect 204562 313398 204646 313634
rect 204882 313398 204914 313634
rect 204294 277954 204914 313398
rect 204294 277718 204326 277954
rect 204562 277718 204646 277954
rect 204882 277718 204914 277954
rect 204294 277634 204914 277718
rect 204294 277398 204326 277634
rect 204562 277398 204646 277634
rect 204882 277398 204914 277634
rect 204294 241954 204914 277398
rect 204294 241718 204326 241954
rect 204562 241718 204646 241954
rect 204882 241718 204914 241954
rect 204294 241634 204914 241718
rect 204294 241398 204326 241634
rect 204562 241398 204646 241634
rect 204882 241398 204914 241634
rect 204294 205954 204914 241398
rect 204294 205718 204326 205954
rect 204562 205718 204646 205954
rect 204882 205718 204914 205954
rect 204294 205634 204914 205718
rect 204294 205398 204326 205634
rect 204562 205398 204646 205634
rect 204882 205398 204914 205634
rect 203011 200836 203077 200837
rect 203011 200772 203012 200836
rect 203076 200772 203077 200836
rect 203011 200771 203077 200772
rect 203014 200293 203074 200771
rect 203011 200292 203077 200293
rect 203011 200228 203012 200292
rect 203076 200228 203077 200292
rect 203011 200227 203077 200228
rect 200987 192540 201053 192541
rect 200987 192476 200988 192540
rect 201052 192476 201053 192540
rect 200987 192475 201053 192476
rect 200619 180300 200685 180301
rect 200619 180236 200620 180300
rect 200684 180236 200685 180300
rect 200619 180235 200685 180236
rect 199794 165218 199826 165454
rect 200062 165218 200146 165454
rect 200382 165218 200414 165454
rect 199794 165134 200414 165218
rect 199794 164898 199826 165134
rect 200062 164898 200146 165134
rect 200382 164898 200414 165134
rect 199794 129454 200414 164898
rect 199794 129218 199826 129454
rect 200062 129218 200146 129454
rect 200382 129218 200414 129454
rect 199794 129134 200414 129218
rect 199794 128898 199826 129134
rect 200062 128898 200146 129134
rect 200382 128898 200414 129134
rect 199794 93454 200414 128898
rect 199794 93218 199826 93454
rect 200062 93218 200146 93454
rect 200382 93218 200414 93454
rect 199794 93134 200414 93218
rect 199794 92898 199826 93134
rect 200062 92898 200146 93134
rect 200382 92898 200414 93134
rect 199331 72452 199397 72453
rect 199331 72388 199332 72452
rect 199396 72388 199397 72452
rect 199331 72387 199397 72388
rect 198963 68372 199029 68373
rect 198963 68308 198964 68372
rect 199028 68308 199029 68372
rect 198963 68307 199029 68308
rect 196203 64564 196269 64565
rect 196203 64500 196204 64564
rect 196268 64500 196269 64564
rect 196203 64499 196269 64500
rect 195294 52718 195326 52954
rect 195562 52718 195646 52954
rect 195882 52718 195914 52954
rect 195294 52634 195914 52718
rect 195294 52398 195326 52634
rect 195562 52398 195646 52634
rect 195882 52398 195914 52634
rect 191787 34508 191853 34509
rect 191787 34444 191788 34508
rect 191852 34444 191853 34508
rect 191787 34443 191853 34444
rect 190794 12218 190826 12454
rect 191062 12218 191146 12454
rect 191382 12218 191414 12454
rect 190794 12134 191414 12218
rect 190794 11898 190826 12134
rect 191062 11898 191146 12134
rect 191382 11898 191414 12134
rect 190794 -2266 191414 11898
rect 190794 -2502 190826 -2266
rect 191062 -2502 191146 -2266
rect 191382 -2502 191414 -2266
rect 190794 -2586 191414 -2502
rect 190794 -2822 190826 -2586
rect 191062 -2822 191146 -2586
rect 191382 -2822 191414 -2586
rect 190794 -7654 191414 -2822
rect 195294 16954 195914 52398
rect 195294 16718 195326 16954
rect 195562 16718 195646 16954
rect 195882 16718 195914 16954
rect 195294 16634 195914 16718
rect 195294 16398 195326 16634
rect 195562 16398 195646 16634
rect 195882 16398 195914 16634
rect 195294 -3226 195914 16398
rect 195294 -3462 195326 -3226
rect 195562 -3462 195646 -3226
rect 195882 -3462 195914 -3226
rect 195294 -3546 195914 -3462
rect 195294 -3782 195326 -3546
rect 195562 -3782 195646 -3546
rect 195882 -3782 195914 -3546
rect 195294 -7654 195914 -3782
rect 199794 57454 200414 92898
rect 200622 64021 200682 180235
rect 200803 180028 200869 180029
rect 200803 179964 200804 180028
rect 200868 179964 200869 180028
rect 200803 179963 200869 179964
rect 200806 64429 200866 179963
rect 200990 76669 201050 192475
rect 201539 191452 201605 191453
rect 201539 191388 201540 191452
rect 201604 191388 201605 191452
rect 201539 191387 201605 191388
rect 200987 76668 201053 76669
rect 200987 76604 200988 76668
rect 201052 76604 201053 76668
rect 200987 76603 201053 76604
rect 201542 75445 201602 191387
rect 203014 190470 203074 200227
rect 202830 190410 203074 190470
rect 201723 138684 201789 138685
rect 201723 138620 201724 138684
rect 201788 138620 201789 138684
rect 201723 138619 201789 138620
rect 201539 75444 201605 75445
rect 201539 75380 201540 75444
rect 201604 75380 201605 75444
rect 201539 75379 201605 75380
rect 200803 64428 200869 64429
rect 200803 64364 200804 64428
rect 200868 64364 200869 64428
rect 200803 64363 200869 64364
rect 201726 64157 201786 138619
rect 202830 81293 202890 190410
rect 203011 185740 203077 185741
rect 203011 185676 203012 185740
rect 203076 185676 203077 185740
rect 203011 185675 203077 185676
rect 202827 81292 202893 81293
rect 202827 81228 202828 81292
rect 202892 81228 202893 81292
rect 202827 81227 202893 81228
rect 203014 68781 203074 185675
rect 203195 180572 203261 180573
rect 203195 180508 203196 180572
rect 203260 180508 203261 180572
rect 203195 180507 203261 180508
rect 204115 180572 204181 180573
rect 204115 180508 204116 180572
rect 204180 180508 204181 180572
rect 204115 180507 204181 180508
rect 203198 76805 203258 180507
rect 204118 180165 204178 180507
rect 204115 180164 204181 180165
rect 204115 180100 204116 180164
rect 204180 180100 204181 180164
rect 204115 180099 204181 180100
rect 204294 169954 204914 205398
rect 208794 710598 209414 711590
rect 208794 710362 208826 710598
rect 209062 710362 209146 710598
rect 209382 710362 209414 710598
rect 208794 710278 209414 710362
rect 208794 710042 208826 710278
rect 209062 710042 209146 710278
rect 209382 710042 209414 710278
rect 208794 678454 209414 710042
rect 208794 678218 208826 678454
rect 209062 678218 209146 678454
rect 209382 678218 209414 678454
rect 208794 678134 209414 678218
rect 208794 677898 208826 678134
rect 209062 677898 209146 678134
rect 209382 677898 209414 678134
rect 208794 642454 209414 677898
rect 208794 642218 208826 642454
rect 209062 642218 209146 642454
rect 209382 642218 209414 642454
rect 208794 642134 209414 642218
rect 208794 641898 208826 642134
rect 209062 641898 209146 642134
rect 209382 641898 209414 642134
rect 208794 606454 209414 641898
rect 208794 606218 208826 606454
rect 209062 606218 209146 606454
rect 209382 606218 209414 606454
rect 208794 606134 209414 606218
rect 208794 605898 208826 606134
rect 209062 605898 209146 606134
rect 209382 605898 209414 606134
rect 208794 570454 209414 605898
rect 208794 570218 208826 570454
rect 209062 570218 209146 570454
rect 209382 570218 209414 570454
rect 208794 570134 209414 570218
rect 208794 569898 208826 570134
rect 209062 569898 209146 570134
rect 209382 569898 209414 570134
rect 208794 534454 209414 569898
rect 208794 534218 208826 534454
rect 209062 534218 209146 534454
rect 209382 534218 209414 534454
rect 208794 534134 209414 534218
rect 208794 533898 208826 534134
rect 209062 533898 209146 534134
rect 209382 533898 209414 534134
rect 208794 498454 209414 533898
rect 208794 498218 208826 498454
rect 209062 498218 209146 498454
rect 209382 498218 209414 498454
rect 208794 498134 209414 498218
rect 208794 497898 208826 498134
rect 209062 497898 209146 498134
rect 209382 497898 209414 498134
rect 208794 462454 209414 497898
rect 208794 462218 208826 462454
rect 209062 462218 209146 462454
rect 209382 462218 209414 462454
rect 208794 462134 209414 462218
rect 208794 461898 208826 462134
rect 209062 461898 209146 462134
rect 209382 461898 209414 462134
rect 208794 426454 209414 461898
rect 208794 426218 208826 426454
rect 209062 426218 209146 426454
rect 209382 426218 209414 426454
rect 208794 426134 209414 426218
rect 208794 425898 208826 426134
rect 209062 425898 209146 426134
rect 209382 425898 209414 426134
rect 208794 390454 209414 425898
rect 208794 390218 208826 390454
rect 209062 390218 209146 390454
rect 209382 390218 209414 390454
rect 208794 390134 209414 390218
rect 208794 389898 208826 390134
rect 209062 389898 209146 390134
rect 209382 389898 209414 390134
rect 208794 354454 209414 389898
rect 208794 354218 208826 354454
rect 209062 354218 209146 354454
rect 209382 354218 209414 354454
rect 208794 354134 209414 354218
rect 208794 353898 208826 354134
rect 209062 353898 209146 354134
rect 209382 353898 209414 354134
rect 208794 318454 209414 353898
rect 208794 318218 208826 318454
rect 209062 318218 209146 318454
rect 209382 318218 209414 318454
rect 208794 318134 209414 318218
rect 208794 317898 208826 318134
rect 209062 317898 209146 318134
rect 209382 317898 209414 318134
rect 208794 282454 209414 317898
rect 208794 282218 208826 282454
rect 209062 282218 209146 282454
rect 209382 282218 209414 282454
rect 208794 282134 209414 282218
rect 208794 281898 208826 282134
rect 209062 281898 209146 282134
rect 209382 281898 209414 282134
rect 208794 246454 209414 281898
rect 208794 246218 208826 246454
rect 209062 246218 209146 246454
rect 209382 246218 209414 246454
rect 208794 246134 209414 246218
rect 208794 245898 208826 246134
rect 209062 245898 209146 246134
rect 209382 245898 209414 246134
rect 208794 210454 209414 245898
rect 208794 210218 208826 210454
rect 209062 210218 209146 210454
rect 209382 210218 209414 210454
rect 208794 210134 209414 210218
rect 208794 209898 208826 210134
rect 209062 209898 209146 210134
rect 209382 209898 209414 210134
rect 207059 200700 207125 200701
rect 207059 200636 207060 200700
rect 207124 200636 207125 200700
rect 207059 200635 207125 200636
rect 207062 200157 207122 200635
rect 207059 200156 207125 200157
rect 207059 200092 207060 200156
rect 207124 200092 207125 200156
rect 207059 200091 207125 200092
rect 205587 194172 205653 194173
rect 205587 194108 205588 194172
rect 205652 194108 205653 194172
rect 205587 194107 205653 194108
rect 204294 169718 204326 169954
rect 204562 169718 204646 169954
rect 204882 169718 204914 169954
rect 204294 169634 204914 169718
rect 204294 169398 204326 169634
rect 204562 169398 204646 169634
rect 204882 169398 204914 169634
rect 204294 133954 204914 169398
rect 204294 133718 204326 133954
rect 204562 133718 204646 133954
rect 204882 133718 204914 133954
rect 204294 133634 204914 133718
rect 204294 133398 204326 133634
rect 204562 133398 204646 133634
rect 204882 133398 204914 133634
rect 204294 97954 204914 133398
rect 204294 97718 204326 97954
rect 204562 97718 204646 97954
rect 204882 97718 204914 97954
rect 204294 97634 204914 97718
rect 204294 97398 204326 97634
rect 204562 97398 204646 97634
rect 204882 97398 204914 97634
rect 203195 76804 203261 76805
rect 203195 76740 203196 76804
rect 203260 76740 203261 76804
rect 203195 76739 203261 76740
rect 203011 68780 203077 68781
rect 203011 68716 203012 68780
rect 203076 68716 203077 68780
rect 203011 68715 203077 68716
rect 201723 64156 201789 64157
rect 201723 64092 201724 64156
rect 201788 64092 201789 64156
rect 201723 64091 201789 64092
rect 200619 64020 200685 64021
rect 200619 63956 200620 64020
rect 200684 63956 200685 64020
rect 200619 63955 200685 63956
rect 199794 57218 199826 57454
rect 200062 57218 200146 57454
rect 200382 57218 200414 57454
rect 199794 57134 200414 57218
rect 199794 56898 199826 57134
rect 200062 56898 200146 57134
rect 200382 56898 200414 57134
rect 199794 21454 200414 56898
rect 199794 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 200414 21454
rect 199794 21134 200414 21218
rect 199794 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 200414 21134
rect 199794 -4186 200414 20898
rect 199794 -4422 199826 -4186
rect 200062 -4422 200146 -4186
rect 200382 -4422 200414 -4186
rect 199794 -4506 200414 -4422
rect 199794 -4742 199826 -4506
rect 200062 -4742 200146 -4506
rect 200382 -4742 200414 -4506
rect 199794 -7654 200414 -4742
rect 204294 61954 204914 97398
rect 205590 70141 205650 194107
rect 205771 189820 205837 189821
rect 205771 189756 205772 189820
rect 205836 189756 205837 189820
rect 205771 189755 205837 189756
rect 205774 188597 205834 189755
rect 205771 188596 205837 188597
rect 205771 188532 205772 188596
rect 205836 188532 205837 188596
rect 205771 188531 205837 188532
rect 205774 71229 205834 188531
rect 205771 71228 205837 71229
rect 205771 71164 205772 71228
rect 205836 71164 205837 71228
rect 205771 71163 205837 71164
rect 205587 70140 205653 70141
rect 205587 70076 205588 70140
rect 205652 70076 205653 70140
rect 205587 70075 205653 70076
rect 207062 69869 207122 200091
rect 207611 189956 207677 189957
rect 207611 189892 207612 189956
rect 207676 189892 207677 189956
rect 207611 189891 207677 189892
rect 207614 74085 207674 189891
rect 208794 174454 209414 209898
rect 213294 711558 213914 711590
rect 213294 711322 213326 711558
rect 213562 711322 213646 711558
rect 213882 711322 213914 711558
rect 213294 711238 213914 711322
rect 213294 711002 213326 711238
rect 213562 711002 213646 711238
rect 213882 711002 213914 711238
rect 213294 682954 213914 711002
rect 213294 682718 213326 682954
rect 213562 682718 213646 682954
rect 213882 682718 213914 682954
rect 213294 682634 213914 682718
rect 213294 682398 213326 682634
rect 213562 682398 213646 682634
rect 213882 682398 213914 682634
rect 213294 646954 213914 682398
rect 213294 646718 213326 646954
rect 213562 646718 213646 646954
rect 213882 646718 213914 646954
rect 213294 646634 213914 646718
rect 213294 646398 213326 646634
rect 213562 646398 213646 646634
rect 213882 646398 213914 646634
rect 213294 610954 213914 646398
rect 213294 610718 213326 610954
rect 213562 610718 213646 610954
rect 213882 610718 213914 610954
rect 213294 610634 213914 610718
rect 213294 610398 213326 610634
rect 213562 610398 213646 610634
rect 213882 610398 213914 610634
rect 213294 574954 213914 610398
rect 213294 574718 213326 574954
rect 213562 574718 213646 574954
rect 213882 574718 213914 574954
rect 213294 574634 213914 574718
rect 213294 574398 213326 574634
rect 213562 574398 213646 574634
rect 213882 574398 213914 574634
rect 213294 538954 213914 574398
rect 213294 538718 213326 538954
rect 213562 538718 213646 538954
rect 213882 538718 213914 538954
rect 213294 538634 213914 538718
rect 213294 538398 213326 538634
rect 213562 538398 213646 538634
rect 213882 538398 213914 538634
rect 213294 502954 213914 538398
rect 213294 502718 213326 502954
rect 213562 502718 213646 502954
rect 213882 502718 213914 502954
rect 213294 502634 213914 502718
rect 213294 502398 213326 502634
rect 213562 502398 213646 502634
rect 213882 502398 213914 502634
rect 213294 466954 213914 502398
rect 213294 466718 213326 466954
rect 213562 466718 213646 466954
rect 213882 466718 213914 466954
rect 213294 466634 213914 466718
rect 213294 466398 213326 466634
rect 213562 466398 213646 466634
rect 213882 466398 213914 466634
rect 213294 430954 213914 466398
rect 213294 430718 213326 430954
rect 213562 430718 213646 430954
rect 213882 430718 213914 430954
rect 213294 430634 213914 430718
rect 213294 430398 213326 430634
rect 213562 430398 213646 430634
rect 213882 430398 213914 430634
rect 213294 394954 213914 430398
rect 213294 394718 213326 394954
rect 213562 394718 213646 394954
rect 213882 394718 213914 394954
rect 213294 394634 213914 394718
rect 213294 394398 213326 394634
rect 213562 394398 213646 394634
rect 213882 394398 213914 394634
rect 213294 358954 213914 394398
rect 213294 358718 213326 358954
rect 213562 358718 213646 358954
rect 213882 358718 213914 358954
rect 213294 358634 213914 358718
rect 213294 358398 213326 358634
rect 213562 358398 213646 358634
rect 213882 358398 213914 358634
rect 213294 322954 213914 358398
rect 213294 322718 213326 322954
rect 213562 322718 213646 322954
rect 213882 322718 213914 322954
rect 213294 322634 213914 322718
rect 213294 322398 213326 322634
rect 213562 322398 213646 322634
rect 213882 322398 213914 322634
rect 213294 286954 213914 322398
rect 213294 286718 213326 286954
rect 213562 286718 213646 286954
rect 213882 286718 213914 286954
rect 213294 286634 213914 286718
rect 213294 286398 213326 286634
rect 213562 286398 213646 286634
rect 213882 286398 213914 286634
rect 213294 250954 213914 286398
rect 213294 250718 213326 250954
rect 213562 250718 213646 250954
rect 213882 250718 213914 250954
rect 213294 250634 213914 250718
rect 213294 250398 213326 250634
rect 213562 250398 213646 250634
rect 213882 250398 213914 250634
rect 213294 214954 213914 250398
rect 213294 214718 213326 214954
rect 213562 214718 213646 214954
rect 213882 214718 213914 214954
rect 213294 214634 213914 214718
rect 213294 214398 213326 214634
rect 213562 214398 213646 214634
rect 213882 214398 213914 214634
rect 211107 199340 211173 199341
rect 211107 199276 211108 199340
rect 211172 199276 211173 199340
rect 211107 199275 211173 199276
rect 208794 174218 208826 174454
rect 209062 174218 209146 174454
rect 209382 174218 209414 174454
rect 208794 174134 209414 174218
rect 208794 173898 208826 174134
rect 209062 173898 209146 174134
rect 209382 173898 209414 174134
rect 208794 138454 209414 173898
rect 208794 138218 208826 138454
rect 209062 138218 209146 138454
rect 209382 138218 209414 138454
rect 208794 138134 209414 138218
rect 208794 137898 208826 138134
rect 209062 137898 209146 138134
rect 209382 137898 209414 138134
rect 208794 102454 209414 137898
rect 208794 102218 208826 102454
rect 209062 102218 209146 102454
rect 209382 102218 209414 102454
rect 208794 102134 209414 102218
rect 208794 101898 208826 102134
rect 209062 101898 209146 102134
rect 209382 101898 209414 102134
rect 207611 74084 207677 74085
rect 207611 74020 207612 74084
rect 207676 74020 207677 74084
rect 207611 74019 207677 74020
rect 207059 69868 207125 69869
rect 207059 69804 207060 69868
rect 207124 69804 207125 69868
rect 207059 69803 207125 69804
rect 204294 61718 204326 61954
rect 204562 61718 204646 61954
rect 204882 61718 204914 61954
rect 204294 61634 204914 61718
rect 204294 61398 204326 61634
rect 204562 61398 204646 61634
rect 204882 61398 204914 61634
rect 204294 25954 204914 61398
rect 204294 25718 204326 25954
rect 204562 25718 204646 25954
rect 204882 25718 204914 25954
rect 204294 25634 204914 25718
rect 204294 25398 204326 25634
rect 204562 25398 204646 25634
rect 204882 25398 204914 25634
rect 204294 -5146 204914 25398
rect 204294 -5382 204326 -5146
rect 204562 -5382 204646 -5146
rect 204882 -5382 204914 -5146
rect 204294 -5466 204914 -5382
rect 204294 -5702 204326 -5466
rect 204562 -5702 204646 -5466
rect 204882 -5702 204914 -5466
rect 204294 -7654 204914 -5702
rect 208794 66454 209414 101898
rect 211110 78301 211170 199275
rect 213294 178954 213914 214398
rect 213294 178718 213326 178954
rect 213562 178718 213646 178954
rect 213882 178718 213914 178954
rect 213294 178634 213914 178718
rect 213294 178398 213326 178634
rect 213562 178398 213646 178634
rect 213882 178398 213914 178634
rect 213294 142954 213914 178398
rect 213294 142718 213326 142954
rect 213562 142718 213646 142954
rect 213882 142718 213914 142954
rect 213294 142634 213914 142718
rect 213294 142398 213326 142634
rect 213562 142398 213646 142634
rect 213882 142398 213914 142634
rect 213294 106954 213914 142398
rect 213294 106718 213326 106954
rect 213562 106718 213646 106954
rect 213882 106718 213914 106954
rect 213294 106634 213914 106718
rect 213294 106398 213326 106634
rect 213562 106398 213646 106634
rect 213882 106398 213914 106634
rect 211107 78300 211173 78301
rect 211107 78236 211108 78300
rect 211172 78236 211173 78300
rect 211107 78235 211173 78236
rect 208794 66218 208826 66454
rect 209062 66218 209146 66454
rect 209382 66218 209414 66454
rect 208794 66134 209414 66218
rect 208794 65898 208826 66134
rect 209062 65898 209146 66134
rect 209382 65898 209414 66134
rect 208794 30454 209414 65898
rect 208794 30218 208826 30454
rect 209062 30218 209146 30454
rect 209382 30218 209414 30454
rect 208794 30134 209414 30218
rect 208794 29898 208826 30134
rect 209062 29898 209146 30134
rect 209382 29898 209414 30134
rect 208794 -6106 209414 29898
rect 208794 -6342 208826 -6106
rect 209062 -6342 209146 -6106
rect 209382 -6342 209414 -6106
rect 208794 -6426 209414 -6342
rect 208794 -6662 208826 -6426
rect 209062 -6662 209146 -6426
rect 209382 -6662 209414 -6426
rect 208794 -7654 209414 -6662
rect 213294 70954 213914 106398
rect 213294 70718 213326 70954
rect 213562 70718 213646 70954
rect 213882 70718 213914 70954
rect 213294 70634 213914 70718
rect 213294 70398 213326 70634
rect 213562 70398 213646 70634
rect 213882 70398 213914 70634
rect 213294 34954 213914 70398
rect 213294 34718 213326 34954
rect 213562 34718 213646 34954
rect 213882 34718 213914 34954
rect 213294 34634 213914 34718
rect 213294 34398 213326 34634
rect 213562 34398 213646 34634
rect 213882 34398 213914 34634
rect 213294 -7066 213914 34398
rect 213294 -7302 213326 -7066
rect 213562 -7302 213646 -7066
rect 213882 -7302 213914 -7066
rect 213294 -7386 213914 -7302
rect 213294 -7622 213326 -7386
rect 213562 -7622 213646 -7386
rect 213882 -7622 213914 -7386
rect 213294 -7654 213914 -7622
rect 217794 704838 218414 711590
rect 217794 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 218414 704838
rect 217794 704518 218414 704602
rect 217794 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 218414 704518
rect 217794 687454 218414 704282
rect 217794 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 218414 687454
rect 217794 687134 218414 687218
rect 217794 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 218414 687134
rect 217794 651454 218414 686898
rect 217794 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 218414 651454
rect 217794 651134 218414 651218
rect 217794 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 218414 651134
rect 217794 615454 218414 650898
rect 217794 615218 217826 615454
rect 218062 615218 218146 615454
rect 218382 615218 218414 615454
rect 217794 615134 218414 615218
rect 217794 614898 217826 615134
rect 218062 614898 218146 615134
rect 218382 614898 218414 615134
rect 217794 579454 218414 614898
rect 217794 579218 217826 579454
rect 218062 579218 218146 579454
rect 218382 579218 218414 579454
rect 217794 579134 218414 579218
rect 217794 578898 217826 579134
rect 218062 578898 218146 579134
rect 218382 578898 218414 579134
rect 217794 543454 218414 578898
rect 217794 543218 217826 543454
rect 218062 543218 218146 543454
rect 218382 543218 218414 543454
rect 217794 543134 218414 543218
rect 217794 542898 217826 543134
rect 218062 542898 218146 543134
rect 218382 542898 218414 543134
rect 217794 507454 218414 542898
rect 217794 507218 217826 507454
rect 218062 507218 218146 507454
rect 218382 507218 218414 507454
rect 217794 507134 218414 507218
rect 217794 506898 217826 507134
rect 218062 506898 218146 507134
rect 218382 506898 218414 507134
rect 217794 471454 218414 506898
rect 217794 471218 217826 471454
rect 218062 471218 218146 471454
rect 218382 471218 218414 471454
rect 217794 471134 218414 471218
rect 217794 470898 217826 471134
rect 218062 470898 218146 471134
rect 218382 470898 218414 471134
rect 217794 435454 218414 470898
rect 217794 435218 217826 435454
rect 218062 435218 218146 435454
rect 218382 435218 218414 435454
rect 217794 435134 218414 435218
rect 217794 434898 217826 435134
rect 218062 434898 218146 435134
rect 218382 434898 218414 435134
rect 217794 399454 218414 434898
rect 217794 399218 217826 399454
rect 218062 399218 218146 399454
rect 218382 399218 218414 399454
rect 217794 399134 218414 399218
rect 217794 398898 217826 399134
rect 218062 398898 218146 399134
rect 218382 398898 218414 399134
rect 217794 363454 218414 398898
rect 217794 363218 217826 363454
rect 218062 363218 218146 363454
rect 218382 363218 218414 363454
rect 217794 363134 218414 363218
rect 217794 362898 217826 363134
rect 218062 362898 218146 363134
rect 218382 362898 218414 363134
rect 217794 327454 218414 362898
rect 217794 327218 217826 327454
rect 218062 327218 218146 327454
rect 218382 327218 218414 327454
rect 217794 327134 218414 327218
rect 217794 326898 217826 327134
rect 218062 326898 218146 327134
rect 218382 326898 218414 327134
rect 217794 291454 218414 326898
rect 217794 291218 217826 291454
rect 218062 291218 218146 291454
rect 218382 291218 218414 291454
rect 217794 291134 218414 291218
rect 217794 290898 217826 291134
rect 218062 290898 218146 291134
rect 218382 290898 218414 291134
rect 217794 255454 218414 290898
rect 217794 255218 217826 255454
rect 218062 255218 218146 255454
rect 218382 255218 218414 255454
rect 217794 255134 218414 255218
rect 217794 254898 217826 255134
rect 218062 254898 218146 255134
rect 218382 254898 218414 255134
rect 217794 219454 218414 254898
rect 217794 219218 217826 219454
rect 218062 219218 218146 219454
rect 218382 219218 218414 219454
rect 217794 219134 218414 219218
rect 217794 218898 217826 219134
rect 218062 218898 218146 219134
rect 218382 218898 218414 219134
rect 217794 183454 218414 218898
rect 217794 183218 217826 183454
rect 218062 183218 218146 183454
rect 218382 183218 218414 183454
rect 217794 183134 218414 183218
rect 217794 182898 217826 183134
rect 218062 182898 218146 183134
rect 218382 182898 218414 183134
rect 217794 147454 218414 182898
rect 217794 147218 217826 147454
rect 218062 147218 218146 147454
rect 218382 147218 218414 147454
rect 217794 147134 218414 147218
rect 217794 146898 217826 147134
rect 218062 146898 218146 147134
rect 218382 146898 218414 147134
rect 217794 111454 218414 146898
rect 217794 111218 217826 111454
rect 218062 111218 218146 111454
rect 218382 111218 218414 111454
rect 217794 111134 218414 111218
rect 217794 110898 217826 111134
rect 218062 110898 218146 111134
rect 218382 110898 218414 111134
rect 217794 75454 218414 110898
rect 217794 75218 217826 75454
rect 218062 75218 218146 75454
rect 218382 75218 218414 75454
rect 217794 75134 218414 75218
rect 217794 74898 217826 75134
rect 218062 74898 218146 75134
rect 218382 74898 218414 75134
rect 217794 39454 218414 74898
rect 217794 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 218414 39454
rect 217794 39134 218414 39218
rect 217794 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 218414 39134
rect 217794 3454 218414 38898
rect 217794 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 218414 3454
rect 217794 3134 218414 3218
rect 217794 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 218414 3134
rect 217794 -346 218414 2898
rect 217794 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 218414 -346
rect 217794 -666 218414 -582
rect 217794 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 218414 -666
rect 217794 -7654 218414 -902
rect 222294 705798 222914 711590
rect 222294 705562 222326 705798
rect 222562 705562 222646 705798
rect 222882 705562 222914 705798
rect 222294 705478 222914 705562
rect 222294 705242 222326 705478
rect 222562 705242 222646 705478
rect 222882 705242 222914 705478
rect 222294 691954 222914 705242
rect 222294 691718 222326 691954
rect 222562 691718 222646 691954
rect 222882 691718 222914 691954
rect 222294 691634 222914 691718
rect 222294 691398 222326 691634
rect 222562 691398 222646 691634
rect 222882 691398 222914 691634
rect 222294 655954 222914 691398
rect 222294 655718 222326 655954
rect 222562 655718 222646 655954
rect 222882 655718 222914 655954
rect 222294 655634 222914 655718
rect 222294 655398 222326 655634
rect 222562 655398 222646 655634
rect 222882 655398 222914 655634
rect 222294 619954 222914 655398
rect 222294 619718 222326 619954
rect 222562 619718 222646 619954
rect 222882 619718 222914 619954
rect 222294 619634 222914 619718
rect 222294 619398 222326 619634
rect 222562 619398 222646 619634
rect 222882 619398 222914 619634
rect 222294 583954 222914 619398
rect 222294 583718 222326 583954
rect 222562 583718 222646 583954
rect 222882 583718 222914 583954
rect 222294 583634 222914 583718
rect 222294 583398 222326 583634
rect 222562 583398 222646 583634
rect 222882 583398 222914 583634
rect 222294 547954 222914 583398
rect 222294 547718 222326 547954
rect 222562 547718 222646 547954
rect 222882 547718 222914 547954
rect 222294 547634 222914 547718
rect 222294 547398 222326 547634
rect 222562 547398 222646 547634
rect 222882 547398 222914 547634
rect 222294 511954 222914 547398
rect 222294 511718 222326 511954
rect 222562 511718 222646 511954
rect 222882 511718 222914 511954
rect 222294 511634 222914 511718
rect 222294 511398 222326 511634
rect 222562 511398 222646 511634
rect 222882 511398 222914 511634
rect 222294 475954 222914 511398
rect 222294 475718 222326 475954
rect 222562 475718 222646 475954
rect 222882 475718 222914 475954
rect 222294 475634 222914 475718
rect 222294 475398 222326 475634
rect 222562 475398 222646 475634
rect 222882 475398 222914 475634
rect 222294 439954 222914 475398
rect 222294 439718 222326 439954
rect 222562 439718 222646 439954
rect 222882 439718 222914 439954
rect 222294 439634 222914 439718
rect 222294 439398 222326 439634
rect 222562 439398 222646 439634
rect 222882 439398 222914 439634
rect 222294 403954 222914 439398
rect 222294 403718 222326 403954
rect 222562 403718 222646 403954
rect 222882 403718 222914 403954
rect 222294 403634 222914 403718
rect 222294 403398 222326 403634
rect 222562 403398 222646 403634
rect 222882 403398 222914 403634
rect 222294 367954 222914 403398
rect 222294 367718 222326 367954
rect 222562 367718 222646 367954
rect 222882 367718 222914 367954
rect 222294 367634 222914 367718
rect 222294 367398 222326 367634
rect 222562 367398 222646 367634
rect 222882 367398 222914 367634
rect 222294 331954 222914 367398
rect 222294 331718 222326 331954
rect 222562 331718 222646 331954
rect 222882 331718 222914 331954
rect 222294 331634 222914 331718
rect 222294 331398 222326 331634
rect 222562 331398 222646 331634
rect 222882 331398 222914 331634
rect 222294 295954 222914 331398
rect 222294 295718 222326 295954
rect 222562 295718 222646 295954
rect 222882 295718 222914 295954
rect 222294 295634 222914 295718
rect 222294 295398 222326 295634
rect 222562 295398 222646 295634
rect 222882 295398 222914 295634
rect 222294 259954 222914 295398
rect 222294 259718 222326 259954
rect 222562 259718 222646 259954
rect 222882 259718 222914 259954
rect 222294 259634 222914 259718
rect 222294 259398 222326 259634
rect 222562 259398 222646 259634
rect 222882 259398 222914 259634
rect 222294 223954 222914 259398
rect 222294 223718 222326 223954
rect 222562 223718 222646 223954
rect 222882 223718 222914 223954
rect 222294 223634 222914 223718
rect 222294 223398 222326 223634
rect 222562 223398 222646 223634
rect 222882 223398 222914 223634
rect 222294 187954 222914 223398
rect 222294 187718 222326 187954
rect 222562 187718 222646 187954
rect 222882 187718 222914 187954
rect 222294 187634 222914 187718
rect 222294 187398 222326 187634
rect 222562 187398 222646 187634
rect 222882 187398 222914 187634
rect 222294 151954 222914 187398
rect 222294 151718 222326 151954
rect 222562 151718 222646 151954
rect 222882 151718 222914 151954
rect 222294 151634 222914 151718
rect 222294 151398 222326 151634
rect 222562 151398 222646 151634
rect 222882 151398 222914 151634
rect 222294 115954 222914 151398
rect 222294 115718 222326 115954
rect 222562 115718 222646 115954
rect 222882 115718 222914 115954
rect 222294 115634 222914 115718
rect 222294 115398 222326 115634
rect 222562 115398 222646 115634
rect 222882 115398 222914 115634
rect 222294 79954 222914 115398
rect 222294 79718 222326 79954
rect 222562 79718 222646 79954
rect 222882 79718 222914 79954
rect 222294 79634 222914 79718
rect 222294 79398 222326 79634
rect 222562 79398 222646 79634
rect 222882 79398 222914 79634
rect 222294 43954 222914 79398
rect 222294 43718 222326 43954
rect 222562 43718 222646 43954
rect 222882 43718 222914 43954
rect 222294 43634 222914 43718
rect 222294 43398 222326 43634
rect 222562 43398 222646 43634
rect 222882 43398 222914 43634
rect 222294 7954 222914 43398
rect 222294 7718 222326 7954
rect 222562 7718 222646 7954
rect 222882 7718 222914 7954
rect 222294 7634 222914 7718
rect 222294 7398 222326 7634
rect 222562 7398 222646 7634
rect 222882 7398 222914 7634
rect 222294 -1306 222914 7398
rect 222294 -1542 222326 -1306
rect 222562 -1542 222646 -1306
rect 222882 -1542 222914 -1306
rect 222294 -1626 222914 -1542
rect 222294 -1862 222326 -1626
rect 222562 -1862 222646 -1626
rect 222882 -1862 222914 -1626
rect 222294 -7654 222914 -1862
rect 226794 706758 227414 711590
rect 226794 706522 226826 706758
rect 227062 706522 227146 706758
rect 227382 706522 227414 706758
rect 226794 706438 227414 706522
rect 226794 706202 226826 706438
rect 227062 706202 227146 706438
rect 227382 706202 227414 706438
rect 226794 696454 227414 706202
rect 226794 696218 226826 696454
rect 227062 696218 227146 696454
rect 227382 696218 227414 696454
rect 226794 696134 227414 696218
rect 226794 695898 226826 696134
rect 227062 695898 227146 696134
rect 227382 695898 227414 696134
rect 226794 660454 227414 695898
rect 226794 660218 226826 660454
rect 227062 660218 227146 660454
rect 227382 660218 227414 660454
rect 226794 660134 227414 660218
rect 226794 659898 226826 660134
rect 227062 659898 227146 660134
rect 227382 659898 227414 660134
rect 226794 624454 227414 659898
rect 226794 624218 226826 624454
rect 227062 624218 227146 624454
rect 227382 624218 227414 624454
rect 226794 624134 227414 624218
rect 226794 623898 226826 624134
rect 227062 623898 227146 624134
rect 227382 623898 227414 624134
rect 226794 588454 227414 623898
rect 226794 588218 226826 588454
rect 227062 588218 227146 588454
rect 227382 588218 227414 588454
rect 226794 588134 227414 588218
rect 226794 587898 226826 588134
rect 227062 587898 227146 588134
rect 227382 587898 227414 588134
rect 226794 552454 227414 587898
rect 226794 552218 226826 552454
rect 227062 552218 227146 552454
rect 227382 552218 227414 552454
rect 226794 552134 227414 552218
rect 226794 551898 226826 552134
rect 227062 551898 227146 552134
rect 227382 551898 227414 552134
rect 226794 516454 227414 551898
rect 226794 516218 226826 516454
rect 227062 516218 227146 516454
rect 227382 516218 227414 516454
rect 226794 516134 227414 516218
rect 226794 515898 226826 516134
rect 227062 515898 227146 516134
rect 227382 515898 227414 516134
rect 226794 480454 227414 515898
rect 226794 480218 226826 480454
rect 227062 480218 227146 480454
rect 227382 480218 227414 480454
rect 226794 480134 227414 480218
rect 226794 479898 226826 480134
rect 227062 479898 227146 480134
rect 227382 479898 227414 480134
rect 226794 444454 227414 479898
rect 226794 444218 226826 444454
rect 227062 444218 227146 444454
rect 227382 444218 227414 444454
rect 226794 444134 227414 444218
rect 226794 443898 226826 444134
rect 227062 443898 227146 444134
rect 227382 443898 227414 444134
rect 226794 408454 227414 443898
rect 226794 408218 226826 408454
rect 227062 408218 227146 408454
rect 227382 408218 227414 408454
rect 226794 408134 227414 408218
rect 226794 407898 226826 408134
rect 227062 407898 227146 408134
rect 227382 407898 227414 408134
rect 226794 372454 227414 407898
rect 226794 372218 226826 372454
rect 227062 372218 227146 372454
rect 227382 372218 227414 372454
rect 226794 372134 227414 372218
rect 226794 371898 226826 372134
rect 227062 371898 227146 372134
rect 227382 371898 227414 372134
rect 226794 336454 227414 371898
rect 226794 336218 226826 336454
rect 227062 336218 227146 336454
rect 227382 336218 227414 336454
rect 226794 336134 227414 336218
rect 226794 335898 226826 336134
rect 227062 335898 227146 336134
rect 227382 335898 227414 336134
rect 226794 300454 227414 335898
rect 226794 300218 226826 300454
rect 227062 300218 227146 300454
rect 227382 300218 227414 300454
rect 226794 300134 227414 300218
rect 226794 299898 226826 300134
rect 227062 299898 227146 300134
rect 227382 299898 227414 300134
rect 226794 264454 227414 299898
rect 226794 264218 226826 264454
rect 227062 264218 227146 264454
rect 227382 264218 227414 264454
rect 226794 264134 227414 264218
rect 226794 263898 226826 264134
rect 227062 263898 227146 264134
rect 227382 263898 227414 264134
rect 226794 228454 227414 263898
rect 226794 228218 226826 228454
rect 227062 228218 227146 228454
rect 227382 228218 227414 228454
rect 226794 228134 227414 228218
rect 226794 227898 226826 228134
rect 227062 227898 227146 228134
rect 227382 227898 227414 228134
rect 226794 192454 227414 227898
rect 226794 192218 226826 192454
rect 227062 192218 227146 192454
rect 227382 192218 227414 192454
rect 226794 192134 227414 192218
rect 226794 191898 226826 192134
rect 227062 191898 227146 192134
rect 227382 191898 227414 192134
rect 226794 156454 227414 191898
rect 226794 156218 226826 156454
rect 227062 156218 227146 156454
rect 227382 156218 227414 156454
rect 226794 156134 227414 156218
rect 226794 155898 226826 156134
rect 227062 155898 227146 156134
rect 227382 155898 227414 156134
rect 226794 120454 227414 155898
rect 226794 120218 226826 120454
rect 227062 120218 227146 120454
rect 227382 120218 227414 120454
rect 226794 120134 227414 120218
rect 226794 119898 226826 120134
rect 227062 119898 227146 120134
rect 227382 119898 227414 120134
rect 226794 84454 227414 119898
rect 226794 84218 226826 84454
rect 227062 84218 227146 84454
rect 227382 84218 227414 84454
rect 226794 84134 227414 84218
rect 226794 83898 226826 84134
rect 227062 83898 227146 84134
rect 227382 83898 227414 84134
rect 226794 48454 227414 83898
rect 226794 48218 226826 48454
rect 227062 48218 227146 48454
rect 227382 48218 227414 48454
rect 226794 48134 227414 48218
rect 226794 47898 226826 48134
rect 227062 47898 227146 48134
rect 227382 47898 227414 48134
rect 226794 12454 227414 47898
rect 226794 12218 226826 12454
rect 227062 12218 227146 12454
rect 227382 12218 227414 12454
rect 226794 12134 227414 12218
rect 226794 11898 226826 12134
rect 227062 11898 227146 12134
rect 227382 11898 227414 12134
rect 226794 -2266 227414 11898
rect 226794 -2502 226826 -2266
rect 227062 -2502 227146 -2266
rect 227382 -2502 227414 -2266
rect 226794 -2586 227414 -2502
rect 226794 -2822 226826 -2586
rect 227062 -2822 227146 -2586
rect 227382 -2822 227414 -2586
rect 226794 -7654 227414 -2822
rect 231294 707718 231914 711590
rect 231294 707482 231326 707718
rect 231562 707482 231646 707718
rect 231882 707482 231914 707718
rect 231294 707398 231914 707482
rect 231294 707162 231326 707398
rect 231562 707162 231646 707398
rect 231882 707162 231914 707398
rect 231294 700954 231914 707162
rect 231294 700718 231326 700954
rect 231562 700718 231646 700954
rect 231882 700718 231914 700954
rect 231294 700634 231914 700718
rect 231294 700398 231326 700634
rect 231562 700398 231646 700634
rect 231882 700398 231914 700634
rect 231294 664954 231914 700398
rect 231294 664718 231326 664954
rect 231562 664718 231646 664954
rect 231882 664718 231914 664954
rect 231294 664634 231914 664718
rect 231294 664398 231326 664634
rect 231562 664398 231646 664634
rect 231882 664398 231914 664634
rect 231294 628954 231914 664398
rect 231294 628718 231326 628954
rect 231562 628718 231646 628954
rect 231882 628718 231914 628954
rect 231294 628634 231914 628718
rect 231294 628398 231326 628634
rect 231562 628398 231646 628634
rect 231882 628398 231914 628634
rect 231294 592954 231914 628398
rect 231294 592718 231326 592954
rect 231562 592718 231646 592954
rect 231882 592718 231914 592954
rect 231294 592634 231914 592718
rect 231294 592398 231326 592634
rect 231562 592398 231646 592634
rect 231882 592398 231914 592634
rect 231294 556954 231914 592398
rect 231294 556718 231326 556954
rect 231562 556718 231646 556954
rect 231882 556718 231914 556954
rect 231294 556634 231914 556718
rect 231294 556398 231326 556634
rect 231562 556398 231646 556634
rect 231882 556398 231914 556634
rect 231294 520954 231914 556398
rect 231294 520718 231326 520954
rect 231562 520718 231646 520954
rect 231882 520718 231914 520954
rect 231294 520634 231914 520718
rect 231294 520398 231326 520634
rect 231562 520398 231646 520634
rect 231882 520398 231914 520634
rect 231294 484954 231914 520398
rect 231294 484718 231326 484954
rect 231562 484718 231646 484954
rect 231882 484718 231914 484954
rect 231294 484634 231914 484718
rect 231294 484398 231326 484634
rect 231562 484398 231646 484634
rect 231882 484398 231914 484634
rect 231294 448954 231914 484398
rect 231294 448718 231326 448954
rect 231562 448718 231646 448954
rect 231882 448718 231914 448954
rect 231294 448634 231914 448718
rect 231294 448398 231326 448634
rect 231562 448398 231646 448634
rect 231882 448398 231914 448634
rect 231294 412954 231914 448398
rect 231294 412718 231326 412954
rect 231562 412718 231646 412954
rect 231882 412718 231914 412954
rect 231294 412634 231914 412718
rect 231294 412398 231326 412634
rect 231562 412398 231646 412634
rect 231882 412398 231914 412634
rect 231294 376954 231914 412398
rect 231294 376718 231326 376954
rect 231562 376718 231646 376954
rect 231882 376718 231914 376954
rect 231294 376634 231914 376718
rect 231294 376398 231326 376634
rect 231562 376398 231646 376634
rect 231882 376398 231914 376634
rect 231294 340954 231914 376398
rect 231294 340718 231326 340954
rect 231562 340718 231646 340954
rect 231882 340718 231914 340954
rect 231294 340634 231914 340718
rect 231294 340398 231326 340634
rect 231562 340398 231646 340634
rect 231882 340398 231914 340634
rect 231294 304954 231914 340398
rect 231294 304718 231326 304954
rect 231562 304718 231646 304954
rect 231882 304718 231914 304954
rect 231294 304634 231914 304718
rect 231294 304398 231326 304634
rect 231562 304398 231646 304634
rect 231882 304398 231914 304634
rect 231294 268954 231914 304398
rect 231294 268718 231326 268954
rect 231562 268718 231646 268954
rect 231882 268718 231914 268954
rect 231294 268634 231914 268718
rect 231294 268398 231326 268634
rect 231562 268398 231646 268634
rect 231882 268398 231914 268634
rect 231294 232954 231914 268398
rect 231294 232718 231326 232954
rect 231562 232718 231646 232954
rect 231882 232718 231914 232954
rect 231294 232634 231914 232718
rect 231294 232398 231326 232634
rect 231562 232398 231646 232634
rect 231882 232398 231914 232634
rect 231294 196954 231914 232398
rect 231294 196718 231326 196954
rect 231562 196718 231646 196954
rect 231882 196718 231914 196954
rect 231294 196634 231914 196718
rect 231294 196398 231326 196634
rect 231562 196398 231646 196634
rect 231882 196398 231914 196634
rect 231294 160954 231914 196398
rect 231294 160718 231326 160954
rect 231562 160718 231646 160954
rect 231882 160718 231914 160954
rect 231294 160634 231914 160718
rect 231294 160398 231326 160634
rect 231562 160398 231646 160634
rect 231882 160398 231914 160634
rect 231294 124954 231914 160398
rect 231294 124718 231326 124954
rect 231562 124718 231646 124954
rect 231882 124718 231914 124954
rect 231294 124634 231914 124718
rect 231294 124398 231326 124634
rect 231562 124398 231646 124634
rect 231882 124398 231914 124634
rect 231294 88954 231914 124398
rect 231294 88718 231326 88954
rect 231562 88718 231646 88954
rect 231882 88718 231914 88954
rect 231294 88634 231914 88718
rect 231294 88398 231326 88634
rect 231562 88398 231646 88634
rect 231882 88398 231914 88634
rect 231294 52954 231914 88398
rect 231294 52718 231326 52954
rect 231562 52718 231646 52954
rect 231882 52718 231914 52954
rect 231294 52634 231914 52718
rect 231294 52398 231326 52634
rect 231562 52398 231646 52634
rect 231882 52398 231914 52634
rect 231294 16954 231914 52398
rect 231294 16718 231326 16954
rect 231562 16718 231646 16954
rect 231882 16718 231914 16954
rect 231294 16634 231914 16718
rect 231294 16398 231326 16634
rect 231562 16398 231646 16634
rect 231882 16398 231914 16634
rect 231294 -3226 231914 16398
rect 231294 -3462 231326 -3226
rect 231562 -3462 231646 -3226
rect 231882 -3462 231914 -3226
rect 231294 -3546 231914 -3462
rect 231294 -3782 231326 -3546
rect 231562 -3782 231646 -3546
rect 231882 -3782 231914 -3546
rect 231294 -7654 231914 -3782
rect 235794 708678 236414 711590
rect 235794 708442 235826 708678
rect 236062 708442 236146 708678
rect 236382 708442 236414 708678
rect 235794 708358 236414 708442
rect 235794 708122 235826 708358
rect 236062 708122 236146 708358
rect 236382 708122 236414 708358
rect 235794 669454 236414 708122
rect 235794 669218 235826 669454
rect 236062 669218 236146 669454
rect 236382 669218 236414 669454
rect 235794 669134 236414 669218
rect 235794 668898 235826 669134
rect 236062 668898 236146 669134
rect 236382 668898 236414 669134
rect 235794 633454 236414 668898
rect 235794 633218 235826 633454
rect 236062 633218 236146 633454
rect 236382 633218 236414 633454
rect 235794 633134 236414 633218
rect 235794 632898 235826 633134
rect 236062 632898 236146 633134
rect 236382 632898 236414 633134
rect 235794 597454 236414 632898
rect 235794 597218 235826 597454
rect 236062 597218 236146 597454
rect 236382 597218 236414 597454
rect 235794 597134 236414 597218
rect 235794 596898 235826 597134
rect 236062 596898 236146 597134
rect 236382 596898 236414 597134
rect 235794 561454 236414 596898
rect 235794 561218 235826 561454
rect 236062 561218 236146 561454
rect 236382 561218 236414 561454
rect 235794 561134 236414 561218
rect 235794 560898 235826 561134
rect 236062 560898 236146 561134
rect 236382 560898 236414 561134
rect 235794 525454 236414 560898
rect 235794 525218 235826 525454
rect 236062 525218 236146 525454
rect 236382 525218 236414 525454
rect 235794 525134 236414 525218
rect 235794 524898 235826 525134
rect 236062 524898 236146 525134
rect 236382 524898 236414 525134
rect 235794 489454 236414 524898
rect 235794 489218 235826 489454
rect 236062 489218 236146 489454
rect 236382 489218 236414 489454
rect 235794 489134 236414 489218
rect 235794 488898 235826 489134
rect 236062 488898 236146 489134
rect 236382 488898 236414 489134
rect 235794 453454 236414 488898
rect 235794 453218 235826 453454
rect 236062 453218 236146 453454
rect 236382 453218 236414 453454
rect 235794 453134 236414 453218
rect 235794 452898 235826 453134
rect 236062 452898 236146 453134
rect 236382 452898 236414 453134
rect 235794 417454 236414 452898
rect 235794 417218 235826 417454
rect 236062 417218 236146 417454
rect 236382 417218 236414 417454
rect 235794 417134 236414 417218
rect 235794 416898 235826 417134
rect 236062 416898 236146 417134
rect 236382 416898 236414 417134
rect 235794 381454 236414 416898
rect 235794 381218 235826 381454
rect 236062 381218 236146 381454
rect 236382 381218 236414 381454
rect 235794 381134 236414 381218
rect 235794 380898 235826 381134
rect 236062 380898 236146 381134
rect 236382 380898 236414 381134
rect 235794 345454 236414 380898
rect 235794 345218 235826 345454
rect 236062 345218 236146 345454
rect 236382 345218 236414 345454
rect 235794 345134 236414 345218
rect 235794 344898 235826 345134
rect 236062 344898 236146 345134
rect 236382 344898 236414 345134
rect 235794 309454 236414 344898
rect 235794 309218 235826 309454
rect 236062 309218 236146 309454
rect 236382 309218 236414 309454
rect 235794 309134 236414 309218
rect 235794 308898 235826 309134
rect 236062 308898 236146 309134
rect 236382 308898 236414 309134
rect 235794 273454 236414 308898
rect 235794 273218 235826 273454
rect 236062 273218 236146 273454
rect 236382 273218 236414 273454
rect 235794 273134 236414 273218
rect 235794 272898 235826 273134
rect 236062 272898 236146 273134
rect 236382 272898 236414 273134
rect 235794 237454 236414 272898
rect 235794 237218 235826 237454
rect 236062 237218 236146 237454
rect 236382 237218 236414 237454
rect 235794 237134 236414 237218
rect 235794 236898 235826 237134
rect 236062 236898 236146 237134
rect 236382 236898 236414 237134
rect 235794 201454 236414 236898
rect 235794 201218 235826 201454
rect 236062 201218 236146 201454
rect 236382 201218 236414 201454
rect 235794 201134 236414 201218
rect 235794 200898 235826 201134
rect 236062 200898 236146 201134
rect 236382 200898 236414 201134
rect 235794 165454 236414 200898
rect 235794 165218 235826 165454
rect 236062 165218 236146 165454
rect 236382 165218 236414 165454
rect 235794 165134 236414 165218
rect 235794 164898 235826 165134
rect 236062 164898 236146 165134
rect 236382 164898 236414 165134
rect 235794 129454 236414 164898
rect 235794 129218 235826 129454
rect 236062 129218 236146 129454
rect 236382 129218 236414 129454
rect 235794 129134 236414 129218
rect 235794 128898 235826 129134
rect 236062 128898 236146 129134
rect 236382 128898 236414 129134
rect 235794 93454 236414 128898
rect 235794 93218 235826 93454
rect 236062 93218 236146 93454
rect 236382 93218 236414 93454
rect 235794 93134 236414 93218
rect 235794 92898 235826 93134
rect 236062 92898 236146 93134
rect 236382 92898 236414 93134
rect 235794 57454 236414 92898
rect 235794 57218 235826 57454
rect 236062 57218 236146 57454
rect 236382 57218 236414 57454
rect 235794 57134 236414 57218
rect 235794 56898 235826 57134
rect 236062 56898 236146 57134
rect 236382 56898 236414 57134
rect 235794 21454 236414 56898
rect 235794 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 236414 21454
rect 235794 21134 236414 21218
rect 235794 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 236414 21134
rect 235794 -4186 236414 20898
rect 235794 -4422 235826 -4186
rect 236062 -4422 236146 -4186
rect 236382 -4422 236414 -4186
rect 235794 -4506 236414 -4422
rect 235794 -4742 235826 -4506
rect 236062 -4742 236146 -4506
rect 236382 -4742 236414 -4506
rect 235794 -7654 236414 -4742
rect 240294 709638 240914 711590
rect 240294 709402 240326 709638
rect 240562 709402 240646 709638
rect 240882 709402 240914 709638
rect 240294 709318 240914 709402
rect 240294 709082 240326 709318
rect 240562 709082 240646 709318
rect 240882 709082 240914 709318
rect 240294 673954 240914 709082
rect 240294 673718 240326 673954
rect 240562 673718 240646 673954
rect 240882 673718 240914 673954
rect 240294 673634 240914 673718
rect 240294 673398 240326 673634
rect 240562 673398 240646 673634
rect 240882 673398 240914 673634
rect 240294 637954 240914 673398
rect 240294 637718 240326 637954
rect 240562 637718 240646 637954
rect 240882 637718 240914 637954
rect 240294 637634 240914 637718
rect 240294 637398 240326 637634
rect 240562 637398 240646 637634
rect 240882 637398 240914 637634
rect 240294 601954 240914 637398
rect 240294 601718 240326 601954
rect 240562 601718 240646 601954
rect 240882 601718 240914 601954
rect 240294 601634 240914 601718
rect 240294 601398 240326 601634
rect 240562 601398 240646 601634
rect 240882 601398 240914 601634
rect 240294 565954 240914 601398
rect 240294 565718 240326 565954
rect 240562 565718 240646 565954
rect 240882 565718 240914 565954
rect 240294 565634 240914 565718
rect 240294 565398 240326 565634
rect 240562 565398 240646 565634
rect 240882 565398 240914 565634
rect 240294 529954 240914 565398
rect 240294 529718 240326 529954
rect 240562 529718 240646 529954
rect 240882 529718 240914 529954
rect 240294 529634 240914 529718
rect 240294 529398 240326 529634
rect 240562 529398 240646 529634
rect 240882 529398 240914 529634
rect 240294 493954 240914 529398
rect 240294 493718 240326 493954
rect 240562 493718 240646 493954
rect 240882 493718 240914 493954
rect 240294 493634 240914 493718
rect 240294 493398 240326 493634
rect 240562 493398 240646 493634
rect 240882 493398 240914 493634
rect 240294 457954 240914 493398
rect 240294 457718 240326 457954
rect 240562 457718 240646 457954
rect 240882 457718 240914 457954
rect 240294 457634 240914 457718
rect 240294 457398 240326 457634
rect 240562 457398 240646 457634
rect 240882 457398 240914 457634
rect 240294 421954 240914 457398
rect 240294 421718 240326 421954
rect 240562 421718 240646 421954
rect 240882 421718 240914 421954
rect 240294 421634 240914 421718
rect 240294 421398 240326 421634
rect 240562 421398 240646 421634
rect 240882 421398 240914 421634
rect 240294 385954 240914 421398
rect 240294 385718 240326 385954
rect 240562 385718 240646 385954
rect 240882 385718 240914 385954
rect 240294 385634 240914 385718
rect 240294 385398 240326 385634
rect 240562 385398 240646 385634
rect 240882 385398 240914 385634
rect 240294 349954 240914 385398
rect 240294 349718 240326 349954
rect 240562 349718 240646 349954
rect 240882 349718 240914 349954
rect 240294 349634 240914 349718
rect 240294 349398 240326 349634
rect 240562 349398 240646 349634
rect 240882 349398 240914 349634
rect 240294 313954 240914 349398
rect 240294 313718 240326 313954
rect 240562 313718 240646 313954
rect 240882 313718 240914 313954
rect 240294 313634 240914 313718
rect 240294 313398 240326 313634
rect 240562 313398 240646 313634
rect 240882 313398 240914 313634
rect 240294 277954 240914 313398
rect 240294 277718 240326 277954
rect 240562 277718 240646 277954
rect 240882 277718 240914 277954
rect 240294 277634 240914 277718
rect 240294 277398 240326 277634
rect 240562 277398 240646 277634
rect 240882 277398 240914 277634
rect 240294 241954 240914 277398
rect 240294 241718 240326 241954
rect 240562 241718 240646 241954
rect 240882 241718 240914 241954
rect 240294 241634 240914 241718
rect 240294 241398 240326 241634
rect 240562 241398 240646 241634
rect 240882 241398 240914 241634
rect 240294 205954 240914 241398
rect 240294 205718 240326 205954
rect 240562 205718 240646 205954
rect 240882 205718 240914 205954
rect 240294 205634 240914 205718
rect 240294 205398 240326 205634
rect 240562 205398 240646 205634
rect 240882 205398 240914 205634
rect 240294 169954 240914 205398
rect 240294 169718 240326 169954
rect 240562 169718 240646 169954
rect 240882 169718 240914 169954
rect 240294 169634 240914 169718
rect 240294 169398 240326 169634
rect 240562 169398 240646 169634
rect 240882 169398 240914 169634
rect 240294 133954 240914 169398
rect 240294 133718 240326 133954
rect 240562 133718 240646 133954
rect 240882 133718 240914 133954
rect 240294 133634 240914 133718
rect 240294 133398 240326 133634
rect 240562 133398 240646 133634
rect 240882 133398 240914 133634
rect 240294 97954 240914 133398
rect 240294 97718 240326 97954
rect 240562 97718 240646 97954
rect 240882 97718 240914 97954
rect 240294 97634 240914 97718
rect 240294 97398 240326 97634
rect 240562 97398 240646 97634
rect 240882 97398 240914 97634
rect 240294 61954 240914 97398
rect 240294 61718 240326 61954
rect 240562 61718 240646 61954
rect 240882 61718 240914 61954
rect 240294 61634 240914 61718
rect 240294 61398 240326 61634
rect 240562 61398 240646 61634
rect 240882 61398 240914 61634
rect 240294 25954 240914 61398
rect 240294 25718 240326 25954
rect 240562 25718 240646 25954
rect 240882 25718 240914 25954
rect 240294 25634 240914 25718
rect 240294 25398 240326 25634
rect 240562 25398 240646 25634
rect 240882 25398 240914 25634
rect 240294 -5146 240914 25398
rect 240294 -5382 240326 -5146
rect 240562 -5382 240646 -5146
rect 240882 -5382 240914 -5146
rect 240294 -5466 240914 -5382
rect 240294 -5702 240326 -5466
rect 240562 -5702 240646 -5466
rect 240882 -5702 240914 -5466
rect 240294 -7654 240914 -5702
rect 244794 710598 245414 711590
rect 244794 710362 244826 710598
rect 245062 710362 245146 710598
rect 245382 710362 245414 710598
rect 244794 710278 245414 710362
rect 244794 710042 244826 710278
rect 245062 710042 245146 710278
rect 245382 710042 245414 710278
rect 244794 678454 245414 710042
rect 244794 678218 244826 678454
rect 245062 678218 245146 678454
rect 245382 678218 245414 678454
rect 244794 678134 245414 678218
rect 244794 677898 244826 678134
rect 245062 677898 245146 678134
rect 245382 677898 245414 678134
rect 244794 642454 245414 677898
rect 244794 642218 244826 642454
rect 245062 642218 245146 642454
rect 245382 642218 245414 642454
rect 244794 642134 245414 642218
rect 244794 641898 244826 642134
rect 245062 641898 245146 642134
rect 245382 641898 245414 642134
rect 244794 606454 245414 641898
rect 244794 606218 244826 606454
rect 245062 606218 245146 606454
rect 245382 606218 245414 606454
rect 244794 606134 245414 606218
rect 244794 605898 244826 606134
rect 245062 605898 245146 606134
rect 245382 605898 245414 606134
rect 244794 570454 245414 605898
rect 244794 570218 244826 570454
rect 245062 570218 245146 570454
rect 245382 570218 245414 570454
rect 244794 570134 245414 570218
rect 244794 569898 244826 570134
rect 245062 569898 245146 570134
rect 245382 569898 245414 570134
rect 244794 534454 245414 569898
rect 244794 534218 244826 534454
rect 245062 534218 245146 534454
rect 245382 534218 245414 534454
rect 244794 534134 245414 534218
rect 244794 533898 244826 534134
rect 245062 533898 245146 534134
rect 245382 533898 245414 534134
rect 244794 498454 245414 533898
rect 244794 498218 244826 498454
rect 245062 498218 245146 498454
rect 245382 498218 245414 498454
rect 244794 498134 245414 498218
rect 244794 497898 244826 498134
rect 245062 497898 245146 498134
rect 245382 497898 245414 498134
rect 244794 462454 245414 497898
rect 244794 462218 244826 462454
rect 245062 462218 245146 462454
rect 245382 462218 245414 462454
rect 244794 462134 245414 462218
rect 244794 461898 244826 462134
rect 245062 461898 245146 462134
rect 245382 461898 245414 462134
rect 244794 426454 245414 461898
rect 244794 426218 244826 426454
rect 245062 426218 245146 426454
rect 245382 426218 245414 426454
rect 244794 426134 245414 426218
rect 244794 425898 244826 426134
rect 245062 425898 245146 426134
rect 245382 425898 245414 426134
rect 244794 390454 245414 425898
rect 244794 390218 244826 390454
rect 245062 390218 245146 390454
rect 245382 390218 245414 390454
rect 244794 390134 245414 390218
rect 244794 389898 244826 390134
rect 245062 389898 245146 390134
rect 245382 389898 245414 390134
rect 244794 354454 245414 389898
rect 244794 354218 244826 354454
rect 245062 354218 245146 354454
rect 245382 354218 245414 354454
rect 244794 354134 245414 354218
rect 244794 353898 244826 354134
rect 245062 353898 245146 354134
rect 245382 353898 245414 354134
rect 244794 318454 245414 353898
rect 244794 318218 244826 318454
rect 245062 318218 245146 318454
rect 245382 318218 245414 318454
rect 244794 318134 245414 318218
rect 244794 317898 244826 318134
rect 245062 317898 245146 318134
rect 245382 317898 245414 318134
rect 244794 282454 245414 317898
rect 244794 282218 244826 282454
rect 245062 282218 245146 282454
rect 245382 282218 245414 282454
rect 244794 282134 245414 282218
rect 244794 281898 244826 282134
rect 245062 281898 245146 282134
rect 245382 281898 245414 282134
rect 244794 246454 245414 281898
rect 244794 246218 244826 246454
rect 245062 246218 245146 246454
rect 245382 246218 245414 246454
rect 244794 246134 245414 246218
rect 244794 245898 244826 246134
rect 245062 245898 245146 246134
rect 245382 245898 245414 246134
rect 244794 210454 245414 245898
rect 244794 210218 244826 210454
rect 245062 210218 245146 210454
rect 245382 210218 245414 210454
rect 244794 210134 245414 210218
rect 244794 209898 244826 210134
rect 245062 209898 245146 210134
rect 245382 209898 245414 210134
rect 244794 174454 245414 209898
rect 244794 174218 244826 174454
rect 245062 174218 245146 174454
rect 245382 174218 245414 174454
rect 244794 174134 245414 174218
rect 244794 173898 244826 174134
rect 245062 173898 245146 174134
rect 245382 173898 245414 174134
rect 244794 138454 245414 173898
rect 244794 138218 244826 138454
rect 245062 138218 245146 138454
rect 245382 138218 245414 138454
rect 244794 138134 245414 138218
rect 244794 137898 244826 138134
rect 245062 137898 245146 138134
rect 245382 137898 245414 138134
rect 244794 102454 245414 137898
rect 244794 102218 244826 102454
rect 245062 102218 245146 102454
rect 245382 102218 245414 102454
rect 244794 102134 245414 102218
rect 244794 101898 244826 102134
rect 245062 101898 245146 102134
rect 245382 101898 245414 102134
rect 244794 66454 245414 101898
rect 244794 66218 244826 66454
rect 245062 66218 245146 66454
rect 245382 66218 245414 66454
rect 244794 66134 245414 66218
rect 244794 65898 244826 66134
rect 245062 65898 245146 66134
rect 245382 65898 245414 66134
rect 244794 30454 245414 65898
rect 244794 30218 244826 30454
rect 245062 30218 245146 30454
rect 245382 30218 245414 30454
rect 244794 30134 245414 30218
rect 244794 29898 244826 30134
rect 245062 29898 245146 30134
rect 245382 29898 245414 30134
rect 244794 -6106 245414 29898
rect 244794 -6342 244826 -6106
rect 245062 -6342 245146 -6106
rect 245382 -6342 245414 -6106
rect 244794 -6426 245414 -6342
rect 244794 -6662 244826 -6426
rect 245062 -6662 245146 -6426
rect 245382 -6662 245414 -6426
rect 244794 -7654 245414 -6662
rect 249294 711558 249914 711590
rect 249294 711322 249326 711558
rect 249562 711322 249646 711558
rect 249882 711322 249914 711558
rect 249294 711238 249914 711322
rect 249294 711002 249326 711238
rect 249562 711002 249646 711238
rect 249882 711002 249914 711238
rect 249294 682954 249914 711002
rect 249294 682718 249326 682954
rect 249562 682718 249646 682954
rect 249882 682718 249914 682954
rect 249294 682634 249914 682718
rect 249294 682398 249326 682634
rect 249562 682398 249646 682634
rect 249882 682398 249914 682634
rect 249294 646954 249914 682398
rect 249294 646718 249326 646954
rect 249562 646718 249646 646954
rect 249882 646718 249914 646954
rect 249294 646634 249914 646718
rect 249294 646398 249326 646634
rect 249562 646398 249646 646634
rect 249882 646398 249914 646634
rect 249294 610954 249914 646398
rect 249294 610718 249326 610954
rect 249562 610718 249646 610954
rect 249882 610718 249914 610954
rect 249294 610634 249914 610718
rect 249294 610398 249326 610634
rect 249562 610398 249646 610634
rect 249882 610398 249914 610634
rect 249294 574954 249914 610398
rect 249294 574718 249326 574954
rect 249562 574718 249646 574954
rect 249882 574718 249914 574954
rect 249294 574634 249914 574718
rect 249294 574398 249326 574634
rect 249562 574398 249646 574634
rect 249882 574398 249914 574634
rect 249294 538954 249914 574398
rect 249294 538718 249326 538954
rect 249562 538718 249646 538954
rect 249882 538718 249914 538954
rect 249294 538634 249914 538718
rect 249294 538398 249326 538634
rect 249562 538398 249646 538634
rect 249882 538398 249914 538634
rect 249294 502954 249914 538398
rect 249294 502718 249326 502954
rect 249562 502718 249646 502954
rect 249882 502718 249914 502954
rect 249294 502634 249914 502718
rect 249294 502398 249326 502634
rect 249562 502398 249646 502634
rect 249882 502398 249914 502634
rect 249294 466954 249914 502398
rect 249294 466718 249326 466954
rect 249562 466718 249646 466954
rect 249882 466718 249914 466954
rect 249294 466634 249914 466718
rect 249294 466398 249326 466634
rect 249562 466398 249646 466634
rect 249882 466398 249914 466634
rect 249294 430954 249914 466398
rect 249294 430718 249326 430954
rect 249562 430718 249646 430954
rect 249882 430718 249914 430954
rect 249294 430634 249914 430718
rect 249294 430398 249326 430634
rect 249562 430398 249646 430634
rect 249882 430398 249914 430634
rect 249294 394954 249914 430398
rect 249294 394718 249326 394954
rect 249562 394718 249646 394954
rect 249882 394718 249914 394954
rect 249294 394634 249914 394718
rect 249294 394398 249326 394634
rect 249562 394398 249646 394634
rect 249882 394398 249914 394634
rect 249294 358954 249914 394398
rect 249294 358718 249326 358954
rect 249562 358718 249646 358954
rect 249882 358718 249914 358954
rect 249294 358634 249914 358718
rect 249294 358398 249326 358634
rect 249562 358398 249646 358634
rect 249882 358398 249914 358634
rect 249294 322954 249914 358398
rect 249294 322718 249326 322954
rect 249562 322718 249646 322954
rect 249882 322718 249914 322954
rect 249294 322634 249914 322718
rect 249294 322398 249326 322634
rect 249562 322398 249646 322634
rect 249882 322398 249914 322634
rect 249294 286954 249914 322398
rect 249294 286718 249326 286954
rect 249562 286718 249646 286954
rect 249882 286718 249914 286954
rect 249294 286634 249914 286718
rect 249294 286398 249326 286634
rect 249562 286398 249646 286634
rect 249882 286398 249914 286634
rect 249294 250954 249914 286398
rect 249294 250718 249326 250954
rect 249562 250718 249646 250954
rect 249882 250718 249914 250954
rect 249294 250634 249914 250718
rect 249294 250398 249326 250634
rect 249562 250398 249646 250634
rect 249882 250398 249914 250634
rect 249294 214954 249914 250398
rect 249294 214718 249326 214954
rect 249562 214718 249646 214954
rect 249882 214718 249914 214954
rect 249294 214634 249914 214718
rect 249294 214398 249326 214634
rect 249562 214398 249646 214634
rect 249882 214398 249914 214634
rect 249294 178954 249914 214398
rect 249294 178718 249326 178954
rect 249562 178718 249646 178954
rect 249882 178718 249914 178954
rect 249294 178634 249914 178718
rect 249294 178398 249326 178634
rect 249562 178398 249646 178634
rect 249882 178398 249914 178634
rect 249294 142954 249914 178398
rect 249294 142718 249326 142954
rect 249562 142718 249646 142954
rect 249882 142718 249914 142954
rect 249294 142634 249914 142718
rect 249294 142398 249326 142634
rect 249562 142398 249646 142634
rect 249882 142398 249914 142634
rect 249294 106954 249914 142398
rect 249294 106718 249326 106954
rect 249562 106718 249646 106954
rect 249882 106718 249914 106954
rect 249294 106634 249914 106718
rect 249294 106398 249326 106634
rect 249562 106398 249646 106634
rect 249882 106398 249914 106634
rect 249294 70954 249914 106398
rect 249294 70718 249326 70954
rect 249562 70718 249646 70954
rect 249882 70718 249914 70954
rect 249294 70634 249914 70718
rect 249294 70398 249326 70634
rect 249562 70398 249646 70634
rect 249882 70398 249914 70634
rect 249294 34954 249914 70398
rect 249294 34718 249326 34954
rect 249562 34718 249646 34954
rect 249882 34718 249914 34954
rect 249294 34634 249914 34718
rect 249294 34398 249326 34634
rect 249562 34398 249646 34634
rect 249882 34398 249914 34634
rect 249294 -7066 249914 34398
rect 249294 -7302 249326 -7066
rect 249562 -7302 249646 -7066
rect 249882 -7302 249914 -7066
rect 249294 -7386 249914 -7302
rect 249294 -7622 249326 -7386
rect 249562 -7622 249646 -7386
rect 249882 -7622 249914 -7386
rect 249294 -7654 249914 -7622
rect 253794 704838 254414 711590
rect 253794 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 254414 704838
rect 253794 704518 254414 704602
rect 253794 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 254414 704518
rect 253794 687454 254414 704282
rect 253794 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 254414 687454
rect 253794 687134 254414 687218
rect 253794 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 254414 687134
rect 253794 651454 254414 686898
rect 253794 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 254414 651454
rect 253794 651134 254414 651218
rect 253794 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 254414 651134
rect 253794 615454 254414 650898
rect 253794 615218 253826 615454
rect 254062 615218 254146 615454
rect 254382 615218 254414 615454
rect 253794 615134 254414 615218
rect 253794 614898 253826 615134
rect 254062 614898 254146 615134
rect 254382 614898 254414 615134
rect 253794 579454 254414 614898
rect 253794 579218 253826 579454
rect 254062 579218 254146 579454
rect 254382 579218 254414 579454
rect 253794 579134 254414 579218
rect 253794 578898 253826 579134
rect 254062 578898 254146 579134
rect 254382 578898 254414 579134
rect 253794 543454 254414 578898
rect 253794 543218 253826 543454
rect 254062 543218 254146 543454
rect 254382 543218 254414 543454
rect 253794 543134 254414 543218
rect 253794 542898 253826 543134
rect 254062 542898 254146 543134
rect 254382 542898 254414 543134
rect 253794 507454 254414 542898
rect 253794 507218 253826 507454
rect 254062 507218 254146 507454
rect 254382 507218 254414 507454
rect 253794 507134 254414 507218
rect 253794 506898 253826 507134
rect 254062 506898 254146 507134
rect 254382 506898 254414 507134
rect 253794 471454 254414 506898
rect 253794 471218 253826 471454
rect 254062 471218 254146 471454
rect 254382 471218 254414 471454
rect 253794 471134 254414 471218
rect 253794 470898 253826 471134
rect 254062 470898 254146 471134
rect 254382 470898 254414 471134
rect 253794 435454 254414 470898
rect 253794 435218 253826 435454
rect 254062 435218 254146 435454
rect 254382 435218 254414 435454
rect 253794 435134 254414 435218
rect 253794 434898 253826 435134
rect 254062 434898 254146 435134
rect 254382 434898 254414 435134
rect 253794 399454 254414 434898
rect 253794 399218 253826 399454
rect 254062 399218 254146 399454
rect 254382 399218 254414 399454
rect 253794 399134 254414 399218
rect 253794 398898 253826 399134
rect 254062 398898 254146 399134
rect 254382 398898 254414 399134
rect 253794 363454 254414 398898
rect 253794 363218 253826 363454
rect 254062 363218 254146 363454
rect 254382 363218 254414 363454
rect 253794 363134 254414 363218
rect 253794 362898 253826 363134
rect 254062 362898 254146 363134
rect 254382 362898 254414 363134
rect 253794 327454 254414 362898
rect 253794 327218 253826 327454
rect 254062 327218 254146 327454
rect 254382 327218 254414 327454
rect 253794 327134 254414 327218
rect 253794 326898 253826 327134
rect 254062 326898 254146 327134
rect 254382 326898 254414 327134
rect 253794 291454 254414 326898
rect 253794 291218 253826 291454
rect 254062 291218 254146 291454
rect 254382 291218 254414 291454
rect 253794 291134 254414 291218
rect 253794 290898 253826 291134
rect 254062 290898 254146 291134
rect 254382 290898 254414 291134
rect 253794 255454 254414 290898
rect 253794 255218 253826 255454
rect 254062 255218 254146 255454
rect 254382 255218 254414 255454
rect 253794 255134 254414 255218
rect 253794 254898 253826 255134
rect 254062 254898 254146 255134
rect 254382 254898 254414 255134
rect 253794 219454 254414 254898
rect 253794 219218 253826 219454
rect 254062 219218 254146 219454
rect 254382 219218 254414 219454
rect 253794 219134 254414 219218
rect 253794 218898 253826 219134
rect 254062 218898 254146 219134
rect 254382 218898 254414 219134
rect 253794 183454 254414 218898
rect 253794 183218 253826 183454
rect 254062 183218 254146 183454
rect 254382 183218 254414 183454
rect 253794 183134 254414 183218
rect 253794 182898 253826 183134
rect 254062 182898 254146 183134
rect 254382 182898 254414 183134
rect 253794 147454 254414 182898
rect 253794 147218 253826 147454
rect 254062 147218 254146 147454
rect 254382 147218 254414 147454
rect 253794 147134 254414 147218
rect 253794 146898 253826 147134
rect 254062 146898 254146 147134
rect 254382 146898 254414 147134
rect 253794 111454 254414 146898
rect 253794 111218 253826 111454
rect 254062 111218 254146 111454
rect 254382 111218 254414 111454
rect 253794 111134 254414 111218
rect 253794 110898 253826 111134
rect 254062 110898 254146 111134
rect 254382 110898 254414 111134
rect 253794 75454 254414 110898
rect 253794 75218 253826 75454
rect 254062 75218 254146 75454
rect 254382 75218 254414 75454
rect 253794 75134 254414 75218
rect 253794 74898 253826 75134
rect 254062 74898 254146 75134
rect 254382 74898 254414 75134
rect 253794 39454 254414 74898
rect 253794 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 254414 39454
rect 253794 39134 254414 39218
rect 253794 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 254414 39134
rect 253794 3454 254414 38898
rect 253794 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 254414 3454
rect 253794 3134 254414 3218
rect 253794 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 254414 3134
rect 253794 -346 254414 2898
rect 253794 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 254414 -346
rect 253794 -666 254414 -582
rect 253794 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 254414 -666
rect 253794 -7654 254414 -902
rect 258294 705798 258914 711590
rect 258294 705562 258326 705798
rect 258562 705562 258646 705798
rect 258882 705562 258914 705798
rect 258294 705478 258914 705562
rect 258294 705242 258326 705478
rect 258562 705242 258646 705478
rect 258882 705242 258914 705478
rect 258294 691954 258914 705242
rect 258294 691718 258326 691954
rect 258562 691718 258646 691954
rect 258882 691718 258914 691954
rect 258294 691634 258914 691718
rect 258294 691398 258326 691634
rect 258562 691398 258646 691634
rect 258882 691398 258914 691634
rect 258294 655954 258914 691398
rect 258294 655718 258326 655954
rect 258562 655718 258646 655954
rect 258882 655718 258914 655954
rect 258294 655634 258914 655718
rect 258294 655398 258326 655634
rect 258562 655398 258646 655634
rect 258882 655398 258914 655634
rect 258294 619954 258914 655398
rect 258294 619718 258326 619954
rect 258562 619718 258646 619954
rect 258882 619718 258914 619954
rect 258294 619634 258914 619718
rect 258294 619398 258326 619634
rect 258562 619398 258646 619634
rect 258882 619398 258914 619634
rect 258294 583954 258914 619398
rect 258294 583718 258326 583954
rect 258562 583718 258646 583954
rect 258882 583718 258914 583954
rect 258294 583634 258914 583718
rect 258294 583398 258326 583634
rect 258562 583398 258646 583634
rect 258882 583398 258914 583634
rect 258294 547954 258914 583398
rect 258294 547718 258326 547954
rect 258562 547718 258646 547954
rect 258882 547718 258914 547954
rect 258294 547634 258914 547718
rect 258294 547398 258326 547634
rect 258562 547398 258646 547634
rect 258882 547398 258914 547634
rect 258294 511954 258914 547398
rect 258294 511718 258326 511954
rect 258562 511718 258646 511954
rect 258882 511718 258914 511954
rect 258294 511634 258914 511718
rect 258294 511398 258326 511634
rect 258562 511398 258646 511634
rect 258882 511398 258914 511634
rect 258294 475954 258914 511398
rect 258294 475718 258326 475954
rect 258562 475718 258646 475954
rect 258882 475718 258914 475954
rect 258294 475634 258914 475718
rect 258294 475398 258326 475634
rect 258562 475398 258646 475634
rect 258882 475398 258914 475634
rect 258294 439954 258914 475398
rect 258294 439718 258326 439954
rect 258562 439718 258646 439954
rect 258882 439718 258914 439954
rect 258294 439634 258914 439718
rect 258294 439398 258326 439634
rect 258562 439398 258646 439634
rect 258882 439398 258914 439634
rect 258294 403954 258914 439398
rect 258294 403718 258326 403954
rect 258562 403718 258646 403954
rect 258882 403718 258914 403954
rect 258294 403634 258914 403718
rect 258294 403398 258326 403634
rect 258562 403398 258646 403634
rect 258882 403398 258914 403634
rect 258294 367954 258914 403398
rect 258294 367718 258326 367954
rect 258562 367718 258646 367954
rect 258882 367718 258914 367954
rect 258294 367634 258914 367718
rect 258294 367398 258326 367634
rect 258562 367398 258646 367634
rect 258882 367398 258914 367634
rect 258294 331954 258914 367398
rect 258294 331718 258326 331954
rect 258562 331718 258646 331954
rect 258882 331718 258914 331954
rect 258294 331634 258914 331718
rect 258294 331398 258326 331634
rect 258562 331398 258646 331634
rect 258882 331398 258914 331634
rect 258294 295954 258914 331398
rect 258294 295718 258326 295954
rect 258562 295718 258646 295954
rect 258882 295718 258914 295954
rect 258294 295634 258914 295718
rect 258294 295398 258326 295634
rect 258562 295398 258646 295634
rect 258882 295398 258914 295634
rect 258294 259954 258914 295398
rect 258294 259718 258326 259954
rect 258562 259718 258646 259954
rect 258882 259718 258914 259954
rect 258294 259634 258914 259718
rect 258294 259398 258326 259634
rect 258562 259398 258646 259634
rect 258882 259398 258914 259634
rect 258294 223954 258914 259398
rect 258294 223718 258326 223954
rect 258562 223718 258646 223954
rect 258882 223718 258914 223954
rect 258294 223634 258914 223718
rect 258294 223398 258326 223634
rect 258562 223398 258646 223634
rect 258882 223398 258914 223634
rect 258294 187954 258914 223398
rect 258294 187718 258326 187954
rect 258562 187718 258646 187954
rect 258882 187718 258914 187954
rect 258294 187634 258914 187718
rect 258294 187398 258326 187634
rect 258562 187398 258646 187634
rect 258882 187398 258914 187634
rect 258294 151954 258914 187398
rect 258294 151718 258326 151954
rect 258562 151718 258646 151954
rect 258882 151718 258914 151954
rect 258294 151634 258914 151718
rect 258294 151398 258326 151634
rect 258562 151398 258646 151634
rect 258882 151398 258914 151634
rect 258294 115954 258914 151398
rect 258294 115718 258326 115954
rect 258562 115718 258646 115954
rect 258882 115718 258914 115954
rect 258294 115634 258914 115718
rect 258294 115398 258326 115634
rect 258562 115398 258646 115634
rect 258882 115398 258914 115634
rect 258294 79954 258914 115398
rect 258294 79718 258326 79954
rect 258562 79718 258646 79954
rect 258882 79718 258914 79954
rect 258294 79634 258914 79718
rect 258294 79398 258326 79634
rect 258562 79398 258646 79634
rect 258882 79398 258914 79634
rect 258294 43954 258914 79398
rect 258294 43718 258326 43954
rect 258562 43718 258646 43954
rect 258882 43718 258914 43954
rect 258294 43634 258914 43718
rect 258294 43398 258326 43634
rect 258562 43398 258646 43634
rect 258882 43398 258914 43634
rect 258294 7954 258914 43398
rect 258294 7718 258326 7954
rect 258562 7718 258646 7954
rect 258882 7718 258914 7954
rect 258294 7634 258914 7718
rect 258294 7398 258326 7634
rect 258562 7398 258646 7634
rect 258882 7398 258914 7634
rect 258294 -1306 258914 7398
rect 258294 -1542 258326 -1306
rect 258562 -1542 258646 -1306
rect 258882 -1542 258914 -1306
rect 258294 -1626 258914 -1542
rect 258294 -1862 258326 -1626
rect 258562 -1862 258646 -1626
rect 258882 -1862 258914 -1626
rect 258294 -7654 258914 -1862
rect 262794 706758 263414 711590
rect 262794 706522 262826 706758
rect 263062 706522 263146 706758
rect 263382 706522 263414 706758
rect 262794 706438 263414 706522
rect 262794 706202 262826 706438
rect 263062 706202 263146 706438
rect 263382 706202 263414 706438
rect 262794 696454 263414 706202
rect 262794 696218 262826 696454
rect 263062 696218 263146 696454
rect 263382 696218 263414 696454
rect 262794 696134 263414 696218
rect 262794 695898 262826 696134
rect 263062 695898 263146 696134
rect 263382 695898 263414 696134
rect 262794 660454 263414 695898
rect 262794 660218 262826 660454
rect 263062 660218 263146 660454
rect 263382 660218 263414 660454
rect 262794 660134 263414 660218
rect 262794 659898 262826 660134
rect 263062 659898 263146 660134
rect 263382 659898 263414 660134
rect 262794 624454 263414 659898
rect 262794 624218 262826 624454
rect 263062 624218 263146 624454
rect 263382 624218 263414 624454
rect 262794 624134 263414 624218
rect 262794 623898 262826 624134
rect 263062 623898 263146 624134
rect 263382 623898 263414 624134
rect 262794 588454 263414 623898
rect 262794 588218 262826 588454
rect 263062 588218 263146 588454
rect 263382 588218 263414 588454
rect 262794 588134 263414 588218
rect 262794 587898 262826 588134
rect 263062 587898 263146 588134
rect 263382 587898 263414 588134
rect 262794 552454 263414 587898
rect 262794 552218 262826 552454
rect 263062 552218 263146 552454
rect 263382 552218 263414 552454
rect 262794 552134 263414 552218
rect 262794 551898 262826 552134
rect 263062 551898 263146 552134
rect 263382 551898 263414 552134
rect 262794 516454 263414 551898
rect 262794 516218 262826 516454
rect 263062 516218 263146 516454
rect 263382 516218 263414 516454
rect 262794 516134 263414 516218
rect 262794 515898 262826 516134
rect 263062 515898 263146 516134
rect 263382 515898 263414 516134
rect 262794 480454 263414 515898
rect 262794 480218 262826 480454
rect 263062 480218 263146 480454
rect 263382 480218 263414 480454
rect 262794 480134 263414 480218
rect 262794 479898 262826 480134
rect 263062 479898 263146 480134
rect 263382 479898 263414 480134
rect 262794 444454 263414 479898
rect 262794 444218 262826 444454
rect 263062 444218 263146 444454
rect 263382 444218 263414 444454
rect 262794 444134 263414 444218
rect 262794 443898 262826 444134
rect 263062 443898 263146 444134
rect 263382 443898 263414 444134
rect 262794 408454 263414 443898
rect 262794 408218 262826 408454
rect 263062 408218 263146 408454
rect 263382 408218 263414 408454
rect 262794 408134 263414 408218
rect 262794 407898 262826 408134
rect 263062 407898 263146 408134
rect 263382 407898 263414 408134
rect 262794 372454 263414 407898
rect 262794 372218 262826 372454
rect 263062 372218 263146 372454
rect 263382 372218 263414 372454
rect 262794 372134 263414 372218
rect 262794 371898 262826 372134
rect 263062 371898 263146 372134
rect 263382 371898 263414 372134
rect 262794 336454 263414 371898
rect 262794 336218 262826 336454
rect 263062 336218 263146 336454
rect 263382 336218 263414 336454
rect 262794 336134 263414 336218
rect 262794 335898 262826 336134
rect 263062 335898 263146 336134
rect 263382 335898 263414 336134
rect 262794 300454 263414 335898
rect 262794 300218 262826 300454
rect 263062 300218 263146 300454
rect 263382 300218 263414 300454
rect 262794 300134 263414 300218
rect 262794 299898 262826 300134
rect 263062 299898 263146 300134
rect 263382 299898 263414 300134
rect 262794 264454 263414 299898
rect 262794 264218 262826 264454
rect 263062 264218 263146 264454
rect 263382 264218 263414 264454
rect 262794 264134 263414 264218
rect 262794 263898 262826 264134
rect 263062 263898 263146 264134
rect 263382 263898 263414 264134
rect 262794 228454 263414 263898
rect 262794 228218 262826 228454
rect 263062 228218 263146 228454
rect 263382 228218 263414 228454
rect 262794 228134 263414 228218
rect 262794 227898 262826 228134
rect 263062 227898 263146 228134
rect 263382 227898 263414 228134
rect 262794 192454 263414 227898
rect 262794 192218 262826 192454
rect 263062 192218 263146 192454
rect 263382 192218 263414 192454
rect 262794 192134 263414 192218
rect 262794 191898 262826 192134
rect 263062 191898 263146 192134
rect 263382 191898 263414 192134
rect 262794 156454 263414 191898
rect 262794 156218 262826 156454
rect 263062 156218 263146 156454
rect 263382 156218 263414 156454
rect 262794 156134 263414 156218
rect 262794 155898 262826 156134
rect 263062 155898 263146 156134
rect 263382 155898 263414 156134
rect 262794 120454 263414 155898
rect 262794 120218 262826 120454
rect 263062 120218 263146 120454
rect 263382 120218 263414 120454
rect 262794 120134 263414 120218
rect 262794 119898 262826 120134
rect 263062 119898 263146 120134
rect 263382 119898 263414 120134
rect 262794 84454 263414 119898
rect 262794 84218 262826 84454
rect 263062 84218 263146 84454
rect 263382 84218 263414 84454
rect 262794 84134 263414 84218
rect 262794 83898 262826 84134
rect 263062 83898 263146 84134
rect 263382 83898 263414 84134
rect 262794 48454 263414 83898
rect 262794 48218 262826 48454
rect 263062 48218 263146 48454
rect 263382 48218 263414 48454
rect 262794 48134 263414 48218
rect 262794 47898 262826 48134
rect 263062 47898 263146 48134
rect 263382 47898 263414 48134
rect 262794 12454 263414 47898
rect 262794 12218 262826 12454
rect 263062 12218 263146 12454
rect 263382 12218 263414 12454
rect 262794 12134 263414 12218
rect 262794 11898 262826 12134
rect 263062 11898 263146 12134
rect 263382 11898 263414 12134
rect 262794 -2266 263414 11898
rect 262794 -2502 262826 -2266
rect 263062 -2502 263146 -2266
rect 263382 -2502 263414 -2266
rect 262794 -2586 263414 -2502
rect 262794 -2822 262826 -2586
rect 263062 -2822 263146 -2586
rect 263382 -2822 263414 -2586
rect 262794 -7654 263414 -2822
rect 267294 707718 267914 711590
rect 267294 707482 267326 707718
rect 267562 707482 267646 707718
rect 267882 707482 267914 707718
rect 267294 707398 267914 707482
rect 267294 707162 267326 707398
rect 267562 707162 267646 707398
rect 267882 707162 267914 707398
rect 267294 700954 267914 707162
rect 267294 700718 267326 700954
rect 267562 700718 267646 700954
rect 267882 700718 267914 700954
rect 267294 700634 267914 700718
rect 267294 700398 267326 700634
rect 267562 700398 267646 700634
rect 267882 700398 267914 700634
rect 267294 664954 267914 700398
rect 267294 664718 267326 664954
rect 267562 664718 267646 664954
rect 267882 664718 267914 664954
rect 267294 664634 267914 664718
rect 267294 664398 267326 664634
rect 267562 664398 267646 664634
rect 267882 664398 267914 664634
rect 267294 628954 267914 664398
rect 267294 628718 267326 628954
rect 267562 628718 267646 628954
rect 267882 628718 267914 628954
rect 267294 628634 267914 628718
rect 267294 628398 267326 628634
rect 267562 628398 267646 628634
rect 267882 628398 267914 628634
rect 267294 592954 267914 628398
rect 267294 592718 267326 592954
rect 267562 592718 267646 592954
rect 267882 592718 267914 592954
rect 267294 592634 267914 592718
rect 267294 592398 267326 592634
rect 267562 592398 267646 592634
rect 267882 592398 267914 592634
rect 267294 556954 267914 592398
rect 267294 556718 267326 556954
rect 267562 556718 267646 556954
rect 267882 556718 267914 556954
rect 267294 556634 267914 556718
rect 267294 556398 267326 556634
rect 267562 556398 267646 556634
rect 267882 556398 267914 556634
rect 267294 520954 267914 556398
rect 267294 520718 267326 520954
rect 267562 520718 267646 520954
rect 267882 520718 267914 520954
rect 267294 520634 267914 520718
rect 267294 520398 267326 520634
rect 267562 520398 267646 520634
rect 267882 520398 267914 520634
rect 267294 484954 267914 520398
rect 267294 484718 267326 484954
rect 267562 484718 267646 484954
rect 267882 484718 267914 484954
rect 267294 484634 267914 484718
rect 267294 484398 267326 484634
rect 267562 484398 267646 484634
rect 267882 484398 267914 484634
rect 267294 448954 267914 484398
rect 267294 448718 267326 448954
rect 267562 448718 267646 448954
rect 267882 448718 267914 448954
rect 267294 448634 267914 448718
rect 267294 448398 267326 448634
rect 267562 448398 267646 448634
rect 267882 448398 267914 448634
rect 267294 412954 267914 448398
rect 267294 412718 267326 412954
rect 267562 412718 267646 412954
rect 267882 412718 267914 412954
rect 267294 412634 267914 412718
rect 267294 412398 267326 412634
rect 267562 412398 267646 412634
rect 267882 412398 267914 412634
rect 267294 376954 267914 412398
rect 267294 376718 267326 376954
rect 267562 376718 267646 376954
rect 267882 376718 267914 376954
rect 267294 376634 267914 376718
rect 267294 376398 267326 376634
rect 267562 376398 267646 376634
rect 267882 376398 267914 376634
rect 267294 340954 267914 376398
rect 267294 340718 267326 340954
rect 267562 340718 267646 340954
rect 267882 340718 267914 340954
rect 267294 340634 267914 340718
rect 267294 340398 267326 340634
rect 267562 340398 267646 340634
rect 267882 340398 267914 340634
rect 267294 304954 267914 340398
rect 267294 304718 267326 304954
rect 267562 304718 267646 304954
rect 267882 304718 267914 304954
rect 267294 304634 267914 304718
rect 267294 304398 267326 304634
rect 267562 304398 267646 304634
rect 267882 304398 267914 304634
rect 267294 268954 267914 304398
rect 267294 268718 267326 268954
rect 267562 268718 267646 268954
rect 267882 268718 267914 268954
rect 267294 268634 267914 268718
rect 267294 268398 267326 268634
rect 267562 268398 267646 268634
rect 267882 268398 267914 268634
rect 267294 232954 267914 268398
rect 267294 232718 267326 232954
rect 267562 232718 267646 232954
rect 267882 232718 267914 232954
rect 267294 232634 267914 232718
rect 267294 232398 267326 232634
rect 267562 232398 267646 232634
rect 267882 232398 267914 232634
rect 267294 196954 267914 232398
rect 267294 196718 267326 196954
rect 267562 196718 267646 196954
rect 267882 196718 267914 196954
rect 267294 196634 267914 196718
rect 267294 196398 267326 196634
rect 267562 196398 267646 196634
rect 267882 196398 267914 196634
rect 267294 160954 267914 196398
rect 267294 160718 267326 160954
rect 267562 160718 267646 160954
rect 267882 160718 267914 160954
rect 267294 160634 267914 160718
rect 267294 160398 267326 160634
rect 267562 160398 267646 160634
rect 267882 160398 267914 160634
rect 267294 124954 267914 160398
rect 267294 124718 267326 124954
rect 267562 124718 267646 124954
rect 267882 124718 267914 124954
rect 267294 124634 267914 124718
rect 267294 124398 267326 124634
rect 267562 124398 267646 124634
rect 267882 124398 267914 124634
rect 267294 88954 267914 124398
rect 267294 88718 267326 88954
rect 267562 88718 267646 88954
rect 267882 88718 267914 88954
rect 267294 88634 267914 88718
rect 267294 88398 267326 88634
rect 267562 88398 267646 88634
rect 267882 88398 267914 88634
rect 267294 52954 267914 88398
rect 267294 52718 267326 52954
rect 267562 52718 267646 52954
rect 267882 52718 267914 52954
rect 267294 52634 267914 52718
rect 267294 52398 267326 52634
rect 267562 52398 267646 52634
rect 267882 52398 267914 52634
rect 267294 16954 267914 52398
rect 267294 16718 267326 16954
rect 267562 16718 267646 16954
rect 267882 16718 267914 16954
rect 267294 16634 267914 16718
rect 267294 16398 267326 16634
rect 267562 16398 267646 16634
rect 267882 16398 267914 16634
rect 267294 -3226 267914 16398
rect 267294 -3462 267326 -3226
rect 267562 -3462 267646 -3226
rect 267882 -3462 267914 -3226
rect 267294 -3546 267914 -3462
rect 267294 -3782 267326 -3546
rect 267562 -3782 267646 -3546
rect 267882 -3782 267914 -3546
rect 267294 -7654 267914 -3782
rect 271794 708678 272414 711590
rect 271794 708442 271826 708678
rect 272062 708442 272146 708678
rect 272382 708442 272414 708678
rect 271794 708358 272414 708442
rect 271794 708122 271826 708358
rect 272062 708122 272146 708358
rect 272382 708122 272414 708358
rect 271794 669454 272414 708122
rect 271794 669218 271826 669454
rect 272062 669218 272146 669454
rect 272382 669218 272414 669454
rect 271794 669134 272414 669218
rect 271794 668898 271826 669134
rect 272062 668898 272146 669134
rect 272382 668898 272414 669134
rect 271794 633454 272414 668898
rect 271794 633218 271826 633454
rect 272062 633218 272146 633454
rect 272382 633218 272414 633454
rect 271794 633134 272414 633218
rect 271794 632898 271826 633134
rect 272062 632898 272146 633134
rect 272382 632898 272414 633134
rect 271794 597454 272414 632898
rect 271794 597218 271826 597454
rect 272062 597218 272146 597454
rect 272382 597218 272414 597454
rect 271794 597134 272414 597218
rect 271794 596898 271826 597134
rect 272062 596898 272146 597134
rect 272382 596898 272414 597134
rect 271794 561454 272414 596898
rect 271794 561218 271826 561454
rect 272062 561218 272146 561454
rect 272382 561218 272414 561454
rect 271794 561134 272414 561218
rect 271794 560898 271826 561134
rect 272062 560898 272146 561134
rect 272382 560898 272414 561134
rect 271794 525454 272414 560898
rect 271794 525218 271826 525454
rect 272062 525218 272146 525454
rect 272382 525218 272414 525454
rect 271794 525134 272414 525218
rect 271794 524898 271826 525134
rect 272062 524898 272146 525134
rect 272382 524898 272414 525134
rect 271794 489454 272414 524898
rect 271794 489218 271826 489454
rect 272062 489218 272146 489454
rect 272382 489218 272414 489454
rect 271794 489134 272414 489218
rect 271794 488898 271826 489134
rect 272062 488898 272146 489134
rect 272382 488898 272414 489134
rect 271794 453454 272414 488898
rect 271794 453218 271826 453454
rect 272062 453218 272146 453454
rect 272382 453218 272414 453454
rect 271794 453134 272414 453218
rect 271794 452898 271826 453134
rect 272062 452898 272146 453134
rect 272382 452898 272414 453134
rect 271794 417454 272414 452898
rect 271794 417218 271826 417454
rect 272062 417218 272146 417454
rect 272382 417218 272414 417454
rect 271794 417134 272414 417218
rect 271794 416898 271826 417134
rect 272062 416898 272146 417134
rect 272382 416898 272414 417134
rect 271794 381454 272414 416898
rect 271794 381218 271826 381454
rect 272062 381218 272146 381454
rect 272382 381218 272414 381454
rect 271794 381134 272414 381218
rect 271794 380898 271826 381134
rect 272062 380898 272146 381134
rect 272382 380898 272414 381134
rect 271794 345454 272414 380898
rect 271794 345218 271826 345454
rect 272062 345218 272146 345454
rect 272382 345218 272414 345454
rect 271794 345134 272414 345218
rect 271794 344898 271826 345134
rect 272062 344898 272146 345134
rect 272382 344898 272414 345134
rect 271794 309454 272414 344898
rect 271794 309218 271826 309454
rect 272062 309218 272146 309454
rect 272382 309218 272414 309454
rect 271794 309134 272414 309218
rect 271794 308898 271826 309134
rect 272062 308898 272146 309134
rect 272382 308898 272414 309134
rect 271794 273454 272414 308898
rect 271794 273218 271826 273454
rect 272062 273218 272146 273454
rect 272382 273218 272414 273454
rect 271794 273134 272414 273218
rect 271794 272898 271826 273134
rect 272062 272898 272146 273134
rect 272382 272898 272414 273134
rect 271794 237454 272414 272898
rect 271794 237218 271826 237454
rect 272062 237218 272146 237454
rect 272382 237218 272414 237454
rect 271794 237134 272414 237218
rect 271794 236898 271826 237134
rect 272062 236898 272146 237134
rect 272382 236898 272414 237134
rect 271794 201454 272414 236898
rect 271794 201218 271826 201454
rect 272062 201218 272146 201454
rect 272382 201218 272414 201454
rect 271794 201134 272414 201218
rect 271794 200898 271826 201134
rect 272062 200898 272146 201134
rect 272382 200898 272414 201134
rect 271794 165454 272414 200898
rect 271794 165218 271826 165454
rect 272062 165218 272146 165454
rect 272382 165218 272414 165454
rect 271794 165134 272414 165218
rect 271794 164898 271826 165134
rect 272062 164898 272146 165134
rect 272382 164898 272414 165134
rect 271794 129454 272414 164898
rect 271794 129218 271826 129454
rect 272062 129218 272146 129454
rect 272382 129218 272414 129454
rect 271794 129134 272414 129218
rect 271794 128898 271826 129134
rect 272062 128898 272146 129134
rect 272382 128898 272414 129134
rect 271794 93454 272414 128898
rect 271794 93218 271826 93454
rect 272062 93218 272146 93454
rect 272382 93218 272414 93454
rect 271794 93134 272414 93218
rect 271794 92898 271826 93134
rect 272062 92898 272146 93134
rect 272382 92898 272414 93134
rect 271794 57454 272414 92898
rect 271794 57218 271826 57454
rect 272062 57218 272146 57454
rect 272382 57218 272414 57454
rect 271794 57134 272414 57218
rect 271794 56898 271826 57134
rect 272062 56898 272146 57134
rect 272382 56898 272414 57134
rect 271794 21454 272414 56898
rect 271794 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 272414 21454
rect 271794 21134 272414 21218
rect 271794 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 272414 21134
rect 271794 -4186 272414 20898
rect 271794 -4422 271826 -4186
rect 272062 -4422 272146 -4186
rect 272382 -4422 272414 -4186
rect 271794 -4506 272414 -4422
rect 271794 -4742 271826 -4506
rect 272062 -4742 272146 -4506
rect 272382 -4742 272414 -4506
rect 271794 -7654 272414 -4742
rect 276294 709638 276914 711590
rect 276294 709402 276326 709638
rect 276562 709402 276646 709638
rect 276882 709402 276914 709638
rect 276294 709318 276914 709402
rect 276294 709082 276326 709318
rect 276562 709082 276646 709318
rect 276882 709082 276914 709318
rect 276294 673954 276914 709082
rect 276294 673718 276326 673954
rect 276562 673718 276646 673954
rect 276882 673718 276914 673954
rect 276294 673634 276914 673718
rect 276294 673398 276326 673634
rect 276562 673398 276646 673634
rect 276882 673398 276914 673634
rect 276294 637954 276914 673398
rect 276294 637718 276326 637954
rect 276562 637718 276646 637954
rect 276882 637718 276914 637954
rect 276294 637634 276914 637718
rect 276294 637398 276326 637634
rect 276562 637398 276646 637634
rect 276882 637398 276914 637634
rect 276294 601954 276914 637398
rect 276294 601718 276326 601954
rect 276562 601718 276646 601954
rect 276882 601718 276914 601954
rect 276294 601634 276914 601718
rect 276294 601398 276326 601634
rect 276562 601398 276646 601634
rect 276882 601398 276914 601634
rect 276294 565954 276914 601398
rect 276294 565718 276326 565954
rect 276562 565718 276646 565954
rect 276882 565718 276914 565954
rect 276294 565634 276914 565718
rect 276294 565398 276326 565634
rect 276562 565398 276646 565634
rect 276882 565398 276914 565634
rect 276294 529954 276914 565398
rect 276294 529718 276326 529954
rect 276562 529718 276646 529954
rect 276882 529718 276914 529954
rect 276294 529634 276914 529718
rect 276294 529398 276326 529634
rect 276562 529398 276646 529634
rect 276882 529398 276914 529634
rect 276294 493954 276914 529398
rect 276294 493718 276326 493954
rect 276562 493718 276646 493954
rect 276882 493718 276914 493954
rect 276294 493634 276914 493718
rect 276294 493398 276326 493634
rect 276562 493398 276646 493634
rect 276882 493398 276914 493634
rect 276294 457954 276914 493398
rect 276294 457718 276326 457954
rect 276562 457718 276646 457954
rect 276882 457718 276914 457954
rect 276294 457634 276914 457718
rect 276294 457398 276326 457634
rect 276562 457398 276646 457634
rect 276882 457398 276914 457634
rect 276294 421954 276914 457398
rect 276294 421718 276326 421954
rect 276562 421718 276646 421954
rect 276882 421718 276914 421954
rect 276294 421634 276914 421718
rect 276294 421398 276326 421634
rect 276562 421398 276646 421634
rect 276882 421398 276914 421634
rect 276294 385954 276914 421398
rect 276294 385718 276326 385954
rect 276562 385718 276646 385954
rect 276882 385718 276914 385954
rect 276294 385634 276914 385718
rect 276294 385398 276326 385634
rect 276562 385398 276646 385634
rect 276882 385398 276914 385634
rect 276294 349954 276914 385398
rect 276294 349718 276326 349954
rect 276562 349718 276646 349954
rect 276882 349718 276914 349954
rect 276294 349634 276914 349718
rect 276294 349398 276326 349634
rect 276562 349398 276646 349634
rect 276882 349398 276914 349634
rect 276294 313954 276914 349398
rect 276294 313718 276326 313954
rect 276562 313718 276646 313954
rect 276882 313718 276914 313954
rect 276294 313634 276914 313718
rect 276294 313398 276326 313634
rect 276562 313398 276646 313634
rect 276882 313398 276914 313634
rect 276294 277954 276914 313398
rect 276294 277718 276326 277954
rect 276562 277718 276646 277954
rect 276882 277718 276914 277954
rect 276294 277634 276914 277718
rect 276294 277398 276326 277634
rect 276562 277398 276646 277634
rect 276882 277398 276914 277634
rect 276294 241954 276914 277398
rect 276294 241718 276326 241954
rect 276562 241718 276646 241954
rect 276882 241718 276914 241954
rect 276294 241634 276914 241718
rect 276294 241398 276326 241634
rect 276562 241398 276646 241634
rect 276882 241398 276914 241634
rect 276294 205954 276914 241398
rect 276294 205718 276326 205954
rect 276562 205718 276646 205954
rect 276882 205718 276914 205954
rect 276294 205634 276914 205718
rect 276294 205398 276326 205634
rect 276562 205398 276646 205634
rect 276882 205398 276914 205634
rect 276294 169954 276914 205398
rect 276294 169718 276326 169954
rect 276562 169718 276646 169954
rect 276882 169718 276914 169954
rect 276294 169634 276914 169718
rect 276294 169398 276326 169634
rect 276562 169398 276646 169634
rect 276882 169398 276914 169634
rect 276294 133954 276914 169398
rect 276294 133718 276326 133954
rect 276562 133718 276646 133954
rect 276882 133718 276914 133954
rect 276294 133634 276914 133718
rect 276294 133398 276326 133634
rect 276562 133398 276646 133634
rect 276882 133398 276914 133634
rect 276294 97954 276914 133398
rect 276294 97718 276326 97954
rect 276562 97718 276646 97954
rect 276882 97718 276914 97954
rect 276294 97634 276914 97718
rect 276294 97398 276326 97634
rect 276562 97398 276646 97634
rect 276882 97398 276914 97634
rect 276294 61954 276914 97398
rect 276294 61718 276326 61954
rect 276562 61718 276646 61954
rect 276882 61718 276914 61954
rect 276294 61634 276914 61718
rect 276294 61398 276326 61634
rect 276562 61398 276646 61634
rect 276882 61398 276914 61634
rect 276294 25954 276914 61398
rect 276294 25718 276326 25954
rect 276562 25718 276646 25954
rect 276882 25718 276914 25954
rect 276294 25634 276914 25718
rect 276294 25398 276326 25634
rect 276562 25398 276646 25634
rect 276882 25398 276914 25634
rect 276294 -5146 276914 25398
rect 276294 -5382 276326 -5146
rect 276562 -5382 276646 -5146
rect 276882 -5382 276914 -5146
rect 276294 -5466 276914 -5382
rect 276294 -5702 276326 -5466
rect 276562 -5702 276646 -5466
rect 276882 -5702 276914 -5466
rect 276294 -7654 276914 -5702
rect 280794 710598 281414 711590
rect 280794 710362 280826 710598
rect 281062 710362 281146 710598
rect 281382 710362 281414 710598
rect 280794 710278 281414 710362
rect 280794 710042 280826 710278
rect 281062 710042 281146 710278
rect 281382 710042 281414 710278
rect 280794 678454 281414 710042
rect 280794 678218 280826 678454
rect 281062 678218 281146 678454
rect 281382 678218 281414 678454
rect 280794 678134 281414 678218
rect 280794 677898 280826 678134
rect 281062 677898 281146 678134
rect 281382 677898 281414 678134
rect 280794 642454 281414 677898
rect 280794 642218 280826 642454
rect 281062 642218 281146 642454
rect 281382 642218 281414 642454
rect 280794 642134 281414 642218
rect 280794 641898 280826 642134
rect 281062 641898 281146 642134
rect 281382 641898 281414 642134
rect 280794 606454 281414 641898
rect 280794 606218 280826 606454
rect 281062 606218 281146 606454
rect 281382 606218 281414 606454
rect 280794 606134 281414 606218
rect 280794 605898 280826 606134
rect 281062 605898 281146 606134
rect 281382 605898 281414 606134
rect 280794 570454 281414 605898
rect 280794 570218 280826 570454
rect 281062 570218 281146 570454
rect 281382 570218 281414 570454
rect 280794 570134 281414 570218
rect 280794 569898 280826 570134
rect 281062 569898 281146 570134
rect 281382 569898 281414 570134
rect 280794 534454 281414 569898
rect 280794 534218 280826 534454
rect 281062 534218 281146 534454
rect 281382 534218 281414 534454
rect 280794 534134 281414 534218
rect 280794 533898 280826 534134
rect 281062 533898 281146 534134
rect 281382 533898 281414 534134
rect 280794 498454 281414 533898
rect 280794 498218 280826 498454
rect 281062 498218 281146 498454
rect 281382 498218 281414 498454
rect 280794 498134 281414 498218
rect 280794 497898 280826 498134
rect 281062 497898 281146 498134
rect 281382 497898 281414 498134
rect 280794 462454 281414 497898
rect 280794 462218 280826 462454
rect 281062 462218 281146 462454
rect 281382 462218 281414 462454
rect 280794 462134 281414 462218
rect 280794 461898 280826 462134
rect 281062 461898 281146 462134
rect 281382 461898 281414 462134
rect 280794 426454 281414 461898
rect 280794 426218 280826 426454
rect 281062 426218 281146 426454
rect 281382 426218 281414 426454
rect 280794 426134 281414 426218
rect 280794 425898 280826 426134
rect 281062 425898 281146 426134
rect 281382 425898 281414 426134
rect 280794 390454 281414 425898
rect 280794 390218 280826 390454
rect 281062 390218 281146 390454
rect 281382 390218 281414 390454
rect 280794 390134 281414 390218
rect 280794 389898 280826 390134
rect 281062 389898 281146 390134
rect 281382 389898 281414 390134
rect 280794 354454 281414 389898
rect 280794 354218 280826 354454
rect 281062 354218 281146 354454
rect 281382 354218 281414 354454
rect 280794 354134 281414 354218
rect 280794 353898 280826 354134
rect 281062 353898 281146 354134
rect 281382 353898 281414 354134
rect 280794 318454 281414 353898
rect 280794 318218 280826 318454
rect 281062 318218 281146 318454
rect 281382 318218 281414 318454
rect 280794 318134 281414 318218
rect 280794 317898 280826 318134
rect 281062 317898 281146 318134
rect 281382 317898 281414 318134
rect 280794 282454 281414 317898
rect 280794 282218 280826 282454
rect 281062 282218 281146 282454
rect 281382 282218 281414 282454
rect 280794 282134 281414 282218
rect 280794 281898 280826 282134
rect 281062 281898 281146 282134
rect 281382 281898 281414 282134
rect 280794 246454 281414 281898
rect 280794 246218 280826 246454
rect 281062 246218 281146 246454
rect 281382 246218 281414 246454
rect 280794 246134 281414 246218
rect 280794 245898 280826 246134
rect 281062 245898 281146 246134
rect 281382 245898 281414 246134
rect 280794 210454 281414 245898
rect 280794 210218 280826 210454
rect 281062 210218 281146 210454
rect 281382 210218 281414 210454
rect 280794 210134 281414 210218
rect 280794 209898 280826 210134
rect 281062 209898 281146 210134
rect 281382 209898 281414 210134
rect 280794 174454 281414 209898
rect 280794 174218 280826 174454
rect 281062 174218 281146 174454
rect 281382 174218 281414 174454
rect 280794 174134 281414 174218
rect 280794 173898 280826 174134
rect 281062 173898 281146 174134
rect 281382 173898 281414 174134
rect 280794 138454 281414 173898
rect 280794 138218 280826 138454
rect 281062 138218 281146 138454
rect 281382 138218 281414 138454
rect 280794 138134 281414 138218
rect 280794 137898 280826 138134
rect 281062 137898 281146 138134
rect 281382 137898 281414 138134
rect 280794 102454 281414 137898
rect 280794 102218 280826 102454
rect 281062 102218 281146 102454
rect 281382 102218 281414 102454
rect 280794 102134 281414 102218
rect 280794 101898 280826 102134
rect 281062 101898 281146 102134
rect 281382 101898 281414 102134
rect 280794 66454 281414 101898
rect 280794 66218 280826 66454
rect 281062 66218 281146 66454
rect 281382 66218 281414 66454
rect 280794 66134 281414 66218
rect 280794 65898 280826 66134
rect 281062 65898 281146 66134
rect 281382 65898 281414 66134
rect 280794 30454 281414 65898
rect 280794 30218 280826 30454
rect 281062 30218 281146 30454
rect 281382 30218 281414 30454
rect 280794 30134 281414 30218
rect 280794 29898 280826 30134
rect 281062 29898 281146 30134
rect 281382 29898 281414 30134
rect 280794 -6106 281414 29898
rect 280794 -6342 280826 -6106
rect 281062 -6342 281146 -6106
rect 281382 -6342 281414 -6106
rect 280794 -6426 281414 -6342
rect 280794 -6662 280826 -6426
rect 281062 -6662 281146 -6426
rect 281382 -6662 281414 -6426
rect 280794 -7654 281414 -6662
rect 285294 711558 285914 711590
rect 285294 711322 285326 711558
rect 285562 711322 285646 711558
rect 285882 711322 285914 711558
rect 285294 711238 285914 711322
rect 285294 711002 285326 711238
rect 285562 711002 285646 711238
rect 285882 711002 285914 711238
rect 285294 682954 285914 711002
rect 285294 682718 285326 682954
rect 285562 682718 285646 682954
rect 285882 682718 285914 682954
rect 285294 682634 285914 682718
rect 285294 682398 285326 682634
rect 285562 682398 285646 682634
rect 285882 682398 285914 682634
rect 285294 646954 285914 682398
rect 285294 646718 285326 646954
rect 285562 646718 285646 646954
rect 285882 646718 285914 646954
rect 285294 646634 285914 646718
rect 285294 646398 285326 646634
rect 285562 646398 285646 646634
rect 285882 646398 285914 646634
rect 285294 610954 285914 646398
rect 285294 610718 285326 610954
rect 285562 610718 285646 610954
rect 285882 610718 285914 610954
rect 285294 610634 285914 610718
rect 285294 610398 285326 610634
rect 285562 610398 285646 610634
rect 285882 610398 285914 610634
rect 285294 574954 285914 610398
rect 285294 574718 285326 574954
rect 285562 574718 285646 574954
rect 285882 574718 285914 574954
rect 285294 574634 285914 574718
rect 285294 574398 285326 574634
rect 285562 574398 285646 574634
rect 285882 574398 285914 574634
rect 285294 538954 285914 574398
rect 285294 538718 285326 538954
rect 285562 538718 285646 538954
rect 285882 538718 285914 538954
rect 285294 538634 285914 538718
rect 285294 538398 285326 538634
rect 285562 538398 285646 538634
rect 285882 538398 285914 538634
rect 285294 502954 285914 538398
rect 285294 502718 285326 502954
rect 285562 502718 285646 502954
rect 285882 502718 285914 502954
rect 285294 502634 285914 502718
rect 285294 502398 285326 502634
rect 285562 502398 285646 502634
rect 285882 502398 285914 502634
rect 285294 466954 285914 502398
rect 285294 466718 285326 466954
rect 285562 466718 285646 466954
rect 285882 466718 285914 466954
rect 285294 466634 285914 466718
rect 285294 466398 285326 466634
rect 285562 466398 285646 466634
rect 285882 466398 285914 466634
rect 285294 430954 285914 466398
rect 285294 430718 285326 430954
rect 285562 430718 285646 430954
rect 285882 430718 285914 430954
rect 285294 430634 285914 430718
rect 285294 430398 285326 430634
rect 285562 430398 285646 430634
rect 285882 430398 285914 430634
rect 285294 394954 285914 430398
rect 285294 394718 285326 394954
rect 285562 394718 285646 394954
rect 285882 394718 285914 394954
rect 285294 394634 285914 394718
rect 285294 394398 285326 394634
rect 285562 394398 285646 394634
rect 285882 394398 285914 394634
rect 285294 358954 285914 394398
rect 285294 358718 285326 358954
rect 285562 358718 285646 358954
rect 285882 358718 285914 358954
rect 285294 358634 285914 358718
rect 285294 358398 285326 358634
rect 285562 358398 285646 358634
rect 285882 358398 285914 358634
rect 285294 322954 285914 358398
rect 285294 322718 285326 322954
rect 285562 322718 285646 322954
rect 285882 322718 285914 322954
rect 285294 322634 285914 322718
rect 285294 322398 285326 322634
rect 285562 322398 285646 322634
rect 285882 322398 285914 322634
rect 285294 286954 285914 322398
rect 285294 286718 285326 286954
rect 285562 286718 285646 286954
rect 285882 286718 285914 286954
rect 285294 286634 285914 286718
rect 285294 286398 285326 286634
rect 285562 286398 285646 286634
rect 285882 286398 285914 286634
rect 285294 250954 285914 286398
rect 285294 250718 285326 250954
rect 285562 250718 285646 250954
rect 285882 250718 285914 250954
rect 285294 250634 285914 250718
rect 285294 250398 285326 250634
rect 285562 250398 285646 250634
rect 285882 250398 285914 250634
rect 285294 214954 285914 250398
rect 285294 214718 285326 214954
rect 285562 214718 285646 214954
rect 285882 214718 285914 214954
rect 285294 214634 285914 214718
rect 285294 214398 285326 214634
rect 285562 214398 285646 214634
rect 285882 214398 285914 214634
rect 285294 178954 285914 214398
rect 285294 178718 285326 178954
rect 285562 178718 285646 178954
rect 285882 178718 285914 178954
rect 285294 178634 285914 178718
rect 285294 178398 285326 178634
rect 285562 178398 285646 178634
rect 285882 178398 285914 178634
rect 285294 142954 285914 178398
rect 285294 142718 285326 142954
rect 285562 142718 285646 142954
rect 285882 142718 285914 142954
rect 285294 142634 285914 142718
rect 285294 142398 285326 142634
rect 285562 142398 285646 142634
rect 285882 142398 285914 142634
rect 285294 106954 285914 142398
rect 285294 106718 285326 106954
rect 285562 106718 285646 106954
rect 285882 106718 285914 106954
rect 285294 106634 285914 106718
rect 285294 106398 285326 106634
rect 285562 106398 285646 106634
rect 285882 106398 285914 106634
rect 285294 70954 285914 106398
rect 285294 70718 285326 70954
rect 285562 70718 285646 70954
rect 285882 70718 285914 70954
rect 285294 70634 285914 70718
rect 285294 70398 285326 70634
rect 285562 70398 285646 70634
rect 285882 70398 285914 70634
rect 285294 34954 285914 70398
rect 285294 34718 285326 34954
rect 285562 34718 285646 34954
rect 285882 34718 285914 34954
rect 285294 34634 285914 34718
rect 285294 34398 285326 34634
rect 285562 34398 285646 34634
rect 285882 34398 285914 34634
rect 285294 -7066 285914 34398
rect 285294 -7302 285326 -7066
rect 285562 -7302 285646 -7066
rect 285882 -7302 285914 -7066
rect 285294 -7386 285914 -7302
rect 285294 -7622 285326 -7386
rect 285562 -7622 285646 -7386
rect 285882 -7622 285914 -7386
rect 285294 -7654 285914 -7622
rect 289794 704838 290414 711590
rect 289794 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 290414 704838
rect 289794 704518 290414 704602
rect 289794 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 290414 704518
rect 289794 687454 290414 704282
rect 289794 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 290414 687454
rect 289794 687134 290414 687218
rect 289794 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 290414 687134
rect 289794 651454 290414 686898
rect 289794 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 290414 651454
rect 289794 651134 290414 651218
rect 289794 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 290414 651134
rect 289794 615454 290414 650898
rect 289794 615218 289826 615454
rect 290062 615218 290146 615454
rect 290382 615218 290414 615454
rect 289794 615134 290414 615218
rect 289794 614898 289826 615134
rect 290062 614898 290146 615134
rect 290382 614898 290414 615134
rect 289794 579454 290414 614898
rect 289794 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 290414 579454
rect 289794 579134 290414 579218
rect 289794 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 290414 579134
rect 289794 543454 290414 578898
rect 289794 543218 289826 543454
rect 290062 543218 290146 543454
rect 290382 543218 290414 543454
rect 289794 543134 290414 543218
rect 289794 542898 289826 543134
rect 290062 542898 290146 543134
rect 290382 542898 290414 543134
rect 289794 507454 290414 542898
rect 289794 507218 289826 507454
rect 290062 507218 290146 507454
rect 290382 507218 290414 507454
rect 289794 507134 290414 507218
rect 289794 506898 289826 507134
rect 290062 506898 290146 507134
rect 290382 506898 290414 507134
rect 289794 471454 290414 506898
rect 289794 471218 289826 471454
rect 290062 471218 290146 471454
rect 290382 471218 290414 471454
rect 289794 471134 290414 471218
rect 289794 470898 289826 471134
rect 290062 470898 290146 471134
rect 290382 470898 290414 471134
rect 289794 435454 290414 470898
rect 289794 435218 289826 435454
rect 290062 435218 290146 435454
rect 290382 435218 290414 435454
rect 289794 435134 290414 435218
rect 289794 434898 289826 435134
rect 290062 434898 290146 435134
rect 290382 434898 290414 435134
rect 289794 399454 290414 434898
rect 289794 399218 289826 399454
rect 290062 399218 290146 399454
rect 290382 399218 290414 399454
rect 289794 399134 290414 399218
rect 289794 398898 289826 399134
rect 290062 398898 290146 399134
rect 290382 398898 290414 399134
rect 289794 363454 290414 398898
rect 289794 363218 289826 363454
rect 290062 363218 290146 363454
rect 290382 363218 290414 363454
rect 289794 363134 290414 363218
rect 289794 362898 289826 363134
rect 290062 362898 290146 363134
rect 290382 362898 290414 363134
rect 289794 327454 290414 362898
rect 289794 327218 289826 327454
rect 290062 327218 290146 327454
rect 290382 327218 290414 327454
rect 289794 327134 290414 327218
rect 289794 326898 289826 327134
rect 290062 326898 290146 327134
rect 290382 326898 290414 327134
rect 289794 291454 290414 326898
rect 289794 291218 289826 291454
rect 290062 291218 290146 291454
rect 290382 291218 290414 291454
rect 289794 291134 290414 291218
rect 289794 290898 289826 291134
rect 290062 290898 290146 291134
rect 290382 290898 290414 291134
rect 289794 255454 290414 290898
rect 289794 255218 289826 255454
rect 290062 255218 290146 255454
rect 290382 255218 290414 255454
rect 289794 255134 290414 255218
rect 289794 254898 289826 255134
rect 290062 254898 290146 255134
rect 290382 254898 290414 255134
rect 289794 219454 290414 254898
rect 289794 219218 289826 219454
rect 290062 219218 290146 219454
rect 290382 219218 290414 219454
rect 289794 219134 290414 219218
rect 289794 218898 289826 219134
rect 290062 218898 290146 219134
rect 290382 218898 290414 219134
rect 289794 183454 290414 218898
rect 289794 183218 289826 183454
rect 290062 183218 290146 183454
rect 290382 183218 290414 183454
rect 289794 183134 290414 183218
rect 289794 182898 289826 183134
rect 290062 182898 290146 183134
rect 290382 182898 290414 183134
rect 289794 147454 290414 182898
rect 289794 147218 289826 147454
rect 290062 147218 290146 147454
rect 290382 147218 290414 147454
rect 289794 147134 290414 147218
rect 289794 146898 289826 147134
rect 290062 146898 290146 147134
rect 290382 146898 290414 147134
rect 289794 111454 290414 146898
rect 289794 111218 289826 111454
rect 290062 111218 290146 111454
rect 290382 111218 290414 111454
rect 289794 111134 290414 111218
rect 289794 110898 289826 111134
rect 290062 110898 290146 111134
rect 290382 110898 290414 111134
rect 289794 75454 290414 110898
rect 289794 75218 289826 75454
rect 290062 75218 290146 75454
rect 290382 75218 290414 75454
rect 289794 75134 290414 75218
rect 289794 74898 289826 75134
rect 290062 74898 290146 75134
rect 290382 74898 290414 75134
rect 289794 39454 290414 74898
rect 289794 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 290414 39454
rect 289794 39134 290414 39218
rect 289794 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 290414 39134
rect 289794 3454 290414 38898
rect 289794 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 290414 3454
rect 289794 3134 290414 3218
rect 289794 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 290414 3134
rect 289794 -346 290414 2898
rect 289794 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 290414 -346
rect 289794 -666 290414 -582
rect 289794 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 290414 -666
rect 289794 -7654 290414 -902
rect 294294 705798 294914 711590
rect 294294 705562 294326 705798
rect 294562 705562 294646 705798
rect 294882 705562 294914 705798
rect 294294 705478 294914 705562
rect 294294 705242 294326 705478
rect 294562 705242 294646 705478
rect 294882 705242 294914 705478
rect 294294 691954 294914 705242
rect 294294 691718 294326 691954
rect 294562 691718 294646 691954
rect 294882 691718 294914 691954
rect 294294 691634 294914 691718
rect 294294 691398 294326 691634
rect 294562 691398 294646 691634
rect 294882 691398 294914 691634
rect 294294 655954 294914 691398
rect 294294 655718 294326 655954
rect 294562 655718 294646 655954
rect 294882 655718 294914 655954
rect 294294 655634 294914 655718
rect 294294 655398 294326 655634
rect 294562 655398 294646 655634
rect 294882 655398 294914 655634
rect 294294 619954 294914 655398
rect 294294 619718 294326 619954
rect 294562 619718 294646 619954
rect 294882 619718 294914 619954
rect 294294 619634 294914 619718
rect 294294 619398 294326 619634
rect 294562 619398 294646 619634
rect 294882 619398 294914 619634
rect 294294 583954 294914 619398
rect 294294 583718 294326 583954
rect 294562 583718 294646 583954
rect 294882 583718 294914 583954
rect 294294 583634 294914 583718
rect 294294 583398 294326 583634
rect 294562 583398 294646 583634
rect 294882 583398 294914 583634
rect 294294 547954 294914 583398
rect 294294 547718 294326 547954
rect 294562 547718 294646 547954
rect 294882 547718 294914 547954
rect 294294 547634 294914 547718
rect 294294 547398 294326 547634
rect 294562 547398 294646 547634
rect 294882 547398 294914 547634
rect 294294 511954 294914 547398
rect 294294 511718 294326 511954
rect 294562 511718 294646 511954
rect 294882 511718 294914 511954
rect 294294 511634 294914 511718
rect 294294 511398 294326 511634
rect 294562 511398 294646 511634
rect 294882 511398 294914 511634
rect 294294 475954 294914 511398
rect 294294 475718 294326 475954
rect 294562 475718 294646 475954
rect 294882 475718 294914 475954
rect 294294 475634 294914 475718
rect 294294 475398 294326 475634
rect 294562 475398 294646 475634
rect 294882 475398 294914 475634
rect 294294 439954 294914 475398
rect 294294 439718 294326 439954
rect 294562 439718 294646 439954
rect 294882 439718 294914 439954
rect 294294 439634 294914 439718
rect 294294 439398 294326 439634
rect 294562 439398 294646 439634
rect 294882 439398 294914 439634
rect 294294 403954 294914 439398
rect 294294 403718 294326 403954
rect 294562 403718 294646 403954
rect 294882 403718 294914 403954
rect 294294 403634 294914 403718
rect 294294 403398 294326 403634
rect 294562 403398 294646 403634
rect 294882 403398 294914 403634
rect 294294 367954 294914 403398
rect 294294 367718 294326 367954
rect 294562 367718 294646 367954
rect 294882 367718 294914 367954
rect 294294 367634 294914 367718
rect 294294 367398 294326 367634
rect 294562 367398 294646 367634
rect 294882 367398 294914 367634
rect 294294 331954 294914 367398
rect 294294 331718 294326 331954
rect 294562 331718 294646 331954
rect 294882 331718 294914 331954
rect 294294 331634 294914 331718
rect 294294 331398 294326 331634
rect 294562 331398 294646 331634
rect 294882 331398 294914 331634
rect 294294 295954 294914 331398
rect 294294 295718 294326 295954
rect 294562 295718 294646 295954
rect 294882 295718 294914 295954
rect 294294 295634 294914 295718
rect 294294 295398 294326 295634
rect 294562 295398 294646 295634
rect 294882 295398 294914 295634
rect 294294 259954 294914 295398
rect 294294 259718 294326 259954
rect 294562 259718 294646 259954
rect 294882 259718 294914 259954
rect 294294 259634 294914 259718
rect 294294 259398 294326 259634
rect 294562 259398 294646 259634
rect 294882 259398 294914 259634
rect 294294 223954 294914 259398
rect 294294 223718 294326 223954
rect 294562 223718 294646 223954
rect 294882 223718 294914 223954
rect 294294 223634 294914 223718
rect 294294 223398 294326 223634
rect 294562 223398 294646 223634
rect 294882 223398 294914 223634
rect 294294 187954 294914 223398
rect 294294 187718 294326 187954
rect 294562 187718 294646 187954
rect 294882 187718 294914 187954
rect 294294 187634 294914 187718
rect 294294 187398 294326 187634
rect 294562 187398 294646 187634
rect 294882 187398 294914 187634
rect 294294 151954 294914 187398
rect 294294 151718 294326 151954
rect 294562 151718 294646 151954
rect 294882 151718 294914 151954
rect 294294 151634 294914 151718
rect 294294 151398 294326 151634
rect 294562 151398 294646 151634
rect 294882 151398 294914 151634
rect 294294 115954 294914 151398
rect 294294 115718 294326 115954
rect 294562 115718 294646 115954
rect 294882 115718 294914 115954
rect 294294 115634 294914 115718
rect 294294 115398 294326 115634
rect 294562 115398 294646 115634
rect 294882 115398 294914 115634
rect 294294 79954 294914 115398
rect 294294 79718 294326 79954
rect 294562 79718 294646 79954
rect 294882 79718 294914 79954
rect 294294 79634 294914 79718
rect 294294 79398 294326 79634
rect 294562 79398 294646 79634
rect 294882 79398 294914 79634
rect 294294 43954 294914 79398
rect 294294 43718 294326 43954
rect 294562 43718 294646 43954
rect 294882 43718 294914 43954
rect 294294 43634 294914 43718
rect 294294 43398 294326 43634
rect 294562 43398 294646 43634
rect 294882 43398 294914 43634
rect 294294 7954 294914 43398
rect 294294 7718 294326 7954
rect 294562 7718 294646 7954
rect 294882 7718 294914 7954
rect 294294 7634 294914 7718
rect 294294 7398 294326 7634
rect 294562 7398 294646 7634
rect 294882 7398 294914 7634
rect 294294 -1306 294914 7398
rect 294294 -1542 294326 -1306
rect 294562 -1542 294646 -1306
rect 294882 -1542 294914 -1306
rect 294294 -1626 294914 -1542
rect 294294 -1862 294326 -1626
rect 294562 -1862 294646 -1626
rect 294882 -1862 294914 -1626
rect 294294 -7654 294914 -1862
rect 298794 706758 299414 711590
rect 298794 706522 298826 706758
rect 299062 706522 299146 706758
rect 299382 706522 299414 706758
rect 298794 706438 299414 706522
rect 298794 706202 298826 706438
rect 299062 706202 299146 706438
rect 299382 706202 299414 706438
rect 298794 696454 299414 706202
rect 298794 696218 298826 696454
rect 299062 696218 299146 696454
rect 299382 696218 299414 696454
rect 298794 696134 299414 696218
rect 298794 695898 298826 696134
rect 299062 695898 299146 696134
rect 299382 695898 299414 696134
rect 298794 660454 299414 695898
rect 298794 660218 298826 660454
rect 299062 660218 299146 660454
rect 299382 660218 299414 660454
rect 298794 660134 299414 660218
rect 298794 659898 298826 660134
rect 299062 659898 299146 660134
rect 299382 659898 299414 660134
rect 298794 624454 299414 659898
rect 298794 624218 298826 624454
rect 299062 624218 299146 624454
rect 299382 624218 299414 624454
rect 298794 624134 299414 624218
rect 298794 623898 298826 624134
rect 299062 623898 299146 624134
rect 299382 623898 299414 624134
rect 298794 588454 299414 623898
rect 298794 588218 298826 588454
rect 299062 588218 299146 588454
rect 299382 588218 299414 588454
rect 298794 588134 299414 588218
rect 298794 587898 298826 588134
rect 299062 587898 299146 588134
rect 299382 587898 299414 588134
rect 298794 552454 299414 587898
rect 298794 552218 298826 552454
rect 299062 552218 299146 552454
rect 299382 552218 299414 552454
rect 298794 552134 299414 552218
rect 298794 551898 298826 552134
rect 299062 551898 299146 552134
rect 299382 551898 299414 552134
rect 298794 516454 299414 551898
rect 298794 516218 298826 516454
rect 299062 516218 299146 516454
rect 299382 516218 299414 516454
rect 298794 516134 299414 516218
rect 298794 515898 298826 516134
rect 299062 515898 299146 516134
rect 299382 515898 299414 516134
rect 298794 480454 299414 515898
rect 298794 480218 298826 480454
rect 299062 480218 299146 480454
rect 299382 480218 299414 480454
rect 298794 480134 299414 480218
rect 298794 479898 298826 480134
rect 299062 479898 299146 480134
rect 299382 479898 299414 480134
rect 298794 444454 299414 479898
rect 298794 444218 298826 444454
rect 299062 444218 299146 444454
rect 299382 444218 299414 444454
rect 298794 444134 299414 444218
rect 298794 443898 298826 444134
rect 299062 443898 299146 444134
rect 299382 443898 299414 444134
rect 298794 408454 299414 443898
rect 298794 408218 298826 408454
rect 299062 408218 299146 408454
rect 299382 408218 299414 408454
rect 298794 408134 299414 408218
rect 298794 407898 298826 408134
rect 299062 407898 299146 408134
rect 299382 407898 299414 408134
rect 298794 372454 299414 407898
rect 298794 372218 298826 372454
rect 299062 372218 299146 372454
rect 299382 372218 299414 372454
rect 298794 372134 299414 372218
rect 298794 371898 298826 372134
rect 299062 371898 299146 372134
rect 299382 371898 299414 372134
rect 298794 336454 299414 371898
rect 298794 336218 298826 336454
rect 299062 336218 299146 336454
rect 299382 336218 299414 336454
rect 298794 336134 299414 336218
rect 298794 335898 298826 336134
rect 299062 335898 299146 336134
rect 299382 335898 299414 336134
rect 298794 300454 299414 335898
rect 298794 300218 298826 300454
rect 299062 300218 299146 300454
rect 299382 300218 299414 300454
rect 298794 300134 299414 300218
rect 298794 299898 298826 300134
rect 299062 299898 299146 300134
rect 299382 299898 299414 300134
rect 298794 264454 299414 299898
rect 298794 264218 298826 264454
rect 299062 264218 299146 264454
rect 299382 264218 299414 264454
rect 298794 264134 299414 264218
rect 298794 263898 298826 264134
rect 299062 263898 299146 264134
rect 299382 263898 299414 264134
rect 298794 228454 299414 263898
rect 298794 228218 298826 228454
rect 299062 228218 299146 228454
rect 299382 228218 299414 228454
rect 298794 228134 299414 228218
rect 298794 227898 298826 228134
rect 299062 227898 299146 228134
rect 299382 227898 299414 228134
rect 298794 192454 299414 227898
rect 298794 192218 298826 192454
rect 299062 192218 299146 192454
rect 299382 192218 299414 192454
rect 298794 192134 299414 192218
rect 298794 191898 298826 192134
rect 299062 191898 299146 192134
rect 299382 191898 299414 192134
rect 298794 156454 299414 191898
rect 298794 156218 298826 156454
rect 299062 156218 299146 156454
rect 299382 156218 299414 156454
rect 298794 156134 299414 156218
rect 298794 155898 298826 156134
rect 299062 155898 299146 156134
rect 299382 155898 299414 156134
rect 298794 120454 299414 155898
rect 298794 120218 298826 120454
rect 299062 120218 299146 120454
rect 299382 120218 299414 120454
rect 298794 120134 299414 120218
rect 298794 119898 298826 120134
rect 299062 119898 299146 120134
rect 299382 119898 299414 120134
rect 298794 84454 299414 119898
rect 298794 84218 298826 84454
rect 299062 84218 299146 84454
rect 299382 84218 299414 84454
rect 298794 84134 299414 84218
rect 298794 83898 298826 84134
rect 299062 83898 299146 84134
rect 299382 83898 299414 84134
rect 298794 48454 299414 83898
rect 298794 48218 298826 48454
rect 299062 48218 299146 48454
rect 299382 48218 299414 48454
rect 298794 48134 299414 48218
rect 298794 47898 298826 48134
rect 299062 47898 299146 48134
rect 299382 47898 299414 48134
rect 298794 12454 299414 47898
rect 298794 12218 298826 12454
rect 299062 12218 299146 12454
rect 299382 12218 299414 12454
rect 298794 12134 299414 12218
rect 298794 11898 298826 12134
rect 299062 11898 299146 12134
rect 299382 11898 299414 12134
rect 298794 -2266 299414 11898
rect 298794 -2502 298826 -2266
rect 299062 -2502 299146 -2266
rect 299382 -2502 299414 -2266
rect 298794 -2586 299414 -2502
rect 298794 -2822 298826 -2586
rect 299062 -2822 299146 -2586
rect 299382 -2822 299414 -2586
rect 298794 -7654 299414 -2822
rect 303294 707718 303914 711590
rect 303294 707482 303326 707718
rect 303562 707482 303646 707718
rect 303882 707482 303914 707718
rect 303294 707398 303914 707482
rect 303294 707162 303326 707398
rect 303562 707162 303646 707398
rect 303882 707162 303914 707398
rect 303294 700954 303914 707162
rect 303294 700718 303326 700954
rect 303562 700718 303646 700954
rect 303882 700718 303914 700954
rect 303294 700634 303914 700718
rect 303294 700398 303326 700634
rect 303562 700398 303646 700634
rect 303882 700398 303914 700634
rect 303294 664954 303914 700398
rect 303294 664718 303326 664954
rect 303562 664718 303646 664954
rect 303882 664718 303914 664954
rect 303294 664634 303914 664718
rect 303294 664398 303326 664634
rect 303562 664398 303646 664634
rect 303882 664398 303914 664634
rect 303294 628954 303914 664398
rect 303294 628718 303326 628954
rect 303562 628718 303646 628954
rect 303882 628718 303914 628954
rect 303294 628634 303914 628718
rect 303294 628398 303326 628634
rect 303562 628398 303646 628634
rect 303882 628398 303914 628634
rect 303294 592954 303914 628398
rect 303294 592718 303326 592954
rect 303562 592718 303646 592954
rect 303882 592718 303914 592954
rect 303294 592634 303914 592718
rect 303294 592398 303326 592634
rect 303562 592398 303646 592634
rect 303882 592398 303914 592634
rect 303294 556954 303914 592398
rect 303294 556718 303326 556954
rect 303562 556718 303646 556954
rect 303882 556718 303914 556954
rect 303294 556634 303914 556718
rect 303294 556398 303326 556634
rect 303562 556398 303646 556634
rect 303882 556398 303914 556634
rect 303294 520954 303914 556398
rect 303294 520718 303326 520954
rect 303562 520718 303646 520954
rect 303882 520718 303914 520954
rect 303294 520634 303914 520718
rect 303294 520398 303326 520634
rect 303562 520398 303646 520634
rect 303882 520398 303914 520634
rect 303294 484954 303914 520398
rect 303294 484718 303326 484954
rect 303562 484718 303646 484954
rect 303882 484718 303914 484954
rect 303294 484634 303914 484718
rect 303294 484398 303326 484634
rect 303562 484398 303646 484634
rect 303882 484398 303914 484634
rect 303294 448954 303914 484398
rect 303294 448718 303326 448954
rect 303562 448718 303646 448954
rect 303882 448718 303914 448954
rect 303294 448634 303914 448718
rect 303294 448398 303326 448634
rect 303562 448398 303646 448634
rect 303882 448398 303914 448634
rect 303294 412954 303914 448398
rect 303294 412718 303326 412954
rect 303562 412718 303646 412954
rect 303882 412718 303914 412954
rect 303294 412634 303914 412718
rect 303294 412398 303326 412634
rect 303562 412398 303646 412634
rect 303882 412398 303914 412634
rect 303294 376954 303914 412398
rect 303294 376718 303326 376954
rect 303562 376718 303646 376954
rect 303882 376718 303914 376954
rect 303294 376634 303914 376718
rect 303294 376398 303326 376634
rect 303562 376398 303646 376634
rect 303882 376398 303914 376634
rect 303294 340954 303914 376398
rect 303294 340718 303326 340954
rect 303562 340718 303646 340954
rect 303882 340718 303914 340954
rect 303294 340634 303914 340718
rect 303294 340398 303326 340634
rect 303562 340398 303646 340634
rect 303882 340398 303914 340634
rect 303294 304954 303914 340398
rect 303294 304718 303326 304954
rect 303562 304718 303646 304954
rect 303882 304718 303914 304954
rect 303294 304634 303914 304718
rect 303294 304398 303326 304634
rect 303562 304398 303646 304634
rect 303882 304398 303914 304634
rect 303294 268954 303914 304398
rect 303294 268718 303326 268954
rect 303562 268718 303646 268954
rect 303882 268718 303914 268954
rect 303294 268634 303914 268718
rect 303294 268398 303326 268634
rect 303562 268398 303646 268634
rect 303882 268398 303914 268634
rect 303294 232954 303914 268398
rect 303294 232718 303326 232954
rect 303562 232718 303646 232954
rect 303882 232718 303914 232954
rect 303294 232634 303914 232718
rect 303294 232398 303326 232634
rect 303562 232398 303646 232634
rect 303882 232398 303914 232634
rect 303294 196954 303914 232398
rect 303294 196718 303326 196954
rect 303562 196718 303646 196954
rect 303882 196718 303914 196954
rect 303294 196634 303914 196718
rect 303294 196398 303326 196634
rect 303562 196398 303646 196634
rect 303882 196398 303914 196634
rect 303294 160954 303914 196398
rect 303294 160718 303326 160954
rect 303562 160718 303646 160954
rect 303882 160718 303914 160954
rect 303294 160634 303914 160718
rect 303294 160398 303326 160634
rect 303562 160398 303646 160634
rect 303882 160398 303914 160634
rect 303294 124954 303914 160398
rect 303294 124718 303326 124954
rect 303562 124718 303646 124954
rect 303882 124718 303914 124954
rect 303294 124634 303914 124718
rect 303294 124398 303326 124634
rect 303562 124398 303646 124634
rect 303882 124398 303914 124634
rect 303294 88954 303914 124398
rect 303294 88718 303326 88954
rect 303562 88718 303646 88954
rect 303882 88718 303914 88954
rect 303294 88634 303914 88718
rect 303294 88398 303326 88634
rect 303562 88398 303646 88634
rect 303882 88398 303914 88634
rect 303294 52954 303914 88398
rect 303294 52718 303326 52954
rect 303562 52718 303646 52954
rect 303882 52718 303914 52954
rect 303294 52634 303914 52718
rect 303294 52398 303326 52634
rect 303562 52398 303646 52634
rect 303882 52398 303914 52634
rect 303294 16954 303914 52398
rect 303294 16718 303326 16954
rect 303562 16718 303646 16954
rect 303882 16718 303914 16954
rect 303294 16634 303914 16718
rect 303294 16398 303326 16634
rect 303562 16398 303646 16634
rect 303882 16398 303914 16634
rect 303294 -3226 303914 16398
rect 303294 -3462 303326 -3226
rect 303562 -3462 303646 -3226
rect 303882 -3462 303914 -3226
rect 303294 -3546 303914 -3462
rect 303294 -3782 303326 -3546
rect 303562 -3782 303646 -3546
rect 303882 -3782 303914 -3546
rect 303294 -7654 303914 -3782
rect 307794 708678 308414 711590
rect 307794 708442 307826 708678
rect 308062 708442 308146 708678
rect 308382 708442 308414 708678
rect 307794 708358 308414 708442
rect 307794 708122 307826 708358
rect 308062 708122 308146 708358
rect 308382 708122 308414 708358
rect 307794 669454 308414 708122
rect 307794 669218 307826 669454
rect 308062 669218 308146 669454
rect 308382 669218 308414 669454
rect 307794 669134 308414 669218
rect 307794 668898 307826 669134
rect 308062 668898 308146 669134
rect 308382 668898 308414 669134
rect 307794 633454 308414 668898
rect 307794 633218 307826 633454
rect 308062 633218 308146 633454
rect 308382 633218 308414 633454
rect 307794 633134 308414 633218
rect 307794 632898 307826 633134
rect 308062 632898 308146 633134
rect 308382 632898 308414 633134
rect 307794 597454 308414 632898
rect 307794 597218 307826 597454
rect 308062 597218 308146 597454
rect 308382 597218 308414 597454
rect 307794 597134 308414 597218
rect 307794 596898 307826 597134
rect 308062 596898 308146 597134
rect 308382 596898 308414 597134
rect 307794 561454 308414 596898
rect 307794 561218 307826 561454
rect 308062 561218 308146 561454
rect 308382 561218 308414 561454
rect 307794 561134 308414 561218
rect 307794 560898 307826 561134
rect 308062 560898 308146 561134
rect 308382 560898 308414 561134
rect 307794 525454 308414 560898
rect 307794 525218 307826 525454
rect 308062 525218 308146 525454
rect 308382 525218 308414 525454
rect 307794 525134 308414 525218
rect 307794 524898 307826 525134
rect 308062 524898 308146 525134
rect 308382 524898 308414 525134
rect 307794 489454 308414 524898
rect 307794 489218 307826 489454
rect 308062 489218 308146 489454
rect 308382 489218 308414 489454
rect 307794 489134 308414 489218
rect 307794 488898 307826 489134
rect 308062 488898 308146 489134
rect 308382 488898 308414 489134
rect 307794 453454 308414 488898
rect 307794 453218 307826 453454
rect 308062 453218 308146 453454
rect 308382 453218 308414 453454
rect 307794 453134 308414 453218
rect 307794 452898 307826 453134
rect 308062 452898 308146 453134
rect 308382 452898 308414 453134
rect 307794 417454 308414 452898
rect 307794 417218 307826 417454
rect 308062 417218 308146 417454
rect 308382 417218 308414 417454
rect 307794 417134 308414 417218
rect 307794 416898 307826 417134
rect 308062 416898 308146 417134
rect 308382 416898 308414 417134
rect 307794 381454 308414 416898
rect 307794 381218 307826 381454
rect 308062 381218 308146 381454
rect 308382 381218 308414 381454
rect 307794 381134 308414 381218
rect 307794 380898 307826 381134
rect 308062 380898 308146 381134
rect 308382 380898 308414 381134
rect 307794 345454 308414 380898
rect 307794 345218 307826 345454
rect 308062 345218 308146 345454
rect 308382 345218 308414 345454
rect 307794 345134 308414 345218
rect 307794 344898 307826 345134
rect 308062 344898 308146 345134
rect 308382 344898 308414 345134
rect 307794 309454 308414 344898
rect 307794 309218 307826 309454
rect 308062 309218 308146 309454
rect 308382 309218 308414 309454
rect 307794 309134 308414 309218
rect 307794 308898 307826 309134
rect 308062 308898 308146 309134
rect 308382 308898 308414 309134
rect 307794 273454 308414 308898
rect 307794 273218 307826 273454
rect 308062 273218 308146 273454
rect 308382 273218 308414 273454
rect 307794 273134 308414 273218
rect 307794 272898 307826 273134
rect 308062 272898 308146 273134
rect 308382 272898 308414 273134
rect 307794 237454 308414 272898
rect 307794 237218 307826 237454
rect 308062 237218 308146 237454
rect 308382 237218 308414 237454
rect 307794 237134 308414 237218
rect 307794 236898 307826 237134
rect 308062 236898 308146 237134
rect 308382 236898 308414 237134
rect 307794 201454 308414 236898
rect 307794 201218 307826 201454
rect 308062 201218 308146 201454
rect 308382 201218 308414 201454
rect 307794 201134 308414 201218
rect 307794 200898 307826 201134
rect 308062 200898 308146 201134
rect 308382 200898 308414 201134
rect 307794 165454 308414 200898
rect 307794 165218 307826 165454
rect 308062 165218 308146 165454
rect 308382 165218 308414 165454
rect 307794 165134 308414 165218
rect 307794 164898 307826 165134
rect 308062 164898 308146 165134
rect 308382 164898 308414 165134
rect 307794 129454 308414 164898
rect 307794 129218 307826 129454
rect 308062 129218 308146 129454
rect 308382 129218 308414 129454
rect 307794 129134 308414 129218
rect 307794 128898 307826 129134
rect 308062 128898 308146 129134
rect 308382 128898 308414 129134
rect 307794 93454 308414 128898
rect 307794 93218 307826 93454
rect 308062 93218 308146 93454
rect 308382 93218 308414 93454
rect 307794 93134 308414 93218
rect 307794 92898 307826 93134
rect 308062 92898 308146 93134
rect 308382 92898 308414 93134
rect 307794 57454 308414 92898
rect 307794 57218 307826 57454
rect 308062 57218 308146 57454
rect 308382 57218 308414 57454
rect 307794 57134 308414 57218
rect 307794 56898 307826 57134
rect 308062 56898 308146 57134
rect 308382 56898 308414 57134
rect 307794 21454 308414 56898
rect 307794 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 308414 21454
rect 307794 21134 308414 21218
rect 307794 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 308414 21134
rect 307794 -4186 308414 20898
rect 307794 -4422 307826 -4186
rect 308062 -4422 308146 -4186
rect 308382 -4422 308414 -4186
rect 307794 -4506 308414 -4422
rect 307794 -4742 307826 -4506
rect 308062 -4742 308146 -4506
rect 308382 -4742 308414 -4506
rect 307794 -7654 308414 -4742
rect 312294 709638 312914 711590
rect 312294 709402 312326 709638
rect 312562 709402 312646 709638
rect 312882 709402 312914 709638
rect 312294 709318 312914 709402
rect 312294 709082 312326 709318
rect 312562 709082 312646 709318
rect 312882 709082 312914 709318
rect 312294 673954 312914 709082
rect 312294 673718 312326 673954
rect 312562 673718 312646 673954
rect 312882 673718 312914 673954
rect 312294 673634 312914 673718
rect 312294 673398 312326 673634
rect 312562 673398 312646 673634
rect 312882 673398 312914 673634
rect 312294 637954 312914 673398
rect 312294 637718 312326 637954
rect 312562 637718 312646 637954
rect 312882 637718 312914 637954
rect 312294 637634 312914 637718
rect 312294 637398 312326 637634
rect 312562 637398 312646 637634
rect 312882 637398 312914 637634
rect 312294 601954 312914 637398
rect 312294 601718 312326 601954
rect 312562 601718 312646 601954
rect 312882 601718 312914 601954
rect 312294 601634 312914 601718
rect 312294 601398 312326 601634
rect 312562 601398 312646 601634
rect 312882 601398 312914 601634
rect 312294 565954 312914 601398
rect 312294 565718 312326 565954
rect 312562 565718 312646 565954
rect 312882 565718 312914 565954
rect 312294 565634 312914 565718
rect 312294 565398 312326 565634
rect 312562 565398 312646 565634
rect 312882 565398 312914 565634
rect 312294 529954 312914 565398
rect 312294 529718 312326 529954
rect 312562 529718 312646 529954
rect 312882 529718 312914 529954
rect 312294 529634 312914 529718
rect 312294 529398 312326 529634
rect 312562 529398 312646 529634
rect 312882 529398 312914 529634
rect 312294 493954 312914 529398
rect 312294 493718 312326 493954
rect 312562 493718 312646 493954
rect 312882 493718 312914 493954
rect 312294 493634 312914 493718
rect 312294 493398 312326 493634
rect 312562 493398 312646 493634
rect 312882 493398 312914 493634
rect 312294 457954 312914 493398
rect 312294 457718 312326 457954
rect 312562 457718 312646 457954
rect 312882 457718 312914 457954
rect 312294 457634 312914 457718
rect 312294 457398 312326 457634
rect 312562 457398 312646 457634
rect 312882 457398 312914 457634
rect 312294 421954 312914 457398
rect 312294 421718 312326 421954
rect 312562 421718 312646 421954
rect 312882 421718 312914 421954
rect 312294 421634 312914 421718
rect 312294 421398 312326 421634
rect 312562 421398 312646 421634
rect 312882 421398 312914 421634
rect 312294 385954 312914 421398
rect 312294 385718 312326 385954
rect 312562 385718 312646 385954
rect 312882 385718 312914 385954
rect 312294 385634 312914 385718
rect 312294 385398 312326 385634
rect 312562 385398 312646 385634
rect 312882 385398 312914 385634
rect 312294 349954 312914 385398
rect 312294 349718 312326 349954
rect 312562 349718 312646 349954
rect 312882 349718 312914 349954
rect 312294 349634 312914 349718
rect 312294 349398 312326 349634
rect 312562 349398 312646 349634
rect 312882 349398 312914 349634
rect 312294 313954 312914 349398
rect 312294 313718 312326 313954
rect 312562 313718 312646 313954
rect 312882 313718 312914 313954
rect 312294 313634 312914 313718
rect 312294 313398 312326 313634
rect 312562 313398 312646 313634
rect 312882 313398 312914 313634
rect 312294 277954 312914 313398
rect 312294 277718 312326 277954
rect 312562 277718 312646 277954
rect 312882 277718 312914 277954
rect 312294 277634 312914 277718
rect 312294 277398 312326 277634
rect 312562 277398 312646 277634
rect 312882 277398 312914 277634
rect 312294 241954 312914 277398
rect 312294 241718 312326 241954
rect 312562 241718 312646 241954
rect 312882 241718 312914 241954
rect 312294 241634 312914 241718
rect 312294 241398 312326 241634
rect 312562 241398 312646 241634
rect 312882 241398 312914 241634
rect 312294 205954 312914 241398
rect 312294 205718 312326 205954
rect 312562 205718 312646 205954
rect 312882 205718 312914 205954
rect 312294 205634 312914 205718
rect 312294 205398 312326 205634
rect 312562 205398 312646 205634
rect 312882 205398 312914 205634
rect 312294 169954 312914 205398
rect 312294 169718 312326 169954
rect 312562 169718 312646 169954
rect 312882 169718 312914 169954
rect 312294 169634 312914 169718
rect 312294 169398 312326 169634
rect 312562 169398 312646 169634
rect 312882 169398 312914 169634
rect 312294 133954 312914 169398
rect 312294 133718 312326 133954
rect 312562 133718 312646 133954
rect 312882 133718 312914 133954
rect 312294 133634 312914 133718
rect 312294 133398 312326 133634
rect 312562 133398 312646 133634
rect 312882 133398 312914 133634
rect 312294 97954 312914 133398
rect 312294 97718 312326 97954
rect 312562 97718 312646 97954
rect 312882 97718 312914 97954
rect 312294 97634 312914 97718
rect 312294 97398 312326 97634
rect 312562 97398 312646 97634
rect 312882 97398 312914 97634
rect 312294 61954 312914 97398
rect 312294 61718 312326 61954
rect 312562 61718 312646 61954
rect 312882 61718 312914 61954
rect 312294 61634 312914 61718
rect 312294 61398 312326 61634
rect 312562 61398 312646 61634
rect 312882 61398 312914 61634
rect 312294 25954 312914 61398
rect 312294 25718 312326 25954
rect 312562 25718 312646 25954
rect 312882 25718 312914 25954
rect 312294 25634 312914 25718
rect 312294 25398 312326 25634
rect 312562 25398 312646 25634
rect 312882 25398 312914 25634
rect 312294 -5146 312914 25398
rect 312294 -5382 312326 -5146
rect 312562 -5382 312646 -5146
rect 312882 -5382 312914 -5146
rect 312294 -5466 312914 -5382
rect 312294 -5702 312326 -5466
rect 312562 -5702 312646 -5466
rect 312882 -5702 312914 -5466
rect 312294 -7654 312914 -5702
rect 316794 710598 317414 711590
rect 316794 710362 316826 710598
rect 317062 710362 317146 710598
rect 317382 710362 317414 710598
rect 316794 710278 317414 710362
rect 316794 710042 316826 710278
rect 317062 710042 317146 710278
rect 317382 710042 317414 710278
rect 316794 678454 317414 710042
rect 316794 678218 316826 678454
rect 317062 678218 317146 678454
rect 317382 678218 317414 678454
rect 316794 678134 317414 678218
rect 316794 677898 316826 678134
rect 317062 677898 317146 678134
rect 317382 677898 317414 678134
rect 316794 642454 317414 677898
rect 316794 642218 316826 642454
rect 317062 642218 317146 642454
rect 317382 642218 317414 642454
rect 316794 642134 317414 642218
rect 316794 641898 316826 642134
rect 317062 641898 317146 642134
rect 317382 641898 317414 642134
rect 316794 606454 317414 641898
rect 316794 606218 316826 606454
rect 317062 606218 317146 606454
rect 317382 606218 317414 606454
rect 316794 606134 317414 606218
rect 316794 605898 316826 606134
rect 317062 605898 317146 606134
rect 317382 605898 317414 606134
rect 316794 570454 317414 605898
rect 316794 570218 316826 570454
rect 317062 570218 317146 570454
rect 317382 570218 317414 570454
rect 316794 570134 317414 570218
rect 316794 569898 316826 570134
rect 317062 569898 317146 570134
rect 317382 569898 317414 570134
rect 316794 534454 317414 569898
rect 316794 534218 316826 534454
rect 317062 534218 317146 534454
rect 317382 534218 317414 534454
rect 316794 534134 317414 534218
rect 316794 533898 316826 534134
rect 317062 533898 317146 534134
rect 317382 533898 317414 534134
rect 316794 498454 317414 533898
rect 316794 498218 316826 498454
rect 317062 498218 317146 498454
rect 317382 498218 317414 498454
rect 316794 498134 317414 498218
rect 316794 497898 316826 498134
rect 317062 497898 317146 498134
rect 317382 497898 317414 498134
rect 316794 462454 317414 497898
rect 316794 462218 316826 462454
rect 317062 462218 317146 462454
rect 317382 462218 317414 462454
rect 316794 462134 317414 462218
rect 316794 461898 316826 462134
rect 317062 461898 317146 462134
rect 317382 461898 317414 462134
rect 316794 426454 317414 461898
rect 316794 426218 316826 426454
rect 317062 426218 317146 426454
rect 317382 426218 317414 426454
rect 316794 426134 317414 426218
rect 316794 425898 316826 426134
rect 317062 425898 317146 426134
rect 317382 425898 317414 426134
rect 316794 390454 317414 425898
rect 316794 390218 316826 390454
rect 317062 390218 317146 390454
rect 317382 390218 317414 390454
rect 316794 390134 317414 390218
rect 316794 389898 316826 390134
rect 317062 389898 317146 390134
rect 317382 389898 317414 390134
rect 316794 354454 317414 389898
rect 316794 354218 316826 354454
rect 317062 354218 317146 354454
rect 317382 354218 317414 354454
rect 316794 354134 317414 354218
rect 316794 353898 316826 354134
rect 317062 353898 317146 354134
rect 317382 353898 317414 354134
rect 316794 318454 317414 353898
rect 316794 318218 316826 318454
rect 317062 318218 317146 318454
rect 317382 318218 317414 318454
rect 316794 318134 317414 318218
rect 316794 317898 316826 318134
rect 317062 317898 317146 318134
rect 317382 317898 317414 318134
rect 316794 282454 317414 317898
rect 316794 282218 316826 282454
rect 317062 282218 317146 282454
rect 317382 282218 317414 282454
rect 316794 282134 317414 282218
rect 316794 281898 316826 282134
rect 317062 281898 317146 282134
rect 317382 281898 317414 282134
rect 316794 246454 317414 281898
rect 316794 246218 316826 246454
rect 317062 246218 317146 246454
rect 317382 246218 317414 246454
rect 316794 246134 317414 246218
rect 316794 245898 316826 246134
rect 317062 245898 317146 246134
rect 317382 245898 317414 246134
rect 316794 210454 317414 245898
rect 316794 210218 316826 210454
rect 317062 210218 317146 210454
rect 317382 210218 317414 210454
rect 316794 210134 317414 210218
rect 316794 209898 316826 210134
rect 317062 209898 317146 210134
rect 317382 209898 317414 210134
rect 316794 174454 317414 209898
rect 316794 174218 316826 174454
rect 317062 174218 317146 174454
rect 317382 174218 317414 174454
rect 316794 174134 317414 174218
rect 316794 173898 316826 174134
rect 317062 173898 317146 174134
rect 317382 173898 317414 174134
rect 316794 138454 317414 173898
rect 316794 138218 316826 138454
rect 317062 138218 317146 138454
rect 317382 138218 317414 138454
rect 316794 138134 317414 138218
rect 316794 137898 316826 138134
rect 317062 137898 317146 138134
rect 317382 137898 317414 138134
rect 316794 102454 317414 137898
rect 316794 102218 316826 102454
rect 317062 102218 317146 102454
rect 317382 102218 317414 102454
rect 316794 102134 317414 102218
rect 316794 101898 316826 102134
rect 317062 101898 317146 102134
rect 317382 101898 317414 102134
rect 316794 66454 317414 101898
rect 316794 66218 316826 66454
rect 317062 66218 317146 66454
rect 317382 66218 317414 66454
rect 316794 66134 317414 66218
rect 316794 65898 316826 66134
rect 317062 65898 317146 66134
rect 317382 65898 317414 66134
rect 316794 30454 317414 65898
rect 316794 30218 316826 30454
rect 317062 30218 317146 30454
rect 317382 30218 317414 30454
rect 316794 30134 317414 30218
rect 316794 29898 316826 30134
rect 317062 29898 317146 30134
rect 317382 29898 317414 30134
rect 316794 -6106 317414 29898
rect 316794 -6342 316826 -6106
rect 317062 -6342 317146 -6106
rect 317382 -6342 317414 -6106
rect 316794 -6426 317414 -6342
rect 316794 -6662 316826 -6426
rect 317062 -6662 317146 -6426
rect 317382 -6662 317414 -6426
rect 316794 -7654 317414 -6662
rect 321294 711558 321914 711590
rect 321294 711322 321326 711558
rect 321562 711322 321646 711558
rect 321882 711322 321914 711558
rect 321294 711238 321914 711322
rect 321294 711002 321326 711238
rect 321562 711002 321646 711238
rect 321882 711002 321914 711238
rect 321294 682954 321914 711002
rect 321294 682718 321326 682954
rect 321562 682718 321646 682954
rect 321882 682718 321914 682954
rect 321294 682634 321914 682718
rect 321294 682398 321326 682634
rect 321562 682398 321646 682634
rect 321882 682398 321914 682634
rect 321294 646954 321914 682398
rect 321294 646718 321326 646954
rect 321562 646718 321646 646954
rect 321882 646718 321914 646954
rect 321294 646634 321914 646718
rect 321294 646398 321326 646634
rect 321562 646398 321646 646634
rect 321882 646398 321914 646634
rect 321294 610954 321914 646398
rect 321294 610718 321326 610954
rect 321562 610718 321646 610954
rect 321882 610718 321914 610954
rect 321294 610634 321914 610718
rect 321294 610398 321326 610634
rect 321562 610398 321646 610634
rect 321882 610398 321914 610634
rect 321294 574954 321914 610398
rect 321294 574718 321326 574954
rect 321562 574718 321646 574954
rect 321882 574718 321914 574954
rect 321294 574634 321914 574718
rect 321294 574398 321326 574634
rect 321562 574398 321646 574634
rect 321882 574398 321914 574634
rect 321294 538954 321914 574398
rect 321294 538718 321326 538954
rect 321562 538718 321646 538954
rect 321882 538718 321914 538954
rect 321294 538634 321914 538718
rect 321294 538398 321326 538634
rect 321562 538398 321646 538634
rect 321882 538398 321914 538634
rect 321294 502954 321914 538398
rect 321294 502718 321326 502954
rect 321562 502718 321646 502954
rect 321882 502718 321914 502954
rect 321294 502634 321914 502718
rect 321294 502398 321326 502634
rect 321562 502398 321646 502634
rect 321882 502398 321914 502634
rect 321294 466954 321914 502398
rect 321294 466718 321326 466954
rect 321562 466718 321646 466954
rect 321882 466718 321914 466954
rect 321294 466634 321914 466718
rect 321294 466398 321326 466634
rect 321562 466398 321646 466634
rect 321882 466398 321914 466634
rect 321294 430954 321914 466398
rect 321294 430718 321326 430954
rect 321562 430718 321646 430954
rect 321882 430718 321914 430954
rect 321294 430634 321914 430718
rect 321294 430398 321326 430634
rect 321562 430398 321646 430634
rect 321882 430398 321914 430634
rect 321294 394954 321914 430398
rect 321294 394718 321326 394954
rect 321562 394718 321646 394954
rect 321882 394718 321914 394954
rect 321294 394634 321914 394718
rect 321294 394398 321326 394634
rect 321562 394398 321646 394634
rect 321882 394398 321914 394634
rect 321294 358954 321914 394398
rect 321294 358718 321326 358954
rect 321562 358718 321646 358954
rect 321882 358718 321914 358954
rect 321294 358634 321914 358718
rect 321294 358398 321326 358634
rect 321562 358398 321646 358634
rect 321882 358398 321914 358634
rect 321294 322954 321914 358398
rect 321294 322718 321326 322954
rect 321562 322718 321646 322954
rect 321882 322718 321914 322954
rect 321294 322634 321914 322718
rect 321294 322398 321326 322634
rect 321562 322398 321646 322634
rect 321882 322398 321914 322634
rect 321294 286954 321914 322398
rect 321294 286718 321326 286954
rect 321562 286718 321646 286954
rect 321882 286718 321914 286954
rect 321294 286634 321914 286718
rect 321294 286398 321326 286634
rect 321562 286398 321646 286634
rect 321882 286398 321914 286634
rect 321294 250954 321914 286398
rect 321294 250718 321326 250954
rect 321562 250718 321646 250954
rect 321882 250718 321914 250954
rect 321294 250634 321914 250718
rect 321294 250398 321326 250634
rect 321562 250398 321646 250634
rect 321882 250398 321914 250634
rect 321294 214954 321914 250398
rect 321294 214718 321326 214954
rect 321562 214718 321646 214954
rect 321882 214718 321914 214954
rect 321294 214634 321914 214718
rect 321294 214398 321326 214634
rect 321562 214398 321646 214634
rect 321882 214398 321914 214634
rect 321294 178954 321914 214398
rect 321294 178718 321326 178954
rect 321562 178718 321646 178954
rect 321882 178718 321914 178954
rect 321294 178634 321914 178718
rect 321294 178398 321326 178634
rect 321562 178398 321646 178634
rect 321882 178398 321914 178634
rect 321294 142954 321914 178398
rect 321294 142718 321326 142954
rect 321562 142718 321646 142954
rect 321882 142718 321914 142954
rect 321294 142634 321914 142718
rect 321294 142398 321326 142634
rect 321562 142398 321646 142634
rect 321882 142398 321914 142634
rect 321294 106954 321914 142398
rect 321294 106718 321326 106954
rect 321562 106718 321646 106954
rect 321882 106718 321914 106954
rect 321294 106634 321914 106718
rect 321294 106398 321326 106634
rect 321562 106398 321646 106634
rect 321882 106398 321914 106634
rect 321294 70954 321914 106398
rect 321294 70718 321326 70954
rect 321562 70718 321646 70954
rect 321882 70718 321914 70954
rect 321294 70634 321914 70718
rect 321294 70398 321326 70634
rect 321562 70398 321646 70634
rect 321882 70398 321914 70634
rect 321294 34954 321914 70398
rect 321294 34718 321326 34954
rect 321562 34718 321646 34954
rect 321882 34718 321914 34954
rect 321294 34634 321914 34718
rect 321294 34398 321326 34634
rect 321562 34398 321646 34634
rect 321882 34398 321914 34634
rect 321294 -7066 321914 34398
rect 321294 -7302 321326 -7066
rect 321562 -7302 321646 -7066
rect 321882 -7302 321914 -7066
rect 321294 -7386 321914 -7302
rect 321294 -7622 321326 -7386
rect 321562 -7622 321646 -7386
rect 321882 -7622 321914 -7386
rect 321294 -7654 321914 -7622
rect 325794 704838 326414 711590
rect 325794 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 326414 704838
rect 325794 704518 326414 704602
rect 325794 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 326414 704518
rect 325794 687454 326414 704282
rect 325794 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 326414 687454
rect 325794 687134 326414 687218
rect 325794 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 326414 687134
rect 325794 651454 326414 686898
rect 325794 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 326414 651454
rect 325794 651134 326414 651218
rect 325794 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 326414 651134
rect 325794 615454 326414 650898
rect 325794 615218 325826 615454
rect 326062 615218 326146 615454
rect 326382 615218 326414 615454
rect 325794 615134 326414 615218
rect 325794 614898 325826 615134
rect 326062 614898 326146 615134
rect 326382 614898 326414 615134
rect 325794 579454 326414 614898
rect 325794 579218 325826 579454
rect 326062 579218 326146 579454
rect 326382 579218 326414 579454
rect 325794 579134 326414 579218
rect 325794 578898 325826 579134
rect 326062 578898 326146 579134
rect 326382 578898 326414 579134
rect 325794 543454 326414 578898
rect 325794 543218 325826 543454
rect 326062 543218 326146 543454
rect 326382 543218 326414 543454
rect 325794 543134 326414 543218
rect 325794 542898 325826 543134
rect 326062 542898 326146 543134
rect 326382 542898 326414 543134
rect 325794 507454 326414 542898
rect 325794 507218 325826 507454
rect 326062 507218 326146 507454
rect 326382 507218 326414 507454
rect 325794 507134 326414 507218
rect 325794 506898 325826 507134
rect 326062 506898 326146 507134
rect 326382 506898 326414 507134
rect 325794 471454 326414 506898
rect 325794 471218 325826 471454
rect 326062 471218 326146 471454
rect 326382 471218 326414 471454
rect 325794 471134 326414 471218
rect 325794 470898 325826 471134
rect 326062 470898 326146 471134
rect 326382 470898 326414 471134
rect 325794 435454 326414 470898
rect 325794 435218 325826 435454
rect 326062 435218 326146 435454
rect 326382 435218 326414 435454
rect 325794 435134 326414 435218
rect 325794 434898 325826 435134
rect 326062 434898 326146 435134
rect 326382 434898 326414 435134
rect 325794 399454 326414 434898
rect 325794 399218 325826 399454
rect 326062 399218 326146 399454
rect 326382 399218 326414 399454
rect 325794 399134 326414 399218
rect 325794 398898 325826 399134
rect 326062 398898 326146 399134
rect 326382 398898 326414 399134
rect 325794 363454 326414 398898
rect 325794 363218 325826 363454
rect 326062 363218 326146 363454
rect 326382 363218 326414 363454
rect 325794 363134 326414 363218
rect 325794 362898 325826 363134
rect 326062 362898 326146 363134
rect 326382 362898 326414 363134
rect 325794 327454 326414 362898
rect 325794 327218 325826 327454
rect 326062 327218 326146 327454
rect 326382 327218 326414 327454
rect 325794 327134 326414 327218
rect 325794 326898 325826 327134
rect 326062 326898 326146 327134
rect 326382 326898 326414 327134
rect 325794 291454 326414 326898
rect 325794 291218 325826 291454
rect 326062 291218 326146 291454
rect 326382 291218 326414 291454
rect 325794 291134 326414 291218
rect 325794 290898 325826 291134
rect 326062 290898 326146 291134
rect 326382 290898 326414 291134
rect 325794 255454 326414 290898
rect 325794 255218 325826 255454
rect 326062 255218 326146 255454
rect 326382 255218 326414 255454
rect 325794 255134 326414 255218
rect 325794 254898 325826 255134
rect 326062 254898 326146 255134
rect 326382 254898 326414 255134
rect 325794 219454 326414 254898
rect 325794 219218 325826 219454
rect 326062 219218 326146 219454
rect 326382 219218 326414 219454
rect 325794 219134 326414 219218
rect 325794 218898 325826 219134
rect 326062 218898 326146 219134
rect 326382 218898 326414 219134
rect 325794 183454 326414 218898
rect 325794 183218 325826 183454
rect 326062 183218 326146 183454
rect 326382 183218 326414 183454
rect 325794 183134 326414 183218
rect 325794 182898 325826 183134
rect 326062 182898 326146 183134
rect 326382 182898 326414 183134
rect 325794 147454 326414 182898
rect 325794 147218 325826 147454
rect 326062 147218 326146 147454
rect 326382 147218 326414 147454
rect 325794 147134 326414 147218
rect 325794 146898 325826 147134
rect 326062 146898 326146 147134
rect 326382 146898 326414 147134
rect 325794 111454 326414 146898
rect 325794 111218 325826 111454
rect 326062 111218 326146 111454
rect 326382 111218 326414 111454
rect 325794 111134 326414 111218
rect 325794 110898 325826 111134
rect 326062 110898 326146 111134
rect 326382 110898 326414 111134
rect 325794 75454 326414 110898
rect 325794 75218 325826 75454
rect 326062 75218 326146 75454
rect 326382 75218 326414 75454
rect 325794 75134 326414 75218
rect 325794 74898 325826 75134
rect 326062 74898 326146 75134
rect 326382 74898 326414 75134
rect 325794 39454 326414 74898
rect 325794 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 326414 39454
rect 325794 39134 326414 39218
rect 325794 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 326414 39134
rect 325794 3454 326414 38898
rect 325794 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 326414 3454
rect 325794 3134 326414 3218
rect 325794 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 326414 3134
rect 325794 -346 326414 2898
rect 325794 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 326414 -346
rect 325794 -666 326414 -582
rect 325794 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 326414 -666
rect 325794 -7654 326414 -902
rect 330294 705798 330914 711590
rect 330294 705562 330326 705798
rect 330562 705562 330646 705798
rect 330882 705562 330914 705798
rect 330294 705478 330914 705562
rect 330294 705242 330326 705478
rect 330562 705242 330646 705478
rect 330882 705242 330914 705478
rect 330294 691954 330914 705242
rect 330294 691718 330326 691954
rect 330562 691718 330646 691954
rect 330882 691718 330914 691954
rect 330294 691634 330914 691718
rect 330294 691398 330326 691634
rect 330562 691398 330646 691634
rect 330882 691398 330914 691634
rect 330294 655954 330914 691398
rect 330294 655718 330326 655954
rect 330562 655718 330646 655954
rect 330882 655718 330914 655954
rect 330294 655634 330914 655718
rect 330294 655398 330326 655634
rect 330562 655398 330646 655634
rect 330882 655398 330914 655634
rect 330294 619954 330914 655398
rect 330294 619718 330326 619954
rect 330562 619718 330646 619954
rect 330882 619718 330914 619954
rect 330294 619634 330914 619718
rect 330294 619398 330326 619634
rect 330562 619398 330646 619634
rect 330882 619398 330914 619634
rect 330294 583954 330914 619398
rect 330294 583718 330326 583954
rect 330562 583718 330646 583954
rect 330882 583718 330914 583954
rect 330294 583634 330914 583718
rect 330294 583398 330326 583634
rect 330562 583398 330646 583634
rect 330882 583398 330914 583634
rect 330294 547954 330914 583398
rect 330294 547718 330326 547954
rect 330562 547718 330646 547954
rect 330882 547718 330914 547954
rect 330294 547634 330914 547718
rect 330294 547398 330326 547634
rect 330562 547398 330646 547634
rect 330882 547398 330914 547634
rect 330294 511954 330914 547398
rect 330294 511718 330326 511954
rect 330562 511718 330646 511954
rect 330882 511718 330914 511954
rect 330294 511634 330914 511718
rect 330294 511398 330326 511634
rect 330562 511398 330646 511634
rect 330882 511398 330914 511634
rect 330294 475954 330914 511398
rect 330294 475718 330326 475954
rect 330562 475718 330646 475954
rect 330882 475718 330914 475954
rect 330294 475634 330914 475718
rect 330294 475398 330326 475634
rect 330562 475398 330646 475634
rect 330882 475398 330914 475634
rect 330294 439954 330914 475398
rect 330294 439718 330326 439954
rect 330562 439718 330646 439954
rect 330882 439718 330914 439954
rect 330294 439634 330914 439718
rect 330294 439398 330326 439634
rect 330562 439398 330646 439634
rect 330882 439398 330914 439634
rect 330294 403954 330914 439398
rect 330294 403718 330326 403954
rect 330562 403718 330646 403954
rect 330882 403718 330914 403954
rect 330294 403634 330914 403718
rect 330294 403398 330326 403634
rect 330562 403398 330646 403634
rect 330882 403398 330914 403634
rect 330294 367954 330914 403398
rect 330294 367718 330326 367954
rect 330562 367718 330646 367954
rect 330882 367718 330914 367954
rect 330294 367634 330914 367718
rect 330294 367398 330326 367634
rect 330562 367398 330646 367634
rect 330882 367398 330914 367634
rect 330294 331954 330914 367398
rect 330294 331718 330326 331954
rect 330562 331718 330646 331954
rect 330882 331718 330914 331954
rect 330294 331634 330914 331718
rect 330294 331398 330326 331634
rect 330562 331398 330646 331634
rect 330882 331398 330914 331634
rect 330294 295954 330914 331398
rect 330294 295718 330326 295954
rect 330562 295718 330646 295954
rect 330882 295718 330914 295954
rect 330294 295634 330914 295718
rect 330294 295398 330326 295634
rect 330562 295398 330646 295634
rect 330882 295398 330914 295634
rect 330294 259954 330914 295398
rect 330294 259718 330326 259954
rect 330562 259718 330646 259954
rect 330882 259718 330914 259954
rect 330294 259634 330914 259718
rect 330294 259398 330326 259634
rect 330562 259398 330646 259634
rect 330882 259398 330914 259634
rect 330294 223954 330914 259398
rect 330294 223718 330326 223954
rect 330562 223718 330646 223954
rect 330882 223718 330914 223954
rect 330294 223634 330914 223718
rect 330294 223398 330326 223634
rect 330562 223398 330646 223634
rect 330882 223398 330914 223634
rect 330294 187954 330914 223398
rect 330294 187718 330326 187954
rect 330562 187718 330646 187954
rect 330882 187718 330914 187954
rect 330294 187634 330914 187718
rect 330294 187398 330326 187634
rect 330562 187398 330646 187634
rect 330882 187398 330914 187634
rect 330294 151954 330914 187398
rect 330294 151718 330326 151954
rect 330562 151718 330646 151954
rect 330882 151718 330914 151954
rect 330294 151634 330914 151718
rect 330294 151398 330326 151634
rect 330562 151398 330646 151634
rect 330882 151398 330914 151634
rect 330294 115954 330914 151398
rect 330294 115718 330326 115954
rect 330562 115718 330646 115954
rect 330882 115718 330914 115954
rect 330294 115634 330914 115718
rect 330294 115398 330326 115634
rect 330562 115398 330646 115634
rect 330882 115398 330914 115634
rect 330294 79954 330914 115398
rect 330294 79718 330326 79954
rect 330562 79718 330646 79954
rect 330882 79718 330914 79954
rect 330294 79634 330914 79718
rect 330294 79398 330326 79634
rect 330562 79398 330646 79634
rect 330882 79398 330914 79634
rect 330294 43954 330914 79398
rect 330294 43718 330326 43954
rect 330562 43718 330646 43954
rect 330882 43718 330914 43954
rect 330294 43634 330914 43718
rect 330294 43398 330326 43634
rect 330562 43398 330646 43634
rect 330882 43398 330914 43634
rect 330294 7954 330914 43398
rect 330294 7718 330326 7954
rect 330562 7718 330646 7954
rect 330882 7718 330914 7954
rect 330294 7634 330914 7718
rect 330294 7398 330326 7634
rect 330562 7398 330646 7634
rect 330882 7398 330914 7634
rect 330294 -1306 330914 7398
rect 330294 -1542 330326 -1306
rect 330562 -1542 330646 -1306
rect 330882 -1542 330914 -1306
rect 330294 -1626 330914 -1542
rect 330294 -1862 330326 -1626
rect 330562 -1862 330646 -1626
rect 330882 -1862 330914 -1626
rect 330294 -7654 330914 -1862
rect 334794 706758 335414 711590
rect 334794 706522 334826 706758
rect 335062 706522 335146 706758
rect 335382 706522 335414 706758
rect 334794 706438 335414 706522
rect 334794 706202 334826 706438
rect 335062 706202 335146 706438
rect 335382 706202 335414 706438
rect 334794 696454 335414 706202
rect 334794 696218 334826 696454
rect 335062 696218 335146 696454
rect 335382 696218 335414 696454
rect 334794 696134 335414 696218
rect 334794 695898 334826 696134
rect 335062 695898 335146 696134
rect 335382 695898 335414 696134
rect 334794 660454 335414 695898
rect 334794 660218 334826 660454
rect 335062 660218 335146 660454
rect 335382 660218 335414 660454
rect 334794 660134 335414 660218
rect 334794 659898 334826 660134
rect 335062 659898 335146 660134
rect 335382 659898 335414 660134
rect 334794 624454 335414 659898
rect 334794 624218 334826 624454
rect 335062 624218 335146 624454
rect 335382 624218 335414 624454
rect 334794 624134 335414 624218
rect 334794 623898 334826 624134
rect 335062 623898 335146 624134
rect 335382 623898 335414 624134
rect 334794 588454 335414 623898
rect 334794 588218 334826 588454
rect 335062 588218 335146 588454
rect 335382 588218 335414 588454
rect 334794 588134 335414 588218
rect 334794 587898 334826 588134
rect 335062 587898 335146 588134
rect 335382 587898 335414 588134
rect 334794 552454 335414 587898
rect 334794 552218 334826 552454
rect 335062 552218 335146 552454
rect 335382 552218 335414 552454
rect 334794 552134 335414 552218
rect 334794 551898 334826 552134
rect 335062 551898 335146 552134
rect 335382 551898 335414 552134
rect 334794 516454 335414 551898
rect 334794 516218 334826 516454
rect 335062 516218 335146 516454
rect 335382 516218 335414 516454
rect 334794 516134 335414 516218
rect 334794 515898 334826 516134
rect 335062 515898 335146 516134
rect 335382 515898 335414 516134
rect 334794 480454 335414 515898
rect 334794 480218 334826 480454
rect 335062 480218 335146 480454
rect 335382 480218 335414 480454
rect 334794 480134 335414 480218
rect 334794 479898 334826 480134
rect 335062 479898 335146 480134
rect 335382 479898 335414 480134
rect 334794 444454 335414 479898
rect 334794 444218 334826 444454
rect 335062 444218 335146 444454
rect 335382 444218 335414 444454
rect 334794 444134 335414 444218
rect 334794 443898 334826 444134
rect 335062 443898 335146 444134
rect 335382 443898 335414 444134
rect 334794 408454 335414 443898
rect 334794 408218 334826 408454
rect 335062 408218 335146 408454
rect 335382 408218 335414 408454
rect 334794 408134 335414 408218
rect 334794 407898 334826 408134
rect 335062 407898 335146 408134
rect 335382 407898 335414 408134
rect 334794 372454 335414 407898
rect 334794 372218 334826 372454
rect 335062 372218 335146 372454
rect 335382 372218 335414 372454
rect 334794 372134 335414 372218
rect 334794 371898 334826 372134
rect 335062 371898 335146 372134
rect 335382 371898 335414 372134
rect 334794 336454 335414 371898
rect 334794 336218 334826 336454
rect 335062 336218 335146 336454
rect 335382 336218 335414 336454
rect 334794 336134 335414 336218
rect 334794 335898 334826 336134
rect 335062 335898 335146 336134
rect 335382 335898 335414 336134
rect 334794 300454 335414 335898
rect 334794 300218 334826 300454
rect 335062 300218 335146 300454
rect 335382 300218 335414 300454
rect 334794 300134 335414 300218
rect 334794 299898 334826 300134
rect 335062 299898 335146 300134
rect 335382 299898 335414 300134
rect 334794 264454 335414 299898
rect 334794 264218 334826 264454
rect 335062 264218 335146 264454
rect 335382 264218 335414 264454
rect 334794 264134 335414 264218
rect 334794 263898 334826 264134
rect 335062 263898 335146 264134
rect 335382 263898 335414 264134
rect 334794 228454 335414 263898
rect 334794 228218 334826 228454
rect 335062 228218 335146 228454
rect 335382 228218 335414 228454
rect 334794 228134 335414 228218
rect 334794 227898 334826 228134
rect 335062 227898 335146 228134
rect 335382 227898 335414 228134
rect 334794 192454 335414 227898
rect 334794 192218 334826 192454
rect 335062 192218 335146 192454
rect 335382 192218 335414 192454
rect 334794 192134 335414 192218
rect 334794 191898 334826 192134
rect 335062 191898 335146 192134
rect 335382 191898 335414 192134
rect 334794 156454 335414 191898
rect 334794 156218 334826 156454
rect 335062 156218 335146 156454
rect 335382 156218 335414 156454
rect 334794 156134 335414 156218
rect 334794 155898 334826 156134
rect 335062 155898 335146 156134
rect 335382 155898 335414 156134
rect 334794 120454 335414 155898
rect 334794 120218 334826 120454
rect 335062 120218 335146 120454
rect 335382 120218 335414 120454
rect 334794 120134 335414 120218
rect 334794 119898 334826 120134
rect 335062 119898 335146 120134
rect 335382 119898 335414 120134
rect 334794 84454 335414 119898
rect 334794 84218 334826 84454
rect 335062 84218 335146 84454
rect 335382 84218 335414 84454
rect 334794 84134 335414 84218
rect 334794 83898 334826 84134
rect 335062 83898 335146 84134
rect 335382 83898 335414 84134
rect 334794 48454 335414 83898
rect 334794 48218 334826 48454
rect 335062 48218 335146 48454
rect 335382 48218 335414 48454
rect 334794 48134 335414 48218
rect 334794 47898 334826 48134
rect 335062 47898 335146 48134
rect 335382 47898 335414 48134
rect 334794 12454 335414 47898
rect 334794 12218 334826 12454
rect 335062 12218 335146 12454
rect 335382 12218 335414 12454
rect 334794 12134 335414 12218
rect 334794 11898 334826 12134
rect 335062 11898 335146 12134
rect 335382 11898 335414 12134
rect 334794 -2266 335414 11898
rect 334794 -2502 334826 -2266
rect 335062 -2502 335146 -2266
rect 335382 -2502 335414 -2266
rect 334794 -2586 335414 -2502
rect 334794 -2822 334826 -2586
rect 335062 -2822 335146 -2586
rect 335382 -2822 335414 -2586
rect 334794 -7654 335414 -2822
rect 339294 707718 339914 711590
rect 339294 707482 339326 707718
rect 339562 707482 339646 707718
rect 339882 707482 339914 707718
rect 339294 707398 339914 707482
rect 339294 707162 339326 707398
rect 339562 707162 339646 707398
rect 339882 707162 339914 707398
rect 339294 700954 339914 707162
rect 339294 700718 339326 700954
rect 339562 700718 339646 700954
rect 339882 700718 339914 700954
rect 339294 700634 339914 700718
rect 339294 700398 339326 700634
rect 339562 700398 339646 700634
rect 339882 700398 339914 700634
rect 339294 664954 339914 700398
rect 339294 664718 339326 664954
rect 339562 664718 339646 664954
rect 339882 664718 339914 664954
rect 339294 664634 339914 664718
rect 339294 664398 339326 664634
rect 339562 664398 339646 664634
rect 339882 664398 339914 664634
rect 339294 628954 339914 664398
rect 339294 628718 339326 628954
rect 339562 628718 339646 628954
rect 339882 628718 339914 628954
rect 339294 628634 339914 628718
rect 339294 628398 339326 628634
rect 339562 628398 339646 628634
rect 339882 628398 339914 628634
rect 339294 592954 339914 628398
rect 339294 592718 339326 592954
rect 339562 592718 339646 592954
rect 339882 592718 339914 592954
rect 339294 592634 339914 592718
rect 339294 592398 339326 592634
rect 339562 592398 339646 592634
rect 339882 592398 339914 592634
rect 339294 556954 339914 592398
rect 339294 556718 339326 556954
rect 339562 556718 339646 556954
rect 339882 556718 339914 556954
rect 339294 556634 339914 556718
rect 339294 556398 339326 556634
rect 339562 556398 339646 556634
rect 339882 556398 339914 556634
rect 339294 520954 339914 556398
rect 339294 520718 339326 520954
rect 339562 520718 339646 520954
rect 339882 520718 339914 520954
rect 339294 520634 339914 520718
rect 339294 520398 339326 520634
rect 339562 520398 339646 520634
rect 339882 520398 339914 520634
rect 339294 484954 339914 520398
rect 339294 484718 339326 484954
rect 339562 484718 339646 484954
rect 339882 484718 339914 484954
rect 339294 484634 339914 484718
rect 339294 484398 339326 484634
rect 339562 484398 339646 484634
rect 339882 484398 339914 484634
rect 339294 448954 339914 484398
rect 339294 448718 339326 448954
rect 339562 448718 339646 448954
rect 339882 448718 339914 448954
rect 339294 448634 339914 448718
rect 339294 448398 339326 448634
rect 339562 448398 339646 448634
rect 339882 448398 339914 448634
rect 339294 412954 339914 448398
rect 339294 412718 339326 412954
rect 339562 412718 339646 412954
rect 339882 412718 339914 412954
rect 339294 412634 339914 412718
rect 339294 412398 339326 412634
rect 339562 412398 339646 412634
rect 339882 412398 339914 412634
rect 339294 376954 339914 412398
rect 339294 376718 339326 376954
rect 339562 376718 339646 376954
rect 339882 376718 339914 376954
rect 339294 376634 339914 376718
rect 339294 376398 339326 376634
rect 339562 376398 339646 376634
rect 339882 376398 339914 376634
rect 339294 340954 339914 376398
rect 339294 340718 339326 340954
rect 339562 340718 339646 340954
rect 339882 340718 339914 340954
rect 339294 340634 339914 340718
rect 339294 340398 339326 340634
rect 339562 340398 339646 340634
rect 339882 340398 339914 340634
rect 339294 304954 339914 340398
rect 339294 304718 339326 304954
rect 339562 304718 339646 304954
rect 339882 304718 339914 304954
rect 339294 304634 339914 304718
rect 339294 304398 339326 304634
rect 339562 304398 339646 304634
rect 339882 304398 339914 304634
rect 339294 268954 339914 304398
rect 339294 268718 339326 268954
rect 339562 268718 339646 268954
rect 339882 268718 339914 268954
rect 339294 268634 339914 268718
rect 339294 268398 339326 268634
rect 339562 268398 339646 268634
rect 339882 268398 339914 268634
rect 339294 232954 339914 268398
rect 339294 232718 339326 232954
rect 339562 232718 339646 232954
rect 339882 232718 339914 232954
rect 339294 232634 339914 232718
rect 339294 232398 339326 232634
rect 339562 232398 339646 232634
rect 339882 232398 339914 232634
rect 339294 196954 339914 232398
rect 339294 196718 339326 196954
rect 339562 196718 339646 196954
rect 339882 196718 339914 196954
rect 339294 196634 339914 196718
rect 339294 196398 339326 196634
rect 339562 196398 339646 196634
rect 339882 196398 339914 196634
rect 339294 160954 339914 196398
rect 339294 160718 339326 160954
rect 339562 160718 339646 160954
rect 339882 160718 339914 160954
rect 339294 160634 339914 160718
rect 339294 160398 339326 160634
rect 339562 160398 339646 160634
rect 339882 160398 339914 160634
rect 339294 124954 339914 160398
rect 339294 124718 339326 124954
rect 339562 124718 339646 124954
rect 339882 124718 339914 124954
rect 339294 124634 339914 124718
rect 339294 124398 339326 124634
rect 339562 124398 339646 124634
rect 339882 124398 339914 124634
rect 339294 88954 339914 124398
rect 339294 88718 339326 88954
rect 339562 88718 339646 88954
rect 339882 88718 339914 88954
rect 339294 88634 339914 88718
rect 339294 88398 339326 88634
rect 339562 88398 339646 88634
rect 339882 88398 339914 88634
rect 339294 52954 339914 88398
rect 339294 52718 339326 52954
rect 339562 52718 339646 52954
rect 339882 52718 339914 52954
rect 339294 52634 339914 52718
rect 339294 52398 339326 52634
rect 339562 52398 339646 52634
rect 339882 52398 339914 52634
rect 339294 16954 339914 52398
rect 339294 16718 339326 16954
rect 339562 16718 339646 16954
rect 339882 16718 339914 16954
rect 339294 16634 339914 16718
rect 339294 16398 339326 16634
rect 339562 16398 339646 16634
rect 339882 16398 339914 16634
rect 339294 -3226 339914 16398
rect 339294 -3462 339326 -3226
rect 339562 -3462 339646 -3226
rect 339882 -3462 339914 -3226
rect 339294 -3546 339914 -3462
rect 339294 -3782 339326 -3546
rect 339562 -3782 339646 -3546
rect 339882 -3782 339914 -3546
rect 339294 -7654 339914 -3782
rect 343794 708678 344414 711590
rect 343794 708442 343826 708678
rect 344062 708442 344146 708678
rect 344382 708442 344414 708678
rect 343794 708358 344414 708442
rect 343794 708122 343826 708358
rect 344062 708122 344146 708358
rect 344382 708122 344414 708358
rect 343794 669454 344414 708122
rect 343794 669218 343826 669454
rect 344062 669218 344146 669454
rect 344382 669218 344414 669454
rect 343794 669134 344414 669218
rect 343794 668898 343826 669134
rect 344062 668898 344146 669134
rect 344382 668898 344414 669134
rect 343794 633454 344414 668898
rect 343794 633218 343826 633454
rect 344062 633218 344146 633454
rect 344382 633218 344414 633454
rect 343794 633134 344414 633218
rect 343794 632898 343826 633134
rect 344062 632898 344146 633134
rect 344382 632898 344414 633134
rect 343794 597454 344414 632898
rect 343794 597218 343826 597454
rect 344062 597218 344146 597454
rect 344382 597218 344414 597454
rect 343794 597134 344414 597218
rect 343794 596898 343826 597134
rect 344062 596898 344146 597134
rect 344382 596898 344414 597134
rect 343794 561454 344414 596898
rect 343794 561218 343826 561454
rect 344062 561218 344146 561454
rect 344382 561218 344414 561454
rect 343794 561134 344414 561218
rect 343794 560898 343826 561134
rect 344062 560898 344146 561134
rect 344382 560898 344414 561134
rect 343794 525454 344414 560898
rect 343794 525218 343826 525454
rect 344062 525218 344146 525454
rect 344382 525218 344414 525454
rect 343794 525134 344414 525218
rect 343794 524898 343826 525134
rect 344062 524898 344146 525134
rect 344382 524898 344414 525134
rect 343794 489454 344414 524898
rect 343794 489218 343826 489454
rect 344062 489218 344146 489454
rect 344382 489218 344414 489454
rect 343794 489134 344414 489218
rect 343794 488898 343826 489134
rect 344062 488898 344146 489134
rect 344382 488898 344414 489134
rect 343794 453454 344414 488898
rect 343794 453218 343826 453454
rect 344062 453218 344146 453454
rect 344382 453218 344414 453454
rect 343794 453134 344414 453218
rect 343794 452898 343826 453134
rect 344062 452898 344146 453134
rect 344382 452898 344414 453134
rect 343794 417454 344414 452898
rect 343794 417218 343826 417454
rect 344062 417218 344146 417454
rect 344382 417218 344414 417454
rect 343794 417134 344414 417218
rect 343794 416898 343826 417134
rect 344062 416898 344146 417134
rect 344382 416898 344414 417134
rect 343794 381454 344414 416898
rect 343794 381218 343826 381454
rect 344062 381218 344146 381454
rect 344382 381218 344414 381454
rect 343794 381134 344414 381218
rect 343794 380898 343826 381134
rect 344062 380898 344146 381134
rect 344382 380898 344414 381134
rect 343794 345454 344414 380898
rect 343794 345218 343826 345454
rect 344062 345218 344146 345454
rect 344382 345218 344414 345454
rect 343794 345134 344414 345218
rect 343794 344898 343826 345134
rect 344062 344898 344146 345134
rect 344382 344898 344414 345134
rect 343794 309454 344414 344898
rect 343794 309218 343826 309454
rect 344062 309218 344146 309454
rect 344382 309218 344414 309454
rect 343794 309134 344414 309218
rect 343794 308898 343826 309134
rect 344062 308898 344146 309134
rect 344382 308898 344414 309134
rect 343794 273454 344414 308898
rect 343794 273218 343826 273454
rect 344062 273218 344146 273454
rect 344382 273218 344414 273454
rect 343794 273134 344414 273218
rect 343794 272898 343826 273134
rect 344062 272898 344146 273134
rect 344382 272898 344414 273134
rect 343794 237454 344414 272898
rect 343794 237218 343826 237454
rect 344062 237218 344146 237454
rect 344382 237218 344414 237454
rect 343794 237134 344414 237218
rect 343794 236898 343826 237134
rect 344062 236898 344146 237134
rect 344382 236898 344414 237134
rect 343794 201454 344414 236898
rect 343794 201218 343826 201454
rect 344062 201218 344146 201454
rect 344382 201218 344414 201454
rect 343794 201134 344414 201218
rect 343794 200898 343826 201134
rect 344062 200898 344146 201134
rect 344382 200898 344414 201134
rect 343794 165454 344414 200898
rect 343794 165218 343826 165454
rect 344062 165218 344146 165454
rect 344382 165218 344414 165454
rect 343794 165134 344414 165218
rect 343794 164898 343826 165134
rect 344062 164898 344146 165134
rect 344382 164898 344414 165134
rect 343794 129454 344414 164898
rect 343794 129218 343826 129454
rect 344062 129218 344146 129454
rect 344382 129218 344414 129454
rect 343794 129134 344414 129218
rect 343794 128898 343826 129134
rect 344062 128898 344146 129134
rect 344382 128898 344414 129134
rect 343794 93454 344414 128898
rect 343794 93218 343826 93454
rect 344062 93218 344146 93454
rect 344382 93218 344414 93454
rect 343794 93134 344414 93218
rect 343794 92898 343826 93134
rect 344062 92898 344146 93134
rect 344382 92898 344414 93134
rect 343794 57454 344414 92898
rect 343794 57218 343826 57454
rect 344062 57218 344146 57454
rect 344382 57218 344414 57454
rect 343794 57134 344414 57218
rect 343794 56898 343826 57134
rect 344062 56898 344146 57134
rect 344382 56898 344414 57134
rect 343794 21454 344414 56898
rect 343794 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 344414 21454
rect 343794 21134 344414 21218
rect 343794 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 344414 21134
rect 343794 -4186 344414 20898
rect 343794 -4422 343826 -4186
rect 344062 -4422 344146 -4186
rect 344382 -4422 344414 -4186
rect 343794 -4506 344414 -4422
rect 343794 -4742 343826 -4506
rect 344062 -4742 344146 -4506
rect 344382 -4742 344414 -4506
rect 343794 -7654 344414 -4742
rect 348294 709638 348914 711590
rect 348294 709402 348326 709638
rect 348562 709402 348646 709638
rect 348882 709402 348914 709638
rect 348294 709318 348914 709402
rect 348294 709082 348326 709318
rect 348562 709082 348646 709318
rect 348882 709082 348914 709318
rect 348294 673954 348914 709082
rect 348294 673718 348326 673954
rect 348562 673718 348646 673954
rect 348882 673718 348914 673954
rect 348294 673634 348914 673718
rect 348294 673398 348326 673634
rect 348562 673398 348646 673634
rect 348882 673398 348914 673634
rect 348294 637954 348914 673398
rect 348294 637718 348326 637954
rect 348562 637718 348646 637954
rect 348882 637718 348914 637954
rect 348294 637634 348914 637718
rect 348294 637398 348326 637634
rect 348562 637398 348646 637634
rect 348882 637398 348914 637634
rect 348294 601954 348914 637398
rect 348294 601718 348326 601954
rect 348562 601718 348646 601954
rect 348882 601718 348914 601954
rect 348294 601634 348914 601718
rect 348294 601398 348326 601634
rect 348562 601398 348646 601634
rect 348882 601398 348914 601634
rect 348294 565954 348914 601398
rect 348294 565718 348326 565954
rect 348562 565718 348646 565954
rect 348882 565718 348914 565954
rect 348294 565634 348914 565718
rect 348294 565398 348326 565634
rect 348562 565398 348646 565634
rect 348882 565398 348914 565634
rect 348294 529954 348914 565398
rect 348294 529718 348326 529954
rect 348562 529718 348646 529954
rect 348882 529718 348914 529954
rect 348294 529634 348914 529718
rect 348294 529398 348326 529634
rect 348562 529398 348646 529634
rect 348882 529398 348914 529634
rect 348294 493954 348914 529398
rect 348294 493718 348326 493954
rect 348562 493718 348646 493954
rect 348882 493718 348914 493954
rect 348294 493634 348914 493718
rect 348294 493398 348326 493634
rect 348562 493398 348646 493634
rect 348882 493398 348914 493634
rect 348294 457954 348914 493398
rect 348294 457718 348326 457954
rect 348562 457718 348646 457954
rect 348882 457718 348914 457954
rect 348294 457634 348914 457718
rect 348294 457398 348326 457634
rect 348562 457398 348646 457634
rect 348882 457398 348914 457634
rect 348294 421954 348914 457398
rect 348294 421718 348326 421954
rect 348562 421718 348646 421954
rect 348882 421718 348914 421954
rect 348294 421634 348914 421718
rect 348294 421398 348326 421634
rect 348562 421398 348646 421634
rect 348882 421398 348914 421634
rect 348294 385954 348914 421398
rect 348294 385718 348326 385954
rect 348562 385718 348646 385954
rect 348882 385718 348914 385954
rect 348294 385634 348914 385718
rect 348294 385398 348326 385634
rect 348562 385398 348646 385634
rect 348882 385398 348914 385634
rect 348294 349954 348914 385398
rect 348294 349718 348326 349954
rect 348562 349718 348646 349954
rect 348882 349718 348914 349954
rect 348294 349634 348914 349718
rect 348294 349398 348326 349634
rect 348562 349398 348646 349634
rect 348882 349398 348914 349634
rect 348294 313954 348914 349398
rect 348294 313718 348326 313954
rect 348562 313718 348646 313954
rect 348882 313718 348914 313954
rect 348294 313634 348914 313718
rect 348294 313398 348326 313634
rect 348562 313398 348646 313634
rect 348882 313398 348914 313634
rect 348294 277954 348914 313398
rect 348294 277718 348326 277954
rect 348562 277718 348646 277954
rect 348882 277718 348914 277954
rect 348294 277634 348914 277718
rect 348294 277398 348326 277634
rect 348562 277398 348646 277634
rect 348882 277398 348914 277634
rect 348294 241954 348914 277398
rect 348294 241718 348326 241954
rect 348562 241718 348646 241954
rect 348882 241718 348914 241954
rect 348294 241634 348914 241718
rect 348294 241398 348326 241634
rect 348562 241398 348646 241634
rect 348882 241398 348914 241634
rect 348294 205954 348914 241398
rect 348294 205718 348326 205954
rect 348562 205718 348646 205954
rect 348882 205718 348914 205954
rect 348294 205634 348914 205718
rect 348294 205398 348326 205634
rect 348562 205398 348646 205634
rect 348882 205398 348914 205634
rect 348294 169954 348914 205398
rect 348294 169718 348326 169954
rect 348562 169718 348646 169954
rect 348882 169718 348914 169954
rect 348294 169634 348914 169718
rect 348294 169398 348326 169634
rect 348562 169398 348646 169634
rect 348882 169398 348914 169634
rect 348294 133954 348914 169398
rect 348294 133718 348326 133954
rect 348562 133718 348646 133954
rect 348882 133718 348914 133954
rect 348294 133634 348914 133718
rect 348294 133398 348326 133634
rect 348562 133398 348646 133634
rect 348882 133398 348914 133634
rect 348294 97954 348914 133398
rect 348294 97718 348326 97954
rect 348562 97718 348646 97954
rect 348882 97718 348914 97954
rect 348294 97634 348914 97718
rect 348294 97398 348326 97634
rect 348562 97398 348646 97634
rect 348882 97398 348914 97634
rect 348294 61954 348914 97398
rect 348294 61718 348326 61954
rect 348562 61718 348646 61954
rect 348882 61718 348914 61954
rect 348294 61634 348914 61718
rect 348294 61398 348326 61634
rect 348562 61398 348646 61634
rect 348882 61398 348914 61634
rect 348294 25954 348914 61398
rect 348294 25718 348326 25954
rect 348562 25718 348646 25954
rect 348882 25718 348914 25954
rect 348294 25634 348914 25718
rect 348294 25398 348326 25634
rect 348562 25398 348646 25634
rect 348882 25398 348914 25634
rect 348294 -5146 348914 25398
rect 348294 -5382 348326 -5146
rect 348562 -5382 348646 -5146
rect 348882 -5382 348914 -5146
rect 348294 -5466 348914 -5382
rect 348294 -5702 348326 -5466
rect 348562 -5702 348646 -5466
rect 348882 -5702 348914 -5466
rect 348294 -7654 348914 -5702
rect 352794 710598 353414 711590
rect 352794 710362 352826 710598
rect 353062 710362 353146 710598
rect 353382 710362 353414 710598
rect 352794 710278 353414 710362
rect 352794 710042 352826 710278
rect 353062 710042 353146 710278
rect 353382 710042 353414 710278
rect 352794 678454 353414 710042
rect 352794 678218 352826 678454
rect 353062 678218 353146 678454
rect 353382 678218 353414 678454
rect 352794 678134 353414 678218
rect 352794 677898 352826 678134
rect 353062 677898 353146 678134
rect 353382 677898 353414 678134
rect 352794 642454 353414 677898
rect 352794 642218 352826 642454
rect 353062 642218 353146 642454
rect 353382 642218 353414 642454
rect 352794 642134 353414 642218
rect 352794 641898 352826 642134
rect 353062 641898 353146 642134
rect 353382 641898 353414 642134
rect 352794 606454 353414 641898
rect 352794 606218 352826 606454
rect 353062 606218 353146 606454
rect 353382 606218 353414 606454
rect 352794 606134 353414 606218
rect 352794 605898 352826 606134
rect 353062 605898 353146 606134
rect 353382 605898 353414 606134
rect 352794 570454 353414 605898
rect 352794 570218 352826 570454
rect 353062 570218 353146 570454
rect 353382 570218 353414 570454
rect 352794 570134 353414 570218
rect 352794 569898 352826 570134
rect 353062 569898 353146 570134
rect 353382 569898 353414 570134
rect 352794 534454 353414 569898
rect 352794 534218 352826 534454
rect 353062 534218 353146 534454
rect 353382 534218 353414 534454
rect 352794 534134 353414 534218
rect 352794 533898 352826 534134
rect 353062 533898 353146 534134
rect 353382 533898 353414 534134
rect 352794 498454 353414 533898
rect 352794 498218 352826 498454
rect 353062 498218 353146 498454
rect 353382 498218 353414 498454
rect 352794 498134 353414 498218
rect 352794 497898 352826 498134
rect 353062 497898 353146 498134
rect 353382 497898 353414 498134
rect 352794 462454 353414 497898
rect 352794 462218 352826 462454
rect 353062 462218 353146 462454
rect 353382 462218 353414 462454
rect 352794 462134 353414 462218
rect 352794 461898 352826 462134
rect 353062 461898 353146 462134
rect 353382 461898 353414 462134
rect 352794 426454 353414 461898
rect 352794 426218 352826 426454
rect 353062 426218 353146 426454
rect 353382 426218 353414 426454
rect 352794 426134 353414 426218
rect 352794 425898 352826 426134
rect 353062 425898 353146 426134
rect 353382 425898 353414 426134
rect 352794 390454 353414 425898
rect 352794 390218 352826 390454
rect 353062 390218 353146 390454
rect 353382 390218 353414 390454
rect 352794 390134 353414 390218
rect 352794 389898 352826 390134
rect 353062 389898 353146 390134
rect 353382 389898 353414 390134
rect 352794 354454 353414 389898
rect 352794 354218 352826 354454
rect 353062 354218 353146 354454
rect 353382 354218 353414 354454
rect 352794 354134 353414 354218
rect 352794 353898 352826 354134
rect 353062 353898 353146 354134
rect 353382 353898 353414 354134
rect 352794 318454 353414 353898
rect 352794 318218 352826 318454
rect 353062 318218 353146 318454
rect 353382 318218 353414 318454
rect 352794 318134 353414 318218
rect 352794 317898 352826 318134
rect 353062 317898 353146 318134
rect 353382 317898 353414 318134
rect 352794 282454 353414 317898
rect 352794 282218 352826 282454
rect 353062 282218 353146 282454
rect 353382 282218 353414 282454
rect 352794 282134 353414 282218
rect 352794 281898 352826 282134
rect 353062 281898 353146 282134
rect 353382 281898 353414 282134
rect 352794 246454 353414 281898
rect 352794 246218 352826 246454
rect 353062 246218 353146 246454
rect 353382 246218 353414 246454
rect 352794 246134 353414 246218
rect 352794 245898 352826 246134
rect 353062 245898 353146 246134
rect 353382 245898 353414 246134
rect 352794 210454 353414 245898
rect 352794 210218 352826 210454
rect 353062 210218 353146 210454
rect 353382 210218 353414 210454
rect 352794 210134 353414 210218
rect 352794 209898 352826 210134
rect 353062 209898 353146 210134
rect 353382 209898 353414 210134
rect 352794 174454 353414 209898
rect 352794 174218 352826 174454
rect 353062 174218 353146 174454
rect 353382 174218 353414 174454
rect 352794 174134 353414 174218
rect 352794 173898 352826 174134
rect 353062 173898 353146 174134
rect 353382 173898 353414 174134
rect 352794 138454 353414 173898
rect 352794 138218 352826 138454
rect 353062 138218 353146 138454
rect 353382 138218 353414 138454
rect 352794 138134 353414 138218
rect 352794 137898 352826 138134
rect 353062 137898 353146 138134
rect 353382 137898 353414 138134
rect 352794 102454 353414 137898
rect 352794 102218 352826 102454
rect 353062 102218 353146 102454
rect 353382 102218 353414 102454
rect 352794 102134 353414 102218
rect 352794 101898 352826 102134
rect 353062 101898 353146 102134
rect 353382 101898 353414 102134
rect 352794 66454 353414 101898
rect 352794 66218 352826 66454
rect 353062 66218 353146 66454
rect 353382 66218 353414 66454
rect 352794 66134 353414 66218
rect 352794 65898 352826 66134
rect 353062 65898 353146 66134
rect 353382 65898 353414 66134
rect 352794 30454 353414 65898
rect 352794 30218 352826 30454
rect 353062 30218 353146 30454
rect 353382 30218 353414 30454
rect 352794 30134 353414 30218
rect 352794 29898 352826 30134
rect 353062 29898 353146 30134
rect 353382 29898 353414 30134
rect 352794 -6106 353414 29898
rect 352794 -6342 352826 -6106
rect 353062 -6342 353146 -6106
rect 353382 -6342 353414 -6106
rect 352794 -6426 353414 -6342
rect 352794 -6662 352826 -6426
rect 353062 -6662 353146 -6426
rect 353382 -6662 353414 -6426
rect 352794 -7654 353414 -6662
rect 357294 711558 357914 711590
rect 357294 711322 357326 711558
rect 357562 711322 357646 711558
rect 357882 711322 357914 711558
rect 357294 711238 357914 711322
rect 357294 711002 357326 711238
rect 357562 711002 357646 711238
rect 357882 711002 357914 711238
rect 357294 682954 357914 711002
rect 357294 682718 357326 682954
rect 357562 682718 357646 682954
rect 357882 682718 357914 682954
rect 357294 682634 357914 682718
rect 357294 682398 357326 682634
rect 357562 682398 357646 682634
rect 357882 682398 357914 682634
rect 357294 646954 357914 682398
rect 357294 646718 357326 646954
rect 357562 646718 357646 646954
rect 357882 646718 357914 646954
rect 357294 646634 357914 646718
rect 357294 646398 357326 646634
rect 357562 646398 357646 646634
rect 357882 646398 357914 646634
rect 357294 610954 357914 646398
rect 357294 610718 357326 610954
rect 357562 610718 357646 610954
rect 357882 610718 357914 610954
rect 357294 610634 357914 610718
rect 357294 610398 357326 610634
rect 357562 610398 357646 610634
rect 357882 610398 357914 610634
rect 357294 574954 357914 610398
rect 357294 574718 357326 574954
rect 357562 574718 357646 574954
rect 357882 574718 357914 574954
rect 357294 574634 357914 574718
rect 357294 574398 357326 574634
rect 357562 574398 357646 574634
rect 357882 574398 357914 574634
rect 357294 538954 357914 574398
rect 357294 538718 357326 538954
rect 357562 538718 357646 538954
rect 357882 538718 357914 538954
rect 357294 538634 357914 538718
rect 357294 538398 357326 538634
rect 357562 538398 357646 538634
rect 357882 538398 357914 538634
rect 357294 502954 357914 538398
rect 357294 502718 357326 502954
rect 357562 502718 357646 502954
rect 357882 502718 357914 502954
rect 357294 502634 357914 502718
rect 357294 502398 357326 502634
rect 357562 502398 357646 502634
rect 357882 502398 357914 502634
rect 357294 466954 357914 502398
rect 357294 466718 357326 466954
rect 357562 466718 357646 466954
rect 357882 466718 357914 466954
rect 357294 466634 357914 466718
rect 357294 466398 357326 466634
rect 357562 466398 357646 466634
rect 357882 466398 357914 466634
rect 357294 430954 357914 466398
rect 357294 430718 357326 430954
rect 357562 430718 357646 430954
rect 357882 430718 357914 430954
rect 357294 430634 357914 430718
rect 357294 430398 357326 430634
rect 357562 430398 357646 430634
rect 357882 430398 357914 430634
rect 357294 394954 357914 430398
rect 357294 394718 357326 394954
rect 357562 394718 357646 394954
rect 357882 394718 357914 394954
rect 357294 394634 357914 394718
rect 357294 394398 357326 394634
rect 357562 394398 357646 394634
rect 357882 394398 357914 394634
rect 357294 358954 357914 394398
rect 357294 358718 357326 358954
rect 357562 358718 357646 358954
rect 357882 358718 357914 358954
rect 357294 358634 357914 358718
rect 357294 358398 357326 358634
rect 357562 358398 357646 358634
rect 357882 358398 357914 358634
rect 357294 322954 357914 358398
rect 357294 322718 357326 322954
rect 357562 322718 357646 322954
rect 357882 322718 357914 322954
rect 357294 322634 357914 322718
rect 357294 322398 357326 322634
rect 357562 322398 357646 322634
rect 357882 322398 357914 322634
rect 357294 286954 357914 322398
rect 357294 286718 357326 286954
rect 357562 286718 357646 286954
rect 357882 286718 357914 286954
rect 357294 286634 357914 286718
rect 357294 286398 357326 286634
rect 357562 286398 357646 286634
rect 357882 286398 357914 286634
rect 357294 250954 357914 286398
rect 357294 250718 357326 250954
rect 357562 250718 357646 250954
rect 357882 250718 357914 250954
rect 357294 250634 357914 250718
rect 357294 250398 357326 250634
rect 357562 250398 357646 250634
rect 357882 250398 357914 250634
rect 357294 214954 357914 250398
rect 357294 214718 357326 214954
rect 357562 214718 357646 214954
rect 357882 214718 357914 214954
rect 357294 214634 357914 214718
rect 357294 214398 357326 214634
rect 357562 214398 357646 214634
rect 357882 214398 357914 214634
rect 357294 178954 357914 214398
rect 357294 178718 357326 178954
rect 357562 178718 357646 178954
rect 357882 178718 357914 178954
rect 357294 178634 357914 178718
rect 357294 178398 357326 178634
rect 357562 178398 357646 178634
rect 357882 178398 357914 178634
rect 357294 142954 357914 178398
rect 357294 142718 357326 142954
rect 357562 142718 357646 142954
rect 357882 142718 357914 142954
rect 357294 142634 357914 142718
rect 357294 142398 357326 142634
rect 357562 142398 357646 142634
rect 357882 142398 357914 142634
rect 357294 106954 357914 142398
rect 357294 106718 357326 106954
rect 357562 106718 357646 106954
rect 357882 106718 357914 106954
rect 357294 106634 357914 106718
rect 357294 106398 357326 106634
rect 357562 106398 357646 106634
rect 357882 106398 357914 106634
rect 357294 70954 357914 106398
rect 357294 70718 357326 70954
rect 357562 70718 357646 70954
rect 357882 70718 357914 70954
rect 357294 70634 357914 70718
rect 357294 70398 357326 70634
rect 357562 70398 357646 70634
rect 357882 70398 357914 70634
rect 357294 34954 357914 70398
rect 357294 34718 357326 34954
rect 357562 34718 357646 34954
rect 357882 34718 357914 34954
rect 357294 34634 357914 34718
rect 357294 34398 357326 34634
rect 357562 34398 357646 34634
rect 357882 34398 357914 34634
rect 357294 -7066 357914 34398
rect 357294 -7302 357326 -7066
rect 357562 -7302 357646 -7066
rect 357882 -7302 357914 -7066
rect 357294 -7386 357914 -7302
rect 357294 -7622 357326 -7386
rect 357562 -7622 357646 -7386
rect 357882 -7622 357914 -7386
rect 357294 -7654 357914 -7622
rect 361794 704838 362414 711590
rect 361794 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 362414 704838
rect 361794 704518 362414 704602
rect 361794 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 362414 704518
rect 361794 687454 362414 704282
rect 361794 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 362414 687454
rect 361794 687134 362414 687218
rect 361794 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 362414 687134
rect 361794 651454 362414 686898
rect 361794 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 362414 651454
rect 361794 651134 362414 651218
rect 361794 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 362414 651134
rect 361794 615454 362414 650898
rect 361794 615218 361826 615454
rect 362062 615218 362146 615454
rect 362382 615218 362414 615454
rect 361794 615134 362414 615218
rect 361794 614898 361826 615134
rect 362062 614898 362146 615134
rect 362382 614898 362414 615134
rect 361794 579454 362414 614898
rect 361794 579218 361826 579454
rect 362062 579218 362146 579454
rect 362382 579218 362414 579454
rect 361794 579134 362414 579218
rect 361794 578898 361826 579134
rect 362062 578898 362146 579134
rect 362382 578898 362414 579134
rect 361794 543454 362414 578898
rect 361794 543218 361826 543454
rect 362062 543218 362146 543454
rect 362382 543218 362414 543454
rect 361794 543134 362414 543218
rect 361794 542898 361826 543134
rect 362062 542898 362146 543134
rect 362382 542898 362414 543134
rect 361794 507454 362414 542898
rect 361794 507218 361826 507454
rect 362062 507218 362146 507454
rect 362382 507218 362414 507454
rect 361794 507134 362414 507218
rect 361794 506898 361826 507134
rect 362062 506898 362146 507134
rect 362382 506898 362414 507134
rect 361794 471454 362414 506898
rect 361794 471218 361826 471454
rect 362062 471218 362146 471454
rect 362382 471218 362414 471454
rect 361794 471134 362414 471218
rect 361794 470898 361826 471134
rect 362062 470898 362146 471134
rect 362382 470898 362414 471134
rect 361794 435454 362414 470898
rect 361794 435218 361826 435454
rect 362062 435218 362146 435454
rect 362382 435218 362414 435454
rect 361794 435134 362414 435218
rect 361794 434898 361826 435134
rect 362062 434898 362146 435134
rect 362382 434898 362414 435134
rect 361794 399454 362414 434898
rect 361794 399218 361826 399454
rect 362062 399218 362146 399454
rect 362382 399218 362414 399454
rect 361794 399134 362414 399218
rect 361794 398898 361826 399134
rect 362062 398898 362146 399134
rect 362382 398898 362414 399134
rect 361794 363454 362414 398898
rect 361794 363218 361826 363454
rect 362062 363218 362146 363454
rect 362382 363218 362414 363454
rect 361794 363134 362414 363218
rect 361794 362898 361826 363134
rect 362062 362898 362146 363134
rect 362382 362898 362414 363134
rect 361794 327454 362414 362898
rect 361794 327218 361826 327454
rect 362062 327218 362146 327454
rect 362382 327218 362414 327454
rect 361794 327134 362414 327218
rect 361794 326898 361826 327134
rect 362062 326898 362146 327134
rect 362382 326898 362414 327134
rect 361794 291454 362414 326898
rect 361794 291218 361826 291454
rect 362062 291218 362146 291454
rect 362382 291218 362414 291454
rect 361794 291134 362414 291218
rect 361794 290898 361826 291134
rect 362062 290898 362146 291134
rect 362382 290898 362414 291134
rect 361794 255454 362414 290898
rect 361794 255218 361826 255454
rect 362062 255218 362146 255454
rect 362382 255218 362414 255454
rect 361794 255134 362414 255218
rect 361794 254898 361826 255134
rect 362062 254898 362146 255134
rect 362382 254898 362414 255134
rect 361794 219454 362414 254898
rect 361794 219218 361826 219454
rect 362062 219218 362146 219454
rect 362382 219218 362414 219454
rect 361794 219134 362414 219218
rect 361794 218898 361826 219134
rect 362062 218898 362146 219134
rect 362382 218898 362414 219134
rect 361794 183454 362414 218898
rect 361794 183218 361826 183454
rect 362062 183218 362146 183454
rect 362382 183218 362414 183454
rect 361794 183134 362414 183218
rect 361794 182898 361826 183134
rect 362062 182898 362146 183134
rect 362382 182898 362414 183134
rect 361794 147454 362414 182898
rect 361794 147218 361826 147454
rect 362062 147218 362146 147454
rect 362382 147218 362414 147454
rect 361794 147134 362414 147218
rect 361794 146898 361826 147134
rect 362062 146898 362146 147134
rect 362382 146898 362414 147134
rect 361794 111454 362414 146898
rect 361794 111218 361826 111454
rect 362062 111218 362146 111454
rect 362382 111218 362414 111454
rect 361794 111134 362414 111218
rect 361794 110898 361826 111134
rect 362062 110898 362146 111134
rect 362382 110898 362414 111134
rect 361794 75454 362414 110898
rect 361794 75218 361826 75454
rect 362062 75218 362146 75454
rect 362382 75218 362414 75454
rect 361794 75134 362414 75218
rect 361794 74898 361826 75134
rect 362062 74898 362146 75134
rect 362382 74898 362414 75134
rect 361794 39454 362414 74898
rect 361794 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 362414 39454
rect 361794 39134 362414 39218
rect 361794 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 362414 39134
rect 361794 3454 362414 38898
rect 361794 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 362414 3454
rect 361794 3134 362414 3218
rect 361794 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 362414 3134
rect 361794 -346 362414 2898
rect 361794 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 362414 -346
rect 361794 -666 362414 -582
rect 361794 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 362414 -666
rect 361794 -7654 362414 -902
rect 366294 705798 366914 711590
rect 366294 705562 366326 705798
rect 366562 705562 366646 705798
rect 366882 705562 366914 705798
rect 366294 705478 366914 705562
rect 366294 705242 366326 705478
rect 366562 705242 366646 705478
rect 366882 705242 366914 705478
rect 366294 691954 366914 705242
rect 366294 691718 366326 691954
rect 366562 691718 366646 691954
rect 366882 691718 366914 691954
rect 366294 691634 366914 691718
rect 366294 691398 366326 691634
rect 366562 691398 366646 691634
rect 366882 691398 366914 691634
rect 366294 655954 366914 691398
rect 366294 655718 366326 655954
rect 366562 655718 366646 655954
rect 366882 655718 366914 655954
rect 366294 655634 366914 655718
rect 366294 655398 366326 655634
rect 366562 655398 366646 655634
rect 366882 655398 366914 655634
rect 366294 619954 366914 655398
rect 366294 619718 366326 619954
rect 366562 619718 366646 619954
rect 366882 619718 366914 619954
rect 366294 619634 366914 619718
rect 366294 619398 366326 619634
rect 366562 619398 366646 619634
rect 366882 619398 366914 619634
rect 366294 583954 366914 619398
rect 366294 583718 366326 583954
rect 366562 583718 366646 583954
rect 366882 583718 366914 583954
rect 366294 583634 366914 583718
rect 366294 583398 366326 583634
rect 366562 583398 366646 583634
rect 366882 583398 366914 583634
rect 366294 547954 366914 583398
rect 366294 547718 366326 547954
rect 366562 547718 366646 547954
rect 366882 547718 366914 547954
rect 366294 547634 366914 547718
rect 366294 547398 366326 547634
rect 366562 547398 366646 547634
rect 366882 547398 366914 547634
rect 366294 511954 366914 547398
rect 366294 511718 366326 511954
rect 366562 511718 366646 511954
rect 366882 511718 366914 511954
rect 366294 511634 366914 511718
rect 366294 511398 366326 511634
rect 366562 511398 366646 511634
rect 366882 511398 366914 511634
rect 366294 475954 366914 511398
rect 366294 475718 366326 475954
rect 366562 475718 366646 475954
rect 366882 475718 366914 475954
rect 366294 475634 366914 475718
rect 366294 475398 366326 475634
rect 366562 475398 366646 475634
rect 366882 475398 366914 475634
rect 366294 439954 366914 475398
rect 366294 439718 366326 439954
rect 366562 439718 366646 439954
rect 366882 439718 366914 439954
rect 366294 439634 366914 439718
rect 366294 439398 366326 439634
rect 366562 439398 366646 439634
rect 366882 439398 366914 439634
rect 366294 403954 366914 439398
rect 366294 403718 366326 403954
rect 366562 403718 366646 403954
rect 366882 403718 366914 403954
rect 366294 403634 366914 403718
rect 366294 403398 366326 403634
rect 366562 403398 366646 403634
rect 366882 403398 366914 403634
rect 366294 367954 366914 403398
rect 366294 367718 366326 367954
rect 366562 367718 366646 367954
rect 366882 367718 366914 367954
rect 366294 367634 366914 367718
rect 366294 367398 366326 367634
rect 366562 367398 366646 367634
rect 366882 367398 366914 367634
rect 366294 331954 366914 367398
rect 366294 331718 366326 331954
rect 366562 331718 366646 331954
rect 366882 331718 366914 331954
rect 366294 331634 366914 331718
rect 366294 331398 366326 331634
rect 366562 331398 366646 331634
rect 366882 331398 366914 331634
rect 366294 295954 366914 331398
rect 366294 295718 366326 295954
rect 366562 295718 366646 295954
rect 366882 295718 366914 295954
rect 366294 295634 366914 295718
rect 366294 295398 366326 295634
rect 366562 295398 366646 295634
rect 366882 295398 366914 295634
rect 366294 259954 366914 295398
rect 366294 259718 366326 259954
rect 366562 259718 366646 259954
rect 366882 259718 366914 259954
rect 366294 259634 366914 259718
rect 366294 259398 366326 259634
rect 366562 259398 366646 259634
rect 366882 259398 366914 259634
rect 366294 223954 366914 259398
rect 366294 223718 366326 223954
rect 366562 223718 366646 223954
rect 366882 223718 366914 223954
rect 366294 223634 366914 223718
rect 366294 223398 366326 223634
rect 366562 223398 366646 223634
rect 366882 223398 366914 223634
rect 366294 187954 366914 223398
rect 366294 187718 366326 187954
rect 366562 187718 366646 187954
rect 366882 187718 366914 187954
rect 366294 187634 366914 187718
rect 366294 187398 366326 187634
rect 366562 187398 366646 187634
rect 366882 187398 366914 187634
rect 366294 151954 366914 187398
rect 366294 151718 366326 151954
rect 366562 151718 366646 151954
rect 366882 151718 366914 151954
rect 366294 151634 366914 151718
rect 366294 151398 366326 151634
rect 366562 151398 366646 151634
rect 366882 151398 366914 151634
rect 366294 115954 366914 151398
rect 366294 115718 366326 115954
rect 366562 115718 366646 115954
rect 366882 115718 366914 115954
rect 366294 115634 366914 115718
rect 366294 115398 366326 115634
rect 366562 115398 366646 115634
rect 366882 115398 366914 115634
rect 366294 79954 366914 115398
rect 366294 79718 366326 79954
rect 366562 79718 366646 79954
rect 366882 79718 366914 79954
rect 366294 79634 366914 79718
rect 366294 79398 366326 79634
rect 366562 79398 366646 79634
rect 366882 79398 366914 79634
rect 366294 43954 366914 79398
rect 366294 43718 366326 43954
rect 366562 43718 366646 43954
rect 366882 43718 366914 43954
rect 366294 43634 366914 43718
rect 366294 43398 366326 43634
rect 366562 43398 366646 43634
rect 366882 43398 366914 43634
rect 366294 7954 366914 43398
rect 366294 7718 366326 7954
rect 366562 7718 366646 7954
rect 366882 7718 366914 7954
rect 366294 7634 366914 7718
rect 366294 7398 366326 7634
rect 366562 7398 366646 7634
rect 366882 7398 366914 7634
rect 366294 -1306 366914 7398
rect 366294 -1542 366326 -1306
rect 366562 -1542 366646 -1306
rect 366882 -1542 366914 -1306
rect 366294 -1626 366914 -1542
rect 366294 -1862 366326 -1626
rect 366562 -1862 366646 -1626
rect 366882 -1862 366914 -1626
rect 366294 -7654 366914 -1862
rect 370794 706758 371414 711590
rect 370794 706522 370826 706758
rect 371062 706522 371146 706758
rect 371382 706522 371414 706758
rect 370794 706438 371414 706522
rect 370794 706202 370826 706438
rect 371062 706202 371146 706438
rect 371382 706202 371414 706438
rect 370794 696454 371414 706202
rect 370794 696218 370826 696454
rect 371062 696218 371146 696454
rect 371382 696218 371414 696454
rect 370794 696134 371414 696218
rect 370794 695898 370826 696134
rect 371062 695898 371146 696134
rect 371382 695898 371414 696134
rect 370794 660454 371414 695898
rect 370794 660218 370826 660454
rect 371062 660218 371146 660454
rect 371382 660218 371414 660454
rect 370794 660134 371414 660218
rect 370794 659898 370826 660134
rect 371062 659898 371146 660134
rect 371382 659898 371414 660134
rect 370794 624454 371414 659898
rect 370794 624218 370826 624454
rect 371062 624218 371146 624454
rect 371382 624218 371414 624454
rect 370794 624134 371414 624218
rect 370794 623898 370826 624134
rect 371062 623898 371146 624134
rect 371382 623898 371414 624134
rect 370794 588454 371414 623898
rect 370794 588218 370826 588454
rect 371062 588218 371146 588454
rect 371382 588218 371414 588454
rect 370794 588134 371414 588218
rect 370794 587898 370826 588134
rect 371062 587898 371146 588134
rect 371382 587898 371414 588134
rect 370794 552454 371414 587898
rect 370794 552218 370826 552454
rect 371062 552218 371146 552454
rect 371382 552218 371414 552454
rect 370794 552134 371414 552218
rect 370794 551898 370826 552134
rect 371062 551898 371146 552134
rect 371382 551898 371414 552134
rect 370794 516454 371414 551898
rect 370794 516218 370826 516454
rect 371062 516218 371146 516454
rect 371382 516218 371414 516454
rect 370794 516134 371414 516218
rect 370794 515898 370826 516134
rect 371062 515898 371146 516134
rect 371382 515898 371414 516134
rect 370794 480454 371414 515898
rect 370794 480218 370826 480454
rect 371062 480218 371146 480454
rect 371382 480218 371414 480454
rect 370794 480134 371414 480218
rect 370794 479898 370826 480134
rect 371062 479898 371146 480134
rect 371382 479898 371414 480134
rect 370794 444454 371414 479898
rect 370794 444218 370826 444454
rect 371062 444218 371146 444454
rect 371382 444218 371414 444454
rect 370794 444134 371414 444218
rect 370794 443898 370826 444134
rect 371062 443898 371146 444134
rect 371382 443898 371414 444134
rect 370794 408454 371414 443898
rect 370794 408218 370826 408454
rect 371062 408218 371146 408454
rect 371382 408218 371414 408454
rect 370794 408134 371414 408218
rect 370794 407898 370826 408134
rect 371062 407898 371146 408134
rect 371382 407898 371414 408134
rect 370794 372454 371414 407898
rect 370794 372218 370826 372454
rect 371062 372218 371146 372454
rect 371382 372218 371414 372454
rect 370794 372134 371414 372218
rect 370794 371898 370826 372134
rect 371062 371898 371146 372134
rect 371382 371898 371414 372134
rect 370794 336454 371414 371898
rect 370794 336218 370826 336454
rect 371062 336218 371146 336454
rect 371382 336218 371414 336454
rect 370794 336134 371414 336218
rect 370794 335898 370826 336134
rect 371062 335898 371146 336134
rect 371382 335898 371414 336134
rect 370794 300454 371414 335898
rect 370794 300218 370826 300454
rect 371062 300218 371146 300454
rect 371382 300218 371414 300454
rect 370794 300134 371414 300218
rect 370794 299898 370826 300134
rect 371062 299898 371146 300134
rect 371382 299898 371414 300134
rect 370794 264454 371414 299898
rect 370794 264218 370826 264454
rect 371062 264218 371146 264454
rect 371382 264218 371414 264454
rect 370794 264134 371414 264218
rect 370794 263898 370826 264134
rect 371062 263898 371146 264134
rect 371382 263898 371414 264134
rect 370794 228454 371414 263898
rect 370794 228218 370826 228454
rect 371062 228218 371146 228454
rect 371382 228218 371414 228454
rect 370794 228134 371414 228218
rect 370794 227898 370826 228134
rect 371062 227898 371146 228134
rect 371382 227898 371414 228134
rect 370794 192454 371414 227898
rect 370794 192218 370826 192454
rect 371062 192218 371146 192454
rect 371382 192218 371414 192454
rect 370794 192134 371414 192218
rect 370794 191898 370826 192134
rect 371062 191898 371146 192134
rect 371382 191898 371414 192134
rect 370794 156454 371414 191898
rect 370794 156218 370826 156454
rect 371062 156218 371146 156454
rect 371382 156218 371414 156454
rect 370794 156134 371414 156218
rect 370794 155898 370826 156134
rect 371062 155898 371146 156134
rect 371382 155898 371414 156134
rect 370794 120454 371414 155898
rect 370794 120218 370826 120454
rect 371062 120218 371146 120454
rect 371382 120218 371414 120454
rect 370794 120134 371414 120218
rect 370794 119898 370826 120134
rect 371062 119898 371146 120134
rect 371382 119898 371414 120134
rect 370794 84454 371414 119898
rect 370794 84218 370826 84454
rect 371062 84218 371146 84454
rect 371382 84218 371414 84454
rect 370794 84134 371414 84218
rect 370794 83898 370826 84134
rect 371062 83898 371146 84134
rect 371382 83898 371414 84134
rect 370794 48454 371414 83898
rect 370794 48218 370826 48454
rect 371062 48218 371146 48454
rect 371382 48218 371414 48454
rect 370794 48134 371414 48218
rect 370794 47898 370826 48134
rect 371062 47898 371146 48134
rect 371382 47898 371414 48134
rect 370794 12454 371414 47898
rect 370794 12218 370826 12454
rect 371062 12218 371146 12454
rect 371382 12218 371414 12454
rect 370794 12134 371414 12218
rect 370794 11898 370826 12134
rect 371062 11898 371146 12134
rect 371382 11898 371414 12134
rect 370794 -2266 371414 11898
rect 370794 -2502 370826 -2266
rect 371062 -2502 371146 -2266
rect 371382 -2502 371414 -2266
rect 370794 -2586 371414 -2502
rect 370794 -2822 370826 -2586
rect 371062 -2822 371146 -2586
rect 371382 -2822 371414 -2586
rect 370794 -7654 371414 -2822
rect 375294 707718 375914 711590
rect 375294 707482 375326 707718
rect 375562 707482 375646 707718
rect 375882 707482 375914 707718
rect 375294 707398 375914 707482
rect 375294 707162 375326 707398
rect 375562 707162 375646 707398
rect 375882 707162 375914 707398
rect 375294 700954 375914 707162
rect 375294 700718 375326 700954
rect 375562 700718 375646 700954
rect 375882 700718 375914 700954
rect 375294 700634 375914 700718
rect 375294 700398 375326 700634
rect 375562 700398 375646 700634
rect 375882 700398 375914 700634
rect 375294 664954 375914 700398
rect 375294 664718 375326 664954
rect 375562 664718 375646 664954
rect 375882 664718 375914 664954
rect 375294 664634 375914 664718
rect 375294 664398 375326 664634
rect 375562 664398 375646 664634
rect 375882 664398 375914 664634
rect 375294 628954 375914 664398
rect 375294 628718 375326 628954
rect 375562 628718 375646 628954
rect 375882 628718 375914 628954
rect 375294 628634 375914 628718
rect 375294 628398 375326 628634
rect 375562 628398 375646 628634
rect 375882 628398 375914 628634
rect 375294 592954 375914 628398
rect 375294 592718 375326 592954
rect 375562 592718 375646 592954
rect 375882 592718 375914 592954
rect 375294 592634 375914 592718
rect 375294 592398 375326 592634
rect 375562 592398 375646 592634
rect 375882 592398 375914 592634
rect 375294 556954 375914 592398
rect 375294 556718 375326 556954
rect 375562 556718 375646 556954
rect 375882 556718 375914 556954
rect 375294 556634 375914 556718
rect 375294 556398 375326 556634
rect 375562 556398 375646 556634
rect 375882 556398 375914 556634
rect 375294 520954 375914 556398
rect 375294 520718 375326 520954
rect 375562 520718 375646 520954
rect 375882 520718 375914 520954
rect 375294 520634 375914 520718
rect 375294 520398 375326 520634
rect 375562 520398 375646 520634
rect 375882 520398 375914 520634
rect 375294 484954 375914 520398
rect 375294 484718 375326 484954
rect 375562 484718 375646 484954
rect 375882 484718 375914 484954
rect 375294 484634 375914 484718
rect 375294 484398 375326 484634
rect 375562 484398 375646 484634
rect 375882 484398 375914 484634
rect 375294 448954 375914 484398
rect 375294 448718 375326 448954
rect 375562 448718 375646 448954
rect 375882 448718 375914 448954
rect 375294 448634 375914 448718
rect 375294 448398 375326 448634
rect 375562 448398 375646 448634
rect 375882 448398 375914 448634
rect 375294 412954 375914 448398
rect 375294 412718 375326 412954
rect 375562 412718 375646 412954
rect 375882 412718 375914 412954
rect 375294 412634 375914 412718
rect 375294 412398 375326 412634
rect 375562 412398 375646 412634
rect 375882 412398 375914 412634
rect 375294 376954 375914 412398
rect 375294 376718 375326 376954
rect 375562 376718 375646 376954
rect 375882 376718 375914 376954
rect 375294 376634 375914 376718
rect 375294 376398 375326 376634
rect 375562 376398 375646 376634
rect 375882 376398 375914 376634
rect 375294 340954 375914 376398
rect 375294 340718 375326 340954
rect 375562 340718 375646 340954
rect 375882 340718 375914 340954
rect 375294 340634 375914 340718
rect 375294 340398 375326 340634
rect 375562 340398 375646 340634
rect 375882 340398 375914 340634
rect 375294 304954 375914 340398
rect 375294 304718 375326 304954
rect 375562 304718 375646 304954
rect 375882 304718 375914 304954
rect 375294 304634 375914 304718
rect 375294 304398 375326 304634
rect 375562 304398 375646 304634
rect 375882 304398 375914 304634
rect 375294 268954 375914 304398
rect 375294 268718 375326 268954
rect 375562 268718 375646 268954
rect 375882 268718 375914 268954
rect 375294 268634 375914 268718
rect 375294 268398 375326 268634
rect 375562 268398 375646 268634
rect 375882 268398 375914 268634
rect 375294 232954 375914 268398
rect 375294 232718 375326 232954
rect 375562 232718 375646 232954
rect 375882 232718 375914 232954
rect 375294 232634 375914 232718
rect 375294 232398 375326 232634
rect 375562 232398 375646 232634
rect 375882 232398 375914 232634
rect 375294 196954 375914 232398
rect 375294 196718 375326 196954
rect 375562 196718 375646 196954
rect 375882 196718 375914 196954
rect 375294 196634 375914 196718
rect 375294 196398 375326 196634
rect 375562 196398 375646 196634
rect 375882 196398 375914 196634
rect 375294 160954 375914 196398
rect 375294 160718 375326 160954
rect 375562 160718 375646 160954
rect 375882 160718 375914 160954
rect 375294 160634 375914 160718
rect 375294 160398 375326 160634
rect 375562 160398 375646 160634
rect 375882 160398 375914 160634
rect 375294 124954 375914 160398
rect 375294 124718 375326 124954
rect 375562 124718 375646 124954
rect 375882 124718 375914 124954
rect 375294 124634 375914 124718
rect 375294 124398 375326 124634
rect 375562 124398 375646 124634
rect 375882 124398 375914 124634
rect 375294 88954 375914 124398
rect 375294 88718 375326 88954
rect 375562 88718 375646 88954
rect 375882 88718 375914 88954
rect 375294 88634 375914 88718
rect 375294 88398 375326 88634
rect 375562 88398 375646 88634
rect 375882 88398 375914 88634
rect 375294 52954 375914 88398
rect 375294 52718 375326 52954
rect 375562 52718 375646 52954
rect 375882 52718 375914 52954
rect 375294 52634 375914 52718
rect 375294 52398 375326 52634
rect 375562 52398 375646 52634
rect 375882 52398 375914 52634
rect 375294 16954 375914 52398
rect 375294 16718 375326 16954
rect 375562 16718 375646 16954
rect 375882 16718 375914 16954
rect 375294 16634 375914 16718
rect 375294 16398 375326 16634
rect 375562 16398 375646 16634
rect 375882 16398 375914 16634
rect 375294 -3226 375914 16398
rect 375294 -3462 375326 -3226
rect 375562 -3462 375646 -3226
rect 375882 -3462 375914 -3226
rect 375294 -3546 375914 -3462
rect 375294 -3782 375326 -3546
rect 375562 -3782 375646 -3546
rect 375882 -3782 375914 -3546
rect 375294 -7654 375914 -3782
rect 379794 708678 380414 711590
rect 379794 708442 379826 708678
rect 380062 708442 380146 708678
rect 380382 708442 380414 708678
rect 379794 708358 380414 708442
rect 379794 708122 379826 708358
rect 380062 708122 380146 708358
rect 380382 708122 380414 708358
rect 379794 669454 380414 708122
rect 379794 669218 379826 669454
rect 380062 669218 380146 669454
rect 380382 669218 380414 669454
rect 379794 669134 380414 669218
rect 379794 668898 379826 669134
rect 380062 668898 380146 669134
rect 380382 668898 380414 669134
rect 379794 633454 380414 668898
rect 379794 633218 379826 633454
rect 380062 633218 380146 633454
rect 380382 633218 380414 633454
rect 379794 633134 380414 633218
rect 379794 632898 379826 633134
rect 380062 632898 380146 633134
rect 380382 632898 380414 633134
rect 379794 597454 380414 632898
rect 379794 597218 379826 597454
rect 380062 597218 380146 597454
rect 380382 597218 380414 597454
rect 379794 597134 380414 597218
rect 379794 596898 379826 597134
rect 380062 596898 380146 597134
rect 380382 596898 380414 597134
rect 379794 561454 380414 596898
rect 379794 561218 379826 561454
rect 380062 561218 380146 561454
rect 380382 561218 380414 561454
rect 379794 561134 380414 561218
rect 379794 560898 379826 561134
rect 380062 560898 380146 561134
rect 380382 560898 380414 561134
rect 379794 525454 380414 560898
rect 379794 525218 379826 525454
rect 380062 525218 380146 525454
rect 380382 525218 380414 525454
rect 379794 525134 380414 525218
rect 379794 524898 379826 525134
rect 380062 524898 380146 525134
rect 380382 524898 380414 525134
rect 379794 489454 380414 524898
rect 379794 489218 379826 489454
rect 380062 489218 380146 489454
rect 380382 489218 380414 489454
rect 379794 489134 380414 489218
rect 379794 488898 379826 489134
rect 380062 488898 380146 489134
rect 380382 488898 380414 489134
rect 379794 453454 380414 488898
rect 379794 453218 379826 453454
rect 380062 453218 380146 453454
rect 380382 453218 380414 453454
rect 379794 453134 380414 453218
rect 379794 452898 379826 453134
rect 380062 452898 380146 453134
rect 380382 452898 380414 453134
rect 379794 417454 380414 452898
rect 379794 417218 379826 417454
rect 380062 417218 380146 417454
rect 380382 417218 380414 417454
rect 379794 417134 380414 417218
rect 379794 416898 379826 417134
rect 380062 416898 380146 417134
rect 380382 416898 380414 417134
rect 379794 381454 380414 416898
rect 379794 381218 379826 381454
rect 380062 381218 380146 381454
rect 380382 381218 380414 381454
rect 379794 381134 380414 381218
rect 379794 380898 379826 381134
rect 380062 380898 380146 381134
rect 380382 380898 380414 381134
rect 379794 345454 380414 380898
rect 379794 345218 379826 345454
rect 380062 345218 380146 345454
rect 380382 345218 380414 345454
rect 379794 345134 380414 345218
rect 379794 344898 379826 345134
rect 380062 344898 380146 345134
rect 380382 344898 380414 345134
rect 379794 309454 380414 344898
rect 379794 309218 379826 309454
rect 380062 309218 380146 309454
rect 380382 309218 380414 309454
rect 379794 309134 380414 309218
rect 379794 308898 379826 309134
rect 380062 308898 380146 309134
rect 380382 308898 380414 309134
rect 379794 273454 380414 308898
rect 379794 273218 379826 273454
rect 380062 273218 380146 273454
rect 380382 273218 380414 273454
rect 379794 273134 380414 273218
rect 379794 272898 379826 273134
rect 380062 272898 380146 273134
rect 380382 272898 380414 273134
rect 379794 237454 380414 272898
rect 379794 237218 379826 237454
rect 380062 237218 380146 237454
rect 380382 237218 380414 237454
rect 379794 237134 380414 237218
rect 379794 236898 379826 237134
rect 380062 236898 380146 237134
rect 380382 236898 380414 237134
rect 379794 201454 380414 236898
rect 379794 201218 379826 201454
rect 380062 201218 380146 201454
rect 380382 201218 380414 201454
rect 379794 201134 380414 201218
rect 379794 200898 379826 201134
rect 380062 200898 380146 201134
rect 380382 200898 380414 201134
rect 379794 165454 380414 200898
rect 379794 165218 379826 165454
rect 380062 165218 380146 165454
rect 380382 165218 380414 165454
rect 379794 165134 380414 165218
rect 379794 164898 379826 165134
rect 380062 164898 380146 165134
rect 380382 164898 380414 165134
rect 379794 129454 380414 164898
rect 379794 129218 379826 129454
rect 380062 129218 380146 129454
rect 380382 129218 380414 129454
rect 379794 129134 380414 129218
rect 379794 128898 379826 129134
rect 380062 128898 380146 129134
rect 380382 128898 380414 129134
rect 379794 93454 380414 128898
rect 379794 93218 379826 93454
rect 380062 93218 380146 93454
rect 380382 93218 380414 93454
rect 379794 93134 380414 93218
rect 379794 92898 379826 93134
rect 380062 92898 380146 93134
rect 380382 92898 380414 93134
rect 379794 57454 380414 92898
rect 379794 57218 379826 57454
rect 380062 57218 380146 57454
rect 380382 57218 380414 57454
rect 379794 57134 380414 57218
rect 379794 56898 379826 57134
rect 380062 56898 380146 57134
rect 380382 56898 380414 57134
rect 379794 21454 380414 56898
rect 379794 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 380414 21454
rect 379794 21134 380414 21218
rect 379794 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 380414 21134
rect 379794 -4186 380414 20898
rect 379794 -4422 379826 -4186
rect 380062 -4422 380146 -4186
rect 380382 -4422 380414 -4186
rect 379794 -4506 380414 -4422
rect 379794 -4742 379826 -4506
rect 380062 -4742 380146 -4506
rect 380382 -4742 380414 -4506
rect 379794 -7654 380414 -4742
rect 384294 709638 384914 711590
rect 384294 709402 384326 709638
rect 384562 709402 384646 709638
rect 384882 709402 384914 709638
rect 384294 709318 384914 709402
rect 384294 709082 384326 709318
rect 384562 709082 384646 709318
rect 384882 709082 384914 709318
rect 384294 673954 384914 709082
rect 384294 673718 384326 673954
rect 384562 673718 384646 673954
rect 384882 673718 384914 673954
rect 384294 673634 384914 673718
rect 384294 673398 384326 673634
rect 384562 673398 384646 673634
rect 384882 673398 384914 673634
rect 384294 637954 384914 673398
rect 384294 637718 384326 637954
rect 384562 637718 384646 637954
rect 384882 637718 384914 637954
rect 384294 637634 384914 637718
rect 384294 637398 384326 637634
rect 384562 637398 384646 637634
rect 384882 637398 384914 637634
rect 384294 601954 384914 637398
rect 384294 601718 384326 601954
rect 384562 601718 384646 601954
rect 384882 601718 384914 601954
rect 384294 601634 384914 601718
rect 384294 601398 384326 601634
rect 384562 601398 384646 601634
rect 384882 601398 384914 601634
rect 384294 565954 384914 601398
rect 384294 565718 384326 565954
rect 384562 565718 384646 565954
rect 384882 565718 384914 565954
rect 384294 565634 384914 565718
rect 384294 565398 384326 565634
rect 384562 565398 384646 565634
rect 384882 565398 384914 565634
rect 384294 529954 384914 565398
rect 384294 529718 384326 529954
rect 384562 529718 384646 529954
rect 384882 529718 384914 529954
rect 384294 529634 384914 529718
rect 384294 529398 384326 529634
rect 384562 529398 384646 529634
rect 384882 529398 384914 529634
rect 384294 493954 384914 529398
rect 384294 493718 384326 493954
rect 384562 493718 384646 493954
rect 384882 493718 384914 493954
rect 384294 493634 384914 493718
rect 384294 493398 384326 493634
rect 384562 493398 384646 493634
rect 384882 493398 384914 493634
rect 384294 457954 384914 493398
rect 384294 457718 384326 457954
rect 384562 457718 384646 457954
rect 384882 457718 384914 457954
rect 384294 457634 384914 457718
rect 384294 457398 384326 457634
rect 384562 457398 384646 457634
rect 384882 457398 384914 457634
rect 384294 421954 384914 457398
rect 384294 421718 384326 421954
rect 384562 421718 384646 421954
rect 384882 421718 384914 421954
rect 384294 421634 384914 421718
rect 384294 421398 384326 421634
rect 384562 421398 384646 421634
rect 384882 421398 384914 421634
rect 384294 385954 384914 421398
rect 384294 385718 384326 385954
rect 384562 385718 384646 385954
rect 384882 385718 384914 385954
rect 384294 385634 384914 385718
rect 384294 385398 384326 385634
rect 384562 385398 384646 385634
rect 384882 385398 384914 385634
rect 384294 349954 384914 385398
rect 384294 349718 384326 349954
rect 384562 349718 384646 349954
rect 384882 349718 384914 349954
rect 384294 349634 384914 349718
rect 384294 349398 384326 349634
rect 384562 349398 384646 349634
rect 384882 349398 384914 349634
rect 384294 313954 384914 349398
rect 384294 313718 384326 313954
rect 384562 313718 384646 313954
rect 384882 313718 384914 313954
rect 384294 313634 384914 313718
rect 384294 313398 384326 313634
rect 384562 313398 384646 313634
rect 384882 313398 384914 313634
rect 384294 277954 384914 313398
rect 384294 277718 384326 277954
rect 384562 277718 384646 277954
rect 384882 277718 384914 277954
rect 384294 277634 384914 277718
rect 384294 277398 384326 277634
rect 384562 277398 384646 277634
rect 384882 277398 384914 277634
rect 384294 241954 384914 277398
rect 384294 241718 384326 241954
rect 384562 241718 384646 241954
rect 384882 241718 384914 241954
rect 384294 241634 384914 241718
rect 384294 241398 384326 241634
rect 384562 241398 384646 241634
rect 384882 241398 384914 241634
rect 384294 205954 384914 241398
rect 384294 205718 384326 205954
rect 384562 205718 384646 205954
rect 384882 205718 384914 205954
rect 384294 205634 384914 205718
rect 384294 205398 384326 205634
rect 384562 205398 384646 205634
rect 384882 205398 384914 205634
rect 384294 169954 384914 205398
rect 384294 169718 384326 169954
rect 384562 169718 384646 169954
rect 384882 169718 384914 169954
rect 384294 169634 384914 169718
rect 384294 169398 384326 169634
rect 384562 169398 384646 169634
rect 384882 169398 384914 169634
rect 384294 133954 384914 169398
rect 384294 133718 384326 133954
rect 384562 133718 384646 133954
rect 384882 133718 384914 133954
rect 384294 133634 384914 133718
rect 384294 133398 384326 133634
rect 384562 133398 384646 133634
rect 384882 133398 384914 133634
rect 384294 97954 384914 133398
rect 384294 97718 384326 97954
rect 384562 97718 384646 97954
rect 384882 97718 384914 97954
rect 384294 97634 384914 97718
rect 384294 97398 384326 97634
rect 384562 97398 384646 97634
rect 384882 97398 384914 97634
rect 384294 61954 384914 97398
rect 384294 61718 384326 61954
rect 384562 61718 384646 61954
rect 384882 61718 384914 61954
rect 384294 61634 384914 61718
rect 384294 61398 384326 61634
rect 384562 61398 384646 61634
rect 384882 61398 384914 61634
rect 384294 25954 384914 61398
rect 384294 25718 384326 25954
rect 384562 25718 384646 25954
rect 384882 25718 384914 25954
rect 384294 25634 384914 25718
rect 384294 25398 384326 25634
rect 384562 25398 384646 25634
rect 384882 25398 384914 25634
rect 384294 -5146 384914 25398
rect 384294 -5382 384326 -5146
rect 384562 -5382 384646 -5146
rect 384882 -5382 384914 -5146
rect 384294 -5466 384914 -5382
rect 384294 -5702 384326 -5466
rect 384562 -5702 384646 -5466
rect 384882 -5702 384914 -5466
rect 384294 -7654 384914 -5702
rect 388794 710598 389414 711590
rect 388794 710362 388826 710598
rect 389062 710362 389146 710598
rect 389382 710362 389414 710598
rect 388794 710278 389414 710362
rect 388794 710042 388826 710278
rect 389062 710042 389146 710278
rect 389382 710042 389414 710278
rect 388794 678454 389414 710042
rect 388794 678218 388826 678454
rect 389062 678218 389146 678454
rect 389382 678218 389414 678454
rect 388794 678134 389414 678218
rect 388794 677898 388826 678134
rect 389062 677898 389146 678134
rect 389382 677898 389414 678134
rect 388794 642454 389414 677898
rect 388794 642218 388826 642454
rect 389062 642218 389146 642454
rect 389382 642218 389414 642454
rect 388794 642134 389414 642218
rect 388794 641898 388826 642134
rect 389062 641898 389146 642134
rect 389382 641898 389414 642134
rect 388794 606454 389414 641898
rect 388794 606218 388826 606454
rect 389062 606218 389146 606454
rect 389382 606218 389414 606454
rect 388794 606134 389414 606218
rect 388794 605898 388826 606134
rect 389062 605898 389146 606134
rect 389382 605898 389414 606134
rect 388794 570454 389414 605898
rect 388794 570218 388826 570454
rect 389062 570218 389146 570454
rect 389382 570218 389414 570454
rect 388794 570134 389414 570218
rect 388794 569898 388826 570134
rect 389062 569898 389146 570134
rect 389382 569898 389414 570134
rect 388794 534454 389414 569898
rect 388794 534218 388826 534454
rect 389062 534218 389146 534454
rect 389382 534218 389414 534454
rect 388794 534134 389414 534218
rect 388794 533898 388826 534134
rect 389062 533898 389146 534134
rect 389382 533898 389414 534134
rect 388794 498454 389414 533898
rect 388794 498218 388826 498454
rect 389062 498218 389146 498454
rect 389382 498218 389414 498454
rect 388794 498134 389414 498218
rect 388794 497898 388826 498134
rect 389062 497898 389146 498134
rect 389382 497898 389414 498134
rect 388794 462454 389414 497898
rect 388794 462218 388826 462454
rect 389062 462218 389146 462454
rect 389382 462218 389414 462454
rect 388794 462134 389414 462218
rect 388794 461898 388826 462134
rect 389062 461898 389146 462134
rect 389382 461898 389414 462134
rect 388794 426454 389414 461898
rect 388794 426218 388826 426454
rect 389062 426218 389146 426454
rect 389382 426218 389414 426454
rect 388794 426134 389414 426218
rect 388794 425898 388826 426134
rect 389062 425898 389146 426134
rect 389382 425898 389414 426134
rect 388794 390454 389414 425898
rect 388794 390218 388826 390454
rect 389062 390218 389146 390454
rect 389382 390218 389414 390454
rect 388794 390134 389414 390218
rect 388794 389898 388826 390134
rect 389062 389898 389146 390134
rect 389382 389898 389414 390134
rect 388794 354454 389414 389898
rect 388794 354218 388826 354454
rect 389062 354218 389146 354454
rect 389382 354218 389414 354454
rect 388794 354134 389414 354218
rect 388794 353898 388826 354134
rect 389062 353898 389146 354134
rect 389382 353898 389414 354134
rect 388794 318454 389414 353898
rect 388794 318218 388826 318454
rect 389062 318218 389146 318454
rect 389382 318218 389414 318454
rect 388794 318134 389414 318218
rect 388794 317898 388826 318134
rect 389062 317898 389146 318134
rect 389382 317898 389414 318134
rect 388794 282454 389414 317898
rect 388794 282218 388826 282454
rect 389062 282218 389146 282454
rect 389382 282218 389414 282454
rect 388794 282134 389414 282218
rect 388794 281898 388826 282134
rect 389062 281898 389146 282134
rect 389382 281898 389414 282134
rect 388794 246454 389414 281898
rect 388794 246218 388826 246454
rect 389062 246218 389146 246454
rect 389382 246218 389414 246454
rect 388794 246134 389414 246218
rect 388794 245898 388826 246134
rect 389062 245898 389146 246134
rect 389382 245898 389414 246134
rect 388794 210454 389414 245898
rect 388794 210218 388826 210454
rect 389062 210218 389146 210454
rect 389382 210218 389414 210454
rect 388794 210134 389414 210218
rect 388794 209898 388826 210134
rect 389062 209898 389146 210134
rect 389382 209898 389414 210134
rect 388794 174454 389414 209898
rect 388794 174218 388826 174454
rect 389062 174218 389146 174454
rect 389382 174218 389414 174454
rect 388794 174134 389414 174218
rect 388794 173898 388826 174134
rect 389062 173898 389146 174134
rect 389382 173898 389414 174134
rect 388794 138454 389414 173898
rect 388794 138218 388826 138454
rect 389062 138218 389146 138454
rect 389382 138218 389414 138454
rect 388794 138134 389414 138218
rect 388794 137898 388826 138134
rect 389062 137898 389146 138134
rect 389382 137898 389414 138134
rect 388794 102454 389414 137898
rect 388794 102218 388826 102454
rect 389062 102218 389146 102454
rect 389382 102218 389414 102454
rect 388794 102134 389414 102218
rect 388794 101898 388826 102134
rect 389062 101898 389146 102134
rect 389382 101898 389414 102134
rect 388794 66454 389414 101898
rect 388794 66218 388826 66454
rect 389062 66218 389146 66454
rect 389382 66218 389414 66454
rect 388794 66134 389414 66218
rect 388794 65898 388826 66134
rect 389062 65898 389146 66134
rect 389382 65898 389414 66134
rect 388794 30454 389414 65898
rect 388794 30218 388826 30454
rect 389062 30218 389146 30454
rect 389382 30218 389414 30454
rect 388794 30134 389414 30218
rect 388794 29898 388826 30134
rect 389062 29898 389146 30134
rect 389382 29898 389414 30134
rect 388794 -6106 389414 29898
rect 388794 -6342 388826 -6106
rect 389062 -6342 389146 -6106
rect 389382 -6342 389414 -6106
rect 388794 -6426 389414 -6342
rect 388794 -6662 388826 -6426
rect 389062 -6662 389146 -6426
rect 389382 -6662 389414 -6426
rect 388794 -7654 389414 -6662
rect 393294 711558 393914 711590
rect 393294 711322 393326 711558
rect 393562 711322 393646 711558
rect 393882 711322 393914 711558
rect 393294 711238 393914 711322
rect 393294 711002 393326 711238
rect 393562 711002 393646 711238
rect 393882 711002 393914 711238
rect 393294 682954 393914 711002
rect 393294 682718 393326 682954
rect 393562 682718 393646 682954
rect 393882 682718 393914 682954
rect 393294 682634 393914 682718
rect 393294 682398 393326 682634
rect 393562 682398 393646 682634
rect 393882 682398 393914 682634
rect 393294 646954 393914 682398
rect 393294 646718 393326 646954
rect 393562 646718 393646 646954
rect 393882 646718 393914 646954
rect 393294 646634 393914 646718
rect 393294 646398 393326 646634
rect 393562 646398 393646 646634
rect 393882 646398 393914 646634
rect 393294 610954 393914 646398
rect 393294 610718 393326 610954
rect 393562 610718 393646 610954
rect 393882 610718 393914 610954
rect 393294 610634 393914 610718
rect 393294 610398 393326 610634
rect 393562 610398 393646 610634
rect 393882 610398 393914 610634
rect 393294 574954 393914 610398
rect 393294 574718 393326 574954
rect 393562 574718 393646 574954
rect 393882 574718 393914 574954
rect 393294 574634 393914 574718
rect 393294 574398 393326 574634
rect 393562 574398 393646 574634
rect 393882 574398 393914 574634
rect 393294 538954 393914 574398
rect 393294 538718 393326 538954
rect 393562 538718 393646 538954
rect 393882 538718 393914 538954
rect 393294 538634 393914 538718
rect 393294 538398 393326 538634
rect 393562 538398 393646 538634
rect 393882 538398 393914 538634
rect 393294 502954 393914 538398
rect 393294 502718 393326 502954
rect 393562 502718 393646 502954
rect 393882 502718 393914 502954
rect 393294 502634 393914 502718
rect 393294 502398 393326 502634
rect 393562 502398 393646 502634
rect 393882 502398 393914 502634
rect 393294 466954 393914 502398
rect 393294 466718 393326 466954
rect 393562 466718 393646 466954
rect 393882 466718 393914 466954
rect 393294 466634 393914 466718
rect 393294 466398 393326 466634
rect 393562 466398 393646 466634
rect 393882 466398 393914 466634
rect 393294 430954 393914 466398
rect 393294 430718 393326 430954
rect 393562 430718 393646 430954
rect 393882 430718 393914 430954
rect 393294 430634 393914 430718
rect 393294 430398 393326 430634
rect 393562 430398 393646 430634
rect 393882 430398 393914 430634
rect 393294 394954 393914 430398
rect 393294 394718 393326 394954
rect 393562 394718 393646 394954
rect 393882 394718 393914 394954
rect 393294 394634 393914 394718
rect 393294 394398 393326 394634
rect 393562 394398 393646 394634
rect 393882 394398 393914 394634
rect 393294 358954 393914 394398
rect 393294 358718 393326 358954
rect 393562 358718 393646 358954
rect 393882 358718 393914 358954
rect 393294 358634 393914 358718
rect 393294 358398 393326 358634
rect 393562 358398 393646 358634
rect 393882 358398 393914 358634
rect 393294 322954 393914 358398
rect 393294 322718 393326 322954
rect 393562 322718 393646 322954
rect 393882 322718 393914 322954
rect 393294 322634 393914 322718
rect 393294 322398 393326 322634
rect 393562 322398 393646 322634
rect 393882 322398 393914 322634
rect 393294 286954 393914 322398
rect 393294 286718 393326 286954
rect 393562 286718 393646 286954
rect 393882 286718 393914 286954
rect 393294 286634 393914 286718
rect 393294 286398 393326 286634
rect 393562 286398 393646 286634
rect 393882 286398 393914 286634
rect 393294 250954 393914 286398
rect 393294 250718 393326 250954
rect 393562 250718 393646 250954
rect 393882 250718 393914 250954
rect 393294 250634 393914 250718
rect 393294 250398 393326 250634
rect 393562 250398 393646 250634
rect 393882 250398 393914 250634
rect 393294 214954 393914 250398
rect 393294 214718 393326 214954
rect 393562 214718 393646 214954
rect 393882 214718 393914 214954
rect 393294 214634 393914 214718
rect 393294 214398 393326 214634
rect 393562 214398 393646 214634
rect 393882 214398 393914 214634
rect 393294 178954 393914 214398
rect 393294 178718 393326 178954
rect 393562 178718 393646 178954
rect 393882 178718 393914 178954
rect 393294 178634 393914 178718
rect 393294 178398 393326 178634
rect 393562 178398 393646 178634
rect 393882 178398 393914 178634
rect 393294 142954 393914 178398
rect 393294 142718 393326 142954
rect 393562 142718 393646 142954
rect 393882 142718 393914 142954
rect 393294 142634 393914 142718
rect 393294 142398 393326 142634
rect 393562 142398 393646 142634
rect 393882 142398 393914 142634
rect 393294 106954 393914 142398
rect 393294 106718 393326 106954
rect 393562 106718 393646 106954
rect 393882 106718 393914 106954
rect 393294 106634 393914 106718
rect 393294 106398 393326 106634
rect 393562 106398 393646 106634
rect 393882 106398 393914 106634
rect 393294 70954 393914 106398
rect 393294 70718 393326 70954
rect 393562 70718 393646 70954
rect 393882 70718 393914 70954
rect 393294 70634 393914 70718
rect 393294 70398 393326 70634
rect 393562 70398 393646 70634
rect 393882 70398 393914 70634
rect 393294 34954 393914 70398
rect 393294 34718 393326 34954
rect 393562 34718 393646 34954
rect 393882 34718 393914 34954
rect 393294 34634 393914 34718
rect 393294 34398 393326 34634
rect 393562 34398 393646 34634
rect 393882 34398 393914 34634
rect 393294 -7066 393914 34398
rect 393294 -7302 393326 -7066
rect 393562 -7302 393646 -7066
rect 393882 -7302 393914 -7066
rect 393294 -7386 393914 -7302
rect 393294 -7622 393326 -7386
rect 393562 -7622 393646 -7386
rect 393882 -7622 393914 -7386
rect 393294 -7654 393914 -7622
rect 397794 704838 398414 711590
rect 397794 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 398414 704838
rect 397794 704518 398414 704602
rect 397794 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 398414 704518
rect 397794 687454 398414 704282
rect 397794 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 398414 687454
rect 397794 687134 398414 687218
rect 397794 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 398414 687134
rect 397794 651454 398414 686898
rect 397794 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 398414 651454
rect 397794 651134 398414 651218
rect 397794 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 398414 651134
rect 397794 615454 398414 650898
rect 397794 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 398414 615454
rect 397794 615134 398414 615218
rect 397794 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 398414 615134
rect 397794 579454 398414 614898
rect 397794 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 398414 579454
rect 397794 579134 398414 579218
rect 397794 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 398414 579134
rect 397794 543454 398414 578898
rect 397794 543218 397826 543454
rect 398062 543218 398146 543454
rect 398382 543218 398414 543454
rect 397794 543134 398414 543218
rect 397794 542898 397826 543134
rect 398062 542898 398146 543134
rect 398382 542898 398414 543134
rect 397794 507454 398414 542898
rect 397794 507218 397826 507454
rect 398062 507218 398146 507454
rect 398382 507218 398414 507454
rect 397794 507134 398414 507218
rect 397794 506898 397826 507134
rect 398062 506898 398146 507134
rect 398382 506898 398414 507134
rect 397794 471454 398414 506898
rect 397794 471218 397826 471454
rect 398062 471218 398146 471454
rect 398382 471218 398414 471454
rect 397794 471134 398414 471218
rect 397794 470898 397826 471134
rect 398062 470898 398146 471134
rect 398382 470898 398414 471134
rect 397794 435454 398414 470898
rect 397794 435218 397826 435454
rect 398062 435218 398146 435454
rect 398382 435218 398414 435454
rect 397794 435134 398414 435218
rect 397794 434898 397826 435134
rect 398062 434898 398146 435134
rect 398382 434898 398414 435134
rect 397794 399454 398414 434898
rect 397794 399218 397826 399454
rect 398062 399218 398146 399454
rect 398382 399218 398414 399454
rect 397794 399134 398414 399218
rect 397794 398898 397826 399134
rect 398062 398898 398146 399134
rect 398382 398898 398414 399134
rect 397794 363454 398414 398898
rect 397794 363218 397826 363454
rect 398062 363218 398146 363454
rect 398382 363218 398414 363454
rect 397794 363134 398414 363218
rect 397794 362898 397826 363134
rect 398062 362898 398146 363134
rect 398382 362898 398414 363134
rect 397794 327454 398414 362898
rect 397794 327218 397826 327454
rect 398062 327218 398146 327454
rect 398382 327218 398414 327454
rect 397794 327134 398414 327218
rect 397794 326898 397826 327134
rect 398062 326898 398146 327134
rect 398382 326898 398414 327134
rect 397794 291454 398414 326898
rect 397794 291218 397826 291454
rect 398062 291218 398146 291454
rect 398382 291218 398414 291454
rect 397794 291134 398414 291218
rect 397794 290898 397826 291134
rect 398062 290898 398146 291134
rect 398382 290898 398414 291134
rect 397794 255454 398414 290898
rect 397794 255218 397826 255454
rect 398062 255218 398146 255454
rect 398382 255218 398414 255454
rect 397794 255134 398414 255218
rect 397794 254898 397826 255134
rect 398062 254898 398146 255134
rect 398382 254898 398414 255134
rect 397794 219454 398414 254898
rect 397794 219218 397826 219454
rect 398062 219218 398146 219454
rect 398382 219218 398414 219454
rect 397794 219134 398414 219218
rect 397794 218898 397826 219134
rect 398062 218898 398146 219134
rect 398382 218898 398414 219134
rect 397794 183454 398414 218898
rect 397794 183218 397826 183454
rect 398062 183218 398146 183454
rect 398382 183218 398414 183454
rect 397794 183134 398414 183218
rect 397794 182898 397826 183134
rect 398062 182898 398146 183134
rect 398382 182898 398414 183134
rect 397794 147454 398414 182898
rect 397794 147218 397826 147454
rect 398062 147218 398146 147454
rect 398382 147218 398414 147454
rect 397794 147134 398414 147218
rect 397794 146898 397826 147134
rect 398062 146898 398146 147134
rect 398382 146898 398414 147134
rect 397794 111454 398414 146898
rect 397794 111218 397826 111454
rect 398062 111218 398146 111454
rect 398382 111218 398414 111454
rect 397794 111134 398414 111218
rect 397794 110898 397826 111134
rect 398062 110898 398146 111134
rect 398382 110898 398414 111134
rect 397794 75454 398414 110898
rect 397794 75218 397826 75454
rect 398062 75218 398146 75454
rect 398382 75218 398414 75454
rect 397794 75134 398414 75218
rect 397794 74898 397826 75134
rect 398062 74898 398146 75134
rect 398382 74898 398414 75134
rect 397794 39454 398414 74898
rect 397794 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 398414 39454
rect 397794 39134 398414 39218
rect 397794 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 398414 39134
rect 397794 3454 398414 38898
rect 397794 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 398414 3454
rect 397794 3134 398414 3218
rect 397794 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 398414 3134
rect 397794 -346 398414 2898
rect 397794 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 398414 -346
rect 397794 -666 398414 -582
rect 397794 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 398414 -666
rect 397794 -7654 398414 -902
rect 402294 705798 402914 711590
rect 402294 705562 402326 705798
rect 402562 705562 402646 705798
rect 402882 705562 402914 705798
rect 402294 705478 402914 705562
rect 402294 705242 402326 705478
rect 402562 705242 402646 705478
rect 402882 705242 402914 705478
rect 402294 691954 402914 705242
rect 402294 691718 402326 691954
rect 402562 691718 402646 691954
rect 402882 691718 402914 691954
rect 402294 691634 402914 691718
rect 402294 691398 402326 691634
rect 402562 691398 402646 691634
rect 402882 691398 402914 691634
rect 402294 655954 402914 691398
rect 402294 655718 402326 655954
rect 402562 655718 402646 655954
rect 402882 655718 402914 655954
rect 402294 655634 402914 655718
rect 402294 655398 402326 655634
rect 402562 655398 402646 655634
rect 402882 655398 402914 655634
rect 402294 619954 402914 655398
rect 402294 619718 402326 619954
rect 402562 619718 402646 619954
rect 402882 619718 402914 619954
rect 402294 619634 402914 619718
rect 402294 619398 402326 619634
rect 402562 619398 402646 619634
rect 402882 619398 402914 619634
rect 402294 583954 402914 619398
rect 402294 583718 402326 583954
rect 402562 583718 402646 583954
rect 402882 583718 402914 583954
rect 402294 583634 402914 583718
rect 402294 583398 402326 583634
rect 402562 583398 402646 583634
rect 402882 583398 402914 583634
rect 402294 547954 402914 583398
rect 402294 547718 402326 547954
rect 402562 547718 402646 547954
rect 402882 547718 402914 547954
rect 402294 547634 402914 547718
rect 402294 547398 402326 547634
rect 402562 547398 402646 547634
rect 402882 547398 402914 547634
rect 402294 511954 402914 547398
rect 402294 511718 402326 511954
rect 402562 511718 402646 511954
rect 402882 511718 402914 511954
rect 402294 511634 402914 511718
rect 402294 511398 402326 511634
rect 402562 511398 402646 511634
rect 402882 511398 402914 511634
rect 402294 475954 402914 511398
rect 402294 475718 402326 475954
rect 402562 475718 402646 475954
rect 402882 475718 402914 475954
rect 402294 475634 402914 475718
rect 402294 475398 402326 475634
rect 402562 475398 402646 475634
rect 402882 475398 402914 475634
rect 402294 439954 402914 475398
rect 402294 439718 402326 439954
rect 402562 439718 402646 439954
rect 402882 439718 402914 439954
rect 402294 439634 402914 439718
rect 402294 439398 402326 439634
rect 402562 439398 402646 439634
rect 402882 439398 402914 439634
rect 402294 403954 402914 439398
rect 402294 403718 402326 403954
rect 402562 403718 402646 403954
rect 402882 403718 402914 403954
rect 402294 403634 402914 403718
rect 402294 403398 402326 403634
rect 402562 403398 402646 403634
rect 402882 403398 402914 403634
rect 402294 367954 402914 403398
rect 402294 367718 402326 367954
rect 402562 367718 402646 367954
rect 402882 367718 402914 367954
rect 402294 367634 402914 367718
rect 402294 367398 402326 367634
rect 402562 367398 402646 367634
rect 402882 367398 402914 367634
rect 402294 331954 402914 367398
rect 402294 331718 402326 331954
rect 402562 331718 402646 331954
rect 402882 331718 402914 331954
rect 402294 331634 402914 331718
rect 402294 331398 402326 331634
rect 402562 331398 402646 331634
rect 402882 331398 402914 331634
rect 402294 295954 402914 331398
rect 402294 295718 402326 295954
rect 402562 295718 402646 295954
rect 402882 295718 402914 295954
rect 402294 295634 402914 295718
rect 402294 295398 402326 295634
rect 402562 295398 402646 295634
rect 402882 295398 402914 295634
rect 402294 259954 402914 295398
rect 402294 259718 402326 259954
rect 402562 259718 402646 259954
rect 402882 259718 402914 259954
rect 402294 259634 402914 259718
rect 402294 259398 402326 259634
rect 402562 259398 402646 259634
rect 402882 259398 402914 259634
rect 402294 223954 402914 259398
rect 402294 223718 402326 223954
rect 402562 223718 402646 223954
rect 402882 223718 402914 223954
rect 402294 223634 402914 223718
rect 402294 223398 402326 223634
rect 402562 223398 402646 223634
rect 402882 223398 402914 223634
rect 402294 187954 402914 223398
rect 402294 187718 402326 187954
rect 402562 187718 402646 187954
rect 402882 187718 402914 187954
rect 402294 187634 402914 187718
rect 402294 187398 402326 187634
rect 402562 187398 402646 187634
rect 402882 187398 402914 187634
rect 402294 151954 402914 187398
rect 402294 151718 402326 151954
rect 402562 151718 402646 151954
rect 402882 151718 402914 151954
rect 402294 151634 402914 151718
rect 402294 151398 402326 151634
rect 402562 151398 402646 151634
rect 402882 151398 402914 151634
rect 402294 115954 402914 151398
rect 402294 115718 402326 115954
rect 402562 115718 402646 115954
rect 402882 115718 402914 115954
rect 402294 115634 402914 115718
rect 402294 115398 402326 115634
rect 402562 115398 402646 115634
rect 402882 115398 402914 115634
rect 402294 79954 402914 115398
rect 402294 79718 402326 79954
rect 402562 79718 402646 79954
rect 402882 79718 402914 79954
rect 402294 79634 402914 79718
rect 402294 79398 402326 79634
rect 402562 79398 402646 79634
rect 402882 79398 402914 79634
rect 402294 43954 402914 79398
rect 402294 43718 402326 43954
rect 402562 43718 402646 43954
rect 402882 43718 402914 43954
rect 402294 43634 402914 43718
rect 402294 43398 402326 43634
rect 402562 43398 402646 43634
rect 402882 43398 402914 43634
rect 402294 7954 402914 43398
rect 402294 7718 402326 7954
rect 402562 7718 402646 7954
rect 402882 7718 402914 7954
rect 402294 7634 402914 7718
rect 402294 7398 402326 7634
rect 402562 7398 402646 7634
rect 402882 7398 402914 7634
rect 402294 -1306 402914 7398
rect 402294 -1542 402326 -1306
rect 402562 -1542 402646 -1306
rect 402882 -1542 402914 -1306
rect 402294 -1626 402914 -1542
rect 402294 -1862 402326 -1626
rect 402562 -1862 402646 -1626
rect 402882 -1862 402914 -1626
rect 402294 -7654 402914 -1862
rect 406794 706758 407414 711590
rect 406794 706522 406826 706758
rect 407062 706522 407146 706758
rect 407382 706522 407414 706758
rect 406794 706438 407414 706522
rect 406794 706202 406826 706438
rect 407062 706202 407146 706438
rect 407382 706202 407414 706438
rect 406794 696454 407414 706202
rect 406794 696218 406826 696454
rect 407062 696218 407146 696454
rect 407382 696218 407414 696454
rect 406794 696134 407414 696218
rect 406794 695898 406826 696134
rect 407062 695898 407146 696134
rect 407382 695898 407414 696134
rect 406794 660454 407414 695898
rect 406794 660218 406826 660454
rect 407062 660218 407146 660454
rect 407382 660218 407414 660454
rect 406794 660134 407414 660218
rect 406794 659898 406826 660134
rect 407062 659898 407146 660134
rect 407382 659898 407414 660134
rect 406794 624454 407414 659898
rect 406794 624218 406826 624454
rect 407062 624218 407146 624454
rect 407382 624218 407414 624454
rect 406794 624134 407414 624218
rect 406794 623898 406826 624134
rect 407062 623898 407146 624134
rect 407382 623898 407414 624134
rect 406794 588454 407414 623898
rect 406794 588218 406826 588454
rect 407062 588218 407146 588454
rect 407382 588218 407414 588454
rect 406794 588134 407414 588218
rect 406794 587898 406826 588134
rect 407062 587898 407146 588134
rect 407382 587898 407414 588134
rect 406794 552454 407414 587898
rect 406794 552218 406826 552454
rect 407062 552218 407146 552454
rect 407382 552218 407414 552454
rect 406794 552134 407414 552218
rect 406794 551898 406826 552134
rect 407062 551898 407146 552134
rect 407382 551898 407414 552134
rect 406794 516454 407414 551898
rect 406794 516218 406826 516454
rect 407062 516218 407146 516454
rect 407382 516218 407414 516454
rect 406794 516134 407414 516218
rect 406794 515898 406826 516134
rect 407062 515898 407146 516134
rect 407382 515898 407414 516134
rect 406794 480454 407414 515898
rect 406794 480218 406826 480454
rect 407062 480218 407146 480454
rect 407382 480218 407414 480454
rect 406794 480134 407414 480218
rect 406794 479898 406826 480134
rect 407062 479898 407146 480134
rect 407382 479898 407414 480134
rect 406794 444454 407414 479898
rect 406794 444218 406826 444454
rect 407062 444218 407146 444454
rect 407382 444218 407414 444454
rect 406794 444134 407414 444218
rect 406794 443898 406826 444134
rect 407062 443898 407146 444134
rect 407382 443898 407414 444134
rect 406794 408454 407414 443898
rect 406794 408218 406826 408454
rect 407062 408218 407146 408454
rect 407382 408218 407414 408454
rect 406794 408134 407414 408218
rect 406794 407898 406826 408134
rect 407062 407898 407146 408134
rect 407382 407898 407414 408134
rect 406794 372454 407414 407898
rect 406794 372218 406826 372454
rect 407062 372218 407146 372454
rect 407382 372218 407414 372454
rect 406794 372134 407414 372218
rect 406794 371898 406826 372134
rect 407062 371898 407146 372134
rect 407382 371898 407414 372134
rect 406794 336454 407414 371898
rect 406794 336218 406826 336454
rect 407062 336218 407146 336454
rect 407382 336218 407414 336454
rect 406794 336134 407414 336218
rect 406794 335898 406826 336134
rect 407062 335898 407146 336134
rect 407382 335898 407414 336134
rect 406794 300454 407414 335898
rect 406794 300218 406826 300454
rect 407062 300218 407146 300454
rect 407382 300218 407414 300454
rect 406794 300134 407414 300218
rect 406794 299898 406826 300134
rect 407062 299898 407146 300134
rect 407382 299898 407414 300134
rect 406794 264454 407414 299898
rect 406794 264218 406826 264454
rect 407062 264218 407146 264454
rect 407382 264218 407414 264454
rect 406794 264134 407414 264218
rect 406794 263898 406826 264134
rect 407062 263898 407146 264134
rect 407382 263898 407414 264134
rect 406794 228454 407414 263898
rect 406794 228218 406826 228454
rect 407062 228218 407146 228454
rect 407382 228218 407414 228454
rect 406794 228134 407414 228218
rect 406794 227898 406826 228134
rect 407062 227898 407146 228134
rect 407382 227898 407414 228134
rect 406794 192454 407414 227898
rect 406794 192218 406826 192454
rect 407062 192218 407146 192454
rect 407382 192218 407414 192454
rect 406794 192134 407414 192218
rect 406794 191898 406826 192134
rect 407062 191898 407146 192134
rect 407382 191898 407414 192134
rect 406794 156454 407414 191898
rect 406794 156218 406826 156454
rect 407062 156218 407146 156454
rect 407382 156218 407414 156454
rect 406794 156134 407414 156218
rect 406794 155898 406826 156134
rect 407062 155898 407146 156134
rect 407382 155898 407414 156134
rect 406794 120454 407414 155898
rect 406794 120218 406826 120454
rect 407062 120218 407146 120454
rect 407382 120218 407414 120454
rect 406794 120134 407414 120218
rect 406794 119898 406826 120134
rect 407062 119898 407146 120134
rect 407382 119898 407414 120134
rect 406794 84454 407414 119898
rect 406794 84218 406826 84454
rect 407062 84218 407146 84454
rect 407382 84218 407414 84454
rect 406794 84134 407414 84218
rect 406794 83898 406826 84134
rect 407062 83898 407146 84134
rect 407382 83898 407414 84134
rect 406794 48454 407414 83898
rect 406794 48218 406826 48454
rect 407062 48218 407146 48454
rect 407382 48218 407414 48454
rect 406794 48134 407414 48218
rect 406794 47898 406826 48134
rect 407062 47898 407146 48134
rect 407382 47898 407414 48134
rect 406794 12454 407414 47898
rect 406794 12218 406826 12454
rect 407062 12218 407146 12454
rect 407382 12218 407414 12454
rect 406794 12134 407414 12218
rect 406794 11898 406826 12134
rect 407062 11898 407146 12134
rect 407382 11898 407414 12134
rect 406794 -2266 407414 11898
rect 406794 -2502 406826 -2266
rect 407062 -2502 407146 -2266
rect 407382 -2502 407414 -2266
rect 406794 -2586 407414 -2502
rect 406794 -2822 406826 -2586
rect 407062 -2822 407146 -2586
rect 407382 -2822 407414 -2586
rect 406794 -7654 407414 -2822
rect 411294 707718 411914 711590
rect 411294 707482 411326 707718
rect 411562 707482 411646 707718
rect 411882 707482 411914 707718
rect 411294 707398 411914 707482
rect 411294 707162 411326 707398
rect 411562 707162 411646 707398
rect 411882 707162 411914 707398
rect 411294 700954 411914 707162
rect 411294 700718 411326 700954
rect 411562 700718 411646 700954
rect 411882 700718 411914 700954
rect 411294 700634 411914 700718
rect 411294 700398 411326 700634
rect 411562 700398 411646 700634
rect 411882 700398 411914 700634
rect 411294 664954 411914 700398
rect 411294 664718 411326 664954
rect 411562 664718 411646 664954
rect 411882 664718 411914 664954
rect 411294 664634 411914 664718
rect 411294 664398 411326 664634
rect 411562 664398 411646 664634
rect 411882 664398 411914 664634
rect 411294 628954 411914 664398
rect 411294 628718 411326 628954
rect 411562 628718 411646 628954
rect 411882 628718 411914 628954
rect 411294 628634 411914 628718
rect 411294 628398 411326 628634
rect 411562 628398 411646 628634
rect 411882 628398 411914 628634
rect 411294 592954 411914 628398
rect 411294 592718 411326 592954
rect 411562 592718 411646 592954
rect 411882 592718 411914 592954
rect 411294 592634 411914 592718
rect 411294 592398 411326 592634
rect 411562 592398 411646 592634
rect 411882 592398 411914 592634
rect 411294 556954 411914 592398
rect 411294 556718 411326 556954
rect 411562 556718 411646 556954
rect 411882 556718 411914 556954
rect 411294 556634 411914 556718
rect 411294 556398 411326 556634
rect 411562 556398 411646 556634
rect 411882 556398 411914 556634
rect 411294 520954 411914 556398
rect 411294 520718 411326 520954
rect 411562 520718 411646 520954
rect 411882 520718 411914 520954
rect 411294 520634 411914 520718
rect 411294 520398 411326 520634
rect 411562 520398 411646 520634
rect 411882 520398 411914 520634
rect 411294 484954 411914 520398
rect 411294 484718 411326 484954
rect 411562 484718 411646 484954
rect 411882 484718 411914 484954
rect 411294 484634 411914 484718
rect 411294 484398 411326 484634
rect 411562 484398 411646 484634
rect 411882 484398 411914 484634
rect 411294 448954 411914 484398
rect 411294 448718 411326 448954
rect 411562 448718 411646 448954
rect 411882 448718 411914 448954
rect 411294 448634 411914 448718
rect 411294 448398 411326 448634
rect 411562 448398 411646 448634
rect 411882 448398 411914 448634
rect 411294 412954 411914 448398
rect 411294 412718 411326 412954
rect 411562 412718 411646 412954
rect 411882 412718 411914 412954
rect 411294 412634 411914 412718
rect 411294 412398 411326 412634
rect 411562 412398 411646 412634
rect 411882 412398 411914 412634
rect 411294 376954 411914 412398
rect 411294 376718 411326 376954
rect 411562 376718 411646 376954
rect 411882 376718 411914 376954
rect 411294 376634 411914 376718
rect 411294 376398 411326 376634
rect 411562 376398 411646 376634
rect 411882 376398 411914 376634
rect 411294 340954 411914 376398
rect 411294 340718 411326 340954
rect 411562 340718 411646 340954
rect 411882 340718 411914 340954
rect 411294 340634 411914 340718
rect 411294 340398 411326 340634
rect 411562 340398 411646 340634
rect 411882 340398 411914 340634
rect 411294 304954 411914 340398
rect 411294 304718 411326 304954
rect 411562 304718 411646 304954
rect 411882 304718 411914 304954
rect 411294 304634 411914 304718
rect 411294 304398 411326 304634
rect 411562 304398 411646 304634
rect 411882 304398 411914 304634
rect 411294 268954 411914 304398
rect 411294 268718 411326 268954
rect 411562 268718 411646 268954
rect 411882 268718 411914 268954
rect 411294 268634 411914 268718
rect 411294 268398 411326 268634
rect 411562 268398 411646 268634
rect 411882 268398 411914 268634
rect 411294 232954 411914 268398
rect 411294 232718 411326 232954
rect 411562 232718 411646 232954
rect 411882 232718 411914 232954
rect 411294 232634 411914 232718
rect 411294 232398 411326 232634
rect 411562 232398 411646 232634
rect 411882 232398 411914 232634
rect 411294 196954 411914 232398
rect 411294 196718 411326 196954
rect 411562 196718 411646 196954
rect 411882 196718 411914 196954
rect 411294 196634 411914 196718
rect 411294 196398 411326 196634
rect 411562 196398 411646 196634
rect 411882 196398 411914 196634
rect 411294 160954 411914 196398
rect 411294 160718 411326 160954
rect 411562 160718 411646 160954
rect 411882 160718 411914 160954
rect 411294 160634 411914 160718
rect 411294 160398 411326 160634
rect 411562 160398 411646 160634
rect 411882 160398 411914 160634
rect 411294 124954 411914 160398
rect 411294 124718 411326 124954
rect 411562 124718 411646 124954
rect 411882 124718 411914 124954
rect 411294 124634 411914 124718
rect 411294 124398 411326 124634
rect 411562 124398 411646 124634
rect 411882 124398 411914 124634
rect 411294 88954 411914 124398
rect 411294 88718 411326 88954
rect 411562 88718 411646 88954
rect 411882 88718 411914 88954
rect 411294 88634 411914 88718
rect 411294 88398 411326 88634
rect 411562 88398 411646 88634
rect 411882 88398 411914 88634
rect 411294 52954 411914 88398
rect 411294 52718 411326 52954
rect 411562 52718 411646 52954
rect 411882 52718 411914 52954
rect 411294 52634 411914 52718
rect 411294 52398 411326 52634
rect 411562 52398 411646 52634
rect 411882 52398 411914 52634
rect 411294 16954 411914 52398
rect 411294 16718 411326 16954
rect 411562 16718 411646 16954
rect 411882 16718 411914 16954
rect 411294 16634 411914 16718
rect 411294 16398 411326 16634
rect 411562 16398 411646 16634
rect 411882 16398 411914 16634
rect 411294 -3226 411914 16398
rect 411294 -3462 411326 -3226
rect 411562 -3462 411646 -3226
rect 411882 -3462 411914 -3226
rect 411294 -3546 411914 -3462
rect 411294 -3782 411326 -3546
rect 411562 -3782 411646 -3546
rect 411882 -3782 411914 -3546
rect 411294 -7654 411914 -3782
rect 415794 708678 416414 711590
rect 415794 708442 415826 708678
rect 416062 708442 416146 708678
rect 416382 708442 416414 708678
rect 415794 708358 416414 708442
rect 415794 708122 415826 708358
rect 416062 708122 416146 708358
rect 416382 708122 416414 708358
rect 415794 669454 416414 708122
rect 415794 669218 415826 669454
rect 416062 669218 416146 669454
rect 416382 669218 416414 669454
rect 415794 669134 416414 669218
rect 415794 668898 415826 669134
rect 416062 668898 416146 669134
rect 416382 668898 416414 669134
rect 415794 633454 416414 668898
rect 415794 633218 415826 633454
rect 416062 633218 416146 633454
rect 416382 633218 416414 633454
rect 415794 633134 416414 633218
rect 415794 632898 415826 633134
rect 416062 632898 416146 633134
rect 416382 632898 416414 633134
rect 415794 597454 416414 632898
rect 415794 597218 415826 597454
rect 416062 597218 416146 597454
rect 416382 597218 416414 597454
rect 415794 597134 416414 597218
rect 415794 596898 415826 597134
rect 416062 596898 416146 597134
rect 416382 596898 416414 597134
rect 415794 561454 416414 596898
rect 415794 561218 415826 561454
rect 416062 561218 416146 561454
rect 416382 561218 416414 561454
rect 415794 561134 416414 561218
rect 415794 560898 415826 561134
rect 416062 560898 416146 561134
rect 416382 560898 416414 561134
rect 415794 525454 416414 560898
rect 415794 525218 415826 525454
rect 416062 525218 416146 525454
rect 416382 525218 416414 525454
rect 415794 525134 416414 525218
rect 415794 524898 415826 525134
rect 416062 524898 416146 525134
rect 416382 524898 416414 525134
rect 415794 489454 416414 524898
rect 415794 489218 415826 489454
rect 416062 489218 416146 489454
rect 416382 489218 416414 489454
rect 415794 489134 416414 489218
rect 415794 488898 415826 489134
rect 416062 488898 416146 489134
rect 416382 488898 416414 489134
rect 415794 453454 416414 488898
rect 415794 453218 415826 453454
rect 416062 453218 416146 453454
rect 416382 453218 416414 453454
rect 415794 453134 416414 453218
rect 415794 452898 415826 453134
rect 416062 452898 416146 453134
rect 416382 452898 416414 453134
rect 415794 417454 416414 452898
rect 415794 417218 415826 417454
rect 416062 417218 416146 417454
rect 416382 417218 416414 417454
rect 415794 417134 416414 417218
rect 415794 416898 415826 417134
rect 416062 416898 416146 417134
rect 416382 416898 416414 417134
rect 415794 381454 416414 416898
rect 415794 381218 415826 381454
rect 416062 381218 416146 381454
rect 416382 381218 416414 381454
rect 415794 381134 416414 381218
rect 415794 380898 415826 381134
rect 416062 380898 416146 381134
rect 416382 380898 416414 381134
rect 415794 345454 416414 380898
rect 415794 345218 415826 345454
rect 416062 345218 416146 345454
rect 416382 345218 416414 345454
rect 415794 345134 416414 345218
rect 415794 344898 415826 345134
rect 416062 344898 416146 345134
rect 416382 344898 416414 345134
rect 415794 309454 416414 344898
rect 415794 309218 415826 309454
rect 416062 309218 416146 309454
rect 416382 309218 416414 309454
rect 415794 309134 416414 309218
rect 415794 308898 415826 309134
rect 416062 308898 416146 309134
rect 416382 308898 416414 309134
rect 415794 273454 416414 308898
rect 415794 273218 415826 273454
rect 416062 273218 416146 273454
rect 416382 273218 416414 273454
rect 415794 273134 416414 273218
rect 415794 272898 415826 273134
rect 416062 272898 416146 273134
rect 416382 272898 416414 273134
rect 415794 237454 416414 272898
rect 415794 237218 415826 237454
rect 416062 237218 416146 237454
rect 416382 237218 416414 237454
rect 415794 237134 416414 237218
rect 415794 236898 415826 237134
rect 416062 236898 416146 237134
rect 416382 236898 416414 237134
rect 415794 201454 416414 236898
rect 415794 201218 415826 201454
rect 416062 201218 416146 201454
rect 416382 201218 416414 201454
rect 415794 201134 416414 201218
rect 415794 200898 415826 201134
rect 416062 200898 416146 201134
rect 416382 200898 416414 201134
rect 415794 165454 416414 200898
rect 415794 165218 415826 165454
rect 416062 165218 416146 165454
rect 416382 165218 416414 165454
rect 415794 165134 416414 165218
rect 415794 164898 415826 165134
rect 416062 164898 416146 165134
rect 416382 164898 416414 165134
rect 415794 129454 416414 164898
rect 415794 129218 415826 129454
rect 416062 129218 416146 129454
rect 416382 129218 416414 129454
rect 415794 129134 416414 129218
rect 415794 128898 415826 129134
rect 416062 128898 416146 129134
rect 416382 128898 416414 129134
rect 415794 93454 416414 128898
rect 415794 93218 415826 93454
rect 416062 93218 416146 93454
rect 416382 93218 416414 93454
rect 415794 93134 416414 93218
rect 415794 92898 415826 93134
rect 416062 92898 416146 93134
rect 416382 92898 416414 93134
rect 415794 57454 416414 92898
rect 415794 57218 415826 57454
rect 416062 57218 416146 57454
rect 416382 57218 416414 57454
rect 415794 57134 416414 57218
rect 415794 56898 415826 57134
rect 416062 56898 416146 57134
rect 416382 56898 416414 57134
rect 415794 21454 416414 56898
rect 415794 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 416414 21454
rect 415794 21134 416414 21218
rect 415794 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 416414 21134
rect 415794 -4186 416414 20898
rect 415794 -4422 415826 -4186
rect 416062 -4422 416146 -4186
rect 416382 -4422 416414 -4186
rect 415794 -4506 416414 -4422
rect 415794 -4742 415826 -4506
rect 416062 -4742 416146 -4506
rect 416382 -4742 416414 -4506
rect 415794 -7654 416414 -4742
rect 420294 709638 420914 711590
rect 420294 709402 420326 709638
rect 420562 709402 420646 709638
rect 420882 709402 420914 709638
rect 420294 709318 420914 709402
rect 420294 709082 420326 709318
rect 420562 709082 420646 709318
rect 420882 709082 420914 709318
rect 420294 673954 420914 709082
rect 420294 673718 420326 673954
rect 420562 673718 420646 673954
rect 420882 673718 420914 673954
rect 420294 673634 420914 673718
rect 420294 673398 420326 673634
rect 420562 673398 420646 673634
rect 420882 673398 420914 673634
rect 420294 637954 420914 673398
rect 420294 637718 420326 637954
rect 420562 637718 420646 637954
rect 420882 637718 420914 637954
rect 420294 637634 420914 637718
rect 420294 637398 420326 637634
rect 420562 637398 420646 637634
rect 420882 637398 420914 637634
rect 420294 601954 420914 637398
rect 420294 601718 420326 601954
rect 420562 601718 420646 601954
rect 420882 601718 420914 601954
rect 420294 601634 420914 601718
rect 420294 601398 420326 601634
rect 420562 601398 420646 601634
rect 420882 601398 420914 601634
rect 420294 565954 420914 601398
rect 420294 565718 420326 565954
rect 420562 565718 420646 565954
rect 420882 565718 420914 565954
rect 420294 565634 420914 565718
rect 420294 565398 420326 565634
rect 420562 565398 420646 565634
rect 420882 565398 420914 565634
rect 420294 529954 420914 565398
rect 420294 529718 420326 529954
rect 420562 529718 420646 529954
rect 420882 529718 420914 529954
rect 420294 529634 420914 529718
rect 420294 529398 420326 529634
rect 420562 529398 420646 529634
rect 420882 529398 420914 529634
rect 420294 493954 420914 529398
rect 420294 493718 420326 493954
rect 420562 493718 420646 493954
rect 420882 493718 420914 493954
rect 420294 493634 420914 493718
rect 420294 493398 420326 493634
rect 420562 493398 420646 493634
rect 420882 493398 420914 493634
rect 420294 457954 420914 493398
rect 420294 457718 420326 457954
rect 420562 457718 420646 457954
rect 420882 457718 420914 457954
rect 420294 457634 420914 457718
rect 420294 457398 420326 457634
rect 420562 457398 420646 457634
rect 420882 457398 420914 457634
rect 420294 421954 420914 457398
rect 420294 421718 420326 421954
rect 420562 421718 420646 421954
rect 420882 421718 420914 421954
rect 420294 421634 420914 421718
rect 420294 421398 420326 421634
rect 420562 421398 420646 421634
rect 420882 421398 420914 421634
rect 420294 385954 420914 421398
rect 420294 385718 420326 385954
rect 420562 385718 420646 385954
rect 420882 385718 420914 385954
rect 420294 385634 420914 385718
rect 420294 385398 420326 385634
rect 420562 385398 420646 385634
rect 420882 385398 420914 385634
rect 420294 349954 420914 385398
rect 420294 349718 420326 349954
rect 420562 349718 420646 349954
rect 420882 349718 420914 349954
rect 420294 349634 420914 349718
rect 420294 349398 420326 349634
rect 420562 349398 420646 349634
rect 420882 349398 420914 349634
rect 420294 313954 420914 349398
rect 420294 313718 420326 313954
rect 420562 313718 420646 313954
rect 420882 313718 420914 313954
rect 420294 313634 420914 313718
rect 420294 313398 420326 313634
rect 420562 313398 420646 313634
rect 420882 313398 420914 313634
rect 420294 277954 420914 313398
rect 420294 277718 420326 277954
rect 420562 277718 420646 277954
rect 420882 277718 420914 277954
rect 420294 277634 420914 277718
rect 420294 277398 420326 277634
rect 420562 277398 420646 277634
rect 420882 277398 420914 277634
rect 420294 241954 420914 277398
rect 420294 241718 420326 241954
rect 420562 241718 420646 241954
rect 420882 241718 420914 241954
rect 420294 241634 420914 241718
rect 420294 241398 420326 241634
rect 420562 241398 420646 241634
rect 420882 241398 420914 241634
rect 420294 205954 420914 241398
rect 420294 205718 420326 205954
rect 420562 205718 420646 205954
rect 420882 205718 420914 205954
rect 420294 205634 420914 205718
rect 420294 205398 420326 205634
rect 420562 205398 420646 205634
rect 420882 205398 420914 205634
rect 420294 169954 420914 205398
rect 420294 169718 420326 169954
rect 420562 169718 420646 169954
rect 420882 169718 420914 169954
rect 420294 169634 420914 169718
rect 420294 169398 420326 169634
rect 420562 169398 420646 169634
rect 420882 169398 420914 169634
rect 420294 133954 420914 169398
rect 420294 133718 420326 133954
rect 420562 133718 420646 133954
rect 420882 133718 420914 133954
rect 420294 133634 420914 133718
rect 420294 133398 420326 133634
rect 420562 133398 420646 133634
rect 420882 133398 420914 133634
rect 420294 97954 420914 133398
rect 420294 97718 420326 97954
rect 420562 97718 420646 97954
rect 420882 97718 420914 97954
rect 420294 97634 420914 97718
rect 420294 97398 420326 97634
rect 420562 97398 420646 97634
rect 420882 97398 420914 97634
rect 420294 61954 420914 97398
rect 420294 61718 420326 61954
rect 420562 61718 420646 61954
rect 420882 61718 420914 61954
rect 420294 61634 420914 61718
rect 420294 61398 420326 61634
rect 420562 61398 420646 61634
rect 420882 61398 420914 61634
rect 420294 25954 420914 61398
rect 420294 25718 420326 25954
rect 420562 25718 420646 25954
rect 420882 25718 420914 25954
rect 420294 25634 420914 25718
rect 420294 25398 420326 25634
rect 420562 25398 420646 25634
rect 420882 25398 420914 25634
rect 420294 -5146 420914 25398
rect 420294 -5382 420326 -5146
rect 420562 -5382 420646 -5146
rect 420882 -5382 420914 -5146
rect 420294 -5466 420914 -5382
rect 420294 -5702 420326 -5466
rect 420562 -5702 420646 -5466
rect 420882 -5702 420914 -5466
rect 420294 -7654 420914 -5702
rect 424794 710598 425414 711590
rect 424794 710362 424826 710598
rect 425062 710362 425146 710598
rect 425382 710362 425414 710598
rect 424794 710278 425414 710362
rect 424794 710042 424826 710278
rect 425062 710042 425146 710278
rect 425382 710042 425414 710278
rect 424794 678454 425414 710042
rect 424794 678218 424826 678454
rect 425062 678218 425146 678454
rect 425382 678218 425414 678454
rect 424794 678134 425414 678218
rect 424794 677898 424826 678134
rect 425062 677898 425146 678134
rect 425382 677898 425414 678134
rect 424794 642454 425414 677898
rect 424794 642218 424826 642454
rect 425062 642218 425146 642454
rect 425382 642218 425414 642454
rect 424794 642134 425414 642218
rect 424794 641898 424826 642134
rect 425062 641898 425146 642134
rect 425382 641898 425414 642134
rect 424794 606454 425414 641898
rect 424794 606218 424826 606454
rect 425062 606218 425146 606454
rect 425382 606218 425414 606454
rect 424794 606134 425414 606218
rect 424794 605898 424826 606134
rect 425062 605898 425146 606134
rect 425382 605898 425414 606134
rect 424794 570454 425414 605898
rect 424794 570218 424826 570454
rect 425062 570218 425146 570454
rect 425382 570218 425414 570454
rect 424794 570134 425414 570218
rect 424794 569898 424826 570134
rect 425062 569898 425146 570134
rect 425382 569898 425414 570134
rect 424794 534454 425414 569898
rect 424794 534218 424826 534454
rect 425062 534218 425146 534454
rect 425382 534218 425414 534454
rect 424794 534134 425414 534218
rect 424794 533898 424826 534134
rect 425062 533898 425146 534134
rect 425382 533898 425414 534134
rect 424794 498454 425414 533898
rect 424794 498218 424826 498454
rect 425062 498218 425146 498454
rect 425382 498218 425414 498454
rect 424794 498134 425414 498218
rect 424794 497898 424826 498134
rect 425062 497898 425146 498134
rect 425382 497898 425414 498134
rect 424794 462454 425414 497898
rect 424794 462218 424826 462454
rect 425062 462218 425146 462454
rect 425382 462218 425414 462454
rect 424794 462134 425414 462218
rect 424794 461898 424826 462134
rect 425062 461898 425146 462134
rect 425382 461898 425414 462134
rect 424794 426454 425414 461898
rect 424794 426218 424826 426454
rect 425062 426218 425146 426454
rect 425382 426218 425414 426454
rect 424794 426134 425414 426218
rect 424794 425898 424826 426134
rect 425062 425898 425146 426134
rect 425382 425898 425414 426134
rect 424794 390454 425414 425898
rect 424794 390218 424826 390454
rect 425062 390218 425146 390454
rect 425382 390218 425414 390454
rect 424794 390134 425414 390218
rect 424794 389898 424826 390134
rect 425062 389898 425146 390134
rect 425382 389898 425414 390134
rect 424794 354454 425414 389898
rect 424794 354218 424826 354454
rect 425062 354218 425146 354454
rect 425382 354218 425414 354454
rect 424794 354134 425414 354218
rect 424794 353898 424826 354134
rect 425062 353898 425146 354134
rect 425382 353898 425414 354134
rect 424794 318454 425414 353898
rect 424794 318218 424826 318454
rect 425062 318218 425146 318454
rect 425382 318218 425414 318454
rect 424794 318134 425414 318218
rect 424794 317898 424826 318134
rect 425062 317898 425146 318134
rect 425382 317898 425414 318134
rect 424794 282454 425414 317898
rect 424794 282218 424826 282454
rect 425062 282218 425146 282454
rect 425382 282218 425414 282454
rect 424794 282134 425414 282218
rect 424794 281898 424826 282134
rect 425062 281898 425146 282134
rect 425382 281898 425414 282134
rect 424794 246454 425414 281898
rect 424794 246218 424826 246454
rect 425062 246218 425146 246454
rect 425382 246218 425414 246454
rect 424794 246134 425414 246218
rect 424794 245898 424826 246134
rect 425062 245898 425146 246134
rect 425382 245898 425414 246134
rect 424794 210454 425414 245898
rect 424794 210218 424826 210454
rect 425062 210218 425146 210454
rect 425382 210218 425414 210454
rect 424794 210134 425414 210218
rect 424794 209898 424826 210134
rect 425062 209898 425146 210134
rect 425382 209898 425414 210134
rect 424794 174454 425414 209898
rect 424794 174218 424826 174454
rect 425062 174218 425146 174454
rect 425382 174218 425414 174454
rect 424794 174134 425414 174218
rect 424794 173898 424826 174134
rect 425062 173898 425146 174134
rect 425382 173898 425414 174134
rect 424794 138454 425414 173898
rect 424794 138218 424826 138454
rect 425062 138218 425146 138454
rect 425382 138218 425414 138454
rect 424794 138134 425414 138218
rect 424794 137898 424826 138134
rect 425062 137898 425146 138134
rect 425382 137898 425414 138134
rect 424794 102454 425414 137898
rect 424794 102218 424826 102454
rect 425062 102218 425146 102454
rect 425382 102218 425414 102454
rect 424794 102134 425414 102218
rect 424794 101898 424826 102134
rect 425062 101898 425146 102134
rect 425382 101898 425414 102134
rect 424794 66454 425414 101898
rect 424794 66218 424826 66454
rect 425062 66218 425146 66454
rect 425382 66218 425414 66454
rect 424794 66134 425414 66218
rect 424794 65898 424826 66134
rect 425062 65898 425146 66134
rect 425382 65898 425414 66134
rect 424794 30454 425414 65898
rect 424794 30218 424826 30454
rect 425062 30218 425146 30454
rect 425382 30218 425414 30454
rect 424794 30134 425414 30218
rect 424794 29898 424826 30134
rect 425062 29898 425146 30134
rect 425382 29898 425414 30134
rect 424794 -6106 425414 29898
rect 424794 -6342 424826 -6106
rect 425062 -6342 425146 -6106
rect 425382 -6342 425414 -6106
rect 424794 -6426 425414 -6342
rect 424794 -6662 424826 -6426
rect 425062 -6662 425146 -6426
rect 425382 -6662 425414 -6426
rect 424794 -7654 425414 -6662
rect 429294 711558 429914 711590
rect 429294 711322 429326 711558
rect 429562 711322 429646 711558
rect 429882 711322 429914 711558
rect 429294 711238 429914 711322
rect 429294 711002 429326 711238
rect 429562 711002 429646 711238
rect 429882 711002 429914 711238
rect 429294 682954 429914 711002
rect 429294 682718 429326 682954
rect 429562 682718 429646 682954
rect 429882 682718 429914 682954
rect 429294 682634 429914 682718
rect 429294 682398 429326 682634
rect 429562 682398 429646 682634
rect 429882 682398 429914 682634
rect 429294 646954 429914 682398
rect 429294 646718 429326 646954
rect 429562 646718 429646 646954
rect 429882 646718 429914 646954
rect 429294 646634 429914 646718
rect 429294 646398 429326 646634
rect 429562 646398 429646 646634
rect 429882 646398 429914 646634
rect 429294 610954 429914 646398
rect 429294 610718 429326 610954
rect 429562 610718 429646 610954
rect 429882 610718 429914 610954
rect 429294 610634 429914 610718
rect 429294 610398 429326 610634
rect 429562 610398 429646 610634
rect 429882 610398 429914 610634
rect 429294 574954 429914 610398
rect 429294 574718 429326 574954
rect 429562 574718 429646 574954
rect 429882 574718 429914 574954
rect 429294 574634 429914 574718
rect 429294 574398 429326 574634
rect 429562 574398 429646 574634
rect 429882 574398 429914 574634
rect 429294 538954 429914 574398
rect 429294 538718 429326 538954
rect 429562 538718 429646 538954
rect 429882 538718 429914 538954
rect 429294 538634 429914 538718
rect 429294 538398 429326 538634
rect 429562 538398 429646 538634
rect 429882 538398 429914 538634
rect 429294 502954 429914 538398
rect 429294 502718 429326 502954
rect 429562 502718 429646 502954
rect 429882 502718 429914 502954
rect 429294 502634 429914 502718
rect 429294 502398 429326 502634
rect 429562 502398 429646 502634
rect 429882 502398 429914 502634
rect 429294 466954 429914 502398
rect 429294 466718 429326 466954
rect 429562 466718 429646 466954
rect 429882 466718 429914 466954
rect 429294 466634 429914 466718
rect 429294 466398 429326 466634
rect 429562 466398 429646 466634
rect 429882 466398 429914 466634
rect 429294 430954 429914 466398
rect 429294 430718 429326 430954
rect 429562 430718 429646 430954
rect 429882 430718 429914 430954
rect 429294 430634 429914 430718
rect 429294 430398 429326 430634
rect 429562 430398 429646 430634
rect 429882 430398 429914 430634
rect 429294 394954 429914 430398
rect 429294 394718 429326 394954
rect 429562 394718 429646 394954
rect 429882 394718 429914 394954
rect 429294 394634 429914 394718
rect 429294 394398 429326 394634
rect 429562 394398 429646 394634
rect 429882 394398 429914 394634
rect 429294 358954 429914 394398
rect 429294 358718 429326 358954
rect 429562 358718 429646 358954
rect 429882 358718 429914 358954
rect 429294 358634 429914 358718
rect 429294 358398 429326 358634
rect 429562 358398 429646 358634
rect 429882 358398 429914 358634
rect 429294 322954 429914 358398
rect 429294 322718 429326 322954
rect 429562 322718 429646 322954
rect 429882 322718 429914 322954
rect 429294 322634 429914 322718
rect 429294 322398 429326 322634
rect 429562 322398 429646 322634
rect 429882 322398 429914 322634
rect 429294 286954 429914 322398
rect 429294 286718 429326 286954
rect 429562 286718 429646 286954
rect 429882 286718 429914 286954
rect 429294 286634 429914 286718
rect 429294 286398 429326 286634
rect 429562 286398 429646 286634
rect 429882 286398 429914 286634
rect 429294 250954 429914 286398
rect 429294 250718 429326 250954
rect 429562 250718 429646 250954
rect 429882 250718 429914 250954
rect 429294 250634 429914 250718
rect 429294 250398 429326 250634
rect 429562 250398 429646 250634
rect 429882 250398 429914 250634
rect 429294 214954 429914 250398
rect 429294 214718 429326 214954
rect 429562 214718 429646 214954
rect 429882 214718 429914 214954
rect 429294 214634 429914 214718
rect 429294 214398 429326 214634
rect 429562 214398 429646 214634
rect 429882 214398 429914 214634
rect 429294 178954 429914 214398
rect 429294 178718 429326 178954
rect 429562 178718 429646 178954
rect 429882 178718 429914 178954
rect 429294 178634 429914 178718
rect 429294 178398 429326 178634
rect 429562 178398 429646 178634
rect 429882 178398 429914 178634
rect 429294 142954 429914 178398
rect 429294 142718 429326 142954
rect 429562 142718 429646 142954
rect 429882 142718 429914 142954
rect 429294 142634 429914 142718
rect 429294 142398 429326 142634
rect 429562 142398 429646 142634
rect 429882 142398 429914 142634
rect 429294 106954 429914 142398
rect 429294 106718 429326 106954
rect 429562 106718 429646 106954
rect 429882 106718 429914 106954
rect 429294 106634 429914 106718
rect 429294 106398 429326 106634
rect 429562 106398 429646 106634
rect 429882 106398 429914 106634
rect 429294 70954 429914 106398
rect 429294 70718 429326 70954
rect 429562 70718 429646 70954
rect 429882 70718 429914 70954
rect 429294 70634 429914 70718
rect 429294 70398 429326 70634
rect 429562 70398 429646 70634
rect 429882 70398 429914 70634
rect 429294 34954 429914 70398
rect 429294 34718 429326 34954
rect 429562 34718 429646 34954
rect 429882 34718 429914 34954
rect 429294 34634 429914 34718
rect 429294 34398 429326 34634
rect 429562 34398 429646 34634
rect 429882 34398 429914 34634
rect 429294 -7066 429914 34398
rect 429294 -7302 429326 -7066
rect 429562 -7302 429646 -7066
rect 429882 -7302 429914 -7066
rect 429294 -7386 429914 -7302
rect 429294 -7622 429326 -7386
rect 429562 -7622 429646 -7386
rect 429882 -7622 429914 -7386
rect 429294 -7654 429914 -7622
rect 433794 704838 434414 711590
rect 433794 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 434414 704838
rect 433794 704518 434414 704602
rect 433794 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 434414 704518
rect 433794 687454 434414 704282
rect 433794 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 434414 687454
rect 433794 687134 434414 687218
rect 433794 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 434414 687134
rect 433794 651454 434414 686898
rect 433794 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 434414 651454
rect 433794 651134 434414 651218
rect 433794 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 434414 651134
rect 433794 615454 434414 650898
rect 433794 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 434414 615454
rect 433794 615134 434414 615218
rect 433794 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 434414 615134
rect 433794 579454 434414 614898
rect 433794 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 434414 579454
rect 433794 579134 434414 579218
rect 433794 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 434414 579134
rect 433794 543454 434414 578898
rect 433794 543218 433826 543454
rect 434062 543218 434146 543454
rect 434382 543218 434414 543454
rect 433794 543134 434414 543218
rect 433794 542898 433826 543134
rect 434062 542898 434146 543134
rect 434382 542898 434414 543134
rect 433794 507454 434414 542898
rect 433794 507218 433826 507454
rect 434062 507218 434146 507454
rect 434382 507218 434414 507454
rect 433794 507134 434414 507218
rect 433794 506898 433826 507134
rect 434062 506898 434146 507134
rect 434382 506898 434414 507134
rect 433794 471454 434414 506898
rect 433794 471218 433826 471454
rect 434062 471218 434146 471454
rect 434382 471218 434414 471454
rect 433794 471134 434414 471218
rect 433794 470898 433826 471134
rect 434062 470898 434146 471134
rect 434382 470898 434414 471134
rect 433794 435454 434414 470898
rect 433794 435218 433826 435454
rect 434062 435218 434146 435454
rect 434382 435218 434414 435454
rect 433794 435134 434414 435218
rect 433794 434898 433826 435134
rect 434062 434898 434146 435134
rect 434382 434898 434414 435134
rect 433794 399454 434414 434898
rect 433794 399218 433826 399454
rect 434062 399218 434146 399454
rect 434382 399218 434414 399454
rect 433794 399134 434414 399218
rect 433794 398898 433826 399134
rect 434062 398898 434146 399134
rect 434382 398898 434414 399134
rect 433794 363454 434414 398898
rect 433794 363218 433826 363454
rect 434062 363218 434146 363454
rect 434382 363218 434414 363454
rect 433794 363134 434414 363218
rect 433794 362898 433826 363134
rect 434062 362898 434146 363134
rect 434382 362898 434414 363134
rect 433794 327454 434414 362898
rect 433794 327218 433826 327454
rect 434062 327218 434146 327454
rect 434382 327218 434414 327454
rect 433794 327134 434414 327218
rect 433794 326898 433826 327134
rect 434062 326898 434146 327134
rect 434382 326898 434414 327134
rect 433794 291454 434414 326898
rect 433794 291218 433826 291454
rect 434062 291218 434146 291454
rect 434382 291218 434414 291454
rect 433794 291134 434414 291218
rect 433794 290898 433826 291134
rect 434062 290898 434146 291134
rect 434382 290898 434414 291134
rect 433794 255454 434414 290898
rect 433794 255218 433826 255454
rect 434062 255218 434146 255454
rect 434382 255218 434414 255454
rect 433794 255134 434414 255218
rect 433794 254898 433826 255134
rect 434062 254898 434146 255134
rect 434382 254898 434414 255134
rect 433794 219454 434414 254898
rect 433794 219218 433826 219454
rect 434062 219218 434146 219454
rect 434382 219218 434414 219454
rect 433794 219134 434414 219218
rect 433794 218898 433826 219134
rect 434062 218898 434146 219134
rect 434382 218898 434414 219134
rect 433794 183454 434414 218898
rect 433794 183218 433826 183454
rect 434062 183218 434146 183454
rect 434382 183218 434414 183454
rect 433794 183134 434414 183218
rect 433794 182898 433826 183134
rect 434062 182898 434146 183134
rect 434382 182898 434414 183134
rect 433794 147454 434414 182898
rect 433794 147218 433826 147454
rect 434062 147218 434146 147454
rect 434382 147218 434414 147454
rect 433794 147134 434414 147218
rect 433794 146898 433826 147134
rect 434062 146898 434146 147134
rect 434382 146898 434414 147134
rect 433794 111454 434414 146898
rect 433794 111218 433826 111454
rect 434062 111218 434146 111454
rect 434382 111218 434414 111454
rect 433794 111134 434414 111218
rect 433794 110898 433826 111134
rect 434062 110898 434146 111134
rect 434382 110898 434414 111134
rect 433794 75454 434414 110898
rect 433794 75218 433826 75454
rect 434062 75218 434146 75454
rect 434382 75218 434414 75454
rect 433794 75134 434414 75218
rect 433794 74898 433826 75134
rect 434062 74898 434146 75134
rect 434382 74898 434414 75134
rect 433794 39454 434414 74898
rect 433794 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 434414 39454
rect 433794 39134 434414 39218
rect 433794 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 434414 39134
rect 433794 3454 434414 38898
rect 433794 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 434414 3454
rect 433794 3134 434414 3218
rect 433794 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 434414 3134
rect 433794 -346 434414 2898
rect 433794 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 434414 -346
rect 433794 -666 434414 -582
rect 433794 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 434414 -666
rect 433794 -7654 434414 -902
rect 438294 705798 438914 711590
rect 438294 705562 438326 705798
rect 438562 705562 438646 705798
rect 438882 705562 438914 705798
rect 438294 705478 438914 705562
rect 438294 705242 438326 705478
rect 438562 705242 438646 705478
rect 438882 705242 438914 705478
rect 438294 691954 438914 705242
rect 438294 691718 438326 691954
rect 438562 691718 438646 691954
rect 438882 691718 438914 691954
rect 438294 691634 438914 691718
rect 438294 691398 438326 691634
rect 438562 691398 438646 691634
rect 438882 691398 438914 691634
rect 438294 655954 438914 691398
rect 438294 655718 438326 655954
rect 438562 655718 438646 655954
rect 438882 655718 438914 655954
rect 438294 655634 438914 655718
rect 438294 655398 438326 655634
rect 438562 655398 438646 655634
rect 438882 655398 438914 655634
rect 438294 619954 438914 655398
rect 438294 619718 438326 619954
rect 438562 619718 438646 619954
rect 438882 619718 438914 619954
rect 438294 619634 438914 619718
rect 438294 619398 438326 619634
rect 438562 619398 438646 619634
rect 438882 619398 438914 619634
rect 438294 583954 438914 619398
rect 438294 583718 438326 583954
rect 438562 583718 438646 583954
rect 438882 583718 438914 583954
rect 438294 583634 438914 583718
rect 438294 583398 438326 583634
rect 438562 583398 438646 583634
rect 438882 583398 438914 583634
rect 438294 547954 438914 583398
rect 438294 547718 438326 547954
rect 438562 547718 438646 547954
rect 438882 547718 438914 547954
rect 438294 547634 438914 547718
rect 438294 547398 438326 547634
rect 438562 547398 438646 547634
rect 438882 547398 438914 547634
rect 438294 511954 438914 547398
rect 438294 511718 438326 511954
rect 438562 511718 438646 511954
rect 438882 511718 438914 511954
rect 438294 511634 438914 511718
rect 438294 511398 438326 511634
rect 438562 511398 438646 511634
rect 438882 511398 438914 511634
rect 438294 475954 438914 511398
rect 438294 475718 438326 475954
rect 438562 475718 438646 475954
rect 438882 475718 438914 475954
rect 438294 475634 438914 475718
rect 438294 475398 438326 475634
rect 438562 475398 438646 475634
rect 438882 475398 438914 475634
rect 438294 439954 438914 475398
rect 438294 439718 438326 439954
rect 438562 439718 438646 439954
rect 438882 439718 438914 439954
rect 438294 439634 438914 439718
rect 438294 439398 438326 439634
rect 438562 439398 438646 439634
rect 438882 439398 438914 439634
rect 438294 403954 438914 439398
rect 438294 403718 438326 403954
rect 438562 403718 438646 403954
rect 438882 403718 438914 403954
rect 438294 403634 438914 403718
rect 438294 403398 438326 403634
rect 438562 403398 438646 403634
rect 438882 403398 438914 403634
rect 438294 367954 438914 403398
rect 438294 367718 438326 367954
rect 438562 367718 438646 367954
rect 438882 367718 438914 367954
rect 438294 367634 438914 367718
rect 438294 367398 438326 367634
rect 438562 367398 438646 367634
rect 438882 367398 438914 367634
rect 438294 331954 438914 367398
rect 438294 331718 438326 331954
rect 438562 331718 438646 331954
rect 438882 331718 438914 331954
rect 438294 331634 438914 331718
rect 438294 331398 438326 331634
rect 438562 331398 438646 331634
rect 438882 331398 438914 331634
rect 438294 295954 438914 331398
rect 438294 295718 438326 295954
rect 438562 295718 438646 295954
rect 438882 295718 438914 295954
rect 438294 295634 438914 295718
rect 438294 295398 438326 295634
rect 438562 295398 438646 295634
rect 438882 295398 438914 295634
rect 438294 259954 438914 295398
rect 438294 259718 438326 259954
rect 438562 259718 438646 259954
rect 438882 259718 438914 259954
rect 438294 259634 438914 259718
rect 438294 259398 438326 259634
rect 438562 259398 438646 259634
rect 438882 259398 438914 259634
rect 438294 223954 438914 259398
rect 438294 223718 438326 223954
rect 438562 223718 438646 223954
rect 438882 223718 438914 223954
rect 438294 223634 438914 223718
rect 438294 223398 438326 223634
rect 438562 223398 438646 223634
rect 438882 223398 438914 223634
rect 438294 187954 438914 223398
rect 438294 187718 438326 187954
rect 438562 187718 438646 187954
rect 438882 187718 438914 187954
rect 438294 187634 438914 187718
rect 438294 187398 438326 187634
rect 438562 187398 438646 187634
rect 438882 187398 438914 187634
rect 438294 151954 438914 187398
rect 438294 151718 438326 151954
rect 438562 151718 438646 151954
rect 438882 151718 438914 151954
rect 438294 151634 438914 151718
rect 438294 151398 438326 151634
rect 438562 151398 438646 151634
rect 438882 151398 438914 151634
rect 438294 115954 438914 151398
rect 438294 115718 438326 115954
rect 438562 115718 438646 115954
rect 438882 115718 438914 115954
rect 438294 115634 438914 115718
rect 438294 115398 438326 115634
rect 438562 115398 438646 115634
rect 438882 115398 438914 115634
rect 438294 79954 438914 115398
rect 438294 79718 438326 79954
rect 438562 79718 438646 79954
rect 438882 79718 438914 79954
rect 438294 79634 438914 79718
rect 438294 79398 438326 79634
rect 438562 79398 438646 79634
rect 438882 79398 438914 79634
rect 438294 43954 438914 79398
rect 438294 43718 438326 43954
rect 438562 43718 438646 43954
rect 438882 43718 438914 43954
rect 438294 43634 438914 43718
rect 438294 43398 438326 43634
rect 438562 43398 438646 43634
rect 438882 43398 438914 43634
rect 438294 7954 438914 43398
rect 438294 7718 438326 7954
rect 438562 7718 438646 7954
rect 438882 7718 438914 7954
rect 438294 7634 438914 7718
rect 438294 7398 438326 7634
rect 438562 7398 438646 7634
rect 438882 7398 438914 7634
rect 438294 -1306 438914 7398
rect 438294 -1542 438326 -1306
rect 438562 -1542 438646 -1306
rect 438882 -1542 438914 -1306
rect 438294 -1626 438914 -1542
rect 438294 -1862 438326 -1626
rect 438562 -1862 438646 -1626
rect 438882 -1862 438914 -1626
rect 438294 -7654 438914 -1862
rect 442794 706758 443414 711590
rect 442794 706522 442826 706758
rect 443062 706522 443146 706758
rect 443382 706522 443414 706758
rect 442794 706438 443414 706522
rect 442794 706202 442826 706438
rect 443062 706202 443146 706438
rect 443382 706202 443414 706438
rect 442794 696454 443414 706202
rect 442794 696218 442826 696454
rect 443062 696218 443146 696454
rect 443382 696218 443414 696454
rect 442794 696134 443414 696218
rect 442794 695898 442826 696134
rect 443062 695898 443146 696134
rect 443382 695898 443414 696134
rect 442794 660454 443414 695898
rect 442794 660218 442826 660454
rect 443062 660218 443146 660454
rect 443382 660218 443414 660454
rect 442794 660134 443414 660218
rect 442794 659898 442826 660134
rect 443062 659898 443146 660134
rect 443382 659898 443414 660134
rect 442794 624454 443414 659898
rect 442794 624218 442826 624454
rect 443062 624218 443146 624454
rect 443382 624218 443414 624454
rect 442794 624134 443414 624218
rect 442794 623898 442826 624134
rect 443062 623898 443146 624134
rect 443382 623898 443414 624134
rect 442794 588454 443414 623898
rect 442794 588218 442826 588454
rect 443062 588218 443146 588454
rect 443382 588218 443414 588454
rect 442794 588134 443414 588218
rect 442794 587898 442826 588134
rect 443062 587898 443146 588134
rect 443382 587898 443414 588134
rect 442794 552454 443414 587898
rect 442794 552218 442826 552454
rect 443062 552218 443146 552454
rect 443382 552218 443414 552454
rect 442794 552134 443414 552218
rect 442794 551898 442826 552134
rect 443062 551898 443146 552134
rect 443382 551898 443414 552134
rect 442794 516454 443414 551898
rect 442794 516218 442826 516454
rect 443062 516218 443146 516454
rect 443382 516218 443414 516454
rect 442794 516134 443414 516218
rect 442794 515898 442826 516134
rect 443062 515898 443146 516134
rect 443382 515898 443414 516134
rect 442794 480454 443414 515898
rect 442794 480218 442826 480454
rect 443062 480218 443146 480454
rect 443382 480218 443414 480454
rect 442794 480134 443414 480218
rect 442794 479898 442826 480134
rect 443062 479898 443146 480134
rect 443382 479898 443414 480134
rect 442794 444454 443414 479898
rect 442794 444218 442826 444454
rect 443062 444218 443146 444454
rect 443382 444218 443414 444454
rect 442794 444134 443414 444218
rect 442794 443898 442826 444134
rect 443062 443898 443146 444134
rect 443382 443898 443414 444134
rect 442794 408454 443414 443898
rect 442794 408218 442826 408454
rect 443062 408218 443146 408454
rect 443382 408218 443414 408454
rect 442794 408134 443414 408218
rect 442794 407898 442826 408134
rect 443062 407898 443146 408134
rect 443382 407898 443414 408134
rect 442794 372454 443414 407898
rect 442794 372218 442826 372454
rect 443062 372218 443146 372454
rect 443382 372218 443414 372454
rect 442794 372134 443414 372218
rect 442794 371898 442826 372134
rect 443062 371898 443146 372134
rect 443382 371898 443414 372134
rect 442794 336454 443414 371898
rect 442794 336218 442826 336454
rect 443062 336218 443146 336454
rect 443382 336218 443414 336454
rect 442794 336134 443414 336218
rect 442794 335898 442826 336134
rect 443062 335898 443146 336134
rect 443382 335898 443414 336134
rect 442794 300454 443414 335898
rect 442794 300218 442826 300454
rect 443062 300218 443146 300454
rect 443382 300218 443414 300454
rect 442794 300134 443414 300218
rect 442794 299898 442826 300134
rect 443062 299898 443146 300134
rect 443382 299898 443414 300134
rect 442794 264454 443414 299898
rect 442794 264218 442826 264454
rect 443062 264218 443146 264454
rect 443382 264218 443414 264454
rect 442794 264134 443414 264218
rect 442794 263898 442826 264134
rect 443062 263898 443146 264134
rect 443382 263898 443414 264134
rect 442794 228454 443414 263898
rect 442794 228218 442826 228454
rect 443062 228218 443146 228454
rect 443382 228218 443414 228454
rect 442794 228134 443414 228218
rect 442794 227898 442826 228134
rect 443062 227898 443146 228134
rect 443382 227898 443414 228134
rect 442794 192454 443414 227898
rect 442794 192218 442826 192454
rect 443062 192218 443146 192454
rect 443382 192218 443414 192454
rect 442794 192134 443414 192218
rect 442794 191898 442826 192134
rect 443062 191898 443146 192134
rect 443382 191898 443414 192134
rect 442794 156454 443414 191898
rect 442794 156218 442826 156454
rect 443062 156218 443146 156454
rect 443382 156218 443414 156454
rect 442794 156134 443414 156218
rect 442794 155898 442826 156134
rect 443062 155898 443146 156134
rect 443382 155898 443414 156134
rect 442794 120454 443414 155898
rect 442794 120218 442826 120454
rect 443062 120218 443146 120454
rect 443382 120218 443414 120454
rect 442794 120134 443414 120218
rect 442794 119898 442826 120134
rect 443062 119898 443146 120134
rect 443382 119898 443414 120134
rect 442794 84454 443414 119898
rect 442794 84218 442826 84454
rect 443062 84218 443146 84454
rect 443382 84218 443414 84454
rect 442794 84134 443414 84218
rect 442794 83898 442826 84134
rect 443062 83898 443146 84134
rect 443382 83898 443414 84134
rect 442794 48454 443414 83898
rect 442794 48218 442826 48454
rect 443062 48218 443146 48454
rect 443382 48218 443414 48454
rect 442794 48134 443414 48218
rect 442794 47898 442826 48134
rect 443062 47898 443146 48134
rect 443382 47898 443414 48134
rect 442794 12454 443414 47898
rect 442794 12218 442826 12454
rect 443062 12218 443146 12454
rect 443382 12218 443414 12454
rect 442794 12134 443414 12218
rect 442794 11898 442826 12134
rect 443062 11898 443146 12134
rect 443382 11898 443414 12134
rect 442794 -2266 443414 11898
rect 442794 -2502 442826 -2266
rect 443062 -2502 443146 -2266
rect 443382 -2502 443414 -2266
rect 442794 -2586 443414 -2502
rect 442794 -2822 442826 -2586
rect 443062 -2822 443146 -2586
rect 443382 -2822 443414 -2586
rect 442794 -7654 443414 -2822
rect 447294 707718 447914 711590
rect 447294 707482 447326 707718
rect 447562 707482 447646 707718
rect 447882 707482 447914 707718
rect 447294 707398 447914 707482
rect 447294 707162 447326 707398
rect 447562 707162 447646 707398
rect 447882 707162 447914 707398
rect 447294 700954 447914 707162
rect 447294 700718 447326 700954
rect 447562 700718 447646 700954
rect 447882 700718 447914 700954
rect 447294 700634 447914 700718
rect 447294 700398 447326 700634
rect 447562 700398 447646 700634
rect 447882 700398 447914 700634
rect 447294 664954 447914 700398
rect 447294 664718 447326 664954
rect 447562 664718 447646 664954
rect 447882 664718 447914 664954
rect 447294 664634 447914 664718
rect 447294 664398 447326 664634
rect 447562 664398 447646 664634
rect 447882 664398 447914 664634
rect 447294 628954 447914 664398
rect 447294 628718 447326 628954
rect 447562 628718 447646 628954
rect 447882 628718 447914 628954
rect 447294 628634 447914 628718
rect 447294 628398 447326 628634
rect 447562 628398 447646 628634
rect 447882 628398 447914 628634
rect 447294 592954 447914 628398
rect 447294 592718 447326 592954
rect 447562 592718 447646 592954
rect 447882 592718 447914 592954
rect 447294 592634 447914 592718
rect 447294 592398 447326 592634
rect 447562 592398 447646 592634
rect 447882 592398 447914 592634
rect 447294 556954 447914 592398
rect 447294 556718 447326 556954
rect 447562 556718 447646 556954
rect 447882 556718 447914 556954
rect 447294 556634 447914 556718
rect 447294 556398 447326 556634
rect 447562 556398 447646 556634
rect 447882 556398 447914 556634
rect 447294 520954 447914 556398
rect 447294 520718 447326 520954
rect 447562 520718 447646 520954
rect 447882 520718 447914 520954
rect 447294 520634 447914 520718
rect 447294 520398 447326 520634
rect 447562 520398 447646 520634
rect 447882 520398 447914 520634
rect 447294 484954 447914 520398
rect 447294 484718 447326 484954
rect 447562 484718 447646 484954
rect 447882 484718 447914 484954
rect 447294 484634 447914 484718
rect 447294 484398 447326 484634
rect 447562 484398 447646 484634
rect 447882 484398 447914 484634
rect 447294 448954 447914 484398
rect 447294 448718 447326 448954
rect 447562 448718 447646 448954
rect 447882 448718 447914 448954
rect 447294 448634 447914 448718
rect 447294 448398 447326 448634
rect 447562 448398 447646 448634
rect 447882 448398 447914 448634
rect 447294 412954 447914 448398
rect 447294 412718 447326 412954
rect 447562 412718 447646 412954
rect 447882 412718 447914 412954
rect 447294 412634 447914 412718
rect 447294 412398 447326 412634
rect 447562 412398 447646 412634
rect 447882 412398 447914 412634
rect 447294 376954 447914 412398
rect 447294 376718 447326 376954
rect 447562 376718 447646 376954
rect 447882 376718 447914 376954
rect 447294 376634 447914 376718
rect 447294 376398 447326 376634
rect 447562 376398 447646 376634
rect 447882 376398 447914 376634
rect 447294 340954 447914 376398
rect 447294 340718 447326 340954
rect 447562 340718 447646 340954
rect 447882 340718 447914 340954
rect 447294 340634 447914 340718
rect 447294 340398 447326 340634
rect 447562 340398 447646 340634
rect 447882 340398 447914 340634
rect 447294 304954 447914 340398
rect 447294 304718 447326 304954
rect 447562 304718 447646 304954
rect 447882 304718 447914 304954
rect 447294 304634 447914 304718
rect 447294 304398 447326 304634
rect 447562 304398 447646 304634
rect 447882 304398 447914 304634
rect 447294 268954 447914 304398
rect 447294 268718 447326 268954
rect 447562 268718 447646 268954
rect 447882 268718 447914 268954
rect 447294 268634 447914 268718
rect 447294 268398 447326 268634
rect 447562 268398 447646 268634
rect 447882 268398 447914 268634
rect 447294 232954 447914 268398
rect 447294 232718 447326 232954
rect 447562 232718 447646 232954
rect 447882 232718 447914 232954
rect 447294 232634 447914 232718
rect 447294 232398 447326 232634
rect 447562 232398 447646 232634
rect 447882 232398 447914 232634
rect 447294 196954 447914 232398
rect 447294 196718 447326 196954
rect 447562 196718 447646 196954
rect 447882 196718 447914 196954
rect 447294 196634 447914 196718
rect 447294 196398 447326 196634
rect 447562 196398 447646 196634
rect 447882 196398 447914 196634
rect 447294 160954 447914 196398
rect 447294 160718 447326 160954
rect 447562 160718 447646 160954
rect 447882 160718 447914 160954
rect 447294 160634 447914 160718
rect 447294 160398 447326 160634
rect 447562 160398 447646 160634
rect 447882 160398 447914 160634
rect 447294 124954 447914 160398
rect 447294 124718 447326 124954
rect 447562 124718 447646 124954
rect 447882 124718 447914 124954
rect 447294 124634 447914 124718
rect 447294 124398 447326 124634
rect 447562 124398 447646 124634
rect 447882 124398 447914 124634
rect 447294 88954 447914 124398
rect 447294 88718 447326 88954
rect 447562 88718 447646 88954
rect 447882 88718 447914 88954
rect 447294 88634 447914 88718
rect 447294 88398 447326 88634
rect 447562 88398 447646 88634
rect 447882 88398 447914 88634
rect 447294 52954 447914 88398
rect 447294 52718 447326 52954
rect 447562 52718 447646 52954
rect 447882 52718 447914 52954
rect 447294 52634 447914 52718
rect 447294 52398 447326 52634
rect 447562 52398 447646 52634
rect 447882 52398 447914 52634
rect 447294 16954 447914 52398
rect 447294 16718 447326 16954
rect 447562 16718 447646 16954
rect 447882 16718 447914 16954
rect 447294 16634 447914 16718
rect 447294 16398 447326 16634
rect 447562 16398 447646 16634
rect 447882 16398 447914 16634
rect 447294 -3226 447914 16398
rect 447294 -3462 447326 -3226
rect 447562 -3462 447646 -3226
rect 447882 -3462 447914 -3226
rect 447294 -3546 447914 -3462
rect 447294 -3782 447326 -3546
rect 447562 -3782 447646 -3546
rect 447882 -3782 447914 -3546
rect 447294 -7654 447914 -3782
rect 451794 708678 452414 711590
rect 451794 708442 451826 708678
rect 452062 708442 452146 708678
rect 452382 708442 452414 708678
rect 451794 708358 452414 708442
rect 451794 708122 451826 708358
rect 452062 708122 452146 708358
rect 452382 708122 452414 708358
rect 451794 669454 452414 708122
rect 451794 669218 451826 669454
rect 452062 669218 452146 669454
rect 452382 669218 452414 669454
rect 451794 669134 452414 669218
rect 451794 668898 451826 669134
rect 452062 668898 452146 669134
rect 452382 668898 452414 669134
rect 451794 633454 452414 668898
rect 451794 633218 451826 633454
rect 452062 633218 452146 633454
rect 452382 633218 452414 633454
rect 451794 633134 452414 633218
rect 451794 632898 451826 633134
rect 452062 632898 452146 633134
rect 452382 632898 452414 633134
rect 451794 597454 452414 632898
rect 451794 597218 451826 597454
rect 452062 597218 452146 597454
rect 452382 597218 452414 597454
rect 451794 597134 452414 597218
rect 451794 596898 451826 597134
rect 452062 596898 452146 597134
rect 452382 596898 452414 597134
rect 451794 561454 452414 596898
rect 451794 561218 451826 561454
rect 452062 561218 452146 561454
rect 452382 561218 452414 561454
rect 451794 561134 452414 561218
rect 451794 560898 451826 561134
rect 452062 560898 452146 561134
rect 452382 560898 452414 561134
rect 451794 525454 452414 560898
rect 451794 525218 451826 525454
rect 452062 525218 452146 525454
rect 452382 525218 452414 525454
rect 451794 525134 452414 525218
rect 451794 524898 451826 525134
rect 452062 524898 452146 525134
rect 452382 524898 452414 525134
rect 451794 489454 452414 524898
rect 451794 489218 451826 489454
rect 452062 489218 452146 489454
rect 452382 489218 452414 489454
rect 451794 489134 452414 489218
rect 451794 488898 451826 489134
rect 452062 488898 452146 489134
rect 452382 488898 452414 489134
rect 451794 453454 452414 488898
rect 451794 453218 451826 453454
rect 452062 453218 452146 453454
rect 452382 453218 452414 453454
rect 451794 453134 452414 453218
rect 451794 452898 451826 453134
rect 452062 452898 452146 453134
rect 452382 452898 452414 453134
rect 451794 417454 452414 452898
rect 451794 417218 451826 417454
rect 452062 417218 452146 417454
rect 452382 417218 452414 417454
rect 451794 417134 452414 417218
rect 451794 416898 451826 417134
rect 452062 416898 452146 417134
rect 452382 416898 452414 417134
rect 451794 381454 452414 416898
rect 451794 381218 451826 381454
rect 452062 381218 452146 381454
rect 452382 381218 452414 381454
rect 451794 381134 452414 381218
rect 451794 380898 451826 381134
rect 452062 380898 452146 381134
rect 452382 380898 452414 381134
rect 451794 345454 452414 380898
rect 451794 345218 451826 345454
rect 452062 345218 452146 345454
rect 452382 345218 452414 345454
rect 451794 345134 452414 345218
rect 451794 344898 451826 345134
rect 452062 344898 452146 345134
rect 452382 344898 452414 345134
rect 451794 309454 452414 344898
rect 451794 309218 451826 309454
rect 452062 309218 452146 309454
rect 452382 309218 452414 309454
rect 451794 309134 452414 309218
rect 451794 308898 451826 309134
rect 452062 308898 452146 309134
rect 452382 308898 452414 309134
rect 451794 273454 452414 308898
rect 451794 273218 451826 273454
rect 452062 273218 452146 273454
rect 452382 273218 452414 273454
rect 451794 273134 452414 273218
rect 451794 272898 451826 273134
rect 452062 272898 452146 273134
rect 452382 272898 452414 273134
rect 451794 237454 452414 272898
rect 451794 237218 451826 237454
rect 452062 237218 452146 237454
rect 452382 237218 452414 237454
rect 451794 237134 452414 237218
rect 451794 236898 451826 237134
rect 452062 236898 452146 237134
rect 452382 236898 452414 237134
rect 451794 201454 452414 236898
rect 451794 201218 451826 201454
rect 452062 201218 452146 201454
rect 452382 201218 452414 201454
rect 451794 201134 452414 201218
rect 451794 200898 451826 201134
rect 452062 200898 452146 201134
rect 452382 200898 452414 201134
rect 451794 165454 452414 200898
rect 451794 165218 451826 165454
rect 452062 165218 452146 165454
rect 452382 165218 452414 165454
rect 451794 165134 452414 165218
rect 451794 164898 451826 165134
rect 452062 164898 452146 165134
rect 452382 164898 452414 165134
rect 451794 129454 452414 164898
rect 451794 129218 451826 129454
rect 452062 129218 452146 129454
rect 452382 129218 452414 129454
rect 451794 129134 452414 129218
rect 451794 128898 451826 129134
rect 452062 128898 452146 129134
rect 452382 128898 452414 129134
rect 451794 93454 452414 128898
rect 451794 93218 451826 93454
rect 452062 93218 452146 93454
rect 452382 93218 452414 93454
rect 451794 93134 452414 93218
rect 451794 92898 451826 93134
rect 452062 92898 452146 93134
rect 452382 92898 452414 93134
rect 451794 57454 452414 92898
rect 451794 57218 451826 57454
rect 452062 57218 452146 57454
rect 452382 57218 452414 57454
rect 451794 57134 452414 57218
rect 451794 56898 451826 57134
rect 452062 56898 452146 57134
rect 452382 56898 452414 57134
rect 451794 21454 452414 56898
rect 451794 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 452414 21454
rect 451794 21134 452414 21218
rect 451794 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 452414 21134
rect 451794 -4186 452414 20898
rect 451794 -4422 451826 -4186
rect 452062 -4422 452146 -4186
rect 452382 -4422 452414 -4186
rect 451794 -4506 452414 -4422
rect 451794 -4742 451826 -4506
rect 452062 -4742 452146 -4506
rect 452382 -4742 452414 -4506
rect 451794 -7654 452414 -4742
rect 456294 709638 456914 711590
rect 456294 709402 456326 709638
rect 456562 709402 456646 709638
rect 456882 709402 456914 709638
rect 456294 709318 456914 709402
rect 456294 709082 456326 709318
rect 456562 709082 456646 709318
rect 456882 709082 456914 709318
rect 456294 673954 456914 709082
rect 456294 673718 456326 673954
rect 456562 673718 456646 673954
rect 456882 673718 456914 673954
rect 456294 673634 456914 673718
rect 456294 673398 456326 673634
rect 456562 673398 456646 673634
rect 456882 673398 456914 673634
rect 456294 637954 456914 673398
rect 456294 637718 456326 637954
rect 456562 637718 456646 637954
rect 456882 637718 456914 637954
rect 456294 637634 456914 637718
rect 456294 637398 456326 637634
rect 456562 637398 456646 637634
rect 456882 637398 456914 637634
rect 456294 601954 456914 637398
rect 456294 601718 456326 601954
rect 456562 601718 456646 601954
rect 456882 601718 456914 601954
rect 456294 601634 456914 601718
rect 456294 601398 456326 601634
rect 456562 601398 456646 601634
rect 456882 601398 456914 601634
rect 456294 565954 456914 601398
rect 456294 565718 456326 565954
rect 456562 565718 456646 565954
rect 456882 565718 456914 565954
rect 456294 565634 456914 565718
rect 456294 565398 456326 565634
rect 456562 565398 456646 565634
rect 456882 565398 456914 565634
rect 456294 529954 456914 565398
rect 456294 529718 456326 529954
rect 456562 529718 456646 529954
rect 456882 529718 456914 529954
rect 456294 529634 456914 529718
rect 456294 529398 456326 529634
rect 456562 529398 456646 529634
rect 456882 529398 456914 529634
rect 456294 493954 456914 529398
rect 456294 493718 456326 493954
rect 456562 493718 456646 493954
rect 456882 493718 456914 493954
rect 456294 493634 456914 493718
rect 456294 493398 456326 493634
rect 456562 493398 456646 493634
rect 456882 493398 456914 493634
rect 456294 457954 456914 493398
rect 456294 457718 456326 457954
rect 456562 457718 456646 457954
rect 456882 457718 456914 457954
rect 456294 457634 456914 457718
rect 456294 457398 456326 457634
rect 456562 457398 456646 457634
rect 456882 457398 456914 457634
rect 456294 421954 456914 457398
rect 456294 421718 456326 421954
rect 456562 421718 456646 421954
rect 456882 421718 456914 421954
rect 456294 421634 456914 421718
rect 456294 421398 456326 421634
rect 456562 421398 456646 421634
rect 456882 421398 456914 421634
rect 456294 385954 456914 421398
rect 456294 385718 456326 385954
rect 456562 385718 456646 385954
rect 456882 385718 456914 385954
rect 456294 385634 456914 385718
rect 456294 385398 456326 385634
rect 456562 385398 456646 385634
rect 456882 385398 456914 385634
rect 456294 349954 456914 385398
rect 456294 349718 456326 349954
rect 456562 349718 456646 349954
rect 456882 349718 456914 349954
rect 456294 349634 456914 349718
rect 456294 349398 456326 349634
rect 456562 349398 456646 349634
rect 456882 349398 456914 349634
rect 456294 313954 456914 349398
rect 456294 313718 456326 313954
rect 456562 313718 456646 313954
rect 456882 313718 456914 313954
rect 456294 313634 456914 313718
rect 456294 313398 456326 313634
rect 456562 313398 456646 313634
rect 456882 313398 456914 313634
rect 456294 277954 456914 313398
rect 456294 277718 456326 277954
rect 456562 277718 456646 277954
rect 456882 277718 456914 277954
rect 456294 277634 456914 277718
rect 456294 277398 456326 277634
rect 456562 277398 456646 277634
rect 456882 277398 456914 277634
rect 456294 241954 456914 277398
rect 456294 241718 456326 241954
rect 456562 241718 456646 241954
rect 456882 241718 456914 241954
rect 456294 241634 456914 241718
rect 456294 241398 456326 241634
rect 456562 241398 456646 241634
rect 456882 241398 456914 241634
rect 456294 205954 456914 241398
rect 456294 205718 456326 205954
rect 456562 205718 456646 205954
rect 456882 205718 456914 205954
rect 456294 205634 456914 205718
rect 456294 205398 456326 205634
rect 456562 205398 456646 205634
rect 456882 205398 456914 205634
rect 456294 169954 456914 205398
rect 456294 169718 456326 169954
rect 456562 169718 456646 169954
rect 456882 169718 456914 169954
rect 456294 169634 456914 169718
rect 456294 169398 456326 169634
rect 456562 169398 456646 169634
rect 456882 169398 456914 169634
rect 456294 133954 456914 169398
rect 456294 133718 456326 133954
rect 456562 133718 456646 133954
rect 456882 133718 456914 133954
rect 456294 133634 456914 133718
rect 456294 133398 456326 133634
rect 456562 133398 456646 133634
rect 456882 133398 456914 133634
rect 456294 97954 456914 133398
rect 456294 97718 456326 97954
rect 456562 97718 456646 97954
rect 456882 97718 456914 97954
rect 456294 97634 456914 97718
rect 456294 97398 456326 97634
rect 456562 97398 456646 97634
rect 456882 97398 456914 97634
rect 456294 61954 456914 97398
rect 456294 61718 456326 61954
rect 456562 61718 456646 61954
rect 456882 61718 456914 61954
rect 456294 61634 456914 61718
rect 456294 61398 456326 61634
rect 456562 61398 456646 61634
rect 456882 61398 456914 61634
rect 456294 25954 456914 61398
rect 456294 25718 456326 25954
rect 456562 25718 456646 25954
rect 456882 25718 456914 25954
rect 456294 25634 456914 25718
rect 456294 25398 456326 25634
rect 456562 25398 456646 25634
rect 456882 25398 456914 25634
rect 456294 -5146 456914 25398
rect 456294 -5382 456326 -5146
rect 456562 -5382 456646 -5146
rect 456882 -5382 456914 -5146
rect 456294 -5466 456914 -5382
rect 456294 -5702 456326 -5466
rect 456562 -5702 456646 -5466
rect 456882 -5702 456914 -5466
rect 456294 -7654 456914 -5702
rect 460794 710598 461414 711590
rect 460794 710362 460826 710598
rect 461062 710362 461146 710598
rect 461382 710362 461414 710598
rect 460794 710278 461414 710362
rect 460794 710042 460826 710278
rect 461062 710042 461146 710278
rect 461382 710042 461414 710278
rect 460794 678454 461414 710042
rect 460794 678218 460826 678454
rect 461062 678218 461146 678454
rect 461382 678218 461414 678454
rect 460794 678134 461414 678218
rect 460794 677898 460826 678134
rect 461062 677898 461146 678134
rect 461382 677898 461414 678134
rect 460794 642454 461414 677898
rect 460794 642218 460826 642454
rect 461062 642218 461146 642454
rect 461382 642218 461414 642454
rect 460794 642134 461414 642218
rect 460794 641898 460826 642134
rect 461062 641898 461146 642134
rect 461382 641898 461414 642134
rect 460794 606454 461414 641898
rect 460794 606218 460826 606454
rect 461062 606218 461146 606454
rect 461382 606218 461414 606454
rect 460794 606134 461414 606218
rect 460794 605898 460826 606134
rect 461062 605898 461146 606134
rect 461382 605898 461414 606134
rect 460794 570454 461414 605898
rect 460794 570218 460826 570454
rect 461062 570218 461146 570454
rect 461382 570218 461414 570454
rect 460794 570134 461414 570218
rect 460794 569898 460826 570134
rect 461062 569898 461146 570134
rect 461382 569898 461414 570134
rect 460794 534454 461414 569898
rect 460794 534218 460826 534454
rect 461062 534218 461146 534454
rect 461382 534218 461414 534454
rect 460794 534134 461414 534218
rect 460794 533898 460826 534134
rect 461062 533898 461146 534134
rect 461382 533898 461414 534134
rect 460794 498454 461414 533898
rect 460794 498218 460826 498454
rect 461062 498218 461146 498454
rect 461382 498218 461414 498454
rect 460794 498134 461414 498218
rect 460794 497898 460826 498134
rect 461062 497898 461146 498134
rect 461382 497898 461414 498134
rect 460794 462454 461414 497898
rect 460794 462218 460826 462454
rect 461062 462218 461146 462454
rect 461382 462218 461414 462454
rect 460794 462134 461414 462218
rect 460794 461898 460826 462134
rect 461062 461898 461146 462134
rect 461382 461898 461414 462134
rect 460794 426454 461414 461898
rect 460794 426218 460826 426454
rect 461062 426218 461146 426454
rect 461382 426218 461414 426454
rect 460794 426134 461414 426218
rect 460794 425898 460826 426134
rect 461062 425898 461146 426134
rect 461382 425898 461414 426134
rect 460794 390454 461414 425898
rect 460794 390218 460826 390454
rect 461062 390218 461146 390454
rect 461382 390218 461414 390454
rect 460794 390134 461414 390218
rect 460794 389898 460826 390134
rect 461062 389898 461146 390134
rect 461382 389898 461414 390134
rect 460794 354454 461414 389898
rect 460794 354218 460826 354454
rect 461062 354218 461146 354454
rect 461382 354218 461414 354454
rect 460794 354134 461414 354218
rect 460794 353898 460826 354134
rect 461062 353898 461146 354134
rect 461382 353898 461414 354134
rect 460794 318454 461414 353898
rect 460794 318218 460826 318454
rect 461062 318218 461146 318454
rect 461382 318218 461414 318454
rect 460794 318134 461414 318218
rect 460794 317898 460826 318134
rect 461062 317898 461146 318134
rect 461382 317898 461414 318134
rect 460794 282454 461414 317898
rect 460794 282218 460826 282454
rect 461062 282218 461146 282454
rect 461382 282218 461414 282454
rect 460794 282134 461414 282218
rect 460794 281898 460826 282134
rect 461062 281898 461146 282134
rect 461382 281898 461414 282134
rect 460794 246454 461414 281898
rect 460794 246218 460826 246454
rect 461062 246218 461146 246454
rect 461382 246218 461414 246454
rect 460794 246134 461414 246218
rect 460794 245898 460826 246134
rect 461062 245898 461146 246134
rect 461382 245898 461414 246134
rect 460794 210454 461414 245898
rect 460794 210218 460826 210454
rect 461062 210218 461146 210454
rect 461382 210218 461414 210454
rect 460794 210134 461414 210218
rect 460794 209898 460826 210134
rect 461062 209898 461146 210134
rect 461382 209898 461414 210134
rect 460794 174454 461414 209898
rect 460794 174218 460826 174454
rect 461062 174218 461146 174454
rect 461382 174218 461414 174454
rect 460794 174134 461414 174218
rect 460794 173898 460826 174134
rect 461062 173898 461146 174134
rect 461382 173898 461414 174134
rect 460794 138454 461414 173898
rect 460794 138218 460826 138454
rect 461062 138218 461146 138454
rect 461382 138218 461414 138454
rect 460794 138134 461414 138218
rect 460794 137898 460826 138134
rect 461062 137898 461146 138134
rect 461382 137898 461414 138134
rect 460794 102454 461414 137898
rect 460794 102218 460826 102454
rect 461062 102218 461146 102454
rect 461382 102218 461414 102454
rect 460794 102134 461414 102218
rect 460794 101898 460826 102134
rect 461062 101898 461146 102134
rect 461382 101898 461414 102134
rect 460794 66454 461414 101898
rect 460794 66218 460826 66454
rect 461062 66218 461146 66454
rect 461382 66218 461414 66454
rect 460794 66134 461414 66218
rect 460794 65898 460826 66134
rect 461062 65898 461146 66134
rect 461382 65898 461414 66134
rect 460794 30454 461414 65898
rect 460794 30218 460826 30454
rect 461062 30218 461146 30454
rect 461382 30218 461414 30454
rect 460794 30134 461414 30218
rect 460794 29898 460826 30134
rect 461062 29898 461146 30134
rect 461382 29898 461414 30134
rect 460794 -6106 461414 29898
rect 460794 -6342 460826 -6106
rect 461062 -6342 461146 -6106
rect 461382 -6342 461414 -6106
rect 460794 -6426 461414 -6342
rect 460794 -6662 460826 -6426
rect 461062 -6662 461146 -6426
rect 461382 -6662 461414 -6426
rect 460794 -7654 461414 -6662
rect 465294 711558 465914 711590
rect 465294 711322 465326 711558
rect 465562 711322 465646 711558
rect 465882 711322 465914 711558
rect 465294 711238 465914 711322
rect 465294 711002 465326 711238
rect 465562 711002 465646 711238
rect 465882 711002 465914 711238
rect 465294 682954 465914 711002
rect 465294 682718 465326 682954
rect 465562 682718 465646 682954
rect 465882 682718 465914 682954
rect 465294 682634 465914 682718
rect 465294 682398 465326 682634
rect 465562 682398 465646 682634
rect 465882 682398 465914 682634
rect 465294 646954 465914 682398
rect 465294 646718 465326 646954
rect 465562 646718 465646 646954
rect 465882 646718 465914 646954
rect 465294 646634 465914 646718
rect 465294 646398 465326 646634
rect 465562 646398 465646 646634
rect 465882 646398 465914 646634
rect 465294 610954 465914 646398
rect 465294 610718 465326 610954
rect 465562 610718 465646 610954
rect 465882 610718 465914 610954
rect 465294 610634 465914 610718
rect 465294 610398 465326 610634
rect 465562 610398 465646 610634
rect 465882 610398 465914 610634
rect 465294 574954 465914 610398
rect 465294 574718 465326 574954
rect 465562 574718 465646 574954
rect 465882 574718 465914 574954
rect 465294 574634 465914 574718
rect 465294 574398 465326 574634
rect 465562 574398 465646 574634
rect 465882 574398 465914 574634
rect 465294 538954 465914 574398
rect 465294 538718 465326 538954
rect 465562 538718 465646 538954
rect 465882 538718 465914 538954
rect 465294 538634 465914 538718
rect 465294 538398 465326 538634
rect 465562 538398 465646 538634
rect 465882 538398 465914 538634
rect 465294 502954 465914 538398
rect 465294 502718 465326 502954
rect 465562 502718 465646 502954
rect 465882 502718 465914 502954
rect 465294 502634 465914 502718
rect 465294 502398 465326 502634
rect 465562 502398 465646 502634
rect 465882 502398 465914 502634
rect 465294 466954 465914 502398
rect 465294 466718 465326 466954
rect 465562 466718 465646 466954
rect 465882 466718 465914 466954
rect 465294 466634 465914 466718
rect 465294 466398 465326 466634
rect 465562 466398 465646 466634
rect 465882 466398 465914 466634
rect 465294 430954 465914 466398
rect 465294 430718 465326 430954
rect 465562 430718 465646 430954
rect 465882 430718 465914 430954
rect 465294 430634 465914 430718
rect 465294 430398 465326 430634
rect 465562 430398 465646 430634
rect 465882 430398 465914 430634
rect 465294 394954 465914 430398
rect 465294 394718 465326 394954
rect 465562 394718 465646 394954
rect 465882 394718 465914 394954
rect 465294 394634 465914 394718
rect 465294 394398 465326 394634
rect 465562 394398 465646 394634
rect 465882 394398 465914 394634
rect 465294 358954 465914 394398
rect 465294 358718 465326 358954
rect 465562 358718 465646 358954
rect 465882 358718 465914 358954
rect 465294 358634 465914 358718
rect 465294 358398 465326 358634
rect 465562 358398 465646 358634
rect 465882 358398 465914 358634
rect 465294 322954 465914 358398
rect 465294 322718 465326 322954
rect 465562 322718 465646 322954
rect 465882 322718 465914 322954
rect 465294 322634 465914 322718
rect 465294 322398 465326 322634
rect 465562 322398 465646 322634
rect 465882 322398 465914 322634
rect 465294 286954 465914 322398
rect 465294 286718 465326 286954
rect 465562 286718 465646 286954
rect 465882 286718 465914 286954
rect 465294 286634 465914 286718
rect 465294 286398 465326 286634
rect 465562 286398 465646 286634
rect 465882 286398 465914 286634
rect 465294 250954 465914 286398
rect 465294 250718 465326 250954
rect 465562 250718 465646 250954
rect 465882 250718 465914 250954
rect 465294 250634 465914 250718
rect 465294 250398 465326 250634
rect 465562 250398 465646 250634
rect 465882 250398 465914 250634
rect 465294 214954 465914 250398
rect 465294 214718 465326 214954
rect 465562 214718 465646 214954
rect 465882 214718 465914 214954
rect 465294 214634 465914 214718
rect 465294 214398 465326 214634
rect 465562 214398 465646 214634
rect 465882 214398 465914 214634
rect 465294 178954 465914 214398
rect 465294 178718 465326 178954
rect 465562 178718 465646 178954
rect 465882 178718 465914 178954
rect 465294 178634 465914 178718
rect 465294 178398 465326 178634
rect 465562 178398 465646 178634
rect 465882 178398 465914 178634
rect 465294 142954 465914 178398
rect 465294 142718 465326 142954
rect 465562 142718 465646 142954
rect 465882 142718 465914 142954
rect 465294 142634 465914 142718
rect 465294 142398 465326 142634
rect 465562 142398 465646 142634
rect 465882 142398 465914 142634
rect 465294 106954 465914 142398
rect 465294 106718 465326 106954
rect 465562 106718 465646 106954
rect 465882 106718 465914 106954
rect 465294 106634 465914 106718
rect 465294 106398 465326 106634
rect 465562 106398 465646 106634
rect 465882 106398 465914 106634
rect 465294 70954 465914 106398
rect 465294 70718 465326 70954
rect 465562 70718 465646 70954
rect 465882 70718 465914 70954
rect 465294 70634 465914 70718
rect 465294 70398 465326 70634
rect 465562 70398 465646 70634
rect 465882 70398 465914 70634
rect 465294 34954 465914 70398
rect 465294 34718 465326 34954
rect 465562 34718 465646 34954
rect 465882 34718 465914 34954
rect 465294 34634 465914 34718
rect 465294 34398 465326 34634
rect 465562 34398 465646 34634
rect 465882 34398 465914 34634
rect 465294 -7066 465914 34398
rect 465294 -7302 465326 -7066
rect 465562 -7302 465646 -7066
rect 465882 -7302 465914 -7066
rect 465294 -7386 465914 -7302
rect 465294 -7622 465326 -7386
rect 465562 -7622 465646 -7386
rect 465882 -7622 465914 -7386
rect 465294 -7654 465914 -7622
rect 469794 704838 470414 711590
rect 469794 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 470414 704838
rect 469794 704518 470414 704602
rect 469794 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 470414 704518
rect 469794 687454 470414 704282
rect 469794 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 470414 687454
rect 469794 687134 470414 687218
rect 469794 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 470414 687134
rect 469794 651454 470414 686898
rect 469794 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 470414 651454
rect 469794 651134 470414 651218
rect 469794 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 470414 651134
rect 469794 615454 470414 650898
rect 469794 615218 469826 615454
rect 470062 615218 470146 615454
rect 470382 615218 470414 615454
rect 469794 615134 470414 615218
rect 469794 614898 469826 615134
rect 470062 614898 470146 615134
rect 470382 614898 470414 615134
rect 469794 579454 470414 614898
rect 469794 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 470414 579454
rect 469794 579134 470414 579218
rect 469794 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 470414 579134
rect 469794 543454 470414 578898
rect 469794 543218 469826 543454
rect 470062 543218 470146 543454
rect 470382 543218 470414 543454
rect 469794 543134 470414 543218
rect 469794 542898 469826 543134
rect 470062 542898 470146 543134
rect 470382 542898 470414 543134
rect 469794 507454 470414 542898
rect 469794 507218 469826 507454
rect 470062 507218 470146 507454
rect 470382 507218 470414 507454
rect 469794 507134 470414 507218
rect 469794 506898 469826 507134
rect 470062 506898 470146 507134
rect 470382 506898 470414 507134
rect 469794 471454 470414 506898
rect 469794 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 470414 471454
rect 469794 471134 470414 471218
rect 469794 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 470414 471134
rect 469794 435454 470414 470898
rect 469794 435218 469826 435454
rect 470062 435218 470146 435454
rect 470382 435218 470414 435454
rect 469794 435134 470414 435218
rect 469794 434898 469826 435134
rect 470062 434898 470146 435134
rect 470382 434898 470414 435134
rect 469794 399454 470414 434898
rect 469794 399218 469826 399454
rect 470062 399218 470146 399454
rect 470382 399218 470414 399454
rect 469794 399134 470414 399218
rect 469794 398898 469826 399134
rect 470062 398898 470146 399134
rect 470382 398898 470414 399134
rect 469794 363454 470414 398898
rect 469794 363218 469826 363454
rect 470062 363218 470146 363454
rect 470382 363218 470414 363454
rect 469794 363134 470414 363218
rect 469794 362898 469826 363134
rect 470062 362898 470146 363134
rect 470382 362898 470414 363134
rect 469794 327454 470414 362898
rect 469794 327218 469826 327454
rect 470062 327218 470146 327454
rect 470382 327218 470414 327454
rect 469794 327134 470414 327218
rect 469794 326898 469826 327134
rect 470062 326898 470146 327134
rect 470382 326898 470414 327134
rect 469794 291454 470414 326898
rect 469794 291218 469826 291454
rect 470062 291218 470146 291454
rect 470382 291218 470414 291454
rect 469794 291134 470414 291218
rect 469794 290898 469826 291134
rect 470062 290898 470146 291134
rect 470382 290898 470414 291134
rect 469794 255454 470414 290898
rect 469794 255218 469826 255454
rect 470062 255218 470146 255454
rect 470382 255218 470414 255454
rect 469794 255134 470414 255218
rect 469794 254898 469826 255134
rect 470062 254898 470146 255134
rect 470382 254898 470414 255134
rect 469794 219454 470414 254898
rect 469794 219218 469826 219454
rect 470062 219218 470146 219454
rect 470382 219218 470414 219454
rect 469794 219134 470414 219218
rect 469794 218898 469826 219134
rect 470062 218898 470146 219134
rect 470382 218898 470414 219134
rect 469794 183454 470414 218898
rect 469794 183218 469826 183454
rect 470062 183218 470146 183454
rect 470382 183218 470414 183454
rect 469794 183134 470414 183218
rect 469794 182898 469826 183134
rect 470062 182898 470146 183134
rect 470382 182898 470414 183134
rect 469794 147454 470414 182898
rect 469794 147218 469826 147454
rect 470062 147218 470146 147454
rect 470382 147218 470414 147454
rect 469794 147134 470414 147218
rect 469794 146898 469826 147134
rect 470062 146898 470146 147134
rect 470382 146898 470414 147134
rect 469794 111454 470414 146898
rect 469794 111218 469826 111454
rect 470062 111218 470146 111454
rect 470382 111218 470414 111454
rect 469794 111134 470414 111218
rect 469794 110898 469826 111134
rect 470062 110898 470146 111134
rect 470382 110898 470414 111134
rect 469794 75454 470414 110898
rect 469794 75218 469826 75454
rect 470062 75218 470146 75454
rect 470382 75218 470414 75454
rect 469794 75134 470414 75218
rect 469794 74898 469826 75134
rect 470062 74898 470146 75134
rect 470382 74898 470414 75134
rect 469794 39454 470414 74898
rect 469794 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 470414 39454
rect 469794 39134 470414 39218
rect 469794 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 470414 39134
rect 469794 3454 470414 38898
rect 469794 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 470414 3454
rect 469794 3134 470414 3218
rect 469794 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 470414 3134
rect 469794 -346 470414 2898
rect 469794 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 470414 -346
rect 469794 -666 470414 -582
rect 469794 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 470414 -666
rect 469794 -7654 470414 -902
rect 474294 705798 474914 711590
rect 474294 705562 474326 705798
rect 474562 705562 474646 705798
rect 474882 705562 474914 705798
rect 474294 705478 474914 705562
rect 474294 705242 474326 705478
rect 474562 705242 474646 705478
rect 474882 705242 474914 705478
rect 474294 691954 474914 705242
rect 474294 691718 474326 691954
rect 474562 691718 474646 691954
rect 474882 691718 474914 691954
rect 474294 691634 474914 691718
rect 474294 691398 474326 691634
rect 474562 691398 474646 691634
rect 474882 691398 474914 691634
rect 474294 655954 474914 691398
rect 474294 655718 474326 655954
rect 474562 655718 474646 655954
rect 474882 655718 474914 655954
rect 474294 655634 474914 655718
rect 474294 655398 474326 655634
rect 474562 655398 474646 655634
rect 474882 655398 474914 655634
rect 474294 619954 474914 655398
rect 474294 619718 474326 619954
rect 474562 619718 474646 619954
rect 474882 619718 474914 619954
rect 474294 619634 474914 619718
rect 474294 619398 474326 619634
rect 474562 619398 474646 619634
rect 474882 619398 474914 619634
rect 474294 583954 474914 619398
rect 474294 583718 474326 583954
rect 474562 583718 474646 583954
rect 474882 583718 474914 583954
rect 474294 583634 474914 583718
rect 474294 583398 474326 583634
rect 474562 583398 474646 583634
rect 474882 583398 474914 583634
rect 474294 547954 474914 583398
rect 474294 547718 474326 547954
rect 474562 547718 474646 547954
rect 474882 547718 474914 547954
rect 474294 547634 474914 547718
rect 474294 547398 474326 547634
rect 474562 547398 474646 547634
rect 474882 547398 474914 547634
rect 474294 511954 474914 547398
rect 474294 511718 474326 511954
rect 474562 511718 474646 511954
rect 474882 511718 474914 511954
rect 474294 511634 474914 511718
rect 474294 511398 474326 511634
rect 474562 511398 474646 511634
rect 474882 511398 474914 511634
rect 474294 475954 474914 511398
rect 474294 475718 474326 475954
rect 474562 475718 474646 475954
rect 474882 475718 474914 475954
rect 474294 475634 474914 475718
rect 474294 475398 474326 475634
rect 474562 475398 474646 475634
rect 474882 475398 474914 475634
rect 474294 439954 474914 475398
rect 474294 439718 474326 439954
rect 474562 439718 474646 439954
rect 474882 439718 474914 439954
rect 474294 439634 474914 439718
rect 474294 439398 474326 439634
rect 474562 439398 474646 439634
rect 474882 439398 474914 439634
rect 474294 403954 474914 439398
rect 474294 403718 474326 403954
rect 474562 403718 474646 403954
rect 474882 403718 474914 403954
rect 474294 403634 474914 403718
rect 474294 403398 474326 403634
rect 474562 403398 474646 403634
rect 474882 403398 474914 403634
rect 474294 367954 474914 403398
rect 474294 367718 474326 367954
rect 474562 367718 474646 367954
rect 474882 367718 474914 367954
rect 474294 367634 474914 367718
rect 474294 367398 474326 367634
rect 474562 367398 474646 367634
rect 474882 367398 474914 367634
rect 474294 331954 474914 367398
rect 474294 331718 474326 331954
rect 474562 331718 474646 331954
rect 474882 331718 474914 331954
rect 474294 331634 474914 331718
rect 474294 331398 474326 331634
rect 474562 331398 474646 331634
rect 474882 331398 474914 331634
rect 474294 295954 474914 331398
rect 474294 295718 474326 295954
rect 474562 295718 474646 295954
rect 474882 295718 474914 295954
rect 474294 295634 474914 295718
rect 474294 295398 474326 295634
rect 474562 295398 474646 295634
rect 474882 295398 474914 295634
rect 474294 259954 474914 295398
rect 474294 259718 474326 259954
rect 474562 259718 474646 259954
rect 474882 259718 474914 259954
rect 474294 259634 474914 259718
rect 474294 259398 474326 259634
rect 474562 259398 474646 259634
rect 474882 259398 474914 259634
rect 474294 223954 474914 259398
rect 474294 223718 474326 223954
rect 474562 223718 474646 223954
rect 474882 223718 474914 223954
rect 474294 223634 474914 223718
rect 474294 223398 474326 223634
rect 474562 223398 474646 223634
rect 474882 223398 474914 223634
rect 474294 187954 474914 223398
rect 474294 187718 474326 187954
rect 474562 187718 474646 187954
rect 474882 187718 474914 187954
rect 474294 187634 474914 187718
rect 474294 187398 474326 187634
rect 474562 187398 474646 187634
rect 474882 187398 474914 187634
rect 474294 151954 474914 187398
rect 474294 151718 474326 151954
rect 474562 151718 474646 151954
rect 474882 151718 474914 151954
rect 474294 151634 474914 151718
rect 474294 151398 474326 151634
rect 474562 151398 474646 151634
rect 474882 151398 474914 151634
rect 474294 115954 474914 151398
rect 474294 115718 474326 115954
rect 474562 115718 474646 115954
rect 474882 115718 474914 115954
rect 474294 115634 474914 115718
rect 474294 115398 474326 115634
rect 474562 115398 474646 115634
rect 474882 115398 474914 115634
rect 474294 79954 474914 115398
rect 474294 79718 474326 79954
rect 474562 79718 474646 79954
rect 474882 79718 474914 79954
rect 474294 79634 474914 79718
rect 474294 79398 474326 79634
rect 474562 79398 474646 79634
rect 474882 79398 474914 79634
rect 474294 43954 474914 79398
rect 474294 43718 474326 43954
rect 474562 43718 474646 43954
rect 474882 43718 474914 43954
rect 474294 43634 474914 43718
rect 474294 43398 474326 43634
rect 474562 43398 474646 43634
rect 474882 43398 474914 43634
rect 474294 7954 474914 43398
rect 474294 7718 474326 7954
rect 474562 7718 474646 7954
rect 474882 7718 474914 7954
rect 474294 7634 474914 7718
rect 474294 7398 474326 7634
rect 474562 7398 474646 7634
rect 474882 7398 474914 7634
rect 474294 -1306 474914 7398
rect 474294 -1542 474326 -1306
rect 474562 -1542 474646 -1306
rect 474882 -1542 474914 -1306
rect 474294 -1626 474914 -1542
rect 474294 -1862 474326 -1626
rect 474562 -1862 474646 -1626
rect 474882 -1862 474914 -1626
rect 474294 -7654 474914 -1862
rect 478794 706758 479414 711590
rect 478794 706522 478826 706758
rect 479062 706522 479146 706758
rect 479382 706522 479414 706758
rect 478794 706438 479414 706522
rect 478794 706202 478826 706438
rect 479062 706202 479146 706438
rect 479382 706202 479414 706438
rect 478794 696454 479414 706202
rect 478794 696218 478826 696454
rect 479062 696218 479146 696454
rect 479382 696218 479414 696454
rect 478794 696134 479414 696218
rect 478794 695898 478826 696134
rect 479062 695898 479146 696134
rect 479382 695898 479414 696134
rect 478794 660454 479414 695898
rect 478794 660218 478826 660454
rect 479062 660218 479146 660454
rect 479382 660218 479414 660454
rect 478794 660134 479414 660218
rect 478794 659898 478826 660134
rect 479062 659898 479146 660134
rect 479382 659898 479414 660134
rect 478794 624454 479414 659898
rect 478794 624218 478826 624454
rect 479062 624218 479146 624454
rect 479382 624218 479414 624454
rect 478794 624134 479414 624218
rect 478794 623898 478826 624134
rect 479062 623898 479146 624134
rect 479382 623898 479414 624134
rect 478794 588454 479414 623898
rect 478794 588218 478826 588454
rect 479062 588218 479146 588454
rect 479382 588218 479414 588454
rect 478794 588134 479414 588218
rect 478794 587898 478826 588134
rect 479062 587898 479146 588134
rect 479382 587898 479414 588134
rect 478794 552454 479414 587898
rect 478794 552218 478826 552454
rect 479062 552218 479146 552454
rect 479382 552218 479414 552454
rect 478794 552134 479414 552218
rect 478794 551898 478826 552134
rect 479062 551898 479146 552134
rect 479382 551898 479414 552134
rect 478794 516454 479414 551898
rect 478794 516218 478826 516454
rect 479062 516218 479146 516454
rect 479382 516218 479414 516454
rect 478794 516134 479414 516218
rect 478794 515898 478826 516134
rect 479062 515898 479146 516134
rect 479382 515898 479414 516134
rect 478794 480454 479414 515898
rect 478794 480218 478826 480454
rect 479062 480218 479146 480454
rect 479382 480218 479414 480454
rect 478794 480134 479414 480218
rect 478794 479898 478826 480134
rect 479062 479898 479146 480134
rect 479382 479898 479414 480134
rect 478794 444454 479414 479898
rect 478794 444218 478826 444454
rect 479062 444218 479146 444454
rect 479382 444218 479414 444454
rect 478794 444134 479414 444218
rect 478794 443898 478826 444134
rect 479062 443898 479146 444134
rect 479382 443898 479414 444134
rect 478794 408454 479414 443898
rect 478794 408218 478826 408454
rect 479062 408218 479146 408454
rect 479382 408218 479414 408454
rect 478794 408134 479414 408218
rect 478794 407898 478826 408134
rect 479062 407898 479146 408134
rect 479382 407898 479414 408134
rect 478794 372454 479414 407898
rect 478794 372218 478826 372454
rect 479062 372218 479146 372454
rect 479382 372218 479414 372454
rect 478794 372134 479414 372218
rect 478794 371898 478826 372134
rect 479062 371898 479146 372134
rect 479382 371898 479414 372134
rect 478794 336454 479414 371898
rect 478794 336218 478826 336454
rect 479062 336218 479146 336454
rect 479382 336218 479414 336454
rect 478794 336134 479414 336218
rect 478794 335898 478826 336134
rect 479062 335898 479146 336134
rect 479382 335898 479414 336134
rect 478794 300454 479414 335898
rect 478794 300218 478826 300454
rect 479062 300218 479146 300454
rect 479382 300218 479414 300454
rect 478794 300134 479414 300218
rect 478794 299898 478826 300134
rect 479062 299898 479146 300134
rect 479382 299898 479414 300134
rect 478794 264454 479414 299898
rect 478794 264218 478826 264454
rect 479062 264218 479146 264454
rect 479382 264218 479414 264454
rect 478794 264134 479414 264218
rect 478794 263898 478826 264134
rect 479062 263898 479146 264134
rect 479382 263898 479414 264134
rect 478794 228454 479414 263898
rect 478794 228218 478826 228454
rect 479062 228218 479146 228454
rect 479382 228218 479414 228454
rect 478794 228134 479414 228218
rect 478794 227898 478826 228134
rect 479062 227898 479146 228134
rect 479382 227898 479414 228134
rect 478794 192454 479414 227898
rect 478794 192218 478826 192454
rect 479062 192218 479146 192454
rect 479382 192218 479414 192454
rect 478794 192134 479414 192218
rect 478794 191898 478826 192134
rect 479062 191898 479146 192134
rect 479382 191898 479414 192134
rect 478794 156454 479414 191898
rect 478794 156218 478826 156454
rect 479062 156218 479146 156454
rect 479382 156218 479414 156454
rect 478794 156134 479414 156218
rect 478794 155898 478826 156134
rect 479062 155898 479146 156134
rect 479382 155898 479414 156134
rect 478794 120454 479414 155898
rect 478794 120218 478826 120454
rect 479062 120218 479146 120454
rect 479382 120218 479414 120454
rect 478794 120134 479414 120218
rect 478794 119898 478826 120134
rect 479062 119898 479146 120134
rect 479382 119898 479414 120134
rect 478794 84454 479414 119898
rect 478794 84218 478826 84454
rect 479062 84218 479146 84454
rect 479382 84218 479414 84454
rect 478794 84134 479414 84218
rect 478794 83898 478826 84134
rect 479062 83898 479146 84134
rect 479382 83898 479414 84134
rect 478794 48454 479414 83898
rect 478794 48218 478826 48454
rect 479062 48218 479146 48454
rect 479382 48218 479414 48454
rect 478794 48134 479414 48218
rect 478794 47898 478826 48134
rect 479062 47898 479146 48134
rect 479382 47898 479414 48134
rect 478794 12454 479414 47898
rect 478794 12218 478826 12454
rect 479062 12218 479146 12454
rect 479382 12218 479414 12454
rect 478794 12134 479414 12218
rect 478794 11898 478826 12134
rect 479062 11898 479146 12134
rect 479382 11898 479414 12134
rect 478794 -2266 479414 11898
rect 478794 -2502 478826 -2266
rect 479062 -2502 479146 -2266
rect 479382 -2502 479414 -2266
rect 478794 -2586 479414 -2502
rect 478794 -2822 478826 -2586
rect 479062 -2822 479146 -2586
rect 479382 -2822 479414 -2586
rect 478794 -7654 479414 -2822
rect 483294 707718 483914 711590
rect 483294 707482 483326 707718
rect 483562 707482 483646 707718
rect 483882 707482 483914 707718
rect 483294 707398 483914 707482
rect 483294 707162 483326 707398
rect 483562 707162 483646 707398
rect 483882 707162 483914 707398
rect 483294 700954 483914 707162
rect 483294 700718 483326 700954
rect 483562 700718 483646 700954
rect 483882 700718 483914 700954
rect 483294 700634 483914 700718
rect 483294 700398 483326 700634
rect 483562 700398 483646 700634
rect 483882 700398 483914 700634
rect 483294 664954 483914 700398
rect 483294 664718 483326 664954
rect 483562 664718 483646 664954
rect 483882 664718 483914 664954
rect 483294 664634 483914 664718
rect 483294 664398 483326 664634
rect 483562 664398 483646 664634
rect 483882 664398 483914 664634
rect 483294 628954 483914 664398
rect 483294 628718 483326 628954
rect 483562 628718 483646 628954
rect 483882 628718 483914 628954
rect 483294 628634 483914 628718
rect 483294 628398 483326 628634
rect 483562 628398 483646 628634
rect 483882 628398 483914 628634
rect 483294 592954 483914 628398
rect 483294 592718 483326 592954
rect 483562 592718 483646 592954
rect 483882 592718 483914 592954
rect 483294 592634 483914 592718
rect 483294 592398 483326 592634
rect 483562 592398 483646 592634
rect 483882 592398 483914 592634
rect 483294 556954 483914 592398
rect 483294 556718 483326 556954
rect 483562 556718 483646 556954
rect 483882 556718 483914 556954
rect 483294 556634 483914 556718
rect 483294 556398 483326 556634
rect 483562 556398 483646 556634
rect 483882 556398 483914 556634
rect 483294 520954 483914 556398
rect 483294 520718 483326 520954
rect 483562 520718 483646 520954
rect 483882 520718 483914 520954
rect 483294 520634 483914 520718
rect 483294 520398 483326 520634
rect 483562 520398 483646 520634
rect 483882 520398 483914 520634
rect 483294 484954 483914 520398
rect 483294 484718 483326 484954
rect 483562 484718 483646 484954
rect 483882 484718 483914 484954
rect 483294 484634 483914 484718
rect 483294 484398 483326 484634
rect 483562 484398 483646 484634
rect 483882 484398 483914 484634
rect 483294 448954 483914 484398
rect 483294 448718 483326 448954
rect 483562 448718 483646 448954
rect 483882 448718 483914 448954
rect 483294 448634 483914 448718
rect 483294 448398 483326 448634
rect 483562 448398 483646 448634
rect 483882 448398 483914 448634
rect 483294 412954 483914 448398
rect 483294 412718 483326 412954
rect 483562 412718 483646 412954
rect 483882 412718 483914 412954
rect 483294 412634 483914 412718
rect 483294 412398 483326 412634
rect 483562 412398 483646 412634
rect 483882 412398 483914 412634
rect 483294 376954 483914 412398
rect 483294 376718 483326 376954
rect 483562 376718 483646 376954
rect 483882 376718 483914 376954
rect 483294 376634 483914 376718
rect 483294 376398 483326 376634
rect 483562 376398 483646 376634
rect 483882 376398 483914 376634
rect 483294 340954 483914 376398
rect 483294 340718 483326 340954
rect 483562 340718 483646 340954
rect 483882 340718 483914 340954
rect 483294 340634 483914 340718
rect 483294 340398 483326 340634
rect 483562 340398 483646 340634
rect 483882 340398 483914 340634
rect 483294 304954 483914 340398
rect 483294 304718 483326 304954
rect 483562 304718 483646 304954
rect 483882 304718 483914 304954
rect 483294 304634 483914 304718
rect 483294 304398 483326 304634
rect 483562 304398 483646 304634
rect 483882 304398 483914 304634
rect 483294 268954 483914 304398
rect 483294 268718 483326 268954
rect 483562 268718 483646 268954
rect 483882 268718 483914 268954
rect 483294 268634 483914 268718
rect 483294 268398 483326 268634
rect 483562 268398 483646 268634
rect 483882 268398 483914 268634
rect 483294 232954 483914 268398
rect 483294 232718 483326 232954
rect 483562 232718 483646 232954
rect 483882 232718 483914 232954
rect 483294 232634 483914 232718
rect 483294 232398 483326 232634
rect 483562 232398 483646 232634
rect 483882 232398 483914 232634
rect 483294 196954 483914 232398
rect 483294 196718 483326 196954
rect 483562 196718 483646 196954
rect 483882 196718 483914 196954
rect 483294 196634 483914 196718
rect 483294 196398 483326 196634
rect 483562 196398 483646 196634
rect 483882 196398 483914 196634
rect 483294 160954 483914 196398
rect 483294 160718 483326 160954
rect 483562 160718 483646 160954
rect 483882 160718 483914 160954
rect 483294 160634 483914 160718
rect 483294 160398 483326 160634
rect 483562 160398 483646 160634
rect 483882 160398 483914 160634
rect 483294 124954 483914 160398
rect 483294 124718 483326 124954
rect 483562 124718 483646 124954
rect 483882 124718 483914 124954
rect 483294 124634 483914 124718
rect 483294 124398 483326 124634
rect 483562 124398 483646 124634
rect 483882 124398 483914 124634
rect 483294 88954 483914 124398
rect 483294 88718 483326 88954
rect 483562 88718 483646 88954
rect 483882 88718 483914 88954
rect 483294 88634 483914 88718
rect 483294 88398 483326 88634
rect 483562 88398 483646 88634
rect 483882 88398 483914 88634
rect 483294 52954 483914 88398
rect 483294 52718 483326 52954
rect 483562 52718 483646 52954
rect 483882 52718 483914 52954
rect 483294 52634 483914 52718
rect 483294 52398 483326 52634
rect 483562 52398 483646 52634
rect 483882 52398 483914 52634
rect 483294 16954 483914 52398
rect 483294 16718 483326 16954
rect 483562 16718 483646 16954
rect 483882 16718 483914 16954
rect 483294 16634 483914 16718
rect 483294 16398 483326 16634
rect 483562 16398 483646 16634
rect 483882 16398 483914 16634
rect 483294 -3226 483914 16398
rect 483294 -3462 483326 -3226
rect 483562 -3462 483646 -3226
rect 483882 -3462 483914 -3226
rect 483294 -3546 483914 -3462
rect 483294 -3782 483326 -3546
rect 483562 -3782 483646 -3546
rect 483882 -3782 483914 -3546
rect 483294 -7654 483914 -3782
rect 487794 708678 488414 711590
rect 487794 708442 487826 708678
rect 488062 708442 488146 708678
rect 488382 708442 488414 708678
rect 487794 708358 488414 708442
rect 487794 708122 487826 708358
rect 488062 708122 488146 708358
rect 488382 708122 488414 708358
rect 487794 669454 488414 708122
rect 487794 669218 487826 669454
rect 488062 669218 488146 669454
rect 488382 669218 488414 669454
rect 487794 669134 488414 669218
rect 487794 668898 487826 669134
rect 488062 668898 488146 669134
rect 488382 668898 488414 669134
rect 487794 633454 488414 668898
rect 487794 633218 487826 633454
rect 488062 633218 488146 633454
rect 488382 633218 488414 633454
rect 487794 633134 488414 633218
rect 487794 632898 487826 633134
rect 488062 632898 488146 633134
rect 488382 632898 488414 633134
rect 487794 597454 488414 632898
rect 487794 597218 487826 597454
rect 488062 597218 488146 597454
rect 488382 597218 488414 597454
rect 487794 597134 488414 597218
rect 487794 596898 487826 597134
rect 488062 596898 488146 597134
rect 488382 596898 488414 597134
rect 487794 561454 488414 596898
rect 487794 561218 487826 561454
rect 488062 561218 488146 561454
rect 488382 561218 488414 561454
rect 487794 561134 488414 561218
rect 487794 560898 487826 561134
rect 488062 560898 488146 561134
rect 488382 560898 488414 561134
rect 487794 525454 488414 560898
rect 487794 525218 487826 525454
rect 488062 525218 488146 525454
rect 488382 525218 488414 525454
rect 487794 525134 488414 525218
rect 487794 524898 487826 525134
rect 488062 524898 488146 525134
rect 488382 524898 488414 525134
rect 487794 489454 488414 524898
rect 487794 489218 487826 489454
rect 488062 489218 488146 489454
rect 488382 489218 488414 489454
rect 487794 489134 488414 489218
rect 487794 488898 487826 489134
rect 488062 488898 488146 489134
rect 488382 488898 488414 489134
rect 487794 453454 488414 488898
rect 487794 453218 487826 453454
rect 488062 453218 488146 453454
rect 488382 453218 488414 453454
rect 487794 453134 488414 453218
rect 487794 452898 487826 453134
rect 488062 452898 488146 453134
rect 488382 452898 488414 453134
rect 487794 417454 488414 452898
rect 487794 417218 487826 417454
rect 488062 417218 488146 417454
rect 488382 417218 488414 417454
rect 487794 417134 488414 417218
rect 487794 416898 487826 417134
rect 488062 416898 488146 417134
rect 488382 416898 488414 417134
rect 487794 381454 488414 416898
rect 487794 381218 487826 381454
rect 488062 381218 488146 381454
rect 488382 381218 488414 381454
rect 487794 381134 488414 381218
rect 487794 380898 487826 381134
rect 488062 380898 488146 381134
rect 488382 380898 488414 381134
rect 487794 345454 488414 380898
rect 487794 345218 487826 345454
rect 488062 345218 488146 345454
rect 488382 345218 488414 345454
rect 487794 345134 488414 345218
rect 487794 344898 487826 345134
rect 488062 344898 488146 345134
rect 488382 344898 488414 345134
rect 487794 309454 488414 344898
rect 487794 309218 487826 309454
rect 488062 309218 488146 309454
rect 488382 309218 488414 309454
rect 487794 309134 488414 309218
rect 487794 308898 487826 309134
rect 488062 308898 488146 309134
rect 488382 308898 488414 309134
rect 487794 273454 488414 308898
rect 487794 273218 487826 273454
rect 488062 273218 488146 273454
rect 488382 273218 488414 273454
rect 487794 273134 488414 273218
rect 487794 272898 487826 273134
rect 488062 272898 488146 273134
rect 488382 272898 488414 273134
rect 487794 237454 488414 272898
rect 487794 237218 487826 237454
rect 488062 237218 488146 237454
rect 488382 237218 488414 237454
rect 487794 237134 488414 237218
rect 487794 236898 487826 237134
rect 488062 236898 488146 237134
rect 488382 236898 488414 237134
rect 487794 201454 488414 236898
rect 487794 201218 487826 201454
rect 488062 201218 488146 201454
rect 488382 201218 488414 201454
rect 487794 201134 488414 201218
rect 487794 200898 487826 201134
rect 488062 200898 488146 201134
rect 488382 200898 488414 201134
rect 487794 165454 488414 200898
rect 487794 165218 487826 165454
rect 488062 165218 488146 165454
rect 488382 165218 488414 165454
rect 487794 165134 488414 165218
rect 487794 164898 487826 165134
rect 488062 164898 488146 165134
rect 488382 164898 488414 165134
rect 487794 129454 488414 164898
rect 487794 129218 487826 129454
rect 488062 129218 488146 129454
rect 488382 129218 488414 129454
rect 487794 129134 488414 129218
rect 487794 128898 487826 129134
rect 488062 128898 488146 129134
rect 488382 128898 488414 129134
rect 487794 93454 488414 128898
rect 487794 93218 487826 93454
rect 488062 93218 488146 93454
rect 488382 93218 488414 93454
rect 487794 93134 488414 93218
rect 487794 92898 487826 93134
rect 488062 92898 488146 93134
rect 488382 92898 488414 93134
rect 487794 57454 488414 92898
rect 487794 57218 487826 57454
rect 488062 57218 488146 57454
rect 488382 57218 488414 57454
rect 487794 57134 488414 57218
rect 487794 56898 487826 57134
rect 488062 56898 488146 57134
rect 488382 56898 488414 57134
rect 487794 21454 488414 56898
rect 487794 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 488414 21454
rect 487794 21134 488414 21218
rect 487794 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 488414 21134
rect 487794 -4186 488414 20898
rect 487794 -4422 487826 -4186
rect 488062 -4422 488146 -4186
rect 488382 -4422 488414 -4186
rect 487794 -4506 488414 -4422
rect 487794 -4742 487826 -4506
rect 488062 -4742 488146 -4506
rect 488382 -4742 488414 -4506
rect 487794 -7654 488414 -4742
rect 492294 709638 492914 711590
rect 492294 709402 492326 709638
rect 492562 709402 492646 709638
rect 492882 709402 492914 709638
rect 492294 709318 492914 709402
rect 492294 709082 492326 709318
rect 492562 709082 492646 709318
rect 492882 709082 492914 709318
rect 492294 673954 492914 709082
rect 492294 673718 492326 673954
rect 492562 673718 492646 673954
rect 492882 673718 492914 673954
rect 492294 673634 492914 673718
rect 492294 673398 492326 673634
rect 492562 673398 492646 673634
rect 492882 673398 492914 673634
rect 492294 637954 492914 673398
rect 492294 637718 492326 637954
rect 492562 637718 492646 637954
rect 492882 637718 492914 637954
rect 492294 637634 492914 637718
rect 492294 637398 492326 637634
rect 492562 637398 492646 637634
rect 492882 637398 492914 637634
rect 492294 601954 492914 637398
rect 492294 601718 492326 601954
rect 492562 601718 492646 601954
rect 492882 601718 492914 601954
rect 492294 601634 492914 601718
rect 492294 601398 492326 601634
rect 492562 601398 492646 601634
rect 492882 601398 492914 601634
rect 492294 565954 492914 601398
rect 492294 565718 492326 565954
rect 492562 565718 492646 565954
rect 492882 565718 492914 565954
rect 492294 565634 492914 565718
rect 492294 565398 492326 565634
rect 492562 565398 492646 565634
rect 492882 565398 492914 565634
rect 492294 529954 492914 565398
rect 492294 529718 492326 529954
rect 492562 529718 492646 529954
rect 492882 529718 492914 529954
rect 492294 529634 492914 529718
rect 492294 529398 492326 529634
rect 492562 529398 492646 529634
rect 492882 529398 492914 529634
rect 492294 493954 492914 529398
rect 492294 493718 492326 493954
rect 492562 493718 492646 493954
rect 492882 493718 492914 493954
rect 492294 493634 492914 493718
rect 492294 493398 492326 493634
rect 492562 493398 492646 493634
rect 492882 493398 492914 493634
rect 492294 457954 492914 493398
rect 492294 457718 492326 457954
rect 492562 457718 492646 457954
rect 492882 457718 492914 457954
rect 492294 457634 492914 457718
rect 492294 457398 492326 457634
rect 492562 457398 492646 457634
rect 492882 457398 492914 457634
rect 492294 421954 492914 457398
rect 492294 421718 492326 421954
rect 492562 421718 492646 421954
rect 492882 421718 492914 421954
rect 492294 421634 492914 421718
rect 492294 421398 492326 421634
rect 492562 421398 492646 421634
rect 492882 421398 492914 421634
rect 492294 385954 492914 421398
rect 492294 385718 492326 385954
rect 492562 385718 492646 385954
rect 492882 385718 492914 385954
rect 492294 385634 492914 385718
rect 492294 385398 492326 385634
rect 492562 385398 492646 385634
rect 492882 385398 492914 385634
rect 492294 349954 492914 385398
rect 492294 349718 492326 349954
rect 492562 349718 492646 349954
rect 492882 349718 492914 349954
rect 492294 349634 492914 349718
rect 492294 349398 492326 349634
rect 492562 349398 492646 349634
rect 492882 349398 492914 349634
rect 492294 313954 492914 349398
rect 492294 313718 492326 313954
rect 492562 313718 492646 313954
rect 492882 313718 492914 313954
rect 492294 313634 492914 313718
rect 492294 313398 492326 313634
rect 492562 313398 492646 313634
rect 492882 313398 492914 313634
rect 492294 277954 492914 313398
rect 492294 277718 492326 277954
rect 492562 277718 492646 277954
rect 492882 277718 492914 277954
rect 492294 277634 492914 277718
rect 492294 277398 492326 277634
rect 492562 277398 492646 277634
rect 492882 277398 492914 277634
rect 492294 241954 492914 277398
rect 492294 241718 492326 241954
rect 492562 241718 492646 241954
rect 492882 241718 492914 241954
rect 492294 241634 492914 241718
rect 492294 241398 492326 241634
rect 492562 241398 492646 241634
rect 492882 241398 492914 241634
rect 492294 205954 492914 241398
rect 492294 205718 492326 205954
rect 492562 205718 492646 205954
rect 492882 205718 492914 205954
rect 492294 205634 492914 205718
rect 492294 205398 492326 205634
rect 492562 205398 492646 205634
rect 492882 205398 492914 205634
rect 492294 169954 492914 205398
rect 492294 169718 492326 169954
rect 492562 169718 492646 169954
rect 492882 169718 492914 169954
rect 492294 169634 492914 169718
rect 492294 169398 492326 169634
rect 492562 169398 492646 169634
rect 492882 169398 492914 169634
rect 492294 133954 492914 169398
rect 492294 133718 492326 133954
rect 492562 133718 492646 133954
rect 492882 133718 492914 133954
rect 492294 133634 492914 133718
rect 492294 133398 492326 133634
rect 492562 133398 492646 133634
rect 492882 133398 492914 133634
rect 492294 97954 492914 133398
rect 492294 97718 492326 97954
rect 492562 97718 492646 97954
rect 492882 97718 492914 97954
rect 492294 97634 492914 97718
rect 492294 97398 492326 97634
rect 492562 97398 492646 97634
rect 492882 97398 492914 97634
rect 492294 61954 492914 97398
rect 492294 61718 492326 61954
rect 492562 61718 492646 61954
rect 492882 61718 492914 61954
rect 492294 61634 492914 61718
rect 492294 61398 492326 61634
rect 492562 61398 492646 61634
rect 492882 61398 492914 61634
rect 492294 25954 492914 61398
rect 492294 25718 492326 25954
rect 492562 25718 492646 25954
rect 492882 25718 492914 25954
rect 492294 25634 492914 25718
rect 492294 25398 492326 25634
rect 492562 25398 492646 25634
rect 492882 25398 492914 25634
rect 492294 -5146 492914 25398
rect 492294 -5382 492326 -5146
rect 492562 -5382 492646 -5146
rect 492882 -5382 492914 -5146
rect 492294 -5466 492914 -5382
rect 492294 -5702 492326 -5466
rect 492562 -5702 492646 -5466
rect 492882 -5702 492914 -5466
rect 492294 -7654 492914 -5702
rect 496794 710598 497414 711590
rect 496794 710362 496826 710598
rect 497062 710362 497146 710598
rect 497382 710362 497414 710598
rect 496794 710278 497414 710362
rect 496794 710042 496826 710278
rect 497062 710042 497146 710278
rect 497382 710042 497414 710278
rect 496794 678454 497414 710042
rect 496794 678218 496826 678454
rect 497062 678218 497146 678454
rect 497382 678218 497414 678454
rect 496794 678134 497414 678218
rect 496794 677898 496826 678134
rect 497062 677898 497146 678134
rect 497382 677898 497414 678134
rect 496794 642454 497414 677898
rect 496794 642218 496826 642454
rect 497062 642218 497146 642454
rect 497382 642218 497414 642454
rect 496794 642134 497414 642218
rect 496794 641898 496826 642134
rect 497062 641898 497146 642134
rect 497382 641898 497414 642134
rect 496794 606454 497414 641898
rect 496794 606218 496826 606454
rect 497062 606218 497146 606454
rect 497382 606218 497414 606454
rect 496794 606134 497414 606218
rect 496794 605898 496826 606134
rect 497062 605898 497146 606134
rect 497382 605898 497414 606134
rect 496794 570454 497414 605898
rect 496794 570218 496826 570454
rect 497062 570218 497146 570454
rect 497382 570218 497414 570454
rect 496794 570134 497414 570218
rect 496794 569898 496826 570134
rect 497062 569898 497146 570134
rect 497382 569898 497414 570134
rect 496794 534454 497414 569898
rect 496794 534218 496826 534454
rect 497062 534218 497146 534454
rect 497382 534218 497414 534454
rect 496794 534134 497414 534218
rect 496794 533898 496826 534134
rect 497062 533898 497146 534134
rect 497382 533898 497414 534134
rect 496794 498454 497414 533898
rect 496794 498218 496826 498454
rect 497062 498218 497146 498454
rect 497382 498218 497414 498454
rect 496794 498134 497414 498218
rect 496794 497898 496826 498134
rect 497062 497898 497146 498134
rect 497382 497898 497414 498134
rect 496794 462454 497414 497898
rect 496794 462218 496826 462454
rect 497062 462218 497146 462454
rect 497382 462218 497414 462454
rect 496794 462134 497414 462218
rect 496794 461898 496826 462134
rect 497062 461898 497146 462134
rect 497382 461898 497414 462134
rect 496794 426454 497414 461898
rect 496794 426218 496826 426454
rect 497062 426218 497146 426454
rect 497382 426218 497414 426454
rect 496794 426134 497414 426218
rect 496794 425898 496826 426134
rect 497062 425898 497146 426134
rect 497382 425898 497414 426134
rect 496794 390454 497414 425898
rect 496794 390218 496826 390454
rect 497062 390218 497146 390454
rect 497382 390218 497414 390454
rect 496794 390134 497414 390218
rect 496794 389898 496826 390134
rect 497062 389898 497146 390134
rect 497382 389898 497414 390134
rect 496794 354454 497414 389898
rect 496794 354218 496826 354454
rect 497062 354218 497146 354454
rect 497382 354218 497414 354454
rect 496794 354134 497414 354218
rect 496794 353898 496826 354134
rect 497062 353898 497146 354134
rect 497382 353898 497414 354134
rect 496794 318454 497414 353898
rect 496794 318218 496826 318454
rect 497062 318218 497146 318454
rect 497382 318218 497414 318454
rect 496794 318134 497414 318218
rect 496794 317898 496826 318134
rect 497062 317898 497146 318134
rect 497382 317898 497414 318134
rect 496794 282454 497414 317898
rect 496794 282218 496826 282454
rect 497062 282218 497146 282454
rect 497382 282218 497414 282454
rect 496794 282134 497414 282218
rect 496794 281898 496826 282134
rect 497062 281898 497146 282134
rect 497382 281898 497414 282134
rect 496794 246454 497414 281898
rect 496794 246218 496826 246454
rect 497062 246218 497146 246454
rect 497382 246218 497414 246454
rect 496794 246134 497414 246218
rect 496794 245898 496826 246134
rect 497062 245898 497146 246134
rect 497382 245898 497414 246134
rect 496794 210454 497414 245898
rect 496794 210218 496826 210454
rect 497062 210218 497146 210454
rect 497382 210218 497414 210454
rect 496794 210134 497414 210218
rect 496794 209898 496826 210134
rect 497062 209898 497146 210134
rect 497382 209898 497414 210134
rect 496794 174454 497414 209898
rect 496794 174218 496826 174454
rect 497062 174218 497146 174454
rect 497382 174218 497414 174454
rect 496794 174134 497414 174218
rect 496794 173898 496826 174134
rect 497062 173898 497146 174134
rect 497382 173898 497414 174134
rect 496794 138454 497414 173898
rect 496794 138218 496826 138454
rect 497062 138218 497146 138454
rect 497382 138218 497414 138454
rect 496794 138134 497414 138218
rect 496794 137898 496826 138134
rect 497062 137898 497146 138134
rect 497382 137898 497414 138134
rect 496794 102454 497414 137898
rect 496794 102218 496826 102454
rect 497062 102218 497146 102454
rect 497382 102218 497414 102454
rect 496794 102134 497414 102218
rect 496794 101898 496826 102134
rect 497062 101898 497146 102134
rect 497382 101898 497414 102134
rect 496794 66454 497414 101898
rect 496794 66218 496826 66454
rect 497062 66218 497146 66454
rect 497382 66218 497414 66454
rect 496794 66134 497414 66218
rect 496794 65898 496826 66134
rect 497062 65898 497146 66134
rect 497382 65898 497414 66134
rect 496794 30454 497414 65898
rect 496794 30218 496826 30454
rect 497062 30218 497146 30454
rect 497382 30218 497414 30454
rect 496794 30134 497414 30218
rect 496794 29898 496826 30134
rect 497062 29898 497146 30134
rect 497382 29898 497414 30134
rect 496794 -6106 497414 29898
rect 496794 -6342 496826 -6106
rect 497062 -6342 497146 -6106
rect 497382 -6342 497414 -6106
rect 496794 -6426 497414 -6342
rect 496794 -6662 496826 -6426
rect 497062 -6662 497146 -6426
rect 497382 -6662 497414 -6426
rect 496794 -7654 497414 -6662
rect 501294 711558 501914 711590
rect 501294 711322 501326 711558
rect 501562 711322 501646 711558
rect 501882 711322 501914 711558
rect 501294 711238 501914 711322
rect 501294 711002 501326 711238
rect 501562 711002 501646 711238
rect 501882 711002 501914 711238
rect 501294 682954 501914 711002
rect 501294 682718 501326 682954
rect 501562 682718 501646 682954
rect 501882 682718 501914 682954
rect 501294 682634 501914 682718
rect 501294 682398 501326 682634
rect 501562 682398 501646 682634
rect 501882 682398 501914 682634
rect 501294 646954 501914 682398
rect 501294 646718 501326 646954
rect 501562 646718 501646 646954
rect 501882 646718 501914 646954
rect 501294 646634 501914 646718
rect 501294 646398 501326 646634
rect 501562 646398 501646 646634
rect 501882 646398 501914 646634
rect 501294 610954 501914 646398
rect 501294 610718 501326 610954
rect 501562 610718 501646 610954
rect 501882 610718 501914 610954
rect 501294 610634 501914 610718
rect 501294 610398 501326 610634
rect 501562 610398 501646 610634
rect 501882 610398 501914 610634
rect 501294 574954 501914 610398
rect 501294 574718 501326 574954
rect 501562 574718 501646 574954
rect 501882 574718 501914 574954
rect 501294 574634 501914 574718
rect 501294 574398 501326 574634
rect 501562 574398 501646 574634
rect 501882 574398 501914 574634
rect 501294 538954 501914 574398
rect 501294 538718 501326 538954
rect 501562 538718 501646 538954
rect 501882 538718 501914 538954
rect 501294 538634 501914 538718
rect 501294 538398 501326 538634
rect 501562 538398 501646 538634
rect 501882 538398 501914 538634
rect 501294 502954 501914 538398
rect 501294 502718 501326 502954
rect 501562 502718 501646 502954
rect 501882 502718 501914 502954
rect 501294 502634 501914 502718
rect 501294 502398 501326 502634
rect 501562 502398 501646 502634
rect 501882 502398 501914 502634
rect 501294 466954 501914 502398
rect 501294 466718 501326 466954
rect 501562 466718 501646 466954
rect 501882 466718 501914 466954
rect 501294 466634 501914 466718
rect 501294 466398 501326 466634
rect 501562 466398 501646 466634
rect 501882 466398 501914 466634
rect 501294 430954 501914 466398
rect 501294 430718 501326 430954
rect 501562 430718 501646 430954
rect 501882 430718 501914 430954
rect 501294 430634 501914 430718
rect 501294 430398 501326 430634
rect 501562 430398 501646 430634
rect 501882 430398 501914 430634
rect 501294 394954 501914 430398
rect 501294 394718 501326 394954
rect 501562 394718 501646 394954
rect 501882 394718 501914 394954
rect 501294 394634 501914 394718
rect 501294 394398 501326 394634
rect 501562 394398 501646 394634
rect 501882 394398 501914 394634
rect 501294 358954 501914 394398
rect 501294 358718 501326 358954
rect 501562 358718 501646 358954
rect 501882 358718 501914 358954
rect 501294 358634 501914 358718
rect 501294 358398 501326 358634
rect 501562 358398 501646 358634
rect 501882 358398 501914 358634
rect 501294 322954 501914 358398
rect 501294 322718 501326 322954
rect 501562 322718 501646 322954
rect 501882 322718 501914 322954
rect 501294 322634 501914 322718
rect 501294 322398 501326 322634
rect 501562 322398 501646 322634
rect 501882 322398 501914 322634
rect 501294 286954 501914 322398
rect 501294 286718 501326 286954
rect 501562 286718 501646 286954
rect 501882 286718 501914 286954
rect 501294 286634 501914 286718
rect 501294 286398 501326 286634
rect 501562 286398 501646 286634
rect 501882 286398 501914 286634
rect 501294 250954 501914 286398
rect 501294 250718 501326 250954
rect 501562 250718 501646 250954
rect 501882 250718 501914 250954
rect 501294 250634 501914 250718
rect 501294 250398 501326 250634
rect 501562 250398 501646 250634
rect 501882 250398 501914 250634
rect 501294 214954 501914 250398
rect 501294 214718 501326 214954
rect 501562 214718 501646 214954
rect 501882 214718 501914 214954
rect 501294 214634 501914 214718
rect 501294 214398 501326 214634
rect 501562 214398 501646 214634
rect 501882 214398 501914 214634
rect 501294 178954 501914 214398
rect 501294 178718 501326 178954
rect 501562 178718 501646 178954
rect 501882 178718 501914 178954
rect 501294 178634 501914 178718
rect 501294 178398 501326 178634
rect 501562 178398 501646 178634
rect 501882 178398 501914 178634
rect 501294 142954 501914 178398
rect 501294 142718 501326 142954
rect 501562 142718 501646 142954
rect 501882 142718 501914 142954
rect 501294 142634 501914 142718
rect 501294 142398 501326 142634
rect 501562 142398 501646 142634
rect 501882 142398 501914 142634
rect 501294 106954 501914 142398
rect 501294 106718 501326 106954
rect 501562 106718 501646 106954
rect 501882 106718 501914 106954
rect 501294 106634 501914 106718
rect 501294 106398 501326 106634
rect 501562 106398 501646 106634
rect 501882 106398 501914 106634
rect 501294 70954 501914 106398
rect 501294 70718 501326 70954
rect 501562 70718 501646 70954
rect 501882 70718 501914 70954
rect 501294 70634 501914 70718
rect 501294 70398 501326 70634
rect 501562 70398 501646 70634
rect 501882 70398 501914 70634
rect 501294 34954 501914 70398
rect 501294 34718 501326 34954
rect 501562 34718 501646 34954
rect 501882 34718 501914 34954
rect 501294 34634 501914 34718
rect 501294 34398 501326 34634
rect 501562 34398 501646 34634
rect 501882 34398 501914 34634
rect 501294 -7066 501914 34398
rect 501294 -7302 501326 -7066
rect 501562 -7302 501646 -7066
rect 501882 -7302 501914 -7066
rect 501294 -7386 501914 -7302
rect 501294 -7622 501326 -7386
rect 501562 -7622 501646 -7386
rect 501882 -7622 501914 -7386
rect 501294 -7654 501914 -7622
rect 505794 704838 506414 711590
rect 505794 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 506414 704838
rect 505794 704518 506414 704602
rect 505794 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 506414 704518
rect 505794 687454 506414 704282
rect 505794 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 506414 687454
rect 505794 687134 506414 687218
rect 505794 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 506414 687134
rect 505794 651454 506414 686898
rect 505794 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 506414 651454
rect 505794 651134 506414 651218
rect 505794 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 506414 651134
rect 505794 615454 506414 650898
rect 505794 615218 505826 615454
rect 506062 615218 506146 615454
rect 506382 615218 506414 615454
rect 505794 615134 506414 615218
rect 505794 614898 505826 615134
rect 506062 614898 506146 615134
rect 506382 614898 506414 615134
rect 505794 579454 506414 614898
rect 505794 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 506414 579454
rect 505794 579134 506414 579218
rect 505794 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 506414 579134
rect 505794 543454 506414 578898
rect 505794 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 506414 543454
rect 505794 543134 506414 543218
rect 505794 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 506414 543134
rect 505794 507454 506414 542898
rect 505794 507218 505826 507454
rect 506062 507218 506146 507454
rect 506382 507218 506414 507454
rect 505794 507134 506414 507218
rect 505794 506898 505826 507134
rect 506062 506898 506146 507134
rect 506382 506898 506414 507134
rect 505794 471454 506414 506898
rect 505794 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 506414 471454
rect 505794 471134 506414 471218
rect 505794 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 506414 471134
rect 505794 435454 506414 470898
rect 505794 435218 505826 435454
rect 506062 435218 506146 435454
rect 506382 435218 506414 435454
rect 505794 435134 506414 435218
rect 505794 434898 505826 435134
rect 506062 434898 506146 435134
rect 506382 434898 506414 435134
rect 505794 399454 506414 434898
rect 505794 399218 505826 399454
rect 506062 399218 506146 399454
rect 506382 399218 506414 399454
rect 505794 399134 506414 399218
rect 505794 398898 505826 399134
rect 506062 398898 506146 399134
rect 506382 398898 506414 399134
rect 505794 363454 506414 398898
rect 505794 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 506414 363454
rect 505794 363134 506414 363218
rect 505794 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 506414 363134
rect 505794 327454 506414 362898
rect 505794 327218 505826 327454
rect 506062 327218 506146 327454
rect 506382 327218 506414 327454
rect 505794 327134 506414 327218
rect 505794 326898 505826 327134
rect 506062 326898 506146 327134
rect 506382 326898 506414 327134
rect 505794 291454 506414 326898
rect 505794 291218 505826 291454
rect 506062 291218 506146 291454
rect 506382 291218 506414 291454
rect 505794 291134 506414 291218
rect 505794 290898 505826 291134
rect 506062 290898 506146 291134
rect 506382 290898 506414 291134
rect 505794 255454 506414 290898
rect 505794 255218 505826 255454
rect 506062 255218 506146 255454
rect 506382 255218 506414 255454
rect 505794 255134 506414 255218
rect 505794 254898 505826 255134
rect 506062 254898 506146 255134
rect 506382 254898 506414 255134
rect 505794 219454 506414 254898
rect 505794 219218 505826 219454
rect 506062 219218 506146 219454
rect 506382 219218 506414 219454
rect 505794 219134 506414 219218
rect 505794 218898 505826 219134
rect 506062 218898 506146 219134
rect 506382 218898 506414 219134
rect 505794 183454 506414 218898
rect 505794 183218 505826 183454
rect 506062 183218 506146 183454
rect 506382 183218 506414 183454
rect 505794 183134 506414 183218
rect 505794 182898 505826 183134
rect 506062 182898 506146 183134
rect 506382 182898 506414 183134
rect 505794 147454 506414 182898
rect 505794 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 506414 147454
rect 505794 147134 506414 147218
rect 505794 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 506414 147134
rect 505794 111454 506414 146898
rect 505794 111218 505826 111454
rect 506062 111218 506146 111454
rect 506382 111218 506414 111454
rect 505794 111134 506414 111218
rect 505794 110898 505826 111134
rect 506062 110898 506146 111134
rect 506382 110898 506414 111134
rect 505794 75454 506414 110898
rect 505794 75218 505826 75454
rect 506062 75218 506146 75454
rect 506382 75218 506414 75454
rect 505794 75134 506414 75218
rect 505794 74898 505826 75134
rect 506062 74898 506146 75134
rect 506382 74898 506414 75134
rect 505794 39454 506414 74898
rect 505794 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 506414 39454
rect 505794 39134 506414 39218
rect 505794 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 506414 39134
rect 505794 3454 506414 38898
rect 505794 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 506414 3454
rect 505794 3134 506414 3218
rect 505794 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 506414 3134
rect 505794 -346 506414 2898
rect 505794 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 506414 -346
rect 505794 -666 506414 -582
rect 505794 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 506414 -666
rect 505794 -7654 506414 -902
rect 510294 705798 510914 711590
rect 510294 705562 510326 705798
rect 510562 705562 510646 705798
rect 510882 705562 510914 705798
rect 510294 705478 510914 705562
rect 510294 705242 510326 705478
rect 510562 705242 510646 705478
rect 510882 705242 510914 705478
rect 510294 691954 510914 705242
rect 510294 691718 510326 691954
rect 510562 691718 510646 691954
rect 510882 691718 510914 691954
rect 510294 691634 510914 691718
rect 510294 691398 510326 691634
rect 510562 691398 510646 691634
rect 510882 691398 510914 691634
rect 510294 655954 510914 691398
rect 510294 655718 510326 655954
rect 510562 655718 510646 655954
rect 510882 655718 510914 655954
rect 510294 655634 510914 655718
rect 510294 655398 510326 655634
rect 510562 655398 510646 655634
rect 510882 655398 510914 655634
rect 510294 619954 510914 655398
rect 510294 619718 510326 619954
rect 510562 619718 510646 619954
rect 510882 619718 510914 619954
rect 510294 619634 510914 619718
rect 510294 619398 510326 619634
rect 510562 619398 510646 619634
rect 510882 619398 510914 619634
rect 510294 583954 510914 619398
rect 510294 583718 510326 583954
rect 510562 583718 510646 583954
rect 510882 583718 510914 583954
rect 510294 583634 510914 583718
rect 510294 583398 510326 583634
rect 510562 583398 510646 583634
rect 510882 583398 510914 583634
rect 510294 547954 510914 583398
rect 510294 547718 510326 547954
rect 510562 547718 510646 547954
rect 510882 547718 510914 547954
rect 510294 547634 510914 547718
rect 510294 547398 510326 547634
rect 510562 547398 510646 547634
rect 510882 547398 510914 547634
rect 510294 511954 510914 547398
rect 510294 511718 510326 511954
rect 510562 511718 510646 511954
rect 510882 511718 510914 511954
rect 510294 511634 510914 511718
rect 510294 511398 510326 511634
rect 510562 511398 510646 511634
rect 510882 511398 510914 511634
rect 510294 475954 510914 511398
rect 510294 475718 510326 475954
rect 510562 475718 510646 475954
rect 510882 475718 510914 475954
rect 510294 475634 510914 475718
rect 510294 475398 510326 475634
rect 510562 475398 510646 475634
rect 510882 475398 510914 475634
rect 510294 439954 510914 475398
rect 510294 439718 510326 439954
rect 510562 439718 510646 439954
rect 510882 439718 510914 439954
rect 510294 439634 510914 439718
rect 510294 439398 510326 439634
rect 510562 439398 510646 439634
rect 510882 439398 510914 439634
rect 510294 403954 510914 439398
rect 510294 403718 510326 403954
rect 510562 403718 510646 403954
rect 510882 403718 510914 403954
rect 510294 403634 510914 403718
rect 510294 403398 510326 403634
rect 510562 403398 510646 403634
rect 510882 403398 510914 403634
rect 510294 367954 510914 403398
rect 510294 367718 510326 367954
rect 510562 367718 510646 367954
rect 510882 367718 510914 367954
rect 510294 367634 510914 367718
rect 510294 367398 510326 367634
rect 510562 367398 510646 367634
rect 510882 367398 510914 367634
rect 510294 331954 510914 367398
rect 510294 331718 510326 331954
rect 510562 331718 510646 331954
rect 510882 331718 510914 331954
rect 510294 331634 510914 331718
rect 510294 331398 510326 331634
rect 510562 331398 510646 331634
rect 510882 331398 510914 331634
rect 510294 295954 510914 331398
rect 510294 295718 510326 295954
rect 510562 295718 510646 295954
rect 510882 295718 510914 295954
rect 510294 295634 510914 295718
rect 510294 295398 510326 295634
rect 510562 295398 510646 295634
rect 510882 295398 510914 295634
rect 510294 259954 510914 295398
rect 510294 259718 510326 259954
rect 510562 259718 510646 259954
rect 510882 259718 510914 259954
rect 510294 259634 510914 259718
rect 510294 259398 510326 259634
rect 510562 259398 510646 259634
rect 510882 259398 510914 259634
rect 510294 223954 510914 259398
rect 510294 223718 510326 223954
rect 510562 223718 510646 223954
rect 510882 223718 510914 223954
rect 510294 223634 510914 223718
rect 510294 223398 510326 223634
rect 510562 223398 510646 223634
rect 510882 223398 510914 223634
rect 510294 187954 510914 223398
rect 510294 187718 510326 187954
rect 510562 187718 510646 187954
rect 510882 187718 510914 187954
rect 510294 187634 510914 187718
rect 510294 187398 510326 187634
rect 510562 187398 510646 187634
rect 510882 187398 510914 187634
rect 510294 151954 510914 187398
rect 510294 151718 510326 151954
rect 510562 151718 510646 151954
rect 510882 151718 510914 151954
rect 510294 151634 510914 151718
rect 510294 151398 510326 151634
rect 510562 151398 510646 151634
rect 510882 151398 510914 151634
rect 510294 115954 510914 151398
rect 510294 115718 510326 115954
rect 510562 115718 510646 115954
rect 510882 115718 510914 115954
rect 510294 115634 510914 115718
rect 510294 115398 510326 115634
rect 510562 115398 510646 115634
rect 510882 115398 510914 115634
rect 510294 79954 510914 115398
rect 510294 79718 510326 79954
rect 510562 79718 510646 79954
rect 510882 79718 510914 79954
rect 510294 79634 510914 79718
rect 510294 79398 510326 79634
rect 510562 79398 510646 79634
rect 510882 79398 510914 79634
rect 510294 43954 510914 79398
rect 510294 43718 510326 43954
rect 510562 43718 510646 43954
rect 510882 43718 510914 43954
rect 510294 43634 510914 43718
rect 510294 43398 510326 43634
rect 510562 43398 510646 43634
rect 510882 43398 510914 43634
rect 510294 7954 510914 43398
rect 510294 7718 510326 7954
rect 510562 7718 510646 7954
rect 510882 7718 510914 7954
rect 510294 7634 510914 7718
rect 510294 7398 510326 7634
rect 510562 7398 510646 7634
rect 510882 7398 510914 7634
rect 510294 -1306 510914 7398
rect 510294 -1542 510326 -1306
rect 510562 -1542 510646 -1306
rect 510882 -1542 510914 -1306
rect 510294 -1626 510914 -1542
rect 510294 -1862 510326 -1626
rect 510562 -1862 510646 -1626
rect 510882 -1862 510914 -1626
rect 510294 -7654 510914 -1862
rect 514794 706758 515414 711590
rect 514794 706522 514826 706758
rect 515062 706522 515146 706758
rect 515382 706522 515414 706758
rect 514794 706438 515414 706522
rect 514794 706202 514826 706438
rect 515062 706202 515146 706438
rect 515382 706202 515414 706438
rect 514794 696454 515414 706202
rect 514794 696218 514826 696454
rect 515062 696218 515146 696454
rect 515382 696218 515414 696454
rect 514794 696134 515414 696218
rect 514794 695898 514826 696134
rect 515062 695898 515146 696134
rect 515382 695898 515414 696134
rect 514794 660454 515414 695898
rect 514794 660218 514826 660454
rect 515062 660218 515146 660454
rect 515382 660218 515414 660454
rect 514794 660134 515414 660218
rect 514794 659898 514826 660134
rect 515062 659898 515146 660134
rect 515382 659898 515414 660134
rect 514794 624454 515414 659898
rect 514794 624218 514826 624454
rect 515062 624218 515146 624454
rect 515382 624218 515414 624454
rect 514794 624134 515414 624218
rect 514794 623898 514826 624134
rect 515062 623898 515146 624134
rect 515382 623898 515414 624134
rect 514794 588454 515414 623898
rect 514794 588218 514826 588454
rect 515062 588218 515146 588454
rect 515382 588218 515414 588454
rect 514794 588134 515414 588218
rect 514794 587898 514826 588134
rect 515062 587898 515146 588134
rect 515382 587898 515414 588134
rect 514794 552454 515414 587898
rect 514794 552218 514826 552454
rect 515062 552218 515146 552454
rect 515382 552218 515414 552454
rect 514794 552134 515414 552218
rect 514794 551898 514826 552134
rect 515062 551898 515146 552134
rect 515382 551898 515414 552134
rect 514794 516454 515414 551898
rect 514794 516218 514826 516454
rect 515062 516218 515146 516454
rect 515382 516218 515414 516454
rect 514794 516134 515414 516218
rect 514794 515898 514826 516134
rect 515062 515898 515146 516134
rect 515382 515898 515414 516134
rect 514794 480454 515414 515898
rect 514794 480218 514826 480454
rect 515062 480218 515146 480454
rect 515382 480218 515414 480454
rect 514794 480134 515414 480218
rect 514794 479898 514826 480134
rect 515062 479898 515146 480134
rect 515382 479898 515414 480134
rect 514794 444454 515414 479898
rect 514794 444218 514826 444454
rect 515062 444218 515146 444454
rect 515382 444218 515414 444454
rect 514794 444134 515414 444218
rect 514794 443898 514826 444134
rect 515062 443898 515146 444134
rect 515382 443898 515414 444134
rect 514794 408454 515414 443898
rect 514794 408218 514826 408454
rect 515062 408218 515146 408454
rect 515382 408218 515414 408454
rect 514794 408134 515414 408218
rect 514794 407898 514826 408134
rect 515062 407898 515146 408134
rect 515382 407898 515414 408134
rect 514794 372454 515414 407898
rect 514794 372218 514826 372454
rect 515062 372218 515146 372454
rect 515382 372218 515414 372454
rect 514794 372134 515414 372218
rect 514794 371898 514826 372134
rect 515062 371898 515146 372134
rect 515382 371898 515414 372134
rect 514794 336454 515414 371898
rect 514794 336218 514826 336454
rect 515062 336218 515146 336454
rect 515382 336218 515414 336454
rect 514794 336134 515414 336218
rect 514794 335898 514826 336134
rect 515062 335898 515146 336134
rect 515382 335898 515414 336134
rect 514794 300454 515414 335898
rect 514794 300218 514826 300454
rect 515062 300218 515146 300454
rect 515382 300218 515414 300454
rect 514794 300134 515414 300218
rect 514794 299898 514826 300134
rect 515062 299898 515146 300134
rect 515382 299898 515414 300134
rect 514794 264454 515414 299898
rect 514794 264218 514826 264454
rect 515062 264218 515146 264454
rect 515382 264218 515414 264454
rect 514794 264134 515414 264218
rect 514794 263898 514826 264134
rect 515062 263898 515146 264134
rect 515382 263898 515414 264134
rect 514794 228454 515414 263898
rect 514794 228218 514826 228454
rect 515062 228218 515146 228454
rect 515382 228218 515414 228454
rect 514794 228134 515414 228218
rect 514794 227898 514826 228134
rect 515062 227898 515146 228134
rect 515382 227898 515414 228134
rect 514794 192454 515414 227898
rect 514794 192218 514826 192454
rect 515062 192218 515146 192454
rect 515382 192218 515414 192454
rect 514794 192134 515414 192218
rect 514794 191898 514826 192134
rect 515062 191898 515146 192134
rect 515382 191898 515414 192134
rect 514794 156454 515414 191898
rect 514794 156218 514826 156454
rect 515062 156218 515146 156454
rect 515382 156218 515414 156454
rect 514794 156134 515414 156218
rect 514794 155898 514826 156134
rect 515062 155898 515146 156134
rect 515382 155898 515414 156134
rect 514794 120454 515414 155898
rect 514794 120218 514826 120454
rect 515062 120218 515146 120454
rect 515382 120218 515414 120454
rect 514794 120134 515414 120218
rect 514794 119898 514826 120134
rect 515062 119898 515146 120134
rect 515382 119898 515414 120134
rect 514794 84454 515414 119898
rect 514794 84218 514826 84454
rect 515062 84218 515146 84454
rect 515382 84218 515414 84454
rect 514794 84134 515414 84218
rect 514794 83898 514826 84134
rect 515062 83898 515146 84134
rect 515382 83898 515414 84134
rect 514794 48454 515414 83898
rect 514794 48218 514826 48454
rect 515062 48218 515146 48454
rect 515382 48218 515414 48454
rect 514794 48134 515414 48218
rect 514794 47898 514826 48134
rect 515062 47898 515146 48134
rect 515382 47898 515414 48134
rect 514794 12454 515414 47898
rect 514794 12218 514826 12454
rect 515062 12218 515146 12454
rect 515382 12218 515414 12454
rect 514794 12134 515414 12218
rect 514794 11898 514826 12134
rect 515062 11898 515146 12134
rect 515382 11898 515414 12134
rect 514794 -2266 515414 11898
rect 514794 -2502 514826 -2266
rect 515062 -2502 515146 -2266
rect 515382 -2502 515414 -2266
rect 514794 -2586 515414 -2502
rect 514794 -2822 514826 -2586
rect 515062 -2822 515146 -2586
rect 515382 -2822 515414 -2586
rect 514794 -7654 515414 -2822
rect 519294 707718 519914 711590
rect 519294 707482 519326 707718
rect 519562 707482 519646 707718
rect 519882 707482 519914 707718
rect 519294 707398 519914 707482
rect 519294 707162 519326 707398
rect 519562 707162 519646 707398
rect 519882 707162 519914 707398
rect 519294 700954 519914 707162
rect 519294 700718 519326 700954
rect 519562 700718 519646 700954
rect 519882 700718 519914 700954
rect 519294 700634 519914 700718
rect 519294 700398 519326 700634
rect 519562 700398 519646 700634
rect 519882 700398 519914 700634
rect 519294 664954 519914 700398
rect 519294 664718 519326 664954
rect 519562 664718 519646 664954
rect 519882 664718 519914 664954
rect 519294 664634 519914 664718
rect 519294 664398 519326 664634
rect 519562 664398 519646 664634
rect 519882 664398 519914 664634
rect 519294 628954 519914 664398
rect 519294 628718 519326 628954
rect 519562 628718 519646 628954
rect 519882 628718 519914 628954
rect 519294 628634 519914 628718
rect 519294 628398 519326 628634
rect 519562 628398 519646 628634
rect 519882 628398 519914 628634
rect 519294 592954 519914 628398
rect 519294 592718 519326 592954
rect 519562 592718 519646 592954
rect 519882 592718 519914 592954
rect 519294 592634 519914 592718
rect 519294 592398 519326 592634
rect 519562 592398 519646 592634
rect 519882 592398 519914 592634
rect 519294 556954 519914 592398
rect 519294 556718 519326 556954
rect 519562 556718 519646 556954
rect 519882 556718 519914 556954
rect 519294 556634 519914 556718
rect 519294 556398 519326 556634
rect 519562 556398 519646 556634
rect 519882 556398 519914 556634
rect 519294 520954 519914 556398
rect 519294 520718 519326 520954
rect 519562 520718 519646 520954
rect 519882 520718 519914 520954
rect 519294 520634 519914 520718
rect 519294 520398 519326 520634
rect 519562 520398 519646 520634
rect 519882 520398 519914 520634
rect 519294 484954 519914 520398
rect 519294 484718 519326 484954
rect 519562 484718 519646 484954
rect 519882 484718 519914 484954
rect 519294 484634 519914 484718
rect 519294 484398 519326 484634
rect 519562 484398 519646 484634
rect 519882 484398 519914 484634
rect 519294 448954 519914 484398
rect 519294 448718 519326 448954
rect 519562 448718 519646 448954
rect 519882 448718 519914 448954
rect 519294 448634 519914 448718
rect 519294 448398 519326 448634
rect 519562 448398 519646 448634
rect 519882 448398 519914 448634
rect 519294 412954 519914 448398
rect 519294 412718 519326 412954
rect 519562 412718 519646 412954
rect 519882 412718 519914 412954
rect 519294 412634 519914 412718
rect 519294 412398 519326 412634
rect 519562 412398 519646 412634
rect 519882 412398 519914 412634
rect 519294 376954 519914 412398
rect 519294 376718 519326 376954
rect 519562 376718 519646 376954
rect 519882 376718 519914 376954
rect 519294 376634 519914 376718
rect 519294 376398 519326 376634
rect 519562 376398 519646 376634
rect 519882 376398 519914 376634
rect 519294 340954 519914 376398
rect 519294 340718 519326 340954
rect 519562 340718 519646 340954
rect 519882 340718 519914 340954
rect 519294 340634 519914 340718
rect 519294 340398 519326 340634
rect 519562 340398 519646 340634
rect 519882 340398 519914 340634
rect 519294 304954 519914 340398
rect 519294 304718 519326 304954
rect 519562 304718 519646 304954
rect 519882 304718 519914 304954
rect 519294 304634 519914 304718
rect 519294 304398 519326 304634
rect 519562 304398 519646 304634
rect 519882 304398 519914 304634
rect 519294 268954 519914 304398
rect 519294 268718 519326 268954
rect 519562 268718 519646 268954
rect 519882 268718 519914 268954
rect 519294 268634 519914 268718
rect 519294 268398 519326 268634
rect 519562 268398 519646 268634
rect 519882 268398 519914 268634
rect 519294 232954 519914 268398
rect 519294 232718 519326 232954
rect 519562 232718 519646 232954
rect 519882 232718 519914 232954
rect 519294 232634 519914 232718
rect 519294 232398 519326 232634
rect 519562 232398 519646 232634
rect 519882 232398 519914 232634
rect 519294 196954 519914 232398
rect 519294 196718 519326 196954
rect 519562 196718 519646 196954
rect 519882 196718 519914 196954
rect 519294 196634 519914 196718
rect 519294 196398 519326 196634
rect 519562 196398 519646 196634
rect 519882 196398 519914 196634
rect 519294 160954 519914 196398
rect 519294 160718 519326 160954
rect 519562 160718 519646 160954
rect 519882 160718 519914 160954
rect 519294 160634 519914 160718
rect 519294 160398 519326 160634
rect 519562 160398 519646 160634
rect 519882 160398 519914 160634
rect 519294 124954 519914 160398
rect 519294 124718 519326 124954
rect 519562 124718 519646 124954
rect 519882 124718 519914 124954
rect 519294 124634 519914 124718
rect 519294 124398 519326 124634
rect 519562 124398 519646 124634
rect 519882 124398 519914 124634
rect 519294 88954 519914 124398
rect 519294 88718 519326 88954
rect 519562 88718 519646 88954
rect 519882 88718 519914 88954
rect 519294 88634 519914 88718
rect 519294 88398 519326 88634
rect 519562 88398 519646 88634
rect 519882 88398 519914 88634
rect 519294 52954 519914 88398
rect 519294 52718 519326 52954
rect 519562 52718 519646 52954
rect 519882 52718 519914 52954
rect 519294 52634 519914 52718
rect 519294 52398 519326 52634
rect 519562 52398 519646 52634
rect 519882 52398 519914 52634
rect 519294 16954 519914 52398
rect 519294 16718 519326 16954
rect 519562 16718 519646 16954
rect 519882 16718 519914 16954
rect 519294 16634 519914 16718
rect 519294 16398 519326 16634
rect 519562 16398 519646 16634
rect 519882 16398 519914 16634
rect 519294 -3226 519914 16398
rect 519294 -3462 519326 -3226
rect 519562 -3462 519646 -3226
rect 519882 -3462 519914 -3226
rect 519294 -3546 519914 -3462
rect 519294 -3782 519326 -3546
rect 519562 -3782 519646 -3546
rect 519882 -3782 519914 -3546
rect 519294 -7654 519914 -3782
rect 523794 708678 524414 711590
rect 523794 708442 523826 708678
rect 524062 708442 524146 708678
rect 524382 708442 524414 708678
rect 523794 708358 524414 708442
rect 523794 708122 523826 708358
rect 524062 708122 524146 708358
rect 524382 708122 524414 708358
rect 523794 669454 524414 708122
rect 523794 669218 523826 669454
rect 524062 669218 524146 669454
rect 524382 669218 524414 669454
rect 523794 669134 524414 669218
rect 523794 668898 523826 669134
rect 524062 668898 524146 669134
rect 524382 668898 524414 669134
rect 523794 633454 524414 668898
rect 523794 633218 523826 633454
rect 524062 633218 524146 633454
rect 524382 633218 524414 633454
rect 523794 633134 524414 633218
rect 523794 632898 523826 633134
rect 524062 632898 524146 633134
rect 524382 632898 524414 633134
rect 523794 597454 524414 632898
rect 523794 597218 523826 597454
rect 524062 597218 524146 597454
rect 524382 597218 524414 597454
rect 523794 597134 524414 597218
rect 523794 596898 523826 597134
rect 524062 596898 524146 597134
rect 524382 596898 524414 597134
rect 523794 561454 524414 596898
rect 523794 561218 523826 561454
rect 524062 561218 524146 561454
rect 524382 561218 524414 561454
rect 523794 561134 524414 561218
rect 523794 560898 523826 561134
rect 524062 560898 524146 561134
rect 524382 560898 524414 561134
rect 523794 525454 524414 560898
rect 523794 525218 523826 525454
rect 524062 525218 524146 525454
rect 524382 525218 524414 525454
rect 523794 525134 524414 525218
rect 523794 524898 523826 525134
rect 524062 524898 524146 525134
rect 524382 524898 524414 525134
rect 523794 489454 524414 524898
rect 523794 489218 523826 489454
rect 524062 489218 524146 489454
rect 524382 489218 524414 489454
rect 523794 489134 524414 489218
rect 523794 488898 523826 489134
rect 524062 488898 524146 489134
rect 524382 488898 524414 489134
rect 523794 453454 524414 488898
rect 523794 453218 523826 453454
rect 524062 453218 524146 453454
rect 524382 453218 524414 453454
rect 523794 453134 524414 453218
rect 523794 452898 523826 453134
rect 524062 452898 524146 453134
rect 524382 452898 524414 453134
rect 523794 417454 524414 452898
rect 523794 417218 523826 417454
rect 524062 417218 524146 417454
rect 524382 417218 524414 417454
rect 523794 417134 524414 417218
rect 523794 416898 523826 417134
rect 524062 416898 524146 417134
rect 524382 416898 524414 417134
rect 523794 381454 524414 416898
rect 523794 381218 523826 381454
rect 524062 381218 524146 381454
rect 524382 381218 524414 381454
rect 523794 381134 524414 381218
rect 523794 380898 523826 381134
rect 524062 380898 524146 381134
rect 524382 380898 524414 381134
rect 523794 345454 524414 380898
rect 523794 345218 523826 345454
rect 524062 345218 524146 345454
rect 524382 345218 524414 345454
rect 523794 345134 524414 345218
rect 523794 344898 523826 345134
rect 524062 344898 524146 345134
rect 524382 344898 524414 345134
rect 523794 309454 524414 344898
rect 523794 309218 523826 309454
rect 524062 309218 524146 309454
rect 524382 309218 524414 309454
rect 523794 309134 524414 309218
rect 523794 308898 523826 309134
rect 524062 308898 524146 309134
rect 524382 308898 524414 309134
rect 523794 273454 524414 308898
rect 523794 273218 523826 273454
rect 524062 273218 524146 273454
rect 524382 273218 524414 273454
rect 523794 273134 524414 273218
rect 523794 272898 523826 273134
rect 524062 272898 524146 273134
rect 524382 272898 524414 273134
rect 523794 237454 524414 272898
rect 523794 237218 523826 237454
rect 524062 237218 524146 237454
rect 524382 237218 524414 237454
rect 523794 237134 524414 237218
rect 523794 236898 523826 237134
rect 524062 236898 524146 237134
rect 524382 236898 524414 237134
rect 523794 201454 524414 236898
rect 523794 201218 523826 201454
rect 524062 201218 524146 201454
rect 524382 201218 524414 201454
rect 523794 201134 524414 201218
rect 523794 200898 523826 201134
rect 524062 200898 524146 201134
rect 524382 200898 524414 201134
rect 523794 165454 524414 200898
rect 523794 165218 523826 165454
rect 524062 165218 524146 165454
rect 524382 165218 524414 165454
rect 523794 165134 524414 165218
rect 523794 164898 523826 165134
rect 524062 164898 524146 165134
rect 524382 164898 524414 165134
rect 523794 129454 524414 164898
rect 523794 129218 523826 129454
rect 524062 129218 524146 129454
rect 524382 129218 524414 129454
rect 523794 129134 524414 129218
rect 523794 128898 523826 129134
rect 524062 128898 524146 129134
rect 524382 128898 524414 129134
rect 523794 93454 524414 128898
rect 523794 93218 523826 93454
rect 524062 93218 524146 93454
rect 524382 93218 524414 93454
rect 523794 93134 524414 93218
rect 523794 92898 523826 93134
rect 524062 92898 524146 93134
rect 524382 92898 524414 93134
rect 523794 57454 524414 92898
rect 523794 57218 523826 57454
rect 524062 57218 524146 57454
rect 524382 57218 524414 57454
rect 523794 57134 524414 57218
rect 523794 56898 523826 57134
rect 524062 56898 524146 57134
rect 524382 56898 524414 57134
rect 523794 21454 524414 56898
rect 523794 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 524414 21454
rect 523794 21134 524414 21218
rect 523794 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 524414 21134
rect 523794 -4186 524414 20898
rect 523794 -4422 523826 -4186
rect 524062 -4422 524146 -4186
rect 524382 -4422 524414 -4186
rect 523794 -4506 524414 -4422
rect 523794 -4742 523826 -4506
rect 524062 -4742 524146 -4506
rect 524382 -4742 524414 -4506
rect 523794 -7654 524414 -4742
rect 528294 709638 528914 711590
rect 528294 709402 528326 709638
rect 528562 709402 528646 709638
rect 528882 709402 528914 709638
rect 528294 709318 528914 709402
rect 528294 709082 528326 709318
rect 528562 709082 528646 709318
rect 528882 709082 528914 709318
rect 528294 673954 528914 709082
rect 528294 673718 528326 673954
rect 528562 673718 528646 673954
rect 528882 673718 528914 673954
rect 528294 673634 528914 673718
rect 528294 673398 528326 673634
rect 528562 673398 528646 673634
rect 528882 673398 528914 673634
rect 528294 637954 528914 673398
rect 528294 637718 528326 637954
rect 528562 637718 528646 637954
rect 528882 637718 528914 637954
rect 528294 637634 528914 637718
rect 528294 637398 528326 637634
rect 528562 637398 528646 637634
rect 528882 637398 528914 637634
rect 528294 601954 528914 637398
rect 528294 601718 528326 601954
rect 528562 601718 528646 601954
rect 528882 601718 528914 601954
rect 528294 601634 528914 601718
rect 528294 601398 528326 601634
rect 528562 601398 528646 601634
rect 528882 601398 528914 601634
rect 528294 565954 528914 601398
rect 528294 565718 528326 565954
rect 528562 565718 528646 565954
rect 528882 565718 528914 565954
rect 528294 565634 528914 565718
rect 528294 565398 528326 565634
rect 528562 565398 528646 565634
rect 528882 565398 528914 565634
rect 528294 529954 528914 565398
rect 528294 529718 528326 529954
rect 528562 529718 528646 529954
rect 528882 529718 528914 529954
rect 528294 529634 528914 529718
rect 528294 529398 528326 529634
rect 528562 529398 528646 529634
rect 528882 529398 528914 529634
rect 528294 493954 528914 529398
rect 528294 493718 528326 493954
rect 528562 493718 528646 493954
rect 528882 493718 528914 493954
rect 528294 493634 528914 493718
rect 528294 493398 528326 493634
rect 528562 493398 528646 493634
rect 528882 493398 528914 493634
rect 528294 457954 528914 493398
rect 528294 457718 528326 457954
rect 528562 457718 528646 457954
rect 528882 457718 528914 457954
rect 528294 457634 528914 457718
rect 528294 457398 528326 457634
rect 528562 457398 528646 457634
rect 528882 457398 528914 457634
rect 528294 421954 528914 457398
rect 528294 421718 528326 421954
rect 528562 421718 528646 421954
rect 528882 421718 528914 421954
rect 528294 421634 528914 421718
rect 528294 421398 528326 421634
rect 528562 421398 528646 421634
rect 528882 421398 528914 421634
rect 528294 385954 528914 421398
rect 528294 385718 528326 385954
rect 528562 385718 528646 385954
rect 528882 385718 528914 385954
rect 528294 385634 528914 385718
rect 528294 385398 528326 385634
rect 528562 385398 528646 385634
rect 528882 385398 528914 385634
rect 528294 349954 528914 385398
rect 528294 349718 528326 349954
rect 528562 349718 528646 349954
rect 528882 349718 528914 349954
rect 528294 349634 528914 349718
rect 528294 349398 528326 349634
rect 528562 349398 528646 349634
rect 528882 349398 528914 349634
rect 528294 313954 528914 349398
rect 528294 313718 528326 313954
rect 528562 313718 528646 313954
rect 528882 313718 528914 313954
rect 528294 313634 528914 313718
rect 528294 313398 528326 313634
rect 528562 313398 528646 313634
rect 528882 313398 528914 313634
rect 528294 277954 528914 313398
rect 528294 277718 528326 277954
rect 528562 277718 528646 277954
rect 528882 277718 528914 277954
rect 528294 277634 528914 277718
rect 528294 277398 528326 277634
rect 528562 277398 528646 277634
rect 528882 277398 528914 277634
rect 528294 241954 528914 277398
rect 528294 241718 528326 241954
rect 528562 241718 528646 241954
rect 528882 241718 528914 241954
rect 528294 241634 528914 241718
rect 528294 241398 528326 241634
rect 528562 241398 528646 241634
rect 528882 241398 528914 241634
rect 528294 205954 528914 241398
rect 528294 205718 528326 205954
rect 528562 205718 528646 205954
rect 528882 205718 528914 205954
rect 528294 205634 528914 205718
rect 528294 205398 528326 205634
rect 528562 205398 528646 205634
rect 528882 205398 528914 205634
rect 528294 169954 528914 205398
rect 528294 169718 528326 169954
rect 528562 169718 528646 169954
rect 528882 169718 528914 169954
rect 528294 169634 528914 169718
rect 528294 169398 528326 169634
rect 528562 169398 528646 169634
rect 528882 169398 528914 169634
rect 528294 133954 528914 169398
rect 528294 133718 528326 133954
rect 528562 133718 528646 133954
rect 528882 133718 528914 133954
rect 528294 133634 528914 133718
rect 528294 133398 528326 133634
rect 528562 133398 528646 133634
rect 528882 133398 528914 133634
rect 528294 97954 528914 133398
rect 528294 97718 528326 97954
rect 528562 97718 528646 97954
rect 528882 97718 528914 97954
rect 528294 97634 528914 97718
rect 528294 97398 528326 97634
rect 528562 97398 528646 97634
rect 528882 97398 528914 97634
rect 528294 61954 528914 97398
rect 528294 61718 528326 61954
rect 528562 61718 528646 61954
rect 528882 61718 528914 61954
rect 528294 61634 528914 61718
rect 528294 61398 528326 61634
rect 528562 61398 528646 61634
rect 528882 61398 528914 61634
rect 528294 25954 528914 61398
rect 528294 25718 528326 25954
rect 528562 25718 528646 25954
rect 528882 25718 528914 25954
rect 528294 25634 528914 25718
rect 528294 25398 528326 25634
rect 528562 25398 528646 25634
rect 528882 25398 528914 25634
rect 528294 -5146 528914 25398
rect 528294 -5382 528326 -5146
rect 528562 -5382 528646 -5146
rect 528882 -5382 528914 -5146
rect 528294 -5466 528914 -5382
rect 528294 -5702 528326 -5466
rect 528562 -5702 528646 -5466
rect 528882 -5702 528914 -5466
rect 528294 -7654 528914 -5702
rect 532794 710598 533414 711590
rect 532794 710362 532826 710598
rect 533062 710362 533146 710598
rect 533382 710362 533414 710598
rect 532794 710278 533414 710362
rect 532794 710042 532826 710278
rect 533062 710042 533146 710278
rect 533382 710042 533414 710278
rect 532794 678454 533414 710042
rect 532794 678218 532826 678454
rect 533062 678218 533146 678454
rect 533382 678218 533414 678454
rect 532794 678134 533414 678218
rect 532794 677898 532826 678134
rect 533062 677898 533146 678134
rect 533382 677898 533414 678134
rect 532794 642454 533414 677898
rect 532794 642218 532826 642454
rect 533062 642218 533146 642454
rect 533382 642218 533414 642454
rect 532794 642134 533414 642218
rect 532794 641898 532826 642134
rect 533062 641898 533146 642134
rect 533382 641898 533414 642134
rect 532794 606454 533414 641898
rect 532794 606218 532826 606454
rect 533062 606218 533146 606454
rect 533382 606218 533414 606454
rect 532794 606134 533414 606218
rect 532794 605898 532826 606134
rect 533062 605898 533146 606134
rect 533382 605898 533414 606134
rect 532794 570454 533414 605898
rect 532794 570218 532826 570454
rect 533062 570218 533146 570454
rect 533382 570218 533414 570454
rect 532794 570134 533414 570218
rect 532794 569898 532826 570134
rect 533062 569898 533146 570134
rect 533382 569898 533414 570134
rect 532794 534454 533414 569898
rect 532794 534218 532826 534454
rect 533062 534218 533146 534454
rect 533382 534218 533414 534454
rect 532794 534134 533414 534218
rect 532794 533898 532826 534134
rect 533062 533898 533146 534134
rect 533382 533898 533414 534134
rect 532794 498454 533414 533898
rect 532794 498218 532826 498454
rect 533062 498218 533146 498454
rect 533382 498218 533414 498454
rect 532794 498134 533414 498218
rect 532794 497898 532826 498134
rect 533062 497898 533146 498134
rect 533382 497898 533414 498134
rect 532794 462454 533414 497898
rect 532794 462218 532826 462454
rect 533062 462218 533146 462454
rect 533382 462218 533414 462454
rect 532794 462134 533414 462218
rect 532794 461898 532826 462134
rect 533062 461898 533146 462134
rect 533382 461898 533414 462134
rect 532794 426454 533414 461898
rect 532794 426218 532826 426454
rect 533062 426218 533146 426454
rect 533382 426218 533414 426454
rect 532794 426134 533414 426218
rect 532794 425898 532826 426134
rect 533062 425898 533146 426134
rect 533382 425898 533414 426134
rect 532794 390454 533414 425898
rect 532794 390218 532826 390454
rect 533062 390218 533146 390454
rect 533382 390218 533414 390454
rect 532794 390134 533414 390218
rect 532794 389898 532826 390134
rect 533062 389898 533146 390134
rect 533382 389898 533414 390134
rect 532794 354454 533414 389898
rect 532794 354218 532826 354454
rect 533062 354218 533146 354454
rect 533382 354218 533414 354454
rect 532794 354134 533414 354218
rect 532794 353898 532826 354134
rect 533062 353898 533146 354134
rect 533382 353898 533414 354134
rect 532794 318454 533414 353898
rect 532794 318218 532826 318454
rect 533062 318218 533146 318454
rect 533382 318218 533414 318454
rect 532794 318134 533414 318218
rect 532794 317898 532826 318134
rect 533062 317898 533146 318134
rect 533382 317898 533414 318134
rect 532794 282454 533414 317898
rect 532794 282218 532826 282454
rect 533062 282218 533146 282454
rect 533382 282218 533414 282454
rect 532794 282134 533414 282218
rect 532794 281898 532826 282134
rect 533062 281898 533146 282134
rect 533382 281898 533414 282134
rect 532794 246454 533414 281898
rect 532794 246218 532826 246454
rect 533062 246218 533146 246454
rect 533382 246218 533414 246454
rect 532794 246134 533414 246218
rect 532794 245898 532826 246134
rect 533062 245898 533146 246134
rect 533382 245898 533414 246134
rect 532794 210454 533414 245898
rect 532794 210218 532826 210454
rect 533062 210218 533146 210454
rect 533382 210218 533414 210454
rect 532794 210134 533414 210218
rect 532794 209898 532826 210134
rect 533062 209898 533146 210134
rect 533382 209898 533414 210134
rect 532794 174454 533414 209898
rect 532794 174218 532826 174454
rect 533062 174218 533146 174454
rect 533382 174218 533414 174454
rect 532794 174134 533414 174218
rect 532794 173898 532826 174134
rect 533062 173898 533146 174134
rect 533382 173898 533414 174134
rect 532794 138454 533414 173898
rect 532794 138218 532826 138454
rect 533062 138218 533146 138454
rect 533382 138218 533414 138454
rect 532794 138134 533414 138218
rect 532794 137898 532826 138134
rect 533062 137898 533146 138134
rect 533382 137898 533414 138134
rect 532794 102454 533414 137898
rect 532794 102218 532826 102454
rect 533062 102218 533146 102454
rect 533382 102218 533414 102454
rect 532794 102134 533414 102218
rect 532794 101898 532826 102134
rect 533062 101898 533146 102134
rect 533382 101898 533414 102134
rect 532794 66454 533414 101898
rect 532794 66218 532826 66454
rect 533062 66218 533146 66454
rect 533382 66218 533414 66454
rect 532794 66134 533414 66218
rect 532794 65898 532826 66134
rect 533062 65898 533146 66134
rect 533382 65898 533414 66134
rect 532794 30454 533414 65898
rect 532794 30218 532826 30454
rect 533062 30218 533146 30454
rect 533382 30218 533414 30454
rect 532794 30134 533414 30218
rect 532794 29898 532826 30134
rect 533062 29898 533146 30134
rect 533382 29898 533414 30134
rect 532794 -6106 533414 29898
rect 532794 -6342 532826 -6106
rect 533062 -6342 533146 -6106
rect 533382 -6342 533414 -6106
rect 532794 -6426 533414 -6342
rect 532794 -6662 532826 -6426
rect 533062 -6662 533146 -6426
rect 533382 -6662 533414 -6426
rect 532794 -7654 533414 -6662
rect 537294 711558 537914 711590
rect 537294 711322 537326 711558
rect 537562 711322 537646 711558
rect 537882 711322 537914 711558
rect 537294 711238 537914 711322
rect 537294 711002 537326 711238
rect 537562 711002 537646 711238
rect 537882 711002 537914 711238
rect 537294 682954 537914 711002
rect 537294 682718 537326 682954
rect 537562 682718 537646 682954
rect 537882 682718 537914 682954
rect 537294 682634 537914 682718
rect 537294 682398 537326 682634
rect 537562 682398 537646 682634
rect 537882 682398 537914 682634
rect 537294 646954 537914 682398
rect 537294 646718 537326 646954
rect 537562 646718 537646 646954
rect 537882 646718 537914 646954
rect 537294 646634 537914 646718
rect 537294 646398 537326 646634
rect 537562 646398 537646 646634
rect 537882 646398 537914 646634
rect 537294 610954 537914 646398
rect 537294 610718 537326 610954
rect 537562 610718 537646 610954
rect 537882 610718 537914 610954
rect 537294 610634 537914 610718
rect 537294 610398 537326 610634
rect 537562 610398 537646 610634
rect 537882 610398 537914 610634
rect 537294 574954 537914 610398
rect 537294 574718 537326 574954
rect 537562 574718 537646 574954
rect 537882 574718 537914 574954
rect 537294 574634 537914 574718
rect 537294 574398 537326 574634
rect 537562 574398 537646 574634
rect 537882 574398 537914 574634
rect 537294 538954 537914 574398
rect 537294 538718 537326 538954
rect 537562 538718 537646 538954
rect 537882 538718 537914 538954
rect 537294 538634 537914 538718
rect 537294 538398 537326 538634
rect 537562 538398 537646 538634
rect 537882 538398 537914 538634
rect 537294 502954 537914 538398
rect 537294 502718 537326 502954
rect 537562 502718 537646 502954
rect 537882 502718 537914 502954
rect 537294 502634 537914 502718
rect 537294 502398 537326 502634
rect 537562 502398 537646 502634
rect 537882 502398 537914 502634
rect 537294 466954 537914 502398
rect 537294 466718 537326 466954
rect 537562 466718 537646 466954
rect 537882 466718 537914 466954
rect 537294 466634 537914 466718
rect 537294 466398 537326 466634
rect 537562 466398 537646 466634
rect 537882 466398 537914 466634
rect 537294 430954 537914 466398
rect 537294 430718 537326 430954
rect 537562 430718 537646 430954
rect 537882 430718 537914 430954
rect 537294 430634 537914 430718
rect 537294 430398 537326 430634
rect 537562 430398 537646 430634
rect 537882 430398 537914 430634
rect 537294 394954 537914 430398
rect 537294 394718 537326 394954
rect 537562 394718 537646 394954
rect 537882 394718 537914 394954
rect 537294 394634 537914 394718
rect 537294 394398 537326 394634
rect 537562 394398 537646 394634
rect 537882 394398 537914 394634
rect 537294 358954 537914 394398
rect 537294 358718 537326 358954
rect 537562 358718 537646 358954
rect 537882 358718 537914 358954
rect 537294 358634 537914 358718
rect 537294 358398 537326 358634
rect 537562 358398 537646 358634
rect 537882 358398 537914 358634
rect 537294 322954 537914 358398
rect 537294 322718 537326 322954
rect 537562 322718 537646 322954
rect 537882 322718 537914 322954
rect 537294 322634 537914 322718
rect 537294 322398 537326 322634
rect 537562 322398 537646 322634
rect 537882 322398 537914 322634
rect 537294 286954 537914 322398
rect 537294 286718 537326 286954
rect 537562 286718 537646 286954
rect 537882 286718 537914 286954
rect 537294 286634 537914 286718
rect 537294 286398 537326 286634
rect 537562 286398 537646 286634
rect 537882 286398 537914 286634
rect 537294 250954 537914 286398
rect 537294 250718 537326 250954
rect 537562 250718 537646 250954
rect 537882 250718 537914 250954
rect 537294 250634 537914 250718
rect 537294 250398 537326 250634
rect 537562 250398 537646 250634
rect 537882 250398 537914 250634
rect 537294 214954 537914 250398
rect 537294 214718 537326 214954
rect 537562 214718 537646 214954
rect 537882 214718 537914 214954
rect 537294 214634 537914 214718
rect 537294 214398 537326 214634
rect 537562 214398 537646 214634
rect 537882 214398 537914 214634
rect 537294 178954 537914 214398
rect 537294 178718 537326 178954
rect 537562 178718 537646 178954
rect 537882 178718 537914 178954
rect 537294 178634 537914 178718
rect 537294 178398 537326 178634
rect 537562 178398 537646 178634
rect 537882 178398 537914 178634
rect 537294 142954 537914 178398
rect 537294 142718 537326 142954
rect 537562 142718 537646 142954
rect 537882 142718 537914 142954
rect 537294 142634 537914 142718
rect 537294 142398 537326 142634
rect 537562 142398 537646 142634
rect 537882 142398 537914 142634
rect 537294 106954 537914 142398
rect 537294 106718 537326 106954
rect 537562 106718 537646 106954
rect 537882 106718 537914 106954
rect 537294 106634 537914 106718
rect 537294 106398 537326 106634
rect 537562 106398 537646 106634
rect 537882 106398 537914 106634
rect 537294 70954 537914 106398
rect 537294 70718 537326 70954
rect 537562 70718 537646 70954
rect 537882 70718 537914 70954
rect 537294 70634 537914 70718
rect 537294 70398 537326 70634
rect 537562 70398 537646 70634
rect 537882 70398 537914 70634
rect 537294 34954 537914 70398
rect 537294 34718 537326 34954
rect 537562 34718 537646 34954
rect 537882 34718 537914 34954
rect 537294 34634 537914 34718
rect 537294 34398 537326 34634
rect 537562 34398 537646 34634
rect 537882 34398 537914 34634
rect 537294 -7066 537914 34398
rect 537294 -7302 537326 -7066
rect 537562 -7302 537646 -7066
rect 537882 -7302 537914 -7066
rect 537294 -7386 537914 -7302
rect 537294 -7622 537326 -7386
rect 537562 -7622 537646 -7386
rect 537882 -7622 537914 -7386
rect 537294 -7654 537914 -7622
rect 541794 704838 542414 711590
rect 541794 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 542414 704838
rect 541794 704518 542414 704602
rect 541794 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 542414 704518
rect 541794 687454 542414 704282
rect 541794 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 542414 687454
rect 541794 687134 542414 687218
rect 541794 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 542414 687134
rect 541794 651454 542414 686898
rect 541794 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 542414 651454
rect 541794 651134 542414 651218
rect 541794 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 542414 651134
rect 541794 615454 542414 650898
rect 541794 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 542414 615454
rect 541794 615134 542414 615218
rect 541794 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 542414 615134
rect 541794 579454 542414 614898
rect 541794 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 542414 579454
rect 541794 579134 542414 579218
rect 541794 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 542414 579134
rect 541794 543454 542414 578898
rect 541794 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 542414 543454
rect 541794 543134 542414 543218
rect 541794 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 542414 543134
rect 541794 507454 542414 542898
rect 541794 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 542414 507454
rect 541794 507134 542414 507218
rect 541794 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 542414 507134
rect 541794 471454 542414 506898
rect 541794 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 542414 471454
rect 541794 471134 542414 471218
rect 541794 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 542414 471134
rect 541794 435454 542414 470898
rect 541794 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 542414 435454
rect 541794 435134 542414 435218
rect 541794 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 542414 435134
rect 541794 399454 542414 434898
rect 541794 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 542414 399454
rect 541794 399134 542414 399218
rect 541794 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 542414 399134
rect 541794 363454 542414 398898
rect 541794 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 542414 363454
rect 541794 363134 542414 363218
rect 541794 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 542414 363134
rect 541794 327454 542414 362898
rect 541794 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 542414 327454
rect 541794 327134 542414 327218
rect 541794 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 542414 327134
rect 541794 291454 542414 326898
rect 541794 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 542414 291454
rect 541794 291134 542414 291218
rect 541794 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 542414 291134
rect 541794 255454 542414 290898
rect 541794 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 542414 255454
rect 541794 255134 542414 255218
rect 541794 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 542414 255134
rect 541794 219454 542414 254898
rect 541794 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 542414 219454
rect 541794 219134 542414 219218
rect 541794 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 542414 219134
rect 541794 183454 542414 218898
rect 541794 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 542414 183454
rect 541794 183134 542414 183218
rect 541794 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 542414 183134
rect 541794 147454 542414 182898
rect 541794 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 542414 147454
rect 541794 147134 542414 147218
rect 541794 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 542414 147134
rect 541794 111454 542414 146898
rect 541794 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 542414 111454
rect 541794 111134 542414 111218
rect 541794 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 542414 111134
rect 541794 75454 542414 110898
rect 541794 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 542414 75454
rect 541794 75134 542414 75218
rect 541794 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 542414 75134
rect 541794 39454 542414 74898
rect 541794 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 542414 39454
rect 541794 39134 542414 39218
rect 541794 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 542414 39134
rect 541794 3454 542414 38898
rect 541794 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 542414 3454
rect 541794 3134 542414 3218
rect 541794 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 542414 3134
rect 541794 -346 542414 2898
rect 541794 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 542414 -346
rect 541794 -666 542414 -582
rect 541794 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 542414 -666
rect 541794 -7654 542414 -902
rect 546294 705798 546914 711590
rect 546294 705562 546326 705798
rect 546562 705562 546646 705798
rect 546882 705562 546914 705798
rect 546294 705478 546914 705562
rect 546294 705242 546326 705478
rect 546562 705242 546646 705478
rect 546882 705242 546914 705478
rect 546294 691954 546914 705242
rect 546294 691718 546326 691954
rect 546562 691718 546646 691954
rect 546882 691718 546914 691954
rect 546294 691634 546914 691718
rect 546294 691398 546326 691634
rect 546562 691398 546646 691634
rect 546882 691398 546914 691634
rect 546294 655954 546914 691398
rect 546294 655718 546326 655954
rect 546562 655718 546646 655954
rect 546882 655718 546914 655954
rect 546294 655634 546914 655718
rect 546294 655398 546326 655634
rect 546562 655398 546646 655634
rect 546882 655398 546914 655634
rect 546294 619954 546914 655398
rect 546294 619718 546326 619954
rect 546562 619718 546646 619954
rect 546882 619718 546914 619954
rect 546294 619634 546914 619718
rect 546294 619398 546326 619634
rect 546562 619398 546646 619634
rect 546882 619398 546914 619634
rect 546294 583954 546914 619398
rect 546294 583718 546326 583954
rect 546562 583718 546646 583954
rect 546882 583718 546914 583954
rect 546294 583634 546914 583718
rect 546294 583398 546326 583634
rect 546562 583398 546646 583634
rect 546882 583398 546914 583634
rect 546294 547954 546914 583398
rect 546294 547718 546326 547954
rect 546562 547718 546646 547954
rect 546882 547718 546914 547954
rect 546294 547634 546914 547718
rect 546294 547398 546326 547634
rect 546562 547398 546646 547634
rect 546882 547398 546914 547634
rect 546294 511954 546914 547398
rect 546294 511718 546326 511954
rect 546562 511718 546646 511954
rect 546882 511718 546914 511954
rect 546294 511634 546914 511718
rect 546294 511398 546326 511634
rect 546562 511398 546646 511634
rect 546882 511398 546914 511634
rect 546294 475954 546914 511398
rect 546294 475718 546326 475954
rect 546562 475718 546646 475954
rect 546882 475718 546914 475954
rect 546294 475634 546914 475718
rect 546294 475398 546326 475634
rect 546562 475398 546646 475634
rect 546882 475398 546914 475634
rect 546294 439954 546914 475398
rect 546294 439718 546326 439954
rect 546562 439718 546646 439954
rect 546882 439718 546914 439954
rect 546294 439634 546914 439718
rect 546294 439398 546326 439634
rect 546562 439398 546646 439634
rect 546882 439398 546914 439634
rect 546294 403954 546914 439398
rect 546294 403718 546326 403954
rect 546562 403718 546646 403954
rect 546882 403718 546914 403954
rect 546294 403634 546914 403718
rect 546294 403398 546326 403634
rect 546562 403398 546646 403634
rect 546882 403398 546914 403634
rect 546294 367954 546914 403398
rect 546294 367718 546326 367954
rect 546562 367718 546646 367954
rect 546882 367718 546914 367954
rect 546294 367634 546914 367718
rect 546294 367398 546326 367634
rect 546562 367398 546646 367634
rect 546882 367398 546914 367634
rect 546294 331954 546914 367398
rect 546294 331718 546326 331954
rect 546562 331718 546646 331954
rect 546882 331718 546914 331954
rect 546294 331634 546914 331718
rect 546294 331398 546326 331634
rect 546562 331398 546646 331634
rect 546882 331398 546914 331634
rect 546294 295954 546914 331398
rect 546294 295718 546326 295954
rect 546562 295718 546646 295954
rect 546882 295718 546914 295954
rect 546294 295634 546914 295718
rect 546294 295398 546326 295634
rect 546562 295398 546646 295634
rect 546882 295398 546914 295634
rect 546294 259954 546914 295398
rect 546294 259718 546326 259954
rect 546562 259718 546646 259954
rect 546882 259718 546914 259954
rect 546294 259634 546914 259718
rect 546294 259398 546326 259634
rect 546562 259398 546646 259634
rect 546882 259398 546914 259634
rect 546294 223954 546914 259398
rect 546294 223718 546326 223954
rect 546562 223718 546646 223954
rect 546882 223718 546914 223954
rect 546294 223634 546914 223718
rect 546294 223398 546326 223634
rect 546562 223398 546646 223634
rect 546882 223398 546914 223634
rect 546294 187954 546914 223398
rect 546294 187718 546326 187954
rect 546562 187718 546646 187954
rect 546882 187718 546914 187954
rect 546294 187634 546914 187718
rect 546294 187398 546326 187634
rect 546562 187398 546646 187634
rect 546882 187398 546914 187634
rect 546294 151954 546914 187398
rect 546294 151718 546326 151954
rect 546562 151718 546646 151954
rect 546882 151718 546914 151954
rect 546294 151634 546914 151718
rect 546294 151398 546326 151634
rect 546562 151398 546646 151634
rect 546882 151398 546914 151634
rect 546294 115954 546914 151398
rect 546294 115718 546326 115954
rect 546562 115718 546646 115954
rect 546882 115718 546914 115954
rect 546294 115634 546914 115718
rect 546294 115398 546326 115634
rect 546562 115398 546646 115634
rect 546882 115398 546914 115634
rect 546294 79954 546914 115398
rect 546294 79718 546326 79954
rect 546562 79718 546646 79954
rect 546882 79718 546914 79954
rect 546294 79634 546914 79718
rect 546294 79398 546326 79634
rect 546562 79398 546646 79634
rect 546882 79398 546914 79634
rect 546294 43954 546914 79398
rect 546294 43718 546326 43954
rect 546562 43718 546646 43954
rect 546882 43718 546914 43954
rect 546294 43634 546914 43718
rect 546294 43398 546326 43634
rect 546562 43398 546646 43634
rect 546882 43398 546914 43634
rect 546294 7954 546914 43398
rect 546294 7718 546326 7954
rect 546562 7718 546646 7954
rect 546882 7718 546914 7954
rect 546294 7634 546914 7718
rect 546294 7398 546326 7634
rect 546562 7398 546646 7634
rect 546882 7398 546914 7634
rect 546294 -1306 546914 7398
rect 546294 -1542 546326 -1306
rect 546562 -1542 546646 -1306
rect 546882 -1542 546914 -1306
rect 546294 -1626 546914 -1542
rect 546294 -1862 546326 -1626
rect 546562 -1862 546646 -1626
rect 546882 -1862 546914 -1626
rect 546294 -7654 546914 -1862
rect 550794 706758 551414 711590
rect 550794 706522 550826 706758
rect 551062 706522 551146 706758
rect 551382 706522 551414 706758
rect 550794 706438 551414 706522
rect 550794 706202 550826 706438
rect 551062 706202 551146 706438
rect 551382 706202 551414 706438
rect 550794 696454 551414 706202
rect 550794 696218 550826 696454
rect 551062 696218 551146 696454
rect 551382 696218 551414 696454
rect 550794 696134 551414 696218
rect 550794 695898 550826 696134
rect 551062 695898 551146 696134
rect 551382 695898 551414 696134
rect 550794 660454 551414 695898
rect 550794 660218 550826 660454
rect 551062 660218 551146 660454
rect 551382 660218 551414 660454
rect 550794 660134 551414 660218
rect 550794 659898 550826 660134
rect 551062 659898 551146 660134
rect 551382 659898 551414 660134
rect 550794 624454 551414 659898
rect 550794 624218 550826 624454
rect 551062 624218 551146 624454
rect 551382 624218 551414 624454
rect 550794 624134 551414 624218
rect 550794 623898 550826 624134
rect 551062 623898 551146 624134
rect 551382 623898 551414 624134
rect 550794 588454 551414 623898
rect 550794 588218 550826 588454
rect 551062 588218 551146 588454
rect 551382 588218 551414 588454
rect 550794 588134 551414 588218
rect 550794 587898 550826 588134
rect 551062 587898 551146 588134
rect 551382 587898 551414 588134
rect 550794 552454 551414 587898
rect 550794 552218 550826 552454
rect 551062 552218 551146 552454
rect 551382 552218 551414 552454
rect 550794 552134 551414 552218
rect 550794 551898 550826 552134
rect 551062 551898 551146 552134
rect 551382 551898 551414 552134
rect 550794 516454 551414 551898
rect 550794 516218 550826 516454
rect 551062 516218 551146 516454
rect 551382 516218 551414 516454
rect 550794 516134 551414 516218
rect 550794 515898 550826 516134
rect 551062 515898 551146 516134
rect 551382 515898 551414 516134
rect 550794 480454 551414 515898
rect 550794 480218 550826 480454
rect 551062 480218 551146 480454
rect 551382 480218 551414 480454
rect 550794 480134 551414 480218
rect 550794 479898 550826 480134
rect 551062 479898 551146 480134
rect 551382 479898 551414 480134
rect 550794 444454 551414 479898
rect 550794 444218 550826 444454
rect 551062 444218 551146 444454
rect 551382 444218 551414 444454
rect 550794 444134 551414 444218
rect 550794 443898 550826 444134
rect 551062 443898 551146 444134
rect 551382 443898 551414 444134
rect 550794 408454 551414 443898
rect 550794 408218 550826 408454
rect 551062 408218 551146 408454
rect 551382 408218 551414 408454
rect 550794 408134 551414 408218
rect 550794 407898 550826 408134
rect 551062 407898 551146 408134
rect 551382 407898 551414 408134
rect 550794 372454 551414 407898
rect 550794 372218 550826 372454
rect 551062 372218 551146 372454
rect 551382 372218 551414 372454
rect 550794 372134 551414 372218
rect 550794 371898 550826 372134
rect 551062 371898 551146 372134
rect 551382 371898 551414 372134
rect 550794 336454 551414 371898
rect 550794 336218 550826 336454
rect 551062 336218 551146 336454
rect 551382 336218 551414 336454
rect 550794 336134 551414 336218
rect 550794 335898 550826 336134
rect 551062 335898 551146 336134
rect 551382 335898 551414 336134
rect 550794 300454 551414 335898
rect 550794 300218 550826 300454
rect 551062 300218 551146 300454
rect 551382 300218 551414 300454
rect 550794 300134 551414 300218
rect 550794 299898 550826 300134
rect 551062 299898 551146 300134
rect 551382 299898 551414 300134
rect 550794 264454 551414 299898
rect 550794 264218 550826 264454
rect 551062 264218 551146 264454
rect 551382 264218 551414 264454
rect 550794 264134 551414 264218
rect 550794 263898 550826 264134
rect 551062 263898 551146 264134
rect 551382 263898 551414 264134
rect 550794 228454 551414 263898
rect 550794 228218 550826 228454
rect 551062 228218 551146 228454
rect 551382 228218 551414 228454
rect 550794 228134 551414 228218
rect 550794 227898 550826 228134
rect 551062 227898 551146 228134
rect 551382 227898 551414 228134
rect 550794 192454 551414 227898
rect 550794 192218 550826 192454
rect 551062 192218 551146 192454
rect 551382 192218 551414 192454
rect 550794 192134 551414 192218
rect 550794 191898 550826 192134
rect 551062 191898 551146 192134
rect 551382 191898 551414 192134
rect 550794 156454 551414 191898
rect 550794 156218 550826 156454
rect 551062 156218 551146 156454
rect 551382 156218 551414 156454
rect 550794 156134 551414 156218
rect 550794 155898 550826 156134
rect 551062 155898 551146 156134
rect 551382 155898 551414 156134
rect 550794 120454 551414 155898
rect 550794 120218 550826 120454
rect 551062 120218 551146 120454
rect 551382 120218 551414 120454
rect 550794 120134 551414 120218
rect 550794 119898 550826 120134
rect 551062 119898 551146 120134
rect 551382 119898 551414 120134
rect 550794 84454 551414 119898
rect 550794 84218 550826 84454
rect 551062 84218 551146 84454
rect 551382 84218 551414 84454
rect 550794 84134 551414 84218
rect 550794 83898 550826 84134
rect 551062 83898 551146 84134
rect 551382 83898 551414 84134
rect 550794 48454 551414 83898
rect 550794 48218 550826 48454
rect 551062 48218 551146 48454
rect 551382 48218 551414 48454
rect 550794 48134 551414 48218
rect 550794 47898 550826 48134
rect 551062 47898 551146 48134
rect 551382 47898 551414 48134
rect 550794 12454 551414 47898
rect 550794 12218 550826 12454
rect 551062 12218 551146 12454
rect 551382 12218 551414 12454
rect 550794 12134 551414 12218
rect 550794 11898 550826 12134
rect 551062 11898 551146 12134
rect 551382 11898 551414 12134
rect 550794 -2266 551414 11898
rect 550794 -2502 550826 -2266
rect 551062 -2502 551146 -2266
rect 551382 -2502 551414 -2266
rect 550794 -2586 551414 -2502
rect 550794 -2822 550826 -2586
rect 551062 -2822 551146 -2586
rect 551382 -2822 551414 -2586
rect 550794 -7654 551414 -2822
rect 555294 707718 555914 711590
rect 555294 707482 555326 707718
rect 555562 707482 555646 707718
rect 555882 707482 555914 707718
rect 555294 707398 555914 707482
rect 555294 707162 555326 707398
rect 555562 707162 555646 707398
rect 555882 707162 555914 707398
rect 555294 700954 555914 707162
rect 555294 700718 555326 700954
rect 555562 700718 555646 700954
rect 555882 700718 555914 700954
rect 555294 700634 555914 700718
rect 555294 700398 555326 700634
rect 555562 700398 555646 700634
rect 555882 700398 555914 700634
rect 555294 664954 555914 700398
rect 555294 664718 555326 664954
rect 555562 664718 555646 664954
rect 555882 664718 555914 664954
rect 555294 664634 555914 664718
rect 555294 664398 555326 664634
rect 555562 664398 555646 664634
rect 555882 664398 555914 664634
rect 555294 628954 555914 664398
rect 555294 628718 555326 628954
rect 555562 628718 555646 628954
rect 555882 628718 555914 628954
rect 555294 628634 555914 628718
rect 555294 628398 555326 628634
rect 555562 628398 555646 628634
rect 555882 628398 555914 628634
rect 555294 592954 555914 628398
rect 555294 592718 555326 592954
rect 555562 592718 555646 592954
rect 555882 592718 555914 592954
rect 555294 592634 555914 592718
rect 555294 592398 555326 592634
rect 555562 592398 555646 592634
rect 555882 592398 555914 592634
rect 555294 556954 555914 592398
rect 555294 556718 555326 556954
rect 555562 556718 555646 556954
rect 555882 556718 555914 556954
rect 555294 556634 555914 556718
rect 555294 556398 555326 556634
rect 555562 556398 555646 556634
rect 555882 556398 555914 556634
rect 555294 520954 555914 556398
rect 555294 520718 555326 520954
rect 555562 520718 555646 520954
rect 555882 520718 555914 520954
rect 555294 520634 555914 520718
rect 555294 520398 555326 520634
rect 555562 520398 555646 520634
rect 555882 520398 555914 520634
rect 555294 484954 555914 520398
rect 555294 484718 555326 484954
rect 555562 484718 555646 484954
rect 555882 484718 555914 484954
rect 555294 484634 555914 484718
rect 555294 484398 555326 484634
rect 555562 484398 555646 484634
rect 555882 484398 555914 484634
rect 555294 448954 555914 484398
rect 555294 448718 555326 448954
rect 555562 448718 555646 448954
rect 555882 448718 555914 448954
rect 555294 448634 555914 448718
rect 555294 448398 555326 448634
rect 555562 448398 555646 448634
rect 555882 448398 555914 448634
rect 555294 412954 555914 448398
rect 555294 412718 555326 412954
rect 555562 412718 555646 412954
rect 555882 412718 555914 412954
rect 555294 412634 555914 412718
rect 555294 412398 555326 412634
rect 555562 412398 555646 412634
rect 555882 412398 555914 412634
rect 555294 376954 555914 412398
rect 555294 376718 555326 376954
rect 555562 376718 555646 376954
rect 555882 376718 555914 376954
rect 555294 376634 555914 376718
rect 555294 376398 555326 376634
rect 555562 376398 555646 376634
rect 555882 376398 555914 376634
rect 555294 340954 555914 376398
rect 555294 340718 555326 340954
rect 555562 340718 555646 340954
rect 555882 340718 555914 340954
rect 555294 340634 555914 340718
rect 555294 340398 555326 340634
rect 555562 340398 555646 340634
rect 555882 340398 555914 340634
rect 555294 304954 555914 340398
rect 555294 304718 555326 304954
rect 555562 304718 555646 304954
rect 555882 304718 555914 304954
rect 555294 304634 555914 304718
rect 555294 304398 555326 304634
rect 555562 304398 555646 304634
rect 555882 304398 555914 304634
rect 555294 268954 555914 304398
rect 555294 268718 555326 268954
rect 555562 268718 555646 268954
rect 555882 268718 555914 268954
rect 555294 268634 555914 268718
rect 555294 268398 555326 268634
rect 555562 268398 555646 268634
rect 555882 268398 555914 268634
rect 555294 232954 555914 268398
rect 555294 232718 555326 232954
rect 555562 232718 555646 232954
rect 555882 232718 555914 232954
rect 555294 232634 555914 232718
rect 555294 232398 555326 232634
rect 555562 232398 555646 232634
rect 555882 232398 555914 232634
rect 555294 196954 555914 232398
rect 555294 196718 555326 196954
rect 555562 196718 555646 196954
rect 555882 196718 555914 196954
rect 555294 196634 555914 196718
rect 555294 196398 555326 196634
rect 555562 196398 555646 196634
rect 555882 196398 555914 196634
rect 555294 160954 555914 196398
rect 555294 160718 555326 160954
rect 555562 160718 555646 160954
rect 555882 160718 555914 160954
rect 555294 160634 555914 160718
rect 555294 160398 555326 160634
rect 555562 160398 555646 160634
rect 555882 160398 555914 160634
rect 555294 124954 555914 160398
rect 555294 124718 555326 124954
rect 555562 124718 555646 124954
rect 555882 124718 555914 124954
rect 555294 124634 555914 124718
rect 555294 124398 555326 124634
rect 555562 124398 555646 124634
rect 555882 124398 555914 124634
rect 555294 88954 555914 124398
rect 555294 88718 555326 88954
rect 555562 88718 555646 88954
rect 555882 88718 555914 88954
rect 555294 88634 555914 88718
rect 555294 88398 555326 88634
rect 555562 88398 555646 88634
rect 555882 88398 555914 88634
rect 555294 52954 555914 88398
rect 555294 52718 555326 52954
rect 555562 52718 555646 52954
rect 555882 52718 555914 52954
rect 555294 52634 555914 52718
rect 555294 52398 555326 52634
rect 555562 52398 555646 52634
rect 555882 52398 555914 52634
rect 555294 16954 555914 52398
rect 555294 16718 555326 16954
rect 555562 16718 555646 16954
rect 555882 16718 555914 16954
rect 555294 16634 555914 16718
rect 555294 16398 555326 16634
rect 555562 16398 555646 16634
rect 555882 16398 555914 16634
rect 555294 -3226 555914 16398
rect 555294 -3462 555326 -3226
rect 555562 -3462 555646 -3226
rect 555882 -3462 555914 -3226
rect 555294 -3546 555914 -3462
rect 555294 -3782 555326 -3546
rect 555562 -3782 555646 -3546
rect 555882 -3782 555914 -3546
rect 555294 -7654 555914 -3782
rect 559794 708678 560414 711590
rect 559794 708442 559826 708678
rect 560062 708442 560146 708678
rect 560382 708442 560414 708678
rect 559794 708358 560414 708442
rect 559794 708122 559826 708358
rect 560062 708122 560146 708358
rect 560382 708122 560414 708358
rect 559794 669454 560414 708122
rect 559794 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 560414 669454
rect 559794 669134 560414 669218
rect 559794 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 560414 669134
rect 559794 633454 560414 668898
rect 559794 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 560414 633454
rect 559794 633134 560414 633218
rect 559794 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 560414 633134
rect 559794 597454 560414 632898
rect 559794 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 560414 597454
rect 559794 597134 560414 597218
rect 559794 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 560414 597134
rect 559794 561454 560414 596898
rect 559794 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 560414 561454
rect 559794 561134 560414 561218
rect 559794 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 560414 561134
rect 559794 525454 560414 560898
rect 559794 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 560414 525454
rect 559794 525134 560414 525218
rect 559794 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 560414 525134
rect 559794 489454 560414 524898
rect 559794 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 560414 489454
rect 559794 489134 560414 489218
rect 559794 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 560414 489134
rect 559794 453454 560414 488898
rect 559794 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 560414 453454
rect 559794 453134 560414 453218
rect 559794 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 560414 453134
rect 559794 417454 560414 452898
rect 559794 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 560414 417454
rect 559794 417134 560414 417218
rect 559794 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 560414 417134
rect 559794 381454 560414 416898
rect 559794 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 560414 381454
rect 559794 381134 560414 381218
rect 559794 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 560414 381134
rect 559794 345454 560414 380898
rect 559794 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 560414 345454
rect 559794 345134 560414 345218
rect 559794 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 560414 345134
rect 559794 309454 560414 344898
rect 559794 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 560414 309454
rect 559794 309134 560414 309218
rect 559794 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 560414 309134
rect 559794 273454 560414 308898
rect 559794 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 560414 273454
rect 559794 273134 560414 273218
rect 559794 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 560414 273134
rect 559794 237454 560414 272898
rect 559794 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 560414 237454
rect 559794 237134 560414 237218
rect 559794 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 560414 237134
rect 559794 201454 560414 236898
rect 559794 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 560414 201454
rect 559794 201134 560414 201218
rect 559794 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 560414 201134
rect 559794 165454 560414 200898
rect 559794 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 560414 165454
rect 559794 165134 560414 165218
rect 559794 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 560414 165134
rect 559794 129454 560414 164898
rect 559794 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 560414 129454
rect 559794 129134 560414 129218
rect 559794 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 560414 129134
rect 559794 93454 560414 128898
rect 559794 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 560414 93454
rect 559794 93134 560414 93218
rect 559794 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 560414 93134
rect 559794 57454 560414 92898
rect 559794 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 560414 57454
rect 559794 57134 560414 57218
rect 559794 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 560414 57134
rect 559794 21454 560414 56898
rect 559794 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 560414 21454
rect 559794 21134 560414 21218
rect 559794 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 560414 21134
rect 559794 -4186 560414 20898
rect 559794 -4422 559826 -4186
rect 560062 -4422 560146 -4186
rect 560382 -4422 560414 -4186
rect 559794 -4506 560414 -4422
rect 559794 -4742 559826 -4506
rect 560062 -4742 560146 -4506
rect 560382 -4742 560414 -4506
rect 559794 -7654 560414 -4742
rect 564294 709638 564914 711590
rect 564294 709402 564326 709638
rect 564562 709402 564646 709638
rect 564882 709402 564914 709638
rect 564294 709318 564914 709402
rect 564294 709082 564326 709318
rect 564562 709082 564646 709318
rect 564882 709082 564914 709318
rect 564294 673954 564914 709082
rect 564294 673718 564326 673954
rect 564562 673718 564646 673954
rect 564882 673718 564914 673954
rect 564294 673634 564914 673718
rect 564294 673398 564326 673634
rect 564562 673398 564646 673634
rect 564882 673398 564914 673634
rect 564294 637954 564914 673398
rect 564294 637718 564326 637954
rect 564562 637718 564646 637954
rect 564882 637718 564914 637954
rect 564294 637634 564914 637718
rect 564294 637398 564326 637634
rect 564562 637398 564646 637634
rect 564882 637398 564914 637634
rect 564294 601954 564914 637398
rect 564294 601718 564326 601954
rect 564562 601718 564646 601954
rect 564882 601718 564914 601954
rect 564294 601634 564914 601718
rect 564294 601398 564326 601634
rect 564562 601398 564646 601634
rect 564882 601398 564914 601634
rect 564294 565954 564914 601398
rect 564294 565718 564326 565954
rect 564562 565718 564646 565954
rect 564882 565718 564914 565954
rect 564294 565634 564914 565718
rect 564294 565398 564326 565634
rect 564562 565398 564646 565634
rect 564882 565398 564914 565634
rect 564294 529954 564914 565398
rect 564294 529718 564326 529954
rect 564562 529718 564646 529954
rect 564882 529718 564914 529954
rect 564294 529634 564914 529718
rect 564294 529398 564326 529634
rect 564562 529398 564646 529634
rect 564882 529398 564914 529634
rect 564294 493954 564914 529398
rect 564294 493718 564326 493954
rect 564562 493718 564646 493954
rect 564882 493718 564914 493954
rect 564294 493634 564914 493718
rect 564294 493398 564326 493634
rect 564562 493398 564646 493634
rect 564882 493398 564914 493634
rect 564294 457954 564914 493398
rect 564294 457718 564326 457954
rect 564562 457718 564646 457954
rect 564882 457718 564914 457954
rect 564294 457634 564914 457718
rect 564294 457398 564326 457634
rect 564562 457398 564646 457634
rect 564882 457398 564914 457634
rect 564294 421954 564914 457398
rect 564294 421718 564326 421954
rect 564562 421718 564646 421954
rect 564882 421718 564914 421954
rect 564294 421634 564914 421718
rect 564294 421398 564326 421634
rect 564562 421398 564646 421634
rect 564882 421398 564914 421634
rect 564294 385954 564914 421398
rect 564294 385718 564326 385954
rect 564562 385718 564646 385954
rect 564882 385718 564914 385954
rect 564294 385634 564914 385718
rect 564294 385398 564326 385634
rect 564562 385398 564646 385634
rect 564882 385398 564914 385634
rect 564294 349954 564914 385398
rect 564294 349718 564326 349954
rect 564562 349718 564646 349954
rect 564882 349718 564914 349954
rect 564294 349634 564914 349718
rect 564294 349398 564326 349634
rect 564562 349398 564646 349634
rect 564882 349398 564914 349634
rect 564294 313954 564914 349398
rect 564294 313718 564326 313954
rect 564562 313718 564646 313954
rect 564882 313718 564914 313954
rect 564294 313634 564914 313718
rect 564294 313398 564326 313634
rect 564562 313398 564646 313634
rect 564882 313398 564914 313634
rect 564294 277954 564914 313398
rect 564294 277718 564326 277954
rect 564562 277718 564646 277954
rect 564882 277718 564914 277954
rect 564294 277634 564914 277718
rect 564294 277398 564326 277634
rect 564562 277398 564646 277634
rect 564882 277398 564914 277634
rect 564294 241954 564914 277398
rect 564294 241718 564326 241954
rect 564562 241718 564646 241954
rect 564882 241718 564914 241954
rect 564294 241634 564914 241718
rect 564294 241398 564326 241634
rect 564562 241398 564646 241634
rect 564882 241398 564914 241634
rect 564294 205954 564914 241398
rect 564294 205718 564326 205954
rect 564562 205718 564646 205954
rect 564882 205718 564914 205954
rect 564294 205634 564914 205718
rect 564294 205398 564326 205634
rect 564562 205398 564646 205634
rect 564882 205398 564914 205634
rect 564294 169954 564914 205398
rect 564294 169718 564326 169954
rect 564562 169718 564646 169954
rect 564882 169718 564914 169954
rect 564294 169634 564914 169718
rect 564294 169398 564326 169634
rect 564562 169398 564646 169634
rect 564882 169398 564914 169634
rect 564294 133954 564914 169398
rect 564294 133718 564326 133954
rect 564562 133718 564646 133954
rect 564882 133718 564914 133954
rect 564294 133634 564914 133718
rect 564294 133398 564326 133634
rect 564562 133398 564646 133634
rect 564882 133398 564914 133634
rect 564294 97954 564914 133398
rect 564294 97718 564326 97954
rect 564562 97718 564646 97954
rect 564882 97718 564914 97954
rect 564294 97634 564914 97718
rect 564294 97398 564326 97634
rect 564562 97398 564646 97634
rect 564882 97398 564914 97634
rect 564294 61954 564914 97398
rect 564294 61718 564326 61954
rect 564562 61718 564646 61954
rect 564882 61718 564914 61954
rect 564294 61634 564914 61718
rect 564294 61398 564326 61634
rect 564562 61398 564646 61634
rect 564882 61398 564914 61634
rect 564294 25954 564914 61398
rect 564294 25718 564326 25954
rect 564562 25718 564646 25954
rect 564882 25718 564914 25954
rect 564294 25634 564914 25718
rect 564294 25398 564326 25634
rect 564562 25398 564646 25634
rect 564882 25398 564914 25634
rect 564294 -5146 564914 25398
rect 564294 -5382 564326 -5146
rect 564562 -5382 564646 -5146
rect 564882 -5382 564914 -5146
rect 564294 -5466 564914 -5382
rect 564294 -5702 564326 -5466
rect 564562 -5702 564646 -5466
rect 564882 -5702 564914 -5466
rect 564294 -7654 564914 -5702
rect 568794 710598 569414 711590
rect 568794 710362 568826 710598
rect 569062 710362 569146 710598
rect 569382 710362 569414 710598
rect 568794 710278 569414 710362
rect 568794 710042 568826 710278
rect 569062 710042 569146 710278
rect 569382 710042 569414 710278
rect 568794 678454 569414 710042
rect 568794 678218 568826 678454
rect 569062 678218 569146 678454
rect 569382 678218 569414 678454
rect 568794 678134 569414 678218
rect 568794 677898 568826 678134
rect 569062 677898 569146 678134
rect 569382 677898 569414 678134
rect 568794 642454 569414 677898
rect 568794 642218 568826 642454
rect 569062 642218 569146 642454
rect 569382 642218 569414 642454
rect 568794 642134 569414 642218
rect 568794 641898 568826 642134
rect 569062 641898 569146 642134
rect 569382 641898 569414 642134
rect 568794 606454 569414 641898
rect 568794 606218 568826 606454
rect 569062 606218 569146 606454
rect 569382 606218 569414 606454
rect 568794 606134 569414 606218
rect 568794 605898 568826 606134
rect 569062 605898 569146 606134
rect 569382 605898 569414 606134
rect 568794 570454 569414 605898
rect 568794 570218 568826 570454
rect 569062 570218 569146 570454
rect 569382 570218 569414 570454
rect 568794 570134 569414 570218
rect 568794 569898 568826 570134
rect 569062 569898 569146 570134
rect 569382 569898 569414 570134
rect 568794 534454 569414 569898
rect 568794 534218 568826 534454
rect 569062 534218 569146 534454
rect 569382 534218 569414 534454
rect 568794 534134 569414 534218
rect 568794 533898 568826 534134
rect 569062 533898 569146 534134
rect 569382 533898 569414 534134
rect 568794 498454 569414 533898
rect 568794 498218 568826 498454
rect 569062 498218 569146 498454
rect 569382 498218 569414 498454
rect 568794 498134 569414 498218
rect 568794 497898 568826 498134
rect 569062 497898 569146 498134
rect 569382 497898 569414 498134
rect 568794 462454 569414 497898
rect 568794 462218 568826 462454
rect 569062 462218 569146 462454
rect 569382 462218 569414 462454
rect 568794 462134 569414 462218
rect 568794 461898 568826 462134
rect 569062 461898 569146 462134
rect 569382 461898 569414 462134
rect 568794 426454 569414 461898
rect 568794 426218 568826 426454
rect 569062 426218 569146 426454
rect 569382 426218 569414 426454
rect 568794 426134 569414 426218
rect 568794 425898 568826 426134
rect 569062 425898 569146 426134
rect 569382 425898 569414 426134
rect 568794 390454 569414 425898
rect 568794 390218 568826 390454
rect 569062 390218 569146 390454
rect 569382 390218 569414 390454
rect 568794 390134 569414 390218
rect 568794 389898 568826 390134
rect 569062 389898 569146 390134
rect 569382 389898 569414 390134
rect 568794 354454 569414 389898
rect 568794 354218 568826 354454
rect 569062 354218 569146 354454
rect 569382 354218 569414 354454
rect 568794 354134 569414 354218
rect 568794 353898 568826 354134
rect 569062 353898 569146 354134
rect 569382 353898 569414 354134
rect 568794 318454 569414 353898
rect 568794 318218 568826 318454
rect 569062 318218 569146 318454
rect 569382 318218 569414 318454
rect 568794 318134 569414 318218
rect 568794 317898 568826 318134
rect 569062 317898 569146 318134
rect 569382 317898 569414 318134
rect 568794 282454 569414 317898
rect 568794 282218 568826 282454
rect 569062 282218 569146 282454
rect 569382 282218 569414 282454
rect 568794 282134 569414 282218
rect 568794 281898 568826 282134
rect 569062 281898 569146 282134
rect 569382 281898 569414 282134
rect 568794 246454 569414 281898
rect 568794 246218 568826 246454
rect 569062 246218 569146 246454
rect 569382 246218 569414 246454
rect 568794 246134 569414 246218
rect 568794 245898 568826 246134
rect 569062 245898 569146 246134
rect 569382 245898 569414 246134
rect 568794 210454 569414 245898
rect 568794 210218 568826 210454
rect 569062 210218 569146 210454
rect 569382 210218 569414 210454
rect 568794 210134 569414 210218
rect 568794 209898 568826 210134
rect 569062 209898 569146 210134
rect 569382 209898 569414 210134
rect 568794 174454 569414 209898
rect 568794 174218 568826 174454
rect 569062 174218 569146 174454
rect 569382 174218 569414 174454
rect 568794 174134 569414 174218
rect 568794 173898 568826 174134
rect 569062 173898 569146 174134
rect 569382 173898 569414 174134
rect 568794 138454 569414 173898
rect 568794 138218 568826 138454
rect 569062 138218 569146 138454
rect 569382 138218 569414 138454
rect 568794 138134 569414 138218
rect 568794 137898 568826 138134
rect 569062 137898 569146 138134
rect 569382 137898 569414 138134
rect 568794 102454 569414 137898
rect 568794 102218 568826 102454
rect 569062 102218 569146 102454
rect 569382 102218 569414 102454
rect 568794 102134 569414 102218
rect 568794 101898 568826 102134
rect 569062 101898 569146 102134
rect 569382 101898 569414 102134
rect 568794 66454 569414 101898
rect 568794 66218 568826 66454
rect 569062 66218 569146 66454
rect 569382 66218 569414 66454
rect 568794 66134 569414 66218
rect 568794 65898 568826 66134
rect 569062 65898 569146 66134
rect 569382 65898 569414 66134
rect 568794 30454 569414 65898
rect 568794 30218 568826 30454
rect 569062 30218 569146 30454
rect 569382 30218 569414 30454
rect 568794 30134 569414 30218
rect 568794 29898 568826 30134
rect 569062 29898 569146 30134
rect 569382 29898 569414 30134
rect 568794 -6106 569414 29898
rect 568794 -6342 568826 -6106
rect 569062 -6342 569146 -6106
rect 569382 -6342 569414 -6106
rect 568794 -6426 569414 -6342
rect 568794 -6662 568826 -6426
rect 569062 -6662 569146 -6426
rect 569382 -6662 569414 -6426
rect 568794 -7654 569414 -6662
rect 573294 711558 573914 711590
rect 573294 711322 573326 711558
rect 573562 711322 573646 711558
rect 573882 711322 573914 711558
rect 573294 711238 573914 711322
rect 573294 711002 573326 711238
rect 573562 711002 573646 711238
rect 573882 711002 573914 711238
rect 573294 682954 573914 711002
rect 573294 682718 573326 682954
rect 573562 682718 573646 682954
rect 573882 682718 573914 682954
rect 573294 682634 573914 682718
rect 573294 682398 573326 682634
rect 573562 682398 573646 682634
rect 573882 682398 573914 682634
rect 573294 646954 573914 682398
rect 573294 646718 573326 646954
rect 573562 646718 573646 646954
rect 573882 646718 573914 646954
rect 573294 646634 573914 646718
rect 573294 646398 573326 646634
rect 573562 646398 573646 646634
rect 573882 646398 573914 646634
rect 573294 610954 573914 646398
rect 573294 610718 573326 610954
rect 573562 610718 573646 610954
rect 573882 610718 573914 610954
rect 573294 610634 573914 610718
rect 573294 610398 573326 610634
rect 573562 610398 573646 610634
rect 573882 610398 573914 610634
rect 573294 574954 573914 610398
rect 573294 574718 573326 574954
rect 573562 574718 573646 574954
rect 573882 574718 573914 574954
rect 573294 574634 573914 574718
rect 573294 574398 573326 574634
rect 573562 574398 573646 574634
rect 573882 574398 573914 574634
rect 573294 538954 573914 574398
rect 573294 538718 573326 538954
rect 573562 538718 573646 538954
rect 573882 538718 573914 538954
rect 573294 538634 573914 538718
rect 573294 538398 573326 538634
rect 573562 538398 573646 538634
rect 573882 538398 573914 538634
rect 573294 502954 573914 538398
rect 573294 502718 573326 502954
rect 573562 502718 573646 502954
rect 573882 502718 573914 502954
rect 573294 502634 573914 502718
rect 573294 502398 573326 502634
rect 573562 502398 573646 502634
rect 573882 502398 573914 502634
rect 573294 466954 573914 502398
rect 573294 466718 573326 466954
rect 573562 466718 573646 466954
rect 573882 466718 573914 466954
rect 573294 466634 573914 466718
rect 573294 466398 573326 466634
rect 573562 466398 573646 466634
rect 573882 466398 573914 466634
rect 573294 430954 573914 466398
rect 573294 430718 573326 430954
rect 573562 430718 573646 430954
rect 573882 430718 573914 430954
rect 573294 430634 573914 430718
rect 573294 430398 573326 430634
rect 573562 430398 573646 430634
rect 573882 430398 573914 430634
rect 573294 394954 573914 430398
rect 573294 394718 573326 394954
rect 573562 394718 573646 394954
rect 573882 394718 573914 394954
rect 573294 394634 573914 394718
rect 573294 394398 573326 394634
rect 573562 394398 573646 394634
rect 573882 394398 573914 394634
rect 573294 358954 573914 394398
rect 573294 358718 573326 358954
rect 573562 358718 573646 358954
rect 573882 358718 573914 358954
rect 573294 358634 573914 358718
rect 573294 358398 573326 358634
rect 573562 358398 573646 358634
rect 573882 358398 573914 358634
rect 573294 322954 573914 358398
rect 573294 322718 573326 322954
rect 573562 322718 573646 322954
rect 573882 322718 573914 322954
rect 573294 322634 573914 322718
rect 573294 322398 573326 322634
rect 573562 322398 573646 322634
rect 573882 322398 573914 322634
rect 573294 286954 573914 322398
rect 573294 286718 573326 286954
rect 573562 286718 573646 286954
rect 573882 286718 573914 286954
rect 573294 286634 573914 286718
rect 573294 286398 573326 286634
rect 573562 286398 573646 286634
rect 573882 286398 573914 286634
rect 573294 250954 573914 286398
rect 573294 250718 573326 250954
rect 573562 250718 573646 250954
rect 573882 250718 573914 250954
rect 573294 250634 573914 250718
rect 573294 250398 573326 250634
rect 573562 250398 573646 250634
rect 573882 250398 573914 250634
rect 573294 214954 573914 250398
rect 573294 214718 573326 214954
rect 573562 214718 573646 214954
rect 573882 214718 573914 214954
rect 573294 214634 573914 214718
rect 573294 214398 573326 214634
rect 573562 214398 573646 214634
rect 573882 214398 573914 214634
rect 573294 178954 573914 214398
rect 573294 178718 573326 178954
rect 573562 178718 573646 178954
rect 573882 178718 573914 178954
rect 573294 178634 573914 178718
rect 573294 178398 573326 178634
rect 573562 178398 573646 178634
rect 573882 178398 573914 178634
rect 573294 142954 573914 178398
rect 573294 142718 573326 142954
rect 573562 142718 573646 142954
rect 573882 142718 573914 142954
rect 573294 142634 573914 142718
rect 573294 142398 573326 142634
rect 573562 142398 573646 142634
rect 573882 142398 573914 142634
rect 573294 106954 573914 142398
rect 573294 106718 573326 106954
rect 573562 106718 573646 106954
rect 573882 106718 573914 106954
rect 573294 106634 573914 106718
rect 573294 106398 573326 106634
rect 573562 106398 573646 106634
rect 573882 106398 573914 106634
rect 573294 70954 573914 106398
rect 573294 70718 573326 70954
rect 573562 70718 573646 70954
rect 573882 70718 573914 70954
rect 573294 70634 573914 70718
rect 573294 70398 573326 70634
rect 573562 70398 573646 70634
rect 573882 70398 573914 70634
rect 573294 34954 573914 70398
rect 573294 34718 573326 34954
rect 573562 34718 573646 34954
rect 573882 34718 573914 34954
rect 573294 34634 573914 34718
rect 573294 34398 573326 34634
rect 573562 34398 573646 34634
rect 573882 34398 573914 34634
rect 573294 -7066 573914 34398
rect 573294 -7302 573326 -7066
rect 573562 -7302 573646 -7066
rect 573882 -7302 573914 -7066
rect 573294 -7386 573914 -7302
rect 573294 -7622 573326 -7386
rect 573562 -7622 573646 -7386
rect 573882 -7622 573914 -7386
rect 573294 -7654 573914 -7622
rect 577794 704838 578414 711590
rect 577794 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 578414 704838
rect 577794 704518 578414 704602
rect 577794 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 578414 704518
rect 577794 687454 578414 704282
rect 577794 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 578414 687454
rect 577794 687134 578414 687218
rect 577794 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 578414 687134
rect 577794 651454 578414 686898
rect 577794 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 578414 651454
rect 577794 651134 578414 651218
rect 577794 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 578414 651134
rect 577794 615454 578414 650898
rect 577794 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 578414 615454
rect 577794 615134 578414 615218
rect 577794 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 578414 615134
rect 577794 579454 578414 614898
rect 577794 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 578414 579454
rect 577794 579134 578414 579218
rect 577794 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 578414 579134
rect 577794 543454 578414 578898
rect 577794 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 578414 543454
rect 577794 543134 578414 543218
rect 577794 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 578414 543134
rect 577794 507454 578414 542898
rect 577794 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 578414 507454
rect 577794 507134 578414 507218
rect 577794 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 578414 507134
rect 577794 471454 578414 506898
rect 577794 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 578414 471454
rect 577794 471134 578414 471218
rect 577794 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 578414 471134
rect 577794 435454 578414 470898
rect 577794 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 578414 435454
rect 577794 435134 578414 435218
rect 577794 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 578414 435134
rect 577794 399454 578414 434898
rect 577794 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 578414 399454
rect 577794 399134 578414 399218
rect 577794 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 578414 399134
rect 577794 363454 578414 398898
rect 577794 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 578414 363454
rect 577794 363134 578414 363218
rect 577794 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 578414 363134
rect 577794 327454 578414 362898
rect 577794 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 578414 327454
rect 577794 327134 578414 327218
rect 577794 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 578414 327134
rect 577794 291454 578414 326898
rect 577794 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 578414 291454
rect 577794 291134 578414 291218
rect 577794 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 578414 291134
rect 577794 255454 578414 290898
rect 577794 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 578414 255454
rect 577794 255134 578414 255218
rect 577794 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 578414 255134
rect 577794 219454 578414 254898
rect 577794 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 578414 219454
rect 577794 219134 578414 219218
rect 577794 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 578414 219134
rect 577794 183454 578414 218898
rect 577794 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 578414 183454
rect 577794 183134 578414 183218
rect 577794 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 578414 183134
rect 577794 147454 578414 182898
rect 577794 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 578414 147454
rect 577794 147134 578414 147218
rect 577794 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 578414 147134
rect 577794 111454 578414 146898
rect 577794 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 578414 111454
rect 577794 111134 578414 111218
rect 577794 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 578414 111134
rect 577794 75454 578414 110898
rect 577794 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 578414 75454
rect 577794 75134 578414 75218
rect 577794 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 578414 75134
rect 577794 39454 578414 74898
rect 577794 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 578414 39454
rect 577794 39134 578414 39218
rect 577794 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 578414 39134
rect 577794 3454 578414 38898
rect 577794 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 578414 3454
rect 577794 3134 578414 3218
rect 577794 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 578414 3134
rect 577794 -346 578414 2898
rect 577794 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 578414 -346
rect 577794 -666 578414 -582
rect 577794 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 578414 -666
rect 577794 -7654 578414 -902
rect 582294 705798 582914 711590
rect 592030 711558 592650 711590
rect 592030 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect 592030 711238 592650 711322
rect 592030 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect 591070 710598 591690 710630
rect 591070 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect 591070 710278 591690 710362
rect 591070 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect 590110 709638 590730 709670
rect 590110 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect 590110 709318 590730 709402
rect 590110 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect 589150 708678 589770 708710
rect 589150 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect 589150 708358 589770 708442
rect 589150 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect 588190 707718 588810 707750
rect 588190 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect 588190 707398 588810 707482
rect 588190 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect 587230 706758 587850 706790
rect 587230 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect 587230 706438 587850 706522
rect 587230 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect 582294 705562 582326 705798
rect 582562 705562 582646 705798
rect 582882 705562 582914 705798
rect 582294 705478 582914 705562
rect 582294 705242 582326 705478
rect 582562 705242 582646 705478
rect 582882 705242 582914 705478
rect 582294 691954 582914 705242
rect 586270 705798 586890 705830
rect 586270 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect 586270 705478 586890 705562
rect 586270 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect 582294 691718 582326 691954
rect 582562 691718 582646 691954
rect 582882 691718 582914 691954
rect 582294 691634 582914 691718
rect 582294 691398 582326 691634
rect 582562 691398 582646 691634
rect 582882 691398 582914 691634
rect 582294 655954 582914 691398
rect 582294 655718 582326 655954
rect 582562 655718 582646 655954
rect 582882 655718 582914 655954
rect 582294 655634 582914 655718
rect 582294 655398 582326 655634
rect 582562 655398 582646 655634
rect 582882 655398 582914 655634
rect 582294 619954 582914 655398
rect 582294 619718 582326 619954
rect 582562 619718 582646 619954
rect 582882 619718 582914 619954
rect 582294 619634 582914 619718
rect 582294 619398 582326 619634
rect 582562 619398 582646 619634
rect 582882 619398 582914 619634
rect 582294 583954 582914 619398
rect 582294 583718 582326 583954
rect 582562 583718 582646 583954
rect 582882 583718 582914 583954
rect 582294 583634 582914 583718
rect 582294 583398 582326 583634
rect 582562 583398 582646 583634
rect 582882 583398 582914 583634
rect 582294 547954 582914 583398
rect 582294 547718 582326 547954
rect 582562 547718 582646 547954
rect 582882 547718 582914 547954
rect 582294 547634 582914 547718
rect 582294 547398 582326 547634
rect 582562 547398 582646 547634
rect 582882 547398 582914 547634
rect 582294 511954 582914 547398
rect 582294 511718 582326 511954
rect 582562 511718 582646 511954
rect 582882 511718 582914 511954
rect 582294 511634 582914 511718
rect 582294 511398 582326 511634
rect 582562 511398 582646 511634
rect 582882 511398 582914 511634
rect 582294 475954 582914 511398
rect 582294 475718 582326 475954
rect 582562 475718 582646 475954
rect 582882 475718 582914 475954
rect 582294 475634 582914 475718
rect 582294 475398 582326 475634
rect 582562 475398 582646 475634
rect 582882 475398 582914 475634
rect 582294 439954 582914 475398
rect 582294 439718 582326 439954
rect 582562 439718 582646 439954
rect 582882 439718 582914 439954
rect 582294 439634 582914 439718
rect 582294 439398 582326 439634
rect 582562 439398 582646 439634
rect 582882 439398 582914 439634
rect 582294 403954 582914 439398
rect 582294 403718 582326 403954
rect 582562 403718 582646 403954
rect 582882 403718 582914 403954
rect 582294 403634 582914 403718
rect 582294 403398 582326 403634
rect 582562 403398 582646 403634
rect 582882 403398 582914 403634
rect 582294 367954 582914 403398
rect 582294 367718 582326 367954
rect 582562 367718 582646 367954
rect 582882 367718 582914 367954
rect 582294 367634 582914 367718
rect 582294 367398 582326 367634
rect 582562 367398 582646 367634
rect 582882 367398 582914 367634
rect 582294 331954 582914 367398
rect 582294 331718 582326 331954
rect 582562 331718 582646 331954
rect 582882 331718 582914 331954
rect 582294 331634 582914 331718
rect 582294 331398 582326 331634
rect 582562 331398 582646 331634
rect 582882 331398 582914 331634
rect 582294 295954 582914 331398
rect 582294 295718 582326 295954
rect 582562 295718 582646 295954
rect 582882 295718 582914 295954
rect 582294 295634 582914 295718
rect 582294 295398 582326 295634
rect 582562 295398 582646 295634
rect 582882 295398 582914 295634
rect 582294 259954 582914 295398
rect 582294 259718 582326 259954
rect 582562 259718 582646 259954
rect 582882 259718 582914 259954
rect 582294 259634 582914 259718
rect 582294 259398 582326 259634
rect 582562 259398 582646 259634
rect 582882 259398 582914 259634
rect 582294 223954 582914 259398
rect 582294 223718 582326 223954
rect 582562 223718 582646 223954
rect 582882 223718 582914 223954
rect 582294 223634 582914 223718
rect 582294 223398 582326 223634
rect 582562 223398 582646 223634
rect 582882 223398 582914 223634
rect 582294 187954 582914 223398
rect 582294 187718 582326 187954
rect 582562 187718 582646 187954
rect 582882 187718 582914 187954
rect 582294 187634 582914 187718
rect 582294 187398 582326 187634
rect 582562 187398 582646 187634
rect 582882 187398 582914 187634
rect 582294 151954 582914 187398
rect 582294 151718 582326 151954
rect 582562 151718 582646 151954
rect 582882 151718 582914 151954
rect 582294 151634 582914 151718
rect 582294 151398 582326 151634
rect 582562 151398 582646 151634
rect 582882 151398 582914 151634
rect 582294 115954 582914 151398
rect 582294 115718 582326 115954
rect 582562 115718 582646 115954
rect 582882 115718 582914 115954
rect 582294 115634 582914 115718
rect 582294 115398 582326 115634
rect 582562 115398 582646 115634
rect 582882 115398 582914 115634
rect 582294 79954 582914 115398
rect 582294 79718 582326 79954
rect 582562 79718 582646 79954
rect 582882 79718 582914 79954
rect 582294 79634 582914 79718
rect 582294 79398 582326 79634
rect 582562 79398 582646 79634
rect 582882 79398 582914 79634
rect 582294 43954 582914 79398
rect 582294 43718 582326 43954
rect 582562 43718 582646 43954
rect 582882 43718 582914 43954
rect 582294 43634 582914 43718
rect 582294 43398 582326 43634
rect 582562 43398 582646 43634
rect 582882 43398 582914 43634
rect 582294 7954 582914 43398
rect 582294 7718 582326 7954
rect 582562 7718 582646 7954
rect 582882 7718 582914 7954
rect 582294 7634 582914 7718
rect 582294 7398 582326 7634
rect 582562 7398 582646 7634
rect 582882 7398 582914 7634
rect 582294 -1306 582914 7398
rect 585310 704838 585930 704870
rect 585310 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect 585310 704518 585930 704602
rect 585310 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect 585310 687454 585930 704282
rect 585310 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 585930 687454
rect 585310 687134 585930 687218
rect 585310 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 585930 687134
rect 585310 651454 585930 686898
rect 585310 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 585930 651454
rect 585310 651134 585930 651218
rect 585310 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 585930 651134
rect 585310 615454 585930 650898
rect 585310 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 585930 615454
rect 585310 615134 585930 615218
rect 585310 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 585930 615134
rect 585310 579454 585930 614898
rect 585310 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 585930 579454
rect 585310 579134 585930 579218
rect 585310 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 585930 579134
rect 585310 543454 585930 578898
rect 585310 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 585930 543454
rect 585310 543134 585930 543218
rect 585310 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 585930 543134
rect 585310 507454 585930 542898
rect 585310 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 585930 507454
rect 585310 507134 585930 507218
rect 585310 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 585930 507134
rect 585310 471454 585930 506898
rect 585310 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 585930 471454
rect 585310 471134 585930 471218
rect 585310 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 585930 471134
rect 585310 435454 585930 470898
rect 585310 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 585930 435454
rect 585310 435134 585930 435218
rect 585310 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 585930 435134
rect 585310 399454 585930 434898
rect 585310 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 585930 399454
rect 585310 399134 585930 399218
rect 585310 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 585930 399134
rect 585310 363454 585930 398898
rect 585310 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 585930 363454
rect 585310 363134 585930 363218
rect 585310 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 585930 363134
rect 585310 327454 585930 362898
rect 585310 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 585930 327454
rect 585310 327134 585930 327218
rect 585310 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 585930 327134
rect 585310 291454 585930 326898
rect 585310 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 585930 291454
rect 585310 291134 585930 291218
rect 585310 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 585930 291134
rect 585310 255454 585930 290898
rect 585310 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 585930 255454
rect 585310 255134 585930 255218
rect 585310 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 585930 255134
rect 585310 219454 585930 254898
rect 585310 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 585930 219454
rect 585310 219134 585930 219218
rect 585310 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 585930 219134
rect 585310 183454 585930 218898
rect 585310 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 585930 183454
rect 585310 183134 585930 183218
rect 585310 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 585930 183134
rect 585310 147454 585930 182898
rect 585310 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 585930 147454
rect 585310 147134 585930 147218
rect 585310 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 585930 147134
rect 585310 111454 585930 146898
rect 585310 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 585930 111454
rect 585310 111134 585930 111218
rect 585310 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 585930 111134
rect 585310 75454 585930 110898
rect 585310 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 585930 75454
rect 585310 75134 585930 75218
rect 585310 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 585930 75134
rect 585310 39454 585930 74898
rect 585310 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 585930 39454
rect 585310 39134 585930 39218
rect 585310 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 585930 39134
rect 585310 3454 585930 38898
rect 585310 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 585930 3454
rect 585310 3134 585930 3218
rect 585310 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 585930 3134
rect 585310 -346 585930 2898
rect 585310 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect 585310 -666 585930 -582
rect 585310 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect 585310 -934 585930 -902
rect 586270 691954 586890 705242
rect 586270 691718 586302 691954
rect 586538 691718 586622 691954
rect 586858 691718 586890 691954
rect 586270 691634 586890 691718
rect 586270 691398 586302 691634
rect 586538 691398 586622 691634
rect 586858 691398 586890 691634
rect 586270 655954 586890 691398
rect 586270 655718 586302 655954
rect 586538 655718 586622 655954
rect 586858 655718 586890 655954
rect 586270 655634 586890 655718
rect 586270 655398 586302 655634
rect 586538 655398 586622 655634
rect 586858 655398 586890 655634
rect 586270 619954 586890 655398
rect 586270 619718 586302 619954
rect 586538 619718 586622 619954
rect 586858 619718 586890 619954
rect 586270 619634 586890 619718
rect 586270 619398 586302 619634
rect 586538 619398 586622 619634
rect 586858 619398 586890 619634
rect 586270 583954 586890 619398
rect 586270 583718 586302 583954
rect 586538 583718 586622 583954
rect 586858 583718 586890 583954
rect 586270 583634 586890 583718
rect 586270 583398 586302 583634
rect 586538 583398 586622 583634
rect 586858 583398 586890 583634
rect 586270 547954 586890 583398
rect 586270 547718 586302 547954
rect 586538 547718 586622 547954
rect 586858 547718 586890 547954
rect 586270 547634 586890 547718
rect 586270 547398 586302 547634
rect 586538 547398 586622 547634
rect 586858 547398 586890 547634
rect 586270 511954 586890 547398
rect 586270 511718 586302 511954
rect 586538 511718 586622 511954
rect 586858 511718 586890 511954
rect 586270 511634 586890 511718
rect 586270 511398 586302 511634
rect 586538 511398 586622 511634
rect 586858 511398 586890 511634
rect 586270 475954 586890 511398
rect 586270 475718 586302 475954
rect 586538 475718 586622 475954
rect 586858 475718 586890 475954
rect 586270 475634 586890 475718
rect 586270 475398 586302 475634
rect 586538 475398 586622 475634
rect 586858 475398 586890 475634
rect 586270 439954 586890 475398
rect 586270 439718 586302 439954
rect 586538 439718 586622 439954
rect 586858 439718 586890 439954
rect 586270 439634 586890 439718
rect 586270 439398 586302 439634
rect 586538 439398 586622 439634
rect 586858 439398 586890 439634
rect 586270 403954 586890 439398
rect 586270 403718 586302 403954
rect 586538 403718 586622 403954
rect 586858 403718 586890 403954
rect 586270 403634 586890 403718
rect 586270 403398 586302 403634
rect 586538 403398 586622 403634
rect 586858 403398 586890 403634
rect 586270 367954 586890 403398
rect 586270 367718 586302 367954
rect 586538 367718 586622 367954
rect 586858 367718 586890 367954
rect 586270 367634 586890 367718
rect 586270 367398 586302 367634
rect 586538 367398 586622 367634
rect 586858 367398 586890 367634
rect 586270 331954 586890 367398
rect 586270 331718 586302 331954
rect 586538 331718 586622 331954
rect 586858 331718 586890 331954
rect 586270 331634 586890 331718
rect 586270 331398 586302 331634
rect 586538 331398 586622 331634
rect 586858 331398 586890 331634
rect 586270 295954 586890 331398
rect 586270 295718 586302 295954
rect 586538 295718 586622 295954
rect 586858 295718 586890 295954
rect 586270 295634 586890 295718
rect 586270 295398 586302 295634
rect 586538 295398 586622 295634
rect 586858 295398 586890 295634
rect 586270 259954 586890 295398
rect 586270 259718 586302 259954
rect 586538 259718 586622 259954
rect 586858 259718 586890 259954
rect 586270 259634 586890 259718
rect 586270 259398 586302 259634
rect 586538 259398 586622 259634
rect 586858 259398 586890 259634
rect 586270 223954 586890 259398
rect 586270 223718 586302 223954
rect 586538 223718 586622 223954
rect 586858 223718 586890 223954
rect 586270 223634 586890 223718
rect 586270 223398 586302 223634
rect 586538 223398 586622 223634
rect 586858 223398 586890 223634
rect 586270 187954 586890 223398
rect 586270 187718 586302 187954
rect 586538 187718 586622 187954
rect 586858 187718 586890 187954
rect 586270 187634 586890 187718
rect 586270 187398 586302 187634
rect 586538 187398 586622 187634
rect 586858 187398 586890 187634
rect 586270 151954 586890 187398
rect 586270 151718 586302 151954
rect 586538 151718 586622 151954
rect 586858 151718 586890 151954
rect 586270 151634 586890 151718
rect 586270 151398 586302 151634
rect 586538 151398 586622 151634
rect 586858 151398 586890 151634
rect 586270 115954 586890 151398
rect 586270 115718 586302 115954
rect 586538 115718 586622 115954
rect 586858 115718 586890 115954
rect 586270 115634 586890 115718
rect 586270 115398 586302 115634
rect 586538 115398 586622 115634
rect 586858 115398 586890 115634
rect 586270 79954 586890 115398
rect 586270 79718 586302 79954
rect 586538 79718 586622 79954
rect 586858 79718 586890 79954
rect 586270 79634 586890 79718
rect 586270 79398 586302 79634
rect 586538 79398 586622 79634
rect 586858 79398 586890 79634
rect 586270 43954 586890 79398
rect 586270 43718 586302 43954
rect 586538 43718 586622 43954
rect 586858 43718 586890 43954
rect 586270 43634 586890 43718
rect 586270 43398 586302 43634
rect 586538 43398 586622 43634
rect 586858 43398 586890 43634
rect 586270 7954 586890 43398
rect 586270 7718 586302 7954
rect 586538 7718 586622 7954
rect 586858 7718 586890 7954
rect 586270 7634 586890 7718
rect 586270 7398 586302 7634
rect 586538 7398 586622 7634
rect 586858 7398 586890 7634
rect 582294 -1542 582326 -1306
rect 582562 -1542 582646 -1306
rect 582882 -1542 582914 -1306
rect 582294 -1626 582914 -1542
rect 582294 -1862 582326 -1626
rect 582562 -1862 582646 -1626
rect 582882 -1862 582914 -1626
rect 582294 -7654 582914 -1862
rect 586270 -1306 586890 7398
rect 586270 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect 586270 -1626 586890 -1542
rect 586270 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect 586270 -1894 586890 -1862
rect 587230 696454 587850 706202
rect 587230 696218 587262 696454
rect 587498 696218 587582 696454
rect 587818 696218 587850 696454
rect 587230 696134 587850 696218
rect 587230 695898 587262 696134
rect 587498 695898 587582 696134
rect 587818 695898 587850 696134
rect 587230 660454 587850 695898
rect 587230 660218 587262 660454
rect 587498 660218 587582 660454
rect 587818 660218 587850 660454
rect 587230 660134 587850 660218
rect 587230 659898 587262 660134
rect 587498 659898 587582 660134
rect 587818 659898 587850 660134
rect 587230 624454 587850 659898
rect 587230 624218 587262 624454
rect 587498 624218 587582 624454
rect 587818 624218 587850 624454
rect 587230 624134 587850 624218
rect 587230 623898 587262 624134
rect 587498 623898 587582 624134
rect 587818 623898 587850 624134
rect 587230 588454 587850 623898
rect 587230 588218 587262 588454
rect 587498 588218 587582 588454
rect 587818 588218 587850 588454
rect 587230 588134 587850 588218
rect 587230 587898 587262 588134
rect 587498 587898 587582 588134
rect 587818 587898 587850 588134
rect 587230 552454 587850 587898
rect 587230 552218 587262 552454
rect 587498 552218 587582 552454
rect 587818 552218 587850 552454
rect 587230 552134 587850 552218
rect 587230 551898 587262 552134
rect 587498 551898 587582 552134
rect 587818 551898 587850 552134
rect 587230 516454 587850 551898
rect 587230 516218 587262 516454
rect 587498 516218 587582 516454
rect 587818 516218 587850 516454
rect 587230 516134 587850 516218
rect 587230 515898 587262 516134
rect 587498 515898 587582 516134
rect 587818 515898 587850 516134
rect 587230 480454 587850 515898
rect 587230 480218 587262 480454
rect 587498 480218 587582 480454
rect 587818 480218 587850 480454
rect 587230 480134 587850 480218
rect 587230 479898 587262 480134
rect 587498 479898 587582 480134
rect 587818 479898 587850 480134
rect 587230 444454 587850 479898
rect 587230 444218 587262 444454
rect 587498 444218 587582 444454
rect 587818 444218 587850 444454
rect 587230 444134 587850 444218
rect 587230 443898 587262 444134
rect 587498 443898 587582 444134
rect 587818 443898 587850 444134
rect 587230 408454 587850 443898
rect 587230 408218 587262 408454
rect 587498 408218 587582 408454
rect 587818 408218 587850 408454
rect 587230 408134 587850 408218
rect 587230 407898 587262 408134
rect 587498 407898 587582 408134
rect 587818 407898 587850 408134
rect 587230 372454 587850 407898
rect 587230 372218 587262 372454
rect 587498 372218 587582 372454
rect 587818 372218 587850 372454
rect 587230 372134 587850 372218
rect 587230 371898 587262 372134
rect 587498 371898 587582 372134
rect 587818 371898 587850 372134
rect 587230 336454 587850 371898
rect 587230 336218 587262 336454
rect 587498 336218 587582 336454
rect 587818 336218 587850 336454
rect 587230 336134 587850 336218
rect 587230 335898 587262 336134
rect 587498 335898 587582 336134
rect 587818 335898 587850 336134
rect 587230 300454 587850 335898
rect 587230 300218 587262 300454
rect 587498 300218 587582 300454
rect 587818 300218 587850 300454
rect 587230 300134 587850 300218
rect 587230 299898 587262 300134
rect 587498 299898 587582 300134
rect 587818 299898 587850 300134
rect 587230 264454 587850 299898
rect 587230 264218 587262 264454
rect 587498 264218 587582 264454
rect 587818 264218 587850 264454
rect 587230 264134 587850 264218
rect 587230 263898 587262 264134
rect 587498 263898 587582 264134
rect 587818 263898 587850 264134
rect 587230 228454 587850 263898
rect 587230 228218 587262 228454
rect 587498 228218 587582 228454
rect 587818 228218 587850 228454
rect 587230 228134 587850 228218
rect 587230 227898 587262 228134
rect 587498 227898 587582 228134
rect 587818 227898 587850 228134
rect 587230 192454 587850 227898
rect 587230 192218 587262 192454
rect 587498 192218 587582 192454
rect 587818 192218 587850 192454
rect 587230 192134 587850 192218
rect 587230 191898 587262 192134
rect 587498 191898 587582 192134
rect 587818 191898 587850 192134
rect 587230 156454 587850 191898
rect 587230 156218 587262 156454
rect 587498 156218 587582 156454
rect 587818 156218 587850 156454
rect 587230 156134 587850 156218
rect 587230 155898 587262 156134
rect 587498 155898 587582 156134
rect 587818 155898 587850 156134
rect 587230 120454 587850 155898
rect 587230 120218 587262 120454
rect 587498 120218 587582 120454
rect 587818 120218 587850 120454
rect 587230 120134 587850 120218
rect 587230 119898 587262 120134
rect 587498 119898 587582 120134
rect 587818 119898 587850 120134
rect 587230 84454 587850 119898
rect 587230 84218 587262 84454
rect 587498 84218 587582 84454
rect 587818 84218 587850 84454
rect 587230 84134 587850 84218
rect 587230 83898 587262 84134
rect 587498 83898 587582 84134
rect 587818 83898 587850 84134
rect 587230 48454 587850 83898
rect 587230 48218 587262 48454
rect 587498 48218 587582 48454
rect 587818 48218 587850 48454
rect 587230 48134 587850 48218
rect 587230 47898 587262 48134
rect 587498 47898 587582 48134
rect 587818 47898 587850 48134
rect 587230 12454 587850 47898
rect 587230 12218 587262 12454
rect 587498 12218 587582 12454
rect 587818 12218 587850 12454
rect 587230 12134 587850 12218
rect 587230 11898 587262 12134
rect 587498 11898 587582 12134
rect 587818 11898 587850 12134
rect 587230 -2266 587850 11898
rect 587230 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect 587230 -2586 587850 -2502
rect 587230 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect 587230 -2854 587850 -2822
rect 588190 700954 588810 707162
rect 588190 700718 588222 700954
rect 588458 700718 588542 700954
rect 588778 700718 588810 700954
rect 588190 700634 588810 700718
rect 588190 700398 588222 700634
rect 588458 700398 588542 700634
rect 588778 700398 588810 700634
rect 588190 664954 588810 700398
rect 588190 664718 588222 664954
rect 588458 664718 588542 664954
rect 588778 664718 588810 664954
rect 588190 664634 588810 664718
rect 588190 664398 588222 664634
rect 588458 664398 588542 664634
rect 588778 664398 588810 664634
rect 588190 628954 588810 664398
rect 588190 628718 588222 628954
rect 588458 628718 588542 628954
rect 588778 628718 588810 628954
rect 588190 628634 588810 628718
rect 588190 628398 588222 628634
rect 588458 628398 588542 628634
rect 588778 628398 588810 628634
rect 588190 592954 588810 628398
rect 588190 592718 588222 592954
rect 588458 592718 588542 592954
rect 588778 592718 588810 592954
rect 588190 592634 588810 592718
rect 588190 592398 588222 592634
rect 588458 592398 588542 592634
rect 588778 592398 588810 592634
rect 588190 556954 588810 592398
rect 588190 556718 588222 556954
rect 588458 556718 588542 556954
rect 588778 556718 588810 556954
rect 588190 556634 588810 556718
rect 588190 556398 588222 556634
rect 588458 556398 588542 556634
rect 588778 556398 588810 556634
rect 588190 520954 588810 556398
rect 588190 520718 588222 520954
rect 588458 520718 588542 520954
rect 588778 520718 588810 520954
rect 588190 520634 588810 520718
rect 588190 520398 588222 520634
rect 588458 520398 588542 520634
rect 588778 520398 588810 520634
rect 588190 484954 588810 520398
rect 588190 484718 588222 484954
rect 588458 484718 588542 484954
rect 588778 484718 588810 484954
rect 588190 484634 588810 484718
rect 588190 484398 588222 484634
rect 588458 484398 588542 484634
rect 588778 484398 588810 484634
rect 588190 448954 588810 484398
rect 588190 448718 588222 448954
rect 588458 448718 588542 448954
rect 588778 448718 588810 448954
rect 588190 448634 588810 448718
rect 588190 448398 588222 448634
rect 588458 448398 588542 448634
rect 588778 448398 588810 448634
rect 588190 412954 588810 448398
rect 588190 412718 588222 412954
rect 588458 412718 588542 412954
rect 588778 412718 588810 412954
rect 588190 412634 588810 412718
rect 588190 412398 588222 412634
rect 588458 412398 588542 412634
rect 588778 412398 588810 412634
rect 588190 376954 588810 412398
rect 588190 376718 588222 376954
rect 588458 376718 588542 376954
rect 588778 376718 588810 376954
rect 588190 376634 588810 376718
rect 588190 376398 588222 376634
rect 588458 376398 588542 376634
rect 588778 376398 588810 376634
rect 588190 340954 588810 376398
rect 588190 340718 588222 340954
rect 588458 340718 588542 340954
rect 588778 340718 588810 340954
rect 588190 340634 588810 340718
rect 588190 340398 588222 340634
rect 588458 340398 588542 340634
rect 588778 340398 588810 340634
rect 588190 304954 588810 340398
rect 588190 304718 588222 304954
rect 588458 304718 588542 304954
rect 588778 304718 588810 304954
rect 588190 304634 588810 304718
rect 588190 304398 588222 304634
rect 588458 304398 588542 304634
rect 588778 304398 588810 304634
rect 588190 268954 588810 304398
rect 588190 268718 588222 268954
rect 588458 268718 588542 268954
rect 588778 268718 588810 268954
rect 588190 268634 588810 268718
rect 588190 268398 588222 268634
rect 588458 268398 588542 268634
rect 588778 268398 588810 268634
rect 588190 232954 588810 268398
rect 588190 232718 588222 232954
rect 588458 232718 588542 232954
rect 588778 232718 588810 232954
rect 588190 232634 588810 232718
rect 588190 232398 588222 232634
rect 588458 232398 588542 232634
rect 588778 232398 588810 232634
rect 588190 196954 588810 232398
rect 588190 196718 588222 196954
rect 588458 196718 588542 196954
rect 588778 196718 588810 196954
rect 588190 196634 588810 196718
rect 588190 196398 588222 196634
rect 588458 196398 588542 196634
rect 588778 196398 588810 196634
rect 588190 160954 588810 196398
rect 588190 160718 588222 160954
rect 588458 160718 588542 160954
rect 588778 160718 588810 160954
rect 588190 160634 588810 160718
rect 588190 160398 588222 160634
rect 588458 160398 588542 160634
rect 588778 160398 588810 160634
rect 588190 124954 588810 160398
rect 588190 124718 588222 124954
rect 588458 124718 588542 124954
rect 588778 124718 588810 124954
rect 588190 124634 588810 124718
rect 588190 124398 588222 124634
rect 588458 124398 588542 124634
rect 588778 124398 588810 124634
rect 588190 88954 588810 124398
rect 588190 88718 588222 88954
rect 588458 88718 588542 88954
rect 588778 88718 588810 88954
rect 588190 88634 588810 88718
rect 588190 88398 588222 88634
rect 588458 88398 588542 88634
rect 588778 88398 588810 88634
rect 588190 52954 588810 88398
rect 588190 52718 588222 52954
rect 588458 52718 588542 52954
rect 588778 52718 588810 52954
rect 588190 52634 588810 52718
rect 588190 52398 588222 52634
rect 588458 52398 588542 52634
rect 588778 52398 588810 52634
rect 588190 16954 588810 52398
rect 588190 16718 588222 16954
rect 588458 16718 588542 16954
rect 588778 16718 588810 16954
rect 588190 16634 588810 16718
rect 588190 16398 588222 16634
rect 588458 16398 588542 16634
rect 588778 16398 588810 16634
rect 588190 -3226 588810 16398
rect 588190 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect 588190 -3546 588810 -3462
rect 588190 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect 588190 -3814 588810 -3782
rect 589150 669454 589770 708122
rect 589150 669218 589182 669454
rect 589418 669218 589502 669454
rect 589738 669218 589770 669454
rect 589150 669134 589770 669218
rect 589150 668898 589182 669134
rect 589418 668898 589502 669134
rect 589738 668898 589770 669134
rect 589150 633454 589770 668898
rect 589150 633218 589182 633454
rect 589418 633218 589502 633454
rect 589738 633218 589770 633454
rect 589150 633134 589770 633218
rect 589150 632898 589182 633134
rect 589418 632898 589502 633134
rect 589738 632898 589770 633134
rect 589150 597454 589770 632898
rect 589150 597218 589182 597454
rect 589418 597218 589502 597454
rect 589738 597218 589770 597454
rect 589150 597134 589770 597218
rect 589150 596898 589182 597134
rect 589418 596898 589502 597134
rect 589738 596898 589770 597134
rect 589150 561454 589770 596898
rect 589150 561218 589182 561454
rect 589418 561218 589502 561454
rect 589738 561218 589770 561454
rect 589150 561134 589770 561218
rect 589150 560898 589182 561134
rect 589418 560898 589502 561134
rect 589738 560898 589770 561134
rect 589150 525454 589770 560898
rect 589150 525218 589182 525454
rect 589418 525218 589502 525454
rect 589738 525218 589770 525454
rect 589150 525134 589770 525218
rect 589150 524898 589182 525134
rect 589418 524898 589502 525134
rect 589738 524898 589770 525134
rect 589150 489454 589770 524898
rect 589150 489218 589182 489454
rect 589418 489218 589502 489454
rect 589738 489218 589770 489454
rect 589150 489134 589770 489218
rect 589150 488898 589182 489134
rect 589418 488898 589502 489134
rect 589738 488898 589770 489134
rect 589150 453454 589770 488898
rect 589150 453218 589182 453454
rect 589418 453218 589502 453454
rect 589738 453218 589770 453454
rect 589150 453134 589770 453218
rect 589150 452898 589182 453134
rect 589418 452898 589502 453134
rect 589738 452898 589770 453134
rect 589150 417454 589770 452898
rect 589150 417218 589182 417454
rect 589418 417218 589502 417454
rect 589738 417218 589770 417454
rect 589150 417134 589770 417218
rect 589150 416898 589182 417134
rect 589418 416898 589502 417134
rect 589738 416898 589770 417134
rect 589150 381454 589770 416898
rect 589150 381218 589182 381454
rect 589418 381218 589502 381454
rect 589738 381218 589770 381454
rect 589150 381134 589770 381218
rect 589150 380898 589182 381134
rect 589418 380898 589502 381134
rect 589738 380898 589770 381134
rect 589150 345454 589770 380898
rect 589150 345218 589182 345454
rect 589418 345218 589502 345454
rect 589738 345218 589770 345454
rect 589150 345134 589770 345218
rect 589150 344898 589182 345134
rect 589418 344898 589502 345134
rect 589738 344898 589770 345134
rect 589150 309454 589770 344898
rect 589150 309218 589182 309454
rect 589418 309218 589502 309454
rect 589738 309218 589770 309454
rect 589150 309134 589770 309218
rect 589150 308898 589182 309134
rect 589418 308898 589502 309134
rect 589738 308898 589770 309134
rect 589150 273454 589770 308898
rect 589150 273218 589182 273454
rect 589418 273218 589502 273454
rect 589738 273218 589770 273454
rect 589150 273134 589770 273218
rect 589150 272898 589182 273134
rect 589418 272898 589502 273134
rect 589738 272898 589770 273134
rect 589150 237454 589770 272898
rect 589150 237218 589182 237454
rect 589418 237218 589502 237454
rect 589738 237218 589770 237454
rect 589150 237134 589770 237218
rect 589150 236898 589182 237134
rect 589418 236898 589502 237134
rect 589738 236898 589770 237134
rect 589150 201454 589770 236898
rect 589150 201218 589182 201454
rect 589418 201218 589502 201454
rect 589738 201218 589770 201454
rect 589150 201134 589770 201218
rect 589150 200898 589182 201134
rect 589418 200898 589502 201134
rect 589738 200898 589770 201134
rect 589150 165454 589770 200898
rect 589150 165218 589182 165454
rect 589418 165218 589502 165454
rect 589738 165218 589770 165454
rect 589150 165134 589770 165218
rect 589150 164898 589182 165134
rect 589418 164898 589502 165134
rect 589738 164898 589770 165134
rect 589150 129454 589770 164898
rect 589150 129218 589182 129454
rect 589418 129218 589502 129454
rect 589738 129218 589770 129454
rect 589150 129134 589770 129218
rect 589150 128898 589182 129134
rect 589418 128898 589502 129134
rect 589738 128898 589770 129134
rect 589150 93454 589770 128898
rect 589150 93218 589182 93454
rect 589418 93218 589502 93454
rect 589738 93218 589770 93454
rect 589150 93134 589770 93218
rect 589150 92898 589182 93134
rect 589418 92898 589502 93134
rect 589738 92898 589770 93134
rect 589150 57454 589770 92898
rect 589150 57218 589182 57454
rect 589418 57218 589502 57454
rect 589738 57218 589770 57454
rect 589150 57134 589770 57218
rect 589150 56898 589182 57134
rect 589418 56898 589502 57134
rect 589738 56898 589770 57134
rect 589150 21454 589770 56898
rect 589150 21218 589182 21454
rect 589418 21218 589502 21454
rect 589738 21218 589770 21454
rect 589150 21134 589770 21218
rect 589150 20898 589182 21134
rect 589418 20898 589502 21134
rect 589738 20898 589770 21134
rect 589150 -4186 589770 20898
rect 589150 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect 589150 -4506 589770 -4422
rect 589150 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect 589150 -4774 589770 -4742
rect 590110 673954 590730 709082
rect 590110 673718 590142 673954
rect 590378 673718 590462 673954
rect 590698 673718 590730 673954
rect 590110 673634 590730 673718
rect 590110 673398 590142 673634
rect 590378 673398 590462 673634
rect 590698 673398 590730 673634
rect 590110 637954 590730 673398
rect 590110 637718 590142 637954
rect 590378 637718 590462 637954
rect 590698 637718 590730 637954
rect 590110 637634 590730 637718
rect 590110 637398 590142 637634
rect 590378 637398 590462 637634
rect 590698 637398 590730 637634
rect 590110 601954 590730 637398
rect 590110 601718 590142 601954
rect 590378 601718 590462 601954
rect 590698 601718 590730 601954
rect 590110 601634 590730 601718
rect 590110 601398 590142 601634
rect 590378 601398 590462 601634
rect 590698 601398 590730 601634
rect 590110 565954 590730 601398
rect 590110 565718 590142 565954
rect 590378 565718 590462 565954
rect 590698 565718 590730 565954
rect 590110 565634 590730 565718
rect 590110 565398 590142 565634
rect 590378 565398 590462 565634
rect 590698 565398 590730 565634
rect 590110 529954 590730 565398
rect 590110 529718 590142 529954
rect 590378 529718 590462 529954
rect 590698 529718 590730 529954
rect 590110 529634 590730 529718
rect 590110 529398 590142 529634
rect 590378 529398 590462 529634
rect 590698 529398 590730 529634
rect 590110 493954 590730 529398
rect 590110 493718 590142 493954
rect 590378 493718 590462 493954
rect 590698 493718 590730 493954
rect 590110 493634 590730 493718
rect 590110 493398 590142 493634
rect 590378 493398 590462 493634
rect 590698 493398 590730 493634
rect 590110 457954 590730 493398
rect 590110 457718 590142 457954
rect 590378 457718 590462 457954
rect 590698 457718 590730 457954
rect 590110 457634 590730 457718
rect 590110 457398 590142 457634
rect 590378 457398 590462 457634
rect 590698 457398 590730 457634
rect 590110 421954 590730 457398
rect 590110 421718 590142 421954
rect 590378 421718 590462 421954
rect 590698 421718 590730 421954
rect 590110 421634 590730 421718
rect 590110 421398 590142 421634
rect 590378 421398 590462 421634
rect 590698 421398 590730 421634
rect 590110 385954 590730 421398
rect 590110 385718 590142 385954
rect 590378 385718 590462 385954
rect 590698 385718 590730 385954
rect 590110 385634 590730 385718
rect 590110 385398 590142 385634
rect 590378 385398 590462 385634
rect 590698 385398 590730 385634
rect 590110 349954 590730 385398
rect 590110 349718 590142 349954
rect 590378 349718 590462 349954
rect 590698 349718 590730 349954
rect 590110 349634 590730 349718
rect 590110 349398 590142 349634
rect 590378 349398 590462 349634
rect 590698 349398 590730 349634
rect 590110 313954 590730 349398
rect 590110 313718 590142 313954
rect 590378 313718 590462 313954
rect 590698 313718 590730 313954
rect 590110 313634 590730 313718
rect 590110 313398 590142 313634
rect 590378 313398 590462 313634
rect 590698 313398 590730 313634
rect 590110 277954 590730 313398
rect 590110 277718 590142 277954
rect 590378 277718 590462 277954
rect 590698 277718 590730 277954
rect 590110 277634 590730 277718
rect 590110 277398 590142 277634
rect 590378 277398 590462 277634
rect 590698 277398 590730 277634
rect 590110 241954 590730 277398
rect 590110 241718 590142 241954
rect 590378 241718 590462 241954
rect 590698 241718 590730 241954
rect 590110 241634 590730 241718
rect 590110 241398 590142 241634
rect 590378 241398 590462 241634
rect 590698 241398 590730 241634
rect 590110 205954 590730 241398
rect 590110 205718 590142 205954
rect 590378 205718 590462 205954
rect 590698 205718 590730 205954
rect 590110 205634 590730 205718
rect 590110 205398 590142 205634
rect 590378 205398 590462 205634
rect 590698 205398 590730 205634
rect 590110 169954 590730 205398
rect 590110 169718 590142 169954
rect 590378 169718 590462 169954
rect 590698 169718 590730 169954
rect 590110 169634 590730 169718
rect 590110 169398 590142 169634
rect 590378 169398 590462 169634
rect 590698 169398 590730 169634
rect 590110 133954 590730 169398
rect 590110 133718 590142 133954
rect 590378 133718 590462 133954
rect 590698 133718 590730 133954
rect 590110 133634 590730 133718
rect 590110 133398 590142 133634
rect 590378 133398 590462 133634
rect 590698 133398 590730 133634
rect 590110 97954 590730 133398
rect 590110 97718 590142 97954
rect 590378 97718 590462 97954
rect 590698 97718 590730 97954
rect 590110 97634 590730 97718
rect 590110 97398 590142 97634
rect 590378 97398 590462 97634
rect 590698 97398 590730 97634
rect 590110 61954 590730 97398
rect 590110 61718 590142 61954
rect 590378 61718 590462 61954
rect 590698 61718 590730 61954
rect 590110 61634 590730 61718
rect 590110 61398 590142 61634
rect 590378 61398 590462 61634
rect 590698 61398 590730 61634
rect 590110 25954 590730 61398
rect 590110 25718 590142 25954
rect 590378 25718 590462 25954
rect 590698 25718 590730 25954
rect 590110 25634 590730 25718
rect 590110 25398 590142 25634
rect 590378 25398 590462 25634
rect 590698 25398 590730 25634
rect 590110 -5146 590730 25398
rect 590110 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect 590110 -5466 590730 -5382
rect 590110 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect 590110 -5734 590730 -5702
rect 591070 678454 591690 710042
rect 591070 678218 591102 678454
rect 591338 678218 591422 678454
rect 591658 678218 591690 678454
rect 591070 678134 591690 678218
rect 591070 677898 591102 678134
rect 591338 677898 591422 678134
rect 591658 677898 591690 678134
rect 591070 642454 591690 677898
rect 591070 642218 591102 642454
rect 591338 642218 591422 642454
rect 591658 642218 591690 642454
rect 591070 642134 591690 642218
rect 591070 641898 591102 642134
rect 591338 641898 591422 642134
rect 591658 641898 591690 642134
rect 591070 606454 591690 641898
rect 591070 606218 591102 606454
rect 591338 606218 591422 606454
rect 591658 606218 591690 606454
rect 591070 606134 591690 606218
rect 591070 605898 591102 606134
rect 591338 605898 591422 606134
rect 591658 605898 591690 606134
rect 591070 570454 591690 605898
rect 591070 570218 591102 570454
rect 591338 570218 591422 570454
rect 591658 570218 591690 570454
rect 591070 570134 591690 570218
rect 591070 569898 591102 570134
rect 591338 569898 591422 570134
rect 591658 569898 591690 570134
rect 591070 534454 591690 569898
rect 591070 534218 591102 534454
rect 591338 534218 591422 534454
rect 591658 534218 591690 534454
rect 591070 534134 591690 534218
rect 591070 533898 591102 534134
rect 591338 533898 591422 534134
rect 591658 533898 591690 534134
rect 591070 498454 591690 533898
rect 591070 498218 591102 498454
rect 591338 498218 591422 498454
rect 591658 498218 591690 498454
rect 591070 498134 591690 498218
rect 591070 497898 591102 498134
rect 591338 497898 591422 498134
rect 591658 497898 591690 498134
rect 591070 462454 591690 497898
rect 591070 462218 591102 462454
rect 591338 462218 591422 462454
rect 591658 462218 591690 462454
rect 591070 462134 591690 462218
rect 591070 461898 591102 462134
rect 591338 461898 591422 462134
rect 591658 461898 591690 462134
rect 591070 426454 591690 461898
rect 591070 426218 591102 426454
rect 591338 426218 591422 426454
rect 591658 426218 591690 426454
rect 591070 426134 591690 426218
rect 591070 425898 591102 426134
rect 591338 425898 591422 426134
rect 591658 425898 591690 426134
rect 591070 390454 591690 425898
rect 591070 390218 591102 390454
rect 591338 390218 591422 390454
rect 591658 390218 591690 390454
rect 591070 390134 591690 390218
rect 591070 389898 591102 390134
rect 591338 389898 591422 390134
rect 591658 389898 591690 390134
rect 591070 354454 591690 389898
rect 591070 354218 591102 354454
rect 591338 354218 591422 354454
rect 591658 354218 591690 354454
rect 591070 354134 591690 354218
rect 591070 353898 591102 354134
rect 591338 353898 591422 354134
rect 591658 353898 591690 354134
rect 591070 318454 591690 353898
rect 591070 318218 591102 318454
rect 591338 318218 591422 318454
rect 591658 318218 591690 318454
rect 591070 318134 591690 318218
rect 591070 317898 591102 318134
rect 591338 317898 591422 318134
rect 591658 317898 591690 318134
rect 591070 282454 591690 317898
rect 591070 282218 591102 282454
rect 591338 282218 591422 282454
rect 591658 282218 591690 282454
rect 591070 282134 591690 282218
rect 591070 281898 591102 282134
rect 591338 281898 591422 282134
rect 591658 281898 591690 282134
rect 591070 246454 591690 281898
rect 591070 246218 591102 246454
rect 591338 246218 591422 246454
rect 591658 246218 591690 246454
rect 591070 246134 591690 246218
rect 591070 245898 591102 246134
rect 591338 245898 591422 246134
rect 591658 245898 591690 246134
rect 591070 210454 591690 245898
rect 591070 210218 591102 210454
rect 591338 210218 591422 210454
rect 591658 210218 591690 210454
rect 591070 210134 591690 210218
rect 591070 209898 591102 210134
rect 591338 209898 591422 210134
rect 591658 209898 591690 210134
rect 591070 174454 591690 209898
rect 591070 174218 591102 174454
rect 591338 174218 591422 174454
rect 591658 174218 591690 174454
rect 591070 174134 591690 174218
rect 591070 173898 591102 174134
rect 591338 173898 591422 174134
rect 591658 173898 591690 174134
rect 591070 138454 591690 173898
rect 591070 138218 591102 138454
rect 591338 138218 591422 138454
rect 591658 138218 591690 138454
rect 591070 138134 591690 138218
rect 591070 137898 591102 138134
rect 591338 137898 591422 138134
rect 591658 137898 591690 138134
rect 591070 102454 591690 137898
rect 591070 102218 591102 102454
rect 591338 102218 591422 102454
rect 591658 102218 591690 102454
rect 591070 102134 591690 102218
rect 591070 101898 591102 102134
rect 591338 101898 591422 102134
rect 591658 101898 591690 102134
rect 591070 66454 591690 101898
rect 591070 66218 591102 66454
rect 591338 66218 591422 66454
rect 591658 66218 591690 66454
rect 591070 66134 591690 66218
rect 591070 65898 591102 66134
rect 591338 65898 591422 66134
rect 591658 65898 591690 66134
rect 591070 30454 591690 65898
rect 591070 30218 591102 30454
rect 591338 30218 591422 30454
rect 591658 30218 591690 30454
rect 591070 30134 591690 30218
rect 591070 29898 591102 30134
rect 591338 29898 591422 30134
rect 591658 29898 591690 30134
rect 591070 -6106 591690 29898
rect 591070 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect 591070 -6426 591690 -6342
rect 591070 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect 591070 -6694 591690 -6662
rect 592030 682954 592650 711002
rect 592030 682718 592062 682954
rect 592298 682718 592382 682954
rect 592618 682718 592650 682954
rect 592030 682634 592650 682718
rect 592030 682398 592062 682634
rect 592298 682398 592382 682634
rect 592618 682398 592650 682634
rect 592030 646954 592650 682398
rect 592030 646718 592062 646954
rect 592298 646718 592382 646954
rect 592618 646718 592650 646954
rect 592030 646634 592650 646718
rect 592030 646398 592062 646634
rect 592298 646398 592382 646634
rect 592618 646398 592650 646634
rect 592030 610954 592650 646398
rect 592030 610718 592062 610954
rect 592298 610718 592382 610954
rect 592618 610718 592650 610954
rect 592030 610634 592650 610718
rect 592030 610398 592062 610634
rect 592298 610398 592382 610634
rect 592618 610398 592650 610634
rect 592030 574954 592650 610398
rect 592030 574718 592062 574954
rect 592298 574718 592382 574954
rect 592618 574718 592650 574954
rect 592030 574634 592650 574718
rect 592030 574398 592062 574634
rect 592298 574398 592382 574634
rect 592618 574398 592650 574634
rect 592030 538954 592650 574398
rect 592030 538718 592062 538954
rect 592298 538718 592382 538954
rect 592618 538718 592650 538954
rect 592030 538634 592650 538718
rect 592030 538398 592062 538634
rect 592298 538398 592382 538634
rect 592618 538398 592650 538634
rect 592030 502954 592650 538398
rect 592030 502718 592062 502954
rect 592298 502718 592382 502954
rect 592618 502718 592650 502954
rect 592030 502634 592650 502718
rect 592030 502398 592062 502634
rect 592298 502398 592382 502634
rect 592618 502398 592650 502634
rect 592030 466954 592650 502398
rect 592030 466718 592062 466954
rect 592298 466718 592382 466954
rect 592618 466718 592650 466954
rect 592030 466634 592650 466718
rect 592030 466398 592062 466634
rect 592298 466398 592382 466634
rect 592618 466398 592650 466634
rect 592030 430954 592650 466398
rect 592030 430718 592062 430954
rect 592298 430718 592382 430954
rect 592618 430718 592650 430954
rect 592030 430634 592650 430718
rect 592030 430398 592062 430634
rect 592298 430398 592382 430634
rect 592618 430398 592650 430634
rect 592030 394954 592650 430398
rect 592030 394718 592062 394954
rect 592298 394718 592382 394954
rect 592618 394718 592650 394954
rect 592030 394634 592650 394718
rect 592030 394398 592062 394634
rect 592298 394398 592382 394634
rect 592618 394398 592650 394634
rect 592030 358954 592650 394398
rect 592030 358718 592062 358954
rect 592298 358718 592382 358954
rect 592618 358718 592650 358954
rect 592030 358634 592650 358718
rect 592030 358398 592062 358634
rect 592298 358398 592382 358634
rect 592618 358398 592650 358634
rect 592030 322954 592650 358398
rect 592030 322718 592062 322954
rect 592298 322718 592382 322954
rect 592618 322718 592650 322954
rect 592030 322634 592650 322718
rect 592030 322398 592062 322634
rect 592298 322398 592382 322634
rect 592618 322398 592650 322634
rect 592030 286954 592650 322398
rect 592030 286718 592062 286954
rect 592298 286718 592382 286954
rect 592618 286718 592650 286954
rect 592030 286634 592650 286718
rect 592030 286398 592062 286634
rect 592298 286398 592382 286634
rect 592618 286398 592650 286634
rect 592030 250954 592650 286398
rect 592030 250718 592062 250954
rect 592298 250718 592382 250954
rect 592618 250718 592650 250954
rect 592030 250634 592650 250718
rect 592030 250398 592062 250634
rect 592298 250398 592382 250634
rect 592618 250398 592650 250634
rect 592030 214954 592650 250398
rect 592030 214718 592062 214954
rect 592298 214718 592382 214954
rect 592618 214718 592650 214954
rect 592030 214634 592650 214718
rect 592030 214398 592062 214634
rect 592298 214398 592382 214634
rect 592618 214398 592650 214634
rect 592030 178954 592650 214398
rect 592030 178718 592062 178954
rect 592298 178718 592382 178954
rect 592618 178718 592650 178954
rect 592030 178634 592650 178718
rect 592030 178398 592062 178634
rect 592298 178398 592382 178634
rect 592618 178398 592650 178634
rect 592030 142954 592650 178398
rect 592030 142718 592062 142954
rect 592298 142718 592382 142954
rect 592618 142718 592650 142954
rect 592030 142634 592650 142718
rect 592030 142398 592062 142634
rect 592298 142398 592382 142634
rect 592618 142398 592650 142634
rect 592030 106954 592650 142398
rect 592030 106718 592062 106954
rect 592298 106718 592382 106954
rect 592618 106718 592650 106954
rect 592030 106634 592650 106718
rect 592030 106398 592062 106634
rect 592298 106398 592382 106634
rect 592618 106398 592650 106634
rect 592030 70954 592650 106398
rect 592030 70718 592062 70954
rect 592298 70718 592382 70954
rect 592618 70718 592650 70954
rect 592030 70634 592650 70718
rect 592030 70398 592062 70634
rect 592298 70398 592382 70634
rect 592618 70398 592650 70634
rect 592030 34954 592650 70398
rect 592030 34718 592062 34954
rect 592298 34718 592382 34954
rect 592618 34718 592650 34954
rect 592030 34634 592650 34718
rect 592030 34398 592062 34634
rect 592298 34398 592382 34634
rect 592618 34398 592650 34634
rect 592030 -7066 592650 34398
rect 592030 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect 592030 -7386 592650 -7302
rect 592030 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect 592030 -7654 592650 -7622
<< via4 >>
rect -8694 711322 -8458 711558
rect -8374 711322 -8138 711558
rect -8694 711002 -8458 711238
rect -8374 711002 -8138 711238
rect -8694 682718 -8458 682954
rect -8374 682718 -8138 682954
rect -8694 682398 -8458 682634
rect -8374 682398 -8138 682634
rect -8694 646718 -8458 646954
rect -8374 646718 -8138 646954
rect -8694 646398 -8458 646634
rect -8374 646398 -8138 646634
rect -8694 610718 -8458 610954
rect -8374 610718 -8138 610954
rect -8694 610398 -8458 610634
rect -8374 610398 -8138 610634
rect -8694 574718 -8458 574954
rect -8374 574718 -8138 574954
rect -8694 574398 -8458 574634
rect -8374 574398 -8138 574634
rect -8694 538718 -8458 538954
rect -8374 538718 -8138 538954
rect -8694 538398 -8458 538634
rect -8374 538398 -8138 538634
rect -8694 502718 -8458 502954
rect -8374 502718 -8138 502954
rect -8694 502398 -8458 502634
rect -8374 502398 -8138 502634
rect -8694 466718 -8458 466954
rect -8374 466718 -8138 466954
rect -8694 466398 -8458 466634
rect -8374 466398 -8138 466634
rect -8694 430718 -8458 430954
rect -8374 430718 -8138 430954
rect -8694 430398 -8458 430634
rect -8374 430398 -8138 430634
rect -8694 394718 -8458 394954
rect -8374 394718 -8138 394954
rect -8694 394398 -8458 394634
rect -8374 394398 -8138 394634
rect -8694 358718 -8458 358954
rect -8374 358718 -8138 358954
rect -8694 358398 -8458 358634
rect -8374 358398 -8138 358634
rect -8694 322718 -8458 322954
rect -8374 322718 -8138 322954
rect -8694 322398 -8458 322634
rect -8374 322398 -8138 322634
rect -8694 286718 -8458 286954
rect -8374 286718 -8138 286954
rect -8694 286398 -8458 286634
rect -8374 286398 -8138 286634
rect -8694 250718 -8458 250954
rect -8374 250718 -8138 250954
rect -8694 250398 -8458 250634
rect -8374 250398 -8138 250634
rect -8694 214718 -8458 214954
rect -8374 214718 -8138 214954
rect -8694 214398 -8458 214634
rect -8374 214398 -8138 214634
rect -8694 178718 -8458 178954
rect -8374 178718 -8138 178954
rect -8694 178398 -8458 178634
rect -8374 178398 -8138 178634
rect -8694 142718 -8458 142954
rect -8374 142718 -8138 142954
rect -8694 142398 -8458 142634
rect -8374 142398 -8138 142634
rect -8694 106718 -8458 106954
rect -8374 106718 -8138 106954
rect -8694 106398 -8458 106634
rect -8374 106398 -8138 106634
rect -8694 70718 -8458 70954
rect -8374 70718 -8138 70954
rect -8694 70398 -8458 70634
rect -8374 70398 -8138 70634
rect -8694 34718 -8458 34954
rect -8374 34718 -8138 34954
rect -8694 34398 -8458 34634
rect -8374 34398 -8138 34634
rect -7734 710362 -7498 710598
rect -7414 710362 -7178 710598
rect -7734 710042 -7498 710278
rect -7414 710042 -7178 710278
rect -7734 678218 -7498 678454
rect -7414 678218 -7178 678454
rect -7734 677898 -7498 678134
rect -7414 677898 -7178 678134
rect -7734 642218 -7498 642454
rect -7414 642218 -7178 642454
rect -7734 641898 -7498 642134
rect -7414 641898 -7178 642134
rect -7734 606218 -7498 606454
rect -7414 606218 -7178 606454
rect -7734 605898 -7498 606134
rect -7414 605898 -7178 606134
rect -7734 570218 -7498 570454
rect -7414 570218 -7178 570454
rect -7734 569898 -7498 570134
rect -7414 569898 -7178 570134
rect -7734 534218 -7498 534454
rect -7414 534218 -7178 534454
rect -7734 533898 -7498 534134
rect -7414 533898 -7178 534134
rect -7734 498218 -7498 498454
rect -7414 498218 -7178 498454
rect -7734 497898 -7498 498134
rect -7414 497898 -7178 498134
rect -7734 462218 -7498 462454
rect -7414 462218 -7178 462454
rect -7734 461898 -7498 462134
rect -7414 461898 -7178 462134
rect -7734 426218 -7498 426454
rect -7414 426218 -7178 426454
rect -7734 425898 -7498 426134
rect -7414 425898 -7178 426134
rect -7734 390218 -7498 390454
rect -7414 390218 -7178 390454
rect -7734 389898 -7498 390134
rect -7414 389898 -7178 390134
rect -7734 354218 -7498 354454
rect -7414 354218 -7178 354454
rect -7734 353898 -7498 354134
rect -7414 353898 -7178 354134
rect -7734 318218 -7498 318454
rect -7414 318218 -7178 318454
rect -7734 317898 -7498 318134
rect -7414 317898 -7178 318134
rect -7734 282218 -7498 282454
rect -7414 282218 -7178 282454
rect -7734 281898 -7498 282134
rect -7414 281898 -7178 282134
rect -7734 246218 -7498 246454
rect -7414 246218 -7178 246454
rect -7734 245898 -7498 246134
rect -7414 245898 -7178 246134
rect -7734 210218 -7498 210454
rect -7414 210218 -7178 210454
rect -7734 209898 -7498 210134
rect -7414 209898 -7178 210134
rect -7734 174218 -7498 174454
rect -7414 174218 -7178 174454
rect -7734 173898 -7498 174134
rect -7414 173898 -7178 174134
rect -7734 138218 -7498 138454
rect -7414 138218 -7178 138454
rect -7734 137898 -7498 138134
rect -7414 137898 -7178 138134
rect -7734 102218 -7498 102454
rect -7414 102218 -7178 102454
rect -7734 101898 -7498 102134
rect -7414 101898 -7178 102134
rect -7734 66218 -7498 66454
rect -7414 66218 -7178 66454
rect -7734 65898 -7498 66134
rect -7414 65898 -7178 66134
rect -7734 30218 -7498 30454
rect -7414 30218 -7178 30454
rect -7734 29898 -7498 30134
rect -7414 29898 -7178 30134
rect -6774 709402 -6538 709638
rect -6454 709402 -6218 709638
rect -6774 709082 -6538 709318
rect -6454 709082 -6218 709318
rect -6774 673718 -6538 673954
rect -6454 673718 -6218 673954
rect -6774 673398 -6538 673634
rect -6454 673398 -6218 673634
rect -6774 637718 -6538 637954
rect -6454 637718 -6218 637954
rect -6774 637398 -6538 637634
rect -6454 637398 -6218 637634
rect -6774 601718 -6538 601954
rect -6454 601718 -6218 601954
rect -6774 601398 -6538 601634
rect -6454 601398 -6218 601634
rect -6774 565718 -6538 565954
rect -6454 565718 -6218 565954
rect -6774 565398 -6538 565634
rect -6454 565398 -6218 565634
rect -6774 529718 -6538 529954
rect -6454 529718 -6218 529954
rect -6774 529398 -6538 529634
rect -6454 529398 -6218 529634
rect -6774 493718 -6538 493954
rect -6454 493718 -6218 493954
rect -6774 493398 -6538 493634
rect -6454 493398 -6218 493634
rect -6774 457718 -6538 457954
rect -6454 457718 -6218 457954
rect -6774 457398 -6538 457634
rect -6454 457398 -6218 457634
rect -6774 421718 -6538 421954
rect -6454 421718 -6218 421954
rect -6774 421398 -6538 421634
rect -6454 421398 -6218 421634
rect -6774 385718 -6538 385954
rect -6454 385718 -6218 385954
rect -6774 385398 -6538 385634
rect -6454 385398 -6218 385634
rect -6774 349718 -6538 349954
rect -6454 349718 -6218 349954
rect -6774 349398 -6538 349634
rect -6454 349398 -6218 349634
rect -6774 313718 -6538 313954
rect -6454 313718 -6218 313954
rect -6774 313398 -6538 313634
rect -6454 313398 -6218 313634
rect -6774 277718 -6538 277954
rect -6454 277718 -6218 277954
rect -6774 277398 -6538 277634
rect -6454 277398 -6218 277634
rect -6774 241718 -6538 241954
rect -6454 241718 -6218 241954
rect -6774 241398 -6538 241634
rect -6454 241398 -6218 241634
rect -6774 205718 -6538 205954
rect -6454 205718 -6218 205954
rect -6774 205398 -6538 205634
rect -6454 205398 -6218 205634
rect -6774 169718 -6538 169954
rect -6454 169718 -6218 169954
rect -6774 169398 -6538 169634
rect -6454 169398 -6218 169634
rect -6774 133718 -6538 133954
rect -6454 133718 -6218 133954
rect -6774 133398 -6538 133634
rect -6454 133398 -6218 133634
rect -6774 97718 -6538 97954
rect -6454 97718 -6218 97954
rect -6774 97398 -6538 97634
rect -6454 97398 -6218 97634
rect -6774 61718 -6538 61954
rect -6454 61718 -6218 61954
rect -6774 61398 -6538 61634
rect -6454 61398 -6218 61634
rect -6774 25718 -6538 25954
rect -6454 25718 -6218 25954
rect -6774 25398 -6538 25634
rect -6454 25398 -6218 25634
rect -5814 708442 -5578 708678
rect -5494 708442 -5258 708678
rect -5814 708122 -5578 708358
rect -5494 708122 -5258 708358
rect -5814 669218 -5578 669454
rect -5494 669218 -5258 669454
rect -5814 668898 -5578 669134
rect -5494 668898 -5258 669134
rect -5814 633218 -5578 633454
rect -5494 633218 -5258 633454
rect -5814 632898 -5578 633134
rect -5494 632898 -5258 633134
rect -5814 597218 -5578 597454
rect -5494 597218 -5258 597454
rect -5814 596898 -5578 597134
rect -5494 596898 -5258 597134
rect -5814 561218 -5578 561454
rect -5494 561218 -5258 561454
rect -5814 560898 -5578 561134
rect -5494 560898 -5258 561134
rect -5814 525218 -5578 525454
rect -5494 525218 -5258 525454
rect -5814 524898 -5578 525134
rect -5494 524898 -5258 525134
rect -5814 489218 -5578 489454
rect -5494 489218 -5258 489454
rect -5814 488898 -5578 489134
rect -5494 488898 -5258 489134
rect -5814 453218 -5578 453454
rect -5494 453218 -5258 453454
rect -5814 452898 -5578 453134
rect -5494 452898 -5258 453134
rect -5814 417218 -5578 417454
rect -5494 417218 -5258 417454
rect -5814 416898 -5578 417134
rect -5494 416898 -5258 417134
rect -5814 381218 -5578 381454
rect -5494 381218 -5258 381454
rect -5814 380898 -5578 381134
rect -5494 380898 -5258 381134
rect -5814 345218 -5578 345454
rect -5494 345218 -5258 345454
rect -5814 344898 -5578 345134
rect -5494 344898 -5258 345134
rect -5814 309218 -5578 309454
rect -5494 309218 -5258 309454
rect -5814 308898 -5578 309134
rect -5494 308898 -5258 309134
rect -5814 273218 -5578 273454
rect -5494 273218 -5258 273454
rect -5814 272898 -5578 273134
rect -5494 272898 -5258 273134
rect -5814 237218 -5578 237454
rect -5494 237218 -5258 237454
rect -5814 236898 -5578 237134
rect -5494 236898 -5258 237134
rect -5814 201218 -5578 201454
rect -5494 201218 -5258 201454
rect -5814 200898 -5578 201134
rect -5494 200898 -5258 201134
rect -5814 165218 -5578 165454
rect -5494 165218 -5258 165454
rect -5814 164898 -5578 165134
rect -5494 164898 -5258 165134
rect -5814 129218 -5578 129454
rect -5494 129218 -5258 129454
rect -5814 128898 -5578 129134
rect -5494 128898 -5258 129134
rect -5814 93218 -5578 93454
rect -5494 93218 -5258 93454
rect -5814 92898 -5578 93134
rect -5494 92898 -5258 93134
rect -5814 57218 -5578 57454
rect -5494 57218 -5258 57454
rect -5814 56898 -5578 57134
rect -5494 56898 -5258 57134
rect -5814 21218 -5578 21454
rect -5494 21218 -5258 21454
rect -5814 20898 -5578 21134
rect -5494 20898 -5258 21134
rect -4854 707482 -4618 707718
rect -4534 707482 -4298 707718
rect -4854 707162 -4618 707398
rect -4534 707162 -4298 707398
rect -4854 700718 -4618 700954
rect -4534 700718 -4298 700954
rect -4854 700398 -4618 700634
rect -4534 700398 -4298 700634
rect -4854 664718 -4618 664954
rect -4534 664718 -4298 664954
rect -4854 664398 -4618 664634
rect -4534 664398 -4298 664634
rect -4854 628718 -4618 628954
rect -4534 628718 -4298 628954
rect -4854 628398 -4618 628634
rect -4534 628398 -4298 628634
rect -4854 592718 -4618 592954
rect -4534 592718 -4298 592954
rect -4854 592398 -4618 592634
rect -4534 592398 -4298 592634
rect -4854 556718 -4618 556954
rect -4534 556718 -4298 556954
rect -4854 556398 -4618 556634
rect -4534 556398 -4298 556634
rect -4854 520718 -4618 520954
rect -4534 520718 -4298 520954
rect -4854 520398 -4618 520634
rect -4534 520398 -4298 520634
rect -4854 484718 -4618 484954
rect -4534 484718 -4298 484954
rect -4854 484398 -4618 484634
rect -4534 484398 -4298 484634
rect -4854 448718 -4618 448954
rect -4534 448718 -4298 448954
rect -4854 448398 -4618 448634
rect -4534 448398 -4298 448634
rect -4854 412718 -4618 412954
rect -4534 412718 -4298 412954
rect -4854 412398 -4618 412634
rect -4534 412398 -4298 412634
rect -4854 376718 -4618 376954
rect -4534 376718 -4298 376954
rect -4854 376398 -4618 376634
rect -4534 376398 -4298 376634
rect -4854 340718 -4618 340954
rect -4534 340718 -4298 340954
rect -4854 340398 -4618 340634
rect -4534 340398 -4298 340634
rect -4854 304718 -4618 304954
rect -4534 304718 -4298 304954
rect -4854 304398 -4618 304634
rect -4534 304398 -4298 304634
rect -4854 268718 -4618 268954
rect -4534 268718 -4298 268954
rect -4854 268398 -4618 268634
rect -4534 268398 -4298 268634
rect -4854 232718 -4618 232954
rect -4534 232718 -4298 232954
rect -4854 232398 -4618 232634
rect -4534 232398 -4298 232634
rect -4854 196718 -4618 196954
rect -4534 196718 -4298 196954
rect -4854 196398 -4618 196634
rect -4534 196398 -4298 196634
rect -4854 160718 -4618 160954
rect -4534 160718 -4298 160954
rect -4854 160398 -4618 160634
rect -4534 160398 -4298 160634
rect -4854 124718 -4618 124954
rect -4534 124718 -4298 124954
rect -4854 124398 -4618 124634
rect -4534 124398 -4298 124634
rect -4854 88718 -4618 88954
rect -4534 88718 -4298 88954
rect -4854 88398 -4618 88634
rect -4534 88398 -4298 88634
rect -4854 52718 -4618 52954
rect -4534 52718 -4298 52954
rect -4854 52398 -4618 52634
rect -4534 52398 -4298 52634
rect -4854 16718 -4618 16954
rect -4534 16718 -4298 16954
rect -4854 16398 -4618 16634
rect -4534 16398 -4298 16634
rect -3894 706522 -3658 706758
rect -3574 706522 -3338 706758
rect -3894 706202 -3658 706438
rect -3574 706202 -3338 706438
rect -3894 696218 -3658 696454
rect -3574 696218 -3338 696454
rect -3894 695898 -3658 696134
rect -3574 695898 -3338 696134
rect -3894 660218 -3658 660454
rect -3574 660218 -3338 660454
rect -3894 659898 -3658 660134
rect -3574 659898 -3338 660134
rect -3894 624218 -3658 624454
rect -3574 624218 -3338 624454
rect -3894 623898 -3658 624134
rect -3574 623898 -3338 624134
rect -3894 588218 -3658 588454
rect -3574 588218 -3338 588454
rect -3894 587898 -3658 588134
rect -3574 587898 -3338 588134
rect -3894 552218 -3658 552454
rect -3574 552218 -3338 552454
rect -3894 551898 -3658 552134
rect -3574 551898 -3338 552134
rect -3894 516218 -3658 516454
rect -3574 516218 -3338 516454
rect -3894 515898 -3658 516134
rect -3574 515898 -3338 516134
rect -3894 480218 -3658 480454
rect -3574 480218 -3338 480454
rect -3894 479898 -3658 480134
rect -3574 479898 -3338 480134
rect -3894 444218 -3658 444454
rect -3574 444218 -3338 444454
rect -3894 443898 -3658 444134
rect -3574 443898 -3338 444134
rect -3894 408218 -3658 408454
rect -3574 408218 -3338 408454
rect -3894 407898 -3658 408134
rect -3574 407898 -3338 408134
rect -3894 372218 -3658 372454
rect -3574 372218 -3338 372454
rect -3894 371898 -3658 372134
rect -3574 371898 -3338 372134
rect -3894 336218 -3658 336454
rect -3574 336218 -3338 336454
rect -3894 335898 -3658 336134
rect -3574 335898 -3338 336134
rect -3894 300218 -3658 300454
rect -3574 300218 -3338 300454
rect -3894 299898 -3658 300134
rect -3574 299898 -3338 300134
rect -3894 264218 -3658 264454
rect -3574 264218 -3338 264454
rect -3894 263898 -3658 264134
rect -3574 263898 -3338 264134
rect -3894 228218 -3658 228454
rect -3574 228218 -3338 228454
rect -3894 227898 -3658 228134
rect -3574 227898 -3338 228134
rect -3894 192218 -3658 192454
rect -3574 192218 -3338 192454
rect -3894 191898 -3658 192134
rect -3574 191898 -3338 192134
rect -3894 156218 -3658 156454
rect -3574 156218 -3338 156454
rect -3894 155898 -3658 156134
rect -3574 155898 -3338 156134
rect -3894 120218 -3658 120454
rect -3574 120218 -3338 120454
rect -3894 119898 -3658 120134
rect -3574 119898 -3338 120134
rect -3894 84218 -3658 84454
rect -3574 84218 -3338 84454
rect -3894 83898 -3658 84134
rect -3574 83898 -3338 84134
rect -3894 48218 -3658 48454
rect -3574 48218 -3338 48454
rect -3894 47898 -3658 48134
rect -3574 47898 -3338 48134
rect -3894 12218 -3658 12454
rect -3574 12218 -3338 12454
rect -3894 11898 -3658 12134
rect -3574 11898 -3338 12134
rect -2934 705562 -2698 705798
rect -2614 705562 -2378 705798
rect -2934 705242 -2698 705478
rect -2614 705242 -2378 705478
rect -2934 691718 -2698 691954
rect -2614 691718 -2378 691954
rect -2934 691398 -2698 691634
rect -2614 691398 -2378 691634
rect -2934 655718 -2698 655954
rect -2614 655718 -2378 655954
rect -2934 655398 -2698 655634
rect -2614 655398 -2378 655634
rect -2934 619718 -2698 619954
rect -2614 619718 -2378 619954
rect -2934 619398 -2698 619634
rect -2614 619398 -2378 619634
rect -2934 583718 -2698 583954
rect -2614 583718 -2378 583954
rect -2934 583398 -2698 583634
rect -2614 583398 -2378 583634
rect -2934 547718 -2698 547954
rect -2614 547718 -2378 547954
rect -2934 547398 -2698 547634
rect -2614 547398 -2378 547634
rect -2934 511718 -2698 511954
rect -2614 511718 -2378 511954
rect -2934 511398 -2698 511634
rect -2614 511398 -2378 511634
rect -2934 475718 -2698 475954
rect -2614 475718 -2378 475954
rect -2934 475398 -2698 475634
rect -2614 475398 -2378 475634
rect -2934 439718 -2698 439954
rect -2614 439718 -2378 439954
rect -2934 439398 -2698 439634
rect -2614 439398 -2378 439634
rect -2934 403718 -2698 403954
rect -2614 403718 -2378 403954
rect -2934 403398 -2698 403634
rect -2614 403398 -2378 403634
rect -2934 367718 -2698 367954
rect -2614 367718 -2378 367954
rect -2934 367398 -2698 367634
rect -2614 367398 -2378 367634
rect -2934 331718 -2698 331954
rect -2614 331718 -2378 331954
rect -2934 331398 -2698 331634
rect -2614 331398 -2378 331634
rect -2934 295718 -2698 295954
rect -2614 295718 -2378 295954
rect -2934 295398 -2698 295634
rect -2614 295398 -2378 295634
rect -2934 259718 -2698 259954
rect -2614 259718 -2378 259954
rect -2934 259398 -2698 259634
rect -2614 259398 -2378 259634
rect -2934 223718 -2698 223954
rect -2614 223718 -2378 223954
rect -2934 223398 -2698 223634
rect -2614 223398 -2378 223634
rect -2934 187718 -2698 187954
rect -2614 187718 -2378 187954
rect -2934 187398 -2698 187634
rect -2614 187398 -2378 187634
rect -2934 151718 -2698 151954
rect -2614 151718 -2378 151954
rect -2934 151398 -2698 151634
rect -2614 151398 -2378 151634
rect -2934 115718 -2698 115954
rect -2614 115718 -2378 115954
rect -2934 115398 -2698 115634
rect -2614 115398 -2378 115634
rect -2934 79718 -2698 79954
rect -2614 79718 -2378 79954
rect -2934 79398 -2698 79634
rect -2614 79398 -2378 79634
rect -2934 43718 -2698 43954
rect -2614 43718 -2378 43954
rect -2934 43398 -2698 43634
rect -2614 43398 -2378 43634
rect -2934 7718 -2698 7954
rect -2614 7718 -2378 7954
rect -2934 7398 -2698 7634
rect -2614 7398 -2378 7634
rect -1974 704602 -1738 704838
rect -1654 704602 -1418 704838
rect -1974 704282 -1738 704518
rect -1654 704282 -1418 704518
rect -1974 687218 -1738 687454
rect -1654 687218 -1418 687454
rect -1974 686898 -1738 687134
rect -1654 686898 -1418 687134
rect -1974 651218 -1738 651454
rect -1654 651218 -1418 651454
rect -1974 650898 -1738 651134
rect -1654 650898 -1418 651134
rect -1974 615218 -1738 615454
rect -1654 615218 -1418 615454
rect -1974 614898 -1738 615134
rect -1654 614898 -1418 615134
rect -1974 579218 -1738 579454
rect -1654 579218 -1418 579454
rect -1974 578898 -1738 579134
rect -1654 578898 -1418 579134
rect -1974 543218 -1738 543454
rect -1654 543218 -1418 543454
rect -1974 542898 -1738 543134
rect -1654 542898 -1418 543134
rect -1974 507218 -1738 507454
rect -1654 507218 -1418 507454
rect -1974 506898 -1738 507134
rect -1654 506898 -1418 507134
rect -1974 471218 -1738 471454
rect -1654 471218 -1418 471454
rect -1974 470898 -1738 471134
rect -1654 470898 -1418 471134
rect -1974 435218 -1738 435454
rect -1654 435218 -1418 435454
rect -1974 434898 -1738 435134
rect -1654 434898 -1418 435134
rect -1974 399218 -1738 399454
rect -1654 399218 -1418 399454
rect -1974 398898 -1738 399134
rect -1654 398898 -1418 399134
rect -1974 363218 -1738 363454
rect -1654 363218 -1418 363454
rect -1974 362898 -1738 363134
rect -1654 362898 -1418 363134
rect -1974 327218 -1738 327454
rect -1654 327218 -1418 327454
rect -1974 326898 -1738 327134
rect -1654 326898 -1418 327134
rect -1974 291218 -1738 291454
rect -1654 291218 -1418 291454
rect -1974 290898 -1738 291134
rect -1654 290898 -1418 291134
rect -1974 255218 -1738 255454
rect -1654 255218 -1418 255454
rect -1974 254898 -1738 255134
rect -1654 254898 -1418 255134
rect -1974 219218 -1738 219454
rect -1654 219218 -1418 219454
rect -1974 218898 -1738 219134
rect -1654 218898 -1418 219134
rect -1974 183218 -1738 183454
rect -1654 183218 -1418 183454
rect -1974 182898 -1738 183134
rect -1654 182898 -1418 183134
rect -1974 147218 -1738 147454
rect -1654 147218 -1418 147454
rect -1974 146898 -1738 147134
rect -1654 146898 -1418 147134
rect -1974 111218 -1738 111454
rect -1654 111218 -1418 111454
rect -1974 110898 -1738 111134
rect -1654 110898 -1418 111134
rect -1974 75218 -1738 75454
rect -1654 75218 -1418 75454
rect -1974 74898 -1738 75134
rect -1654 74898 -1418 75134
rect -1974 39218 -1738 39454
rect -1654 39218 -1418 39454
rect -1974 38898 -1738 39134
rect -1654 38898 -1418 39134
rect -1974 3218 -1738 3454
rect -1654 3218 -1418 3454
rect -1974 2898 -1738 3134
rect -1654 2898 -1418 3134
rect -1974 -582 -1738 -346
rect -1654 -582 -1418 -346
rect -1974 -902 -1738 -666
rect -1654 -902 -1418 -666
rect 1826 704602 2062 704838
rect 2146 704602 2382 704838
rect 1826 704282 2062 704518
rect 2146 704282 2382 704518
rect 1826 687218 2062 687454
rect 2146 687218 2382 687454
rect 1826 686898 2062 687134
rect 2146 686898 2382 687134
rect 1826 651218 2062 651454
rect 2146 651218 2382 651454
rect 1826 650898 2062 651134
rect 2146 650898 2382 651134
rect 1826 615218 2062 615454
rect 2146 615218 2382 615454
rect 1826 614898 2062 615134
rect 2146 614898 2382 615134
rect 1826 579218 2062 579454
rect 2146 579218 2382 579454
rect 1826 578898 2062 579134
rect 2146 578898 2382 579134
rect 1826 543218 2062 543454
rect 2146 543218 2382 543454
rect 1826 542898 2062 543134
rect 2146 542898 2382 543134
rect 1826 507218 2062 507454
rect 2146 507218 2382 507454
rect 1826 506898 2062 507134
rect 2146 506898 2382 507134
rect 1826 471218 2062 471454
rect 2146 471218 2382 471454
rect 1826 470898 2062 471134
rect 2146 470898 2382 471134
rect 1826 435218 2062 435454
rect 2146 435218 2382 435454
rect 1826 434898 2062 435134
rect 2146 434898 2382 435134
rect 1826 399218 2062 399454
rect 2146 399218 2382 399454
rect 1826 398898 2062 399134
rect 2146 398898 2382 399134
rect 1826 363218 2062 363454
rect 2146 363218 2382 363454
rect 1826 362898 2062 363134
rect 2146 362898 2382 363134
rect 1826 327218 2062 327454
rect 2146 327218 2382 327454
rect 1826 326898 2062 327134
rect 2146 326898 2382 327134
rect 1826 291218 2062 291454
rect 2146 291218 2382 291454
rect 1826 290898 2062 291134
rect 2146 290898 2382 291134
rect 1826 255218 2062 255454
rect 2146 255218 2382 255454
rect 1826 254898 2062 255134
rect 2146 254898 2382 255134
rect 1826 219218 2062 219454
rect 2146 219218 2382 219454
rect 1826 218898 2062 219134
rect 2146 218898 2382 219134
rect 1826 183218 2062 183454
rect 2146 183218 2382 183454
rect 1826 182898 2062 183134
rect 2146 182898 2382 183134
rect 1826 147218 2062 147454
rect 2146 147218 2382 147454
rect 1826 146898 2062 147134
rect 2146 146898 2382 147134
rect 1826 111218 2062 111454
rect 2146 111218 2382 111454
rect 1826 110898 2062 111134
rect 2146 110898 2382 111134
rect 1826 75218 2062 75454
rect 2146 75218 2382 75454
rect 1826 74898 2062 75134
rect 2146 74898 2382 75134
rect 1826 39218 2062 39454
rect 2146 39218 2382 39454
rect 1826 38898 2062 39134
rect 2146 38898 2382 39134
rect 1826 3218 2062 3454
rect 2146 3218 2382 3454
rect 1826 2898 2062 3134
rect 2146 2898 2382 3134
rect 1826 -582 2062 -346
rect 2146 -582 2382 -346
rect 1826 -902 2062 -666
rect 2146 -902 2382 -666
rect -2934 -1542 -2698 -1306
rect -2614 -1542 -2378 -1306
rect -2934 -1862 -2698 -1626
rect -2614 -1862 -2378 -1626
rect -3894 -2502 -3658 -2266
rect -3574 -2502 -3338 -2266
rect -3894 -2822 -3658 -2586
rect -3574 -2822 -3338 -2586
rect -4854 -3462 -4618 -3226
rect -4534 -3462 -4298 -3226
rect -4854 -3782 -4618 -3546
rect -4534 -3782 -4298 -3546
rect -5814 -4422 -5578 -4186
rect -5494 -4422 -5258 -4186
rect -5814 -4742 -5578 -4506
rect -5494 -4742 -5258 -4506
rect -6774 -5382 -6538 -5146
rect -6454 -5382 -6218 -5146
rect -6774 -5702 -6538 -5466
rect -6454 -5702 -6218 -5466
rect -7734 -6342 -7498 -6106
rect -7414 -6342 -7178 -6106
rect -7734 -6662 -7498 -6426
rect -7414 -6662 -7178 -6426
rect -8694 -7302 -8458 -7066
rect -8374 -7302 -8138 -7066
rect -8694 -7622 -8458 -7386
rect -8374 -7622 -8138 -7386
rect 6326 705562 6562 705798
rect 6646 705562 6882 705798
rect 6326 705242 6562 705478
rect 6646 705242 6882 705478
rect 6326 691718 6562 691954
rect 6646 691718 6882 691954
rect 6326 691398 6562 691634
rect 6646 691398 6882 691634
rect 6326 655718 6562 655954
rect 6646 655718 6882 655954
rect 6326 655398 6562 655634
rect 6646 655398 6882 655634
rect 6326 619718 6562 619954
rect 6646 619718 6882 619954
rect 6326 619398 6562 619634
rect 6646 619398 6882 619634
rect 6326 583718 6562 583954
rect 6646 583718 6882 583954
rect 6326 583398 6562 583634
rect 6646 583398 6882 583634
rect 6326 547718 6562 547954
rect 6646 547718 6882 547954
rect 6326 547398 6562 547634
rect 6646 547398 6882 547634
rect 6326 511718 6562 511954
rect 6646 511718 6882 511954
rect 6326 511398 6562 511634
rect 6646 511398 6882 511634
rect 6326 475718 6562 475954
rect 6646 475718 6882 475954
rect 6326 475398 6562 475634
rect 6646 475398 6882 475634
rect 6326 439718 6562 439954
rect 6646 439718 6882 439954
rect 6326 439398 6562 439634
rect 6646 439398 6882 439634
rect 6326 403718 6562 403954
rect 6646 403718 6882 403954
rect 6326 403398 6562 403634
rect 6646 403398 6882 403634
rect 6326 367718 6562 367954
rect 6646 367718 6882 367954
rect 6326 367398 6562 367634
rect 6646 367398 6882 367634
rect 6326 331718 6562 331954
rect 6646 331718 6882 331954
rect 6326 331398 6562 331634
rect 6646 331398 6882 331634
rect 6326 295718 6562 295954
rect 6646 295718 6882 295954
rect 6326 295398 6562 295634
rect 6646 295398 6882 295634
rect 6326 259718 6562 259954
rect 6646 259718 6882 259954
rect 6326 259398 6562 259634
rect 6646 259398 6882 259634
rect 6326 223718 6562 223954
rect 6646 223718 6882 223954
rect 6326 223398 6562 223634
rect 6646 223398 6882 223634
rect 6326 187718 6562 187954
rect 6646 187718 6882 187954
rect 6326 187398 6562 187634
rect 6646 187398 6882 187634
rect 6326 151718 6562 151954
rect 6646 151718 6882 151954
rect 6326 151398 6562 151634
rect 6646 151398 6882 151634
rect 6326 115718 6562 115954
rect 6646 115718 6882 115954
rect 6326 115398 6562 115634
rect 6646 115398 6882 115634
rect 6326 79718 6562 79954
rect 6646 79718 6882 79954
rect 6326 79398 6562 79634
rect 6646 79398 6882 79634
rect 6326 43718 6562 43954
rect 6646 43718 6882 43954
rect 6326 43398 6562 43634
rect 6646 43398 6882 43634
rect 6326 7718 6562 7954
rect 6646 7718 6882 7954
rect 6326 7398 6562 7634
rect 6646 7398 6882 7634
rect 6326 -1542 6562 -1306
rect 6646 -1542 6882 -1306
rect 6326 -1862 6562 -1626
rect 6646 -1862 6882 -1626
rect 10826 706522 11062 706758
rect 11146 706522 11382 706758
rect 10826 706202 11062 706438
rect 11146 706202 11382 706438
rect 10826 696218 11062 696454
rect 11146 696218 11382 696454
rect 10826 695898 11062 696134
rect 11146 695898 11382 696134
rect 10826 660218 11062 660454
rect 11146 660218 11382 660454
rect 10826 659898 11062 660134
rect 11146 659898 11382 660134
rect 10826 624218 11062 624454
rect 11146 624218 11382 624454
rect 10826 623898 11062 624134
rect 11146 623898 11382 624134
rect 10826 588218 11062 588454
rect 11146 588218 11382 588454
rect 10826 587898 11062 588134
rect 11146 587898 11382 588134
rect 10826 552218 11062 552454
rect 11146 552218 11382 552454
rect 10826 551898 11062 552134
rect 11146 551898 11382 552134
rect 10826 516218 11062 516454
rect 11146 516218 11382 516454
rect 10826 515898 11062 516134
rect 11146 515898 11382 516134
rect 10826 480218 11062 480454
rect 11146 480218 11382 480454
rect 10826 479898 11062 480134
rect 11146 479898 11382 480134
rect 10826 444218 11062 444454
rect 11146 444218 11382 444454
rect 10826 443898 11062 444134
rect 11146 443898 11382 444134
rect 10826 408218 11062 408454
rect 11146 408218 11382 408454
rect 10826 407898 11062 408134
rect 11146 407898 11382 408134
rect 10826 372218 11062 372454
rect 11146 372218 11382 372454
rect 10826 371898 11062 372134
rect 11146 371898 11382 372134
rect 10826 336218 11062 336454
rect 11146 336218 11382 336454
rect 10826 335898 11062 336134
rect 11146 335898 11382 336134
rect 10826 300218 11062 300454
rect 11146 300218 11382 300454
rect 10826 299898 11062 300134
rect 11146 299898 11382 300134
rect 10826 264218 11062 264454
rect 11146 264218 11382 264454
rect 10826 263898 11062 264134
rect 11146 263898 11382 264134
rect 10826 228218 11062 228454
rect 11146 228218 11382 228454
rect 10826 227898 11062 228134
rect 11146 227898 11382 228134
rect 10826 192218 11062 192454
rect 11146 192218 11382 192454
rect 10826 191898 11062 192134
rect 11146 191898 11382 192134
rect 10826 156218 11062 156454
rect 11146 156218 11382 156454
rect 10826 155898 11062 156134
rect 11146 155898 11382 156134
rect 10826 120218 11062 120454
rect 11146 120218 11382 120454
rect 10826 119898 11062 120134
rect 11146 119898 11382 120134
rect 10826 84218 11062 84454
rect 11146 84218 11382 84454
rect 10826 83898 11062 84134
rect 11146 83898 11382 84134
rect 10826 48218 11062 48454
rect 11146 48218 11382 48454
rect 10826 47898 11062 48134
rect 11146 47898 11382 48134
rect 10826 12218 11062 12454
rect 11146 12218 11382 12454
rect 10826 11898 11062 12134
rect 11146 11898 11382 12134
rect 10826 -2502 11062 -2266
rect 11146 -2502 11382 -2266
rect 10826 -2822 11062 -2586
rect 11146 -2822 11382 -2586
rect 15326 707482 15562 707718
rect 15646 707482 15882 707718
rect 15326 707162 15562 707398
rect 15646 707162 15882 707398
rect 15326 700718 15562 700954
rect 15646 700718 15882 700954
rect 15326 700398 15562 700634
rect 15646 700398 15882 700634
rect 15326 664718 15562 664954
rect 15646 664718 15882 664954
rect 15326 664398 15562 664634
rect 15646 664398 15882 664634
rect 15326 628718 15562 628954
rect 15646 628718 15882 628954
rect 15326 628398 15562 628634
rect 15646 628398 15882 628634
rect 15326 592718 15562 592954
rect 15646 592718 15882 592954
rect 15326 592398 15562 592634
rect 15646 592398 15882 592634
rect 15326 556718 15562 556954
rect 15646 556718 15882 556954
rect 15326 556398 15562 556634
rect 15646 556398 15882 556634
rect 15326 520718 15562 520954
rect 15646 520718 15882 520954
rect 15326 520398 15562 520634
rect 15646 520398 15882 520634
rect 15326 484718 15562 484954
rect 15646 484718 15882 484954
rect 15326 484398 15562 484634
rect 15646 484398 15882 484634
rect 15326 448718 15562 448954
rect 15646 448718 15882 448954
rect 15326 448398 15562 448634
rect 15646 448398 15882 448634
rect 15326 412718 15562 412954
rect 15646 412718 15882 412954
rect 15326 412398 15562 412634
rect 15646 412398 15882 412634
rect 15326 376718 15562 376954
rect 15646 376718 15882 376954
rect 15326 376398 15562 376634
rect 15646 376398 15882 376634
rect 15326 340718 15562 340954
rect 15646 340718 15882 340954
rect 15326 340398 15562 340634
rect 15646 340398 15882 340634
rect 15326 304718 15562 304954
rect 15646 304718 15882 304954
rect 15326 304398 15562 304634
rect 15646 304398 15882 304634
rect 15326 268718 15562 268954
rect 15646 268718 15882 268954
rect 15326 268398 15562 268634
rect 15646 268398 15882 268634
rect 15326 232718 15562 232954
rect 15646 232718 15882 232954
rect 15326 232398 15562 232634
rect 15646 232398 15882 232634
rect 15326 196718 15562 196954
rect 15646 196718 15882 196954
rect 15326 196398 15562 196634
rect 15646 196398 15882 196634
rect 15326 160718 15562 160954
rect 15646 160718 15882 160954
rect 15326 160398 15562 160634
rect 15646 160398 15882 160634
rect 15326 124718 15562 124954
rect 15646 124718 15882 124954
rect 15326 124398 15562 124634
rect 15646 124398 15882 124634
rect 15326 88718 15562 88954
rect 15646 88718 15882 88954
rect 15326 88398 15562 88634
rect 15646 88398 15882 88634
rect 15326 52718 15562 52954
rect 15646 52718 15882 52954
rect 15326 52398 15562 52634
rect 15646 52398 15882 52634
rect 15326 16718 15562 16954
rect 15646 16718 15882 16954
rect 15326 16398 15562 16634
rect 15646 16398 15882 16634
rect 15326 -3462 15562 -3226
rect 15646 -3462 15882 -3226
rect 15326 -3782 15562 -3546
rect 15646 -3782 15882 -3546
rect 19826 708442 20062 708678
rect 20146 708442 20382 708678
rect 19826 708122 20062 708358
rect 20146 708122 20382 708358
rect 19826 669218 20062 669454
rect 20146 669218 20382 669454
rect 19826 668898 20062 669134
rect 20146 668898 20382 669134
rect 19826 633218 20062 633454
rect 20146 633218 20382 633454
rect 19826 632898 20062 633134
rect 20146 632898 20382 633134
rect 19826 597218 20062 597454
rect 20146 597218 20382 597454
rect 19826 596898 20062 597134
rect 20146 596898 20382 597134
rect 19826 561218 20062 561454
rect 20146 561218 20382 561454
rect 19826 560898 20062 561134
rect 20146 560898 20382 561134
rect 19826 525218 20062 525454
rect 20146 525218 20382 525454
rect 19826 524898 20062 525134
rect 20146 524898 20382 525134
rect 19826 489218 20062 489454
rect 20146 489218 20382 489454
rect 19826 488898 20062 489134
rect 20146 488898 20382 489134
rect 19826 453218 20062 453454
rect 20146 453218 20382 453454
rect 19826 452898 20062 453134
rect 20146 452898 20382 453134
rect 19826 417218 20062 417454
rect 20146 417218 20382 417454
rect 19826 416898 20062 417134
rect 20146 416898 20382 417134
rect 19826 381218 20062 381454
rect 20146 381218 20382 381454
rect 19826 380898 20062 381134
rect 20146 380898 20382 381134
rect 19826 345218 20062 345454
rect 20146 345218 20382 345454
rect 19826 344898 20062 345134
rect 20146 344898 20382 345134
rect 19826 309218 20062 309454
rect 20146 309218 20382 309454
rect 19826 308898 20062 309134
rect 20146 308898 20382 309134
rect 19826 273218 20062 273454
rect 20146 273218 20382 273454
rect 19826 272898 20062 273134
rect 20146 272898 20382 273134
rect 19826 237218 20062 237454
rect 20146 237218 20382 237454
rect 19826 236898 20062 237134
rect 20146 236898 20382 237134
rect 19826 201218 20062 201454
rect 20146 201218 20382 201454
rect 19826 200898 20062 201134
rect 20146 200898 20382 201134
rect 19826 165218 20062 165454
rect 20146 165218 20382 165454
rect 19826 164898 20062 165134
rect 20146 164898 20382 165134
rect 19826 129218 20062 129454
rect 20146 129218 20382 129454
rect 19826 128898 20062 129134
rect 20146 128898 20382 129134
rect 19826 93218 20062 93454
rect 20146 93218 20382 93454
rect 19826 92898 20062 93134
rect 20146 92898 20382 93134
rect 19826 57218 20062 57454
rect 20146 57218 20382 57454
rect 19826 56898 20062 57134
rect 20146 56898 20382 57134
rect 19826 21218 20062 21454
rect 20146 21218 20382 21454
rect 19826 20898 20062 21134
rect 20146 20898 20382 21134
rect 19826 -4422 20062 -4186
rect 20146 -4422 20382 -4186
rect 19826 -4742 20062 -4506
rect 20146 -4742 20382 -4506
rect 24326 709402 24562 709638
rect 24646 709402 24882 709638
rect 24326 709082 24562 709318
rect 24646 709082 24882 709318
rect 24326 673718 24562 673954
rect 24646 673718 24882 673954
rect 24326 673398 24562 673634
rect 24646 673398 24882 673634
rect 24326 637718 24562 637954
rect 24646 637718 24882 637954
rect 24326 637398 24562 637634
rect 24646 637398 24882 637634
rect 24326 601718 24562 601954
rect 24646 601718 24882 601954
rect 24326 601398 24562 601634
rect 24646 601398 24882 601634
rect 24326 565718 24562 565954
rect 24646 565718 24882 565954
rect 24326 565398 24562 565634
rect 24646 565398 24882 565634
rect 24326 529718 24562 529954
rect 24646 529718 24882 529954
rect 24326 529398 24562 529634
rect 24646 529398 24882 529634
rect 24326 493718 24562 493954
rect 24646 493718 24882 493954
rect 24326 493398 24562 493634
rect 24646 493398 24882 493634
rect 24326 457718 24562 457954
rect 24646 457718 24882 457954
rect 24326 457398 24562 457634
rect 24646 457398 24882 457634
rect 24326 421718 24562 421954
rect 24646 421718 24882 421954
rect 24326 421398 24562 421634
rect 24646 421398 24882 421634
rect 24326 385718 24562 385954
rect 24646 385718 24882 385954
rect 24326 385398 24562 385634
rect 24646 385398 24882 385634
rect 24326 349718 24562 349954
rect 24646 349718 24882 349954
rect 24326 349398 24562 349634
rect 24646 349398 24882 349634
rect 24326 313718 24562 313954
rect 24646 313718 24882 313954
rect 24326 313398 24562 313634
rect 24646 313398 24882 313634
rect 24326 277718 24562 277954
rect 24646 277718 24882 277954
rect 24326 277398 24562 277634
rect 24646 277398 24882 277634
rect 24326 241718 24562 241954
rect 24646 241718 24882 241954
rect 24326 241398 24562 241634
rect 24646 241398 24882 241634
rect 24326 205718 24562 205954
rect 24646 205718 24882 205954
rect 24326 205398 24562 205634
rect 24646 205398 24882 205634
rect 24326 169718 24562 169954
rect 24646 169718 24882 169954
rect 24326 169398 24562 169634
rect 24646 169398 24882 169634
rect 24326 133718 24562 133954
rect 24646 133718 24882 133954
rect 24326 133398 24562 133634
rect 24646 133398 24882 133634
rect 24326 97718 24562 97954
rect 24646 97718 24882 97954
rect 24326 97398 24562 97634
rect 24646 97398 24882 97634
rect 24326 61718 24562 61954
rect 24646 61718 24882 61954
rect 24326 61398 24562 61634
rect 24646 61398 24882 61634
rect 24326 25718 24562 25954
rect 24646 25718 24882 25954
rect 24326 25398 24562 25634
rect 24646 25398 24882 25634
rect 24326 -5382 24562 -5146
rect 24646 -5382 24882 -5146
rect 24326 -5702 24562 -5466
rect 24646 -5702 24882 -5466
rect 28826 710362 29062 710598
rect 29146 710362 29382 710598
rect 28826 710042 29062 710278
rect 29146 710042 29382 710278
rect 28826 678218 29062 678454
rect 29146 678218 29382 678454
rect 28826 677898 29062 678134
rect 29146 677898 29382 678134
rect 28826 642218 29062 642454
rect 29146 642218 29382 642454
rect 28826 641898 29062 642134
rect 29146 641898 29382 642134
rect 28826 606218 29062 606454
rect 29146 606218 29382 606454
rect 28826 605898 29062 606134
rect 29146 605898 29382 606134
rect 28826 570218 29062 570454
rect 29146 570218 29382 570454
rect 28826 569898 29062 570134
rect 29146 569898 29382 570134
rect 28826 534218 29062 534454
rect 29146 534218 29382 534454
rect 28826 533898 29062 534134
rect 29146 533898 29382 534134
rect 28826 498218 29062 498454
rect 29146 498218 29382 498454
rect 28826 497898 29062 498134
rect 29146 497898 29382 498134
rect 28826 462218 29062 462454
rect 29146 462218 29382 462454
rect 28826 461898 29062 462134
rect 29146 461898 29382 462134
rect 28826 426218 29062 426454
rect 29146 426218 29382 426454
rect 28826 425898 29062 426134
rect 29146 425898 29382 426134
rect 28826 390218 29062 390454
rect 29146 390218 29382 390454
rect 28826 389898 29062 390134
rect 29146 389898 29382 390134
rect 28826 354218 29062 354454
rect 29146 354218 29382 354454
rect 28826 353898 29062 354134
rect 29146 353898 29382 354134
rect 28826 318218 29062 318454
rect 29146 318218 29382 318454
rect 28826 317898 29062 318134
rect 29146 317898 29382 318134
rect 28826 282218 29062 282454
rect 29146 282218 29382 282454
rect 28826 281898 29062 282134
rect 29146 281898 29382 282134
rect 28826 246218 29062 246454
rect 29146 246218 29382 246454
rect 28826 245898 29062 246134
rect 29146 245898 29382 246134
rect 28826 210218 29062 210454
rect 29146 210218 29382 210454
rect 28826 209898 29062 210134
rect 29146 209898 29382 210134
rect 28826 174218 29062 174454
rect 29146 174218 29382 174454
rect 28826 173898 29062 174134
rect 29146 173898 29382 174134
rect 28826 138218 29062 138454
rect 29146 138218 29382 138454
rect 28826 137898 29062 138134
rect 29146 137898 29382 138134
rect 28826 102218 29062 102454
rect 29146 102218 29382 102454
rect 28826 101898 29062 102134
rect 29146 101898 29382 102134
rect 28826 66218 29062 66454
rect 29146 66218 29382 66454
rect 28826 65898 29062 66134
rect 29146 65898 29382 66134
rect 28826 30218 29062 30454
rect 29146 30218 29382 30454
rect 28826 29898 29062 30134
rect 29146 29898 29382 30134
rect 28826 -6342 29062 -6106
rect 29146 -6342 29382 -6106
rect 28826 -6662 29062 -6426
rect 29146 -6662 29382 -6426
rect 33326 711322 33562 711558
rect 33646 711322 33882 711558
rect 33326 711002 33562 711238
rect 33646 711002 33882 711238
rect 33326 682718 33562 682954
rect 33646 682718 33882 682954
rect 33326 682398 33562 682634
rect 33646 682398 33882 682634
rect 33326 646718 33562 646954
rect 33646 646718 33882 646954
rect 33326 646398 33562 646634
rect 33646 646398 33882 646634
rect 33326 610718 33562 610954
rect 33646 610718 33882 610954
rect 33326 610398 33562 610634
rect 33646 610398 33882 610634
rect 33326 574718 33562 574954
rect 33646 574718 33882 574954
rect 33326 574398 33562 574634
rect 33646 574398 33882 574634
rect 33326 538718 33562 538954
rect 33646 538718 33882 538954
rect 33326 538398 33562 538634
rect 33646 538398 33882 538634
rect 33326 502718 33562 502954
rect 33646 502718 33882 502954
rect 33326 502398 33562 502634
rect 33646 502398 33882 502634
rect 33326 466718 33562 466954
rect 33646 466718 33882 466954
rect 33326 466398 33562 466634
rect 33646 466398 33882 466634
rect 33326 430718 33562 430954
rect 33646 430718 33882 430954
rect 33326 430398 33562 430634
rect 33646 430398 33882 430634
rect 33326 394718 33562 394954
rect 33646 394718 33882 394954
rect 33326 394398 33562 394634
rect 33646 394398 33882 394634
rect 33326 358718 33562 358954
rect 33646 358718 33882 358954
rect 33326 358398 33562 358634
rect 33646 358398 33882 358634
rect 33326 322718 33562 322954
rect 33646 322718 33882 322954
rect 33326 322398 33562 322634
rect 33646 322398 33882 322634
rect 33326 286718 33562 286954
rect 33646 286718 33882 286954
rect 33326 286398 33562 286634
rect 33646 286398 33882 286634
rect 33326 250718 33562 250954
rect 33646 250718 33882 250954
rect 33326 250398 33562 250634
rect 33646 250398 33882 250634
rect 33326 214718 33562 214954
rect 33646 214718 33882 214954
rect 33326 214398 33562 214634
rect 33646 214398 33882 214634
rect 33326 178718 33562 178954
rect 33646 178718 33882 178954
rect 33326 178398 33562 178634
rect 33646 178398 33882 178634
rect 33326 142718 33562 142954
rect 33646 142718 33882 142954
rect 33326 142398 33562 142634
rect 33646 142398 33882 142634
rect 33326 106718 33562 106954
rect 33646 106718 33882 106954
rect 33326 106398 33562 106634
rect 33646 106398 33882 106634
rect 33326 70718 33562 70954
rect 33646 70718 33882 70954
rect 33326 70398 33562 70634
rect 33646 70398 33882 70634
rect 33326 34718 33562 34954
rect 33646 34718 33882 34954
rect 33326 34398 33562 34634
rect 33646 34398 33882 34634
rect 33326 -7302 33562 -7066
rect 33646 -7302 33882 -7066
rect 33326 -7622 33562 -7386
rect 33646 -7622 33882 -7386
rect 37826 704602 38062 704838
rect 38146 704602 38382 704838
rect 37826 704282 38062 704518
rect 38146 704282 38382 704518
rect 37826 687218 38062 687454
rect 38146 687218 38382 687454
rect 37826 686898 38062 687134
rect 38146 686898 38382 687134
rect 37826 651218 38062 651454
rect 38146 651218 38382 651454
rect 37826 650898 38062 651134
rect 38146 650898 38382 651134
rect 37826 615218 38062 615454
rect 38146 615218 38382 615454
rect 37826 614898 38062 615134
rect 38146 614898 38382 615134
rect 37826 579218 38062 579454
rect 38146 579218 38382 579454
rect 37826 578898 38062 579134
rect 38146 578898 38382 579134
rect 37826 543218 38062 543454
rect 38146 543218 38382 543454
rect 37826 542898 38062 543134
rect 38146 542898 38382 543134
rect 37826 507218 38062 507454
rect 38146 507218 38382 507454
rect 37826 506898 38062 507134
rect 38146 506898 38382 507134
rect 37826 471218 38062 471454
rect 38146 471218 38382 471454
rect 37826 470898 38062 471134
rect 38146 470898 38382 471134
rect 37826 435218 38062 435454
rect 38146 435218 38382 435454
rect 37826 434898 38062 435134
rect 38146 434898 38382 435134
rect 37826 399218 38062 399454
rect 38146 399218 38382 399454
rect 37826 398898 38062 399134
rect 38146 398898 38382 399134
rect 37826 363218 38062 363454
rect 38146 363218 38382 363454
rect 37826 362898 38062 363134
rect 38146 362898 38382 363134
rect 37826 327218 38062 327454
rect 38146 327218 38382 327454
rect 37826 326898 38062 327134
rect 38146 326898 38382 327134
rect 37826 291218 38062 291454
rect 38146 291218 38382 291454
rect 37826 290898 38062 291134
rect 38146 290898 38382 291134
rect 37826 255218 38062 255454
rect 38146 255218 38382 255454
rect 37826 254898 38062 255134
rect 38146 254898 38382 255134
rect 37826 219218 38062 219454
rect 38146 219218 38382 219454
rect 37826 218898 38062 219134
rect 38146 218898 38382 219134
rect 37826 183218 38062 183454
rect 38146 183218 38382 183454
rect 37826 182898 38062 183134
rect 38146 182898 38382 183134
rect 37826 147218 38062 147454
rect 38146 147218 38382 147454
rect 37826 146898 38062 147134
rect 38146 146898 38382 147134
rect 37826 111218 38062 111454
rect 38146 111218 38382 111454
rect 37826 110898 38062 111134
rect 38146 110898 38382 111134
rect 37826 75218 38062 75454
rect 38146 75218 38382 75454
rect 37826 74898 38062 75134
rect 38146 74898 38382 75134
rect 37826 39218 38062 39454
rect 38146 39218 38382 39454
rect 37826 38898 38062 39134
rect 38146 38898 38382 39134
rect 37826 3218 38062 3454
rect 38146 3218 38382 3454
rect 37826 2898 38062 3134
rect 38146 2898 38382 3134
rect 37826 -582 38062 -346
rect 38146 -582 38382 -346
rect 37826 -902 38062 -666
rect 38146 -902 38382 -666
rect 42326 705562 42562 705798
rect 42646 705562 42882 705798
rect 42326 705242 42562 705478
rect 42646 705242 42882 705478
rect 42326 691718 42562 691954
rect 42646 691718 42882 691954
rect 42326 691398 42562 691634
rect 42646 691398 42882 691634
rect 42326 655718 42562 655954
rect 42646 655718 42882 655954
rect 42326 655398 42562 655634
rect 42646 655398 42882 655634
rect 42326 619718 42562 619954
rect 42646 619718 42882 619954
rect 42326 619398 42562 619634
rect 42646 619398 42882 619634
rect 42326 583718 42562 583954
rect 42646 583718 42882 583954
rect 42326 583398 42562 583634
rect 42646 583398 42882 583634
rect 42326 547718 42562 547954
rect 42646 547718 42882 547954
rect 42326 547398 42562 547634
rect 42646 547398 42882 547634
rect 42326 511718 42562 511954
rect 42646 511718 42882 511954
rect 42326 511398 42562 511634
rect 42646 511398 42882 511634
rect 42326 475718 42562 475954
rect 42646 475718 42882 475954
rect 42326 475398 42562 475634
rect 42646 475398 42882 475634
rect 42326 439718 42562 439954
rect 42646 439718 42882 439954
rect 42326 439398 42562 439634
rect 42646 439398 42882 439634
rect 42326 403718 42562 403954
rect 42646 403718 42882 403954
rect 42326 403398 42562 403634
rect 42646 403398 42882 403634
rect 42326 367718 42562 367954
rect 42646 367718 42882 367954
rect 42326 367398 42562 367634
rect 42646 367398 42882 367634
rect 42326 331718 42562 331954
rect 42646 331718 42882 331954
rect 42326 331398 42562 331634
rect 42646 331398 42882 331634
rect 42326 295718 42562 295954
rect 42646 295718 42882 295954
rect 42326 295398 42562 295634
rect 42646 295398 42882 295634
rect 42326 259718 42562 259954
rect 42646 259718 42882 259954
rect 42326 259398 42562 259634
rect 42646 259398 42882 259634
rect 42326 223718 42562 223954
rect 42646 223718 42882 223954
rect 42326 223398 42562 223634
rect 42646 223398 42882 223634
rect 42326 187718 42562 187954
rect 42646 187718 42882 187954
rect 42326 187398 42562 187634
rect 42646 187398 42882 187634
rect 42326 151718 42562 151954
rect 42646 151718 42882 151954
rect 42326 151398 42562 151634
rect 42646 151398 42882 151634
rect 42326 115718 42562 115954
rect 42646 115718 42882 115954
rect 42326 115398 42562 115634
rect 42646 115398 42882 115634
rect 42326 79718 42562 79954
rect 42646 79718 42882 79954
rect 42326 79398 42562 79634
rect 42646 79398 42882 79634
rect 42326 43718 42562 43954
rect 42646 43718 42882 43954
rect 42326 43398 42562 43634
rect 42646 43398 42882 43634
rect 42326 7718 42562 7954
rect 42646 7718 42882 7954
rect 42326 7398 42562 7634
rect 42646 7398 42882 7634
rect 42326 -1542 42562 -1306
rect 42646 -1542 42882 -1306
rect 42326 -1862 42562 -1626
rect 42646 -1862 42882 -1626
rect 46826 706522 47062 706758
rect 47146 706522 47382 706758
rect 46826 706202 47062 706438
rect 47146 706202 47382 706438
rect 46826 696218 47062 696454
rect 47146 696218 47382 696454
rect 46826 695898 47062 696134
rect 47146 695898 47382 696134
rect 46826 660218 47062 660454
rect 47146 660218 47382 660454
rect 46826 659898 47062 660134
rect 47146 659898 47382 660134
rect 46826 624218 47062 624454
rect 47146 624218 47382 624454
rect 46826 623898 47062 624134
rect 47146 623898 47382 624134
rect 46826 588218 47062 588454
rect 47146 588218 47382 588454
rect 46826 587898 47062 588134
rect 47146 587898 47382 588134
rect 46826 552218 47062 552454
rect 47146 552218 47382 552454
rect 46826 551898 47062 552134
rect 47146 551898 47382 552134
rect 46826 516218 47062 516454
rect 47146 516218 47382 516454
rect 46826 515898 47062 516134
rect 47146 515898 47382 516134
rect 46826 480218 47062 480454
rect 47146 480218 47382 480454
rect 46826 479898 47062 480134
rect 47146 479898 47382 480134
rect 46826 444218 47062 444454
rect 47146 444218 47382 444454
rect 46826 443898 47062 444134
rect 47146 443898 47382 444134
rect 46826 408218 47062 408454
rect 47146 408218 47382 408454
rect 46826 407898 47062 408134
rect 47146 407898 47382 408134
rect 46826 372218 47062 372454
rect 47146 372218 47382 372454
rect 46826 371898 47062 372134
rect 47146 371898 47382 372134
rect 46826 336218 47062 336454
rect 47146 336218 47382 336454
rect 46826 335898 47062 336134
rect 47146 335898 47382 336134
rect 46826 300218 47062 300454
rect 47146 300218 47382 300454
rect 46826 299898 47062 300134
rect 47146 299898 47382 300134
rect 46826 264218 47062 264454
rect 47146 264218 47382 264454
rect 46826 263898 47062 264134
rect 47146 263898 47382 264134
rect 46826 228218 47062 228454
rect 47146 228218 47382 228454
rect 46826 227898 47062 228134
rect 47146 227898 47382 228134
rect 46826 192218 47062 192454
rect 47146 192218 47382 192454
rect 46826 191898 47062 192134
rect 47146 191898 47382 192134
rect 46826 156218 47062 156454
rect 47146 156218 47382 156454
rect 46826 155898 47062 156134
rect 47146 155898 47382 156134
rect 46826 120218 47062 120454
rect 47146 120218 47382 120454
rect 46826 119898 47062 120134
rect 47146 119898 47382 120134
rect 46826 84218 47062 84454
rect 47146 84218 47382 84454
rect 46826 83898 47062 84134
rect 47146 83898 47382 84134
rect 46826 48218 47062 48454
rect 47146 48218 47382 48454
rect 46826 47898 47062 48134
rect 47146 47898 47382 48134
rect 46826 12218 47062 12454
rect 47146 12218 47382 12454
rect 46826 11898 47062 12134
rect 47146 11898 47382 12134
rect 46826 -2502 47062 -2266
rect 47146 -2502 47382 -2266
rect 46826 -2822 47062 -2586
rect 47146 -2822 47382 -2586
rect 51326 707482 51562 707718
rect 51646 707482 51882 707718
rect 51326 707162 51562 707398
rect 51646 707162 51882 707398
rect 51326 700718 51562 700954
rect 51646 700718 51882 700954
rect 51326 700398 51562 700634
rect 51646 700398 51882 700634
rect 51326 664718 51562 664954
rect 51646 664718 51882 664954
rect 51326 664398 51562 664634
rect 51646 664398 51882 664634
rect 51326 628718 51562 628954
rect 51646 628718 51882 628954
rect 51326 628398 51562 628634
rect 51646 628398 51882 628634
rect 51326 592718 51562 592954
rect 51646 592718 51882 592954
rect 51326 592398 51562 592634
rect 51646 592398 51882 592634
rect 51326 556718 51562 556954
rect 51646 556718 51882 556954
rect 51326 556398 51562 556634
rect 51646 556398 51882 556634
rect 51326 520718 51562 520954
rect 51646 520718 51882 520954
rect 51326 520398 51562 520634
rect 51646 520398 51882 520634
rect 51326 484718 51562 484954
rect 51646 484718 51882 484954
rect 51326 484398 51562 484634
rect 51646 484398 51882 484634
rect 51326 448718 51562 448954
rect 51646 448718 51882 448954
rect 51326 448398 51562 448634
rect 51646 448398 51882 448634
rect 51326 412718 51562 412954
rect 51646 412718 51882 412954
rect 51326 412398 51562 412634
rect 51646 412398 51882 412634
rect 51326 376718 51562 376954
rect 51646 376718 51882 376954
rect 51326 376398 51562 376634
rect 51646 376398 51882 376634
rect 51326 340718 51562 340954
rect 51646 340718 51882 340954
rect 51326 340398 51562 340634
rect 51646 340398 51882 340634
rect 51326 304718 51562 304954
rect 51646 304718 51882 304954
rect 51326 304398 51562 304634
rect 51646 304398 51882 304634
rect 51326 268718 51562 268954
rect 51646 268718 51882 268954
rect 51326 268398 51562 268634
rect 51646 268398 51882 268634
rect 51326 232718 51562 232954
rect 51646 232718 51882 232954
rect 51326 232398 51562 232634
rect 51646 232398 51882 232634
rect 51326 196718 51562 196954
rect 51646 196718 51882 196954
rect 51326 196398 51562 196634
rect 51646 196398 51882 196634
rect 51326 160718 51562 160954
rect 51646 160718 51882 160954
rect 51326 160398 51562 160634
rect 51646 160398 51882 160634
rect 51326 124718 51562 124954
rect 51646 124718 51882 124954
rect 51326 124398 51562 124634
rect 51646 124398 51882 124634
rect 51326 88718 51562 88954
rect 51646 88718 51882 88954
rect 51326 88398 51562 88634
rect 51646 88398 51882 88634
rect 51326 52718 51562 52954
rect 51646 52718 51882 52954
rect 51326 52398 51562 52634
rect 51646 52398 51882 52634
rect 51326 16718 51562 16954
rect 51646 16718 51882 16954
rect 51326 16398 51562 16634
rect 51646 16398 51882 16634
rect 51326 -3462 51562 -3226
rect 51646 -3462 51882 -3226
rect 51326 -3782 51562 -3546
rect 51646 -3782 51882 -3546
rect 55826 708442 56062 708678
rect 56146 708442 56382 708678
rect 55826 708122 56062 708358
rect 56146 708122 56382 708358
rect 55826 669218 56062 669454
rect 56146 669218 56382 669454
rect 55826 668898 56062 669134
rect 56146 668898 56382 669134
rect 55826 633218 56062 633454
rect 56146 633218 56382 633454
rect 55826 632898 56062 633134
rect 56146 632898 56382 633134
rect 55826 597218 56062 597454
rect 56146 597218 56382 597454
rect 55826 596898 56062 597134
rect 56146 596898 56382 597134
rect 55826 561218 56062 561454
rect 56146 561218 56382 561454
rect 55826 560898 56062 561134
rect 56146 560898 56382 561134
rect 55826 525218 56062 525454
rect 56146 525218 56382 525454
rect 55826 524898 56062 525134
rect 56146 524898 56382 525134
rect 55826 489218 56062 489454
rect 56146 489218 56382 489454
rect 55826 488898 56062 489134
rect 56146 488898 56382 489134
rect 55826 453218 56062 453454
rect 56146 453218 56382 453454
rect 55826 452898 56062 453134
rect 56146 452898 56382 453134
rect 55826 417218 56062 417454
rect 56146 417218 56382 417454
rect 55826 416898 56062 417134
rect 56146 416898 56382 417134
rect 55826 381218 56062 381454
rect 56146 381218 56382 381454
rect 55826 380898 56062 381134
rect 56146 380898 56382 381134
rect 55826 345218 56062 345454
rect 56146 345218 56382 345454
rect 55826 344898 56062 345134
rect 56146 344898 56382 345134
rect 55826 309218 56062 309454
rect 56146 309218 56382 309454
rect 55826 308898 56062 309134
rect 56146 308898 56382 309134
rect 55826 273218 56062 273454
rect 56146 273218 56382 273454
rect 55826 272898 56062 273134
rect 56146 272898 56382 273134
rect 55826 237218 56062 237454
rect 56146 237218 56382 237454
rect 55826 236898 56062 237134
rect 56146 236898 56382 237134
rect 55826 201218 56062 201454
rect 56146 201218 56382 201454
rect 55826 200898 56062 201134
rect 56146 200898 56382 201134
rect 55826 165218 56062 165454
rect 56146 165218 56382 165454
rect 55826 164898 56062 165134
rect 56146 164898 56382 165134
rect 55826 129218 56062 129454
rect 56146 129218 56382 129454
rect 55826 128898 56062 129134
rect 56146 128898 56382 129134
rect 55826 93218 56062 93454
rect 56146 93218 56382 93454
rect 55826 92898 56062 93134
rect 56146 92898 56382 93134
rect 55826 57218 56062 57454
rect 56146 57218 56382 57454
rect 55826 56898 56062 57134
rect 56146 56898 56382 57134
rect 55826 21218 56062 21454
rect 56146 21218 56382 21454
rect 55826 20898 56062 21134
rect 56146 20898 56382 21134
rect 55826 -4422 56062 -4186
rect 56146 -4422 56382 -4186
rect 55826 -4742 56062 -4506
rect 56146 -4742 56382 -4506
rect 60326 709402 60562 709638
rect 60646 709402 60882 709638
rect 60326 709082 60562 709318
rect 60646 709082 60882 709318
rect 60326 673718 60562 673954
rect 60646 673718 60882 673954
rect 60326 673398 60562 673634
rect 60646 673398 60882 673634
rect 60326 637718 60562 637954
rect 60646 637718 60882 637954
rect 60326 637398 60562 637634
rect 60646 637398 60882 637634
rect 60326 601718 60562 601954
rect 60646 601718 60882 601954
rect 60326 601398 60562 601634
rect 60646 601398 60882 601634
rect 60326 565718 60562 565954
rect 60646 565718 60882 565954
rect 60326 565398 60562 565634
rect 60646 565398 60882 565634
rect 60326 529718 60562 529954
rect 60646 529718 60882 529954
rect 60326 529398 60562 529634
rect 60646 529398 60882 529634
rect 60326 493718 60562 493954
rect 60646 493718 60882 493954
rect 60326 493398 60562 493634
rect 60646 493398 60882 493634
rect 60326 457718 60562 457954
rect 60646 457718 60882 457954
rect 60326 457398 60562 457634
rect 60646 457398 60882 457634
rect 60326 421718 60562 421954
rect 60646 421718 60882 421954
rect 60326 421398 60562 421634
rect 60646 421398 60882 421634
rect 60326 385718 60562 385954
rect 60646 385718 60882 385954
rect 60326 385398 60562 385634
rect 60646 385398 60882 385634
rect 60326 349718 60562 349954
rect 60646 349718 60882 349954
rect 60326 349398 60562 349634
rect 60646 349398 60882 349634
rect 60326 313718 60562 313954
rect 60646 313718 60882 313954
rect 60326 313398 60562 313634
rect 60646 313398 60882 313634
rect 60326 277718 60562 277954
rect 60646 277718 60882 277954
rect 60326 277398 60562 277634
rect 60646 277398 60882 277634
rect 60326 241718 60562 241954
rect 60646 241718 60882 241954
rect 60326 241398 60562 241634
rect 60646 241398 60882 241634
rect 60326 205718 60562 205954
rect 60646 205718 60882 205954
rect 60326 205398 60562 205634
rect 60646 205398 60882 205634
rect 60326 169718 60562 169954
rect 60646 169718 60882 169954
rect 60326 169398 60562 169634
rect 60646 169398 60882 169634
rect 60326 133718 60562 133954
rect 60646 133718 60882 133954
rect 60326 133398 60562 133634
rect 60646 133398 60882 133634
rect 60326 97718 60562 97954
rect 60646 97718 60882 97954
rect 60326 97398 60562 97634
rect 60646 97398 60882 97634
rect 60326 61718 60562 61954
rect 60646 61718 60882 61954
rect 60326 61398 60562 61634
rect 60646 61398 60882 61634
rect 60326 25718 60562 25954
rect 60646 25718 60882 25954
rect 60326 25398 60562 25634
rect 60646 25398 60882 25634
rect 60326 -5382 60562 -5146
rect 60646 -5382 60882 -5146
rect 60326 -5702 60562 -5466
rect 60646 -5702 60882 -5466
rect 64826 710362 65062 710598
rect 65146 710362 65382 710598
rect 64826 710042 65062 710278
rect 65146 710042 65382 710278
rect 64826 678218 65062 678454
rect 65146 678218 65382 678454
rect 64826 677898 65062 678134
rect 65146 677898 65382 678134
rect 64826 642218 65062 642454
rect 65146 642218 65382 642454
rect 64826 641898 65062 642134
rect 65146 641898 65382 642134
rect 64826 606218 65062 606454
rect 65146 606218 65382 606454
rect 64826 605898 65062 606134
rect 65146 605898 65382 606134
rect 64826 570218 65062 570454
rect 65146 570218 65382 570454
rect 64826 569898 65062 570134
rect 65146 569898 65382 570134
rect 64826 534218 65062 534454
rect 65146 534218 65382 534454
rect 64826 533898 65062 534134
rect 65146 533898 65382 534134
rect 64826 498218 65062 498454
rect 65146 498218 65382 498454
rect 64826 497898 65062 498134
rect 65146 497898 65382 498134
rect 64826 462218 65062 462454
rect 65146 462218 65382 462454
rect 64826 461898 65062 462134
rect 65146 461898 65382 462134
rect 64826 426218 65062 426454
rect 65146 426218 65382 426454
rect 64826 425898 65062 426134
rect 65146 425898 65382 426134
rect 64826 390218 65062 390454
rect 65146 390218 65382 390454
rect 64826 389898 65062 390134
rect 65146 389898 65382 390134
rect 64826 354218 65062 354454
rect 65146 354218 65382 354454
rect 64826 353898 65062 354134
rect 65146 353898 65382 354134
rect 64826 318218 65062 318454
rect 65146 318218 65382 318454
rect 64826 317898 65062 318134
rect 65146 317898 65382 318134
rect 64826 282218 65062 282454
rect 65146 282218 65382 282454
rect 64826 281898 65062 282134
rect 65146 281898 65382 282134
rect 64826 246218 65062 246454
rect 65146 246218 65382 246454
rect 64826 245898 65062 246134
rect 65146 245898 65382 246134
rect 64826 210218 65062 210454
rect 65146 210218 65382 210454
rect 64826 209898 65062 210134
rect 65146 209898 65382 210134
rect 64826 174218 65062 174454
rect 65146 174218 65382 174454
rect 64826 173898 65062 174134
rect 65146 173898 65382 174134
rect 64826 138218 65062 138454
rect 65146 138218 65382 138454
rect 64826 137898 65062 138134
rect 65146 137898 65382 138134
rect 64826 102218 65062 102454
rect 65146 102218 65382 102454
rect 64826 101898 65062 102134
rect 65146 101898 65382 102134
rect 64826 66218 65062 66454
rect 65146 66218 65382 66454
rect 64826 65898 65062 66134
rect 65146 65898 65382 66134
rect 64826 30218 65062 30454
rect 65146 30218 65382 30454
rect 64826 29898 65062 30134
rect 65146 29898 65382 30134
rect 64826 -6342 65062 -6106
rect 65146 -6342 65382 -6106
rect 64826 -6662 65062 -6426
rect 65146 -6662 65382 -6426
rect 69326 711322 69562 711558
rect 69646 711322 69882 711558
rect 69326 711002 69562 711238
rect 69646 711002 69882 711238
rect 69326 682718 69562 682954
rect 69646 682718 69882 682954
rect 69326 682398 69562 682634
rect 69646 682398 69882 682634
rect 69326 646718 69562 646954
rect 69646 646718 69882 646954
rect 69326 646398 69562 646634
rect 69646 646398 69882 646634
rect 69326 610718 69562 610954
rect 69646 610718 69882 610954
rect 69326 610398 69562 610634
rect 69646 610398 69882 610634
rect 69326 574718 69562 574954
rect 69646 574718 69882 574954
rect 69326 574398 69562 574634
rect 69646 574398 69882 574634
rect 69326 538718 69562 538954
rect 69646 538718 69882 538954
rect 69326 538398 69562 538634
rect 69646 538398 69882 538634
rect 69326 502718 69562 502954
rect 69646 502718 69882 502954
rect 69326 502398 69562 502634
rect 69646 502398 69882 502634
rect 69326 466718 69562 466954
rect 69646 466718 69882 466954
rect 69326 466398 69562 466634
rect 69646 466398 69882 466634
rect 69326 430718 69562 430954
rect 69646 430718 69882 430954
rect 69326 430398 69562 430634
rect 69646 430398 69882 430634
rect 69326 394718 69562 394954
rect 69646 394718 69882 394954
rect 69326 394398 69562 394634
rect 69646 394398 69882 394634
rect 69326 358718 69562 358954
rect 69646 358718 69882 358954
rect 69326 358398 69562 358634
rect 69646 358398 69882 358634
rect 69326 322718 69562 322954
rect 69646 322718 69882 322954
rect 69326 322398 69562 322634
rect 69646 322398 69882 322634
rect 69326 286718 69562 286954
rect 69646 286718 69882 286954
rect 69326 286398 69562 286634
rect 69646 286398 69882 286634
rect 69326 250718 69562 250954
rect 69646 250718 69882 250954
rect 69326 250398 69562 250634
rect 69646 250398 69882 250634
rect 69326 214718 69562 214954
rect 69646 214718 69882 214954
rect 69326 214398 69562 214634
rect 69646 214398 69882 214634
rect 69326 178718 69562 178954
rect 69646 178718 69882 178954
rect 69326 178398 69562 178634
rect 69646 178398 69882 178634
rect 69326 142718 69562 142954
rect 69646 142718 69882 142954
rect 69326 142398 69562 142634
rect 69646 142398 69882 142634
rect 69326 106718 69562 106954
rect 69646 106718 69882 106954
rect 69326 106398 69562 106634
rect 69646 106398 69882 106634
rect 69326 70718 69562 70954
rect 69646 70718 69882 70954
rect 69326 70398 69562 70634
rect 69646 70398 69882 70634
rect 69326 34718 69562 34954
rect 69646 34718 69882 34954
rect 69326 34398 69562 34634
rect 69646 34398 69882 34634
rect 69326 -7302 69562 -7066
rect 69646 -7302 69882 -7066
rect 69326 -7622 69562 -7386
rect 69646 -7622 69882 -7386
rect 73826 704602 74062 704838
rect 74146 704602 74382 704838
rect 73826 704282 74062 704518
rect 74146 704282 74382 704518
rect 73826 687218 74062 687454
rect 74146 687218 74382 687454
rect 73826 686898 74062 687134
rect 74146 686898 74382 687134
rect 73826 651218 74062 651454
rect 74146 651218 74382 651454
rect 73826 650898 74062 651134
rect 74146 650898 74382 651134
rect 73826 615218 74062 615454
rect 74146 615218 74382 615454
rect 73826 614898 74062 615134
rect 74146 614898 74382 615134
rect 73826 579218 74062 579454
rect 74146 579218 74382 579454
rect 73826 578898 74062 579134
rect 74146 578898 74382 579134
rect 73826 543218 74062 543454
rect 74146 543218 74382 543454
rect 73826 542898 74062 543134
rect 74146 542898 74382 543134
rect 73826 507218 74062 507454
rect 74146 507218 74382 507454
rect 73826 506898 74062 507134
rect 74146 506898 74382 507134
rect 73826 471218 74062 471454
rect 74146 471218 74382 471454
rect 73826 470898 74062 471134
rect 74146 470898 74382 471134
rect 73826 435218 74062 435454
rect 74146 435218 74382 435454
rect 73826 434898 74062 435134
rect 74146 434898 74382 435134
rect 73826 399218 74062 399454
rect 74146 399218 74382 399454
rect 73826 398898 74062 399134
rect 74146 398898 74382 399134
rect 73826 363218 74062 363454
rect 74146 363218 74382 363454
rect 73826 362898 74062 363134
rect 74146 362898 74382 363134
rect 73826 327218 74062 327454
rect 74146 327218 74382 327454
rect 73826 326898 74062 327134
rect 74146 326898 74382 327134
rect 73826 291218 74062 291454
rect 74146 291218 74382 291454
rect 73826 290898 74062 291134
rect 74146 290898 74382 291134
rect 73826 255218 74062 255454
rect 74146 255218 74382 255454
rect 73826 254898 74062 255134
rect 74146 254898 74382 255134
rect 73826 219218 74062 219454
rect 74146 219218 74382 219454
rect 73826 218898 74062 219134
rect 74146 218898 74382 219134
rect 73826 183218 74062 183454
rect 74146 183218 74382 183454
rect 73826 182898 74062 183134
rect 74146 182898 74382 183134
rect 73826 147218 74062 147454
rect 74146 147218 74382 147454
rect 73826 146898 74062 147134
rect 74146 146898 74382 147134
rect 73826 111218 74062 111454
rect 74146 111218 74382 111454
rect 73826 110898 74062 111134
rect 74146 110898 74382 111134
rect 73826 75218 74062 75454
rect 74146 75218 74382 75454
rect 73826 74898 74062 75134
rect 74146 74898 74382 75134
rect 73826 39218 74062 39454
rect 74146 39218 74382 39454
rect 73826 38898 74062 39134
rect 74146 38898 74382 39134
rect 73826 3218 74062 3454
rect 74146 3218 74382 3454
rect 73826 2898 74062 3134
rect 74146 2898 74382 3134
rect 73826 -582 74062 -346
rect 74146 -582 74382 -346
rect 73826 -902 74062 -666
rect 74146 -902 74382 -666
rect 78326 705562 78562 705798
rect 78646 705562 78882 705798
rect 78326 705242 78562 705478
rect 78646 705242 78882 705478
rect 78326 691718 78562 691954
rect 78646 691718 78882 691954
rect 78326 691398 78562 691634
rect 78646 691398 78882 691634
rect 78326 655718 78562 655954
rect 78646 655718 78882 655954
rect 78326 655398 78562 655634
rect 78646 655398 78882 655634
rect 78326 619718 78562 619954
rect 78646 619718 78882 619954
rect 78326 619398 78562 619634
rect 78646 619398 78882 619634
rect 78326 583718 78562 583954
rect 78646 583718 78882 583954
rect 78326 583398 78562 583634
rect 78646 583398 78882 583634
rect 78326 547718 78562 547954
rect 78646 547718 78882 547954
rect 78326 547398 78562 547634
rect 78646 547398 78882 547634
rect 78326 511718 78562 511954
rect 78646 511718 78882 511954
rect 78326 511398 78562 511634
rect 78646 511398 78882 511634
rect 78326 475718 78562 475954
rect 78646 475718 78882 475954
rect 78326 475398 78562 475634
rect 78646 475398 78882 475634
rect 78326 439718 78562 439954
rect 78646 439718 78882 439954
rect 78326 439398 78562 439634
rect 78646 439398 78882 439634
rect 78326 403718 78562 403954
rect 78646 403718 78882 403954
rect 78326 403398 78562 403634
rect 78646 403398 78882 403634
rect 78326 367718 78562 367954
rect 78646 367718 78882 367954
rect 78326 367398 78562 367634
rect 78646 367398 78882 367634
rect 78326 331718 78562 331954
rect 78646 331718 78882 331954
rect 78326 331398 78562 331634
rect 78646 331398 78882 331634
rect 78326 295718 78562 295954
rect 78646 295718 78882 295954
rect 78326 295398 78562 295634
rect 78646 295398 78882 295634
rect 78326 259718 78562 259954
rect 78646 259718 78882 259954
rect 78326 259398 78562 259634
rect 78646 259398 78882 259634
rect 78326 223718 78562 223954
rect 78646 223718 78882 223954
rect 78326 223398 78562 223634
rect 78646 223398 78882 223634
rect 78326 187718 78562 187954
rect 78646 187718 78882 187954
rect 78326 187398 78562 187634
rect 78646 187398 78882 187634
rect 78326 151718 78562 151954
rect 78646 151718 78882 151954
rect 78326 151398 78562 151634
rect 78646 151398 78882 151634
rect 78326 115718 78562 115954
rect 78646 115718 78882 115954
rect 78326 115398 78562 115634
rect 78646 115398 78882 115634
rect 78326 79718 78562 79954
rect 78646 79718 78882 79954
rect 78326 79398 78562 79634
rect 78646 79398 78882 79634
rect 78326 43718 78562 43954
rect 78646 43718 78882 43954
rect 78326 43398 78562 43634
rect 78646 43398 78882 43634
rect 78326 7718 78562 7954
rect 78646 7718 78882 7954
rect 78326 7398 78562 7634
rect 78646 7398 78882 7634
rect 78326 -1542 78562 -1306
rect 78646 -1542 78882 -1306
rect 78326 -1862 78562 -1626
rect 78646 -1862 78882 -1626
rect 82826 706522 83062 706758
rect 83146 706522 83382 706758
rect 82826 706202 83062 706438
rect 83146 706202 83382 706438
rect 82826 696218 83062 696454
rect 83146 696218 83382 696454
rect 82826 695898 83062 696134
rect 83146 695898 83382 696134
rect 82826 660218 83062 660454
rect 83146 660218 83382 660454
rect 82826 659898 83062 660134
rect 83146 659898 83382 660134
rect 82826 624218 83062 624454
rect 83146 624218 83382 624454
rect 82826 623898 83062 624134
rect 83146 623898 83382 624134
rect 82826 588218 83062 588454
rect 83146 588218 83382 588454
rect 82826 587898 83062 588134
rect 83146 587898 83382 588134
rect 82826 552218 83062 552454
rect 83146 552218 83382 552454
rect 82826 551898 83062 552134
rect 83146 551898 83382 552134
rect 82826 516218 83062 516454
rect 83146 516218 83382 516454
rect 82826 515898 83062 516134
rect 83146 515898 83382 516134
rect 82826 480218 83062 480454
rect 83146 480218 83382 480454
rect 82826 479898 83062 480134
rect 83146 479898 83382 480134
rect 82826 444218 83062 444454
rect 83146 444218 83382 444454
rect 82826 443898 83062 444134
rect 83146 443898 83382 444134
rect 82826 408218 83062 408454
rect 83146 408218 83382 408454
rect 82826 407898 83062 408134
rect 83146 407898 83382 408134
rect 82826 372218 83062 372454
rect 83146 372218 83382 372454
rect 82826 371898 83062 372134
rect 83146 371898 83382 372134
rect 82826 336218 83062 336454
rect 83146 336218 83382 336454
rect 82826 335898 83062 336134
rect 83146 335898 83382 336134
rect 82826 300218 83062 300454
rect 83146 300218 83382 300454
rect 82826 299898 83062 300134
rect 83146 299898 83382 300134
rect 82826 264218 83062 264454
rect 83146 264218 83382 264454
rect 82826 263898 83062 264134
rect 83146 263898 83382 264134
rect 82826 228218 83062 228454
rect 83146 228218 83382 228454
rect 82826 227898 83062 228134
rect 83146 227898 83382 228134
rect 82826 192218 83062 192454
rect 83146 192218 83382 192454
rect 82826 191898 83062 192134
rect 83146 191898 83382 192134
rect 82826 156218 83062 156454
rect 83146 156218 83382 156454
rect 82826 155898 83062 156134
rect 83146 155898 83382 156134
rect 82826 120218 83062 120454
rect 83146 120218 83382 120454
rect 82826 119898 83062 120134
rect 83146 119898 83382 120134
rect 82826 84218 83062 84454
rect 83146 84218 83382 84454
rect 82826 83898 83062 84134
rect 83146 83898 83382 84134
rect 82826 48218 83062 48454
rect 83146 48218 83382 48454
rect 82826 47898 83062 48134
rect 83146 47898 83382 48134
rect 82826 12218 83062 12454
rect 83146 12218 83382 12454
rect 82826 11898 83062 12134
rect 83146 11898 83382 12134
rect 82826 -2502 83062 -2266
rect 83146 -2502 83382 -2266
rect 82826 -2822 83062 -2586
rect 83146 -2822 83382 -2586
rect 87326 707482 87562 707718
rect 87646 707482 87882 707718
rect 87326 707162 87562 707398
rect 87646 707162 87882 707398
rect 87326 700718 87562 700954
rect 87646 700718 87882 700954
rect 87326 700398 87562 700634
rect 87646 700398 87882 700634
rect 87326 664718 87562 664954
rect 87646 664718 87882 664954
rect 87326 664398 87562 664634
rect 87646 664398 87882 664634
rect 87326 628718 87562 628954
rect 87646 628718 87882 628954
rect 87326 628398 87562 628634
rect 87646 628398 87882 628634
rect 87326 592718 87562 592954
rect 87646 592718 87882 592954
rect 87326 592398 87562 592634
rect 87646 592398 87882 592634
rect 87326 556718 87562 556954
rect 87646 556718 87882 556954
rect 87326 556398 87562 556634
rect 87646 556398 87882 556634
rect 87326 520718 87562 520954
rect 87646 520718 87882 520954
rect 87326 520398 87562 520634
rect 87646 520398 87882 520634
rect 87326 484718 87562 484954
rect 87646 484718 87882 484954
rect 87326 484398 87562 484634
rect 87646 484398 87882 484634
rect 87326 448718 87562 448954
rect 87646 448718 87882 448954
rect 87326 448398 87562 448634
rect 87646 448398 87882 448634
rect 87326 412718 87562 412954
rect 87646 412718 87882 412954
rect 87326 412398 87562 412634
rect 87646 412398 87882 412634
rect 87326 376718 87562 376954
rect 87646 376718 87882 376954
rect 87326 376398 87562 376634
rect 87646 376398 87882 376634
rect 87326 340718 87562 340954
rect 87646 340718 87882 340954
rect 87326 340398 87562 340634
rect 87646 340398 87882 340634
rect 87326 304718 87562 304954
rect 87646 304718 87882 304954
rect 87326 304398 87562 304634
rect 87646 304398 87882 304634
rect 87326 268718 87562 268954
rect 87646 268718 87882 268954
rect 87326 268398 87562 268634
rect 87646 268398 87882 268634
rect 87326 232718 87562 232954
rect 87646 232718 87882 232954
rect 87326 232398 87562 232634
rect 87646 232398 87882 232634
rect 87326 196718 87562 196954
rect 87646 196718 87882 196954
rect 87326 196398 87562 196634
rect 87646 196398 87882 196634
rect 87326 160718 87562 160954
rect 87646 160718 87882 160954
rect 87326 160398 87562 160634
rect 87646 160398 87882 160634
rect 87326 124718 87562 124954
rect 87646 124718 87882 124954
rect 87326 124398 87562 124634
rect 87646 124398 87882 124634
rect 87326 88718 87562 88954
rect 87646 88718 87882 88954
rect 87326 88398 87562 88634
rect 87646 88398 87882 88634
rect 87326 52718 87562 52954
rect 87646 52718 87882 52954
rect 87326 52398 87562 52634
rect 87646 52398 87882 52634
rect 87326 16718 87562 16954
rect 87646 16718 87882 16954
rect 87326 16398 87562 16634
rect 87646 16398 87882 16634
rect 87326 -3462 87562 -3226
rect 87646 -3462 87882 -3226
rect 87326 -3782 87562 -3546
rect 87646 -3782 87882 -3546
rect 91826 708442 92062 708678
rect 92146 708442 92382 708678
rect 91826 708122 92062 708358
rect 92146 708122 92382 708358
rect 91826 669218 92062 669454
rect 92146 669218 92382 669454
rect 91826 668898 92062 669134
rect 92146 668898 92382 669134
rect 96326 709402 96562 709638
rect 96646 709402 96882 709638
rect 96326 709082 96562 709318
rect 96646 709082 96882 709318
rect 96326 673718 96562 673954
rect 96646 673718 96882 673954
rect 96326 673398 96562 673634
rect 96646 673398 96882 673634
rect 91826 633218 92062 633454
rect 92146 633218 92382 633454
rect 91826 632898 92062 633134
rect 92146 632898 92382 633134
rect 91826 597218 92062 597454
rect 92146 597218 92382 597454
rect 91826 596898 92062 597134
rect 92146 596898 92382 597134
rect 91826 561218 92062 561454
rect 92146 561218 92382 561454
rect 91826 560898 92062 561134
rect 92146 560898 92382 561134
rect 91826 525218 92062 525454
rect 92146 525218 92382 525454
rect 91826 524898 92062 525134
rect 92146 524898 92382 525134
rect 91826 489218 92062 489454
rect 92146 489218 92382 489454
rect 91826 488898 92062 489134
rect 92146 488898 92382 489134
rect 91826 453218 92062 453454
rect 92146 453218 92382 453454
rect 91826 452898 92062 453134
rect 92146 452898 92382 453134
rect 91826 417218 92062 417454
rect 92146 417218 92382 417454
rect 91826 416898 92062 417134
rect 92146 416898 92382 417134
rect 91826 381218 92062 381454
rect 92146 381218 92382 381454
rect 91826 380898 92062 381134
rect 92146 380898 92382 381134
rect 91826 345218 92062 345454
rect 92146 345218 92382 345454
rect 91826 344898 92062 345134
rect 92146 344898 92382 345134
rect 91826 309218 92062 309454
rect 92146 309218 92382 309454
rect 91826 308898 92062 309134
rect 92146 308898 92382 309134
rect 91826 273218 92062 273454
rect 92146 273218 92382 273454
rect 91826 272898 92062 273134
rect 92146 272898 92382 273134
rect 91826 237218 92062 237454
rect 92146 237218 92382 237454
rect 91826 236898 92062 237134
rect 92146 236898 92382 237134
rect 91826 201218 92062 201454
rect 92146 201218 92382 201454
rect 91826 200898 92062 201134
rect 92146 200898 92382 201134
rect 96326 637718 96562 637954
rect 96646 637718 96882 637954
rect 96326 637398 96562 637634
rect 96646 637398 96882 637634
rect 96326 601718 96562 601954
rect 96646 601718 96882 601954
rect 96326 601398 96562 601634
rect 96646 601398 96882 601634
rect 96326 565718 96562 565954
rect 96646 565718 96882 565954
rect 96326 565398 96562 565634
rect 96646 565398 96882 565634
rect 96326 529718 96562 529954
rect 96646 529718 96882 529954
rect 96326 529398 96562 529634
rect 96646 529398 96882 529634
rect 96326 493718 96562 493954
rect 96646 493718 96882 493954
rect 96326 493398 96562 493634
rect 96646 493398 96882 493634
rect 96326 457718 96562 457954
rect 96646 457718 96882 457954
rect 96326 457398 96562 457634
rect 96646 457398 96882 457634
rect 96326 421718 96562 421954
rect 96646 421718 96882 421954
rect 96326 421398 96562 421634
rect 96646 421398 96882 421634
rect 96326 385718 96562 385954
rect 96646 385718 96882 385954
rect 96326 385398 96562 385634
rect 96646 385398 96882 385634
rect 96326 349718 96562 349954
rect 96646 349718 96882 349954
rect 96326 349398 96562 349634
rect 96646 349398 96882 349634
rect 96326 313718 96562 313954
rect 96646 313718 96882 313954
rect 96326 313398 96562 313634
rect 96646 313398 96882 313634
rect 96326 277718 96562 277954
rect 96646 277718 96882 277954
rect 96326 277398 96562 277634
rect 96646 277398 96882 277634
rect 96326 241718 96562 241954
rect 96646 241718 96882 241954
rect 96326 241398 96562 241634
rect 96646 241398 96882 241634
rect 96326 205718 96562 205954
rect 96646 205718 96882 205954
rect 96326 205398 96562 205634
rect 96646 205398 96882 205634
rect 91826 165218 92062 165454
rect 92146 165218 92382 165454
rect 91826 164898 92062 165134
rect 92146 164898 92382 165134
rect 91826 129218 92062 129454
rect 92146 129218 92382 129454
rect 91826 128898 92062 129134
rect 92146 128898 92382 129134
rect 91826 93218 92062 93454
rect 92146 93218 92382 93454
rect 91826 92898 92062 93134
rect 92146 92898 92382 93134
rect 91826 57218 92062 57454
rect 92146 57218 92382 57454
rect 91826 56898 92062 57134
rect 92146 56898 92382 57134
rect 91826 21218 92062 21454
rect 92146 21218 92382 21454
rect 91826 20898 92062 21134
rect 92146 20898 92382 21134
rect 91826 -4422 92062 -4186
rect 92146 -4422 92382 -4186
rect 91826 -4742 92062 -4506
rect 92146 -4742 92382 -4506
rect 100826 710362 101062 710598
rect 101146 710362 101382 710598
rect 100826 710042 101062 710278
rect 101146 710042 101382 710278
rect 100826 678218 101062 678454
rect 101146 678218 101382 678454
rect 100826 677898 101062 678134
rect 101146 677898 101382 678134
rect 100826 642218 101062 642454
rect 101146 642218 101382 642454
rect 100826 641898 101062 642134
rect 101146 641898 101382 642134
rect 100826 606218 101062 606454
rect 101146 606218 101382 606454
rect 100826 605898 101062 606134
rect 101146 605898 101382 606134
rect 100826 570218 101062 570454
rect 101146 570218 101382 570454
rect 100826 569898 101062 570134
rect 101146 569898 101382 570134
rect 100826 534218 101062 534454
rect 101146 534218 101382 534454
rect 100826 533898 101062 534134
rect 101146 533898 101382 534134
rect 100826 498218 101062 498454
rect 101146 498218 101382 498454
rect 100826 497898 101062 498134
rect 101146 497898 101382 498134
rect 100826 462218 101062 462454
rect 101146 462218 101382 462454
rect 100826 461898 101062 462134
rect 101146 461898 101382 462134
rect 100826 426218 101062 426454
rect 101146 426218 101382 426454
rect 100826 425898 101062 426134
rect 101146 425898 101382 426134
rect 100826 390218 101062 390454
rect 101146 390218 101382 390454
rect 100826 389898 101062 390134
rect 101146 389898 101382 390134
rect 100826 354218 101062 354454
rect 101146 354218 101382 354454
rect 100826 353898 101062 354134
rect 101146 353898 101382 354134
rect 100826 318218 101062 318454
rect 101146 318218 101382 318454
rect 100826 317898 101062 318134
rect 101146 317898 101382 318134
rect 100826 282218 101062 282454
rect 101146 282218 101382 282454
rect 100826 281898 101062 282134
rect 101146 281898 101382 282134
rect 100826 246218 101062 246454
rect 101146 246218 101382 246454
rect 100826 245898 101062 246134
rect 101146 245898 101382 246134
rect 100826 210218 101062 210454
rect 101146 210218 101382 210454
rect 100826 209898 101062 210134
rect 101146 209898 101382 210134
rect 96326 169718 96562 169954
rect 96646 169718 96882 169954
rect 96326 169398 96562 169634
rect 96646 169398 96882 169634
rect 96326 133718 96562 133954
rect 96646 133718 96882 133954
rect 96326 133398 96562 133634
rect 96646 133398 96882 133634
rect 96326 97718 96562 97954
rect 96646 97718 96882 97954
rect 96326 97398 96562 97634
rect 96646 97398 96882 97634
rect 105326 711322 105562 711558
rect 105646 711322 105882 711558
rect 105326 711002 105562 711238
rect 105646 711002 105882 711238
rect 105326 682718 105562 682954
rect 105646 682718 105882 682954
rect 105326 682398 105562 682634
rect 105646 682398 105882 682634
rect 105326 646718 105562 646954
rect 105646 646718 105882 646954
rect 105326 646398 105562 646634
rect 105646 646398 105882 646634
rect 105326 610718 105562 610954
rect 105646 610718 105882 610954
rect 105326 610398 105562 610634
rect 105646 610398 105882 610634
rect 105326 574718 105562 574954
rect 105646 574718 105882 574954
rect 105326 574398 105562 574634
rect 105646 574398 105882 574634
rect 105326 538718 105562 538954
rect 105646 538718 105882 538954
rect 105326 538398 105562 538634
rect 105646 538398 105882 538634
rect 105326 502718 105562 502954
rect 105646 502718 105882 502954
rect 105326 502398 105562 502634
rect 105646 502398 105882 502634
rect 105326 466718 105562 466954
rect 105646 466718 105882 466954
rect 105326 466398 105562 466634
rect 105646 466398 105882 466634
rect 105326 430718 105562 430954
rect 105646 430718 105882 430954
rect 105326 430398 105562 430634
rect 105646 430398 105882 430634
rect 105326 394718 105562 394954
rect 105646 394718 105882 394954
rect 105326 394398 105562 394634
rect 105646 394398 105882 394634
rect 105326 358718 105562 358954
rect 105646 358718 105882 358954
rect 105326 358398 105562 358634
rect 105646 358398 105882 358634
rect 105326 322718 105562 322954
rect 105646 322718 105882 322954
rect 105326 322398 105562 322634
rect 105646 322398 105882 322634
rect 105326 286718 105562 286954
rect 105646 286718 105882 286954
rect 105326 286398 105562 286634
rect 105646 286398 105882 286634
rect 105326 250718 105562 250954
rect 105646 250718 105882 250954
rect 105326 250398 105562 250634
rect 105646 250398 105882 250634
rect 105326 214718 105562 214954
rect 105646 214718 105882 214954
rect 105326 214398 105562 214634
rect 105646 214398 105882 214634
rect 100826 174218 101062 174454
rect 101146 174218 101382 174454
rect 100826 173898 101062 174134
rect 101146 173898 101382 174134
rect 100826 138218 101062 138454
rect 101146 138218 101382 138454
rect 100826 137898 101062 138134
rect 101146 137898 101382 138134
rect 100826 102218 101062 102454
rect 101146 102218 101382 102454
rect 100826 101898 101062 102134
rect 101146 101898 101382 102134
rect 96326 61718 96562 61954
rect 96646 61718 96882 61954
rect 96326 61398 96562 61634
rect 96646 61398 96882 61634
rect 96326 25718 96562 25954
rect 96646 25718 96882 25954
rect 96326 25398 96562 25634
rect 96646 25398 96882 25634
rect 96326 -5382 96562 -5146
rect 96646 -5382 96882 -5146
rect 96326 -5702 96562 -5466
rect 96646 -5702 96882 -5466
rect 109826 704602 110062 704838
rect 110146 704602 110382 704838
rect 109826 704282 110062 704518
rect 110146 704282 110382 704518
rect 109826 687218 110062 687454
rect 110146 687218 110382 687454
rect 109826 686898 110062 687134
rect 110146 686898 110382 687134
rect 109826 651218 110062 651454
rect 110146 651218 110382 651454
rect 109826 650898 110062 651134
rect 110146 650898 110382 651134
rect 109826 615218 110062 615454
rect 110146 615218 110382 615454
rect 109826 614898 110062 615134
rect 110146 614898 110382 615134
rect 109826 579218 110062 579454
rect 110146 579218 110382 579454
rect 109826 578898 110062 579134
rect 110146 578898 110382 579134
rect 109826 543218 110062 543454
rect 110146 543218 110382 543454
rect 109826 542898 110062 543134
rect 110146 542898 110382 543134
rect 109826 507218 110062 507454
rect 110146 507218 110382 507454
rect 109826 506898 110062 507134
rect 110146 506898 110382 507134
rect 109826 471218 110062 471454
rect 110146 471218 110382 471454
rect 109826 470898 110062 471134
rect 110146 470898 110382 471134
rect 109826 435218 110062 435454
rect 110146 435218 110382 435454
rect 109826 434898 110062 435134
rect 110146 434898 110382 435134
rect 109826 399218 110062 399454
rect 110146 399218 110382 399454
rect 109826 398898 110062 399134
rect 110146 398898 110382 399134
rect 109826 363218 110062 363454
rect 110146 363218 110382 363454
rect 109826 362898 110062 363134
rect 110146 362898 110382 363134
rect 109826 327218 110062 327454
rect 110146 327218 110382 327454
rect 109826 326898 110062 327134
rect 110146 326898 110382 327134
rect 109826 291218 110062 291454
rect 110146 291218 110382 291454
rect 109826 290898 110062 291134
rect 110146 290898 110382 291134
rect 109826 255218 110062 255454
rect 110146 255218 110382 255454
rect 109826 254898 110062 255134
rect 110146 254898 110382 255134
rect 109826 219218 110062 219454
rect 110146 219218 110382 219454
rect 109826 218898 110062 219134
rect 110146 218898 110382 219134
rect 105326 178718 105562 178954
rect 105646 178718 105882 178954
rect 105326 178398 105562 178634
rect 105646 178398 105882 178634
rect 105326 142718 105562 142954
rect 105646 142718 105882 142954
rect 105326 142398 105562 142634
rect 105646 142398 105882 142634
rect 105326 106718 105562 106954
rect 105646 106718 105882 106954
rect 105326 106398 105562 106634
rect 105646 106398 105882 106634
rect 100826 66218 101062 66454
rect 101146 66218 101382 66454
rect 100826 65898 101062 66134
rect 101146 65898 101382 66134
rect 100826 30218 101062 30454
rect 101146 30218 101382 30454
rect 100826 29898 101062 30134
rect 101146 29898 101382 30134
rect 100826 -6342 101062 -6106
rect 101146 -6342 101382 -6106
rect 100826 -6662 101062 -6426
rect 101146 -6662 101382 -6426
rect 105326 70718 105562 70954
rect 105646 70718 105882 70954
rect 105326 70398 105562 70634
rect 105646 70398 105882 70634
rect 114326 705562 114562 705798
rect 114646 705562 114882 705798
rect 114326 705242 114562 705478
rect 114646 705242 114882 705478
rect 114326 691718 114562 691954
rect 114646 691718 114882 691954
rect 114326 691398 114562 691634
rect 114646 691398 114882 691634
rect 114326 655718 114562 655954
rect 114646 655718 114882 655954
rect 114326 655398 114562 655634
rect 114646 655398 114882 655634
rect 114326 619718 114562 619954
rect 114646 619718 114882 619954
rect 114326 619398 114562 619634
rect 114646 619398 114882 619634
rect 114326 583718 114562 583954
rect 114646 583718 114882 583954
rect 114326 583398 114562 583634
rect 114646 583398 114882 583634
rect 114326 547718 114562 547954
rect 114646 547718 114882 547954
rect 114326 547398 114562 547634
rect 114646 547398 114882 547634
rect 114326 511718 114562 511954
rect 114646 511718 114882 511954
rect 114326 511398 114562 511634
rect 114646 511398 114882 511634
rect 114326 475718 114562 475954
rect 114646 475718 114882 475954
rect 114326 475398 114562 475634
rect 114646 475398 114882 475634
rect 114326 439718 114562 439954
rect 114646 439718 114882 439954
rect 114326 439398 114562 439634
rect 114646 439398 114882 439634
rect 114326 403718 114562 403954
rect 114646 403718 114882 403954
rect 114326 403398 114562 403634
rect 114646 403398 114882 403634
rect 114326 367718 114562 367954
rect 114646 367718 114882 367954
rect 114326 367398 114562 367634
rect 114646 367398 114882 367634
rect 114326 331718 114562 331954
rect 114646 331718 114882 331954
rect 114326 331398 114562 331634
rect 114646 331398 114882 331634
rect 114326 295718 114562 295954
rect 114646 295718 114882 295954
rect 114326 295398 114562 295634
rect 114646 295398 114882 295634
rect 118826 706522 119062 706758
rect 119146 706522 119382 706758
rect 118826 706202 119062 706438
rect 119146 706202 119382 706438
rect 118826 696218 119062 696454
rect 119146 696218 119382 696454
rect 118826 695898 119062 696134
rect 119146 695898 119382 696134
rect 118826 660218 119062 660454
rect 119146 660218 119382 660454
rect 118826 659898 119062 660134
rect 119146 659898 119382 660134
rect 118826 624218 119062 624454
rect 119146 624218 119382 624454
rect 118826 623898 119062 624134
rect 119146 623898 119382 624134
rect 118826 588218 119062 588454
rect 119146 588218 119382 588454
rect 118826 587898 119062 588134
rect 119146 587898 119382 588134
rect 118826 552218 119062 552454
rect 119146 552218 119382 552454
rect 118826 551898 119062 552134
rect 119146 551898 119382 552134
rect 118826 516218 119062 516454
rect 119146 516218 119382 516454
rect 118826 515898 119062 516134
rect 119146 515898 119382 516134
rect 118826 480218 119062 480454
rect 119146 480218 119382 480454
rect 118826 479898 119062 480134
rect 119146 479898 119382 480134
rect 118826 444218 119062 444454
rect 119146 444218 119382 444454
rect 118826 443898 119062 444134
rect 119146 443898 119382 444134
rect 118826 408218 119062 408454
rect 119146 408218 119382 408454
rect 118826 407898 119062 408134
rect 119146 407898 119382 408134
rect 118826 372218 119062 372454
rect 119146 372218 119382 372454
rect 118826 371898 119062 372134
rect 119146 371898 119382 372134
rect 118826 336218 119062 336454
rect 119146 336218 119382 336454
rect 118826 335898 119062 336134
rect 119146 335898 119382 336134
rect 118826 300218 119062 300454
rect 119146 300218 119382 300454
rect 118826 299898 119062 300134
rect 119146 299898 119382 300134
rect 118826 264218 119062 264454
rect 119146 264218 119382 264454
rect 118826 263898 119062 264134
rect 119146 263898 119382 264134
rect 114326 259718 114562 259954
rect 114646 259718 114882 259954
rect 114326 259398 114562 259634
rect 114646 259398 114882 259634
rect 114326 223718 114562 223954
rect 114646 223718 114882 223954
rect 114326 223398 114562 223634
rect 114646 223398 114882 223634
rect 109826 183218 110062 183454
rect 110146 183218 110382 183454
rect 109826 182898 110062 183134
rect 110146 182898 110382 183134
rect 109826 147218 110062 147454
rect 110146 147218 110382 147454
rect 109826 146898 110062 147134
rect 110146 146898 110382 147134
rect 109826 111218 110062 111454
rect 110146 111218 110382 111454
rect 109826 110898 110062 111134
rect 110146 110898 110382 111134
rect 109826 75218 110062 75454
rect 110146 75218 110382 75454
rect 109826 74898 110062 75134
rect 110146 74898 110382 75134
rect 105326 34718 105562 34954
rect 105646 34718 105882 34954
rect 105326 34398 105562 34634
rect 105646 34398 105882 34634
rect 105326 -7302 105562 -7066
rect 105646 -7302 105882 -7066
rect 105326 -7622 105562 -7386
rect 105646 -7622 105882 -7386
rect 114326 187718 114562 187954
rect 114646 187718 114882 187954
rect 114326 187398 114562 187634
rect 114646 187398 114882 187634
rect 114326 151718 114562 151954
rect 114646 151718 114882 151954
rect 114326 151398 114562 151634
rect 114646 151398 114882 151634
rect 114326 115718 114562 115954
rect 114646 115718 114882 115954
rect 114326 115398 114562 115634
rect 114646 115398 114882 115634
rect 114326 79718 114562 79954
rect 114646 79718 114882 79954
rect 114326 79398 114562 79634
rect 114646 79398 114882 79634
rect 109826 39218 110062 39454
rect 110146 39218 110382 39454
rect 109826 38898 110062 39134
rect 110146 38898 110382 39134
rect 109826 3218 110062 3454
rect 110146 3218 110382 3454
rect 109826 2898 110062 3134
rect 110146 2898 110382 3134
rect 109826 -582 110062 -346
rect 110146 -582 110382 -346
rect 109826 -902 110062 -666
rect 110146 -902 110382 -666
rect 123326 707482 123562 707718
rect 123646 707482 123882 707718
rect 123326 707162 123562 707398
rect 123646 707162 123882 707398
rect 123326 700718 123562 700954
rect 123646 700718 123882 700954
rect 123326 700398 123562 700634
rect 123646 700398 123882 700634
rect 123326 664718 123562 664954
rect 123646 664718 123882 664954
rect 123326 664398 123562 664634
rect 123646 664398 123882 664634
rect 123326 628718 123562 628954
rect 123646 628718 123882 628954
rect 123326 628398 123562 628634
rect 123646 628398 123882 628634
rect 123326 592718 123562 592954
rect 123646 592718 123882 592954
rect 123326 592398 123562 592634
rect 123646 592398 123882 592634
rect 123326 556718 123562 556954
rect 123646 556718 123882 556954
rect 123326 556398 123562 556634
rect 123646 556398 123882 556634
rect 123326 520718 123562 520954
rect 123646 520718 123882 520954
rect 123326 520398 123562 520634
rect 123646 520398 123882 520634
rect 123326 484718 123562 484954
rect 123646 484718 123882 484954
rect 123326 484398 123562 484634
rect 123646 484398 123882 484634
rect 123326 448718 123562 448954
rect 123646 448718 123882 448954
rect 123326 448398 123562 448634
rect 123646 448398 123882 448634
rect 123326 412718 123562 412954
rect 123646 412718 123882 412954
rect 123326 412398 123562 412634
rect 123646 412398 123882 412634
rect 123326 376718 123562 376954
rect 123646 376718 123882 376954
rect 123326 376398 123562 376634
rect 123646 376398 123882 376634
rect 123326 340718 123562 340954
rect 123646 340718 123882 340954
rect 123326 340398 123562 340634
rect 123646 340398 123882 340634
rect 123326 304718 123562 304954
rect 123646 304718 123882 304954
rect 123326 304398 123562 304634
rect 123646 304398 123882 304634
rect 123326 268718 123562 268954
rect 123646 268718 123882 268954
rect 123326 268398 123562 268634
rect 123646 268398 123882 268634
rect 127826 708442 128062 708678
rect 128146 708442 128382 708678
rect 127826 708122 128062 708358
rect 128146 708122 128382 708358
rect 127826 669218 128062 669454
rect 128146 669218 128382 669454
rect 127826 668898 128062 669134
rect 128146 668898 128382 669134
rect 127826 633218 128062 633454
rect 128146 633218 128382 633454
rect 127826 632898 128062 633134
rect 128146 632898 128382 633134
rect 127826 597218 128062 597454
rect 128146 597218 128382 597454
rect 127826 596898 128062 597134
rect 128146 596898 128382 597134
rect 127826 561218 128062 561454
rect 128146 561218 128382 561454
rect 127826 560898 128062 561134
rect 128146 560898 128382 561134
rect 127826 525218 128062 525454
rect 128146 525218 128382 525454
rect 127826 524898 128062 525134
rect 128146 524898 128382 525134
rect 127826 489218 128062 489454
rect 128146 489218 128382 489454
rect 127826 488898 128062 489134
rect 128146 488898 128382 489134
rect 127826 453218 128062 453454
rect 128146 453218 128382 453454
rect 127826 452898 128062 453134
rect 128146 452898 128382 453134
rect 127826 417218 128062 417454
rect 128146 417218 128382 417454
rect 127826 416898 128062 417134
rect 128146 416898 128382 417134
rect 127826 381218 128062 381454
rect 128146 381218 128382 381454
rect 127826 380898 128062 381134
rect 128146 380898 128382 381134
rect 127826 345218 128062 345454
rect 128146 345218 128382 345454
rect 127826 344898 128062 345134
rect 128146 344898 128382 345134
rect 127826 309218 128062 309454
rect 128146 309218 128382 309454
rect 127826 308898 128062 309134
rect 128146 308898 128382 309134
rect 127826 273218 128062 273454
rect 128146 273218 128382 273454
rect 127826 272898 128062 273134
rect 128146 272898 128382 273134
rect 132326 709402 132562 709638
rect 132646 709402 132882 709638
rect 132326 709082 132562 709318
rect 132646 709082 132882 709318
rect 132326 673718 132562 673954
rect 132646 673718 132882 673954
rect 132326 673398 132562 673634
rect 132646 673398 132882 673634
rect 132326 637718 132562 637954
rect 132646 637718 132882 637954
rect 132326 637398 132562 637634
rect 132646 637398 132882 637634
rect 132326 601718 132562 601954
rect 132646 601718 132882 601954
rect 132326 601398 132562 601634
rect 132646 601398 132882 601634
rect 132326 565718 132562 565954
rect 132646 565718 132882 565954
rect 132326 565398 132562 565634
rect 132646 565398 132882 565634
rect 132326 529718 132562 529954
rect 132646 529718 132882 529954
rect 132326 529398 132562 529634
rect 132646 529398 132882 529634
rect 132326 493718 132562 493954
rect 132646 493718 132882 493954
rect 132326 493398 132562 493634
rect 132646 493398 132882 493634
rect 132326 457718 132562 457954
rect 132646 457718 132882 457954
rect 132326 457398 132562 457634
rect 132646 457398 132882 457634
rect 132326 421718 132562 421954
rect 132646 421718 132882 421954
rect 132326 421398 132562 421634
rect 132646 421398 132882 421634
rect 132326 385718 132562 385954
rect 132646 385718 132882 385954
rect 132326 385398 132562 385634
rect 132646 385398 132882 385634
rect 132326 349718 132562 349954
rect 132646 349718 132882 349954
rect 132326 349398 132562 349634
rect 132646 349398 132882 349634
rect 132326 313718 132562 313954
rect 132646 313718 132882 313954
rect 132326 313398 132562 313634
rect 132646 313398 132882 313634
rect 132326 277718 132562 277954
rect 132646 277718 132882 277954
rect 132326 277398 132562 277634
rect 132646 277398 132882 277634
rect 136826 710362 137062 710598
rect 137146 710362 137382 710598
rect 136826 710042 137062 710278
rect 137146 710042 137382 710278
rect 136826 678218 137062 678454
rect 137146 678218 137382 678454
rect 136826 677898 137062 678134
rect 137146 677898 137382 678134
rect 136826 642218 137062 642454
rect 137146 642218 137382 642454
rect 136826 641898 137062 642134
rect 137146 641898 137382 642134
rect 136826 606218 137062 606454
rect 137146 606218 137382 606454
rect 136826 605898 137062 606134
rect 137146 605898 137382 606134
rect 136826 570218 137062 570454
rect 137146 570218 137382 570454
rect 136826 569898 137062 570134
rect 137146 569898 137382 570134
rect 136826 534218 137062 534454
rect 137146 534218 137382 534454
rect 136826 533898 137062 534134
rect 137146 533898 137382 534134
rect 136826 498218 137062 498454
rect 137146 498218 137382 498454
rect 136826 497898 137062 498134
rect 137146 497898 137382 498134
rect 136826 462218 137062 462454
rect 137146 462218 137382 462454
rect 136826 461898 137062 462134
rect 137146 461898 137382 462134
rect 136826 426218 137062 426454
rect 137146 426218 137382 426454
rect 136826 425898 137062 426134
rect 137146 425898 137382 426134
rect 136826 390218 137062 390454
rect 137146 390218 137382 390454
rect 136826 389898 137062 390134
rect 137146 389898 137382 390134
rect 136826 354218 137062 354454
rect 137146 354218 137382 354454
rect 136826 353898 137062 354134
rect 137146 353898 137382 354134
rect 136826 318218 137062 318454
rect 137146 318218 137382 318454
rect 136826 317898 137062 318134
rect 137146 317898 137382 318134
rect 136826 282218 137062 282454
rect 137146 282218 137382 282454
rect 136826 281898 137062 282134
rect 137146 281898 137382 282134
rect 141326 711322 141562 711558
rect 141646 711322 141882 711558
rect 141326 711002 141562 711238
rect 141646 711002 141882 711238
rect 141326 682718 141562 682954
rect 141646 682718 141882 682954
rect 141326 682398 141562 682634
rect 141646 682398 141882 682634
rect 141326 646718 141562 646954
rect 141646 646718 141882 646954
rect 141326 646398 141562 646634
rect 141646 646398 141882 646634
rect 141326 610718 141562 610954
rect 141646 610718 141882 610954
rect 141326 610398 141562 610634
rect 141646 610398 141882 610634
rect 141326 574718 141562 574954
rect 141646 574718 141882 574954
rect 141326 574398 141562 574634
rect 141646 574398 141882 574634
rect 141326 538718 141562 538954
rect 141646 538718 141882 538954
rect 141326 538398 141562 538634
rect 141646 538398 141882 538634
rect 141326 502718 141562 502954
rect 141646 502718 141882 502954
rect 141326 502398 141562 502634
rect 141646 502398 141882 502634
rect 141326 466718 141562 466954
rect 141646 466718 141882 466954
rect 141326 466398 141562 466634
rect 141646 466398 141882 466634
rect 141326 430718 141562 430954
rect 141646 430718 141882 430954
rect 141326 430398 141562 430634
rect 141646 430398 141882 430634
rect 141326 394718 141562 394954
rect 141646 394718 141882 394954
rect 141326 394398 141562 394634
rect 141646 394398 141882 394634
rect 141326 358718 141562 358954
rect 141646 358718 141882 358954
rect 141326 358398 141562 358634
rect 141646 358398 141882 358634
rect 141326 322718 141562 322954
rect 141646 322718 141882 322954
rect 141326 322398 141562 322634
rect 141646 322398 141882 322634
rect 141326 286718 141562 286954
rect 141646 286718 141882 286954
rect 141326 286398 141562 286634
rect 141646 286398 141882 286634
rect 145826 704602 146062 704838
rect 146146 704602 146382 704838
rect 145826 704282 146062 704518
rect 146146 704282 146382 704518
rect 145826 687218 146062 687454
rect 146146 687218 146382 687454
rect 145826 686898 146062 687134
rect 146146 686898 146382 687134
rect 145826 651218 146062 651454
rect 146146 651218 146382 651454
rect 145826 650898 146062 651134
rect 146146 650898 146382 651134
rect 145826 615218 146062 615454
rect 146146 615218 146382 615454
rect 145826 614898 146062 615134
rect 146146 614898 146382 615134
rect 145826 579218 146062 579454
rect 146146 579218 146382 579454
rect 145826 578898 146062 579134
rect 146146 578898 146382 579134
rect 145826 543218 146062 543454
rect 146146 543218 146382 543454
rect 145826 542898 146062 543134
rect 146146 542898 146382 543134
rect 145826 507218 146062 507454
rect 146146 507218 146382 507454
rect 145826 506898 146062 507134
rect 146146 506898 146382 507134
rect 145826 471218 146062 471454
rect 146146 471218 146382 471454
rect 145826 470898 146062 471134
rect 146146 470898 146382 471134
rect 145826 435218 146062 435454
rect 146146 435218 146382 435454
rect 145826 434898 146062 435134
rect 146146 434898 146382 435134
rect 145826 399218 146062 399454
rect 146146 399218 146382 399454
rect 145826 398898 146062 399134
rect 146146 398898 146382 399134
rect 145826 363218 146062 363454
rect 146146 363218 146382 363454
rect 145826 362898 146062 363134
rect 146146 362898 146382 363134
rect 145826 327218 146062 327454
rect 146146 327218 146382 327454
rect 145826 326898 146062 327134
rect 146146 326898 146382 327134
rect 145826 291218 146062 291454
rect 146146 291218 146382 291454
rect 145826 290898 146062 291134
rect 146146 290898 146382 291134
rect 150326 705562 150562 705798
rect 150646 705562 150882 705798
rect 150326 705242 150562 705478
rect 150646 705242 150882 705478
rect 150326 691718 150562 691954
rect 150646 691718 150882 691954
rect 150326 691398 150562 691634
rect 150646 691398 150882 691634
rect 150326 655718 150562 655954
rect 150646 655718 150882 655954
rect 150326 655398 150562 655634
rect 150646 655398 150882 655634
rect 150326 619718 150562 619954
rect 150646 619718 150882 619954
rect 150326 619398 150562 619634
rect 150646 619398 150882 619634
rect 150326 583718 150562 583954
rect 150646 583718 150882 583954
rect 150326 583398 150562 583634
rect 150646 583398 150882 583634
rect 150326 547718 150562 547954
rect 150646 547718 150882 547954
rect 150326 547398 150562 547634
rect 150646 547398 150882 547634
rect 150326 511718 150562 511954
rect 150646 511718 150882 511954
rect 150326 511398 150562 511634
rect 150646 511398 150882 511634
rect 150326 475718 150562 475954
rect 150646 475718 150882 475954
rect 150326 475398 150562 475634
rect 150646 475398 150882 475634
rect 150326 439718 150562 439954
rect 150646 439718 150882 439954
rect 150326 439398 150562 439634
rect 150646 439398 150882 439634
rect 150326 403718 150562 403954
rect 150646 403718 150882 403954
rect 150326 403398 150562 403634
rect 150646 403398 150882 403634
rect 150326 367718 150562 367954
rect 150646 367718 150882 367954
rect 150326 367398 150562 367634
rect 150646 367398 150882 367634
rect 150326 331718 150562 331954
rect 150646 331718 150882 331954
rect 150326 331398 150562 331634
rect 150646 331398 150882 331634
rect 150326 295718 150562 295954
rect 150646 295718 150882 295954
rect 150326 295398 150562 295634
rect 150646 295398 150882 295634
rect 154826 706522 155062 706758
rect 155146 706522 155382 706758
rect 154826 706202 155062 706438
rect 155146 706202 155382 706438
rect 154826 696218 155062 696454
rect 155146 696218 155382 696454
rect 154826 695898 155062 696134
rect 155146 695898 155382 696134
rect 154826 660218 155062 660454
rect 155146 660218 155382 660454
rect 154826 659898 155062 660134
rect 155146 659898 155382 660134
rect 154826 624218 155062 624454
rect 155146 624218 155382 624454
rect 154826 623898 155062 624134
rect 155146 623898 155382 624134
rect 154826 588218 155062 588454
rect 155146 588218 155382 588454
rect 154826 587898 155062 588134
rect 155146 587898 155382 588134
rect 154826 552218 155062 552454
rect 155146 552218 155382 552454
rect 154826 551898 155062 552134
rect 155146 551898 155382 552134
rect 154826 516218 155062 516454
rect 155146 516218 155382 516454
rect 154826 515898 155062 516134
rect 155146 515898 155382 516134
rect 154826 480218 155062 480454
rect 155146 480218 155382 480454
rect 154826 479898 155062 480134
rect 155146 479898 155382 480134
rect 154826 444218 155062 444454
rect 155146 444218 155382 444454
rect 154826 443898 155062 444134
rect 155146 443898 155382 444134
rect 154826 408218 155062 408454
rect 155146 408218 155382 408454
rect 154826 407898 155062 408134
rect 155146 407898 155382 408134
rect 154826 372218 155062 372454
rect 155146 372218 155382 372454
rect 154826 371898 155062 372134
rect 155146 371898 155382 372134
rect 154826 336218 155062 336454
rect 155146 336218 155382 336454
rect 154826 335898 155062 336134
rect 155146 335898 155382 336134
rect 154826 300218 155062 300454
rect 155146 300218 155382 300454
rect 154826 299898 155062 300134
rect 155146 299898 155382 300134
rect 154826 264218 155062 264454
rect 155146 264218 155382 264454
rect 154826 263898 155062 264134
rect 155146 263898 155382 264134
rect 159326 707482 159562 707718
rect 159646 707482 159882 707718
rect 159326 707162 159562 707398
rect 159646 707162 159882 707398
rect 159326 700718 159562 700954
rect 159646 700718 159882 700954
rect 159326 700398 159562 700634
rect 159646 700398 159882 700634
rect 159326 664718 159562 664954
rect 159646 664718 159882 664954
rect 159326 664398 159562 664634
rect 159646 664398 159882 664634
rect 159326 628718 159562 628954
rect 159646 628718 159882 628954
rect 159326 628398 159562 628634
rect 159646 628398 159882 628634
rect 159326 592718 159562 592954
rect 159646 592718 159882 592954
rect 159326 592398 159562 592634
rect 159646 592398 159882 592634
rect 159326 556718 159562 556954
rect 159646 556718 159882 556954
rect 159326 556398 159562 556634
rect 159646 556398 159882 556634
rect 159326 520718 159562 520954
rect 159646 520718 159882 520954
rect 159326 520398 159562 520634
rect 159646 520398 159882 520634
rect 159326 484718 159562 484954
rect 159646 484718 159882 484954
rect 159326 484398 159562 484634
rect 159646 484398 159882 484634
rect 159326 448718 159562 448954
rect 159646 448718 159882 448954
rect 159326 448398 159562 448634
rect 159646 448398 159882 448634
rect 159326 412718 159562 412954
rect 159646 412718 159882 412954
rect 159326 412398 159562 412634
rect 159646 412398 159882 412634
rect 159326 376718 159562 376954
rect 159646 376718 159882 376954
rect 159326 376398 159562 376634
rect 159646 376398 159882 376634
rect 159326 340718 159562 340954
rect 159646 340718 159882 340954
rect 159326 340398 159562 340634
rect 159646 340398 159882 340634
rect 159326 304718 159562 304954
rect 159646 304718 159882 304954
rect 159326 304398 159562 304634
rect 159646 304398 159882 304634
rect 159326 268718 159562 268954
rect 159646 268718 159882 268954
rect 159326 268398 159562 268634
rect 159646 268398 159882 268634
rect 163826 708442 164062 708678
rect 164146 708442 164382 708678
rect 163826 708122 164062 708358
rect 164146 708122 164382 708358
rect 163826 669218 164062 669454
rect 164146 669218 164382 669454
rect 163826 668898 164062 669134
rect 164146 668898 164382 669134
rect 163826 633218 164062 633454
rect 164146 633218 164382 633454
rect 163826 632898 164062 633134
rect 164146 632898 164382 633134
rect 163826 597218 164062 597454
rect 164146 597218 164382 597454
rect 163826 596898 164062 597134
rect 164146 596898 164382 597134
rect 163826 561218 164062 561454
rect 164146 561218 164382 561454
rect 163826 560898 164062 561134
rect 164146 560898 164382 561134
rect 163826 525218 164062 525454
rect 164146 525218 164382 525454
rect 163826 524898 164062 525134
rect 164146 524898 164382 525134
rect 163826 489218 164062 489454
rect 164146 489218 164382 489454
rect 163826 488898 164062 489134
rect 164146 488898 164382 489134
rect 163826 453218 164062 453454
rect 164146 453218 164382 453454
rect 163826 452898 164062 453134
rect 164146 452898 164382 453134
rect 163826 417218 164062 417454
rect 164146 417218 164382 417454
rect 163826 416898 164062 417134
rect 164146 416898 164382 417134
rect 163826 381218 164062 381454
rect 164146 381218 164382 381454
rect 163826 380898 164062 381134
rect 164146 380898 164382 381134
rect 163826 345218 164062 345454
rect 164146 345218 164382 345454
rect 163826 344898 164062 345134
rect 164146 344898 164382 345134
rect 163826 309218 164062 309454
rect 164146 309218 164382 309454
rect 163826 308898 164062 309134
rect 164146 308898 164382 309134
rect 163826 273218 164062 273454
rect 164146 273218 164382 273454
rect 163826 272898 164062 273134
rect 164146 272898 164382 273134
rect 168326 709402 168562 709638
rect 168646 709402 168882 709638
rect 168326 709082 168562 709318
rect 168646 709082 168882 709318
rect 168326 673718 168562 673954
rect 168646 673718 168882 673954
rect 168326 673398 168562 673634
rect 168646 673398 168882 673634
rect 168326 637718 168562 637954
rect 168646 637718 168882 637954
rect 168326 637398 168562 637634
rect 168646 637398 168882 637634
rect 168326 601718 168562 601954
rect 168646 601718 168882 601954
rect 168326 601398 168562 601634
rect 168646 601398 168882 601634
rect 168326 565718 168562 565954
rect 168646 565718 168882 565954
rect 168326 565398 168562 565634
rect 168646 565398 168882 565634
rect 168326 529718 168562 529954
rect 168646 529718 168882 529954
rect 168326 529398 168562 529634
rect 168646 529398 168882 529634
rect 168326 493718 168562 493954
rect 168646 493718 168882 493954
rect 168326 493398 168562 493634
rect 168646 493398 168882 493634
rect 168326 457718 168562 457954
rect 168646 457718 168882 457954
rect 168326 457398 168562 457634
rect 168646 457398 168882 457634
rect 168326 421718 168562 421954
rect 168646 421718 168882 421954
rect 168326 421398 168562 421634
rect 168646 421398 168882 421634
rect 168326 385718 168562 385954
rect 168646 385718 168882 385954
rect 168326 385398 168562 385634
rect 168646 385398 168882 385634
rect 168326 349718 168562 349954
rect 168646 349718 168882 349954
rect 168326 349398 168562 349634
rect 168646 349398 168882 349634
rect 168326 313718 168562 313954
rect 168646 313718 168882 313954
rect 168326 313398 168562 313634
rect 168646 313398 168882 313634
rect 168326 277718 168562 277954
rect 168646 277718 168882 277954
rect 168326 277398 168562 277634
rect 168646 277398 168882 277634
rect 172826 710362 173062 710598
rect 173146 710362 173382 710598
rect 172826 710042 173062 710278
rect 173146 710042 173382 710278
rect 172826 678218 173062 678454
rect 173146 678218 173382 678454
rect 172826 677898 173062 678134
rect 173146 677898 173382 678134
rect 172826 642218 173062 642454
rect 173146 642218 173382 642454
rect 172826 641898 173062 642134
rect 173146 641898 173382 642134
rect 172826 606218 173062 606454
rect 173146 606218 173382 606454
rect 172826 605898 173062 606134
rect 173146 605898 173382 606134
rect 172826 570218 173062 570454
rect 173146 570218 173382 570454
rect 172826 569898 173062 570134
rect 173146 569898 173382 570134
rect 172826 534218 173062 534454
rect 173146 534218 173382 534454
rect 172826 533898 173062 534134
rect 173146 533898 173382 534134
rect 172826 498218 173062 498454
rect 173146 498218 173382 498454
rect 172826 497898 173062 498134
rect 173146 497898 173382 498134
rect 172826 462218 173062 462454
rect 173146 462218 173382 462454
rect 172826 461898 173062 462134
rect 173146 461898 173382 462134
rect 172826 426218 173062 426454
rect 173146 426218 173382 426454
rect 172826 425898 173062 426134
rect 173146 425898 173382 426134
rect 172826 390218 173062 390454
rect 173146 390218 173382 390454
rect 172826 389898 173062 390134
rect 173146 389898 173382 390134
rect 172826 354218 173062 354454
rect 173146 354218 173382 354454
rect 172826 353898 173062 354134
rect 173146 353898 173382 354134
rect 172826 318218 173062 318454
rect 173146 318218 173382 318454
rect 172826 317898 173062 318134
rect 173146 317898 173382 318134
rect 172826 282218 173062 282454
rect 173146 282218 173382 282454
rect 172826 281898 173062 282134
rect 173146 281898 173382 282134
rect 177326 711322 177562 711558
rect 177646 711322 177882 711558
rect 177326 711002 177562 711238
rect 177646 711002 177882 711238
rect 177326 682718 177562 682954
rect 177646 682718 177882 682954
rect 177326 682398 177562 682634
rect 177646 682398 177882 682634
rect 177326 646718 177562 646954
rect 177646 646718 177882 646954
rect 177326 646398 177562 646634
rect 177646 646398 177882 646634
rect 177326 610718 177562 610954
rect 177646 610718 177882 610954
rect 177326 610398 177562 610634
rect 177646 610398 177882 610634
rect 177326 574718 177562 574954
rect 177646 574718 177882 574954
rect 177326 574398 177562 574634
rect 177646 574398 177882 574634
rect 177326 538718 177562 538954
rect 177646 538718 177882 538954
rect 177326 538398 177562 538634
rect 177646 538398 177882 538634
rect 177326 502718 177562 502954
rect 177646 502718 177882 502954
rect 177326 502398 177562 502634
rect 177646 502398 177882 502634
rect 177326 466718 177562 466954
rect 177646 466718 177882 466954
rect 177326 466398 177562 466634
rect 177646 466398 177882 466634
rect 177326 430718 177562 430954
rect 177646 430718 177882 430954
rect 177326 430398 177562 430634
rect 177646 430398 177882 430634
rect 177326 394718 177562 394954
rect 177646 394718 177882 394954
rect 177326 394398 177562 394634
rect 177646 394398 177882 394634
rect 177326 358718 177562 358954
rect 177646 358718 177882 358954
rect 177326 358398 177562 358634
rect 177646 358398 177882 358634
rect 177326 322718 177562 322954
rect 177646 322718 177882 322954
rect 177326 322398 177562 322634
rect 177646 322398 177882 322634
rect 177326 286718 177562 286954
rect 177646 286718 177882 286954
rect 177326 286398 177562 286634
rect 177646 286398 177882 286634
rect 181826 704602 182062 704838
rect 182146 704602 182382 704838
rect 181826 704282 182062 704518
rect 182146 704282 182382 704518
rect 181826 687218 182062 687454
rect 182146 687218 182382 687454
rect 181826 686898 182062 687134
rect 182146 686898 182382 687134
rect 181826 651218 182062 651454
rect 182146 651218 182382 651454
rect 181826 650898 182062 651134
rect 182146 650898 182382 651134
rect 181826 615218 182062 615454
rect 182146 615218 182382 615454
rect 181826 614898 182062 615134
rect 182146 614898 182382 615134
rect 181826 579218 182062 579454
rect 182146 579218 182382 579454
rect 181826 578898 182062 579134
rect 182146 578898 182382 579134
rect 181826 543218 182062 543454
rect 182146 543218 182382 543454
rect 181826 542898 182062 543134
rect 182146 542898 182382 543134
rect 181826 507218 182062 507454
rect 182146 507218 182382 507454
rect 181826 506898 182062 507134
rect 182146 506898 182382 507134
rect 181826 471218 182062 471454
rect 182146 471218 182382 471454
rect 181826 470898 182062 471134
rect 182146 470898 182382 471134
rect 181826 435218 182062 435454
rect 182146 435218 182382 435454
rect 181826 434898 182062 435134
rect 182146 434898 182382 435134
rect 181826 399218 182062 399454
rect 182146 399218 182382 399454
rect 181826 398898 182062 399134
rect 182146 398898 182382 399134
rect 181826 363218 182062 363454
rect 182146 363218 182382 363454
rect 181826 362898 182062 363134
rect 182146 362898 182382 363134
rect 181826 327218 182062 327454
rect 182146 327218 182382 327454
rect 181826 326898 182062 327134
rect 182146 326898 182382 327134
rect 181826 291218 182062 291454
rect 182146 291218 182382 291454
rect 181826 290898 182062 291134
rect 182146 290898 182382 291134
rect 186326 705562 186562 705798
rect 186646 705562 186882 705798
rect 186326 705242 186562 705478
rect 186646 705242 186882 705478
rect 186326 691718 186562 691954
rect 186646 691718 186882 691954
rect 186326 691398 186562 691634
rect 186646 691398 186882 691634
rect 186326 655718 186562 655954
rect 186646 655718 186882 655954
rect 186326 655398 186562 655634
rect 186646 655398 186882 655634
rect 186326 619718 186562 619954
rect 186646 619718 186882 619954
rect 186326 619398 186562 619634
rect 186646 619398 186882 619634
rect 186326 583718 186562 583954
rect 186646 583718 186882 583954
rect 186326 583398 186562 583634
rect 186646 583398 186882 583634
rect 186326 547718 186562 547954
rect 186646 547718 186882 547954
rect 186326 547398 186562 547634
rect 186646 547398 186882 547634
rect 186326 511718 186562 511954
rect 186646 511718 186882 511954
rect 186326 511398 186562 511634
rect 186646 511398 186882 511634
rect 186326 475718 186562 475954
rect 186646 475718 186882 475954
rect 186326 475398 186562 475634
rect 186646 475398 186882 475634
rect 186326 439718 186562 439954
rect 186646 439718 186882 439954
rect 186326 439398 186562 439634
rect 186646 439398 186882 439634
rect 186326 403718 186562 403954
rect 186646 403718 186882 403954
rect 186326 403398 186562 403634
rect 186646 403398 186882 403634
rect 186326 367718 186562 367954
rect 186646 367718 186882 367954
rect 186326 367398 186562 367634
rect 186646 367398 186882 367634
rect 186326 331718 186562 331954
rect 186646 331718 186882 331954
rect 186326 331398 186562 331634
rect 186646 331398 186882 331634
rect 186326 295718 186562 295954
rect 186646 295718 186882 295954
rect 186326 295398 186562 295634
rect 186646 295398 186882 295634
rect 190826 706522 191062 706758
rect 191146 706522 191382 706758
rect 190826 706202 191062 706438
rect 191146 706202 191382 706438
rect 190826 696218 191062 696454
rect 191146 696218 191382 696454
rect 190826 695898 191062 696134
rect 191146 695898 191382 696134
rect 190826 660218 191062 660454
rect 191146 660218 191382 660454
rect 190826 659898 191062 660134
rect 191146 659898 191382 660134
rect 190826 624218 191062 624454
rect 191146 624218 191382 624454
rect 190826 623898 191062 624134
rect 191146 623898 191382 624134
rect 190826 588218 191062 588454
rect 191146 588218 191382 588454
rect 190826 587898 191062 588134
rect 191146 587898 191382 588134
rect 190826 552218 191062 552454
rect 191146 552218 191382 552454
rect 190826 551898 191062 552134
rect 191146 551898 191382 552134
rect 190826 516218 191062 516454
rect 191146 516218 191382 516454
rect 190826 515898 191062 516134
rect 191146 515898 191382 516134
rect 190826 480218 191062 480454
rect 191146 480218 191382 480454
rect 190826 479898 191062 480134
rect 191146 479898 191382 480134
rect 190826 444218 191062 444454
rect 191146 444218 191382 444454
rect 190826 443898 191062 444134
rect 191146 443898 191382 444134
rect 190826 408218 191062 408454
rect 191146 408218 191382 408454
rect 190826 407898 191062 408134
rect 191146 407898 191382 408134
rect 190826 372218 191062 372454
rect 191146 372218 191382 372454
rect 190826 371898 191062 372134
rect 191146 371898 191382 372134
rect 190826 336218 191062 336454
rect 191146 336218 191382 336454
rect 190826 335898 191062 336134
rect 191146 335898 191382 336134
rect 190826 300218 191062 300454
rect 191146 300218 191382 300454
rect 190826 299898 191062 300134
rect 191146 299898 191382 300134
rect 190826 264218 191062 264454
rect 191146 264218 191382 264454
rect 190826 263898 191062 264134
rect 191146 263898 191382 264134
rect 195326 707482 195562 707718
rect 195646 707482 195882 707718
rect 195326 707162 195562 707398
rect 195646 707162 195882 707398
rect 195326 700718 195562 700954
rect 195646 700718 195882 700954
rect 195326 700398 195562 700634
rect 195646 700398 195882 700634
rect 195326 664718 195562 664954
rect 195646 664718 195882 664954
rect 195326 664398 195562 664634
rect 195646 664398 195882 664634
rect 195326 628718 195562 628954
rect 195646 628718 195882 628954
rect 195326 628398 195562 628634
rect 195646 628398 195882 628634
rect 195326 592718 195562 592954
rect 195646 592718 195882 592954
rect 195326 592398 195562 592634
rect 195646 592398 195882 592634
rect 195326 556718 195562 556954
rect 195646 556718 195882 556954
rect 195326 556398 195562 556634
rect 195646 556398 195882 556634
rect 195326 520718 195562 520954
rect 195646 520718 195882 520954
rect 195326 520398 195562 520634
rect 195646 520398 195882 520634
rect 195326 484718 195562 484954
rect 195646 484718 195882 484954
rect 195326 484398 195562 484634
rect 195646 484398 195882 484634
rect 195326 448718 195562 448954
rect 195646 448718 195882 448954
rect 195326 448398 195562 448634
rect 195646 448398 195882 448634
rect 195326 412718 195562 412954
rect 195646 412718 195882 412954
rect 195326 412398 195562 412634
rect 195646 412398 195882 412634
rect 195326 376718 195562 376954
rect 195646 376718 195882 376954
rect 195326 376398 195562 376634
rect 195646 376398 195882 376634
rect 195326 340718 195562 340954
rect 195646 340718 195882 340954
rect 195326 340398 195562 340634
rect 195646 340398 195882 340634
rect 195326 304718 195562 304954
rect 195646 304718 195882 304954
rect 195326 304398 195562 304634
rect 195646 304398 195882 304634
rect 195326 268718 195562 268954
rect 195646 268718 195882 268954
rect 195326 268398 195562 268634
rect 195646 268398 195882 268634
rect 118826 192218 119062 192454
rect 119146 192218 119382 192454
rect 118826 191898 119062 192134
rect 119146 191898 119382 192134
rect 118826 156218 119062 156454
rect 119146 156218 119382 156454
rect 118826 155898 119062 156134
rect 119146 155898 119382 156134
rect 114326 43718 114562 43954
rect 114646 43718 114882 43954
rect 114326 43398 114562 43634
rect 114646 43398 114882 43634
rect 114326 7718 114562 7954
rect 114646 7718 114882 7954
rect 114326 7398 114562 7634
rect 114646 7398 114882 7634
rect 114326 -1542 114562 -1306
rect 114646 -1542 114882 -1306
rect 114326 -1862 114562 -1626
rect 114646 -1862 114882 -1626
rect 124250 255218 124486 255454
rect 124250 254898 124486 255134
rect 154970 255218 155206 255454
rect 154970 254898 155206 255134
rect 185690 255218 185926 255454
rect 185690 254898 185926 255134
rect 139610 223718 139846 223954
rect 139610 223398 139846 223634
rect 170330 223718 170566 223954
rect 170330 223398 170566 223634
rect 124250 219218 124486 219454
rect 124250 218898 124486 219134
rect 154970 219218 155206 219454
rect 154970 218898 155206 219134
rect 185690 219218 185926 219454
rect 185690 218898 185926 219134
rect 123326 196718 123562 196954
rect 123646 196718 123882 196954
rect 123326 196398 123562 196634
rect 123646 196398 123882 196634
rect 123326 160718 123562 160954
rect 123646 160718 123882 160954
rect 123326 160398 123562 160634
rect 123646 160398 123882 160634
rect 141326 178718 141562 178954
rect 141646 178718 141882 178954
rect 141326 178398 141562 178634
rect 141646 178398 141882 178634
rect 145826 183218 146062 183454
rect 146146 183218 146382 183454
rect 145826 182898 146062 183134
rect 146146 182898 146382 183134
rect 141326 142718 141562 142954
rect 141646 142718 141882 142954
rect 141326 142398 141562 142634
rect 141646 142398 141882 142634
rect 150326 187718 150562 187954
rect 150646 187718 150882 187954
rect 150326 187398 150562 187634
rect 150646 187398 150882 187634
rect 145826 147218 146062 147454
rect 146146 147218 146382 147454
rect 145826 146898 146062 147134
rect 146146 146898 146382 147134
rect 150326 151718 150562 151954
rect 150646 151718 150882 151954
rect 150326 151398 150562 151634
rect 150646 151398 150882 151634
rect 154826 192218 155062 192454
rect 155146 192218 155382 192454
rect 154826 191898 155062 192134
rect 155146 191898 155382 192134
rect 159326 196718 159562 196954
rect 159646 196718 159882 196954
rect 159326 196398 159562 196634
rect 159646 196398 159882 196634
rect 154826 156218 155062 156454
rect 155146 156218 155382 156454
rect 154826 155898 155062 156134
rect 155146 155898 155382 156134
rect 159326 160718 159562 160954
rect 159646 160718 159882 160954
rect 159326 160398 159562 160634
rect 159646 160398 159882 160634
rect 177326 178718 177562 178954
rect 177646 178718 177882 178954
rect 177326 178398 177562 178634
rect 177646 178398 177882 178634
rect 177326 142718 177562 142954
rect 177646 142718 177882 142954
rect 177326 142398 177562 142634
rect 177646 142398 177882 142634
rect 181826 183218 182062 183454
rect 182146 183218 182382 183454
rect 181826 182898 182062 183134
rect 182146 182898 182382 183134
rect 181826 147218 182062 147454
rect 182146 147218 182382 147454
rect 181826 146898 182062 147134
rect 182146 146898 182382 147134
rect 186326 187718 186562 187954
rect 186646 187718 186882 187954
rect 186326 187398 186562 187634
rect 186646 187398 186882 187634
rect 186326 151718 186562 151954
rect 186646 151718 186882 151954
rect 186326 151398 186562 151634
rect 186646 151398 186882 151634
rect 139610 115718 139846 115954
rect 139610 115398 139846 115634
rect 170330 115718 170566 115954
rect 170330 115398 170566 115634
rect 124250 111218 124486 111454
rect 124250 110898 124486 111134
rect 154970 111218 155206 111454
rect 154970 110898 155206 111134
rect 185690 111218 185926 111454
rect 185690 110898 185926 111134
rect 118826 48218 119062 48454
rect 119146 48218 119382 48454
rect 118826 47898 119062 48134
rect 119146 47898 119382 48134
rect 118826 12218 119062 12454
rect 119146 12218 119382 12454
rect 118826 11898 119062 12134
rect 119146 11898 119382 12134
rect 118826 -2502 119062 -2266
rect 119146 -2502 119382 -2266
rect 118826 -2822 119062 -2586
rect 119146 -2822 119382 -2586
rect 123326 52718 123562 52954
rect 123646 52718 123882 52954
rect 123326 52398 123562 52634
rect 123646 52398 123882 52634
rect 123326 16718 123562 16954
rect 123646 16718 123882 16954
rect 123326 16398 123562 16634
rect 123646 16398 123882 16634
rect 123326 -3462 123562 -3226
rect 123646 -3462 123882 -3226
rect 123326 -3782 123562 -3546
rect 123646 -3782 123882 -3546
rect 127826 57218 128062 57454
rect 128146 57218 128382 57454
rect 127826 56898 128062 57134
rect 128146 56898 128382 57134
rect 127826 21218 128062 21454
rect 128146 21218 128382 21454
rect 127826 20898 128062 21134
rect 128146 20898 128382 21134
rect 127826 -4422 128062 -4186
rect 128146 -4422 128382 -4186
rect 127826 -4742 128062 -4506
rect 128146 -4742 128382 -4506
rect 141326 70718 141562 70954
rect 141646 70718 141882 70954
rect 141326 70398 141562 70634
rect 141646 70398 141882 70634
rect 136826 66218 137062 66454
rect 137146 66218 137382 66454
rect 136826 65898 137062 66134
rect 137146 65898 137382 66134
rect 132326 61718 132562 61954
rect 132646 61718 132882 61954
rect 132326 61398 132562 61634
rect 132646 61398 132882 61634
rect 132326 25718 132562 25954
rect 132646 25718 132882 25954
rect 132326 25398 132562 25634
rect 132646 25398 132882 25634
rect 132326 -5382 132562 -5146
rect 132646 -5382 132882 -5146
rect 132326 -5702 132562 -5466
rect 132646 -5702 132882 -5466
rect 136826 30218 137062 30454
rect 137146 30218 137382 30454
rect 136826 29898 137062 30134
rect 137146 29898 137382 30134
rect 136826 -6342 137062 -6106
rect 137146 -6342 137382 -6106
rect 136826 -6662 137062 -6426
rect 137146 -6662 137382 -6426
rect 145826 75218 146062 75454
rect 146146 75218 146382 75454
rect 145826 74898 146062 75134
rect 146146 74898 146382 75134
rect 141326 34718 141562 34954
rect 141646 34718 141882 34954
rect 141326 34398 141562 34634
rect 141646 34398 141882 34634
rect 141326 -7302 141562 -7066
rect 141646 -7302 141882 -7066
rect 141326 -7622 141562 -7386
rect 141646 -7622 141882 -7386
rect 145826 39218 146062 39454
rect 146146 39218 146382 39454
rect 145826 38898 146062 39134
rect 146146 38898 146382 39134
rect 145826 3218 146062 3454
rect 146146 3218 146382 3454
rect 145826 2898 146062 3134
rect 146146 2898 146382 3134
rect 145826 -582 146062 -346
rect 146146 -582 146382 -346
rect 145826 -902 146062 -666
rect 146146 -902 146382 -666
rect 150326 43718 150562 43954
rect 150646 43718 150882 43954
rect 150326 43398 150562 43634
rect 150646 43398 150882 43634
rect 150326 7718 150562 7954
rect 150646 7718 150882 7954
rect 150326 7398 150562 7634
rect 150646 7398 150882 7634
rect 150326 -1542 150562 -1306
rect 150646 -1542 150882 -1306
rect 150326 -1862 150562 -1626
rect 150646 -1862 150882 -1626
rect 154826 48218 155062 48454
rect 155146 48218 155382 48454
rect 154826 47898 155062 48134
rect 155146 47898 155382 48134
rect 154826 12218 155062 12454
rect 155146 12218 155382 12454
rect 154826 11898 155062 12134
rect 155146 11898 155382 12134
rect 154826 -2502 155062 -2266
rect 155146 -2502 155382 -2266
rect 154826 -2822 155062 -2586
rect 155146 -2822 155382 -2586
rect 159326 52718 159562 52954
rect 159646 52718 159882 52954
rect 159326 52398 159562 52634
rect 159646 52398 159882 52634
rect 159326 16718 159562 16954
rect 159646 16718 159882 16954
rect 159326 16398 159562 16634
rect 159646 16398 159882 16634
rect 159326 -3462 159562 -3226
rect 159646 -3462 159882 -3226
rect 159326 -3782 159562 -3546
rect 159646 -3782 159882 -3546
rect 163826 57218 164062 57454
rect 164146 57218 164382 57454
rect 163826 56898 164062 57134
rect 164146 56898 164382 57134
rect 163826 21218 164062 21454
rect 164146 21218 164382 21454
rect 163826 20898 164062 21134
rect 164146 20898 164382 21134
rect 163826 -4422 164062 -4186
rect 164146 -4422 164382 -4186
rect 163826 -4742 164062 -4506
rect 164146 -4742 164382 -4506
rect 172826 66218 173062 66454
rect 173146 66218 173382 66454
rect 172826 65898 173062 66134
rect 173146 65898 173382 66134
rect 168326 61718 168562 61954
rect 168646 61718 168882 61954
rect 168326 61398 168562 61634
rect 168646 61398 168882 61634
rect 168326 25718 168562 25954
rect 168646 25718 168882 25954
rect 168326 25398 168562 25634
rect 168646 25398 168882 25634
rect 168326 -5382 168562 -5146
rect 168646 -5382 168882 -5146
rect 168326 -5702 168562 -5466
rect 168646 -5702 168882 -5466
rect 177326 70718 177562 70954
rect 177646 70718 177882 70954
rect 177326 70398 177562 70634
rect 177646 70398 177882 70634
rect 172826 30218 173062 30454
rect 173146 30218 173382 30454
rect 172826 29898 173062 30134
rect 173146 29898 173382 30134
rect 172826 -6342 173062 -6106
rect 173146 -6342 173382 -6106
rect 172826 -6662 173062 -6426
rect 173146 -6662 173382 -6426
rect 177326 34718 177562 34954
rect 177646 34718 177882 34954
rect 177326 34398 177562 34634
rect 177646 34398 177882 34634
rect 177326 -7302 177562 -7066
rect 177646 -7302 177882 -7066
rect 177326 -7622 177562 -7386
rect 177646 -7622 177882 -7386
rect 181826 75218 182062 75454
rect 182146 75218 182382 75454
rect 181826 74898 182062 75134
rect 182146 74898 182382 75134
rect 181826 39218 182062 39454
rect 182146 39218 182382 39454
rect 181826 38898 182062 39134
rect 182146 38898 182382 39134
rect 181826 3218 182062 3454
rect 182146 3218 182382 3454
rect 181826 2898 182062 3134
rect 182146 2898 182382 3134
rect 181826 -582 182062 -346
rect 182146 -582 182382 -346
rect 181826 -902 182062 -666
rect 182146 -902 182382 -666
rect 190826 192218 191062 192454
rect 191146 192218 191382 192454
rect 190826 191898 191062 192134
rect 191146 191898 191382 192134
rect 190826 156218 191062 156454
rect 191146 156218 191382 156454
rect 190826 155898 191062 156134
rect 191146 155898 191382 156134
rect 195326 232718 195562 232954
rect 195646 232718 195882 232954
rect 195326 232398 195562 232634
rect 195646 232398 195882 232634
rect 195326 196718 195562 196954
rect 195646 196718 195882 196954
rect 195326 196398 195562 196634
rect 195646 196398 195882 196634
rect 199826 708442 200062 708678
rect 200146 708442 200382 708678
rect 199826 708122 200062 708358
rect 200146 708122 200382 708358
rect 199826 669218 200062 669454
rect 200146 669218 200382 669454
rect 199826 668898 200062 669134
rect 200146 668898 200382 669134
rect 199826 633218 200062 633454
rect 200146 633218 200382 633454
rect 199826 632898 200062 633134
rect 200146 632898 200382 633134
rect 199826 597218 200062 597454
rect 200146 597218 200382 597454
rect 199826 596898 200062 597134
rect 200146 596898 200382 597134
rect 199826 561218 200062 561454
rect 200146 561218 200382 561454
rect 199826 560898 200062 561134
rect 200146 560898 200382 561134
rect 199826 525218 200062 525454
rect 200146 525218 200382 525454
rect 199826 524898 200062 525134
rect 200146 524898 200382 525134
rect 199826 489218 200062 489454
rect 200146 489218 200382 489454
rect 199826 488898 200062 489134
rect 200146 488898 200382 489134
rect 199826 453218 200062 453454
rect 200146 453218 200382 453454
rect 199826 452898 200062 453134
rect 200146 452898 200382 453134
rect 199826 417218 200062 417454
rect 200146 417218 200382 417454
rect 199826 416898 200062 417134
rect 200146 416898 200382 417134
rect 199826 381218 200062 381454
rect 200146 381218 200382 381454
rect 199826 380898 200062 381134
rect 200146 380898 200382 381134
rect 199826 345218 200062 345454
rect 200146 345218 200382 345454
rect 199826 344898 200062 345134
rect 200146 344898 200382 345134
rect 199826 309218 200062 309454
rect 200146 309218 200382 309454
rect 199826 308898 200062 309134
rect 200146 308898 200382 309134
rect 199826 273218 200062 273454
rect 200146 273218 200382 273454
rect 199826 272898 200062 273134
rect 200146 272898 200382 273134
rect 199826 237218 200062 237454
rect 200146 237218 200382 237454
rect 199826 236898 200062 237134
rect 200146 236898 200382 237134
rect 199826 201218 200062 201454
rect 200146 201218 200382 201454
rect 199826 200898 200062 201134
rect 200146 200898 200382 201134
rect 186326 43718 186562 43954
rect 186646 43718 186882 43954
rect 186326 43398 186562 43634
rect 186646 43398 186882 43634
rect 186326 7718 186562 7954
rect 186646 7718 186882 7954
rect 186326 7398 186562 7634
rect 186646 7398 186882 7634
rect 186326 -1542 186562 -1306
rect 186646 -1542 186882 -1306
rect 186326 -1862 186562 -1626
rect 186646 -1862 186882 -1626
rect 195326 160718 195562 160954
rect 195646 160718 195882 160954
rect 195326 160398 195562 160634
rect 195646 160398 195882 160634
rect 195326 124718 195562 124954
rect 195646 124718 195882 124954
rect 195326 124398 195562 124634
rect 195646 124398 195882 124634
rect 195326 88718 195562 88954
rect 195646 88718 195882 88954
rect 195326 88398 195562 88634
rect 195646 88398 195882 88634
rect 190826 48218 191062 48454
rect 191146 48218 191382 48454
rect 190826 47898 191062 48134
rect 191146 47898 191382 48134
rect 204326 709402 204562 709638
rect 204646 709402 204882 709638
rect 204326 709082 204562 709318
rect 204646 709082 204882 709318
rect 204326 673718 204562 673954
rect 204646 673718 204882 673954
rect 204326 673398 204562 673634
rect 204646 673398 204882 673634
rect 204326 637718 204562 637954
rect 204646 637718 204882 637954
rect 204326 637398 204562 637634
rect 204646 637398 204882 637634
rect 204326 601718 204562 601954
rect 204646 601718 204882 601954
rect 204326 601398 204562 601634
rect 204646 601398 204882 601634
rect 204326 565718 204562 565954
rect 204646 565718 204882 565954
rect 204326 565398 204562 565634
rect 204646 565398 204882 565634
rect 204326 529718 204562 529954
rect 204646 529718 204882 529954
rect 204326 529398 204562 529634
rect 204646 529398 204882 529634
rect 204326 493718 204562 493954
rect 204646 493718 204882 493954
rect 204326 493398 204562 493634
rect 204646 493398 204882 493634
rect 204326 457718 204562 457954
rect 204646 457718 204882 457954
rect 204326 457398 204562 457634
rect 204646 457398 204882 457634
rect 204326 421718 204562 421954
rect 204646 421718 204882 421954
rect 204326 421398 204562 421634
rect 204646 421398 204882 421634
rect 204326 385718 204562 385954
rect 204646 385718 204882 385954
rect 204326 385398 204562 385634
rect 204646 385398 204882 385634
rect 204326 349718 204562 349954
rect 204646 349718 204882 349954
rect 204326 349398 204562 349634
rect 204646 349398 204882 349634
rect 204326 313718 204562 313954
rect 204646 313718 204882 313954
rect 204326 313398 204562 313634
rect 204646 313398 204882 313634
rect 204326 277718 204562 277954
rect 204646 277718 204882 277954
rect 204326 277398 204562 277634
rect 204646 277398 204882 277634
rect 204326 241718 204562 241954
rect 204646 241718 204882 241954
rect 204326 241398 204562 241634
rect 204646 241398 204882 241634
rect 204326 205718 204562 205954
rect 204646 205718 204882 205954
rect 204326 205398 204562 205634
rect 204646 205398 204882 205634
rect 199826 165218 200062 165454
rect 200146 165218 200382 165454
rect 199826 164898 200062 165134
rect 200146 164898 200382 165134
rect 199826 129218 200062 129454
rect 200146 129218 200382 129454
rect 199826 128898 200062 129134
rect 200146 128898 200382 129134
rect 199826 93218 200062 93454
rect 200146 93218 200382 93454
rect 199826 92898 200062 93134
rect 200146 92898 200382 93134
rect 195326 52718 195562 52954
rect 195646 52718 195882 52954
rect 195326 52398 195562 52634
rect 195646 52398 195882 52634
rect 190826 12218 191062 12454
rect 191146 12218 191382 12454
rect 190826 11898 191062 12134
rect 191146 11898 191382 12134
rect 190826 -2502 191062 -2266
rect 191146 -2502 191382 -2266
rect 190826 -2822 191062 -2586
rect 191146 -2822 191382 -2586
rect 195326 16718 195562 16954
rect 195646 16718 195882 16954
rect 195326 16398 195562 16634
rect 195646 16398 195882 16634
rect 195326 -3462 195562 -3226
rect 195646 -3462 195882 -3226
rect 195326 -3782 195562 -3546
rect 195646 -3782 195882 -3546
rect 208826 710362 209062 710598
rect 209146 710362 209382 710598
rect 208826 710042 209062 710278
rect 209146 710042 209382 710278
rect 208826 678218 209062 678454
rect 209146 678218 209382 678454
rect 208826 677898 209062 678134
rect 209146 677898 209382 678134
rect 208826 642218 209062 642454
rect 209146 642218 209382 642454
rect 208826 641898 209062 642134
rect 209146 641898 209382 642134
rect 208826 606218 209062 606454
rect 209146 606218 209382 606454
rect 208826 605898 209062 606134
rect 209146 605898 209382 606134
rect 208826 570218 209062 570454
rect 209146 570218 209382 570454
rect 208826 569898 209062 570134
rect 209146 569898 209382 570134
rect 208826 534218 209062 534454
rect 209146 534218 209382 534454
rect 208826 533898 209062 534134
rect 209146 533898 209382 534134
rect 208826 498218 209062 498454
rect 209146 498218 209382 498454
rect 208826 497898 209062 498134
rect 209146 497898 209382 498134
rect 208826 462218 209062 462454
rect 209146 462218 209382 462454
rect 208826 461898 209062 462134
rect 209146 461898 209382 462134
rect 208826 426218 209062 426454
rect 209146 426218 209382 426454
rect 208826 425898 209062 426134
rect 209146 425898 209382 426134
rect 208826 390218 209062 390454
rect 209146 390218 209382 390454
rect 208826 389898 209062 390134
rect 209146 389898 209382 390134
rect 208826 354218 209062 354454
rect 209146 354218 209382 354454
rect 208826 353898 209062 354134
rect 209146 353898 209382 354134
rect 208826 318218 209062 318454
rect 209146 318218 209382 318454
rect 208826 317898 209062 318134
rect 209146 317898 209382 318134
rect 208826 282218 209062 282454
rect 209146 282218 209382 282454
rect 208826 281898 209062 282134
rect 209146 281898 209382 282134
rect 208826 246218 209062 246454
rect 209146 246218 209382 246454
rect 208826 245898 209062 246134
rect 209146 245898 209382 246134
rect 208826 210218 209062 210454
rect 209146 210218 209382 210454
rect 208826 209898 209062 210134
rect 209146 209898 209382 210134
rect 204326 169718 204562 169954
rect 204646 169718 204882 169954
rect 204326 169398 204562 169634
rect 204646 169398 204882 169634
rect 204326 133718 204562 133954
rect 204646 133718 204882 133954
rect 204326 133398 204562 133634
rect 204646 133398 204882 133634
rect 204326 97718 204562 97954
rect 204646 97718 204882 97954
rect 204326 97398 204562 97634
rect 204646 97398 204882 97634
rect 199826 57218 200062 57454
rect 200146 57218 200382 57454
rect 199826 56898 200062 57134
rect 200146 56898 200382 57134
rect 199826 21218 200062 21454
rect 200146 21218 200382 21454
rect 199826 20898 200062 21134
rect 200146 20898 200382 21134
rect 199826 -4422 200062 -4186
rect 200146 -4422 200382 -4186
rect 199826 -4742 200062 -4506
rect 200146 -4742 200382 -4506
rect 213326 711322 213562 711558
rect 213646 711322 213882 711558
rect 213326 711002 213562 711238
rect 213646 711002 213882 711238
rect 213326 682718 213562 682954
rect 213646 682718 213882 682954
rect 213326 682398 213562 682634
rect 213646 682398 213882 682634
rect 213326 646718 213562 646954
rect 213646 646718 213882 646954
rect 213326 646398 213562 646634
rect 213646 646398 213882 646634
rect 213326 610718 213562 610954
rect 213646 610718 213882 610954
rect 213326 610398 213562 610634
rect 213646 610398 213882 610634
rect 213326 574718 213562 574954
rect 213646 574718 213882 574954
rect 213326 574398 213562 574634
rect 213646 574398 213882 574634
rect 213326 538718 213562 538954
rect 213646 538718 213882 538954
rect 213326 538398 213562 538634
rect 213646 538398 213882 538634
rect 213326 502718 213562 502954
rect 213646 502718 213882 502954
rect 213326 502398 213562 502634
rect 213646 502398 213882 502634
rect 213326 466718 213562 466954
rect 213646 466718 213882 466954
rect 213326 466398 213562 466634
rect 213646 466398 213882 466634
rect 213326 430718 213562 430954
rect 213646 430718 213882 430954
rect 213326 430398 213562 430634
rect 213646 430398 213882 430634
rect 213326 394718 213562 394954
rect 213646 394718 213882 394954
rect 213326 394398 213562 394634
rect 213646 394398 213882 394634
rect 213326 358718 213562 358954
rect 213646 358718 213882 358954
rect 213326 358398 213562 358634
rect 213646 358398 213882 358634
rect 213326 322718 213562 322954
rect 213646 322718 213882 322954
rect 213326 322398 213562 322634
rect 213646 322398 213882 322634
rect 213326 286718 213562 286954
rect 213646 286718 213882 286954
rect 213326 286398 213562 286634
rect 213646 286398 213882 286634
rect 213326 250718 213562 250954
rect 213646 250718 213882 250954
rect 213326 250398 213562 250634
rect 213646 250398 213882 250634
rect 213326 214718 213562 214954
rect 213646 214718 213882 214954
rect 213326 214398 213562 214634
rect 213646 214398 213882 214634
rect 208826 174218 209062 174454
rect 209146 174218 209382 174454
rect 208826 173898 209062 174134
rect 209146 173898 209382 174134
rect 208826 138218 209062 138454
rect 209146 138218 209382 138454
rect 208826 137898 209062 138134
rect 209146 137898 209382 138134
rect 208826 102218 209062 102454
rect 209146 102218 209382 102454
rect 208826 101898 209062 102134
rect 209146 101898 209382 102134
rect 204326 61718 204562 61954
rect 204646 61718 204882 61954
rect 204326 61398 204562 61634
rect 204646 61398 204882 61634
rect 204326 25718 204562 25954
rect 204646 25718 204882 25954
rect 204326 25398 204562 25634
rect 204646 25398 204882 25634
rect 204326 -5382 204562 -5146
rect 204646 -5382 204882 -5146
rect 204326 -5702 204562 -5466
rect 204646 -5702 204882 -5466
rect 213326 178718 213562 178954
rect 213646 178718 213882 178954
rect 213326 178398 213562 178634
rect 213646 178398 213882 178634
rect 213326 142718 213562 142954
rect 213646 142718 213882 142954
rect 213326 142398 213562 142634
rect 213646 142398 213882 142634
rect 213326 106718 213562 106954
rect 213646 106718 213882 106954
rect 213326 106398 213562 106634
rect 213646 106398 213882 106634
rect 208826 66218 209062 66454
rect 209146 66218 209382 66454
rect 208826 65898 209062 66134
rect 209146 65898 209382 66134
rect 208826 30218 209062 30454
rect 209146 30218 209382 30454
rect 208826 29898 209062 30134
rect 209146 29898 209382 30134
rect 208826 -6342 209062 -6106
rect 209146 -6342 209382 -6106
rect 208826 -6662 209062 -6426
rect 209146 -6662 209382 -6426
rect 213326 70718 213562 70954
rect 213646 70718 213882 70954
rect 213326 70398 213562 70634
rect 213646 70398 213882 70634
rect 213326 34718 213562 34954
rect 213646 34718 213882 34954
rect 213326 34398 213562 34634
rect 213646 34398 213882 34634
rect 213326 -7302 213562 -7066
rect 213646 -7302 213882 -7066
rect 213326 -7622 213562 -7386
rect 213646 -7622 213882 -7386
rect 217826 704602 218062 704838
rect 218146 704602 218382 704838
rect 217826 704282 218062 704518
rect 218146 704282 218382 704518
rect 217826 687218 218062 687454
rect 218146 687218 218382 687454
rect 217826 686898 218062 687134
rect 218146 686898 218382 687134
rect 217826 651218 218062 651454
rect 218146 651218 218382 651454
rect 217826 650898 218062 651134
rect 218146 650898 218382 651134
rect 217826 615218 218062 615454
rect 218146 615218 218382 615454
rect 217826 614898 218062 615134
rect 218146 614898 218382 615134
rect 217826 579218 218062 579454
rect 218146 579218 218382 579454
rect 217826 578898 218062 579134
rect 218146 578898 218382 579134
rect 217826 543218 218062 543454
rect 218146 543218 218382 543454
rect 217826 542898 218062 543134
rect 218146 542898 218382 543134
rect 217826 507218 218062 507454
rect 218146 507218 218382 507454
rect 217826 506898 218062 507134
rect 218146 506898 218382 507134
rect 217826 471218 218062 471454
rect 218146 471218 218382 471454
rect 217826 470898 218062 471134
rect 218146 470898 218382 471134
rect 217826 435218 218062 435454
rect 218146 435218 218382 435454
rect 217826 434898 218062 435134
rect 218146 434898 218382 435134
rect 217826 399218 218062 399454
rect 218146 399218 218382 399454
rect 217826 398898 218062 399134
rect 218146 398898 218382 399134
rect 217826 363218 218062 363454
rect 218146 363218 218382 363454
rect 217826 362898 218062 363134
rect 218146 362898 218382 363134
rect 217826 327218 218062 327454
rect 218146 327218 218382 327454
rect 217826 326898 218062 327134
rect 218146 326898 218382 327134
rect 217826 291218 218062 291454
rect 218146 291218 218382 291454
rect 217826 290898 218062 291134
rect 218146 290898 218382 291134
rect 217826 255218 218062 255454
rect 218146 255218 218382 255454
rect 217826 254898 218062 255134
rect 218146 254898 218382 255134
rect 217826 219218 218062 219454
rect 218146 219218 218382 219454
rect 217826 218898 218062 219134
rect 218146 218898 218382 219134
rect 217826 183218 218062 183454
rect 218146 183218 218382 183454
rect 217826 182898 218062 183134
rect 218146 182898 218382 183134
rect 217826 147218 218062 147454
rect 218146 147218 218382 147454
rect 217826 146898 218062 147134
rect 218146 146898 218382 147134
rect 217826 111218 218062 111454
rect 218146 111218 218382 111454
rect 217826 110898 218062 111134
rect 218146 110898 218382 111134
rect 217826 75218 218062 75454
rect 218146 75218 218382 75454
rect 217826 74898 218062 75134
rect 218146 74898 218382 75134
rect 217826 39218 218062 39454
rect 218146 39218 218382 39454
rect 217826 38898 218062 39134
rect 218146 38898 218382 39134
rect 217826 3218 218062 3454
rect 218146 3218 218382 3454
rect 217826 2898 218062 3134
rect 218146 2898 218382 3134
rect 217826 -582 218062 -346
rect 218146 -582 218382 -346
rect 217826 -902 218062 -666
rect 218146 -902 218382 -666
rect 222326 705562 222562 705798
rect 222646 705562 222882 705798
rect 222326 705242 222562 705478
rect 222646 705242 222882 705478
rect 222326 691718 222562 691954
rect 222646 691718 222882 691954
rect 222326 691398 222562 691634
rect 222646 691398 222882 691634
rect 222326 655718 222562 655954
rect 222646 655718 222882 655954
rect 222326 655398 222562 655634
rect 222646 655398 222882 655634
rect 222326 619718 222562 619954
rect 222646 619718 222882 619954
rect 222326 619398 222562 619634
rect 222646 619398 222882 619634
rect 222326 583718 222562 583954
rect 222646 583718 222882 583954
rect 222326 583398 222562 583634
rect 222646 583398 222882 583634
rect 222326 547718 222562 547954
rect 222646 547718 222882 547954
rect 222326 547398 222562 547634
rect 222646 547398 222882 547634
rect 222326 511718 222562 511954
rect 222646 511718 222882 511954
rect 222326 511398 222562 511634
rect 222646 511398 222882 511634
rect 222326 475718 222562 475954
rect 222646 475718 222882 475954
rect 222326 475398 222562 475634
rect 222646 475398 222882 475634
rect 222326 439718 222562 439954
rect 222646 439718 222882 439954
rect 222326 439398 222562 439634
rect 222646 439398 222882 439634
rect 222326 403718 222562 403954
rect 222646 403718 222882 403954
rect 222326 403398 222562 403634
rect 222646 403398 222882 403634
rect 222326 367718 222562 367954
rect 222646 367718 222882 367954
rect 222326 367398 222562 367634
rect 222646 367398 222882 367634
rect 222326 331718 222562 331954
rect 222646 331718 222882 331954
rect 222326 331398 222562 331634
rect 222646 331398 222882 331634
rect 222326 295718 222562 295954
rect 222646 295718 222882 295954
rect 222326 295398 222562 295634
rect 222646 295398 222882 295634
rect 222326 259718 222562 259954
rect 222646 259718 222882 259954
rect 222326 259398 222562 259634
rect 222646 259398 222882 259634
rect 222326 223718 222562 223954
rect 222646 223718 222882 223954
rect 222326 223398 222562 223634
rect 222646 223398 222882 223634
rect 222326 187718 222562 187954
rect 222646 187718 222882 187954
rect 222326 187398 222562 187634
rect 222646 187398 222882 187634
rect 222326 151718 222562 151954
rect 222646 151718 222882 151954
rect 222326 151398 222562 151634
rect 222646 151398 222882 151634
rect 222326 115718 222562 115954
rect 222646 115718 222882 115954
rect 222326 115398 222562 115634
rect 222646 115398 222882 115634
rect 222326 79718 222562 79954
rect 222646 79718 222882 79954
rect 222326 79398 222562 79634
rect 222646 79398 222882 79634
rect 222326 43718 222562 43954
rect 222646 43718 222882 43954
rect 222326 43398 222562 43634
rect 222646 43398 222882 43634
rect 222326 7718 222562 7954
rect 222646 7718 222882 7954
rect 222326 7398 222562 7634
rect 222646 7398 222882 7634
rect 222326 -1542 222562 -1306
rect 222646 -1542 222882 -1306
rect 222326 -1862 222562 -1626
rect 222646 -1862 222882 -1626
rect 226826 706522 227062 706758
rect 227146 706522 227382 706758
rect 226826 706202 227062 706438
rect 227146 706202 227382 706438
rect 226826 696218 227062 696454
rect 227146 696218 227382 696454
rect 226826 695898 227062 696134
rect 227146 695898 227382 696134
rect 226826 660218 227062 660454
rect 227146 660218 227382 660454
rect 226826 659898 227062 660134
rect 227146 659898 227382 660134
rect 226826 624218 227062 624454
rect 227146 624218 227382 624454
rect 226826 623898 227062 624134
rect 227146 623898 227382 624134
rect 226826 588218 227062 588454
rect 227146 588218 227382 588454
rect 226826 587898 227062 588134
rect 227146 587898 227382 588134
rect 226826 552218 227062 552454
rect 227146 552218 227382 552454
rect 226826 551898 227062 552134
rect 227146 551898 227382 552134
rect 226826 516218 227062 516454
rect 227146 516218 227382 516454
rect 226826 515898 227062 516134
rect 227146 515898 227382 516134
rect 226826 480218 227062 480454
rect 227146 480218 227382 480454
rect 226826 479898 227062 480134
rect 227146 479898 227382 480134
rect 226826 444218 227062 444454
rect 227146 444218 227382 444454
rect 226826 443898 227062 444134
rect 227146 443898 227382 444134
rect 226826 408218 227062 408454
rect 227146 408218 227382 408454
rect 226826 407898 227062 408134
rect 227146 407898 227382 408134
rect 226826 372218 227062 372454
rect 227146 372218 227382 372454
rect 226826 371898 227062 372134
rect 227146 371898 227382 372134
rect 226826 336218 227062 336454
rect 227146 336218 227382 336454
rect 226826 335898 227062 336134
rect 227146 335898 227382 336134
rect 226826 300218 227062 300454
rect 227146 300218 227382 300454
rect 226826 299898 227062 300134
rect 227146 299898 227382 300134
rect 226826 264218 227062 264454
rect 227146 264218 227382 264454
rect 226826 263898 227062 264134
rect 227146 263898 227382 264134
rect 226826 228218 227062 228454
rect 227146 228218 227382 228454
rect 226826 227898 227062 228134
rect 227146 227898 227382 228134
rect 226826 192218 227062 192454
rect 227146 192218 227382 192454
rect 226826 191898 227062 192134
rect 227146 191898 227382 192134
rect 226826 156218 227062 156454
rect 227146 156218 227382 156454
rect 226826 155898 227062 156134
rect 227146 155898 227382 156134
rect 226826 120218 227062 120454
rect 227146 120218 227382 120454
rect 226826 119898 227062 120134
rect 227146 119898 227382 120134
rect 226826 84218 227062 84454
rect 227146 84218 227382 84454
rect 226826 83898 227062 84134
rect 227146 83898 227382 84134
rect 226826 48218 227062 48454
rect 227146 48218 227382 48454
rect 226826 47898 227062 48134
rect 227146 47898 227382 48134
rect 226826 12218 227062 12454
rect 227146 12218 227382 12454
rect 226826 11898 227062 12134
rect 227146 11898 227382 12134
rect 226826 -2502 227062 -2266
rect 227146 -2502 227382 -2266
rect 226826 -2822 227062 -2586
rect 227146 -2822 227382 -2586
rect 231326 707482 231562 707718
rect 231646 707482 231882 707718
rect 231326 707162 231562 707398
rect 231646 707162 231882 707398
rect 231326 700718 231562 700954
rect 231646 700718 231882 700954
rect 231326 700398 231562 700634
rect 231646 700398 231882 700634
rect 231326 664718 231562 664954
rect 231646 664718 231882 664954
rect 231326 664398 231562 664634
rect 231646 664398 231882 664634
rect 231326 628718 231562 628954
rect 231646 628718 231882 628954
rect 231326 628398 231562 628634
rect 231646 628398 231882 628634
rect 231326 592718 231562 592954
rect 231646 592718 231882 592954
rect 231326 592398 231562 592634
rect 231646 592398 231882 592634
rect 231326 556718 231562 556954
rect 231646 556718 231882 556954
rect 231326 556398 231562 556634
rect 231646 556398 231882 556634
rect 231326 520718 231562 520954
rect 231646 520718 231882 520954
rect 231326 520398 231562 520634
rect 231646 520398 231882 520634
rect 231326 484718 231562 484954
rect 231646 484718 231882 484954
rect 231326 484398 231562 484634
rect 231646 484398 231882 484634
rect 231326 448718 231562 448954
rect 231646 448718 231882 448954
rect 231326 448398 231562 448634
rect 231646 448398 231882 448634
rect 231326 412718 231562 412954
rect 231646 412718 231882 412954
rect 231326 412398 231562 412634
rect 231646 412398 231882 412634
rect 231326 376718 231562 376954
rect 231646 376718 231882 376954
rect 231326 376398 231562 376634
rect 231646 376398 231882 376634
rect 231326 340718 231562 340954
rect 231646 340718 231882 340954
rect 231326 340398 231562 340634
rect 231646 340398 231882 340634
rect 231326 304718 231562 304954
rect 231646 304718 231882 304954
rect 231326 304398 231562 304634
rect 231646 304398 231882 304634
rect 231326 268718 231562 268954
rect 231646 268718 231882 268954
rect 231326 268398 231562 268634
rect 231646 268398 231882 268634
rect 231326 232718 231562 232954
rect 231646 232718 231882 232954
rect 231326 232398 231562 232634
rect 231646 232398 231882 232634
rect 231326 196718 231562 196954
rect 231646 196718 231882 196954
rect 231326 196398 231562 196634
rect 231646 196398 231882 196634
rect 231326 160718 231562 160954
rect 231646 160718 231882 160954
rect 231326 160398 231562 160634
rect 231646 160398 231882 160634
rect 231326 124718 231562 124954
rect 231646 124718 231882 124954
rect 231326 124398 231562 124634
rect 231646 124398 231882 124634
rect 231326 88718 231562 88954
rect 231646 88718 231882 88954
rect 231326 88398 231562 88634
rect 231646 88398 231882 88634
rect 231326 52718 231562 52954
rect 231646 52718 231882 52954
rect 231326 52398 231562 52634
rect 231646 52398 231882 52634
rect 231326 16718 231562 16954
rect 231646 16718 231882 16954
rect 231326 16398 231562 16634
rect 231646 16398 231882 16634
rect 231326 -3462 231562 -3226
rect 231646 -3462 231882 -3226
rect 231326 -3782 231562 -3546
rect 231646 -3782 231882 -3546
rect 235826 708442 236062 708678
rect 236146 708442 236382 708678
rect 235826 708122 236062 708358
rect 236146 708122 236382 708358
rect 235826 669218 236062 669454
rect 236146 669218 236382 669454
rect 235826 668898 236062 669134
rect 236146 668898 236382 669134
rect 235826 633218 236062 633454
rect 236146 633218 236382 633454
rect 235826 632898 236062 633134
rect 236146 632898 236382 633134
rect 235826 597218 236062 597454
rect 236146 597218 236382 597454
rect 235826 596898 236062 597134
rect 236146 596898 236382 597134
rect 235826 561218 236062 561454
rect 236146 561218 236382 561454
rect 235826 560898 236062 561134
rect 236146 560898 236382 561134
rect 235826 525218 236062 525454
rect 236146 525218 236382 525454
rect 235826 524898 236062 525134
rect 236146 524898 236382 525134
rect 235826 489218 236062 489454
rect 236146 489218 236382 489454
rect 235826 488898 236062 489134
rect 236146 488898 236382 489134
rect 235826 453218 236062 453454
rect 236146 453218 236382 453454
rect 235826 452898 236062 453134
rect 236146 452898 236382 453134
rect 235826 417218 236062 417454
rect 236146 417218 236382 417454
rect 235826 416898 236062 417134
rect 236146 416898 236382 417134
rect 235826 381218 236062 381454
rect 236146 381218 236382 381454
rect 235826 380898 236062 381134
rect 236146 380898 236382 381134
rect 235826 345218 236062 345454
rect 236146 345218 236382 345454
rect 235826 344898 236062 345134
rect 236146 344898 236382 345134
rect 235826 309218 236062 309454
rect 236146 309218 236382 309454
rect 235826 308898 236062 309134
rect 236146 308898 236382 309134
rect 235826 273218 236062 273454
rect 236146 273218 236382 273454
rect 235826 272898 236062 273134
rect 236146 272898 236382 273134
rect 235826 237218 236062 237454
rect 236146 237218 236382 237454
rect 235826 236898 236062 237134
rect 236146 236898 236382 237134
rect 235826 201218 236062 201454
rect 236146 201218 236382 201454
rect 235826 200898 236062 201134
rect 236146 200898 236382 201134
rect 235826 165218 236062 165454
rect 236146 165218 236382 165454
rect 235826 164898 236062 165134
rect 236146 164898 236382 165134
rect 235826 129218 236062 129454
rect 236146 129218 236382 129454
rect 235826 128898 236062 129134
rect 236146 128898 236382 129134
rect 235826 93218 236062 93454
rect 236146 93218 236382 93454
rect 235826 92898 236062 93134
rect 236146 92898 236382 93134
rect 235826 57218 236062 57454
rect 236146 57218 236382 57454
rect 235826 56898 236062 57134
rect 236146 56898 236382 57134
rect 235826 21218 236062 21454
rect 236146 21218 236382 21454
rect 235826 20898 236062 21134
rect 236146 20898 236382 21134
rect 235826 -4422 236062 -4186
rect 236146 -4422 236382 -4186
rect 235826 -4742 236062 -4506
rect 236146 -4742 236382 -4506
rect 240326 709402 240562 709638
rect 240646 709402 240882 709638
rect 240326 709082 240562 709318
rect 240646 709082 240882 709318
rect 240326 673718 240562 673954
rect 240646 673718 240882 673954
rect 240326 673398 240562 673634
rect 240646 673398 240882 673634
rect 240326 637718 240562 637954
rect 240646 637718 240882 637954
rect 240326 637398 240562 637634
rect 240646 637398 240882 637634
rect 240326 601718 240562 601954
rect 240646 601718 240882 601954
rect 240326 601398 240562 601634
rect 240646 601398 240882 601634
rect 240326 565718 240562 565954
rect 240646 565718 240882 565954
rect 240326 565398 240562 565634
rect 240646 565398 240882 565634
rect 240326 529718 240562 529954
rect 240646 529718 240882 529954
rect 240326 529398 240562 529634
rect 240646 529398 240882 529634
rect 240326 493718 240562 493954
rect 240646 493718 240882 493954
rect 240326 493398 240562 493634
rect 240646 493398 240882 493634
rect 240326 457718 240562 457954
rect 240646 457718 240882 457954
rect 240326 457398 240562 457634
rect 240646 457398 240882 457634
rect 240326 421718 240562 421954
rect 240646 421718 240882 421954
rect 240326 421398 240562 421634
rect 240646 421398 240882 421634
rect 240326 385718 240562 385954
rect 240646 385718 240882 385954
rect 240326 385398 240562 385634
rect 240646 385398 240882 385634
rect 240326 349718 240562 349954
rect 240646 349718 240882 349954
rect 240326 349398 240562 349634
rect 240646 349398 240882 349634
rect 240326 313718 240562 313954
rect 240646 313718 240882 313954
rect 240326 313398 240562 313634
rect 240646 313398 240882 313634
rect 240326 277718 240562 277954
rect 240646 277718 240882 277954
rect 240326 277398 240562 277634
rect 240646 277398 240882 277634
rect 240326 241718 240562 241954
rect 240646 241718 240882 241954
rect 240326 241398 240562 241634
rect 240646 241398 240882 241634
rect 240326 205718 240562 205954
rect 240646 205718 240882 205954
rect 240326 205398 240562 205634
rect 240646 205398 240882 205634
rect 240326 169718 240562 169954
rect 240646 169718 240882 169954
rect 240326 169398 240562 169634
rect 240646 169398 240882 169634
rect 240326 133718 240562 133954
rect 240646 133718 240882 133954
rect 240326 133398 240562 133634
rect 240646 133398 240882 133634
rect 240326 97718 240562 97954
rect 240646 97718 240882 97954
rect 240326 97398 240562 97634
rect 240646 97398 240882 97634
rect 240326 61718 240562 61954
rect 240646 61718 240882 61954
rect 240326 61398 240562 61634
rect 240646 61398 240882 61634
rect 240326 25718 240562 25954
rect 240646 25718 240882 25954
rect 240326 25398 240562 25634
rect 240646 25398 240882 25634
rect 240326 -5382 240562 -5146
rect 240646 -5382 240882 -5146
rect 240326 -5702 240562 -5466
rect 240646 -5702 240882 -5466
rect 244826 710362 245062 710598
rect 245146 710362 245382 710598
rect 244826 710042 245062 710278
rect 245146 710042 245382 710278
rect 244826 678218 245062 678454
rect 245146 678218 245382 678454
rect 244826 677898 245062 678134
rect 245146 677898 245382 678134
rect 244826 642218 245062 642454
rect 245146 642218 245382 642454
rect 244826 641898 245062 642134
rect 245146 641898 245382 642134
rect 244826 606218 245062 606454
rect 245146 606218 245382 606454
rect 244826 605898 245062 606134
rect 245146 605898 245382 606134
rect 244826 570218 245062 570454
rect 245146 570218 245382 570454
rect 244826 569898 245062 570134
rect 245146 569898 245382 570134
rect 244826 534218 245062 534454
rect 245146 534218 245382 534454
rect 244826 533898 245062 534134
rect 245146 533898 245382 534134
rect 244826 498218 245062 498454
rect 245146 498218 245382 498454
rect 244826 497898 245062 498134
rect 245146 497898 245382 498134
rect 244826 462218 245062 462454
rect 245146 462218 245382 462454
rect 244826 461898 245062 462134
rect 245146 461898 245382 462134
rect 244826 426218 245062 426454
rect 245146 426218 245382 426454
rect 244826 425898 245062 426134
rect 245146 425898 245382 426134
rect 244826 390218 245062 390454
rect 245146 390218 245382 390454
rect 244826 389898 245062 390134
rect 245146 389898 245382 390134
rect 244826 354218 245062 354454
rect 245146 354218 245382 354454
rect 244826 353898 245062 354134
rect 245146 353898 245382 354134
rect 244826 318218 245062 318454
rect 245146 318218 245382 318454
rect 244826 317898 245062 318134
rect 245146 317898 245382 318134
rect 244826 282218 245062 282454
rect 245146 282218 245382 282454
rect 244826 281898 245062 282134
rect 245146 281898 245382 282134
rect 244826 246218 245062 246454
rect 245146 246218 245382 246454
rect 244826 245898 245062 246134
rect 245146 245898 245382 246134
rect 244826 210218 245062 210454
rect 245146 210218 245382 210454
rect 244826 209898 245062 210134
rect 245146 209898 245382 210134
rect 244826 174218 245062 174454
rect 245146 174218 245382 174454
rect 244826 173898 245062 174134
rect 245146 173898 245382 174134
rect 244826 138218 245062 138454
rect 245146 138218 245382 138454
rect 244826 137898 245062 138134
rect 245146 137898 245382 138134
rect 244826 102218 245062 102454
rect 245146 102218 245382 102454
rect 244826 101898 245062 102134
rect 245146 101898 245382 102134
rect 244826 66218 245062 66454
rect 245146 66218 245382 66454
rect 244826 65898 245062 66134
rect 245146 65898 245382 66134
rect 244826 30218 245062 30454
rect 245146 30218 245382 30454
rect 244826 29898 245062 30134
rect 245146 29898 245382 30134
rect 244826 -6342 245062 -6106
rect 245146 -6342 245382 -6106
rect 244826 -6662 245062 -6426
rect 245146 -6662 245382 -6426
rect 249326 711322 249562 711558
rect 249646 711322 249882 711558
rect 249326 711002 249562 711238
rect 249646 711002 249882 711238
rect 249326 682718 249562 682954
rect 249646 682718 249882 682954
rect 249326 682398 249562 682634
rect 249646 682398 249882 682634
rect 249326 646718 249562 646954
rect 249646 646718 249882 646954
rect 249326 646398 249562 646634
rect 249646 646398 249882 646634
rect 249326 610718 249562 610954
rect 249646 610718 249882 610954
rect 249326 610398 249562 610634
rect 249646 610398 249882 610634
rect 249326 574718 249562 574954
rect 249646 574718 249882 574954
rect 249326 574398 249562 574634
rect 249646 574398 249882 574634
rect 249326 538718 249562 538954
rect 249646 538718 249882 538954
rect 249326 538398 249562 538634
rect 249646 538398 249882 538634
rect 249326 502718 249562 502954
rect 249646 502718 249882 502954
rect 249326 502398 249562 502634
rect 249646 502398 249882 502634
rect 249326 466718 249562 466954
rect 249646 466718 249882 466954
rect 249326 466398 249562 466634
rect 249646 466398 249882 466634
rect 249326 430718 249562 430954
rect 249646 430718 249882 430954
rect 249326 430398 249562 430634
rect 249646 430398 249882 430634
rect 249326 394718 249562 394954
rect 249646 394718 249882 394954
rect 249326 394398 249562 394634
rect 249646 394398 249882 394634
rect 249326 358718 249562 358954
rect 249646 358718 249882 358954
rect 249326 358398 249562 358634
rect 249646 358398 249882 358634
rect 249326 322718 249562 322954
rect 249646 322718 249882 322954
rect 249326 322398 249562 322634
rect 249646 322398 249882 322634
rect 249326 286718 249562 286954
rect 249646 286718 249882 286954
rect 249326 286398 249562 286634
rect 249646 286398 249882 286634
rect 249326 250718 249562 250954
rect 249646 250718 249882 250954
rect 249326 250398 249562 250634
rect 249646 250398 249882 250634
rect 249326 214718 249562 214954
rect 249646 214718 249882 214954
rect 249326 214398 249562 214634
rect 249646 214398 249882 214634
rect 249326 178718 249562 178954
rect 249646 178718 249882 178954
rect 249326 178398 249562 178634
rect 249646 178398 249882 178634
rect 249326 142718 249562 142954
rect 249646 142718 249882 142954
rect 249326 142398 249562 142634
rect 249646 142398 249882 142634
rect 249326 106718 249562 106954
rect 249646 106718 249882 106954
rect 249326 106398 249562 106634
rect 249646 106398 249882 106634
rect 249326 70718 249562 70954
rect 249646 70718 249882 70954
rect 249326 70398 249562 70634
rect 249646 70398 249882 70634
rect 249326 34718 249562 34954
rect 249646 34718 249882 34954
rect 249326 34398 249562 34634
rect 249646 34398 249882 34634
rect 249326 -7302 249562 -7066
rect 249646 -7302 249882 -7066
rect 249326 -7622 249562 -7386
rect 249646 -7622 249882 -7386
rect 253826 704602 254062 704838
rect 254146 704602 254382 704838
rect 253826 704282 254062 704518
rect 254146 704282 254382 704518
rect 253826 687218 254062 687454
rect 254146 687218 254382 687454
rect 253826 686898 254062 687134
rect 254146 686898 254382 687134
rect 253826 651218 254062 651454
rect 254146 651218 254382 651454
rect 253826 650898 254062 651134
rect 254146 650898 254382 651134
rect 253826 615218 254062 615454
rect 254146 615218 254382 615454
rect 253826 614898 254062 615134
rect 254146 614898 254382 615134
rect 253826 579218 254062 579454
rect 254146 579218 254382 579454
rect 253826 578898 254062 579134
rect 254146 578898 254382 579134
rect 253826 543218 254062 543454
rect 254146 543218 254382 543454
rect 253826 542898 254062 543134
rect 254146 542898 254382 543134
rect 253826 507218 254062 507454
rect 254146 507218 254382 507454
rect 253826 506898 254062 507134
rect 254146 506898 254382 507134
rect 253826 471218 254062 471454
rect 254146 471218 254382 471454
rect 253826 470898 254062 471134
rect 254146 470898 254382 471134
rect 253826 435218 254062 435454
rect 254146 435218 254382 435454
rect 253826 434898 254062 435134
rect 254146 434898 254382 435134
rect 253826 399218 254062 399454
rect 254146 399218 254382 399454
rect 253826 398898 254062 399134
rect 254146 398898 254382 399134
rect 253826 363218 254062 363454
rect 254146 363218 254382 363454
rect 253826 362898 254062 363134
rect 254146 362898 254382 363134
rect 253826 327218 254062 327454
rect 254146 327218 254382 327454
rect 253826 326898 254062 327134
rect 254146 326898 254382 327134
rect 253826 291218 254062 291454
rect 254146 291218 254382 291454
rect 253826 290898 254062 291134
rect 254146 290898 254382 291134
rect 253826 255218 254062 255454
rect 254146 255218 254382 255454
rect 253826 254898 254062 255134
rect 254146 254898 254382 255134
rect 253826 219218 254062 219454
rect 254146 219218 254382 219454
rect 253826 218898 254062 219134
rect 254146 218898 254382 219134
rect 253826 183218 254062 183454
rect 254146 183218 254382 183454
rect 253826 182898 254062 183134
rect 254146 182898 254382 183134
rect 253826 147218 254062 147454
rect 254146 147218 254382 147454
rect 253826 146898 254062 147134
rect 254146 146898 254382 147134
rect 253826 111218 254062 111454
rect 254146 111218 254382 111454
rect 253826 110898 254062 111134
rect 254146 110898 254382 111134
rect 253826 75218 254062 75454
rect 254146 75218 254382 75454
rect 253826 74898 254062 75134
rect 254146 74898 254382 75134
rect 253826 39218 254062 39454
rect 254146 39218 254382 39454
rect 253826 38898 254062 39134
rect 254146 38898 254382 39134
rect 253826 3218 254062 3454
rect 254146 3218 254382 3454
rect 253826 2898 254062 3134
rect 254146 2898 254382 3134
rect 253826 -582 254062 -346
rect 254146 -582 254382 -346
rect 253826 -902 254062 -666
rect 254146 -902 254382 -666
rect 258326 705562 258562 705798
rect 258646 705562 258882 705798
rect 258326 705242 258562 705478
rect 258646 705242 258882 705478
rect 258326 691718 258562 691954
rect 258646 691718 258882 691954
rect 258326 691398 258562 691634
rect 258646 691398 258882 691634
rect 258326 655718 258562 655954
rect 258646 655718 258882 655954
rect 258326 655398 258562 655634
rect 258646 655398 258882 655634
rect 258326 619718 258562 619954
rect 258646 619718 258882 619954
rect 258326 619398 258562 619634
rect 258646 619398 258882 619634
rect 258326 583718 258562 583954
rect 258646 583718 258882 583954
rect 258326 583398 258562 583634
rect 258646 583398 258882 583634
rect 258326 547718 258562 547954
rect 258646 547718 258882 547954
rect 258326 547398 258562 547634
rect 258646 547398 258882 547634
rect 258326 511718 258562 511954
rect 258646 511718 258882 511954
rect 258326 511398 258562 511634
rect 258646 511398 258882 511634
rect 258326 475718 258562 475954
rect 258646 475718 258882 475954
rect 258326 475398 258562 475634
rect 258646 475398 258882 475634
rect 258326 439718 258562 439954
rect 258646 439718 258882 439954
rect 258326 439398 258562 439634
rect 258646 439398 258882 439634
rect 258326 403718 258562 403954
rect 258646 403718 258882 403954
rect 258326 403398 258562 403634
rect 258646 403398 258882 403634
rect 258326 367718 258562 367954
rect 258646 367718 258882 367954
rect 258326 367398 258562 367634
rect 258646 367398 258882 367634
rect 258326 331718 258562 331954
rect 258646 331718 258882 331954
rect 258326 331398 258562 331634
rect 258646 331398 258882 331634
rect 258326 295718 258562 295954
rect 258646 295718 258882 295954
rect 258326 295398 258562 295634
rect 258646 295398 258882 295634
rect 258326 259718 258562 259954
rect 258646 259718 258882 259954
rect 258326 259398 258562 259634
rect 258646 259398 258882 259634
rect 258326 223718 258562 223954
rect 258646 223718 258882 223954
rect 258326 223398 258562 223634
rect 258646 223398 258882 223634
rect 258326 187718 258562 187954
rect 258646 187718 258882 187954
rect 258326 187398 258562 187634
rect 258646 187398 258882 187634
rect 258326 151718 258562 151954
rect 258646 151718 258882 151954
rect 258326 151398 258562 151634
rect 258646 151398 258882 151634
rect 258326 115718 258562 115954
rect 258646 115718 258882 115954
rect 258326 115398 258562 115634
rect 258646 115398 258882 115634
rect 258326 79718 258562 79954
rect 258646 79718 258882 79954
rect 258326 79398 258562 79634
rect 258646 79398 258882 79634
rect 258326 43718 258562 43954
rect 258646 43718 258882 43954
rect 258326 43398 258562 43634
rect 258646 43398 258882 43634
rect 258326 7718 258562 7954
rect 258646 7718 258882 7954
rect 258326 7398 258562 7634
rect 258646 7398 258882 7634
rect 258326 -1542 258562 -1306
rect 258646 -1542 258882 -1306
rect 258326 -1862 258562 -1626
rect 258646 -1862 258882 -1626
rect 262826 706522 263062 706758
rect 263146 706522 263382 706758
rect 262826 706202 263062 706438
rect 263146 706202 263382 706438
rect 262826 696218 263062 696454
rect 263146 696218 263382 696454
rect 262826 695898 263062 696134
rect 263146 695898 263382 696134
rect 262826 660218 263062 660454
rect 263146 660218 263382 660454
rect 262826 659898 263062 660134
rect 263146 659898 263382 660134
rect 262826 624218 263062 624454
rect 263146 624218 263382 624454
rect 262826 623898 263062 624134
rect 263146 623898 263382 624134
rect 262826 588218 263062 588454
rect 263146 588218 263382 588454
rect 262826 587898 263062 588134
rect 263146 587898 263382 588134
rect 262826 552218 263062 552454
rect 263146 552218 263382 552454
rect 262826 551898 263062 552134
rect 263146 551898 263382 552134
rect 262826 516218 263062 516454
rect 263146 516218 263382 516454
rect 262826 515898 263062 516134
rect 263146 515898 263382 516134
rect 262826 480218 263062 480454
rect 263146 480218 263382 480454
rect 262826 479898 263062 480134
rect 263146 479898 263382 480134
rect 262826 444218 263062 444454
rect 263146 444218 263382 444454
rect 262826 443898 263062 444134
rect 263146 443898 263382 444134
rect 262826 408218 263062 408454
rect 263146 408218 263382 408454
rect 262826 407898 263062 408134
rect 263146 407898 263382 408134
rect 262826 372218 263062 372454
rect 263146 372218 263382 372454
rect 262826 371898 263062 372134
rect 263146 371898 263382 372134
rect 262826 336218 263062 336454
rect 263146 336218 263382 336454
rect 262826 335898 263062 336134
rect 263146 335898 263382 336134
rect 262826 300218 263062 300454
rect 263146 300218 263382 300454
rect 262826 299898 263062 300134
rect 263146 299898 263382 300134
rect 262826 264218 263062 264454
rect 263146 264218 263382 264454
rect 262826 263898 263062 264134
rect 263146 263898 263382 264134
rect 262826 228218 263062 228454
rect 263146 228218 263382 228454
rect 262826 227898 263062 228134
rect 263146 227898 263382 228134
rect 262826 192218 263062 192454
rect 263146 192218 263382 192454
rect 262826 191898 263062 192134
rect 263146 191898 263382 192134
rect 262826 156218 263062 156454
rect 263146 156218 263382 156454
rect 262826 155898 263062 156134
rect 263146 155898 263382 156134
rect 262826 120218 263062 120454
rect 263146 120218 263382 120454
rect 262826 119898 263062 120134
rect 263146 119898 263382 120134
rect 262826 84218 263062 84454
rect 263146 84218 263382 84454
rect 262826 83898 263062 84134
rect 263146 83898 263382 84134
rect 262826 48218 263062 48454
rect 263146 48218 263382 48454
rect 262826 47898 263062 48134
rect 263146 47898 263382 48134
rect 262826 12218 263062 12454
rect 263146 12218 263382 12454
rect 262826 11898 263062 12134
rect 263146 11898 263382 12134
rect 262826 -2502 263062 -2266
rect 263146 -2502 263382 -2266
rect 262826 -2822 263062 -2586
rect 263146 -2822 263382 -2586
rect 267326 707482 267562 707718
rect 267646 707482 267882 707718
rect 267326 707162 267562 707398
rect 267646 707162 267882 707398
rect 267326 700718 267562 700954
rect 267646 700718 267882 700954
rect 267326 700398 267562 700634
rect 267646 700398 267882 700634
rect 267326 664718 267562 664954
rect 267646 664718 267882 664954
rect 267326 664398 267562 664634
rect 267646 664398 267882 664634
rect 267326 628718 267562 628954
rect 267646 628718 267882 628954
rect 267326 628398 267562 628634
rect 267646 628398 267882 628634
rect 267326 592718 267562 592954
rect 267646 592718 267882 592954
rect 267326 592398 267562 592634
rect 267646 592398 267882 592634
rect 267326 556718 267562 556954
rect 267646 556718 267882 556954
rect 267326 556398 267562 556634
rect 267646 556398 267882 556634
rect 267326 520718 267562 520954
rect 267646 520718 267882 520954
rect 267326 520398 267562 520634
rect 267646 520398 267882 520634
rect 267326 484718 267562 484954
rect 267646 484718 267882 484954
rect 267326 484398 267562 484634
rect 267646 484398 267882 484634
rect 267326 448718 267562 448954
rect 267646 448718 267882 448954
rect 267326 448398 267562 448634
rect 267646 448398 267882 448634
rect 267326 412718 267562 412954
rect 267646 412718 267882 412954
rect 267326 412398 267562 412634
rect 267646 412398 267882 412634
rect 267326 376718 267562 376954
rect 267646 376718 267882 376954
rect 267326 376398 267562 376634
rect 267646 376398 267882 376634
rect 267326 340718 267562 340954
rect 267646 340718 267882 340954
rect 267326 340398 267562 340634
rect 267646 340398 267882 340634
rect 267326 304718 267562 304954
rect 267646 304718 267882 304954
rect 267326 304398 267562 304634
rect 267646 304398 267882 304634
rect 267326 268718 267562 268954
rect 267646 268718 267882 268954
rect 267326 268398 267562 268634
rect 267646 268398 267882 268634
rect 267326 232718 267562 232954
rect 267646 232718 267882 232954
rect 267326 232398 267562 232634
rect 267646 232398 267882 232634
rect 267326 196718 267562 196954
rect 267646 196718 267882 196954
rect 267326 196398 267562 196634
rect 267646 196398 267882 196634
rect 267326 160718 267562 160954
rect 267646 160718 267882 160954
rect 267326 160398 267562 160634
rect 267646 160398 267882 160634
rect 267326 124718 267562 124954
rect 267646 124718 267882 124954
rect 267326 124398 267562 124634
rect 267646 124398 267882 124634
rect 267326 88718 267562 88954
rect 267646 88718 267882 88954
rect 267326 88398 267562 88634
rect 267646 88398 267882 88634
rect 267326 52718 267562 52954
rect 267646 52718 267882 52954
rect 267326 52398 267562 52634
rect 267646 52398 267882 52634
rect 267326 16718 267562 16954
rect 267646 16718 267882 16954
rect 267326 16398 267562 16634
rect 267646 16398 267882 16634
rect 267326 -3462 267562 -3226
rect 267646 -3462 267882 -3226
rect 267326 -3782 267562 -3546
rect 267646 -3782 267882 -3546
rect 271826 708442 272062 708678
rect 272146 708442 272382 708678
rect 271826 708122 272062 708358
rect 272146 708122 272382 708358
rect 271826 669218 272062 669454
rect 272146 669218 272382 669454
rect 271826 668898 272062 669134
rect 272146 668898 272382 669134
rect 271826 633218 272062 633454
rect 272146 633218 272382 633454
rect 271826 632898 272062 633134
rect 272146 632898 272382 633134
rect 271826 597218 272062 597454
rect 272146 597218 272382 597454
rect 271826 596898 272062 597134
rect 272146 596898 272382 597134
rect 271826 561218 272062 561454
rect 272146 561218 272382 561454
rect 271826 560898 272062 561134
rect 272146 560898 272382 561134
rect 271826 525218 272062 525454
rect 272146 525218 272382 525454
rect 271826 524898 272062 525134
rect 272146 524898 272382 525134
rect 271826 489218 272062 489454
rect 272146 489218 272382 489454
rect 271826 488898 272062 489134
rect 272146 488898 272382 489134
rect 271826 453218 272062 453454
rect 272146 453218 272382 453454
rect 271826 452898 272062 453134
rect 272146 452898 272382 453134
rect 271826 417218 272062 417454
rect 272146 417218 272382 417454
rect 271826 416898 272062 417134
rect 272146 416898 272382 417134
rect 271826 381218 272062 381454
rect 272146 381218 272382 381454
rect 271826 380898 272062 381134
rect 272146 380898 272382 381134
rect 271826 345218 272062 345454
rect 272146 345218 272382 345454
rect 271826 344898 272062 345134
rect 272146 344898 272382 345134
rect 271826 309218 272062 309454
rect 272146 309218 272382 309454
rect 271826 308898 272062 309134
rect 272146 308898 272382 309134
rect 271826 273218 272062 273454
rect 272146 273218 272382 273454
rect 271826 272898 272062 273134
rect 272146 272898 272382 273134
rect 271826 237218 272062 237454
rect 272146 237218 272382 237454
rect 271826 236898 272062 237134
rect 272146 236898 272382 237134
rect 271826 201218 272062 201454
rect 272146 201218 272382 201454
rect 271826 200898 272062 201134
rect 272146 200898 272382 201134
rect 271826 165218 272062 165454
rect 272146 165218 272382 165454
rect 271826 164898 272062 165134
rect 272146 164898 272382 165134
rect 271826 129218 272062 129454
rect 272146 129218 272382 129454
rect 271826 128898 272062 129134
rect 272146 128898 272382 129134
rect 271826 93218 272062 93454
rect 272146 93218 272382 93454
rect 271826 92898 272062 93134
rect 272146 92898 272382 93134
rect 271826 57218 272062 57454
rect 272146 57218 272382 57454
rect 271826 56898 272062 57134
rect 272146 56898 272382 57134
rect 271826 21218 272062 21454
rect 272146 21218 272382 21454
rect 271826 20898 272062 21134
rect 272146 20898 272382 21134
rect 271826 -4422 272062 -4186
rect 272146 -4422 272382 -4186
rect 271826 -4742 272062 -4506
rect 272146 -4742 272382 -4506
rect 276326 709402 276562 709638
rect 276646 709402 276882 709638
rect 276326 709082 276562 709318
rect 276646 709082 276882 709318
rect 276326 673718 276562 673954
rect 276646 673718 276882 673954
rect 276326 673398 276562 673634
rect 276646 673398 276882 673634
rect 276326 637718 276562 637954
rect 276646 637718 276882 637954
rect 276326 637398 276562 637634
rect 276646 637398 276882 637634
rect 276326 601718 276562 601954
rect 276646 601718 276882 601954
rect 276326 601398 276562 601634
rect 276646 601398 276882 601634
rect 276326 565718 276562 565954
rect 276646 565718 276882 565954
rect 276326 565398 276562 565634
rect 276646 565398 276882 565634
rect 276326 529718 276562 529954
rect 276646 529718 276882 529954
rect 276326 529398 276562 529634
rect 276646 529398 276882 529634
rect 276326 493718 276562 493954
rect 276646 493718 276882 493954
rect 276326 493398 276562 493634
rect 276646 493398 276882 493634
rect 276326 457718 276562 457954
rect 276646 457718 276882 457954
rect 276326 457398 276562 457634
rect 276646 457398 276882 457634
rect 276326 421718 276562 421954
rect 276646 421718 276882 421954
rect 276326 421398 276562 421634
rect 276646 421398 276882 421634
rect 276326 385718 276562 385954
rect 276646 385718 276882 385954
rect 276326 385398 276562 385634
rect 276646 385398 276882 385634
rect 276326 349718 276562 349954
rect 276646 349718 276882 349954
rect 276326 349398 276562 349634
rect 276646 349398 276882 349634
rect 276326 313718 276562 313954
rect 276646 313718 276882 313954
rect 276326 313398 276562 313634
rect 276646 313398 276882 313634
rect 276326 277718 276562 277954
rect 276646 277718 276882 277954
rect 276326 277398 276562 277634
rect 276646 277398 276882 277634
rect 276326 241718 276562 241954
rect 276646 241718 276882 241954
rect 276326 241398 276562 241634
rect 276646 241398 276882 241634
rect 276326 205718 276562 205954
rect 276646 205718 276882 205954
rect 276326 205398 276562 205634
rect 276646 205398 276882 205634
rect 276326 169718 276562 169954
rect 276646 169718 276882 169954
rect 276326 169398 276562 169634
rect 276646 169398 276882 169634
rect 276326 133718 276562 133954
rect 276646 133718 276882 133954
rect 276326 133398 276562 133634
rect 276646 133398 276882 133634
rect 276326 97718 276562 97954
rect 276646 97718 276882 97954
rect 276326 97398 276562 97634
rect 276646 97398 276882 97634
rect 276326 61718 276562 61954
rect 276646 61718 276882 61954
rect 276326 61398 276562 61634
rect 276646 61398 276882 61634
rect 276326 25718 276562 25954
rect 276646 25718 276882 25954
rect 276326 25398 276562 25634
rect 276646 25398 276882 25634
rect 276326 -5382 276562 -5146
rect 276646 -5382 276882 -5146
rect 276326 -5702 276562 -5466
rect 276646 -5702 276882 -5466
rect 280826 710362 281062 710598
rect 281146 710362 281382 710598
rect 280826 710042 281062 710278
rect 281146 710042 281382 710278
rect 280826 678218 281062 678454
rect 281146 678218 281382 678454
rect 280826 677898 281062 678134
rect 281146 677898 281382 678134
rect 280826 642218 281062 642454
rect 281146 642218 281382 642454
rect 280826 641898 281062 642134
rect 281146 641898 281382 642134
rect 280826 606218 281062 606454
rect 281146 606218 281382 606454
rect 280826 605898 281062 606134
rect 281146 605898 281382 606134
rect 280826 570218 281062 570454
rect 281146 570218 281382 570454
rect 280826 569898 281062 570134
rect 281146 569898 281382 570134
rect 280826 534218 281062 534454
rect 281146 534218 281382 534454
rect 280826 533898 281062 534134
rect 281146 533898 281382 534134
rect 280826 498218 281062 498454
rect 281146 498218 281382 498454
rect 280826 497898 281062 498134
rect 281146 497898 281382 498134
rect 280826 462218 281062 462454
rect 281146 462218 281382 462454
rect 280826 461898 281062 462134
rect 281146 461898 281382 462134
rect 280826 426218 281062 426454
rect 281146 426218 281382 426454
rect 280826 425898 281062 426134
rect 281146 425898 281382 426134
rect 280826 390218 281062 390454
rect 281146 390218 281382 390454
rect 280826 389898 281062 390134
rect 281146 389898 281382 390134
rect 280826 354218 281062 354454
rect 281146 354218 281382 354454
rect 280826 353898 281062 354134
rect 281146 353898 281382 354134
rect 280826 318218 281062 318454
rect 281146 318218 281382 318454
rect 280826 317898 281062 318134
rect 281146 317898 281382 318134
rect 280826 282218 281062 282454
rect 281146 282218 281382 282454
rect 280826 281898 281062 282134
rect 281146 281898 281382 282134
rect 280826 246218 281062 246454
rect 281146 246218 281382 246454
rect 280826 245898 281062 246134
rect 281146 245898 281382 246134
rect 280826 210218 281062 210454
rect 281146 210218 281382 210454
rect 280826 209898 281062 210134
rect 281146 209898 281382 210134
rect 280826 174218 281062 174454
rect 281146 174218 281382 174454
rect 280826 173898 281062 174134
rect 281146 173898 281382 174134
rect 280826 138218 281062 138454
rect 281146 138218 281382 138454
rect 280826 137898 281062 138134
rect 281146 137898 281382 138134
rect 280826 102218 281062 102454
rect 281146 102218 281382 102454
rect 280826 101898 281062 102134
rect 281146 101898 281382 102134
rect 280826 66218 281062 66454
rect 281146 66218 281382 66454
rect 280826 65898 281062 66134
rect 281146 65898 281382 66134
rect 280826 30218 281062 30454
rect 281146 30218 281382 30454
rect 280826 29898 281062 30134
rect 281146 29898 281382 30134
rect 280826 -6342 281062 -6106
rect 281146 -6342 281382 -6106
rect 280826 -6662 281062 -6426
rect 281146 -6662 281382 -6426
rect 285326 711322 285562 711558
rect 285646 711322 285882 711558
rect 285326 711002 285562 711238
rect 285646 711002 285882 711238
rect 285326 682718 285562 682954
rect 285646 682718 285882 682954
rect 285326 682398 285562 682634
rect 285646 682398 285882 682634
rect 285326 646718 285562 646954
rect 285646 646718 285882 646954
rect 285326 646398 285562 646634
rect 285646 646398 285882 646634
rect 285326 610718 285562 610954
rect 285646 610718 285882 610954
rect 285326 610398 285562 610634
rect 285646 610398 285882 610634
rect 285326 574718 285562 574954
rect 285646 574718 285882 574954
rect 285326 574398 285562 574634
rect 285646 574398 285882 574634
rect 285326 538718 285562 538954
rect 285646 538718 285882 538954
rect 285326 538398 285562 538634
rect 285646 538398 285882 538634
rect 285326 502718 285562 502954
rect 285646 502718 285882 502954
rect 285326 502398 285562 502634
rect 285646 502398 285882 502634
rect 285326 466718 285562 466954
rect 285646 466718 285882 466954
rect 285326 466398 285562 466634
rect 285646 466398 285882 466634
rect 285326 430718 285562 430954
rect 285646 430718 285882 430954
rect 285326 430398 285562 430634
rect 285646 430398 285882 430634
rect 285326 394718 285562 394954
rect 285646 394718 285882 394954
rect 285326 394398 285562 394634
rect 285646 394398 285882 394634
rect 285326 358718 285562 358954
rect 285646 358718 285882 358954
rect 285326 358398 285562 358634
rect 285646 358398 285882 358634
rect 285326 322718 285562 322954
rect 285646 322718 285882 322954
rect 285326 322398 285562 322634
rect 285646 322398 285882 322634
rect 285326 286718 285562 286954
rect 285646 286718 285882 286954
rect 285326 286398 285562 286634
rect 285646 286398 285882 286634
rect 285326 250718 285562 250954
rect 285646 250718 285882 250954
rect 285326 250398 285562 250634
rect 285646 250398 285882 250634
rect 285326 214718 285562 214954
rect 285646 214718 285882 214954
rect 285326 214398 285562 214634
rect 285646 214398 285882 214634
rect 285326 178718 285562 178954
rect 285646 178718 285882 178954
rect 285326 178398 285562 178634
rect 285646 178398 285882 178634
rect 285326 142718 285562 142954
rect 285646 142718 285882 142954
rect 285326 142398 285562 142634
rect 285646 142398 285882 142634
rect 285326 106718 285562 106954
rect 285646 106718 285882 106954
rect 285326 106398 285562 106634
rect 285646 106398 285882 106634
rect 285326 70718 285562 70954
rect 285646 70718 285882 70954
rect 285326 70398 285562 70634
rect 285646 70398 285882 70634
rect 285326 34718 285562 34954
rect 285646 34718 285882 34954
rect 285326 34398 285562 34634
rect 285646 34398 285882 34634
rect 285326 -7302 285562 -7066
rect 285646 -7302 285882 -7066
rect 285326 -7622 285562 -7386
rect 285646 -7622 285882 -7386
rect 289826 704602 290062 704838
rect 290146 704602 290382 704838
rect 289826 704282 290062 704518
rect 290146 704282 290382 704518
rect 289826 687218 290062 687454
rect 290146 687218 290382 687454
rect 289826 686898 290062 687134
rect 290146 686898 290382 687134
rect 289826 651218 290062 651454
rect 290146 651218 290382 651454
rect 289826 650898 290062 651134
rect 290146 650898 290382 651134
rect 289826 615218 290062 615454
rect 290146 615218 290382 615454
rect 289826 614898 290062 615134
rect 290146 614898 290382 615134
rect 289826 579218 290062 579454
rect 290146 579218 290382 579454
rect 289826 578898 290062 579134
rect 290146 578898 290382 579134
rect 289826 543218 290062 543454
rect 290146 543218 290382 543454
rect 289826 542898 290062 543134
rect 290146 542898 290382 543134
rect 289826 507218 290062 507454
rect 290146 507218 290382 507454
rect 289826 506898 290062 507134
rect 290146 506898 290382 507134
rect 289826 471218 290062 471454
rect 290146 471218 290382 471454
rect 289826 470898 290062 471134
rect 290146 470898 290382 471134
rect 289826 435218 290062 435454
rect 290146 435218 290382 435454
rect 289826 434898 290062 435134
rect 290146 434898 290382 435134
rect 289826 399218 290062 399454
rect 290146 399218 290382 399454
rect 289826 398898 290062 399134
rect 290146 398898 290382 399134
rect 289826 363218 290062 363454
rect 290146 363218 290382 363454
rect 289826 362898 290062 363134
rect 290146 362898 290382 363134
rect 289826 327218 290062 327454
rect 290146 327218 290382 327454
rect 289826 326898 290062 327134
rect 290146 326898 290382 327134
rect 289826 291218 290062 291454
rect 290146 291218 290382 291454
rect 289826 290898 290062 291134
rect 290146 290898 290382 291134
rect 289826 255218 290062 255454
rect 290146 255218 290382 255454
rect 289826 254898 290062 255134
rect 290146 254898 290382 255134
rect 289826 219218 290062 219454
rect 290146 219218 290382 219454
rect 289826 218898 290062 219134
rect 290146 218898 290382 219134
rect 289826 183218 290062 183454
rect 290146 183218 290382 183454
rect 289826 182898 290062 183134
rect 290146 182898 290382 183134
rect 289826 147218 290062 147454
rect 290146 147218 290382 147454
rect 289826 146898 290062 147134
rect 290146 146898 290382 147134
rect 289826 111218 290062 111454
rect 290146 111218 290382 111454
rect 289826 110898 290062 111134
rect 290146 110898 290382 111134
rect 289826 75218 290062 75454
rect 290146 75218 290382 75454
rect 289826 74898 290062 75134
rect 290146 74898 290382 75134
rect 289826 39218 290062 39454
rect 290146 39218 290382 39454
rect 289826 38898 290062 39134
rect 290146 38898 290382 39134
rect 289826 3218 290062 3454
rect 290146 3218 290382 3454
rect 289826 2898 290062 3134
rect 290146 2898 290382 3134
rect 289826 -582 290062 -346
rect 290146 -582 290382 -346
rect 289826 -902 290062 -666
rect 290146 -902 290382 -666
rect 294326 705562 294562 705798
rect 294646 705562 294882 705798
rect 294326 705242 294562 705478
rect 294646 705242 294882 705478
rect 294326 691718 294562 691954
rect 294646 691718 294882 691954
rect 294326 691398 294562 691634
rect 294646 691398 294882 691634
rect 294326 655718 294562 655954
rect 294646 655718 294882 655954
rect 294326 655398 294562 655634
rect 294646 655398 294882 655634
rect 294326 619718 294562 619954
rect 294646 619718 294882 619954
rect 294326 619398 294562 619634
rect 294646 619398 294882 619634
rect 294326 583718 294562 583954
rect 294646 583718 294882 583954
rect 294326 583398 294562 583634
rect 294646 583398 294882 583634
rect 294326 547718 294562 547954
rect 294646 547718 294882 547954
rect 294326 547398 294562 547634
rect 294646 547398 294882 547634
rect 294326 511718 294562 511954
rect 294646 511718 294882 511954
rect 294326 511398 294562 511634
rect 294646 511398 294882 511634
rect 294326 475718 294562 475954
rect 294646 475718 294882 475954
rect 294326 475398 294562 475634
rect 294646 475398 294882 475634
rect 294326 439718 294562 439954
rect 294646 439718 294882 439954
rect 294326 439398 294562 439634
rect 294646 439398 294882 439634
rect 294326 403718 294562 403954
rect 294646 403718 294882 403954
rect 294326 403398 294562 403634
rect 294646 403398 294882 403634
rect 294326 367718 294562 367954
rect 294646 367718 294882 367954
rect 294326 367398 294562 367634
rect 294646 367398 294882 367634
rect 294326 331718 294562 331954
rect 294646 331718 294882 331954
rect 294326 331398 294562 331634
rect 294646 331398 294882 331634
rect 294326 295718 294562 295954
rect 294646 295718 294882 295954
rect 294326 295398 294562 295634
rect 294646 295398 294882 295634
rect 294326 259718 294562 259954
rect 294646 259718 294882 259954
rect 294326 259398 294562 259634
rect 294646 259398 294882 259634
rect 294326 223718 294562 223954
rect 294646 223718 294882 223954
rect 294326 223398 294562 223634
rect 294646 223398 294882 223634
rect 294326 187718 294562 187954
rect 294646 187718 294882 187954
rect 294326 187398 294562 187634
rect 294646 187398 294882 187634
rect 294326 151718 294562 151954
rect 294646 151718 294882 151954
rect 294326 151398 294562 151634
rect 294646 151398 294882 151634
rect 294326 115718 294562 115954
rect 294646 115718 294882 115954
rect 294326 115398 294562 115634
rect 294646 115398 294882 115634
rect 294326 79718 294562 79954
rect 294646 79718 294882 79954
rect 294326 79398 294562 79634
rect 294646 79398 294882 79634
rect 294326 43718 294562 43954
rect 294646 43718 294882 43954
rect 294326 43398 294562 43634
rect 294646 43398 294882 43634
rect 294326 7718 294562 7954
rect 294646 7718 294882 7954
rect 294326 7398 294562 7634
rect 294646 7398 294882 7634
rect 294326 -1542 294562 -1306
rect 294646 -1542 294882 -1306
rect 294326 -1862 294562 -1626
rect 294646 -1862 294882 -1626
rect 298826 706522 299062 706758
rect 299146 706522 299382 706758
rect 298826 706202 299062 706438
rect 299146 706202 299382 706438
rect 298826 696218 299062 696454
rect 299146 696218 299382 696454
rect 298826 695898 299062 696134
rect 299146 695898 299382 696134
rect 298826 660218 299062 660454
rect 299146 660218 299382 660454
rect 298826 659898 299062 660134
rect 299146 659898 299382 660134
rect 298826 624218 299062 624454
rect 299146 624218 299382 624454
rect 298826 623898 299062 624134
rect 299146 623898 299382 624134
rect 298826 588218 299062 588454
rect 299146 588218 299382 588454
rect 298826 587898 299062 588134
rect 299146 587898 299382 588134
rect 298826 552218 299062 552454
rect 299146 552218 299382 552454
rect 298826 551898 299062 552134
rect 299146 551898 299382 552134
rect 298826 516218 299062 516454
rect 299146 516218 299382 516454
rect 298826 515898 299062 516134
rect 299146 515898 299382 516134
rect 298826 480218 299062 480454
rect 299146 480218 299382 480454
rect 298826 479898 299062 480134
rect 299146 479898 299382 480134
rect 298826 444218 299062 444454
rect 299146 444218 299382 444454
rect 298826 443898 299062 444134
rect 299146 443898 299382 444134
rect 298826 408218 299062 408454
rect 299146 408218 299382 408454
rect 298826 407898 299062 408134
rect 299146 407898 299382 408134
rect 298826 372218 299062 372454
rect 299146 372218 299382 372454
rect 298826 371898 299062 372134
rect 299146 371898 299382 372134
rect 298826 336218 299062 336454
rect 299146 336218 299382 336454
rect 298826 335898 299062 336134
rect 299146 335898 299382 336134
rect 298826 300218 299062 300454
rect 299146 300218 299382 300454
rect 298826 299898 299062 300134
rect 299146 299898 299382 300134
rect 298826 264218 299062 264454
rect 299146 264218 299382 264454
rect 298826 263898 299062 264134
rect 299146 263898 299382 264134
rect 298826 228218 299062 228454
rect 299146 228218 299382 228454
rect 298826 227898 299062 228134
rect 299146 227898 299382 228134
rect 298826 192218 299062 192454
rect 299146 192218 299382 192454
rect 298826 191898 299062 192134
rect 299146 191898 299382 192134
rect 298826 156218 299062 156454
rect 299146 156218 299382 156454
rect 298826 155898 299062 156134
rect 299146 155898 299382 156134
rect 298826 120218 299062 120454
rect 299146 120218 299382 120454
rect 298826 119898 299062 120134
rect 299146 119898 299382 120134
rect 298826 84218 299062 84454
rect 299146 84218 299382 84454
rect 298826 83898 299062 84134
rect 299146 83898 299382 84134
rect 298826 48218 299062 48454
rect 299146 48218 299382 48454
rect 298826 47898 299062 48134
rect 299146 47898 299382 48134
rect 298826 12218 299062 12454
rect 299146 12218 299382 12454
rect 298826 11898 299062 12134
rect 299146 11898 299382 12134
rect 298826 -2502 299062 -2266
rect 299146 -2502 299382 -2266
rect 298826 -2822 299062 -2586
rect 299146 -2822 299382 -2586
rect 303326 707482 303562 707718
rect 303646 707482 303882 707718
rect 303326 707162 303562 707398
rect 303646 707162 303882 707398
rect 303326 700718 303562 700954
rect 303646 700718 303882 700954
rect 303326 700398 303562 700634
rect 303646 700398 303882 700634
rect 303326 664718 303562 664954
rect 303646 664718 303882 664954
rect 303326 664398 303562 664634
rect 303646 664398 303882 664634
rect 303326 628718 303562 628954
rect 303646 628718 303882 628954
rect 303326 628398 303562 628634
rect 303646 628398 303882 628634
rect 303326 592718 303562 592954
rect 303646 592718 303882 592954
rect 303326 592398 303562 592634
rect 303646 592398 303882 592634
rect 303326 556718 303562 556954
rect 303646 556718 303882 556954
rect 303326 556398 303562 556634
rect 303646 556398 303882 556634
rect 303326 520718 303562 520954
rect 303646 520718 303882 520954
rect 303326 520398 303562 520634
rect 303646 520398 303882 520634
rect 303326 484718 303562 484954
rect 303646 484718 303882 484954
rect 303326 484398 303562 484634
rect 303646 484398 303882 484634
rect 303326 448718 303562 448954
rect 303646 448718 303882 448954
rect 303326 448398 303562 448634
rect 303646 448398 303882 448634
rect 303326 412718 303562 412954
rect 303646 412718 303882 412954
rect 303326 412398 303562 412634
rect 303646 412398 303882 412634
rect 303326 376718 303562 376954
rect 303646 376718 303882 376954
rect 303326 376398 303562 376634
rect 303646 376398 303882 376634
rect 303326 340718 303562 340954
rect 303646 340718 303882 340954
rect 303326 340398 303562 340634
rect 303646 340398 303882 340634
rect 303326 304718 303562 304954
rect 303646 304718 303882 304954
rect 303326 304398 303562 304634
rect 303646 304398 303882 304634
rect 303326 268718 303562 268954
rect 303646 268718 303882 268954
rect 303326 268398 303562 268634
rect 303646 268398 303882 268634
rect 303326 232718 303562 232954
rect 303646 232718 303882 232954
rect 303326 232398 303562 232634
rect 303646 232398 303882 232634
rect 303326 196718 303562 196954
rect 303646 196718 303882 196954
rect 303326 196398 303562 196634
rect 303646 196398 303882 196634
rect 303326 160718 303562 160954
rect 303646 160718 303882 160954
rect 303326 160398 303562 160634
rect 303646 160398 303882 160634
rect 303326 124718 303562 124954
rect 303646 124718 303882 124954
rect 303326 124398 303562 124634
rect 303646 124398 303882 124634
rect 303326 88718 303562 88954
rect 303646 88718 303882 88954
rect 303326 88398 303562 88634
rect 303646 88398 303882 88634
rect 303326 52718 303562 52954
rect 303646 52718 303882 52954
rect 303326 52398 303562 52634
rect 303646 52398 303882 52634
rect 303326 16718 303562 16954
rect 303646 16718 303882 16954
rect 303326 16398 303562 16634
rect 303646 16398 303882 16634
rect 303326 -3462 303562 -3226
rect 303646 -3462 303882 -3226
rect 303326 -3782 303562 -3546
rect 303646 -3782 303882 -3546
rect 307826 708442 308062 708678
rect 308146 708442 308382 708678
rect 307826 708122 308062 708358
rect 308146 708122 308382 708358
rect 307826 669218 308062 669454
rect 308146 669218 308382 669454
rect 307826 668898 308062 669134
rect 308146 668898 308382 669134
rect 307826 633218 308062 633454
rect 308146 633218 308382 633454
rect 307826 632898 308062 633134
rect 308146 632898 308382 633134
rect 307826 597218 308062 597454
rect 308146 597218 308382 597454
rect 307826 596898 308062 597134
rect 308146 596898 308382 597134
rect 307826 561218 308062 561454
rect 308146 561218 308382 561454
rect 307826 560898 308062 561134
rect 308146 560898 308382 561134
rect 307826 525218 308062 525454
rect 308146 525218 308382 525454
rect 307826 524898 308062 525134
rect 308146 524898 308382 525134
rect 307826 489218 308062 489454
rect 308146 489218 308382 489454
rect 307826 488898 308062 489134
rect 308146 488898 308382 489134
rect 307826 453218 308062 453454
rect 308146 453218 308382 453454
rect 307826 452898 308062 453134
rect 308146 452898 308382 453134
rect 307826 417218 308062 417454
rect 308146 417218 308382 417454
rect 307826 416898 308062 417134
rect 308146 416898 308382 417134
rect 307826 381218 308062 381454
rect 308146 381218 308382 381454
rect 307826 380898 308062 381134
rect 308146 380898 308382 381134
rect 307826 345218 308062 345454
rect 308146 345218 308382 345454
rect 307826 344898 308062 345134
rect 308146 344898 308382 345134
rect 307826 309218 308062 309454
rect 308146 309218 308382 309454
rect 307826 308898 308062 309134
rect 308146 308898 308382 309134
rect 307826 273218 308062 273454
rect 308146 273218 308382 273454
rect 307826 272898 308062 273134
rect 308146 272898 308382 273134
rect 307826 237218 308062 237454
rect 308146 237218 308382 237454
rect 307826 236898 308062 237134
rect 308146 236898 308382 237134
rect 307826 201218 308062 201454
rect 308146 201218 308382 201454
rect 307826 200898 308062 201134
rect 308146 200898 308382 201134
rect 307826 165218 308062 165454
rect 308146 165218 308382 165454
rect 307826 164898 308062 165134
rect 308146 164898 308382 165134
rect 307826 129218 308062 129454
rect 308146 129218 308382 129454
rect 307826 128898 308062 129134
rect 308146 128898 308382 129134
rect 307826 93218 308062 93454
rect 308146 93218 308382 93454
rect 307826 92898 308062 93134
rect 308146 92898 308382 93134
rect 307826 57218 308062 57454
rect 308146 57218 308382 57454
rect 307826 56898 308062 57134
rect 308146 56898 308382 57134
rect 307826 21218 308062 21454
rect 308146 21218 308382 21454
rect 307826 20898 308062 21134
rect 308146 20898 308382 21134
rect 307826 -4422 308062 -4186
rect 308146 -4422 308382 -4186
rect 307826 -4742 308062 -4506
rect 308146 -4742 308382 -4506
rect 312326 709402 312562 709638
rect 312646 709402 312882 709638
rect 312326 709082 312562 709318
rect 312646 709082 312882 709318
rect 312326 673718 312562 673954
rect 312646 673718 312882 673954
rect 312326 673398 312562 673634
rect 312646 673398 312882 673634
rect 312326 637718 312562 637954
rect 312646 637718 312882 637954
rect 312326 637398 312562 637634
rect 312646 637398 312882 637634
rect 312326 601718 312562 601954
rect 312646 601718 312882 601954
rect 312326 601398 312562 601634
rect 312646 601398 312882 601634
rect 312326 565718 312562 565954
rect 312646 565718 312882 565954
rect 312326 565398 312562 565634
rect 312646 565398 312882 565634
rect 312326 529718 312562 529954
rect 312646 529718 312882 529954
rect 312326 529398 312562 529634
rect 312646 529398 312882 529634
rect 312326 493718 312562 493954
rect 312646 493718 312882 493954
rect 312326 493398 312562 493634
rect 312646 493398 312882 493634
rect 312326 457718 312562 457954
rect 312646 457718 312882 457954
rect 312326 457398 312562 457634
rect 312646 457398 312882 457634
rect 312326 421718 312562 421954
rect 312646 421718 312882 421954
rect 312326 421398 312562 421634
rect 312646 421398 312882 421634
rect 312326 385718 312562 385954
rect 312646 385718 312882 385954
rect 312326 385398 312562 385634
rect 312646 385398 312882 385634
rect 312326 349718 312562 349954
rect 312646 349718 312882 349954
rect 312326 349398 312562 349634
rect 312646 349398 312882 349634
rect 312326 313718 312562 313954
rect 312646 313718 312882 313954
rect 312326 313398 312562 313634
rect 312646 313398 312882 313634
rect 312326 277718 312562 277954
rect 312646 277718 312882 277954
rect 312326 277398 312562 277634
rect 312646 277398 312882 277634
rect 312326 241718 312562 241954
rect 312646 241718 312882 241954
rect 312326 241398 312562 241634
rect 312646 241398 312882 241634
rect 312326 205718 312562 205954
rect 312646 205718 312882 205954
rect 312326 205398 312562 205634
rect 312646 205398 312882 205634
rect 312326 169718 312562 169954
rect 312646 169718 312882 169954
rect 312326 169398 312562 169634
rect 312646 169398 312882 169634
rect 312326 133718 312562 133954
rect 312646 133718 312882 133954
rect 312326 133398 312562 133634
rect 312646 133398 312882 133634
rect 312326 97718 312562 97954
rect 312646 97718 312882 97954
rect 312326 97398 312562 97634
rect 312646 97398 312882 97634
rect 312326 61718 312562 61954
rect 312646 61718 312882 61954
rect 312326 61398 312562 61634
rect 312646 61398 312882 61634
rect 312326 25718 312562 25954
rect 312646 25718 312882 25954
rect 312326 25398 312562 25634
rect 312646 25398 312882 25634
rect 312326 -5382 312562 -5146
rect 312646 -5382 312882 -5146
rect 312326 -5702 312562 -5466
rect 312646 -5702 312882 -5466
rect 316826 710362 317062 710598
rect 317146 710362 317382 710598
rect 316826 710042 317062 710278
rect 317146 710042 317382 710278
rect 316826 678218 317062 678454
rect 317146 678218 317382 678454
rect 316826 677898 317062 678134
rect 317146 677898 317382 678134
rect 316826 642218 317062 642454
rect 317146 642218 317382 642454
rect 316826 641898 317062 642134
rect 317146 641898 317382 642134
rect 316826 606218 317062 606454
rect 317146 606218 317382 606454
rect 316826 605898 317062 606134
rect 317146 605898 317382 606134
rect 316826 570218 317062 570454
rect 317146 570218 317382 570454
rect 316826 569898 317062 570134
rect 317146 569898 317382 570134
rect 316826 534218 317062 534454
rect 317146 534218 317382 534454
rect 316826 533898 317062 534134
rect 317146 533898 317382 534134
rect 316826 498218 317062 498454
rect 317146 498218 317382 498454
rect 316826 497898 317062 498134
rect 317146 497898 317382 498134
rect 316826 462218 317062 462454
rect 317146 462218 317382 462454
rect 316826 461898 317062 462134
rect 317146 461898 317382 462134
rect 316826 426218 317062 426454
rect 317146 426218 317382 426454
rect 316826 425898 317062 426134
rect 317146 425898 317382 426134
rect 316826 390218 317062 390454
rect 317146 390218 317382 390454
rect 316826 389898 317062 390134
rect 317146 389898 317382 390134
rect 316826 354218 317062 354454
rect 317146 354218 317382 354454
rect 316826 353898 317062 354134
rect 317146 353898 317382 354134
rect 316826 318218 317062 318454
rect 317146 318218 317382 318454
rect 316826 317898 317062 318134
rect 317146 317898 317382 318134
rect 316826 282218 317062 282454
rect 317146 282218 317382 282454
rect 316826 281898 317062 282134
rect 317146 281898 317382 282134
rect 316826 246218 317062 246454
rect 317146 246218 317382 246454
rect 316826 245898 317062 246134
rect 317146 245898 317382 246134
rect 316826 210218 317062 210454
rect 317146 210218 317382 210454
rect 316826 209898 317062 210134
rect 317146 209898 317382 210134
rect 316826 174218 317062 174454
rect 317146 174218 317382 174454
rect 316826 173898 317062 174134
rect 317146 173898 317382 174134
rect 316826 138218 317062 138454
rect 317146 138218 317382 138454
rect 316826 137898 317062 138134
rect 317146 137898 317382 138134
rect 316826 102218 317062 102454
rect 317146 102218 317382 102454
rect 316826 101898 317062 102134
rect 317146 101898 317382 102134
rect 316826 66218 317062 66454
rect 317146 66218 317382 66454
rect 316826 65898 317062 66134
rect 317146 65898 317382 66134
rect 316826 30218 317062 30454
rect 317146 30218 317382 30454
rect 316826 29898 317062 30134
rect 317146 29898 317382 30134
rect 316826 -6342 317062 -6106
rect 317146 -6342 317382 -6106
rect 316826 -6662 317062 -6426
rect 317146 -6662 317382 -6426
rect 321326 711322 321562 711558
rect 321646 711322 321882 711558
rect 321326 711002 321562 711238
rect 321646 711002 321882 711238
rect 321326 682718 321562 682954
rect 321646 682718 321882 682954
rect 321326 682398 321562 682634
rect 321646 682398 321882 682634
rect 321326 646718 321562 646954
rect 321646 646718 321882 646954
rect 321326 646398 321562 646634
rect 321646 646398 321882 646634
rect 321326 610718 321562 610954
rect 321646 610718 321882 610954
rect 321326 610398 321562 610634
rect 321646 610398 321882 610634
rect 321326 574718 321562 574954
rect 321646 574718 321882 574954
rect 321326 574398 321562 574634
rect 321646 574398 321882 574634
rect 321326 538718 321562 538954
rect 321646 538718 321882 538954
rect 321326 538398 321562 538634
rect 321646 538398 321882 538634
rect 321326 502718 321562 502954
rect 321646 502718 321882 502954
rect 321326 502398 321562 502634
rect 321646 502398 321882 502634
rect 321326 466718 321562 466954
rect 321646 466718 321882 466954
rect 321326 466398 321562 466634
rect 321646 466398 321882 466634
rect 321326 430718 321562 430954
rect 321646 430718 321882 430954
rect 321326 430398 321562 430634
rect 321646 430398 321882 430634
rect 321326 394718 321562 394954
rect 321646 394718 321882 394954
rect 321326 394398 321562 394634
rect 321646 394398 321882 394634
rect 321326 358718 321562 358954
rect 321646 358718 321882 358954
rect 321326 358398 321562 358634
rect 321646 358398 321882 358634
rect 321326 322718 321562 322954
rect 321646 322718 321882 322954
rect 321326 322398 321562 322634
rect 321646 322398 321882 322634
rect 321326 286718 321562 286954
rect 321646 286718 321882 286954
rect 321326 286398 321562 286634
rect 321646 286398 321882 286634
rect 321326 250718 321562 250954
rect 321646 250718 321882 250954
rect 321326 250398 321562 250634
rect 321646 250398 321882 250634
rect 321326 214718 321562 214954
rect 321646 214718 321882 214954
rect 321326 214398 321562 214634
rect 321646 214398 321882 214634
rect 321326 178718 321562 178954
rect 321646 178718 321882 178954
rect 321326 178398 321562 178634
rect 321646 178398 321882 178634
rect 321326 142718 321562 142954
rect 321646 142718 321882 142954
rect 321326 142398 321562 142634
rect 321646 142398 321882 142634
rect 321326 106718 321562 106954
rect 321646 106718 321882 106954
rect 321326 106398 321562 106634
rect 321646 106398 321882 106634
rect 321326 70718 321562 70954
rect 321646 70718 321882 70954
rect 321326 70398 321562 70634
rect 321646 70398 321882 70634
rect 321326 34718 321562 34954
rect 321646 34718 321882 34954
rect 321326 34398 321562 34634
rect 321646 34398 321882 34634
rect 321326 -7302 321562 -7066
rect 321646 -7302 321882 -7066
rect 321326 -7622 321562 -7386
rect 321646 -7622 321882 -7386
rect 325826 704602 326062 704838
rect 326146 704602 326382 704838
rect 325826 704282 326062 704518
rect 326146 704282 326382 704518
rect 325826 687218 326062 687454
rect 326146 687218 326382 687454
rect 325826 686898 326062 687134
rect 326146 686898 326382 687134
rect 325826 651218 326062 651454
rect 326146 651218 326382 651454
rect 325826 650898 326062 651134
rect 326146 650898 326382 651134
rect 325826 615218 326062 615454
rect 326146 615218 326382 615454
rect 325826 614898 326062 615134
rect 326146 614898 326382 615134
rect 325826 579218 326062 579454
rect 326146 579218 326382 579454
rect 325826 578898 326062 579134
rect 326146 578898 326382 579134
rect 325826 543218 326062 543454
rect 326146 543218 326382 543454
rect 325826 542898 326062 543134
rect 326146 542898 326382 543134
rect 325826 507218 326062 507454
rect 326146 507218 326382 507454
rect 325826 506898 326062 507134
rect 326146 506898 326382 507134
rect 325826 471218 326062 471454
rect 326146 471218 326382 471454
rect 325826 470898 326062 471134
rect 326146 470898 326382 471134
rect 325826 435218 326062 435454
rect 326146 435218 326382 435454
rect 325826 434898 326062 435134
rect 326146 434898 326382 435134
rect 325826 399218 326062 399454
rect 326146 399218 326382 399454
rect 325826 398898 326062 399134
rect 326146 398898 326382 399134
rect 325826 363218 326062 363454
rect 326146 363218 326382 363454
rect 325826 362898 326062 363134
rect 326146 362898 326382 363134
rect 325826 327218 326062 327454
rect 326146 327218 326382 327454
rect 325826 326898 326062 327134
rect 326146 326898 326382 327134
rect 325826 291218 326062 291454
rect 326146 291218 326382 291454
rect 325826 290898 326062 291134
rect 326146 290898 326382 291134
rect 325826 255218 326062 255454
rect 326146 255218 326382 255454
rect 325826 254898 326062 255134
rect 326146 254898 326382 255134
rect 325826 219218 326062 219454
rect 326146 219218 326382 219454
rect 325826 218898 326062 219134
rect 326146 218898 326382 219134
rect 325826 183218 326062 183454
rect 326146 183218 326382 183454
rect 325826 182898 326062 183134
rect 326146 182898 326382 183134
rect 325826 147218 326062 147454
rect 326146 147218 326382 147454
rect 325826 146898 326062 147134
rect 326146 146898 326382 147134
rect 325826 111218 326062 111454
rect 326146 111218 326382 111454
rect 325826 110898 326062 111134
rect 326146 110898 326382 111134
rect 325826 75218 326062 75454
rect 326146 75218 326382 75454
rect 325826 74898 326062 75134
rect 326146 74898 326382 75134
rect 325826 39218 326062 39454
rect 326146 39218 326382 39454
rect 325826 38898 326062 39134
rect 326146 38898 326382 39134
rect 325826 3218 326062 3454
rect 326146 3218 326382 3454
rect 325826 2898 326062 3134
rect 326146 2898 326382 3134
rect 325826 -582 326062 -346
rect 326146 -582 326382 -346
rect 325826 -902 326062 -666
rect 326146 -902 326382 -666
rect 330326 705562 330562 705798
rect 330646 705562 330882 705798
rect 330326 705242 330562 705478
rect 330646 705242 330882 705478
rect 330326 691718 330562 691954
rect 330646 691718 330882 691954
rect 330326 691398 330562 691634
rect 330646 691398 330882 691634
rect 330326 655718 330562 655954
rect 330646 655718 330882 655954
rect 330326 655398 330562 655634
rect 330646 655398 330882 655634
rect 330326 619718 330562 619954
rect 330646 619718 330882 619954
rect 330326 619398 330562 619634
rect 330646 619398 330882 619634
rect 330326 583718 330562 583954
rect 330646 583718 330882 583954
rect 330326 583398 330562 583634
rect 330646 583398 330882 583634
rect 330326 547718 330562 547954
rect 330646 547718 330882 547954
rect 330326 547398 330562 547634
rect 330646 547398 330882 547634
rect 330326 511718 330562 511954
rect 330646 511718 330882 511954
rect 330326 511398 330562 511634
rect 330646 511398 330882 511634
rect 330326 475718 330562 475954
rect 330646 475718 330882 475954
rect 330326 475398 330562 475634
rect 330646 475398 330882 475634
rect 330326 439718 330562 439954
rect 330646 439718 330882 439954
rect 330326 439398 330562 439634
rect 330646 439398 330882 439634
rect 330326 403718 330562 403954
rect 330646 403718 330882 403954
rect 330326 403398 330562 403634
rect 330646 403398 330882 403634
rect 330326 367718 330562 367954
rect 330646 367718 330882 367954
rect 330326 367398 330562 367634
rect 330646 367398 330882 367634
rect 330326 331718 330562 331954
rect 330646 331718 330882 331954
rect 330326 331398 330562 331634
rect 330646 331398 330882 331634
rect 330326 295718 330562 295954
rect 330646 295718 330882 295954
rect 330326 295398 330562 295634
rect 330646 295398 330882 295634
rect 330326 259718 330562 259954
rect 330646 259718 330882 259954
rect 330326 259398 330562 259634
rect 330646 259398 330882 259634
rect 330326 223718 330562 223954
rect 330646 223718 330882 223954
rect 330326 223398 330562 223634
rect 330646 223398 330882 223634
rect 330326 187718 330562 187954
rect 330646 187718 330882 187954
rect 330326 187398 330562 187634
rect 330646 187398 330882 187634
rect 330326 151718 330562 151954
rect 330646 151718 330882 151954
rect 330326 151398 330562 151634
rect 330646 151398 330882 151634
rect 330326 115718 330562 115954
rect 330646 115718 330882 115954
rect 330326 115398 330562 115634
rect 330646 115398 330882 115634
rect 330326 79718 330562 79954
rect 330646 79718 330882 79954
rect 330326 79398 330562 79634
rect 330646 79398 330882 79634
rect 330326 43718 330562 43954
rect 330646 43718 330882 43954
rect 330326 43398 330562 43634
rect 330646 43398 330882 43634
rect 330326 7718 330562 7954
rect 330646 7718 330882 7954
rect 330326 7398 330562 7634
rect 330646 7398 330882 7634
rect 330326 -1542 330562 -1306
rect 330646 -1542 330882 -1306
rect 330326 -1862 330562 -1626
rect 330646 -1862 330882 -1626
rect 334826 706522 335062 706758
rect 335146 706522 335382 706758
rect 334826 706202 335062 706438
rect 335146 706202 335382 706438
rect 334826 696218 335062 696454
rect 335146 696218 335382 696454
rect 334826 695898 335062 696134
rect 335146 695898 335382 696134
rect 334826 660218 335062 660454
rect 335146 660218 335382 660454
rect 334826 659898 335062 660134
rect 335146 659898 335382 660134
rect 334826 624218 335062 624454
rect 335146 624218 335382 624454
rect 334826 623898 335062 624134
rect 335146 623898 335382 624134
rect 334826 588218 335062 588454
rect 335146 588218 335382 588454
rect 334826 587898 335062 588134
rect 335146 587898 335382 588134
rect 334826 552218 335062 552454
rect 335146 552218 335382 552454
rect 334826 551898 335062 552134
rect 335146 551898 335382 552134
rect 334826 516218 335062 516454
rect 335146 516218 335382 516454
rect 334826 515898 335062 516134
rect 335146 515898 335382 516134
rect 334826 480218 335062 480454
rect 335146 480218 335382 480454
rect 334826 479898 335062 480134
rect 335146 479898 335382 480134
rect 334826 444218 335062 444454
rect 335146 444218 335382 444454
rect 334826 443898 335062 444134
rect 335146 443898 335382 444134
rect 334826 408218 335062 408454
rect 335146 408218 335382 408454
rect 334826 407898 335062 408134
rect 335146 407898 335382 408134
rect 334826 372218 335062 372454
rect 335146 372218 335382 372454
rect 334826 371898 335062 372134
rect 335146 371898 335382 372134
rect 334826 336218 335062 336454
rect 335146 336218 335382 336454
rect 334826 335898 335062 336134
rect 335146 335898 335382 336134
rect 334826 300218 335062 300454
rect 335146 300218 335382 300454
rect 334826 299898 335062 300134
rect 335146 299898 335382 300134
rect 334826 264218 335062 264454
rect 335146 264218 335382 264454
rect 334826 263898 335062 264134
rect 335146 263898 335382 264134
rect 334826 228218 335062 228454
rect 335146 228218 335382 228454
rect 334826 227898 335062 228134
rect 335146 227898 335382 228134
rect 334826 192218 335062 192454
rect 335146 192218 335382 192454
rect 334826 191898 335062 192134
rect 335146 191898 335382 192134
rect 334826 156218 335062 156454
rect 335146 156218 335382 156454
rect 334826 155898 335062 156134
rect 335146 155898 335382 156134
rect 334826 120218 335062 120454
rect 335146 120218 335382 120454
rect 334826 119898 335062 120134
rect 335146 119898 335382 120134
rect 334826 84218 335062 84454
rect 335146 84218 335382 84454
rect 334826 83898 335062 84134
rect 335146 83898 335382 84134
rect 334826 48218 335062 48454
rect 335146 48218 335382 48454
rect 334826 47898 335062 48134
rect 335146 47898 335382 48134
rect 334826 12218 335062 12454
rect 335146 12218 335382 12454
rect 334826 11898 335062 12134
rect 335146 11898 335382 12134
rect 334826 -2502 335062 -2266
rect 335146 -2502 335382 -2266
rect 334826 -2822 335062 -2586
rect 335146 -2822 335382 -2586
rect 339326 707482 339562 707718
rect 339646 707482 339882 707718
rect 339326 707162 339562 707398
rect 339646 707162 339882 707398
rect 339326 700718 339562 700954
rect 339646 700718 339882 700954
rect 339326 700398 339562 700634
rect 339646 700398 339882 700634
rect 339326 664718 339562 664954
rect 339646 664718 339882 664954
rect 339326 664398 339562 664634
rect 339646 664398 339882 664634
rect 339326 628718 339562 628954
rect 339646 628718 339882 628954
rect 339326 628398 339562 628634
rect 339646 628398 339882 628634
rect 339326 592718 339562 592954
rect 339646 592718 339882 592954
rect 339326 592398 339562 592634
rect 339646 592398 339882 592634
rect 339326 556718 339562 556954
rect 339646 556718 339882 556954
rect 339326 556398 339562 556634
rect 339646 556398 339882 556634
rect 339326 520718 339562 520954
rect 339646 520718 339882 520954
rect 339326 520398 339562 520634
rect 339646 520398 339882 520634
rect 339326 484718 339562 484954
rect 339646 484718 339882 484954
rect 339326 484398 339562 484634
rect 339646 484398 339882 484634
rect 339326 448718 339562 448954
rect 339646 448718 339882 448954
rect 339326 448398 339562 448634
rect 339646 448398 339882 448634
rect 339326 412718 339562 412954
rect 339646 412718 339882 412954
rect 339326 412398 339562 412634
rect 339646 412398 339882 412634
rect 339326 376718 339562 376954
rect 339646 376718 339882 376954
rect 339326 376398 339562 376634
rect 339646 376398 339882 376634
rect 339326 340718 339562 340954
rect 339646 340718 339882 340954
rect 339326 340398 339562 340634
rect 339646 340398 339882 340634
rect 339326 304718 339562 304954
rect 339646 304718 339882 304954
rect 339326 304398 339562 304634
rect 339646 304398 339882 304634
rect 339326 268718 339562 268954
rect 339646 268718 339882 268954
rect 339326 268398 339562 268634
rect 339646 268398 339882 268634
rect 339326 232718 339562 232954
rect 339646 232718 339882 232954
rect 339326 232398 339562 232634
rect 339646 232398 339882 232634
rect 339326 196718 339562 196954
rect 339646 196718 339882 196954
rect 339326 196398 339562 196634
rect 339646 196398 339882 196634
rect 339326 160718 339562 160954
rect 339646 160718 339882 160954
rect 339326 160398 339562 160634
rect 339646 160398 339882 160634
rect 339326 124718 339562 124954
rect 339646 124718 339882 124954
rect 339326 124398 339562 124634
rect 339646 124398 339882 124634
rect 339326 88718 339562 88954
rect 339646 88718 339882 88954
rect 339326 88398 339562 88634
rect 339646 88398 339882 88634
rect 339326 52718 339562 52954
rect 339646 52718 339882 52954
rect 339326 52398 339562 52634
rect 339646 52398 339882 52634
rect 339326 16718 339562 16954
rect 339646 16718 339882 16954
rect 339326 16398 339562 16634
rect 339646 16398 339882 16634
rect 339326 -3462 339562 -3226
rect 339646 -3462 339882 -3226
rect 339326 -3782 339562 -3546
rect 339646 -3782 339882 -3546
rect 343826 708442 344062 708678
rect 344146 708442 344382 708678
rect 343826 708122 344062 708358
rect 344146 708122 344382 708358
rect 343826 669218 344062 669454
rect 344146 669218 344382 669454
rect 343826 668898 344062 669134
rect 344146 668898 344382 669134
rect 343826 633218 344062 633454
rect 344146 633218 344382 633454
rect 343826 632898 344062 633134
rect 344146 632898 344382 633134
rect 343826 597218 344062 597454
rect 344146 597218 344382 597454
rect 343826 596898 344062 597134
rect 344146 596898 344382 597134
rect 343826 561218 344062 561454
rect 344146 561218 344382 561454
rect 343826 560898 344062 561134
rect 344146 560898 344382 561134
rect 343826 525218 344062 525454
rect 344146 525218 344382 525454
rect 343826 524898 344062 525134
rect 344146 524898 344382 525134
rect 343826 489218 344062 489454
rect 344146 489218 344382 489454
rect 343826 488898 344062 489134
rect 344146 488898 344382 489134
rect 343826 453218 344062 453454
rect 344146 453218 344382 453454
rect 343826 452898 344062 453134
rect 344146 452898 344382 453134
rect 343826 417218 344062 417454
rect 344146 417218 344382 417454
rect 343826 416898 344062 417134
rect 344146 416898 344382 417134
rect 343826 381218 344062 381454
rect 344146 381218 344382 381454
rect 343826 380898 344062 381134
rect 344146 380898 344382 381134
rect 343826 345218 344062 345454
rect 344146 345218 344382 345454
rect 343826 344898 344062 345134
rect 344146 344898 344382 345134
rect 343826 309218 344062 309454
rect 344146 309218 344382 309454
rect 343826 308898 344062 309134
rect 344146 308898 344382 309134
rect 343826 273218 344062 273454
rect 344146 273218 344382 273454
rect 343826 272898 344062 273134
rect 344146 272898 344382 273134
rect 343826 237218 344062 237454
rect 344146 237218 344382 237454
rect 343826 236898 344062 237134
rect 344146 236898 344382 237134
rect 343826 201218 344062 201454
rect 344146 201218 344382 201454
rect 343826 200898 344062 201134
rect 344146 200898 344382 201134
rect 343826 165218 344062 165454
rect 344146 165218 344382 165454
rect 343826 164898 344062 165134
rect 344146 164898 344382 165134
rect 343826 129218 344062 129454
rect 344146 129218 344382 129454
rect 343826 128898 344062 129134
rect 344146 128898 344382 129134
rect 343826 93218 344062 93454
rect 344146 93218 344382 93454
rect 343826 92898 344062 93134
rect 344146 92898 344382 93134
rect 343826 57218 344062 57454
rect 344146 57218 344382 57454
rect 343826 56898 344062 57134
rect 344146 56898 344382 57134
rect 343826 21218 344062 21454
rect 344146 21218 344382 21454
rect 343826 20898 344062 21134
rect 344146 20898 344382 21134
rect 343826 -4422 344062 -4186
rect 344146 -4422 344382 -4186
rect 343826 -4742 344062 -4506
rect 344146 -4742 344382 -4506
rect 348326 709402 348562 709638
rect 348646 709402 348882 709638
rect 348326 709082 348562 709318
rect 348646 709082 348882 709318
rect 348326 673718 348562 673954
rect 348646 673718 348882 673954
rect 348326 673398 348562 673634
rect 348646 673398 348882 673634
rect 348326 637718 348562 637954
rect 348646 637718 348882 637954
rect 348326 637398 348562 637634
rect 348646 637398 348882 637634
rect 348326 601718 348562 601954
rect 348646 601718 348882 601954
rect 348326 601398 348562 601634
rect 348646 601398 348882 601634
rect 348326 565718 348562 565954
rect 348646 565718 348882 565954
rect 348326 565398 348562 565634
rect 348646 565398 348882 565634
rect 348326 529718 348562 529954
rect 348646 529718 348882 529954
rect 348326 529398 348562 529634
rect 348646 529398 348882 529634
rect 348326 493718 348562 493954
rect 348646 493718 348882 493954
rect 348326 493398 348562 493634
rect 348646 493398 348882 493634
rect 348326 457718 348562 457954
rect 348646 457718 348882 457954
rect 348326 457398 348562 457634
rect 348646 457398 348882 457634
rect 348326 421718 348562 421954
rect 348646 421718 348882 421954
rect 348326 421398 348562 421634
rect 348646 421398 348882 421634
rect 348326 385718 348562 385954
rect 348646 385718 348882 385954
rect 348326 385398 348562 385634
rect 348646 385398 348882 385634
rect 348326 349718 348562 349954
rect 348646 349718 348882 349954
rect 348326 349398 348562 349634
rect 348646 349398 348882 349634
rect 348326 313718 348562 313954
rect 348646 313718 348882 313954
rect 348326 313398 348562 313634
rect 348646 313398 348882 313634
rect 348326 277718 348562 277954
rect 348646 277718 348882 277954
rect 348326 277398 348562 277634
rect 348646 277398 348882 277634
rect 348326 241718 348562 241954
rect 348646 241718 348882 241954
rect 348326 241398 348562 241634
rect 348646 241398 348882 241634
rect 348326 205718 348562 205954
rect 348646 205718 348882 205954
rect 348326 205398 348562 205634
rect 348646 205398 348882 205634
rect 348326 169718 348562 169954
rect 348646 169718 348882 169954
rect 348326 169398 348562 169634
rect 348646 169398 348882 169634
rect 348326 133718 348562 133954
rect 348646 133718 348882 133954
rect 348326 133398 348562 133634
rect 348646 133398 348882 133634
rect 348326 97718 348562 97954
rect 348646 97718 348882 97954
rect 348326 97398 348562 97634
rect 348646 97398 348882 97634
rect 348326 61718 348562 61954
rect 348646 61718 348882 61954
rect 348326 61398 348562 61634
rect 348646 61398 348882 61634
rect 348326 25718 348562 25954
rect 348646 25718 348882 25954
rect 348326 25398 348562 25634
rect 348646 25398 348882 25634
rect 348326 -5382 348562 -5146
rect 348646 -5382 348882 -5146
rect 348326 -5702 348562 -5466
rect 348646 -5702 348882 -5466
rect 352826 710362 353062 710598
rect 353146 710362 353382 710598
rect 352826 710042 353062 710278
rect 353146 710042 353382 710278
rect 352826 678218 353062 678454
rect 353146 678218 353382 678454
rect 352826 677898 353062 678134
rect 353146 677898 353382 678134
rect 352826 642218 353062 642454
rect 353146 642218 353382 642454
rect 352826 641898 353062 642134
rect 353146 641898 353382 642134
rect 352826 606218 353062 606454
rect 353146 606218 353382 606454
rect 352826 605898 353062 606134
rect 353146 605898 353382 606134
rect 352826 570218 353062 570454
rect 353146 570218 353382 570454
rect 352826 569898 353062 570134
rect 353146 569898 353382 570134
rect 352826 534218 353062 534454
rect 353146 534218 353382 534454
rect 352826 533898 353062 534134
rect 353146 533898 353382 534134
rect 352826 498218 353062 498454
rect 353146 498218 353382 498454
rect 352826 497898 353062 498134
rect 353146 497898 353382 498134
rect 352826 462218 353062 462454
rect 353146 462218 353382 462454
rect 352826 461898 353062 462134
rect 353146 461898 353382 462134
rect 352826 426218 353062 426454
rect 353146 426218 353382 426454
rect 352826 425898 353062 426134
rect 353146 425898 353382 426134
rect 352826 390218 353062 390454
rect 353146 390218 353382 390454
rect 352826 389898 353062 390134
rect 353146 389898 353382 390134
rect 352826 354218 353062 354454
rect 353146 354218 353382 354454
rect 352826 353898 353062 354134
rect 353146 353898 353382 354134
rect 352826 318218 353062 318454
rect 353146 318218 353382 318454
rect 352826 317898 353062 318134
rect 353146 317898 353382 318134
rect 352826 282218 353062 282454
rect 353146 282218 353382 282454
rect 352826 281898 353062 282134
rect 353146 281898 353382 282134
rect 352826 246218 353062 246454
rect 353146 246218 353382 246454
rect 352826 245898 353062 246134
rect 353146 245898 353382 246134
rect 352826 210218 353062 210454
rect 353146 210218 353382 210454
rect 352826 209898 353062 210134
rect 353146 209898 353382 210134
rect 352826 174218 353062 174454
rect 353146 174218 353382 174454
rect 352826 173898 353062 174134
rect 353146 173898 353382 174134
rect 352826 138218 353062 138454
rect 353146 138218 353382 138454
rect 352826 137898 353062 138134
rect 353146 137898 353382 138134
rect 352826 102218 353062 102454
rect 353146 102218 353382 102454
rect 352826 101898 353062 102134
rect 353146 101898 353382 102134
rect 352826 66218 353062 66454
rect 353146 66218 353382 66454
rect 352826 65898 353062 66134
rect 353146 65898 353382 66134
rect 352826 30218 353062 30454
rect 353146 30218 353382 30454
rect 352826 29898 353062 30134
rect 353146 29898 353382 30134
rect 352826 -6342 353062 -6106
rect 353146 -6342 353382 -6106
rect 352826 -6662 353062 -6426
rect 353146 -6662 353382 -6426
rect 357326 711322 357562 711558
rect 357646 711322 357882 711558
rect 357326 711002 357562 711238
rect 357646 711002 357882 711238
rect 357326 682718 357562 682954
rect 357646 682718 357882 682954
rect 357326 682398 357562 682634
rect 357646 682398 357882 682634
rect 357326 646718 357562 646954
rect 357646 646718 357882 646954
rect 357326 646398 357562 646634
rect 357646 646398 357882 646634
rect 357326 610718 357562 610954
rect 357646 610718 357882 610954
rect 357326 610398 357562 610634
rect 357646 610398 357882 610634
rect 357326 574718 357562 574954
rect 357646 574718 357882 574954
rect 357326 574398 357562 574634
rect 357646 574398 357882 574634
rect 357326 538718 357562 538954
rect 357646 538718 357882 538954
rect 357326 538398 357562 538634
rect 357646 538398 357882 538634
rect 357326 502718 357562 502954
rect 357646 502718 357882 502954
rect 357326 502398 357562 502634
rect 357646 502398 357882 502634
rect 357326 466718 357562 466954
rect 357646 466718 357882 466954
rect 357326 466398 357562 466634
rect 357646 466398 357882 466634
rect 357326 430718 357562 430954
rect 357646 430718 357882 430954
rect 357326 430398 357562 430634
rect 357646 430398 357882 430634
rect 357326 394718 357562 394954
rect 357646 394718 357882 394954
rect 357326 394398 357562 394634
rect 357646 394398 357882 394634
rect 357326 358718 357562 358954
rect 357646 358718 357882 358954
rect 357326 358398 357562 358634
rect 357646 358398 357882 358634
rect 357326 322718 357562 322954
rect 357646 322718 357882 322954
rect 357326 322398 357562 322634
rect 357646 322398 357882 322634
rect 357326 286718 357562 286954
rect 357646 286718 357882 286954
rect 357326 286398 357562 286634
rect 357646 286398 357882 286634
rect 357326 250718 357562 250954
rect 357646 250718 357882 250954
rect 357326 250398 357562 250634
rect 357646 250398 357882 250634
rect 357326 214718 357562 214954
rect 357646 214718 357882 214954
rect 357326 214398 357562 214634
rect 357646 214398 357882 214634
rect 357326 178718 357562 178954
rect 357646 178718 357882 178954
rect 357326 178398 357562 178634
rect 357646 178398 357882 178634
rect 357326 142718 357562 142954
rect 357646 142718 357882 142954
rect 357326 142398 357562 142634
rect 357646 142398 357882 142634
rect 357326 106718 357562 106954
rect 357646 106718 357882 106954
rect 357326 106398 357562 106634
rect 357646 106398 357882 106634
rect 357326 70718 357562 70954
rect 357646 70718 357882 70954
rect 357326 70398 357562 70634
rect 357646 70398 357882 70634
rect 357326 34718 357562 34954
rect 357646 34718 357882 34954
rect 357326 34398 357562 34634
rect 357646 34398 357882 34634
rect 357326 -7302 357562 -7066
rect 357646 -7302 357882 -7066
rect 357326 -7622 357562 -7386
rect 357646 -7622 357882 -7386
rect 361826 704602 362062 704838
rect 362146 704602 362382 704838
rect 361826 704282 362062 704518
rect 362146 704282 362382 704518
rect 361826 687218 362062 687454
rect 362146 687218 362382 687454
rect 361826 686898 362062 687134
rect 362146 686898 362382 687134
rect 361826 651218 362062 651454
rect 362146 651218 362382 651454
rect 361826 650898 362062 651134
rect 362146 650898 362382 651134
rect 361826 615218 362062 615454
rect 362146 615218 362382 615454
rect 361826 614898 362062 615134
rect 362146 614898 362382 615134
rect 361826 579218 362062 579454
rect 362146 579218 362382 579454
rect 361826 578898 362062 579134
rect 362146 578898 362382 579134
rect 361826 543218 362062 543454
rect 362146 543218 362382 543454
rect 361826 542898 362062 543134
rect 362146 542898 362382 543134
rect 361826 507218 362062 507454
rect 362146 507218 362382 507454
rect 361826 506898 362062 507134
rect 362146 506898 362382 507134
rect 361826 471218 362062 471454
rect 362146 471218 362382 471454
rect 361826 470898 362062 471134
rect 362146 470898 362382 471134
rect 361826 435218 362062 435454
rect 362146 435218 362382 435454
rect 361826 434898 362062 435134
rect 362146 434898 362382 435134
rect 361826 399218 362062 399454
rect 362146 399218 362382 399454
rect 361826 398898 362062 399134
rect 362146 398898 362382 399134
rect 361826 363218 362062 363454
rect 362146 363218 362382 363454
rect 361826 362898 362062 363134
rect 362146 362898 362382 363134
rect 361826 327218 362062 327454
rect 362146 327218 362382 327454
rect 361826 326898 362062 327134
rect 362146 326898 362382 327134
rect 361826 291218 362062 291454
rect 362146 291218 362382 291454
rect 361826 290898 362062 291134
rect 362146 290898 362382 291134
rect 361826 255218 362062 255454
rect 362146 255218 362382 255454
rect 361826 254898 362062 255134
rect 362146 254898 362382 255134
rect 361826 219218 362062 219454
rect 362146 219218 362382 219454
rect 361826 218898 362062 219134
rect 362146 218898 362382 219134
rect 361826 183218 362062 183454
rect 362146 183218 362382 183454
rect 361826 182898 362062 183134
rect 362146 182898 362382 183134
rect 361826 147218 362062 147454
rect 362146 147218 362382 147454
rect 361826 146898 362062 147134
rect 362146 146898 362382 147134
rect 361826 111218 362062 111454
rect 362146 111218 362382 111454
rect 361826 110898 362062 111134
rect 362146 110898 362382 111134
rect 361826 75218 362062 75454
rect 362146 75218 362382 75454
rect 361826 74898 362062 75134
rect 362146 74898 362382 75134
rect 361826 39218 362062 39454
rect 362146 39218 362382 39454
rect 361826 38898 362062 39134
rect 362146 38898 362382 39134
rect 361826 3218 362062 3454
rect 362146 3218 362382 3454
rect 361826 2898 362062 3134
rect 362146 2898 362382 3134
rect 361826 -582 362062 -346
rect 362146 -582 362382 -346
rect 361826 -902 362062 -666
rect 362146 -902 362382 -666
rect 366326 705562 366562 705798
rect 366646 705562 366882 705798
rect 366326 705242 366562 705478
rect 366646 705242 366882 705478
rect 366326 691718 366562 691954
rect 366646 691718 366882 691954
rect 366326 691398 366562 691634
rect 366646 691398 366882 691634
rect 366326 655718 366562 655954
rect 366646 655718 366882 655954
rect 366326 655398 366562 655634
rect 366646 655398 366882 655634
rect 366326 619718 366562 619954
rect 366646 619718 366882 619954
rect 366326 619398 366562 619634
rect 366646 619398 366882 619634
rect 366326 583718 366562 583954
rect 366646 583718 366882 583954
rect 366326 583398 366562 583634
rect 366646 583398 366882 583634
rect 366326 547718 366562 547954
rect 366646 547718 366882 547954
rect 366326 547398 366562 547634
rect 366646 547398 366882 547634
rect 366326 511718 366562 511954
rect 366646 511718 366882 511954
rect 366326 511398 366562 511634
rect 366646 511398 366882 511634
rect 366326 475718 366562 475954
rect 366646 475718 366882 475954
rect 366326 475398 366562 475634
rect 366646 475398 366882 475634
rect 366326 439718 366562 439954
rect 366646 439718 366882 439954
rect 366326 439398 366562 439634
rect 366646 439398 366882 439634
rect 366326 403718 366562 403954
rect 366646 403718 366882 403954
rect 366326 403398 366562 403634
rect 366646 403398 366882 403634
rect 366326 367718 366562 367954
rect 366646 367718 366882 367954
rect 366326 367398 366562 367634
rect 366646 367398 366882 367634
rect 366326 331718 366562 331954
rect 366646 331718 366882 331954
rect 366326 331398 366562 331634
rect 366646 331398 366882 331634
rect 366326 295718 366562 295954
rect 366646 295718 366882 295954
rect 366326 295398 366562 295634
rect 366646 295398 366882 295634
rect 366326 259718 366562 259954
rect 366646 259718 366882 259954
rect 366326 259398 366562 259634
rect 366646 259398 366882 259634
rect 366326 223718 366562 223954
rect 366646 223718 366882 223954
rect 366326 223398 366562 223634
rect 366646 223398 366882 223634
rect 366326 187718 366562 187954
rect 366646 187718 366882 187954
rect 366326 187398 366562 187634
rect 366646 187398 366882 187634
rect 366326 151718 366562 151954
rect 366646 151718 366882 151954
rect 366326 151398 366562 151634
rect 366646 151398 366882 151634
rect 366326 115718 366562 115954
rect 366646 115718 366882 115954
rect 366326 115398 366562 115634
rect 366646 115398 366882 115634
rect 366326 79718 366562 79954
rect 366646 79718 366882 79954
rect 366326 79398 366562 79634
rect 366646 79398 366882 79634
rect 366326 43718 366562 43954
rect 366646 43718 366882 43954
rect 366326 43398 366562 43634
rect 366646 43398 366882 43634
rect 366326 7718 366562 7954
rect 366646 7718 366882 7954
rect 366326 7398 366562 7634
rect 366646 7398 366882 7634
rect 366326 -1542 366562 -1306
rect 366646 -1542 366882 -1306
rect 366326 -1862 366562 -1626
rect 366646 -1862 366882 -1626
rect 370826 706522 371062 706758
rect 371146 706522 371382 706758
rect 370826 706202 371062 706438
rect 371146 706202 371382 706438
rect 370826 696218 371062 696454
rect 371146 696218 371382 696454
rect 370826 695898 371062 696134
rect 371146 695898 371382 696134
rect 370826 660218 371062 660454
rect 371146 660218 371382 660454
rect 370826 659898 371062 660134
rect 371146 659898 371382 660134
rect 370826 624218 371062 624454
rect 371146 624218 371382 624454
rect 370826 623898 371062 624134
rect 371146 623898 371382 624134
rect 370826 588218 371062 588454
rect 371146 588218 371382 588454
rect 370826 587898 371062 588134
rect 371146 587898 371382 588134
rect 370826 552218 371062 552454
rect 371146 552218 371382 552454
rect 370826 551898 371062 552134
rect 371146 551898 371382 552134
rect 370826 516218 371062 516454
rect 371146 516218 371382 516454
rect 370826 515898 371062 516134
rect 371146 515898 371382 516134
rect 370826 480218 371062 480454
rect 371146 480218 371382 480454
rect 370826 479898 371062 480134
rect 371146 479898 371382 480134
rect 370826 444218 371062 444454
rect 371146 444218 371382 444454
rect 370826 443898 371062 444134
rect 371146 443898 371382 444134
rect 370826 408218 371062 408454
rect 371146 408218 371382 408454
rect 370826 407898 371062 408134
rect 371146 407898 371382 408134
rect 370826 372218 371062 372454
rect 371146 372218 371382 372454
rect 370826 371898 371062 372134
rect 371146 371898 371382 372134
rect 370826 336218 371062 336454
rect 371146 336218 371382 336454
rect 370826 335898 371062 336134
rect 371146 335898 371382 336134
rect 370826 300218 371062 300454
rect 371146 300218 371382 300454
rect 370826 299898 371062 300134
rect 371146 299898 371382 300134
rect 370826 264218 371062 264454
rect 371146 264218 371382 264454
rect 370826 263898 371062 264134
rect 371146 263898 371382 264134
rect 370826 228218 371062 228454
rect 371146 228218 371382 228454
rect 370826 227898 371062 228134
rect 371146 227898 371382 228134
rect 370826 192218 371062 192454
rect 371146 192218 371382 192454
rect 370826 191898 371062 192134
rect 371146 191898 371382 192134
rect 370826 156218 371062 156454
rect 371146 156218 371382 156454
rect 370826 155898 371062 156134
rect 371146 155898 371382 156134
rect 370826 120218 371062 120454
rect 371146 120218 371382 120454
rect 370826 119898 371062 120134
rect 371146 119898 371382 120134
rect 370826 84218 371062 84454
rect 371146 84218 371382 84454
rect 370826 83898 371062 84134
rect 371146 83898 371382 84134
rect 370826 48218 371062 48454
rect 371146 48218 371382 48454
rect 370826 47898 371062 48134
rect 371146 47898 371382 48134
rect 370826 12218 371062 12454
rect 371146 12218 371382 12454
rect 370826 11898 371062 12134
rect 371146 11898 371382 12134
rect 370826 -2502 371062 -2266
rect 371146 -2502 371382 -2266
rect 370826 -2822 371062 -2586
rect 371146 -2822 371382 -2586
rect 375326 707482 375562 707718
rect 375646 707482 375882 707718
rect 375326 707162 375562 707398
rect 375646 707162 375882 707398
rect 375326 700718 375562 700954
rect 375646 700718 375882 700954
rect 375326 700398 375562 700634
rect 375646 700398 375882 700634
rect 375326 664718 375562 664954
rect 375646 664718 375882 664954
rect 375326 664398 375562 664634
rect 375646 664398 375882 664634
rect 375326 628718 375562 628954
rect 375646 628718 375882 628954
rect 375326 628398 375562 628634
rect 375646 628398 375882 628634
rect 375326 592718 375562 592954
rect 375646 592718 375882 592954
rect 375326 592398 375562 592634
rect 375646 592398 375882 592634
rect 375326 556718 375562 556954
rect 375646 556718 375882 556954
rect 375326 556398 375562 556634
rect 375646 556398 375882 556634
rect 375326 520718 375562 520954
rect 375646 520718 375882 520954
rect 375326 520398 375562 520634
rect 375646 520398 375882 520634
rect 375326 484718 375562 484954
rect 375646 484718 375882 484954
rect 375326 484398 375562 484634
rect 375646 484398 375882 484634
rect 375326 448718 375562 448954
rect 375646 448718 375882 448954
rect 375326 448398 375562 448634
rect 375646 448398 375882 448634
rect 375326 412718 375562 412954
rect 375646 412718 375882 412954
rect 375326 412398 375562 412634
rect 375646 412398 375882 412634
rect 375326 376718 375562 376954
rect 375646 376718 375882 376954
rect 375326 376398 375562 376634
rect 375646 376398 375882 376634
rect 375326 340718 375562 340954
rect 375646 340718 375882 340954
rect 375326 340398 375562 340634
rect 375646 340398 375882 340634
rect 375326 304718 375562 304954
rect 375646 304718 375882 304954
rect 375326 304398 375562 304634
rect 375646 304398 375882 304634
rect 375326 268718 375562 268954
rect 375646 268718 375882 268954
rect 375326 268398 375562 268634
rect 375646 268398 375882 268634
rect 375326 232718 375562 232954
rect 375646 232718 375882 232954
rect 375326 232398 375562 232634
rect 375646 232398 375882 232634
rect 375326 196718 375562 196954
rect 375646 196718 375882 196954
rect 375326 196398 375562 196634
rect 375646 196398 375882 196634
rect 375326 160718 375562 160954
rect 375646 160718 375882 160954
rect 375326 160398 375562 160634
rect 375646 160398 375882 160634
rect 375326 124718 375562 124954
rect 375646 124718 375882 124954
rect 375326 124398 375562 124634
rect 375646 124398 375882 124634
rect 375326 88718 375562 88954
rect 375646 88718 375882 88954
rect 375326 88398 375562 88634
rect 375646 88398 375882 88634
rect 375326 52718 375562 52954
rect 375646 52718 375882 52954
rect 375326 52398 375562 52634
rect 375646 52398 375882 52634
rect 375326 16718 375562 16954
rect 375646 16718 375882 16954
rect 375326 16398 375562 16634
rect 375646 16398 375882 16634
rect 375326 -3462 375562 -3226
rect 375646 -3462 375882 -3226
rect 375326 -3782 375562 -3546
rect 375646 -3782 375882 -3546
rect 379826 708442 380062 708678
rect 380146 708442 380382 708678
rect 379826 708122 380062 708358
rect 380146 708122 380382 708358
rect 379826 669218 380062 669454
rect 380146 669218 380382 669454
rect 379826 668898 380062 669134
rect 380146 668898 380382 669134
rect 379826 633218 380062 633454
rect 380146 633218 380382 633454
rect 379826 632898 380062 633134
rect 380146 632898 380382 633134
rect 379826 597218 380062 597454
rect 380146 597218 380382 597454
rect 379826 596898 380062 597134
rect 380146 596898 380382 597134
rect 379826 561218 380062 561454
rect 380146 561218 380382 561454
rect 379826 560898 380062 561134
rect 380146 560898 380382 561134
rect 379826 525218 380062 525454
rect 380146 525218 380382 525454
rect 379826 524898 380062 525134
rect 380146 524898 380382 525134
rect 379826 489218 380062 489454
rect 380146 489218 380382 489454
rect 379826 488898 380062 489134
rect 380146 488898 380382 489134
rect 379826 453218 380062 453454
rect 380146 453218 380382 453454
rect 379826 452898 380062 453134
rect 380146 452898 380382 453134
rect 379826 417218 380062 417454
rect 380146 417218 380382 417454
rect 379826 416898 380062 417134
rect 380146 416898 380382 417134
rect 379826 381218 380062 381454
rect 380146 381218 380382 381454
rect 379826 380898 380062 381134
rect 380146 380898 380382 381134
rect 379826 345218 380062 345454
rect 380146 345218 380382 345454
rect 379826 344898 380062 345134
rect 380146 344898 380382 345134
rect 379826 309218 380062 309454
rect 380146 309218 380382 309454
rect 379826 308898 380062 309134
rect 380146 308898 380382 309134
rect 379826 273218 380062 273454
rect 380146 273218 380382 273454
rect 379826 272898 380062 273134
rect 380146 272898 380382 273134
rect 379826 237218 380062 237454
rect 380146 237218 380382 237454
rect 379826 236898 380062 237134
rect 380146 236898 380382 237134
rect 379826 201218 380062 201454
rect 380146 201218 380382 201454
rect 379826 200898 380062 201134
rect 380146 200898 380382 201134
rect 379826 165218 380062 165454
rect 380146 165218 380382 165454
rect 379826 164898 380062 165134
rect 380146 164898 380382 165134
rect 379826 129218 380062 129454
rect 380146 129218 380382 129454
rect 379826 128898 380062 129134
rect 380146 128898 380382 129134
rect 379826 93218 380062 93454
rect 380146 93218 380382 93454
rect 379826 92898 380062 93134
rect 380146 92898 380382 93134
rect 379826 57218 380062 57454
rect 380146 57218 380382 57454
rect 379826 56898 380062 57134
rect 380146 56898 380382 57134
rect 379826 21218 380062 21454
rect 380146 21218 380382 21454
rect 379826 20898 380062 21134
rect 380146 20898 380382 21134
rect 379826 -4422 380062 -4186
rect 380146 -4422 380382 -4186
rect 379826 -4742 380062 -4506
rect 380146 -4742 380382 -4506
rect 384326 709402 384562 709638
rect 384646 709402 384882 709638
rect 384326 709082 384562 709318
rect 384646 709082 384882 709318
rect 384326 673718 384562 673954
rect 384646 673718 384882 673954
rect 384326 673398 384562 673634
rect 384646 673398 384882 673634
rect 384326 637718 384562 637954
rect 384646 637718 384882 637954
rect 384326 637398 384562 637634
rect 384646 637398 384882 637634
rect 384326 601718 384562 601954
rect 384646 601718 384882 601954
rect 384326 601398 384562 601634
rect 384646 601398 384882 601634
rect 384326 565718 384562 565954
rect 384646 565718 384882 565954
rect 384326 565398 384562 565634
rect 384646 565398 384882 565634
rect 384326 529718 384562 529954
rect 384646 529718 384882 529954
rect 384326 529398 384562 529634
rect 384646 529398 384882 529634
rect 384326 493718 384562 493954
rect 384646 493718 384882 493954
rect 384326 493398 384562 493634
rect 384646 493398 384882 493634
rect 384326 457718 384562 457954
rect 384646 457718 384882 457954
rect 384326 457398 384562 457634
rect 384646 457398 384882 457634
rect 384326 421718 384562 421954
rect 384646 421718 384882 421954
rect 384326 421398 384562 421634
rect 384646 421398 384882 421634
rect 384326 385718 384562 385954
rect 384646 385718 384882 385954
rect 384326 385398 384562 385634
rect 384646 385398 384882 385634
rect 384326 349718 384562 349954
rect 384646 349718 384882 349954
rect 384326 349398 384562 349634
rect 384646 349398 384882 349634
rect 384326 313718 384562 313954
rect 384646 313718 384882 313954
rect 384326 313398 384562 313634
rect 384646 313398 384882 313634
rect 384326 277718 384562 277954
rect 384646 277718 384882 277954
rect 384326 277398 384562 277634
rect 384646 277398 384882 277634
rect 384326 241718 384562 241954
rect 384646 241718 384882 241954
rect 384326 241398 384562 241634
rect 384646 241398 384882 241634
rect 384326 205718 384562 205954
rect 384646 205718 384882 205954
rect 384326 205398 384562 205634
rect 384646 205398 384882 205634
rect 384326 169718 384562 169954
rect 384646 169718 384882 169954
rect 384326 169398 384562 169634
rect 384646 169398 384882 169634
rect 384326 133718 384562 133954
rect 384646 133718 384882 133954
rect 384326 133398 384562 133634
rect 384646 133398 384882 133634
rect 384326 97718 384562 97954
rect 384646 97718 384882 97954
rect 384326 97398 384562 97634
rect 384646 97398 384882 97634
rect 384326 61718 384562 61954
rect 384646 61718 384882 61954
rect 384326 61398 384562 61634
rect 384646 61398 384882 61634
rect 384326 25718 384562 25954
rect 384646 25718 384882 25954
rect 384326 25398 384562 25634
rect 384646 25398 384882 25634
rect 384326 -5382 384562 -5146
rect 384646 -5382 384882 -5146
rect 384326 -5702 384562 -5466
rect 384646 -5702 384882 -5466
rect 388826 710362 389062 710598
rect 389146 710362 389382 710598
rect 388826 710042 389062 710278
rect 389146 710042 389382 710278
rect 388826 678218 389062 678454
rect 389146 678218 389382 678454
rect 388826 677898 389062 678134
rect 389146 677898 389382 678134
rect 388826 642218 389062 642454
rect 389146 642218 389382 642454
rect 388826 641898 389062 642134
rect 389146 641898 389382 642134
rect 388826 606218 389062 606454
rect 389146 606218 389382 606454
rect 388826 605898 389062 606134
rect 389146 605898 389382 606134
rect 388826 570218 389062 570454
rect 389146 570218 389382 570454
rect 388826 569898 389062 570134
rect 389146 569898 389382 570134
rect 388826 534218 389062 534454
rect 389146 534218 389382 534454
rect 388826 533898 389062 534134
rect 389146 533898 389382 534134
rect 388826 498218 389062 498454
rect 389146 498218 389382 498454
rect 388826 497898 389062 498134
rect 389146 497898 389382 498134
rect 388826 462218 389062 462454
rect 389146 462218 389382 462454
rect 388826 461898 389062 462134
rect 389146 461898 389382 462134
rect 388826 426218 389062 426454
rect 389146 426218 389382 426454
rect 388826 425898 389062 426134
rect 389146 425898 389382 426134
rect 388826 390218 389062 390454
rect 389146 390218 389382 390454
rect 388826 389898 389062 390134
rect 389146 389898 389382 390134
rect 388826 354218 389062 354454
rect 389146 354218 389382 354454
rect 388826 353898 389062 354134
rect 389146 353898 389382 354134
rect 388826 318218 389062 318454
rect 389146 318218 389382 318454
rect 388826 317898 389062 318134
rect 389146 317898 389382 318134
rect 388826 282218 389062 282454
rect 389146 282218 389382 282454
rect 388826 281898 389062 282134
rect 389146 281898 389382 282134
rect 388826 246218 389062 246454
rect 389146 246218 389382 246454
rect 388826 245898 389062 246134
rect 389146 245898 389382 246134
rect 388826 210218 389062 210454
rect 389146 210218 389382 210454
rect 388826 209898 389062 210134
rect 389146 209898 389382 210134
rect 388826 174218 389062 174454
rect 389146 174218 389382 174454
rect 388826 173898 389062 174134
rect 389146 173898 389382 174134
rect 388826 138218 389062 138454
rect 389146 138218 389382 138454
rect 388826 137898 389062 138134
rect 389146 137898 389382 138134
rect 388826 102218 389062 102454
rect 389146 102218 389382 102454
rect 388826 101898 389062 102134
rect 389146 101898 389382 102134
rect 388826 66218 389062 66454
rect 389146 66218 389382 66454
rect 388826 65898 389062 66134
rect 389146 65898 389382 66134
rect 388826 30218 389062 30454
rect 389146 30218 389382 30454
rect 388826 29898 389062 30134
rect 389146 29898 389382 30134
rect 388826 -6342 389062 -6106
rect 389146 -6342 389382 -6106
rect 388826 -6662 389062 -6426
rect 389146 -6662 389382 -6426
rect 393326 711322 393562 711558
rect 393646 711322 393882 711558
rect 393326 711002 393562 711238
rect 393646 711002 393882 711238
rect 393326 682718 393562 682954
rect 393646 682718 393882 682954
rect 393326 682398 393562 682634
rect 393646 682398 393882 682634
rect 393326 646718 393562 646954
rect 393646 646718 393882 646954
rect 393326 646398 393562 646634
rect 393646 646398 393882 646634
rect 393326 610718 393562 610954
rect 393646 610718 393882 610954
rect 393326 610398 393562 610634
rect 393646 610398 393882 610634
rect 393326 574718 393562 574954
rect 393646 574718 393882 574954
rect 393326 574398 393562 574634
rect 393646 574398 393882 574634
rect 393326 538718 393562 538954
rect 393646 538718 393882 538954
rect 393326 538398 393562 538634
rect 393646 538398 393882 538634
rect 393326 502718 393562 502954
rect 393646 502718 393882 502954
rect 393326 502398 393562 502634
rect 393646 502398 393882 502634
rect 393326 466718 393562 466954
rect 393646 466718 393882 466954
rect 393326 466398 393562 466634
rect 393646 466398 393882 466634
rect 393326 430718 393562 430954
rect 393646 430718 393882 430954
rect 393326 430398 393562 430634
rect 393646 430398 393882 430634
rect 393326 394718 393562 394954
rect 393646 394718 393882 394954
rect 393326 394398 393562 394634
rect 393646 394398 393882 394634
rect 393326 358718 393562 358954
rect 393646 358718 393882 358954
rect 393326 358398 393562 358634
rect 393646 358398 393882 358634
rect 393326 322718 393562 322954
rect 393646 322718 393882 322954
rect 393326 322398 393562 322634
rect 393646 322398 393882 322634
rect 393326 286718 393562 286954
rect 393646 286718 393882 286954
rect 393326 286398 393562 286634
rect 393646 286398 393882 286634
rect 393326 250718 393562 250954
rect 393646 250718 393882 250954
rect 393326 250398 393562 250634
rect 393646 250398 393882 250634
rect 393326 214718 393562 214954
rect 393646 214718 393882 214954
rect 393326 214398 393562 214634
rect 393646 214398 393882 214634
rect 393326 178718 393562 178954
rect 393646 178718 393882 178954
rect 393326 178398 393562 178634
rect 393646 178398 393882 178634
rect 393326 142718 393562 142954
rect 393646 142718 393882 142954
rect 393326 142398 393562 142634
rect 393646 142398 393882 142634
rect 393326 106718 393562 106954
rect 393646 106718 393882 106954
rect 393326 106398 393562 106634
rect 393646 106398 393882 106634
rect 393326 70718 393562 70954
rect 393646 70718 393882 70954
rect 393326 70398 393562 70634
rect 393646 70398 393882 70634
rect 393326 34718 393562 34954
rect 393646 34718 393882 34954
rect 393326 34398 393562 34634
rect 393646 34398 393882 34634
rect 393326 -7302 393562 -7066
rect 393646 -7302 393882 -7066
rect 393326 -7622 393562 -7386
rect 393646 -7622 393882 -7386
rect 397826 704602 398062 704838
rect 398146 704602 398382 704838
rect 397826 704282 398062 704518
rect 398146 704282 398382 704518
rect 397826 687218 398062 687454
rect 398146 687218 398382 687454
rect 397826 686898 398062 687134
rect 398146 686898 398382 687134
rect 397826 651218 398062 651454
rect 398146 651218 398382 651454
rect 397826 650898 398062 651134
rect 398146 650898 398382 651134
rect 397826 615218 398062 615454
rect 398146 615218 398382 615454
rect 397826 614898 398062 615134
rect 398146 614898 398382 615134
rect 397826 579218 398062 579454
rect 398146 579218 398382 579454
rect 397826 578898 398062 579134
rect 398146 578898 398382 579134
rect 397826 543218 398062 543454
rect 398146 543218 398382 543454
rect 397826 542898 398062 543134
rect 398146 542898 398382 543134
rect 397826 507218 398062 507454
rect 398146 507218 398382 507454
rect 397826 506898 398062 507134
rect 398146 506898 398382 507134
rect 397826 471218 398062 471454
rect 398146 471218 398382 471454
rect 397826 470898 398062 471134
rect 398146 470898 398382 471134
rect 397826 435218 398062 435454
rect 398146 435218 398382 435454
rect 397826 434898 398062 435134
rect 398146 434898 398382 435134
rect 397826 399218 398062 399454
rect 398146 399218 398382 399454
rect 397826 398898 398062 399134
rect 398146 398898 398382 399134
rect 397826 363218 398062 363454
rect 398146 363218 398382 363454
rect 397826 362898 398062 363134
rect 398146 362898 398382 363134
rect 397826 327218 398062 327454
rect 398146 327218 398382 327454
rect 397826 326898 398062 327134
rect 398146 326898 398382 327134
rect 397826 291218 398062 291454
rect 398146 291218 398382 291454
rect 397826 290898 398062 291134
rect 398146 290898 398382 291134
rect 397826 255218 398062 255454
rect 398146 255218 398382 255454
rect 397826 254898 398062 255134
rect 398146 254898 398382 255134
rect 397826 219218 398062 219454
rect 398146 219218 398382 219454
rect 397826 218898 398062 219134
rect 398146 218898 398382 219134
rect 397826 183218 398062 183454
rect 398146 183218 398382 183454
rect 397826 182898 398062 183134
rect 398146 182898 398382 183134
rect 397826 147218 398062 147454
rect 398146 147218 398382 147454
rect 397826 146898 398062 147134
rect 398146 146898 398382 147134
rect 397826 111218 398062 111454
rect 398146 111218 398382 111454
rect 397826 110898 398062 111134
rect 398146 110898 398382 111134
rect 397826 75218 398062 75454
rect 398146 75218 398382 75454
rect 397826 74898 398062 75134
rect 398146 74898 398382 75134
rect 397826 39218 398062 39454
rect 398146 39218 398382 39454
rect 397826 38898 398062 39134
rect 398146 38898 398382 39134
rect 397826 3218 398062 3454
rect 398146 3218 398382 3454
rect 397826 2898 398062 3134
rect 398146 2898 398382 3134
rect 397826 -582 398062 -346
rect 398146 -582 398382 -346
rect 397826 -902 398062 -666
rect 398146 -902 398382 -666
rect 402326 705562 402562 705798
rect 402646 705562 402882 705798
rect 402326 705242 402562 705478
rect 402646 705242 402882 705478
rect 402326 691718 402562 691954
rect 402646 691718 402882 691954
rect 402326 691398 402562 691634
rect 402646 691398 402882 691634
rect 402326 655718 402562 655954
rect 402646 655718 402882 655954
rect 402326 655398 402562 655634
rect 402646 655398 402882 655634
rect 402326 619718 402562 619954
rect 402646 619718 402882 619954
rect 402326 619398 402562 619634
rect 402646 619398 402882 619634
rect 402326 583718 402562 583954
rect 402646 583718 402882 583954
rect 402326 583398 402562 583634
rect 402646 583398 402882 583634
rect 402326 547718 402562 547954
rect 402646 547718 402882 547954
rect 402326 547398 402562 547634
rect 402646 547398 402882 547634
rect 402326 511718 402562 511954
rect 402646 511718 402882 511954
rect 402326 511398 402562 511634
rect 402646 511398 402882 511634
rect 402326 475718 402562 475954
rect 402646 475718 402882 475954
rect 402326 475398 402562 475634
rect 402646 475398 402882 475634
rect 402326 439718 402562 439954
rect 402646 439718 402882 439954
rect 402326 439398 402562 439634
rect 402646 439398 402882 439634
rect 402326 403718 402562 403954
rect 402646 403718 402882 403954
rect 402326 403398 402562 403634
rect 402646 403398 402882 403634
rect 402326 367718 402562 367954
rect 402646 367718 402882 367954
rect 402326 367398 402562 367634
rect 402646 367398 402882 367634
rect 402326 331718 402562 331954
rect 402646 331718 402882 331954
rect 402326 331398 402562 331634
rect 402646 331398 402882 331634
rect 402326 295718 402562 295954
rect 402646 295718 402882 295954
rect 402326 295398 402562 295634
rect 402646 295398 402882 295634
rect 402326 259718 402562 259954
rect 402646 259718 402882 259954
rect 402326 259398 402562 259634
rect 402646 259398 402882 259634
rect 402326 223718 402562 223954
rect 402646 223718 402882 223954
rect 402326 223398 402562 223634
rect 402646 223398 402882 223634
rect 402326 187718 402562 187954
rect 402646 187718 402882 187954
rect 402326 187398 402562 187634
rect 402646 187398 402882 187634
rect 402326 151718 402562 151954
rect 402646 151718 402882 151954
rect 402326 151398 402562 151634
rect 402646 151398 402882 151634
rect 402326 115718 402562 115954
rect 402646 115718 402882 115954
rect 402326 115398 402562 115634
rect 402646 115398 402882 115634
rect 402326 79718 402562 79954
rect 402646 79718 402882 79954
rect 402326 79398 402562 79634
rect 402646 79398 402882 79634
rect 402326 43718 402562 43954
rect 402646 43718 402882 43954
rect 402326 43398 402562 43634
rect 402646 43398 402882 43634
rect 402326 7718 402562 7954
rect 402646 7718 402882 7954
rect 402326 7398 402562 7634
rect 402646 7398 402882 7634
rect 402326 -1542 402562 -1306
rect 402646 -1542 402882 -1306
rect 402326 -1862 402562 -1626
rect 402646 -1862 402882 -1626
rect 406826 706522 407062 706758
rect 407146 706522 407382 706758
rect 406826 706202 407062 706438
rect 407146 706202 407382 706438
rect 406826 696218 407062 696454
rect 407146 696218 407382 696454
rect 406826 695898 407062 696134
rect 407146 695898 407382 696134
rect 406826 660218 407062 660454
rect 407146 660218 407382 660454
rect 406826 659898 407062 660134
rect 407146 659898 407382 660134
rect 406826 624218 407062 624454
rect 407146 624218 407382 624454
rect 406826 623898 407062 624134
rect 407146 623898 407382 624134
rect 406826 588218 407062 588454
rect 407146 588218 407382 588454
rect 406826 587898 407062 588134
rect 407146 587898 407382 588134
rect 406826 552218 407062 552454
rect 407146 552218 407382 552454
rect 406826 551898 407062 552134
rect 407146 551898 407382 552134
rect 406826 516218 407062 516454
rect 407146 516218 407382 516454
rect 406826 515898 407062 516134
rect 407146 515898 407382 516134
rect 406826 480218 407062 480454
rect 407146 480218 407382 480454
rect 406826 479898 407062 480134
rect 407146 479898 407382 480134
rect 406826 444218 407062 444454
rect 407146 444218 407382 444454
rect 406826 443898 407062 444134
rect 407146 443898 407382 444134
rect 406826 408218 407062 408454
rect 407146 408218 407382 408454
rect 406826 407898 407062 408134
rect 407146 407898 407382 408134
rect 406826 372218 407062 372454
rect 407146 372218 407382 372454
rect 406826 371898 407062 372134
rect 407146 371898 407382 372134
rect 406826 336218 407062 336454
rect 407146 336218 407382 336454
rect 406826 335898 407062 336134
rect 407146 335898 407382 336134
rect 406826 300218 407062 300454
rect 407146 300218 407382 300454
rect 406826 299898 407062 300134
rect 407146 299898 407382 300134
rect 406826 264218 407062 264454
rect 407146 264218 407382 264454
rect 406826 263898 407062 264134
rect 407146 263898 407382 264134
rect 406826 228218 407062 228454
rect 407146 228218 407382 228454
rect 406826 227898 407062 228134
rect 407146 227898 407382 228134
rect 406826 192218 407062 192454
rect 407146 192218 407382 192454
rect 406826 191898 407062 192134
rect 407146 191898 407382 192134
rect 406826 156218 407062 156454
rect 407146 156218 407382 156454
rect 406826 155898 407062 156134
rect 407146 155898 407382 156134
rect 406826 120218 407062 120454
rect 407146 120218 407382 120454
rect 406826 119898 407062 120134
rect 407146 119898 407382 120134
rect 406826 84218 407062 84454
rect 407146 84218 407382 84454
rect 406826 83898 407062 84134
rect 407146 83898 407382 84134
rect 406826 48218 407062 48454
rect 407146 48218 407382 48454
rect 406826 47898 407062 48134
rect 407146 47898 407382 48134
rect 406826 12218 407062 12454
rect 407146 12218 407382 12454
rect 406826 11898 407062 12134
rect 407146 11898 407382 12134
rect 406826 -2502 407062 -2266
rect 407146 -2502 407382 -2266
rect 406826 -2822 407062 -2586
rect 407146 -2822 407382 -2586
rect 411326 707482 411562 707718
rect 411646 707482 411882 707718
rect 411326 707162 411562 707398
rect 411646 707162 411882 707398
rect 411326 700718 411562 700954
rect 411646 700718 411882 700954
rect 411326 700398 411562 700634
rect 411646 700398 411882 700634
rect 411326 664718 411562 664954
rect 411646 664718 411882 664954
rect 411326 664398 411562 664634
rect 411646 664398 411882 664634
rect 411326 628718 411562 628954
rect 411646 628718 411882 628954
rect 411326 628398 411562 628634
rect 411646 628398 411882 628634
rect 411326 592718 411562 592954
rect 411646 592718 411882 592954
rect 411326 592398 411562 592634
rect 411646 592398 411882 592634
rect 411326 556718 411562 556954
rect 411646 556718 411882 556954
rect 411326 556398 411562 556634
rect 411646 556398 411882 556634
rect 411326 520718 411562 520954
rect 411646 520718 411882 520954
rect 411326 520398 411562 520634
rect 411646 520398 411882 520634
rect 411326 484718 411562 484954
rect 411646 484718 411882 484954
rect 411326 484398 411562 484634
rect 411646 484398 411882 484634
rect 411326 448718 411562 448954
rect 411646 448718 411882 448954
rect 411326 448398 411562 448634
rect 411646 448398 411882 448634
rect 411326 412718 411562 412954
rect 411646 412718 411882 412954
rect 411326 412398 411562 412634
rect 411646 412398 411882 412634
rect 411326 376718 411562 376954
rect 411646 376718 411882 376954
rect 411326 376398 411562 376634
rect 411646 376398 411882 376634
rect 411326 340718 411562 340954
rect 411646 340718 411882 340954
rect 411326 340398 411562 340634
rect 411646 340398 411882 340634
rect 411326 304718 411562 304954
rect 411646 304718 411882 304954
rect 411326 304398 411562 304634
rect 411646 304398 411882 304634
rect 411326 268718 411562 268954
rect 411646 268718 411882 268954
rect 411326 268398 411562 268634
rect 411646 268398 411882 268634
rect 411326 232718 411562 232954
rect 411646 232718 411882 232954
rect 411326 232398 411562 232634
rect 411646 232398 411882 232634
rect 411326 196718 411562 196954
rect 411646 196718 411882 196954
rect 411326 196398 411562 196634
rect 411646 196398 411882 196634
rect 411326 160718 411562 160954
rect 411646 160718 411882 160954
rect 411326 160398 411562 160634
rect 411646 160398 411882 160634
rect 411326 124718 411562 124954
rect 411646 124718 411882 124954
rect 411326 124398 411562 124634
rect 411646 124398 411882 124634
rect 411326 88718 411562 88954
rect 411646 88718 411882 88954
rect 411326 88398 411562 88634
rect 411646 88398 411882 88634
rect 411326 52718 411562 52954
rect 411646 52718 411882 52954
rect 411326 52398 411562 52634
rect 411646 52398 411882 52634
rect 411326 16718 411562 16954
rect 411646 16718 411882 16954
rect 411326 16398 411562 16634
rect 411646 16398 411882 16634
rect 411326 -3462 411562 -3226
rect 411646 -3462 411882 -3226
rect 411326 -3782 411562 -3546
rect 411646 -3782 411882 -3546
rect 415826 708442 416062 708678
rect 416146 708442 416382 708678
rect 415826 708122 416062 708358
rect 416146 708122 416382 708358
rect 415826 669218 416062 669454
rect 416146 669218 416382 669454
rect 415826 668898 416062 669134
rect 416146 668898 416382 669134
rect 415826 633218 416062 633454
rect 416146 633218 416382 633454
rect 415826 632898 416062 633134
rect 416146 632898 416382 633134
rect 415826 597218 416062 597454
rect 416146 597218 416382 597454
rect 415826 596898 416062 597134
rect 416146 596898 416382 597134
rect 415826 561218 416062 561454
rect 416146 561218 416382 561454
rect 415826 560898 416062 561134
rect 416146 560898 416382 561134
rect 415826 525218 416062 525454
rect 416146 525218 416382 525454
rect 415826 524898 416062 525134
rect 416146 524898 416382 525134
rect 415826 489218 416062 489454
rect 416146 489218 416382 489454
rect 415826 488898 416062 489134
rect 416146 488898 416382 489134
rect 415826 453218 416062 453454
rect 416146 453218 416382 453454
rect 415826 452898 416062 453134
rect 416146 452898 416382 453134
rect 415826 417218 416062 417454
rect 416146 417218 416382 417454
rect 415826 416898 416062 417134
rect 416146 416898 416382 417134
rect 415826 381218 416062 381454
rect 416146 381218 416382 381454
rect 415826 380898 416062 381134
rect 416146 380898 416382 381134
rect 415826 345218 416062 345454
rect 416146 345218 416382 345454
rect 415826 344898 416062 345134
rect 416146 344898 416382 345134
rect 415826 309218 416062 309454
rect 416146 309218 416382 309454
rect 415826 308898 416062 309134
rect 416146 308898 416382 309134
rect 415826 273218 416062 273454
rect 416146 273218 416382 273454
rect 415826 272898 416062 273134
rect 416146 272898 416382 273134
rect 415826 237218 416062 237454
rect 416146 237218 416382 237454
rect 415826 236898 416062 237134
rect 416146 236898 416382 237134
rect 415826 201218 416062 201454
rect 416146 201218 416382 201454
rect 415826 200898 416062 201134
rect 416146 200898 416382 201134
rect 415826 165218 416062 165454
rect 416146 165218 416382 165454
rect 415826 164898 416062 165134
rect 416146 164898 416382 165134
rect 415826 129218 416062 129454
rect 416146 129218 416382 129454
rect 415826 128898 416062 129134
rect 416146 128898 416382 129134
rect 415826 93218 416062 93454
rect 416146 93218 416382 93454
rect 415826 92898 416062 93134
rect 416146 92898 416382 93134
rect 415826 57218 416062 57454
rect 416146 57218 416382 57454
rect 415826 56898 416062 57134
rect 416146 56898 416382 57134
rect 415826 21218 416062 21454
rect 416146 21218 416382 21454
rect 415826 20898 416062 21134
rect 416146 20898 416382 21134
rect 415826 -4422 416062 -4186
rect 416146 -4422 416382 -4186
rect 415826 -4742 416062 -4506
rect 416146 -4742 416382 -4506
rect 420326 709402 420562 709638
rect 420646 709402 420882 709638
rect 420326 709082 420562 709318
rect 420646 709082 420882 709318
rect 420326 673718 420562 673954
rect 420646 673718 420882 673954
rect 420326 673398 420562 673634
rect 420646 673398 420882 673634
rect 420326 637718 420562 637954
rect 420646 637718 420882 637954
rect 420326 637398 420562 637634
rect 420646 637398 420882 637634
rect 420326 601718 420562 601954
rect 420646 601718 420882 601954
rect 420326 601398 420562 601634
rect 420646 601398 420882 601634
rect 420326 565718 420562 565954
rect 420646 565718 420882 565954
rect 420326 565398 420562 565634
rect 420646 565398 420882 565634
rect 420326 529718 420562 529954
rect 420646 529718 420882 529954
rect 420326 529398 420562 529634
rect 420646 529398 420882 529634
rect 420326 493718 420562 493954
rect 420646 493718 420882 493954
rect 420326 493398 420562 493634
rect 420646 493398 420882 493634
rect 420326 457718 420562 457954
rect 420646 457718 420882 457954
rect 420326 457398 420562 457634
rect 420646 457398 420882 457634
rect 420326 421718 420562 421954
rect 420646 421718 420882 421954
rect 420326 421398 420562 421634
rect 420646 421398 420882 421634
rect 420326 385718 420562 385954
rect 420646 385718 420882 385954
rect 420326 385398 420562 385634
rect 420646 385398 420882 385634
rect 420326 349718 420562 349954
rect 420646 349718 420882 349954
rect 420326 349398 420562 349634
rect 420646 349398 420882 349634
rect 420326 313718 420562 313954
rect 420646 313718 420882 313954
rect 420326 313398 420562 313634
rect 420646 313398 420882 313634
rect 420326 277718 420562 277954
rect 420646 277718 420882 277954
rect 420326 277398 420562 277634
rect 420646 277398 420882 277634
rect 420326 241718 420562 241954
rect 420646 241718 420882 241954
rect 420326 241398 420562 241634
rect 420646 241398 420882 241634
rect 420326 205718 420562 205954
rect 420646 205718 420882 205954
rect 420326 205398 420562 205634
rect 420646 205398 420882 205634
rect 420326 169718 420562 169954
rect 420646 169718 420882 169954
rect 420326 169398 420562 169634
rect 420646 169398 420882 169634
rect 420326 133718 420562 133954
rect 420646 133718 420882 133954
rect 420326 133398 420562 133634
rect 420646 133398 420882 133634
rect 420326 97718 420562 97954
rect 420646 97718 420882 97954
rect 420326 97398 420562 97634
rect 420646 97398 420882 97634
rect 420326 61718 420562 61954
rect 420646 61718 420882 61954
rect 420326 61398 420562 61634
rect 420646 61398 420882 61634
rect 420326 25718 420562 25954
rect 420646 25718 420882 25954
rect 420326 25398 420562 25634
rect 420646 25398 420882 25634
rect 420326 -5382 420562 -5146
rect 420646 -5382 420882 -5146
rect 420326 -5702 420562 -5466
rect 420646 -5702 420882 -5466
rect 424826 710362 425062 710598
rect 425146 710362 425382 710598
rect 424826 710042 425062 710278
rect 425146 710042 425382 710278
rect 424826 678218 425062 678454
rect 425146 678218 425382 678454
rect 424826 677898 425062 678134
rect 425146 677898 425382 678134
rect 424826 642218 425062 642454
rect 425146 642218 425382 642454
rect 424826 641898 425062 642134
rect 425146 641898 425382 642134
rect 424826 606218 425062 606454
rect 425146 606218 425382 606454
rect 424826 605898 425062 606134
rect 425146 605898 425382 606134
rect 424826 570218 425062 570454
rect 425146 570218 425382 570454
rect 424826 569898 425062 570134
rect 425146 569898 425382 570134
rect 424826 534218 425062 534454
rect 425146 534218 425382 534454
rect 424826 533898 425062 534134
rect 425146 533898 425382 534134
rect 424826 498218 425062 498454
rect 425146 498218 425382 498454
rect 424826 497898 425062 498134
rect 425146 497898 425382 498134
rect 424826 462218 425062 462454
rect 425146 462218 425382 462454
rect 424826 461898 425062 462134
rect 425146 461898 425382 462134
rect 424826 426218 425062 426454
rect 425146 426218 425382 426454
rect 424826 425898 425062 426134
rect 425146 425898 425382 426134
rect 424826 390218 425062 390454
rect 425146 390218 425382 390454
rect 424826 389898 425062 390134
rect 425146 389898 425382 390134
rect 424826 354218 425062 354454
rect 425146 354218 425382 354454
rect 424826 353898 425062 354134
rect 425146 353898 425382 354134
rect 424826 318218 425062 318454
rect 425146 318218 425382 318454
rect 424826 317898 425062 318134
rect 425146 317898 425382 318134
rect 424826 282218 425062 282454
rect 425146 282218 425382 282454
rect 424826 281898 425062 282134
rect 425146 281898 425382 282134
rect 424826 246218 425062 246454
rect 425146 246218 425382 246454
rect 424826 245898 425062 246134
rect 425146 245898 425382 246134
rect 424826 210218 425062 210454
rect 425146 210218 425382 210454
rect 424826 209898 425062 210134
rect 425146 209898 425382 210134
rect 424826 174218 425062 174454
rect 425146 174218 425382 174454
rect 424826 173898 425062 174134
rect 425146 173898 425382 174134
rect 424826 138218 425062 138454
rect 425146 138218 425382 138454
rect 424826 137898 425062 138134
rect 425146 137898 425382 138134
rect 424826 102218 425062 102454
rect 425146 102218 425382 102454
rect 424826 101898 425062 102134
rect 425146 101898 425382 102134
rect 424826 66218 425062 66454
rect 425146 66218 425382 66454
rect 424826 65898 425062 66134
rect 425146 65898 425382 66134
rect 424826 30218 425062 30454
rect 425146 30218 425382 30454
rect 424826 29898 425062 30134
rect 425146 29898 425382 30134
rect 424826 -6342 425062 -6106
rect 425146 -6342 425382 -6106
rect 424826 -6662 425062 -6426
rect 425146 -6662 425382 -6426
rect 429326 711322 429562 711558
rect 429646 711322 429882 711558
rect 429326 711002 429562 711238
rect 429646 711002 429882 711238
rect 429326 682718 429562 682954
rect 429646 682718 429882 682954
rect 429326 682398 429562 682634
rect 429646 682398 429882 682634
rect 429326 646718 429562 646954
rect 429646 646718 429882 646954
rect 429326 646398 429562 646634
rect 429646 646398 429882 646634
rect 429326 610718 429562 610954
rect 429646 610718 429882 610954
rect 429326 610398 429562 610634
rect 429646 610398 429882 610634
rect 429326 574718 429562 574954
rect 429646 574718 429882 574954
rect 429326 574398 429562 574634
rect 429646 574398 429882 574634
rect 429326 538718 429562 538954
rect 429646 538718 429882 538954
rect 429326 538398 429562 538634
rect 429646 538398 429882 538634
rect 429326 502718 429562 502954
rect 429646 502718 429882 502954
rect 429326 502398 429562 502634
rect 429646 502398 429882 502634
rect 429326 466718 429562 466954
rect 429646 466718 429882 466954
rect 429326 466398 429562 466634
rect 429646 466398 429882 466634
rect 429326 430718 429562 430954
rect 429646 430718 429882 430954
rect 429326 430398 429562 430634
rect 429646 430398 429882 430634
rect 429326 394718 429562 394954
rect 429646 394718 429882 394954
rect 429326 394398 429562 394634
rect 429646 394398 429882 394634
rect 429326 358718 429562 358954
rect 429646 358718 429882 358954
rect 429326 358398 429562 358634
rect 429646 358398 429882 358634
rect 429326 322718 429562 322954
rect 429646 322718 429882 322954
rect 429326 322398 429562 322634
rect 429646 322398 429882 322634
rect 429326 286718 429562 286954
rect 429646 286718 429882 286954
rect 429326 286398 429562 286634
rect 429646 286398 429882 286634
rect 429326 250718 429562 250954
rect 429646 250718 429882 250954
rect 429326 250398 429562 250634
rect 429646 250398 429882 250634
rect 429326 214718 429562 214954
rect 429646 214718 429882 214954
rect 429326 214398 429562 214634
rect 429646 214398 429882 214634
rect 429326 178718 429562 178954
rect 429646 178718 429882 178954
rect 429326 178398 429562 178634
rect 429646 178398 429882 178634
rect 429326 142718 429562 142954
rect 429646 142718 429882 142954
rect 429326 142398 429562 142634
rect 429646 142398 429882 142634
rect 429326 106718 429562 106954
rect 429646 106718 429882 106954
rect 429326 106398 429562 106634
rect 429646 106398 429882 106634
rect 429326 70718 429562 70954
rect 429646 70718 429882 70954
rect 429326 70398 429562 70634
rect 429646 70398 429882 70634
rect 429326 34718 429562 34954
rect 429646 34718 429882 34954
rect 429326 34398 429562 34634
rect 429646 34398 429882 34634
rect 429326 -7302 429562 -7066
rect 429646 -7302 429882 -7066
rect 429326 -7622 429562 -7386
rect 429646 -7622 429882 -7386
rect 433826 704602 434062 704838
rect 434146 704602 434382 704838
rect 433826 704282 434062 704518
rect 434146 704282 434382 704518
rect 433826 687218 434062 687454
rect 434146 687218 434382 687454
rect 433826 686898 434062 687134
rect 434146 686898 434382 687134
rect 433826 651218 434062 651454
rect 434146 651218 434382 651454
rect 433826 650898 434062 651134
rect 434146 650898 434382 651134
rect 433826 615218 434062 615454
rect 434146 615218 434382 615454
rect 433826 614898 434062 615134
rect 434146 614898 434382 615134
rect 433826 579218 434062 579454
rect 434146 579218 434382 579454
rect 433826 578898 434062 579134
rect 434146 578898 434382 579134
rect 433826 543218 434062 543454
rect 434146 543218 434382 543454
rect 433826 542898 434062 543134
rect 434146 542898 434382 543134
rect 433826 507218 434062 507454
rect 434146 507218 434382 507454
rect 433826 506898 434062 507134
rect 434146 506898 434382 507134
rect 433826 471218 434062 471454
rect 434146 471218 434382 471454
rect 433826 470898 434062 471134
rect 434146 470898 434382 471134
rect 433826 435218 434062 435454
rect 434146 435218 434382 435454
rect 433826 434898 434062 435134
rect 434146 434898 434382 435134
rect 433826 399218 434062 399454
rect 434146 399218 434382 399454
rect 433826 398898 434062 399134
rect 434146 398898 434382 399134
rect 433826 363218 434062 363454
rect 434146 363218 434382 363454
rect 433826 362898 434062 363134
rect 434146 362898 434382 363134
rect 433826 327218 434062 327454
rect 434146 327218 434382 327454
rect 433826 326898 434062 327134
rect 434146 326898 434382 327134
rect 433826 291218 434062 291454
rect 434146 291218 434382 291454
rect 433826 290898 434062 291134
rect 434146 290898 434382 291134
rect 433826 255218 434062 255454
rect 434146 255218 434382 255454
rect 433826 254898 434062 255134
rect 434146 254898 434382 255134
rect 433826 219218 434062 219454
rect 434146 219218 434382 219454
rect 433826 218898 434062 219134
rect 434146 218898 434382 219134
rect 433826 183218 434062 183454
rect 434146 183218 434382 183454
rect 433826 182898 434062 183134
rect 434146 182898 434382 183134
rect 433826 147218 434062 147454
rect 434146 147218 434382 147454
rect 433826 146898 434062 147134
rect 434146 146898 434382 147134
rect 433826 111218 434062 111454
rect 434146 111218 434382 111454
rect 433826 110898 434062 111134
rect 434146 110898 434382 111134
rect 433826 75218 434062 75454
rect 434146 75218 434382 75454
rect 433826 74898 434062 75134
rect 434146 74898 434382 75134
rect 433826 39218 434062 39454
rect 434146 39218 434382 39454
rect 433826 38898 434062 39134
rect 434146 38898 434382 39134
rect 433826 3218 434062 3454
rect 434146 3218 434382 3454
rect 433826 2898 434062 3134
rect 434146 2898 434382 3134
rect 433826 -582 434062 -346
rect 434146 -582 434382 -346
rect 433826 -902 434062 -666
rect 434146 -902 434382 -666
rect 438326 705562 438562 705798
rect 438646 705562 438882 705798
rect 438326 705242 438562 705478
rect 438646 705242 438882 705478
rect 438326 691718 438562 691954
rect 438646 691718 438882 691954
rect 438326 691398 438562 691634
rect 438646 691398 438882 691634
rect 438326 655718 438562 655954
rect 438646 655718 438882 655954
rect 438326 655398 438562 655634
rect 438646 655398 438882 655634
rect 438326 619718 438562 619954
rect 438646 619718 438882 619954
rect 438326 619398 438562 619634
rect 438646 619398 438882 619634
rect 438326 583718 438562 583954
rect 438646 583718 438882 583954
rect 438326 583398 438562 583634
rect 438646 583398 438882 583634
rect 438326 547718 438562 547954
rect 438646 547718 438882 547954
rect 438326 547398 438562 547634
rect 438646 547398 438882 547634
rect 438326 511718 438562 511954
rect 438646 511718 438882 511954
rect 438326 511398 438562 511634
rect 438646 511398 438882 511634
rect 438326 475718 438562 475954
rect 438646 475718 438882 475954
rect 438326 475398 438562 475634
rect 438646 475398 438882 475634
rect 438326 439718 438562 439954
rect 438646 439718 438882 439954
rect 438326 439398 438562 439634
rect 438646 439398 438882 439634
rect 438326 403718 438562 403954
rect 438646 403718 438882 403954
rect 438326 403398 438562 403634
rect 438646 403398 438882 403634
rect 438326 367718 438562 367954
rect 438646 367718 438882 367954
rect 438326 367398 438562 367634
rect 438646 367398 438882 367634
rect 438326 331718 438562 331954
rect 438646 331718 438882 331954
rect 438326 331398 438562 331634
rect 438646 331398 438882 331634
rect 438326 295718 438562 295954
rect 438646 295718 438882 295954
rect 438326 295398 438562 295634
rect 438646 295398 438882 295634
rect 438326 259718 438562 259954
rect 438646 259718 438882 259954
rect 438326 259398 438562 259634
rect 438646 259398 438882 259634
rect 438326 223718 438562 223954
rect 438646 223718 438882 223954
rect 438326 223398 438562 223634
rect 438646 223398 438882 223634
rect 438326 187718 438562 187954
rect 438646 187718 438882 187954
rect 438326 187398 438562 187634
rect 438646 187398 438882 187634
rect 438326 151718 438562 151954
rect 438646 151718 438882 151954
rect 438326 151398 438562 151634
rect 438646 151398 438882 151634
rect 438326 115718 438562 115954
rect 438646 115718 438882 115954
rect 438326 115398 438562 115634
rect 438646 115398 438882 115634
rect 438326 79718 438562 79954
rect 438646 79718 438882 79954
rect 438326 79398 438562 79634
rect 438646 79398 438882 79634
rect 438326 43718 438562 43954
rect 438646 43718 438882 43954
rect 438326 43398 438562 43634
rect 438646 43398 438882 43634
rect 438326 7718 438562 7954
rect 438646 7718 438882 7954
rect 438326 7398 438562 7634
rect 438646 7398 438882 7634
rect 438326 -1542 438562 -1306
rect 438646 -1542 438882 -1306
rect 438326 -1862 438562 -1626
rect 438646 -1862 438882 -1626
rect 442826 706522 443062 706758
rect 443146 706522 443382 706758
rect 442826 706202 443062 706438
rect 443146 706202 443382 706438
rect 442826 696218 443062 696454
rect 443146 696218 443382 696454
rect 442826 695898 443062 696134
rect 443146 695898 443382 696134
rect 442826 660218 443062 660454
rect 443146 660218 443382 660454
rect 442826 659898 443062 660134
rect 443146 659898 443382 660134
rect 442826 624218 443062 624454
rect 443146 624218 443382 624454
rect 442826 623898 443062 624134
rect 443146 623898 443382 624134
rect 442826 588218 443062 588454
rect 443146 588218 443382 588454
rect 442826 587898 443062 588134
rect 443146 587898 443382 588134
rect 442826 552218 443062 552454
rect 443146 552218 443382 552454
rect 442826 551898 443062 552134
rect 443146 551898 443382 552134
rect 442826 516218 443062 516454
rect 443146 516218 443382 516454
rect 442826 515898 443062 516134
rect 443146 515898 443382 516134
rect 442826 480218 443062 480454
rect 443146 480218 443382 480454
rect 442826 479898 443062 480134
rect 443146 479898 443382 480134
rect 442826 444218 443062 444454
rect 443146 444218 443382 444454
rect 442826 443898 443062 444134
rect 443146 443898 443382 444134
rect 442826 408218 443062 408454
rect 443146 408218 443382 408454
rect 442826 407898 443062 408134
rect 443146 407898 443382 408134
rect 442826 372218 443062 372454
rect 443146 372218 443382 372454
rect 442826 371898 443062 372134
rect 443146 371898 443382 372134
rect 442826 336218 443062 336454
rect 443146 336218 443382 336454
rect 442826 335898 443062 336134
rect 443146 335898 443382 336134
rect 442826 300218 443062 300454
rect 443146 300218 443382 300454
rect 442826 299898 443062 300134
rect 443146 299898 443382 300134
rect 442826 264218 443062 264454
rect 443146 264218 443382 264454
rect 442826 263898 443062 264134
rect 443146 263898 443382 264134
rect 442826 228218 443062 228454
rect 443146 228218 443382 228454
rect 442826 227898 443062 228134
rect 443146 227898 443382 228134
rect 442826 192218 443062 192454
rect 443146 192218 443382 192454
rect 442826 191898 443062 192134
rect 443146 191898 443382 192134
rect 442826 156218 443062 156454
rect 443146 156218 443382 156454
rect 442826 155898 443062 156134
rect 443146 155898 443382 156134
rect 442826 120218 443062 120454
rect 443146 120218 443382 120454
rect 442826 119898 443062 120134
rect 443146 119898 443382 120134
rect 442826 84218 443062 84454
rect 443146 84218 443382 84454
rect 442826 83898 443062 84134
rect 443146 83898 443382 84134
rect 442826 48218 443062 48454
rect 443146 48218 443382 48454
rect 442826 47898 443062 48134
rect 443146 47898 443382 48134
rect 442826 12218 443062 12454
rect 443146 12218 443382 12454
rect 442826 11898 443062 12134
rect 443146 11898 443382 12134
rect 442826 -2502 443062 -2266
rect 443146 -2502 443382 -2266
rect 442826 -2822 443062 -2586
rect 443146 -2822 443382 -2586
rect 447326 707482 447562 707718
rect 447646 707482 447882 707718
rect 447326 707162 447562 707398
rect 447646 707162 447882 707398
rect 447326 700718 447562 700954
rect 447646 700718 447882 700954
rect 447326 700398 447562 700634
rect 447646 700398 447882 700634
rect 447326 664718 447562 664954
rect 447646 664718 447882 664954
rect 447326 664398 447562 664634
rect 447646 664398 447882 664634
rect 447326 628718 447562 628954
rect 447646 628718 447882 628954
rect 447326 628398 447562 628634
rect 447646 628398 447882 628634
rect 447326 592718 447562 592954
rect 447646 592718 447882 592954
rect 447326 592398 447562 592634
rect 447646 592398 447882 592634
rect 447326 556718 447562 556954
rect 447646 556718 447882 556954
rect 447326 556398 447562 556634
rect 447646 556398 447882 556634
rect 447326 520718 447562 520954
rect 447646 520718 447882 520954
rect 447326 520398 447562 520634
rect 447646 520398 447882 520634
rect 447326 484718 447562 484954
rect 447646 484718 447882 484954
rect 447326 484398 447562 484634
rect 447646 484398 447882 484634
rect 447326 448718 447562 448954
rect 447646 448718 447882 448954
rect 447326 448398 447562 448634
rect 447646 448398 447882 448634
rect 447326 412718 447562 412954
rect 447646 412718 447882 412954
rect 447326 412398 447562 412634
rect 447646 412398 447882 412634
rect 447326 376718 447562 376954
rect 447646 376718 447882 376954
rect 447326 376398 447562 376634
rect 447646 376398 447882 376634
rect 447326 340718 447562 340954
rect 447646 340718 447882 340954
rect 447326 340398 447562 340634
rect 447646 340398 447882 340634
rect 447326 304718 447562 304954
rect 447646 304718 447882 304954
rect 447326 304398 447562 304634
rect 447646 304398 447882 304634
rect 447326 268718 447562 268954
rect 447646 268718 447882 268954
rect 447326 268398 447562 268634
rect 447646 268398 447882 268634
rect 447326 232718 447562 232954
rect 447646 232718 447882 232954
rect 447326 232398 447562 232634
rect 447646 232398 447882 232634
rect 447326 196718 447562 196954
rect 447646 196718 447882 196954
rect 447326 196398 447562 196634
rect 447646 196398 447882 196634
rect 447326 160718 447562 160954
rect 447646 160718 447882 160954
rect 447326 160398 447562 160634
rect 447646 160398 447882 160634
rect 447326 124718 447562 124954
rect 447646 124718 447882 124954
rect 447326 124398 447562 124634
rect 447646 124398 447882 124634
rect 447326 88718 447562 88954
rect 447646 88718 447882 88954
rect 447326 88398 447562 88634
rect 447646 88398 447882 88634
rect 447326 52718 447562 52954
rect 447646 52718 447882 52954
rect 447326 52398 447562 52634
rect 447646 52398 447882 52634
rect 447326 16718 447562 16954
rect 447646 16718 447882 16954
rect 447326 16398 447562 16634
rect 447646 16398 447882 16634
rect 447326 -3462 447562 -3226
rect 447646 -3462 447882 -3226
rect 447326 -3782 447562 -3546
rect 447646 -3782 447882 -3546
rect 451826 708442 452062 708678
rect 452146 708442 452382 708678
rect 451826 708122 452062 708358
rect 452146 708122 452382 708358
rect 451826 669218 452062 669454
rect 452146 669218 452382 669454
rect 451826 668898 452062 669134
rect 452146 668898 452382 669134
rect 451826 633218 452062 633454
rect 452146 633218 452382 633454
rect 451826 632898 452062 633134
rect 452146 632898 452382 633134
rect 451826 597218 452062 597454
rect 452146 597218 452382 597454
rect 451826 596898 452062 597134
rect 452146 596898 452382 597134
rect 451826 561218 452062 561454
rect 452146 561218 452382 561454
rect 451826 560898 452062 561134
rect 452146 560898 452382 561134
rect 451826 525218 452062 525454
rect 452146 525218 452382 525454
rect 451826 524898 452062 525134
rect 452146 524898 452382 525134
rect 451826 489218 452062 489454
rect 452146 489218 452382 489454
rect 451826 488898 452062 489134
rect 452146 488898 452382 489134
rect 451826 453218 452062 453454
rect 452146 453218 452382 453454
rect 451826 452898 452062 453134
rect 452146 452898 452382 453134
rect 451826 417218 452062 417454
rect 452146 417218 452382 417454
rect 451826 416898 452062 417134
rect 452146 416898 452382 417134
rect 451826 381218 452062 381454
rect 452146 381218 452382 381454
rect 451826 380898 452062 381134
rect 452146 380898 452382 381134
rect 451826 345218 452062 345454
rect 452146 345218 452382 345454
rect 451826 344898 452062 345134
rect 452146 344898 452382 345134
rect 451826 309218 452062 309454
rect 452146 309218 452382 309454
rect 451826 308898 452062 309134
rect 452146 308898 452382 309134
rect 451826 273218 452062 273454
rect 452146 273218 452382 273454
rect 451826 272898 452062 273134
rect 452146 272898 452382 273134
rect 451826 237218 452062 237454
rect 452146 237218 452382 237454
rect 451826 236898 452062 237134
rect 452146 236898 452382 237134
rect 451826 201218 452062 201454
rect 452146 201218 452382 201454
rect 451826 200898 452062 201134
rect 452146 200898 452382 201134
rect 451826 165218 452062 165454
rect 452146 165218 452382 165454
rect 451826 164898 452062 165134
rect 452146 164898 452382 165134
rect 451826 129218 452062 129454
rect 452146 129218 452382 129454
rect 451826 128898 452062 129134
rect 452146 128898 452382 129134
rect 451826 93218 452062 93454
rect 452146 93218 452382 93454
rect 451826 92898 452062 93134
rect 452146 92898 452382 93134
rect 451826 57218 452062 57454
rect 452146 57218 452382 57454
rect 451826 56898 452062 57134
rect 452146 56898 452382 57134
rect 451826 21218 452062 21454
rect 452146 21218 452382 21454
rect 451826 20898 452062 21134
rect 452146 20898 452382 21134
rect 451826 -4422 452062 -4186
rect 452146 -4422 452382 -4186
rect 451826 -4742 452062 -4506
rect 452146 -4742 452382 -4506
rect 456326 709402 456562 709638
rect 456646 709402 456882 709638
rect 456326 709082 456562 709318
rect 456646 709082 456882 709318
rect 456326 673718 456562 673954
rect 456646 673718 456882 673954
rect 456326 673398 456562 673634
rect 456646 673398 456882 673634
rect 456326 637718 456562 637954
rect 456646 637718 456882 637954
rect 456326 637398 456562 637634
rect 456646 637398 456882 637634
rect 456326 601718 456562 601954
rect 456646 601718 456882 601954
rect 456326 601398 456562 601634
rect 456646 601398 456882 601634
rect 456326 565718 456562 565954
rect 456646 565718 456882 565954
rect 456326 565398 456562 565634
rect 456646 565398 456882 565634
rect 456326 529718 456562 529954
rect 456646 529718 456882 529954
rect 456326 529398 456562 529634
rect 456646 529398 456882 529634
rect 456326 493718 456562 493954
rect 456646 493718 456882 493954
rect 456326 493398 456562 493634
rect 456646 493398 456882 493634
rect 456326 457718 456562 457954
rect 456646 457718 456882 457954
rect 456326 457398 456562 457634
rect 456646 457398 456882 457634
rect 456326 421718 456562 421954
rect 456646 421718 456882 421954
rect 456326 421398 456562 421634
rect 456646 421398 456882 421634
rect 456326 385718 456562 385954
rect 456646 385718 456882 385954
rect 456326 385398 456562 385634
rect 456646 385398 456882 385634
rect 456326 349718 456562 349954
rect 456646 349718 456882 349954
rect 456326 349398 456562 349634
rect 456646 349398 456882 349634
rect 456326 313718 456562 313954
rect 456646 313718 456882 313954
rect 456326 313398 456562 313634
rect 456646 313398 456882 313634
rect 456326 277718 456562 277954
rect 456646 277718 456882 277954
rect 456326 277398 456562 277634
rect 456646 277398 456882 277634
rect 456326 241718 456562 241954
rect 456646 241718 456882 241954
rect 456326 241398 456562 241634
rect 456646 241398 456882 241634
rect 456326 205718 456562 205954
rect 456646 205718 456882 205954
rect 456326 205398 456562 205634
rect 456646 205398 456882 205634
rect 456326 169718 456562 169954
rect 456646 169718 456882 169954
rect 456326 169398 456562 169634
rect 456646 169398 456882 169634
rect 456326 133718 456562 133954
rect 456646 133718 456882 133954
rect 456326 133398 456562 133634
rect 456646 133398 456882 133634
rect 456326 97718 456562 97954
rect 456646 97718 456882 97954
rect 456326 97398 456562 97634
rect 456646 97398 456882 97634
rect 456326 61718 456562 61954
rect 456646 61718 456882 61954
rect 456326 61398 456562 61634
rect 456646 61398 456882 61634
rect 456326 25718 456562 25954
rect 456646 25718 456882 25954
rect 456326 25398 456562 25634
rect 456646 25398 456882 25634
rect 456326 -5382 456562 -5146
rect 456646 -5382 456882 -5146
rect 456326 -5702 456562 -5466
rect 456646 -5702 456882 -5466
rect 460826 710362 461062 710598
rect 461146 710362 461382 710598
rect 460826 710042 461062 710278
rect 461146 710042 461382 710278
rect 460826 678218 461062 678454
rect 461146 678218 461382 678454
rect 460826 677898 461062 678134
rect 461146 677898 461382 678134
rect 460826 642218 461062 642454
rect 461146 642218 461382 642454
rect 460826 641898 461062 642134
rect 461146 641898 461382 642134
rect 460826 606218 461062 606454
rect 461146 606218 461382 606454
rect 460826 605898 461062 606134
rect 461146 605898 461382 606134
rect 460826 570218 461062 570454
rect 461146 570218 461382 570454
rect 460826 569898 461062 570134
rect 461146 569898 461382 570134
rect 460826 534218 461062 534454
rect 461146 534218 461382 534454
rect 460826 533898 461062 534134
rect 461146 533898 461382 534134
rect 460826 498218 461062 498454
rect 461146 498218 461382 498454
rect 460826 497898 461062 498134
rect 461146 497898 461382 498134
rect 460826 462218 461062 462454
rect 461146 462218 461382 462454
rect 460826 461898 461062 462134
rect 461146 461898 461382 462134
rect 460826 426218 461062 426454
rect 461146 426218 461382 426454
rect 460826 425898 461062 426134
rect 461146 425898 461382 426134
rect 460826 390218 461062 390454
rect 461146 390218 461382 390454
rect 460826 389898 461062 390134
rect 461146 389898 461382 390134
rect 460826 354218 461062 354454
rect 461146 354218 461382 354454
rect 460826 353898 461062 354134
rect 461146 353898 461382 354134
rect 460826 318218 461062 318454
rect 461146 318218 461382 318454
rect 460826 317898 461062 318134
rect 461146 317898 461382 318134
rect 460826 282218 461062 282454
rect 461146 282218 461382 282454
rect 460826 281898 461062 282134
rect 461146 281898 461382 282134
rect 460826 246218 461062 246454
rect 461146 246218 461382 246454
rect 460826 245898 461062 246134
rect 461146 245898 461382 246134
rect 460826 210218 461062 210454
rect 461146 210218 461382 210454
rect 460826 209898 461062 210134
rect 461146 209898 461382 210134
rect 460826 174218 461062 174454
rect 461146 174218 461382 174454
rect 460826 173898 461062 174134
rect 461146 173898 461382 174134
rect 460826 138218 461062 138454
rect 461146 138218 461382 138454
rect 460826 137898 461062 138134
rect 461146 137898 461382 138134
rect 460826 102218 461062 102454
rect 461146 102218 461382 102454
rect 460826 101898 461062 102134
rect 461146 101898 461382 102134
rect 460826 66218 461062 66454
rect 461146 66218 461382 66454
rect 460826 65898 461062 66134
rect 461146 65898 461382 66134
rect 460826 30218 461062 30454
rect 461146 30218 461382 30454
rect 460826 29898 461062 30134
rect 461146 29898 461382 30134
rect 460826 -6342 461062 -6106
rect 461146 -6342 461382 -6106
rect 460826 -6662 461062 -6426
rect 461146 -6662 461382 -6426
rect 465326 711322 465562 711558
rect 465646 711322 465882 711558
rect 465326 711002 465562 711238
rect 465646 711002 465882 711238
rect 465326 682718 465562 682954
rect 465646 682718 465882 682954
rect 465326 682398 465562 682634
rect 465646 682398 465882 682634
rect 465326 646718 465562 646954
rect 465646 646718 465882 646954
rect 465326 646398 465562 646634
rect 465646 646398 465882 646634
rect 465326 610718 465562 610954
rect 465646 610718 465882 610954
rect 465326 610398 465562 610634
rect 465646 610398 465882 610634
rect 465326 574718 465562 574954
rect 465646 574718 465882 574954
rect 465326 574398 465562 574634
rect 465646 574398 465882 574634
rect 465326 538718 465562 538954
rect 465646 538718 465882 538954
rect 465326 538398 465562 538634
rect 465646 538398 465882 538634
rect 465326 502718 465562 502954
rect 465646 502718 465882 502954
rect 465326 502398 465562 502634
rect 465646 502398 465882 502634
rect 465326 466718 465562 466954
rect 465646 466718 465882 466954
rect 465326 466398 465562 466634
rect 465646 466398 465882 466634
rect 465326 430718 465562 430954
rect 465646 430718 465882 430954
rect 465326 430398 465562 430634
rect 465646 430398 465882 430634
rect 465326 394718 465562 394954
rect 465646 394718 465882 394954
rect 465326 394398 465562 394634
rect 465646 394398 465882 394634
rect 465326 358718 465562 358954
rect 465646 358718 465882 358954
rect 465326 358398 465562 358634
rect 465646 358398 465882 358634
rect 465326 322718 465562 322954
rect 465646 322718 465882 322954
rect 465326 322398 465562 322634
rect 465646 322398 465882 322634
rect 465326 286718 465562 286954
rect 465646 286718 465882 286954
rect 465326 286398 465562 286634
rect 465646 286398 465882 286634
rect 465326 250718 465562 250954
rect 465646 250718 465882 250954
rect 465326 250398 465562 250634
rect 465646 250398 465882 250634
rect 465326 214718 465562 214954
rect 465646 214718 465882 214954
rect 465326 214398 465562 214634
rect 465646 214398 465882 214634
rect 465326 178718 465562 178954
rect 465646 178718 465882 178954
rect 465326 178398 465562 178634
rect 465646 178398 465882 178634
rect 465326 142718 465562 142954
rect 465646 142718 465882 142954
rect 465326 142398 465562 142634
rect 465646 142398 465882 142634
rect 465326 106718 465562 106954
rect 465646 106718 465882 106954
rect 465326 106398 465562 106634
rect 465646 106398 465882 106634
rect 465326 70718 465562 70954
rect 465646 70718 465882 70954
rect 465326 70398 465562 70634
rect 465646 70398 465882 70634
rect 465326 34718 465562 34954
rect 465646 34718 465882 34954
rect 465326 34398 465562 34634
rect 465646 34398 465882 34634
rect 465326 -7302 465562 -7066
rect 465646 -7302 465882 -7066
rect 465326 -7622 465562 -7386
rect 465646 -7622 465882 -7386
rect 469826 704602 470062 704838
rect 470146 704602 470382 704838
rect 469826 704282 470062 704518
rect 470146 704282 470382 704518
rect 469826 687218 470062 687454
rect 470146 687218 470382 687454
rect 469826 686898 470062 687134
rect 470146 686898 470382 687134
rect 469826 651218 470062 651454
rect 470146 651218 470382 651454
rect 469826 650898 470062 651134
rect 470146 650898 470382 651134
rect 469826 615218 470062 615454
rect 470146 615218 470382 615454
rect 469826 614898 470062 615134
rect 470146 614898 470382 615134
rect 469826 579218 470062 579454
rect 470146 579218 470382 579454
rect 469826 578898 470062 579134
rect 470146 578898 470382 579134
rect 469826 543218 470062 543454
rect 470146 543218 470382 543454
rect 469826 542898 470062 543134
rect 470146 542898 470382 543134
rect 469826 507218 470062 507454
rect 470146 507218 470382 507454
rect 469826 506898 470062 507134
rect 470146 506898 470382 507134
rect 469826 471218 470062 471454
rect 470146 471218 470382 471454
rect 469826 470898 470062 471134
rect 470146 470898 470382 471134
rect 469826 435218 470062 435454
rect 470146 435218 470382 435454
rect 469826 434898 470062 435134
rect 470146 434898 470382 435134
rect 469826 399218 470062 399454
rect 470146 399218 470382 399454
rect 469826 398898 470062 399134
rect 470146 398898 470382 399134
rect 469826 363218 470062 363454
rect 470146 363218 470382 363454
rect 469826 362898 470062 363134
rect 470146 362898 470382 363134
rect 469826 327218 470062 327454
rect 470146 327218 470382 327454
rect 469826 326898 470062 327134
rect 470146 326898 470382 327134
rect 469826 291218 470062 291454
rect 470146 291218 470382 291454
rect 469826 290898 470062 291134
rect 470146 290898 470382 291134
rect 469826 255218 470062 255454
rect 470146 255218 470382 255454
rect 469826 254898 470062 255134
rect 470146 254898 470382 255134
rect 469826 219218 470062 219454
rect 470146 219218 470382 219454
rect 469826 218898 470062 219134
rect 470146 218898 470382 219134
rect 469826 183218 470062 183454
rect 470146 183218 470382 183454
rect 469826 182898 470062 183134
rect 470146 182898 470382 183134
rect 469826 147218 470062 147454
rect 470146 147218 470382 147454
rect 469826 146898 470062 147134
rect 470146 146898 470382 147134
rect 469826 111218 470062 111454
rect 470146 111218 470382 111454
rect 469826 110898 470062 111134
rect 470146 110898 470382 111134
rect 469826 75218 470062 75454
rect 470146 75218 470382 75454
rect 469826 74898 470062 75134
rect 470146 74898 470382 75134
rect 469826 39218 470062 39454
rect 470146 39218 470382 39454
rect 469826 38898 470062 39134
rect 470146 38898 470382 39134
rect 469826 3218 470062 3454
rect 470146 3218 470382 3454
rect 469826 2898 470062 3134
rect 470146 2898 470382 3134
rect 469826 -582 470062 -346
rect 470146 -582 470382 -346
rect 469826 -902 470062 -666
rect 470146 -902 470382 -666
rect 474326 705562 474562 705798
rect 474646 705562 474882 705798
rect 474326 705242 474562 705478
rect 474646 705242 474882 705478
rect 474326 691718 474562 691954
rect 474646 691718 474882 691954
rect 474326 691398 474562 691634
rect 474646 691398 474882 691634
rect 474326 655718 474562 655954
rect 474646 655718 474882 655954
rect 474326 655398 474562 655634
rect 474646 655398 474882 655634
rect 474326 619718 474562 619954
rect 474646 619718 474882 619954
rect 474326 619398 474562 619634
rect 474646 619398 474882 619634
rect 474326 583718 474562 583954
rect 474646 583718 474882 583954
rect 474326 583398 474562 583634
rect 474646 583398 474882 583634
rect 474326 547718 474562 547954
rect 474646 547718 474882 547954
rect 474326 547398 474562 547634
rect 474646 547398 474882 547634
rect 474326 511718 474562 511954
rect 474646 511718 474882 511954
rect 474326 511398 474562 511634
rect 474646 511398 474882 511634
rect 474326 475718 474562 475954
rect 474646 475718 474882 475954
rect 474326 475398 474562 475634
rect 474646 475398 474882 475634
rect 474326 439718 474562 439954
rect 474646 439718 474882 439954
rect 474326 439398 474562 439634
rect 474646 439398 474882 439634
rect 474326 403718 474562 403954
rect 474646 403718 474882 403954
rect 474326 403398 474562 403634
rect 474646 403398 474882 403634
rect 474326 367718 474562 367954
rect 474646 367718 474882 367954
rect 474326 367398 474562 367634
rect 474646 367398 474882 367634
rect 474326 331718 474562 331954
rect 474646 331718 474882 331954
rect 474326 331398 474562 331634
rect 474646 331398 474882 331634
rect 474326 295718 474562 295954
rect 474646 295718 474882 295954
rect 474326 295398 474562 295634
rect 474646 295398 474882 295634
rect 474326 259718 474562 259954
rect 474646 259718 474882 259954
rect 474326 259398 474562 259634
rect 474646 259398 474882 259634
rect 474326 223718 474562 223954
rect 474646 223718 474882 223954
rect 474326 223398 474562 223634
rect 474646 223398 474882 223634
rect 474326 187718 474562 187954
rect 474646 187718 474882 187954
rect 474326 187398 474562 187634
rect 474646 187398 474882 187634
rect 474326 151718 474562 151954
rect 474646 151718 474882 151954
rect 474326 151398 474562 151634
rect 474646 151398 474882 151634
rect 474326 115718 474562 115954
rect 474646 115718 474882 115954
rect 474326 115398 474562 115634
rect 474646 115398 474882 115634
rect 474326 79718 474562 79954
rect 474646 79718 474882 79954
rect 474326 79398 474562 79634
rect 474646 79398 474882 79634
rect 474326 43718 474562 43954
rect 474646 43718 474882 43954
rect 474326 43398 474562 43634
rect 474646 43398 474882 43634
rect 474326 7718 474562 7954
rect 474646 7718 474882 7954
rect 474326 7398 474562 7634
rect 474646 7398 474882 7634
rect 474326 -1542 474562 -1306
rect 474646 -1542 474882 -1306
rect 474326 -1862 474562 -1626
rect 474646 -1862 474882 -1626
rect 478826 706522 479062 706758
rect 479146 706522 479382 706758
rect 478826 706202 479062 706438
rect 479146 706202 479382 706438
rect 478826 696218 479062 696454
rect 479146 696218 479382 696454
rect 478826 695898 479062 696134
rect 479146 695898 479382 696134
rect 478826 660218 479062 660454
rect 479146 660218 479382 660454
rect 478826 659898 479062 660134
rect 479146 659898 479382 660134
rect 478826 624218 479062 624454
rect 479146 624218 479382 624454
rect 478826 623898 479062 624134
rect 479146 623898 479382 624134
rect 478826 588218 479062 588454
rect 479146 588218 479382 588454
rect 478826 587898 479062 588134
rect 479146 587898 479382 588134
rect 478826 552218 479062 552454
rect 479146 552218 479382 552454
rect 478826 551898 479062 552134
rect 479146 551898 479382 552134
rect 478826 516218 479062 516454
rect 479146 516218 479382 516454
rect 478826 515898 479062 516134
rect 479146 515898 479382 516134
rect 478826 480218 479062 480454
rect 479146 480218 479382 480454
rect 478826 479898 479062 480134
rect 479146 479898 479382 480134
rect 478826 444218 479062 444454
rect 479146 444218 479382 444454
rect 478826 443898 479062 444134
rect 479146 443898 479382 444134
rect 478826 408218 479062 408454
rect 479146 408218 479382 408454
rect 478826 407898 479062 408134
rect 479146 407898 479382 408134
rect 478826 372218 479062 372454
rect 479146 372218 479382 372454
rect 478826 371898 479062 372134
rect 479146 371898 479382 372134
rect 478826 336218 479062 336454
rect 479146 336218 479382 336454
rect 478826 335898 479062 336134
rect 479146 335898 479382 336134
rect 478826 300218 479062 300454
rect 479146 300218 479382 300454
rect 478826 299898 479062 300134
rect 479146 299898 479382 300134
rect 478826 264218 479062 264454
rect 479146 264218 479382 264454
rect 478826 263898 479062 264134
rect 479146 263898 479382 264134
rect 478826 228218 479062 228454
rect 479146 228218 479382 228454
rect 478826 227898 479062 228134
rect 479146 227898 479382 228134
rect 478826 192218 479062 192454
rect 479146 192218 479382 192454
rect 478826 191898 479062 192134
rect 479146 191898 479382 192134
rect 478826 156218 479062 156454
rect 479146 156218 479382 156454
rect 478826 155898 479062 156134
rect 479146 155898 479382 156134
rect 478826 120218 479062 120454
rect 479146 120218 479382 120454
rect 478826 119898 479062 120134
rect 479146 119898 479382 120134
rect 478826 84218 479062 84454
rect 479146 84218 479382 84454
rect 478826 83898 479062 84134
rect 479146 83898 479382 84134
rect 478826 48218 479062 48454
rect 479146 48218 479382 48454
rect 478826 47898 479062 48134
rect 479146 47898 479382 48134
rect 478826 12218 479062 12454
rect 479146 12218 479382 12454
rect 478826 11898 479062 12134
rect 479146 11898 479382 12134
rect 478826 -2502 479062 -2266
rect 479146 -2502 479382 -2266
rect 478826 -2822 479062 -2586
rect 479146 -2822 479382 -2586
rect 483326 707482 483562 707718
rect 483646 707482 483882 707718
rect 483326 707162 483562 707398
rect 483646 707162 483882 707398
rect 483326 700718 483562 700954
rect 483646 700718 483882 700954
rect 483326 700398 483562 700634
rect 483646 700398 483882 700634
rect 483326 664718 483562 664954
rect 483646 664718 483882 664954
rect 483326 664398 483562 664634
rect 483646 664398 483882 664634
rect 483326 628718 483562 628954
rect 483646 628718 483882 628954
rect 483326 628398 483562 628634
rect 483646 628398 483882 628634
rect 483326 592718 483562 592954
rect 483646 592718 483882 592954
rect 483326 592398 483562 592634
rect 483646 592398 483882 592634
rect 483326 556718 483562 556954
rect 483646 556718 483882 556954
rect 483326 556398 483562 556634
rect 483646 556398 483882 556634
rect 483326 520718 483562 520954
rect 483646 520718 483882 520954
rect 483326 520398 483562 520634
rect 483646 520398 483882 520634
rect 483326 484718 483562 484954
rect 483646 484718 483882 484954
rect 483326 484398 483562 484634
rect 483646 484398 483882 484634
rect 483326 448718 483562 448954
rect 483646 448718 483882 448954
rect 483326 448398 483562 448634
rect 483646 448398 483882 448634
rect 483326 412718 483562 412954
rect 483646 412718 483882 412954
rect 483326 412398 483562 412634
rect 483646 412398 483882 412634
rect 483326 376718 483562 376954
rect 483646 376718 483882 376954
rect 483326 376398 483562 376634
rect 483646 376398 483882 376634
rect 483326 340718 483562 340954
rect 483646 340718 483882 340954
rect 483326 340398 483562 340634
rect 483646 340398 483882 340634
rect 483326 304718 483562 304954
rect 483646 304718 483882 304954
rect 483326 304398 483562 304634
rect 483646 304398 483882 304634
rect 483326 268718 483562 268954
rect 483646 268718 483882 268954
rect 483326 268398 483562 268634
rect 483646 268398 483882 268634
rect 483326 232718 483562 232954
rect 483646 232718 483882 232954
rect 483326 232398 483562 232634
rect 483646 232398 483882 232634
rect 483326 196718 483562 196954
rect 483646 196718 483882 196954
rect 483326 196398 483562 196634
rect 483646 196398 483882 196634
rect 483326 160718 483562 160954
rect 483646 160718 483882 160954
rect 483326 160398 483562 160634
rect 483646 160398 483882 160634
rect 483326 124718 483562 124954
rect 483646 124718 483882 124954
rect 483326 124398 483562 124634
rect 483646 124398 483882 124634
rect 483326 88718 483562 88954
rect 483646 88718 483882 88954
rect 483326 88398 483562 88634
rect 483646 88398 483882 88634
rect 483326 52718 483562 52954
rect 483646 52718 483882 52954
rect 483326 52398 483562 52634
rect 483646 52398 483882 52634
rect 483326 16718 483562 16954
rect 483646 16718 483882 16954
rect 483326 16398 483562 16634
rect 483646 16398 483882 16634
rect 483326 -3462 483562 -3226
rect 483646 -3462 483882 -3226
rect 483326 -3782 483562 -3546
rect 483646 -3782 483882 -3546
rect 487826 708442 488062 708678
rect 488146 708442 488382 708678
rect 487826 708122 488062 708358
rect 488146 708122 488382 708358
rect 487826 669218 488062 669454
rect 488146 669218 488382 669454
rect 487826 668898 488062 669134
rect 488146 668898 488382 669134
rect 487826 633218 488062 633454
rect 488146 633218 488382 633454
rect 487826 632898 488062 633134
rect 488146 632898 488382 633134
rect 487826 597218 488062 597454
rect 488146 597218 488382 597454
rect 487826 596898 488062 597134
rect 488146 596898 488382 597134
rect 487826 561218 488062 561454
rect 488146 561218 488382 561454
rect 487826 560898 488062 561134
rect 488146 560898 488382 561134
rect 487826 525218 488062 525454
rect 488146 525218 488382 525454
rect 487826 524898 488062 525134
rect 488146 524898 488382 525134
rect 487826 489218 488062 489454
rect 488146 489218 488382 489454
rect 487826 488898 488062 489134
rect 488146 488898 488382 489134
rect 487826 453218 488062 453454
rect 488146 453218 488382 453454
rect 487826 452898 488062 453134
rect 488146 452898 488382 453134
rect 487826 417218 488062 417454
rect 488146 417218 488382 417454
rect 487826 416898 488062 417134
rect 488146 416898 488382 417134
rect 487826 381218 488062 381454
rect 488146 381218 488382 381454
rect 487826 380898 488062 381134
rect 488146 380898 488382 381134
rect 487826 345218 488062 345454
rect 488146 345218 488382 345454
rect 487826 344898 488062 345134
rect 488146 344898 488382 345134
rect 487826 309218 488062 309454
rect 488146 309218 488382 309454
rect 487826 308898 488062 309134
rect 488146 308898 488382 309134
rect 487826 273218 488062 273454
rect 488146 273218 488382 273454
rect 487826 272898 488062 273134
rect 488146 272898 488382 273134
rect 487826 237218 488062 237454
rect 488146 237218 488382 237454
rect 487826 236898 488062 237134
rect 488146 236898 488382 237134
rect 487826 201218 488062 201454
rect 488146 201218 488382 201454
rect 487826 200898 488062 201134
rect 488146 200898 488382 201134
rect 487826 165218 488062 165454
rect 488146 165218 488382 165454
rect 487826 164898 488062 165134
rect 488146 164898 488382 165134
rect 487826 129218 488062 129454
rect 488146 129218 488382 129454
rect 487826 128898 488062 129134
rect 488146 128898 488382 129134
rect 487826 93218 488062 93454
rect 488146 93218 488382 93454
rect 487826 92898 488062 93134
rect 488146 92898 488382 93134
rect 487826 57218 488062 57454
rect 488146 57218 488382 57454
rect 487826 56898 488062 57134
rect 488146 56898 488382 57134
rect 487826 21218 488062 21454
rect 488146 21218 488382 21454
rect 487826 20898 488062 21134
rect 488146 20898 488382 21134
rect 487826 -4422 488062 -4186
rect 488146 -4422 488382 -4186
rect 487826 -4742 488062 -4506
rect 488146 -4742 488382 -4506
rect 492326 709402 492562 709638
rect 492646 709402 492882 709638
rect 492326 709082 492562 709318
rect 492646 709082 492882 709318
rect 492326 673718 492562 673954
rect 492646 673718 492882 673954
rect 492326 673398 492562 673634
rect 492646 673398 492882 673634
rect 492326 637718 492562 637954
rect 492646 637718 492882 637954
rect 492326 637398 492562 637634
rect 492646 637398 492882 637634
rect 492326 601718 492562 601954
rect 492646 601718 492882 601954
rect 492326 601398 492562 601634
rect 492646 601398 492882 601634
rect 492326 565718 492562 565954
rect 492646 565718 492882 565954
rect 492326 565398 492562 565634
rect 492646 565398 492882 565634
rect 492326 529718 492562 529954
rect 492646 529718 492882 529954
rect 492326 529398 492562 529634
rect 492646 529398 492882 529634
rect 492326 493718 492562 493954
rect 492646 493718 492882 493954
rect 492326 493398 492562 493634
rect 492646 493398 492882 493634
rect 492326 457718 492562 457954
rect 492646 457718 492882 457954
rect 492326 457398 492562 457634
rect 492646 457398 492882 457634
rect 492326 421718 492562 421954
rect 492646 421718 492882 421954
rect 492326 421398 492562 421634
rect 492646 421398 492882 421634
rect 492326 385718 492562 385954
rect 492646 385718 492882 385954
rect 492326 385398 492562 385634
rect 492646 385398 492882 385634
rect 492326 349718 492562 349954
rect 492646 349718 492882 349954
rect 492326 349398 492562 349634
rect 492646 349398 492882 349634
rect 492326 313718 492562 313954
rect 492646 313718 492882 313954
rect 492326 313398 492562 313634
rect 492646 313398 492882 313634
rect 492326 277718 492562 277954
rect 492646 277718 492882 277954
rect 492326 277398 492562 277634
rect 492646 277398 492882 277634
rect 492326 241718 492562 241954
rect 492646 241718 492882 241954
rect 492326 241398 492562 241634
rect 492646 241398 492882 241634
rect 492326 205718 492562 205954
rect 492646 205718 492882 205954
rect 492326 205398 492562 205634
rect 492646 205398 492882 205634
rect 492326 169718 492562 169954
rect 492646 169718 492882 169954
rect 492326 169398 492562 169634
rect 492646 169398 492882 169634
rect 492326 133718 492562 133954
rect 492646 133718 492882 133954
rect 492326 133398 492562 133634
rect 492646 133398 492882 133634
rect 492326 97718 492562 97954
rect 492646 97718 492882 97954
rect 492326 97398 492562 97634
rect 492646 97398 492882 97634
rect 492326 61718 492562 61954
rect 492646 61718 492882 61954
rect 492326 61398 492562 61634
rect 492646 61398 492882 61634
rect 492326 25718 492562 25954
rect 492646 25718 492882 25954
rect 492326 25398 492562 25634
rect 492646 25398 492882 25634
rect 492326 -5382 492562 -5146
rect 492646 -5382 492882 -5146
rect 492326 -5702 492562 -5466
rect 492646 -5702 492882 -5466
rect 496826 710362 497062 710598
rect 497146 710362 497382 710598
rect 496826 710042 497062 710278
rect 497146 710042 497382 710278
rect 496826 678218 497062 678454
rect 497146 678218 497382 678454
rect 496826 677898 497062 678134
rect 497146 677898 497382 678134
rect 496826 642218 497062 642454
rect 497146 642218 497382 642454
rect 496826 641898 497062 642134
rect 497146 641898 497382 642134
rect 496826 606218 497062 606454
rect 497146 606218 497382 606454
rect 496826 605898 497062 606134
rect 497146 605898 497382 606134
rect 496826 570218 497062 570454
rect 497146 570218 497382 570454
rect 496826 569898 497062 570134
rect 497146 569898 497382 570134
rect 496826 534218 497062 534454
rect 497146 534218 497382 534454
rect 496826 533898 497062 534134
rect 497146 533898 497382 534134
rect 496826 498218 497062 498454
rect 497146 498218 497382 498454
rect 496826 497898 497062 498134
rect 497146 497898 497382 498134
rect 496826 462218 497062 462454
rect 497146 462218 497382 462454
rect 496826 461898 497062 462134
rect 497146 461898 497382 462134
rect 496826 426218 497062 426454
rect 497146 426218 497382 426454
rect 496826 425898 497062 426134
rect 497146 425898 497382 426134
rect 496826 390218 497062 390454
rect 497146 390218 497382 390454
rect 496826 389898 497062 390134
rect 497146 389898 497382 390134
rect 496826 354218 497062 354454
rect 497146 354218 497382 354454
rect 496826 353898 497062 354134
rect 497146 353898 497382 354134
rect 496826 318218 497062 318454
rect 497146 318218 497382 318454
rect 496826 317898 497062 318134
rect 497146 317898 497382 318134
rect 496826 282218 497062 282454
rect 497146 282218 497382 282454
rect 496826 281898 497062 282134
rect 497146 281898 497382 282134
rect 496826 246218 497062 246454
rect 497146 246218 497382 246454
rect 496826 245898 497062 246134
rect 497146 245898 497382 246134
rect 496826 210218 497062 210454
rect 497146 210218 497382 210454
rect 496826 209898 497062 210134
rect 497146 209898 497382 210134
rect 496826 174218 497062 174454
rect 497146 174218 497382 174454
rect 496826 173898 497062 174134
rect 497146 173898 497382 174134
rect 496826 138218 497062 138454
rect 497146 138218 497382 138454
rect 496826 137898 497062 138134
rect 497146 137898 497382 138134
rect 496826 102218 497062 102454
rect 497146 102218 497382 102454
rect 496826 101898 497062 102134
rect 497146 101898 497382 102134
rect 496826 66218 497062 66454
rect 497146 66218 497382 66454
rect 496826 65898 497062 66134
rect 497146 65898 497382 66134
rect 496826 30218 497062 30454
rect 497146 30218 497382 30454
rect 496826 29898 497062 30134
rect 497146 29898 497382 30134
rect 496826 -6342 497062 -6106
rect 497146 -6342 497382 -6106
rect 496826 -6662 497062 -6426
rect 497146 -6662 497382 -6426
rect 501326 711322 501562 711558
rect 501646 711322 501882 711558
rect 501326 711002 501562 711238
rect 501646 711002 501882 711238
rect 501326 682718 501562 682954
rect 501646 682718 501882 682954
rect 501326 682398 501562 682634
rect 501646 682398 501882 682634
rect 501326 646718 501562 646954
rect 501646 646718 501882 646954
rect 501326 646398 501562 646634
rect 501646 646398 501882 646634
rect 501326 610718 501562 610954
rect 501646 610718 501882 610954
rect 501326 610398 501562 610634
rect 501646 610398 501882 610634
rect 501326 574718 501562 574954
rect 501646 574718 501882 574954
rect 501326 574398 501562 574634
rect 501646 574398 501882 574634
rect 501326 538718 501562 538954
rect 501646 538718 501882 538954
rect 501326 538398 501562 538634
rect 501646 538398 501882 538634
rect 501326 502718 501562 502954
rect 501646 502718 501882 502954
rect 501326 502398 501562 502634
rect 501646 502398 501882 502634
rect 501326 466718 501562 466954
rect 501646 466718 501882 466954
rect 501326 466398 501562 466634
rect 501646 466398 501882 466634
rect 501326 430718 501562 430954
rect 501646 430718 501882 430954
rect 501326 430398 501562 430634
rect 501646 430398 501882 430634
rect 501326 394718 501562 394954
rect 501646 394718 501882 394954
rect 501326 394398 501562 394634
rect 501646 394398 501882 394634
rect 501326 358718 501562 358954
rect 501646 358718 501882 358954
rect 501326 358398 501562 358634
rect 501646 358398 501882 358634
rect 501326 322718 501562 322954
rect 501646 322718 501882 322954
rect 501326 322398 501562 322634
rect 501646 322398 501882 322634
rect 501326 286718 501562 286954
rect 501646 286718 501882 286954
rect 501326 286398 501562 286634
rect 501646 286398 501882 286634
rect 501326 250718 501562 250954
rect 501646 250718 501882 250954
rect 501326 250398 501562 250634
rect 501646 250398 501882 250634
rect 501326 214718 501562 214954
rect 501646 214718 501882 214954
rect 501326 214398 501562 214634
rect 501646 214398 501882 214634
rect 501326 178718 501562 178954
rect 501646 178718 501882 178954
rect 501326 178398 501562 178634
rect 501646 178398 501882 178634
rect 501326 142718 501562 142954
rect 501646 142718 501882 142954
rect 501326 142398 501562 142634
rect 501646 142398 501882 142634
rect 501326 106718 501562 106954
rect 501646 106718 501882 106954
rect 501326 106398 501562 106634
rect 501646 106398 501882 106634
rect 501326 70718 501562 70954
rect 501646 70718 501882 70954
rect 501326 70398 501562 70634
rect 501646 70398 501882 70634
rect 501326 34718 501562 34954
rect 501646 34718 501882 34954
rect 501326 34398 501562 34634
rect 501646 34398 501882 34634
rect 501326 -7302 501562 -7066
rect 501646 -7302 501882 -7066
rect 501326 -7622 501562 -7386
rect 501646 -7622 501882 -7386
rect 505826 704602 506062 704838
rect 506146 704602 506382 704838
rect 505826 704282 506062 704518
rect 506146 704282 506382 704518
rect 505826 687218 506062 687454
rect 506146 687218 506382 687454
rect 505826 686898 506062 687134
rect 506146 686898 506382 687134
rect 505826 651218 506062 651454
rect 506146 651218 506382 651454
rect 505826 650898 506062 651134
rect 506146 650898 506382 651134
rect 505826 615218 506062 615454
rect 506146 615218 506382 615454
rect 505826 614898 506062 615134
rect 506146 614898 506382 615134
rect 505826 579218 506062 579454
rect 506146 579218 506382 579454
rect 505826 578898 506062 579134
rect 506146 578898 506382 579134
rect 505826 543218 506062 543454
rect 506146 543218 506382 543454
rect 505826 542898 506062 543134
rect 506146 542898 506382 543134
rect 505826 507218 506062 507454
rect 506146 507218 506382 507454
rect 505826 506898 506062 507134
rect 506146 506898 506382 507134
rect 505826 471218 506062 471454
rect 506146 471218 506382 471454
rect 505826 470898 506062 471134
rect 506146 470898 506382 471134
rect 505826 435218 506062 435454
rect 506146 435218 506382 435454
rect 505826 434898 506062 435134
rect 506146 434898 506382 435134
rect 505826 399218 506062 399454
rect 506146 399218 506382 399454
rect 505826 398898 506062 399134
rect 506146 398898 506382 399134
rect 505826 363218 506062 363454
rect 506146 363218 506382 363454
rect 505826 362898 506062 363134
rect 506146 362898 506382 363134
rect 505826 327218 506062 327454
rect 506146 327218 506382 327454
rect 505826 326898 506062 327134
rect 506146 326898 506382 327134
rect 505826 291218 506062 291454
rect 506146 291218 506382 291454
rect 505826 290898 506062 291134
rect 506146 290898 506382 291134
rect 505826 255218 506062 255454
rect 506146 255218 506382 255454
rect 505826 254898 506062 255134
rect 506146 254898 506382 255134
rect 505826 219218 506062 219454
rect 506146 219218 506382 219454
rect 505826 218898 506062 219134
rect 506146 218898 506382 219134
rect 505826 183218 506062 183454
rect 506146 183218 506382 183454
rect 505826 182898 506062 183134
rect 506146 182898 506382 183134
rect 505826 147218 506062 147454
rect 506146 147218 506382 147454
rect 505826 146898 506062 147134
rect 506146 146898 506382 147134
rect 505826 111218 506062 111454
rect 506146 111218 506382 111454
rect 505826 110898 506062 111134
rect 506146 110898 506382 111134
rect 505826 75218 506062 75454
rect 506146 75218 506382 75454
rect 505826 74898 506062 75134
rect 506146 74898 506382 75134
rect 505826 39218 506062 39454
rect 506146 39218 506382 39454
rect 505826 38898 506062 39134
rect 506146 38898 506382 39134
rect 505826 3218 506062 3454
rect 506146 3218 506382 3454
rect 505826 2898 506062 3134
rect 506146 2898 506382 3134
rect 505826 -582 506062 -346
rect 506146 -582 506382 -346
rect 505826 -902 506062 -666
rect 506146 -902 506382 -666
rect 510326 705562 510562 705798
rect 510646 705562 510882 705798
rect 510326 705242 510562 705478
rect 510646 705242 510882 705478
rect 510326 691718 510562 691954
rect 510646 691718 510882 691954
rect 510326 691398 510562 691634
rect 510646 691398 510882 691634
rect 510326 655718 510562 655954
rect 510646 655718 510882 655954
rect 510326 655398 510562 655634
rect 510646 655398 510882 655634
rect 510326 619718 510562 619954
rect 510646 619718 510882 619954
rect 510326 619398 510562 619634
rect 510646 619398 510882 619634
rect 510326 583718 510562 583954
rect 510646 583718 510882 583954
rect 510326 583398 510562 583634
rect 510646 583398 510882 583634
rect 510326 547718 510562 547954
rect 510646 547718 510882 547954
rect 510326 547398 510562 547634
rect 510646 547398 510882 547634
rect 510326 511718 510562 511954
rect 510646 511718 510882 511954
rect 510326 511398 510562 511634
rect 510646 511398 510882 511634
rect 510326 475718 510562 475954
rect 510646 475718 510882 475954
rect 510326 475398 510562 475634
rect 510646 475398 510882 475634
rect 510326 439718 510562 439954
rect 510646 439718 510882 439954
rect 510326 439398 510562 439634
rect 510646 439398 510882 439634
rect 510326 403718 510562 403954
rect 510646 403718 510882 403954
rect 510326 403398 510562 403634
rect 510646 403398 510882 403634
rect 510326 367718 510562 367954
rect 510646 367718 510882 367954
rect 510326 367398 510562 367634
rect 510646 367398 510882 367634
rect 510326 331718 510562 331954
rect 510646 331718 510882 331954
rect 510326 331398 510562 331634
rect 510646 331398 510882 331634
rect 510326 295718 510562 295954
rect 510646 295718 510882 295954
rect 510326 295398 510562 295634
rect 510646 295398 510882 295634
rect 510326 259718 510562 259954
rect 510646 259718 510882 259954
rect 510326 259398 510562 259634
rect 510646 259398 510882 259634
rect 510326 223718 510562 223954
rect 510646 223718 510882 223954
rect 510326 223398 510562 223634
rect 510646 223398 510882 223634
rect 510326 187718 510562 187954
rect 510646 187718 510882 187954
rect 510326 187398 510562 187634
rect 510646 187398 510882 187634
rect 510326 151718 510562 151954
rect 510646 151718 510882 151954
rect 510326 151398 510562 151634
rect 510646 151398 510882 151634
rect 510326 115718 510562 115954
rect 510646 115718 510882 115954
rect 510326 115398 510562 115634
rect 510646 115398 510882 115634
rect 510326 79718 510562 79954
rect 510646 79718 510882 79954
rect 510326 79398 510562 79634
rect 510646 79398 510882 79634
rect 510326 43718 510562 43954
rect 510646 43718 510882 43954
rect 510326 43398 510562 43634
rect 510646 43398 510882 43634
rect 510326 7718 510562 7954
rect 510646 7718 510882 7954
rect 510326 7398 510562 7634
rect 510646 7398 510882 7634
rect 510326 -1542 510562 -1306
rect 510646 -1542 510882 -1306
rect 510326 -1862 510562 -1626
rect 510646 -1862 510882 -1626
rect 514826 706522 515062 706758
rect 515146 706522 515382 706758
rect 514826 706202 515062 706438
rect 515146 706202 515382 706438
rect 514826 696218 515062 696454
rect 515146 696218 515382 696454
rect 514826 695898 515062 696134
rect 515146 695898 515382 696134
rect 514826 660218 515062 660454
rect 515146 660218 515382 660454
rect 514826 659898 515062 660134
rect 515146 659898 515382 660134
rect 514826 624218 515062 624454
rect 515146 624218 515382 624454
rect 514826 623898 515062 624134
rect 515146 623898 515382 624134
rect 514826 588218 515062 588454
rect 515146 588218 515382 588454
rect 514826 587898 515062 588134
rect 515146 587898 515382 588134
rect 514826 552218 515062 552454
rect 515146 552218 515382 552454
rect 514826 551898 515062 552134
rect 515146 551898 515382 552134
rect 514826 516218 515062 516454
rect 515146 516218 515382 516454
rect 514826 515898 515062 516134
rect 515146 515898 515382 516134
rect 514826 480218 515062 480454
rect 515146 480218 515382 480454
rect 514826 479898 515062 480134
rect 515146 479898 515382 480134
rect 514826 444218 515062 444454
rect 515146 444218 515382 444454
rect 514826 443898 515062 444134
rect 515146 443898 515382 444134
rect 514826 408218 515062 408454
rect 515146 408218 515382 408454
rect 514826 407898 515062 408134
rect 515146 407898 515382 408134
rect 514826 372218 515062 372454
rect 515146 372218 515382 372454
rect 514826 371898 515062 372134
rect 515146 371898 515382 372134
rect 514826 336218 515062 336454
rect 515146 336218 515382 336454
rect 514826 335898 515062 336134
rect 515146 335898 515382 336134
rect 514826 300218 515062 300454
rect 515146 300218 515382 300454
rect 514826 299898 515062 300134
rect 515146 299898 515382 300134
rect 514826 264218 515062 264454
rect 515146 264218 515382 264454
rect 514826 263898 515062 264134
rect 515146 263898 515382 264134
rect 514826 228218 515062 228454
rect 515146 228218 515382 228454
rect 514826 227898 515062 228134
rect 515146 227898 515382 228134
rect 514826 192218 515062 192454
rect 515146 192218 515382 192454
rect 514826 191898 515062 192134
rect 515146 191898 515382 192134
rect 514826 156218 515062 156454
rect 515146 156218 515382 156454
rect 514826 155898 515062 156134
rect 515146 155898 515382 156134
rect 514826 120218 515062 120454
rect 515146 120218 515382 120454
rect 514826 119898 515062 120134
rect 515146 119898 515382 120134
rect 514826 84218 515062 84454
rect 515146 84218 515382 84454
rect 514826 83898 515062 84134
rect 515146 83898 515382 84134
rect 514826 48218 515062 48454
rect 515146 48218 515382 48454
rect 514826 47898 515062 48134
rect 515146 47898 515382 48134
rect 514826 12218 515062 12454
rect 515146 12218 515382 12454
rect 514826 11898 515062 12134
rect 515146 11898 515382 12134
rect 514826 -2502 515062 -2266
rect 515146 -2502 515382 -2266
rect 514826 -2822 515062 -2586
rect 515146 -2822 515382 -2586
rect 519326 707482 519562 707718
rect 519646 707482 519882 707718
rect 519326 707162 519562 707398
rect 519646 707162 519882 707398
rect 519326 700718 519562 700954
rect 519646 700718 519882 700954
rect 519326 700398 519562 700634
rect 519646 700398 519882 700634
rect 519326 664718 519562 664954
rect 519646 664718 519882 664954
rect 519326 664398 519562 664634
rect 519646 664398 519882 664634
rect 519326 628718 519562 628954
rect 519646 628718 519882 628954
rect 519326 628398 519562 628634
rect 519646 628398 519882 628634
rect 519326 592718 519562 592954
rect 519646 592718 519882 592954
rect 519326 592398 519562 592634
rect 519646 592398 519882 592634
rect 519326 556718 519562 556954
rect 519646 556718 519882 556954
rect 519326 556398 519562 556634
rect 519646 556398 519882 556634
rect 519326 520718 519562 520954
rect 519646 520718 519882 520954
rect 519326 520398 519562 520634
rect 519646 520398 519882 520634
rect 519326 484718 519562 484954
rect 519646 484718 519882 484954
rect 519326 484398 519562 484634
rect 519646 484398 519882 484634
rect 519326 448718 519562 448954
rect 519646 448718 519882 448954
rect 519326 448398 519562 448634
rect 519646 448398 519882 448634
rect 519326 412718 519562 412954
rect 519646 412718 519882 412954
rect 519326 412398 519562 412634
rect 519646 412398 519882 412634
rect 519326 376718 519562 376954
rect 519646 376718 519882 376954
rect 519326 376398 519562 376634
rect 519646 376398 519882 376634
rect 519326 340718 519562 340954
rect 519646 340718 519882 340954
rect 519326 340398 519562 340634
rect 519646 340398 519882 340634
rect 519326 304718 519562 304954
rect 519646 304718 519882 304954
rect 519326 304398 519562 304634
rect 519646 304398 519882 304634
rect 519326 268718 519562 268954
rect 519646 268718 519882 268954
rect 519326 268398 519562 268634
rect 519646 268398 519882 268634
rect 519326 232718 519562 232954
rect 519646 232718 519882 232954
rect 519326 232398 519562 232634
rect 519646 232398 519882 232634
rect 519326 196718 519562 196954
rect 519646 196718 519882 196954
rect 519326 196398 519562 196634
rect 519646 196398 519882 196634
rect 519326 160718 519562 160954
rect 519646 160718 519882 160954
rect 519326 160398 519562 160634
rect 519646 160398 519882 160634
rect 519326 124718 519562 124954
rect 519646 124718 519882 124954
rect 519326 124398 519562 124634
rect 519646 124398 519882 124634
rect 519326 88718 519562 88954
rect 519646 88718 519882 88954
rect 519326 88398 519562 88634
rect 519646 88398 519882 88634
rect 519326 52718 519562 52954
rect 519646 52718 519882 52954
rect 519326 52398 519562 52634
rect 519646 52398 519882 52634
rect 519326 16718 519562 16954
rect 519646 16718 519882 16954
rect 519326 16398 519562 16634
rect 519646 16398 519882 16634
rect 519326 -3462 519562 -3226
rect 519646 -3462 519882 -3226
rect 519326 -3782 519562 -3546
rect 519646 -3782 519882 -3546
rect 523826 708442 524062 708678
rect 524146 708442 524382 708678
rect 523826 708122 524062 708358
rect 524146 708122 524382 708358
rect 523826 669218 524062 669454
rect 524146 669218 524382 669454
rect 523826 668898 524062 669134
rect 524146 668898 524382 669134
rect 523826 633218 524062 633454
rect 524146 633218 524382 633454
rect 523826 632898 524062 633134
rect 524146 632898 524382 633134
rect 523826 597218 524062 597454
rect 524146 597218 524382 597454
rect 523826 596898 524062 597134
rect 524146 596898 524382 597134
rect 523826 561218 524062 561454
rect 524146 561218 524382 561454
rect 523826 560898 524062 561134
rect 524146 560898 524382 561134
rect 523826 525218 524062 525454
rect 524146 525218 524382 525454
rect 523826 524898 524062 525134
rect 524146 524898 524382 525134
rect 523826 489218 524062 489454
rect 524146 489218 524382 489454
rect 523826 488898 524062 489134
rect 524146 488898 524382 489134
rect 523826 453218 524062 453454
rect 524146 453218 524382 453454
rect 523826 452898 524062 453134
rect 524146 452898 524382 453134
rect 523826 417218 524062 417454
rect 524146 417218 524382 417454
rect 523826 416898 524062 417134
rect 524146 416898 524382 417134
rect 523826 381218 524062 381454
rect 524146 381218 524382 381454
rect 523826 380898 524062 381134
rect 524146 380898 524382 381134
rect 523826 345218 524062 345454
rect 524146 345218 524382 345454
rect 523826 344898 524062 345134
rect 524146 344898 524382 345134
rect 523826 309218 524062 309454
rect 524146 309218 524382 309454
rect 523826 308898 524062 309134
rect 524146 308898 524382 309134
rect 523826 273218 524062 273454
rect 524146 273218 524382 273454
rect 523826 272898 524062 273134
rect 524146 272898 524382 273134
rect 523826 237218 524062 237454
rect 524146 237218 524382 237454
rect 523826 236898 524062 237134
rect 524146 236898 524382 237134
rect 523826 201218 524062 201454
rect 524146 201218 524382 201454
rect 523826 200898 524062 201134
rect 524146 200898 524382 201134
rect 523826 165218 524062 165454
rect 524146 165218 524382 165454
rect 523826 164898 524062 165134
rect 524146 164898 524382 165134
rect 523826 129218 524062 129454
rect 524146 129218 524382 129454
rect 523826 128898 524062 129134
rect 524146 128898 524382 129134
rect 523826 93218 524062 93454
rect 524146 93218 524382 93454
rect 523826 92898 524062 93134
rect 524146 92898 524382 93134
rect 523826 57218 524062 57454
rect 524146 57218 524382 57454
rect 523826 56898 524062 57134
rect 524146 56898 524382 57134
rect 523826 21218 524062 21454
rect 524146 21218 524382 21454
rect 523826 20898 524062 21134
rect 524146 20898 524382 21134
rect 523826 -4422 524062 -4186
rect 524146 -4422 524382 -4186
rect 523826 -4742 524062 -4506
rect 524146 -4742 524382 -4506
rect 528326 709402 528562 709638
rect 528646 709402 528882 709638
rect 528326 709082 528562 709318
rect 528646 709082 528882 709318
rect 528326 673718 528562 673954
rect 528646 673718 528882 673954
rect 528326 673398 528562 673634
rect 528646 673398 528882 673634
rect 528326 637718 528562 637954
rect 528646 637718 528882 637954
rect 528326 637398 528562 637634
rect 528646 637398 528882 637634
rect 528326 601718 528562 601954
rect 528646 601718 528882 601954
rect 528326 601398 528562 601634
rect 528646 601398 528882 601634
rect 528326 565718 528562 565954
rect 528646 565718 528882 565954
rect 528326 565398 528562 565634
rect 528646 565398 528882 565634
rect 528326 529718 528562 529954
rect 528646 529718 528882 529954
rect 528326 529398 528562 529634
rect 528646 529398 528882 529634
rect 528326 493718 528562 493954
rect 528646 493718 528882 493954
rect 528326 493398 528562 493634
rect 528646 493398 528882 493634
rect 528326 457718 528562 457954
rect 528646 457718 528882 457954
rect 528326 457398 528562 457634
rect 528646 457398 528882 457634
rect 528326 421718 528562 421954
rect 528646 421718 528882 421954
rect 528326 421398 528562 421634
rect 528646 421398 528882 421634
rect 528326 385718 528562 385954
rect 528646 385718 528882 385954
rect 528326 385398 528562 385634
rect 528646 385398 528882 385634
rect 528326 349718 528562 349954
rect 528646 349718 528882 349954
rect 528326 349398 528562 349634
rect 528646 349398 528882 349634
rect 528326 313718 528562 313954
rect 528646 313718 528882 313954
rect 528326 313398 528562 313634
rect 528646 313398 528882 313634
rect 528326 277718 528562 277954
rect 528646 277718 528882 277954
rect 528326 277398 528562 277634
rect 528646 277398 528882 277634
rect 528326 241718 528562 241954
rect 528646 241718 528882 241954
rect 528326 241398 528562 241634
rect 528646 241398 528882 241634
rect 528326 205718 528562 205954
rect 528646 205718 528882 205954
rect 528326 205398 528562 205634
rect 528646 205398 528882 205634
rect 528326 169718 528562 169954
rect 528646 169718 528882 169954
rect 528326 169398 528562 169634
rect 528646 169398 528882 169634
rect 528326 133718 528562 133954
rect 528646 133718 528882 133954
rect 528326 133398 528562 133634
rect 528646 133398 528882 133634
rect 528326 97718 528562 97954
rect 528646 97718 528882 97954
rect 528326 97398 528562 97634
rect 528646 97398 528882 97634
rect 528326 61718 528562 61954
rect 528646 61718 528882 61954
rect 528326 61398 528562 61634
rect 528646 61398 528882 61634
rect 528326 25718 528562 25954
rect 528646 25718 528882 25954
rect 528326 25398 528562 25634
rect 528646 25398 528882 25634
rect 528326 -5382 528562 -5146
rect 528646 -5382 528882 -5146
rect 528326 -5702 528562 -5466
rect 528646 -5702 528882 -5466
rect 532826 710362 533062 710598
rect 533146 710362 533382 710598
rect 532826 710042 533062 710278
rect 533146 710042 533382 710278
rect 532826 678218 533062 678454
rect 533146 678218 533382 678454
rect 532826 677898 533062 678134
rect 533146 677898 533382 678134
rect 532826 642218 533062 642454
rect 533146 642218 533382 642454
rect 532826 641898 533062 642134
rect 533146 641898 533382 642134
rect 532826 606218 533062 606454
rect 533146 606218 533382 606454
rect 532826 605898 533062 606134
rect 533146 605898 533382 606134
rect 532826 570218 533062 570454
rect 533146 570218 533382 570454
rect 532826 569898 533062 570134
rect 533146 569898 533382 570134
rect 532826 534218 533062 534454
rect 533146 534218 533382 534454
rect 532826 533898 533062 534134
rect 533146 533898 533382 534134
rect 532826 498218 533062 498454
rect 533146 498218 533382 498454
rect 532826 497898 533062 498134
rect 533146 497898 533382 498134
rect 532826 462218 533062 462454
rect 533146 462218 533382 462454
rect 532826 461898 533062 462134
rect 533146 461898 533382 462134
rect 532826 426218 533062 426454
rect 533146 426218 533382 426454
rect 532826 425898 533062 426134
rect 533146 425898 533382 426134
rect 532826 390218 533062 390454
rect 533146 390218 533382 390454
rect 532826 389898 533062 390134
rect 533146 389898 533382 390134
rect 532826 354218 533062 354454
rect 533146 354218 533382 354454
rect 532826 353898 533062 354134
rect 533146 353898 533382 354134
rect 532826 318218 533062 318454
rect 533146 318218 533382 318454
rect 532826 317898 533062 318134
rect 533146 317898 533382 318134
rect 532826 282218 533062 282454
rect 533146 282218 533382 282454
rect 532826 281898 533062 282134
rect 533146 281898 533382 282134
rect 532826 246218 533062 246454
rect 533146 246218 533382 246454
rect 532826 245898 533062 246134
rect 533146 245898 533382 246134
rect 532826 210218 533062 210454
rect 533146 210218 533382 210454
rect 532826 209898 533062 210134
rect 533146 209898 533382 210134
rect 532826 174218 533062 174454
rect 533146 174218 533382 174454
rect 532826 173898 533062 174134
rect 533146 173898 533382 174134
rect 532826 138218 533062 138454
rect 533146 138218 533382 138454
rect 532826 137898 533062 138134
rect 533146 137898 533382 138134
rect 532826 102218 533062 102454
rect 533146 102218 533382 102454
rect 532826 101898 533062 102134
rect 533146 101898 533382 102134
rect 532826 66218 533062 66454
rect 533146 66218 533382 66454
rect 532826 65898 533062 66134
rect 533146 65898 533382 66134
rect 532826 30218 533062 30454
rect 533146 30218 533382 30454
rect 532826 29898 533062 30134
rect 533146 29898 533382 30134
rect 532826 -6342 533062 -6106
rect 533146 -6342 533382 -6106
rect 532826 -6662 533062 -6426
rect 533146 -6662 533382 -6426
rect 537326 711322 537562 711558
rect 537646 711322 537882 711558
rect 537326 711002 537562 711238
rect 537646 711002 537882 711238
rect 537326 682718 537562 682954
rect 537646 682718 537882 682954
rect 537326 682398 537562 682634
rect 537646 682398 537882 682634
rect 537326 646718 537562 646954
rect 537646 646718 537882 646954
rect 537326 646398 537562 646634
rect 537646 646398 537882 646634
rect 537326 610718 537562 610954
rect 537646 610718 537882 610954
rect 537326 610398 537562 610634
rect 537646 610398 537882 610634
rect 537326 574718 537562 574954
rect 537646 574718 537882 574954
rect 537326 574398 537562 574634
rect 537646 574398 537882 574634
rect 537326 538718 537562 538954
rect 537646 538718 537882 538954
rect 537326 538398 537562 538634
rect 537646 538398 537882 538634
rect 537326 502718 537562 502954
rect 537646 502718 537882 502954
rect 537326 502398 537562 502634
rect 537646 502398 537882 502634
rect 537326 466718 537562 466954
rect 537646 466718 537882 466954
rect 537326 466398 537562 466634
rect 537646 466398 537882 466634
rect 537326 430718 537562 430954
rect 537646 430718 537882 430954
rect 537326 430398 537562 430634
rect 537646 430398 537882 430634
rect 537326 394718 537562 394954
rect 537646 394718 537882 394954
rect 537326 394398 537562 394634
rect 537646 394398 537882 394634
rect 537326 358718 537562 358954
rect 537646 358718 537882 358954
rect 537326 358398 537562 358634
rect 537646 358398 537882 358634
rect 537326 322718 537562 322954
rect 537646 322718 537882 322954
rect 537326 322398 537562 322634
rect 537646 322398 537882 322634
rect 537326 286718 537562 286954
rect 537646 286718 537882 286954
rect 537326 286398 537562 286634
rect 537646 286398 537882 286634
rect 537326 250718 537562 250954
rect 537646 250718 537882 250954
rect 537326 250398 537562 250634
rect 537646 250398 537882 250634
rect 537326 214718 537562 214954
rect 537646 214718 537882 214954
rect 537326 214398 537562 214634
rect 537646 214398 537882 214634
rect 537326 178718 537562 178954
rect 537646 178718 537882 178954
rect 537326 178398 537562 178634
rect 537646 178398 537882 178634
rect 537326 142718 537562 142954
rect 537646 142718 537882 142954
rect 537326 142398 537562 142634
rect 537646 142398 537882 142634
rect 537326 106718 537562 106954
rect 537646 106718 537882 106954
rect 537326 106398 537562 106634
rect 537646 106398 537882 106634
rect 537326 70718 537562 70954
rect 537646 70718 537882 70954
rect 537326 70398 537562 70634
rect 537646 70398 537882 70634
rect 537326 34718 537562 34954
rect 537646 34718 537882 34954
rect 537326 34398 537562 34634
rect 537646 34398 537882 34634
rect 537326 -7302 537562 -7066
rect 537646 -7302 537882 -7066
rect 537326 -7622 537562 -7386
rect 537646 -7622 537882 -7386
rect 541826 704602 542062 704838
rect 542146 704602 542382 704838
rect 541826 704282 542062 704518
rect 542146 704282 542382 704518
rect 541826 687218 542062 687454
rect 542146 687218 542382 687454
rect 541826 686898 542062 687134
rect 542146 686898 542382 687134
rect 541826 651218 542062 651454
rect 542146 651218 542382 651454
rect 541826 650898 542062 651134
rect 542146 650898 542382 651134
rect 541826 615218 542062 615454
rect 542146 615218 542382 615454
rect 541826 614898 542062 615134
rect 542146 614898 542382 615134
rect 541826 579218 542062 579454
rect 542146 579218 542382 579454
rect 541826 578898 542062 579134
rect 542146 578898 542382 579134
rect 541826 543218 542062 543454
rect 542146 543218 542382 543454
rect 541826 542898 542062 543134
rect 542146 542898 542382 543134
rect 541826 507218 542062 507454
rect 542146 507218 542382 507454
rect 541826 506898 542062 507134
rect 542146 506898 542382 507134
rect 541826 471218 542062 471454
rect 542146 471218 542382 471454
rect 541826 470898 542062 471134
rect 542146 470898 542382 471134
rect 541826 435218 542062 435454
rect 542146 435218 542382 435454
rect 541826 434898 542062 435134
rect 542146 434898 542382 435134
rect 541826 399218 542062 399454
rect 542146 399218 542382 399454
rect 541826 398898 542062 399134
rect 542146 398898 542382 399134
rect 541826 363218 542062 363454
rect 542146 363218 542382 363454
rect 541826 362898 542062 363134
rect 542146 362898 542382 363134
rect 541826 327218 542062 327454
rect 542146 327218 542382 327454
rect 541826 326898 542062 327134
rect 542146 326898 542382 327134
rect 541826 291218 542062 291454
rect 542146 291218 542382 291454
rect 541826 290898 542062 291134
rect 542146 290898 542382 291134
rect 541826 255218 542062 255454
rect 542146 255218 542382 255454
rect 541826 254898 542062 255134
rect 542146 254898 542382 255134
rect 541826 219218 542062 219454
rect 542146 219218 542382 219454
rect 541826 218898 542062 219134
rect 542146 218898 542382 219134
rect 541826 183218 542062 183454
rect 542146 183218 542382 183454
rect 541826 182898 542062 183134
rect 542146 182898 542382 183134
rect 541826 147218 542062 147454
rect 542146 147218 542382 147454
rect 541826 146898 542062 147134
rect 542146 146898 542382 147134
rect 541826 111218 542062 111454
rect 542146 111218 542382 111454
rect 541826 110898 542062 111134
rect 542146 110898 542382 111134
rect 541826 75218 542062 75454
rect 542146 75218 542382 75454
rect 541826 74898 542062 75134
rect 542146 74898 542382 75134
rect 541826 39218 542062 39454
rect 542146 39218 542382 39454
rect 541826 38898 542062 39134
rect 542146 38898 542382 39134
rect 541826 3218 542062 3454
rect 542146 3218 542382 3454
rect 541826 2898 542062 3134
rect 542146 2898 542382 3134
rect 541826 -582 542062 -346
rect 542146 -582 542382 -346
rect 541826 -902 542062 -666
rect 542146 -902 542382 -666
rect 546326 705562 546562 705798
rect 546646 705562 546882 705798
rect 546326 705242 546562 705478
rect 546646 705242 546882 705478
rect 546326 691718 546562 691954
rect 546646 691718 546882 691954
rect 546326 691398 546562 691634
rect 546646 691398 546882 691634
rect 546326 655718 546562 655954
rect 546646 655718 546882 655954
rect 546326 655398 546562 655634
rect 546646 655398 546882 655634
rect 546326 619718 546562 619954
rect 546646 619718 546882 619954
rect 546326 619398 546562 619634
rect 546646 619398 546882 619634
rect 546326 583718 546562 583954
rect 546646 583718 546882 583954
rect 546326 583398 546562 583634
rect 546646 583398 546882 583634
rect 546326 547718 546562 547954
rect 546646 547718 546882 547954
rect 546326 547398 546562 547634
rect 546646 547398 546882 547634
rect 546326 511718 546562 511954
rect 546646 511718 546882 511954
rect 546326 511398 546562 511634
rect 546646 511398 546882 511634
rect 546326 475718 546562 475954
rect 546646 475718 546882 475954
rect 546326 475398 546562 475634
rect 546646 475398 546882 475634
rect 546326 439718 546562 439954
rect 546646 439718 546882 439954
rect 546326 439398 546562 439634
rect 546646 439398 546882 439634
rect 546326 403718 546562 403954
rect 546646 403718 546882 403954
rect 546326 403398 546562 403634
rect 546646 403398 546882 403634
rect 546326 367718 546562 367954
rect 546646 367718 546882 367954
rect 546326 367398 546562 367634
rect 546646 367398 546882 367634
rect 546326 331718 546562 331954
rect 546646 331718 546882 331954
rect 546326 331398 546562 331634
rect 546646 331398 546882 331634
rect 546326 295718 546562 295954
rect 546646 295718 546882 295954
rect 546326 295398 546562 295634
rect 546646 295398 546882 295634
rect 546326 259718 546562 259954
rect 546646 259718 546882 259954
rect 546326 259398 546562 259634
rect 546646 259398 546882 259634
rect 546326 223718 546562 223954
rect 546646 223718 546882 223954
rect 546326 223398 546562 223634
rect 546646 223398 546882 223634
rect 546326 187718 546562 187954
rect 546646 187718 546882 187954
rect 546326 187398 546562 187634
rect 546646 187398 546882 187634
rect 546326 151718 546562 151954
rect 546646 151718 546882 151954
rect 546326 151398 546562 151634
rect 546646 151398 546882 151634
rect 546326 115718 546562 115954
rect 546646 115718 546882 115954
rect 546326 115398 546562 115634
rect 546646 115398 546882 115634
rect 546326 79718 546562 79954
rect 546646 79718 546882 79954
rect 546326 79398 546562 79634
rect 546646 79398 546882 79634
rect 546326 43718 546562 43954
rect 546646 43718 546882 43954
rect 546326 43398 546562 43634
rect 546646 43398 546882 43634
rect 546326 7718 546562 7954
rect 546646 7718 546882 7954
rect 546326 7398 546562 7634
rect 546646 7398 546882 7634
rect 546326 -1542 546562 -1306
rect 546646 -1542 546882 -1306
rect 546326 -1862 546562 -1626
rect 546646 -1862 546882 -1626
rect 550826 706522 551062 706758
rect 551146 706522 551382 706758
rect 550826 706202 551062 706438
rect 551146 706202 551382 706438
rect 550826 696218 551062 696454
rect 551146 696218 551382 696454
rect 550826 695898 551062 696134
rect 551146 695898 551382 696134
rect 550826 660218 551062 660454
rect 551146 660218 551382 660454
rect 550826 659898 551062 660134
rect 551146 659898 551382 660134
rect 550826 624218 551062 624454
rect 551146 624218 551382 624454
rect 550826 623898 551062 624134
rect 551146 623898 551382 624134
rect 550826 588218 551062 588454
rect 551146 588218 551382 588454
rect 550826 587898 551062 588134
rect 551146 587898 551382 588134
rect 550826 552218 551062 552454
rect 551146 552218 551382 552454
rect 550826 551898 551062 552134
rect 551146 551898 551382 552134
rect 550826 516218 551062 516454
rect 551146 516218 551382 516454
rect 550826 515898 551062 516134
rect 551146 515898 551382 516134
rect 550826 480218 551062 480454
rect 551146 480218 551382 480454
rect 550826 479898 551062 480134
rect 551146 479898 551382 480134
rect 550826 444218 551062 444454
rect 551146 444218 551382 444454
rect 550826 443898 551062 444134
rect 551146 443898 551382 444134
rect 550826 408218 551062 408454
rect 551146 408218 551382 408454
rect 550826 407898 551062 408134
rect 551146 407898 551382 408134
rect 550826 372218 551062 372454
rect 551146 372218 551382 372454
rect 550826 371898 551062 372134
rect 551146 371898 551382 372134
rect 550826 336218 551062 336454
rect 551146 336218 551382 336454
rect 550826 335898 551062 336134
rect 551146 335898 551382 336134
rect 550826 300218 551062 300454
rect 551146 300218 551382 300454
rect 550826 299898 551062 300134
rect 551146 299898 551382 300134
rect 550826 264218 551062 264454
rect 551146 264218 551382 264454
rect 550826 263898 551062 264134
rect 551146 263898 551382 264134
rect 550826 228218 551062 228454
rect 551146 228218 551382 228454
rect 550826 227898 551062 228134
rect 551146 227898 551382 228134
rect 550826 192218 551062 192454
rect 551146 192218 551382 192454
rect 550826 191898 551062 192134
rect 551146 191898 551382 192134
rect 550826 156218 551062 156454
rect 551146 156218 551382 156454
rect 550826 155898 551062 156134
rect 551146 155898 551382 156134
rect 550826 120218 551062 120454
rect 551146 120218 551382 120454
rect 550826 119898 551062 120134
rect 551146 119898 551382 120134
rect 550826 84218 551062 84454
rect 551146 84218 551382 84454
rect 550826 83898 551062 84134
rect 551146 83898 551382 84134
rect 550826 48218 551062 48454
rect 551146 48218 551382 48454
rect 550826 47898 551062 48134
rect 551146 47898 551382 48134
rect 550826 12218 551062 12454
rect 551146 12218 551382 12454
rect 550826 11898 551062 12134
rect 551146 11898 551382 12134
rect 550826 -2502 551062 -2266
rect 551146 -2502 551382 -2266
rect 550826 -2822 551062 -2586
rect 551146 -2822 551382 -2586
rect 555326 707482 555562 707718
rect 555646 707482 555882 707718
rect 555326 707162 555562 707398
rect 555646 707162 555882 707398
rect 555326 700718 555562 700954
rect 555646 700718 555882 700954
rect 555326 700398 555562 700634
rect 555646 700398 555882 700634
rect 555326 664718 555562 664954
rect 555646 664718 555882 664954
rect 555326 664398 555562 664634
rect 555646 664398 555882 664634
rect 555326 628718 555562 628954
rect 555646 628718 555882 628954
rect 555326 628398 555562 628634
rect 555646 628398 555882 628634
rect 555326 592718 555562 592954
rect 555646 592718 555882 592954
rect 555326 592398 555562 592634
rect 555646 592398 555882 592634
rect 555326 556718 555562 556954
rect 555646 556718 555882 556954
rect 555326 556398 555562 556634
rect 555646 556398 555882 556634
rect 555326 520718 555562 520954
rect 555646 520718 555882 520954
rect 555326 520398 555562 520634
rect 555646 520398 555882 520634
rect 555326 484718 555562 484954
rect 555646 484718 555882 484954
rect 555326 484398 555562 484634
rect 555646 484398 555882 484634
rect 555326 448718 555562 448954
rect 555646 448718 555882 448954
rect 555326 448398 555562 448634
rect 555646 448398 555882 448634
rect 555326 412718 555562 412954
rect 555646 412718 555882 412954
rect 555326 412398 555562 412634
rect 555646 412398 555882 412634
rect 555326 376718 555562 376954
rect 555646 376718 555882 376954
rect 555326 376398 555562 376634
rect 555646 376398 555882 376634
rect 555326 340718 555562 340954
rect 555646 340718 555882 340954
rect 555326 340398 555562 340634
rect 555646 340398 555882 340634
rect 555326 304718 555562 304954
rect 555646 304718 555882 304954
rect 555326 304398 555562 304634
rect 555646 304398 555882 304634
rect 555326 268718 555562 268954
rect 555646 268718 555882 268954
rect 555326 268398 555562 268634
rect 555646 268398 555882 268634
rect 555326 232718 555562 232954
rect 555646 232718 555882 232954
rect 555326 232398 555562 232634
rect 555646 232398 555882 232634
rect 555326 196718 555562 196954
rect 555646 196718 555882 196954
rect 555326 196398 555562 196634
rect 555646 196398 555882 196634
rect 555326 160718 555562 160954
rect 555646 160718 555882 160954
rect 555326 160398 555562 160634
rect 555646 160398 555882 160634
rect 555326 124718 555562 124954
rect 555646 124718 555882 124954
rect 555326 124398 555562 124634
rect 555646 124398 555882 124634
rect 555326 88718 555562 88954
rect 555646 88718 555882 88954
rect 555326 88398 555562 88634
rect 555646 88398 555882 88634
rect 555326 52718 555562 52954
rect 555646 52718 555882 52954
rect 555326 52398 555562 52634
rect 555646 52398 555882 52634
rect 555326 16718 555562 16954
rect 555646 16718 555882 16954
rect 555326 16398 555562 16634
rect 555646 16398 555882 16634
rect 555326 -3462 555562 -3226
rect 555646 -3462 555882 -3226
rect 555326 -3782 555562 -3546
rect 555646 -3782 555882 -3546
rect 559826 708442 560062 708678
rect 560146 708442 560382 708678
rect 559826 708122 560062 708358
rect 560146 708122 560382 708358
rect 559826 669218 560062 669454
rect 560146 669218 560382 669454
rect 559826 668898 560062 669134
rect 560146 668898 560382 669134
rect 559826 633218 560062 633454
rect 560146 633218 560382 633454
rect 559826 632898 560062 633134
rect 560146 632898 560382 633134
rect 559826 597218 560062 597454
rect 560146 597218 560382 597454
rect 559826 596898 560062 597134
rect 560146 596898 560382 597134
rect 559826 561218 560062 561454
rect 560146 561218 560382 561454
rect 559826 560898 560062 561134
rect 560146 560898 560382 561134
rect 559826 525218 560062 525454
rect 560146 525218 560382 525454
rect 559826 524898 560062 525134
rect 560146 524898 560382 525134
rect 559826 489218 560062 489454
rect 560146 489218 560382 489454
rect 559826 488898 560062 489134
rect 560146 488898 560382 489134
rect 559826 453218 560062 453454
rect 560146 453218 560382 453454
rect 559826 452898 560062 453134
rect 560146 452898 560382 453134
rect 559826 417218 560062 417454
rect 560146 417218 560382 417454
rect 559826 416898 560062 417134
rect 560146 416898 560382 417134
rect 559826 381218 560062 381454
rect 560146 381218 560382 381454
rect 559826 380898 560062 381134
rect 560146 380898 560382 381134
rect 559826 345218 560062 345454
rect 560146 345218 560382 345454
rect 559826 344898 560062 345134
rect 560146 344898 560382 345134
rect 559826 309218 560062 309454
rect 560146 309218 560382 309454
rect 559826 308898 560062 309134
rect 560146 308898 560382 309134
rect 559826 273218 560062 273454
rect 560146 273218 560382 273454
rect 559826 272898 560062 273134
rect 560146 272898 560382 273134
rect 559826 237218 560062 237454
rect 560146 237218 560382 237454
rect 559826 236898 560062 237134
rect 560146 236898 560382 237134
rect 559826 201218 560062 201454
rect 560146 201218 560382 201454
rect 559826 200898 560062 201134
rect 560146 200898 560382 201134
rect 559826 165218 560062 165454
rect 560146 165218 560382 165454
rect 559826 164898 560062 165134
rect 560146 164898 560382 165134
rect 559826 129218 560062 129454
rect 560146 129218 560382 129454
rect 559826 128898 560062 129134
rect 560146 128898 560382 129134
rect 559826 93218 560062 93454
rect 560146 93218 560382 93454
rect 559826 92898 560062 93134
rect 560146 92898 560382 93134
rect 559826 57218 560062 57454
rect 560146 57218 560382 57454
rect 559826 56898 560062 57134
rect 560146 56898 560382 57134
rect 559826 21218 560062 21454
rect 560146 21218 560382 21454
rect 559826 20898 560062 21134
rect 560146 20898 560382 21134
rect 559826 -4422 560062 -4186
rect 560146 -4422 560382 -4186
rect 559826 -4742 560062 -4506
rect 560146 -4742 560382 -4506
rect 564326 709402 564562 709638
rect 564646 709402 564882 709638
rect 564326 709082 564562 709318
rect 564646 709082 564882 709318
rect 564326 673718 564562 673954
rect 564646 673718 564882 673954
rect 564326 673398 564562 673634
rect 564646 673398 564882 673634
rect 564326 637718 564562 637954
rect 564646 637718 564882 637954
rect 564326 637398 564562 637634
rect 564646 637398 564882 637634
rect 564326 601718 564562 601954
rect 564646 601718 564882 601954
rect 564326 601398 564562 601634
rect 564646 601398 564882 601634
rect 564326 565718 564562 565954
rect 564646 565718 564882 565954
rect 564326 565398 564562 565634
rect 564646 565398 564882 565634
rect 564326 529718 564562 529954
rect 564646 529718 564882 529954
rect 564326 529398 564562 529634
rect 564646 529398 564882 529634
rect 564326 493718 564562 493954
rect 564646 493718 564882 493954
rect 564326 493398 564562 493634
rect 564646 493398 564882 493634
rect 564326 457718 564562 457954
rect 564646 457718 564882 457954
rect 564326 457398 564562 457634
rect 564646 457398 564882 457634
rect 564326 421718 564562 421954
rect 564646 421718 564882 421954
rect 564326 421398 564562 421634
rect 564646 421398 564882 421634
rect 564326 385718 564562 385954
rect 564646 385718 564882 385954
rect 564326 385398 564562 385634
rect 564646 385398 564882 385634
rect 564326 349718 564562 349954
rect 564646 349718 564882 349954
rect 564326 349398 564562 349634
rect 564646 349398 564882 349634
rect 564326 313718 564562 313954
rect 564646 313718 564882 313954
rect 564326 313398 564562 313634
rect 564646 313398 564882 313634
rect 564326 277718 564562 277954
rect 564646 277718 564882 277954
rect 564326 277398 564562 277634
rect 564646 277398 564882 277634
rect 564326 241718 564562 241954
rect 564646 241718 564882 241954
rect 564326 241398 564562 241634
rect 564646 241398 564882 241634
rect 564326 205718 564562 205954
rect 564646 205718 564882 205954
rect 564326 205398 564562 205634
rect 564646 205398 564882 205634
rect 564326 169718 564562 169954
rect 564646 169718 564882 169954
rect 564326 169398 564562 169634
rect 564646 169398 564882 169634
rect 564326 133718 564562 133954
rect 564646 133718 564882 133954
rect 564326 133398 564562 133634
rect 564646 133398 564882 133634
rect 564326 97718 564562 97954
rect 564646 97718 564882 97954
rect 564326 97398 564562 97634
rect 564646 97398 564882 97634
rect 564326 61718 564562 61954
rect 564646 61718 564882 61954
rect 564326 61398 564562 61634
rect 564646 61398 564882 61634
rect 564326 25718 564562 25954
rect 564646 25718 564882 25954
rect 564326 25398 564562 25634
rect 564646 25398 564882 25634
rect 564326 -5382 564562 -5146
rect 564646 -5382 564882 -5146
rect 564326 -5702 564562 -5466
rect 564646 -5702 564882 -5466
rect 568826 710362 569062 710598
rect 569146 710362 569382 710598
rect 568826 710042 569062 710278
rect 569146 710042 569382 710278
rect 568826 678218 569062 678454
rect 569146 678218 569382 678454
rect 568826 677898 569062 678134
rect 569146 677898 569382 678134
rect 568826 642218 569062 642454
rect 569146 642218 569382 642454
rect 568826 641898 569062 642134
rect 569146 641898 569382 642134
rect 568826 606218 569062 606454
rect 569146 606218 569382 606454
rect 568826 605898 569062 606134
rect 569146 605898 569382 606134
rect 568826 570218 569062 570454
rect 569146 570218 569382 570454
rect 568826 569898 569062 570134
rect 569146 569898 569382 570134
rect 568826 534218 569062 534454
rect 569146 534218 569382 534454
rect 568826 533898 569062 534134
rect 569146 533898 569382 534134
rect 568826 498218 569062 498454
rect 569146 498218 569382 498454
rect 568826 497898 569062 498134
rect 569146 497898 569382 498134
rect 568826 462218 569062 462454
rect 569146 462218 569382 462454
rect 568826 461898 569062 462134
rect 569146 461898 569382 462134
rect 568826 426218 569062 426454
rect 569146 426218 569382 426454
rect 568826 425898 569062 426134
rect 569146 425898 569382 426134
rect 568826 390218 569062 390454
rect 569146 390218 569382 390454
rect 568826 389898 569062 390134
rect 569146 389898 569382 390134
rect 568826 354218 569062 354454
rect 569146 354218 569382 354454
rect 568826 353898 569062 354134
rect 569146 353898 569382 354134
rect 568826 318218 569062 318454
rect 569146 318218 569382 318454
rect 568826 317898 569062 318134
rect 569146 317898 569382 318134
rect 568826 282218 569062 282454
rect 569146 282218 569382 282454
rect 568826 281898 569062 282134
rect 569146 281898 569382 282134
rect 568826 246218 569062 246454
rect 569146 246218 569382 246454
rect 568826 245898 569062 246134
rect 569146 245898 569382 246134
rect 568826 210218 569062 210454
rect 569146 210218 569382 210454
rect 568826 209898 569062 210134
rect 569146 209898 569382 210134
rect 568826 174218 569062 174454
rect 569146 174218 569382 174454
rect 568826 173898 569062 174134
rect 569146 173898 569382 174134
rect 568826 138218 569062 138454
rect 569146 138218 569382 138454
rect 568826 137898 569062 138134
rect 569146 137898 569382 138134
rect 568826 102218 569062 102454
rect 569146 102218 569382 102454
rect 568826 101898 569062 102134
rect 569146 101898 569382 102134
rect 568826 66218 569062 66454
rect 569146 66218 569382 66454
rect 568826 65898 569062 66134
rect 569146 65898 569382 66134
rect 568826 30218 569062 30454
rect 569146 30218 569382 30454
rect 568826 29898 569062 30134
rect 569146 29898 569382 30134
rect 568826 -6342 569062 -6106
rect 569146 -6342 569382 -6106
rect 568826 -6662 569062 -6426
rect 569146 -6662 569382 -6426
rect 573326 711322 573562 711558
rect 573646 711322 573882 711558
rect 573326 711002 573562 711238
rect 573646 711002 573882 711238
rect 573326 682718 573562 682954
rect 573646 682718 573882 682954
rect 573326 682398 573562 682634
rect 573646 682398 573882 682634
rect 573326 646718 573562 646954
rect 573646 646718 573882 646954
rect 573326 646398 573562 646634
rect 573646 646398 573882 646634
rect 573326 610718 573562 610954
rect 573646 610718 573882 610954
rect 573326 610398 573562 610634
rect 573646 610398 573882 610634
rect 573326 574718 573562 574954
rect 573646 574718 573882 574954
rect 573326 574398 573562 574634
rect 573646 574398 573882 574634
rect 573326 538718 573562 538954
rect 573646 538718 573882 538954
rect 573326 538398 573562 538634
rect 573646 538398 573882 538634
rect 573326 502718 573562 502954
rect 573646 502718 573882 502954
rect 573326 502398 573562 502634
rect 573646 502398 573882 502634
rect 573326 466718 573562 466954
rect 573646 466718 573882 466954
rect 573326 466398 573562 466634
rect 573646 466398 573882 466634
rect 573326 430718 573562 430954
rect 573646 430718 573882 430954
rect 573326 430398 573562 430634
rect 573646 430398 573882 430634
rect 573326 394718 573562 394954
rect 573646 394718 573882 394954
rect 573326 394398 573562 394634
rect 573646 394398 573882 394634
rect 573326 358718 573562 358954
rect 573646 358718 573882 358954
rect 573326 358398 573562 358634
rect 573646 358398 573882 358634
rect 573326 322718 573562 322954
rect 573646 322718 573882 322954
rect 573326 322398 573562 322634
rect 573646 322398 573882 322634
rect 573326 286718 573562 286954
rect 573646 286718 573882 286954
rect 573326 286398 573562 286634
rect 573646 286398 573882 286634
rect 573326 250718 573562 250954
rect 573646 250718 573882 250954
rect 573326 250398 573562 250634
rect 573646 250398 573882 250634
rect 573326 214718 573562 214954
rect 573646 214718 573882 214954
rect 573326 214398 573562 214634
rect 573646 214398 573882 214634
rect 573326 178718 573562 178954
rect 573646 178718 573882 178954
rect 573326 178398 573562 178634
rect 573646 178398 573882 178634
rect 573326 142718 573562 142954
rect 573646 142718 573882 142954
rect 573326 142398 573562 142634
rect 573646 142398 573882 142634
rect 573326 106718 573562 106954
rect 573646 106718 573882 106954
rect 573326 106398 573562 106634
rect 573646 106398 573882 106634
rect 573326 70718 573562 70954
rect 573646 70718 573882 70954
rect 573326 70398 573562 70634
rect 573646 70398 573882 70634
rect 573326 34718 573562 34954
rect 573646 34718 573882 34954
rect 573326 34398 573562 34634
rect 573646 34398 573882 34634
rect 573326 -7302 573562 -7066
rect 573646 -7302 573882 -7066
rect 573326 -7622 573562 -7386
rect 573646 -7622 573882 -7386
rect 577826 704602 578062 704838
rect 578146 704602 578382 704838
rect 577826 704282 578062 704518
rect 578146 704282 578382 704518
rect 577826 687218 578062 687454
rect 578146 687218 578382 687454
rect 577826 686898 578062 687134
rect 578146 686898 578382 687134
rect 577826 651218 578062 651454
rect 578146 651218 578382 651454
rect 577826 650898 578062 651134
rect 578146 650898 578382 651134
rect 577826 615218 578062 615454
rect 578146 615218 578382 615454
rect 577826 614898 578062 615134
rect 578146 614898 578382 615134
rect 577826 579218 578062 579454
rect 578146 579218 578382 579454
rect 577826 578898 578062 579134
rect 578146 578898 578382 579134
rect 577826 543218 578062 543454
rect 578146 543218 578382 543454
rect 577826 542898 578062 543134
rect 578146 542898 578382 543134
rect 577826 507218 578062 507454
rect 578146 507218 578382 507454
rect 577826 506898 578062 507134
rect 578146 506898 578382 507134
rect 577826 471218 578062 471454
rect 578146 471218 578382 471454
rect 577826 470898 578062 471134
rect 578146 470898 578382 471134
rect 577826 435218 578062 435454
rect 578146 435218 578382 435454
rect 577826 434898 578062 435134
rect 578146 434898 578382 435134
rect 577826 399218 578062 399454
rect 578146 399218 578382 399454
rect 577826 398898 578062 399134
rect 578146 398898 578382 399134
rect 577826 363218 578062 363454
rect 578146 363218 578382 363454
rect 577826 362898 578062 363134
rect 578146 362898 578382 363134
rect 577826 327218 578062 327454
rect 578146 327218 578382 327454
rect 577826 326898 578062 327134
rect 578146 326898 578382 327134
rect 577826 291218 578062 291454
rect 578146 291218 578382 291454
rect 577826 290898 578062 291134
rect 578146 290898 578382 291134
rect 577826 255218 578062 255454
rect 578146 255218 578382 255454
rect 577826 254898 578062 255134
rect 578146 254898 578382 255134
rect 577826 219218 578062 219454
rect 578146 219218 578382 219454
rect 577826 218898 578062 219134
rect 578146 218898 578382 219134
rect 577826 183218 578062 183454
rect 578146 183218 578382 183454
rect 577826 182898 578062 183134
rect 578146 182898 578382 183134
rect 577826 147218 578062 147454
rect 578146 147218 578382 147454
rect 577826 146898 578062 147134
rect 578146 146898 578382 147134
rect 577826 111218 578062 111454
rect 578146 111218 578382 111454
rect 577826 110898 578062 111134
rect 578146 110898 578382 111134
rect 577826 75218 578062 75454
rect 578146 75218 578382 75454
rect 577826 74898 578062 75134
rect 578146 74898 578382 75134
rect 577826 39218 578062 39454
rect 578146 39218 578382 39454
rect 577826 38898 578062 39134
rect 578146 38898 578382 39134
rect 577826 3218 578062 3454
rect 578146 3218 578382 3454
rect 577826 2898 578062 3134
rect 578146 2898 578382 3134
rect 577826 -582 578062 -346
rect 578146 -582 578382 -346
rect 577826 -902 578062 -666
rect 578146 -902 578382 -666
rect 592062 711322 592298 711558
rect 592382 711322 592618 711558
rect 592062 711002 592298 711238
rect 592382 711002 592618 711238
rect 591102 710362 591338 710598
rect 591422 710362 591658 710598
rect 591102 710042 591338 710278
rect 591422 710042 591658 710278
rect 590142 709402 590378 709638
rect 590462 709402 590698 709638
rect 590142 709082 590378 709318
rect 590462 709082 590698 709318
rect 589182 708442 589418 708678
rect 589502 708442 589738 708678
rect 589182 708122 589418 708358
rect 589502 708122 589738 708358
rect 588222 707482 588458 707718
rect 588542 707482 588778 707718
rect 588222 707162 588458 707398
rect 588542 707162 588778 707398
rect 587262 706522 587498 706758
rect 587582 706522 587818 706758
rect 587262 706202 587498 706438
rect 587582 706202 587818 706438
rect 582326 705562 582562 705798
rect 582646 705562 582882 705798
rect 582326 705242 582562 705478
rect 582646 705242 582882 705478
rect 586302 705562 586538 705798
rect 586622 705562 586858 705798
rect 586302 705242 586538 705478
rect 586622 705242 586858 705478
rect 582326 691718 582562 691954
rect 582646 691718 582882 691954
rect 582326 691398 582562 691634
rect 582646 691398 582882 691634
rect 582326 655718 582562 655954
rect 582646 655718 582882 655954
rect 582326 655398 582562 655634
rect 582646 655398 582882 655634
rect 582326 619718 582562 619954
rect 582646 619718 582882 619954
rect 582326 619398 582562 619634
rect 582646 619398 582882 619634
rect 582326 583718 582562 583954
rect 582646 583718 582882 583954
rect 582326 583398 582562 583634
rect 582646 583398 582882 583634
rect 582326 547718 582562 547954
rect 582646 547718 582882 547954
rect 582326 547398 582562 547634
rect 582646 547398 582882 547634
rect 582326 511718 582562 511954
rect 582646 511718 582882 511954
rect 582326 511398 582562 511634
rect 582646 511398 582882 511634
rect 582326 475718 582562 475954
rect 582646 475718 582882 475954
rect 582326 475398 582562 475634
rect 582646 475398 582882 475634
rect 582326 439718 582562 439954
rect 582646 439718 582882 439954
rect 582326 439398 582562 439634
rect 582646 439398 582882 439634
rect 582326 403718 582562 403954
rect 582646 403718 582882 403954
rect 582326 403398 582562 403634
rect 582646 403398 582882 403634
rect 582326 367718 582562 367954
rect 582646 367718 582882 367954
rect 582326 367398 582562 367634
rect 582646 367398 582882 367634
rect 582326 331718 582562 331954
rect 582646 331718 582882 331954
rect 582326 331398 582562 331634
rect 582646 331398 582882 331634
rect 582326 295718 582562 295954
rect 582646 295718 582882 295954
rect 582326 295398 582562 295634
rect 582646 295398 582882 295634
rect 582326 259718 582562 259954
rect 582646 259718 582882 259954
rect 582326 259398 582562 259634
rect 582646 259398 582882 259634
rect 582326 223718 582562 223954
rect 582646 223718 582882 223954
rect 582326 223398 582562 223634
rect 582646 223398 582882 223634
rect 582326 187718 582562 187954
rect 582646 187718 582882 187954
rect 582326 187398 582562 187634
rect 582646 187398 582882 187634
rect 582326 151718 582562 151954
rect 582646 151718 582882 151954
rect 582326 151398 582562 151634
rect 582646 151398 582882 151634
rect 582326 115718 582562 115954
rect 582646 115718 582882 115954
rect 582326 115398 582562 115634
rect 582646 115398 582882 115634
rect 582326 79718 582562 79954
rect 582646 79718 582882 79954
rect 582326 79398 582562 79634
rect 582646 79398 582882 79634
rect 582326 43718 582562 43954
rect 582646 43718 582882 43954
rect 582326 43398 582562 43634
rect 582646 43398 582882 43634
rect 582326 7718 582562 7954
rect 582646 7718 582882 7954
rect 582326 7398 582562 7634
rect 582646 7398 582882 7634
rect 585342 704602 585578 704838
rect 585662 704602 585898 704838
rect 585342 704282 585578 704518
rect 585662 704282 585898 704518
rect 585342 687218 585578 687454
rect 585662 687218 585898 687454
rect 585342 686898 585578 687134
rect 585662 686898 585898 687134
rect 585342 651218 585578 651454
rect 585662 651218 585898 651454
rect 585342 650898 585578 651134
rect 585662 650898 585898 651134
rect 585342 615218 585578 615454
rect 585662 615218 585898 615454
rect 585342 614898 585578 615134
rect 585662 614898 585898 615134
rect 585342 579218 585578 579454
rect 585662 579218 585898 579454
rect 585342 578898 585578 579134
rect 585662 578898 585898 579134
rect 585342 543218 585578 543454
rect 585662 543218 585898 543454
rect 585342 542898 585578 543134
rect 585662 542898 585898 543134
rect 585342 507218 585578 507454
rect 585662 507218 585898 507454
rect 585342 506898 585578 507134
rect 585662 506898 585898 507134
rect 585342 471218 585578 471454
rect 585662 471218 585898 471454
rect 585342 470898 585578 471134
rect 585662 470898 585898 471134
rect 585342 435218 585578 435454
rect 585662 435218 585898 435454
rect 585342 434898 585578 435134
rect 585662 434898 585898 435134
rect 585342 399218 585578 399454
rect 585662 399218 585898 399454
rect 585342 398898 585578 399134
rect 585662 398898 585898 399134
rect 585342 363218 585578 363454
rect 585662 363218 585898 363454
rect 585342 362898 585578 363134
rect 585662 362898 585898 363134
rect 585342 327218 585578 327454
rect 585662 327218 585898 327454
rect 585342 326898 585578 327134
rect 585662 326898 585898 327134
rect 585342 291218 585578 291454
rect 585662 291218 585898 291454
rect 585342 290898 585578 291134
rect 585662 290898 585898 291134
rect 585342 255218 585578 255454
rect 585662 255218 585898 255454
rect 585342 254898 585578 255134
rect 585662 254898 585898 255134
rect 585342 219218 585578 219454
rect 585662 219218 585898 219454
rect 585342 218898 585578 219134
rect 585662 218898 585898 219134
rect 585342 183218 585578 183454
rect 585662 183218 585898 183454
rect 585342 182898 585578 183134
rect 585662 182898 585898 183134
rect 585342 147218 585578 147454
rect 585662 147218 585898 147454
rect 585342 146898 585578 147134
rect 585662 146898 585898 147134
rect 585342 111218 585578 111454
rect 585662 111218 585898 111454
rect 585342 110898 585578 111134
rect 585662 110898 585898 111134
rect 585342 75218 585578 75454
rect 585662 75218 585898 75454
rect 585342 74898 585578 75134
rect 585662 74898 585898 75134
rect 585342 39218 585578 39454
rect 585662 39218 585898 39454
rect 585342 38898 585578 39134
rect 585662 38898 585898 39134
rect 585342 3218 585578 3454
rect 585662 3218 585898 3454
rect 585342 2898 585578 3134
rect 585662 2898 585898 3134
rect 585342 -582 585578 -346
rect 585662 -582 585898 -346
rect 585342 -902 585578 -666
rect 585662 -902 585898 -666
rect 586302 691718 586538 691954
rect 586622 691718 586858 691954
rect 586302 691398 586538 691634
rect 586622 691398 586858 691634
rect 586302 655718 586538 655954
rect 586622 655718 586858 655954
rect 586302 655398 586538 655634
rect 586622 655398 586858 655634
rect 586302 619718 586538 619954
rect 586622 619718 586858 619954
rect 586302 619398 586538 619634
rect 586622 619398 586858 619634
rect 586302 583718 586538 583954
rect 586622 583718 586858 583954
rect 586302 583398 586538 583634
rect 586622 583398 586858 583634
rect 586302 547718 586538 547954
rect 586622 547718 586858 547954
rect 586302 547398 586538 547634
rect 586622 547398 586858 547634
rect 586302 511718 586538 511954
rect 586622 511718 586858 511954
rect 586302 511398 586538 511634
rect 586622 511398 586858 511634
rect 586302 475718 586538 475954
rect 586622 475718 586858 475954
rect 586302 475398 586538 475634
rect 586622 475398 586858 475634
rect 586302 439718 586538 439954
rect 586622 439718 586858 439954
rect 586302 439398 586538 439634
rect 586622 439398 586858 439634
rect 586302 403718 586538 403954
rect 586622 403718 586858 403954
rect 586302 403398 586538 403634
rect 586622 403398 586858 403634
rect 586302 367718 586538 367954
rect 586622 367718 586858 367954
rect 586302 367398 586538 367634
rect 586622 367398 586858 367634
rect 586302 331718 586538 331954
rect 586622 331718 586858 331954
rect 586302 331398 586538 331634
rect 586622 331398 586858 331634
rect 586302 295718 586538 295954
rect 586622 295718 586858 295954
rect 586302 295398 586538 295634
rect 586622 295398 586858 295634
rect 586302 259718 586538 259954
rect 586622 259718 586858 259954
rect 586302 259398 586538 259634
rect 586622 259398 586858 259634
rect 586302 223718 586538 223954
rect 586622 223718 586858 223954
rect 586302 223398 586538 223634
rect 586622 223398 586858 223634
rect 586302 187718 586538 187954
rect 586622 187718 586858 187954
rect 586302 187398 586538 187634
rect 586622 187398 586858 187634
rect 586302 151718 586538 151954
rect 586622 151718 586858 151954
rect 586302 151398 586538 151634
rect 586622 151398 586858 151634
rect 586302 115718 586538 115954
rect 586622 115718 586858 115954
rect 586302 115398 586538 115634
rect 586622 115398 586858 115634
rect 586302 79718 586538 79954
rect 586622 79718 586858 79954
rect 586302 79398 586538 79634
rect 586622 79398 586858 79634
rect 586302 43718 586538 43954
rect 586622 43718 586858 43954
rect 586302 43398 586538 43634
rect 586622 43398 586858 43634
rect 586302 7718 586538 7954
rect 586622 7718 586858 7954
rect 586302 7398 586538 7634
rect 586622 7398 586858 7634
rect 582326 -1542 582562 -1306
rect 582646 -1542 582882 -1306
rect 582326 -1862 582562 -1626
rect 582646 -1862 582882 -1626
rect 586302 -1542 586538 -1306
rect 586622 -1542 586858 -1306
rect 586302 -1862 586538 -1626
rect 586622 -1862 586858 -1626
rect 587262 696218 587498 696454
rect 587582 696218 587818 696454
rect 587262 695898 587498 696134
rect 587582 695898 587818 696134
rect 587262 660218 587498 660454
rect 587582 660218 587818 660454
rect 587262 659898 587498 660134
rect 587582 659898 587818 660134
rect 587262 624218 587498 624454
rect 587582 624218 587818 624454
rect 587262 623898 587498 624134
rect 587582 623898 587818 624134
rect 587262 588218 587498 588454
rect 587582 588218 587818 588454
rect 587262 587898 587498 588134
rect 587582 587898 587818 588134
rect 587262 552218 587498 552454
rect 587582 552218 587818 552454
rect 587262 551898 587498 552134
rect 587582 551898 587818 552134
rect 587262 516218 587498 516454
rect 587582 516218 587818 516454
rect 587262 515898 587498 516134
rect 587582 515898 587818 516134
rect 587262 480218 587498 480454
rect 587582 480218 587818 480454
rect 587262 479898 587498 480134
rect 587582 479898 587818 480134
rect 587262 444218 587498 444454
rect 587582 444218 587818 444454
rect 587262 443898 587498 444134
rect 587582 443898 587818 444134
rect 587262 408218 587498 408454
rect 587582 408218 587818 408454
rect 587262 407898 587498 408134
rect 587582 407898 587818 408134
rect 587262 372218 587498 372454
rect 587582 372218 587818 372454
rect 587262 371898 587498 372134
rect 587582 371898 587818 372134
rect 587262 336218 587498 336454
rect 587582 336218 587818 336454
rect 587262 335898 587498 336134
rect 587582 335898 587818 336134
rect 587262 300218 587498 300454
rect 587582 300218 587818 300454
rect 587262 299898 587498 300134
rect 587582 299898 587818 300134
rect 587262 264218 587498 264454
rect 587582 264218 587818 264454
rect 587262 263898 587498 264134
rect 587582 263898 587818 264134
rect 587262 228218 587498 228454
rect 587582 228218 587818 228454
rect 587262 227898 587498 228134
rect 587582 227898 587818 228134
rect 587262 192218 587498 192454
rect 587582 192218 587818 192454
rect 587262 191898 587498 192134
rect 587582 191898 587818 192134
rect 587262 156218 587498 156454
rect 587582 156218 587818 156454
rect 587262 155898 587498 156134
rect 587582 155898 587818 156134
rect 587262 120218 587498 120454
rect 587582 120218 587818 120454
rect 587262 119898 587498 120134
rect 587582 119898 587818 120134
rect 587262 84218 587498 84454
rect 587582 84218 587818 84454
rect 587262 83898 587498 84134
rect 587582 83898 587818 84134
rect 587262 48218 587498 48454
rect 587582 48218 587818 48454
rect 587262 47898 587498 48134
rect 587582 47898 587818 48134
rect 587262 12218 587498 12454
rect 587582 12218 587818 12454
rect 587262 11898 587498 12134
rect 587582 11898 587818 12134
rect 587262 -2502 587498 -2266
rect 587582 -2502 587818 -2266
rect 587262 -2822 587498 -2586
rect 587582 -2822 587818 -2586
rect 588222 700718 588458 700954
rect 588542 700718 588778 700954
rect 588222 700398 588458 700634
rect 588542 700398 588778 700634
rect 588222 664718 588458 664954
rect 588542 664718 588778 664954
rect 588222 664398 588458 664634
rect 588542 664398 588778 664634
rect 588222 628718 588458 628954
rect 588542 628718 588778 628954
rect 588222 628398 588458 628634
rect 588542 628398 588778 628634
rect 588222 592718 588458 592954
rect 588542 592718 588778 592954
rect 588222 592398 588458 592634
rect 588542 592398 588778 592634
rect 588222 556718 588458 556954
rect 588542 556718 588778 556954
rect 588222 556398 588458 556634
rect 588542 556398 588778 556634
rect 588222 520718 588458 520954
rect 588542 520718 588778 520954
rect 588222 520398 588458 520634
rect 588542 520398 588778 520634
rect 588222 484718 588458 484954
rect 588542 484718 588778 484954
rect 588222 484398 588458 484634
rect 588542 484398 588778 484634
rect 588222 448718 588458 448954
rect 588542 448718 588778 448954
rect 588222 448398 588458 448634
rect 588542 448398 588778 448634
rect 588222 412718 588458 412954
rect 588542 412718 588778 412954
rect 588222 412398 588458 412634
rect 588542 412398 588778 412634
rect 588222 376718 588458 376954
rect 588542 376718 588778 376954
rect 588222 376398 588458 376634
rect 588542 376398 588778 376634
rect 588222 340718 588458 340954
rect 588542 340718 588778 340954
rect 588222 340398 588458 340634
rect 588542 340398 588778 340634
rect 588222 304718 588458 304954
rect 588542 304718 588778 304954
rect 588222 304398 588458 304634
rect 588542 304398 588778 304634
rect 588222 268718 588458 268954
rect 588542 268718 588778 268954
rect 588222 268398 588458 268634
rect 588542 268398 588778 268634
rect 588222 232718 588458 232954
rect 588542 232718 588778 232954
rect 588222 232398 588458 232634
rect 588542 232398 588778 232634
rect 588222 196718 588458 196954
rect 588542 196718 588778 196954
rect 588222 196398 588458 196634
rect 588542 196398 588778 196634
rect 588222 160718 588458 160954
rect 588542 160718 588778 160954
rect 588222 160398 588458 160634
rect 588542 160398 588778 160634
rect 588222 124718 588458 124954
rect 588542 124718 588778 124954
rect 588222 124398 588458 124634
rect 588542 124398 588778 124634
rect 588222 88718 588458 88954
rect 588542 88718 588778 88954
rect 588222 88398 588458 88634
rect 588542 88398 588778 88634
rect 588222 52718 588458 52954
rect 588542 52718 588778 52954
rect 588222 52398 588458 52634
rect 588542 52398 588778 52634
rect 588222 16718 588458 16954
rect 588542 16718 588778 16954
rect 588222 16398 588458 16634
rect 588542 16398 588778 16634
rect 588222 -3462 588458 -3226
rect 588542 -3462 588778 -3226
rect 588222 -3782 588458 -3546
rect 588542 -3782 588778 -3546
rect 589182 669218 589418 669454
rect 589502 669218 589738 669454
rect 589182 668898 589418 669134
rect 589502 668898 589738 669134
rect 589182 633218 589418 633454
rect 589502 633218 589738 633454
rect 589182 632898 589418 633134
rect 589502 632898 589738 633134
rect 589182 597218 589418 597454
rect 589502 597218 589738 597454
rect 589182 596898 589418 597134
rect 589502 596898 589738 597134
rect 589182 561218 589418 561454
rect 589502 561218 589738 561454
rect 589182 560898 589418 561134
rect 589502 560898 589738 561134
rect 589182 525218 589418 525454
rect 589502 525218 589738 525454
rect 589182 524898 589418 525134
rect 589502 524898 589738 525134
rect 589182 489218 589418 489454
rect 589502 489218 589738 489454
rect 589182 488898 589418 489134
rect 589502 488898 589738 489134
rect 589182 453218 589418 453454
rect 589502 453218 589738 453454
rect 589182 452898 589418 453134
rect 589502 452898 589738 453134
rect 589182 417218 589418 417454
rect 589502 417218 589738 417454
rect 589182 416898 589418 417134
rect 589502 416898 589738 417134
rect 589182 381218 589418 381454
rect 589502 381218 589738 381454
rect 589182 380898 589418 381134
rect 589502 380898 589738 381134
rect 589182 345218 589418 345454
rect 589502 345218 589738 345454
rect 589182 344898 589418 345134
rect 589502 344898 589738 345134
rect 589182 309218 589418 309454
rect 589502 309218 589738 309454
rect 589182 308898 589418 309134
rect 589502 308898 589738 309134
rect 589182 273218 589418 273454
rect 589502 273218 589738 273454
rect 589182 272898 589418 273134
rect 589502 272898 589738 273134
rect 589182 237218 589418 237454
rect 589502 237218 589738 237454
rect 589182 236898 589418 237134
rect 589502 236898 589738 237134
rect 589182 201218 589418 201454
rect 589502 201218 589738 201454
rect 589182 200898 589418 201134
rect 589502 200898 589738 201134
rect 589182 165218 589418 165454
rect 589502 165218 589738 165454
rect 589182 164898 589418 165134
rect 589502 164898 589738 165134
rect 589182 129218 589418 129454
rect 589502 129218 589738 129454
rect 589182 128898 589418 129134
rect 589502 128898 589738 129134
rect 589182 93218 589418 93454
rect 589502 93218 589738 93454
rect 589182 92898 589418 93134
rect 589502 92898 589738 93134
rect 589182 57218 589418 57454
rect 589502 57218 589738 57454
rect 589182 56898 589418 57134
rect 589502 56898 589738 57134
rect 589182 21218 589418 21454
rect 589502 21218 589738 21454
rect 589182 20898 589418 21134
rect 589502 20898 589738 21134
rect 589182 -4422 589418 -4186
rect 589502 -4422 589738 -4186
rect 589182 -4742 589418 -4506
rect 589502 -4742 589738 -4506
rect 590142 673718 590378 673954
rect 590462 673718 590698 673954
rect 590142 673398 590378 673634
rect 590462 673398 590698 673634
rect 590142 637718 590378 637954
rect 590462 637718 590698 637954
rect 590142 637398 590378 637634
rect 590462 637398 590698 637634
rect 590142 601718 590378 601954
rect 590462 601718 590698 601954
rect 590142 601398 590378 601634
rect 590462 601398 590698 601634
rect 590142 565718 590378 565954
rect 590462 565718 590698 565954
rect 590142 565398 590378 565634
rect 590462 565398 590698 565634
rect 590142 529718 590378 529954
rect 590462 529718 590698 529954
rect 590142 529398 590378 529634
rect 590462 529398 590698 529634
rect 590142 493718 590378 493954
rect 590462 493718 590698 493954
rect 590142 493398 590378 493634
rect 590462 493398 590698 493634
rect 590142 457718 590378 457954
rect 590462 457718 590698 457954
rect 590142 457398 590378 457634
rect 590462 457398 590698 457634
rect 590142 421718 590378 421954
rect 590462 421718 590698 421954
rect 590142 421398 590378 421634
rect 590462 421398 590698 421634
rect 590142 385718 590378 385954
rect 590462 385718 590698 385954
rect 590142 385398 590378 385634
rect 590462 385398 590698 385634
rect 590142 349718 590378 349954
rect 590462 349718 590698 349954
rect 590142 349398 590378 349634
rect 590462 349398 590698 349634
rect 590142 313718 590378 313954
rect 590462 313718 590698 313954
rect 590142 313398 590378 313634
rect 590462 313398 590698 313634
rect 590142 277718 590378 277954
rect 590462 277718 590698 277954
rect 590142 277398 590378 277634
rect 590462 277398 590698 277634
rect 590142 241718 590378 241954
rect 590462 241718 590698 241954
rect 590142 241398 590378 241634
rect 590462 241398 590698 241634
rect 590142 205718 590378 205954
rect 590462 205718 590698 205954
rect 590142 205398 590378 205634
rect 590462 205398 590698 205634
rect 590142 169718 590378 169954
rect 590462 169718 590698 169954
rect 590142 169398 590378 169634
rect 590462 169398 590698 169634
rect 590142 133718 590378 133954
rect 590462 133718 590698 133954
rect 590142 133398 590378 133634
rect 590462 133398 590698 133634
rect 590142 97718 590378 97954
rect 590462 97718 590698 97954
rect 590142 97398 590378 97634
rect 590462 97398 590698 97634
rect 590142 61718 590378 61954
rect 590462 61718 590698 61954
rect 590142 61398 590378 61634
rect 590462 61398 590698 61634
rect 590142 25718 590378 25954
rect 590462 25718 590698 25954
rect 590142 25398 590378 25634
rect 590462 25398 590698 25634
rect 590142 -5382 590378 -5146
rect 590462 -5382 590698 -5146
rect 590142 -5702 590378 -5466
rect 590462 -5702 590698 -5466
rect 591102 678218 591338 678454
rect 591422 678218 591658 678454
rect 591102 677898 591338 678134
rect 591422 677898 591658 678134
rect 591102 642218 591338 642454
rect 591422 642218 591658 642454
rect 591102 641898 591338 642134
rect 591422 641898 591658 642134
rect 591102 606218 591338 606454
rect 591422 606218 591658 606454
rect 591102 605898 591338 606134
rect 591422 605898 591658 606134
rect 591102 570218 591338 570454
rect 591422 570218 591658 570454
rect 591102 569898 591338 570134
rect 591422 569898 591658 570134
rect 591102 534218 591338 534454
rect 591422 534218 591658 534454
rect 591102 533898 591338 534134
rect 591422 533898 591658 534134
rect 591102 498218 591338 498454
rect 591422 498218 591658 498454
rect 591102 497898 591338 498134
rect 591422 497898 591658 498134
rect 591102 462218 591338 462454
rect 591422 462218 591658 462454
rect 591102 461898 591338 462134
rect 591422 461898 591658 462134
rect 591102 426218 591338 426454
rect 591422 426218 591658 426454
rect 591102 425898 591338 426134
rect 591422 425898 591658 426134
rect 591102 390218 591338 390454
rect 591422 390218 591658 390454
rect 591102 389898 591338 390134
rect 591422 389898 591658 390134
rect 591102 354218 591338 354454
rect 591422 354218 591658 354454
rect 591102 353898 591338 354134
rect 591422 353898 591658 354134
rect 591102 318218 591338 318454
rect 591422 318218 591658 318454
rect 591102 317898 591338 318134
rect 591422 317898 591658 318134
rect 591102 282218 591338 282454
rect 591422 282218 591658 282454
rect 591102 281898 591338 282134
rect 591422 281898 591658 282134
rect 591102 246218 591338 246454
rect 591422 246218 591658 246454
rect 591102 245898 591338 246134
rect 591422 245898 591658 246134
rect 591102 210218 591338 210454
rect 591422 210218 591658 210454
rect 591102 209898 591338 210134
rect 591422 209898 591658 210134
rect 591102 174218 591338 174454
rect 591422 174218 591658 174454
rect 591102 173898 591338 174134
rect 591422 173898 591658 174134
rect 591102 138218 591338 138454
rect 591422 138218 591658 138454
rect 591102 137898 591338 138134
rect 591422 137898 591658 138134
rect 591102 102218 591338 102454
rect 591422 102218 591658 102454
rect 591102 101898 591338 102134
rect 591422 101898 591658 102134
rect 591102 66218 591338 66454
rect 591422 66218 591658 66454
rect 591102 65898 591338 66134
rect 591422 65898 591658 66134
rect 591102 30218 591338 30454
rect 591422 30218 591658 30454
rect 591102 29898 591338 30134
rect 591422 29898 591658 30134
rect 591102 -6342 591338 -6106
rect 591422 -6342 591658 -6106
rect 591102 -6662 591338 -6426
rect 591422 -6662 591658 -6426
rect 592062 682718 592298 682954
rect 592382 682718 592618 682954
rect 592062 682398 592298 682634
rect 592382 682398 592618 682634
rect 592062 646718 592298 646954
rect 592382 646718 592618 646954
rect 592062 646398 592298 646634
rect 592382 646398 592618 646634
rect 592062 610718 592298 610954
rect 592382 610718 592618 610954
rect 592062 610398 592298 610634
rect 592382 610398 592618 610634
rect 592062 574718 592298 574954
rect 592382 574718 592618 574954
rect 592062 574398 592298 574634
rect 592382 574398 592618 574634
rect 592062 538718 592298 538954
rect 592382 538718 592618 538954
rect 592062 538398 592298 538634
rect 592382 538398 592618 538634
rect 592062 502718 592298 502954
rect 592382 502718 592618 502954
rect 592062 502398 592298 502634
rect 592382 502398 592618 502634
rect 592062 466718 592298 466954
rect 592382 466718 592618 466954
rect 592062 466398 592298 466634
rect 592382 466398 592618 466634
rect 592062 430718 592298 430954
rect 592382 430718 592618 430954
rect 592062 430398 592298 430634
rect 592382 430398 592618 430634
rect 592062 394718 592298 394954
rect 592382 394718 592618 394954
rect 592062 394398 592298 394634
rect 592382 394398 592618 394634
rect 592062 358718 592298 358954
rect 592382 358718 592618 358954
rect 592062 358398 592298 358634
rect 592382 358398 592618 358634
rect 592062 322718 592298 322954
rect 592382 322718 592618 322954
rect 592062 322398 592298 322634
rect 592382 322398 592618 322634
rect 592062 286718 592298 286954
rect 592382 286718 592618 286954
rect 592062 286398 592298 286634
rect 592382 286398 592618 286634
rect 592062 250718 592298 250954
rect 592382 250718 592618 250954
rect 592062 250398 592298 250634
rect 592382 250398 592618 250634
rect 592062 214718 592298 214954
rect 592382 214718 592618 214954
rect 592062 214398 592298 214634
rect 592382 214398 592618 214634
rect 592062 178718 592298 178954
rect 592382 178718 592618 178954
rect 592062 178398 592298 178634
rect 592382 178398 592618 178634
rect 592062 142718 592298 142954
rect 592382 142718 592618 142954
rect 592062 142398 592298 142634
rect 592382 142398 592618 142634
rect 592062 106718 592298 106954
rect 592382 106718 592618 106954
rect 592062 106398 592298 106634
rect 592382 106398 592618 106634
rect 592062 70718 592298 70954
rect 592382 70718 592618 70954
rect 592062 70398 592298 70634
rect 592382 70398 592618 70634
rect 592062 34718 592298 34954
rect 592382 34718 592618 34954
rect 592062 34398 592298 34634
rect 592382 34398 592618 34634
rect 592062 -7302 592298 -7066
rect 592382 -7302 592618 -7066
rect 592062 -7622 592298 -7386
rect 592382 -7622 592618 -7386
<< metal5 >>
rect -8726 711558 592650 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 33326 711558
rect 33562 711322 33646 711558
rect 33882 711322 69326 711558
rect 69562 711322 69646 711558
rect 69882 711322 105326 711558
rect 105562 711322 105646 711558
rect 105882 711322 141326 711558
rect 141562 711322 141646 711558
rect 141882 711322 177326 711558
rect 177562 711322 177646 711558
rect 177882 711322 213326 711558
rect 213562 711322 213646 711558
rect 213882 711322 249326 711558
rect 249562 711322 249646 711558
rect 249882 711322 285326 711558
rect 285562 711322 285646 711558
rect 285882 711322 321326 711558
rect 321562 711322 321646 711558
rect 321882 711322 357326 711558
rect 357562 711322 357646 711558
rect 357882 711322 393326 711558
rect 393562 711322 393646 711558
rect 393882 711322 429326 711558
rect 429562 711322 429646 711558
rect 429882 711322 465326 711558
rect 465562 711322 465646 711558
rect 465882 711322 501326 711558
rect 501562 711322 501646 711558
rect 501882 711322 537326 711558
rect 537562 711322 537646 711558
rect 537882 711322 573326 711558
rect 573562 711322 573646 711558
rect 573882 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect -8726 711238 592650 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 33326 711238
rect 33562 711002 33646 711238
rect 33882 711002 69326 711238
rect 69562 711002 69646 711238
rect 69882 711002 105326 711238
rect 105562 711002 105646 711238
rect 105882 711002 141326 711238
rect 141562 711002 141646 711238
rect 141882 711002 177326 711238
rect 177562 711002 177646 711238
rect 177882 711002 213326 711238
rect 213562 711002 213646 711238
rect 213882 711002 249326 711238
rect 249562 711002 249646 711238
rect 249882 711002 285326 711238
rect 285562 711002 285646 711238
rect 285882 711002 321326 711238
rect 321562 711002 321646 711238
rect 321882 711002 357326 711238
rect 357562 711002 357646 711238
rect 357882 711002 393326 711238
rect 393562 711002 393646 711238
rect 393882 711002 429326 711238
rect 429562 711002 429646 711238
rect 429882 711002 465326 711238
rect 465562 711002 465646 711238
rect 465882 711002 501326 711238
rect 501562 711002 501646 711238
rect 501882 711002 537326 711238
rect 537562 711002 537646 711238
rect 537882 711002 573326 711238
rect 573562 711002 573646 711238
rect 573882 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect -8726 710970 592650 711002
rect -7766 710598 591690 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 28826 710598
rect 29062 710362 29146 710598
rect 29382 710362 64826 710598
rect 65062 710362 65146 710598
rect 65382 710362 100826 710598
rect 101062 710362 101146 710598
rect 101382 710362 136826 710598
rect 137062 710362 137146 710598
rect 137382 710362 172826 710598
rect 173062 710362 173146 710598
rect 173382 710362 208826 710598
rect 209062 710362 209146 710598
rect 209382 710362 244826 710598
rect 245062 710362 245146 710598
rect 245382 710362 280826 710598
rect 281062 710362 281146 710598
rect 281382 710362 316826 710598
rect 317062 710362 317146 710598
rect 317382 710362 352826 710598
rect 353062 710362 353146 710598
rect 353382 710362 388826 710598
rect 389062 710362 389146 710598
rect 389382 710362 424826 710598
rect 425062 710362 425146 710598
rect 425382 710362 460826 710598
rect 461062 710362 461146 710598
rect 461382 710362 496826 710598
rect 497062 710362 497146 710598
rect 497382 710362 532826 710598
rect 533062 710362 533146 710598
rect 533382 710362 568826 710598
rect 569062 710362 569146 710598
rect 569382 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect -7766 710278 591690 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 28826 710278
rect 29062 710042 29146 710278
rect 29382 710042 64826 710278
rect 65062 710042 65146 710278
rect 65382 710042 100826 710278
rect 101062 710042 101146 710278
rect 101382 710042 136826 710278
rect 137062 710042 137146 710278
rect 137382 710042 172826 710278
rect 173062 710042 173146 710278
rect 173382 710042 208826 710278
rect 209062 710042 209146 710278
rect 209382 710042 244826 710278
rect 245062 710042 245146 710278
rect 245382 710042 280826 710278
rect 281062 710042 281146 710278
rect 281382 710042 316826 710278
rect 317062 710042 317146 710278
rect 317382 710042 352826 710278
rect 353062 710042 353146 710278
rect 353382 710042 388826 710278
rect 389062 710042 389146 710278
rect 389382 710042 424826 710278
rect 425062 710042 425146 710278
rect 425382 710042 460826 710278
rect 461062 710042 461146 710278
rect 461382 710042 496826 710278
rect 497062 710042 497146 710278
rect 497382 710042 532826 710278
rect 533062 710042 533146 710278
rect 533382 710042 568826 710278
rect 569062 710042 569146 710278
rect 569382 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect -7766 710010 591690 710042
rect -6806 709638 590730 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 24326 709638
rect 24562 709402 24646 709638
rect 24882 709402 60326 709638
rect 60562 709402 60646 709638
rect 60882 709402 96326 709638
rect 96562 709402 96646 709638
rect 96882 709402 132326 709638
rect 132562 709402 132646 709638
rect 132882 709402 168326 709638
rect 168562 709402 168646 709638
rect 168882 709402 204326 709638
rect 204562 709402 204646 709638
rect 204882 709402 240326 709638
rect 240562 709402 240646 709638
rect 240882 709402 276326 709638
rect 276562 709402 276646 709638
rect 276882 709402 312326 709638
rect 312562 709402 312646 709638
rect 312882 709402 348326 709638
rect 348562 709402 348646 709638
rect 348882 709402 384326 709638
rect 384562 709402 384646 709638
rect 384882 709402 420326 709638
rect 420562 709402 420646 709638
rect 420882 709402 456326 709638
rect 456562 709402 456646 709638
rect 456882 709402 492326 709638
rect 492562 709402 492646 709638
rect 492882 709402 528326 709638
rect 528562 709402 528646 709638
rect 528882 709402 564326 709638
rect 564562 709402 564646 709638
rect 564882 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect -6806 709318 590730 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 24326 709318
rect 24562 709082 24646 709318
rect 24882 709082 60326 709318
rect 60562 709082 60646 709318
rect 60882 709082 96326 709318
rect 96562 709082 96646 709318
rect 96882 709082 132326 709318
rect 132562 709082 132646 709318
rect 132882 709082 168326 709318
rect 168562 709082 168646 709318
rect 168882 709082 204326 709318
rect 204562 709082 204646 709318
rect 204882 709082 240326 709318
rect 240562 709082 240646 709318
rect 240882 709082 276326 709318
rect 276562 709082 276646 709318
rect 276882 709082 312326 709318
rect 312562 709082 312646 709318
rect 312882 709082 348326 709318
rect 348562 709082 348646 709318
rect 348882 709082 384326 709318
rect 384562 709082 384646 709318
rect 384882 709082 420326 709318
rect 420562 709082 420646 709318
rect 420882 709082 456326 709318
rect 456562 709082 456646 709318
rect 456882 709082 492326 709318
rect 492562 709082 492646 709318
rect 492882 709082 528326 709318
rect 528562 709082 528646 709318
rect 528882 709082 564326 709318
rect 564562 709082 564646 709318
rect 564882 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect -6806 709050 590730 709082
rect -5846 708678 589770 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 19826 708678
rect 20062 708442 20146 708678
rect 20382 708442 55826 708678
rect 56062 708442 56146 708678
rect 56382 708442 91826 708678
rect 92062 708442 92146 708678
rect 92382 708442 127826 708678
rect 128062 708442 128146 708678
rect 128382 708442 163826 708678
rect 164062 708442 164146 708678
rect 164382 708442 199826 708678
rect 200062 708442 200146 708678
rect 200382 708442 235826 708678
rect 236062 708442 236146 708678
rect 236382 708442 271826 708678
rect 272062 708442 272146 708678
rect 272382 708442 307826 708678
rect 308062 708442 308146 708678
rect 308382 708442 343826 708678
rect 344062 708442 344146 708678
rect 344382 708442 379826 708678
rect 380062 708442 380146 708678
rect 380382 708442 415826 708678
rect 416062 708442 416146 708678
rect 416382 708442 451826 708678
rect 452062 708442 452146 708678
rect 452382 708442 487826 708678
rect 488062 708442 488146 708678
rect 488382 708442 523826 708678
rect 524062 708442 524146 708678
rect 524382 708442 559826 708678
rect 560062 708442 560146 708678
rect 560382 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect -5846 708358 589770 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 19826 708358
rect 20062 708122 20146 708358
rect 20382 708122 55826 708358
rect 56062 708122 56146 708358
rect 56382 708122 91826 708358
rect 92062 708122 92146 708358
rect 92382 708122 127826 708358
rect 128062 708122 128146 708358
rect 128382 708122 163826 708358
rect 164062 708122 164146 708358
rect 164382 708122 199826 708358
rect 200062 708122 200146 708358
rect 200382 708122 235826 708358
rect 236062 708122 236146 708358
rect 236382 708122 271826 708358
rect 272062 708122 272146 708358
rect 272382 708122 307826 708358
rect 308062 708122 308146 708358
rect 308382 708122 343826 708358
rect 344062 708122 344146 708358
rect 344382 708122 379826 708358
rect 380062 708122 380146 708358
rect 380382 708122 415826 708358
rect 416062 708122 416146 708358
rect 416382 708122 451826 708358
rect 452062 708122 452146 708358
rect 452382 708122 487826 708358
rect 488062 708122 488146 708358
rect 488382 708122 523826 708358
rect 524062 708122 524146 708358
rect 524382 708122 559826 708358
rect 560062 708122 560146 708358
rect 560382 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect -5846 708090 589770 708122
rect -4886 707718 588810 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 15326 707718
rect 15562 707482 15646 707718
rect 15882 707482 51326 707718
rect 51562 707482 51646 707718
rect 51882 707482 87326 707718
rect 87562 707482 87646 707718
rect 87882 707482 123326 707718
rect 123562 707482 123646 707718
rect 123882 707482 159326 707718
rect 159562 707482 159646 707718
rect 159882 707482 195326 707718
rect 195562 707482 195646 707718
rect 195882 707482 231326 707718
rect 231562 707482 231646 707718
rect 231882 707482 267326 707718
rect 267562 707482 267646 707718
rect 267882 707482 303326 707718
rect 303562 707482 303646 707718
rect 303882 707482 339326 707718
rect 339562 707482 339646 707718
rect 339882 707482 375326 707718
rect 375562 707482 375646 707718
rect 375882 707482 411326 707718
rect 411562 707482 411646 707718
rect 411882 707482 447326 707718
rect 447562 707482 447646 707718
rect 447882 707482 483326 707718
rect 483562 707482 483646 707718
rect 483882 707482 519326 707718
rect 519562 707482 519646 707718
rect 519882 707482 555326 707718
rect 555562 707482 555646 707718
rect 555882 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect -4886 707398 588810 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 15326 707398
rect 15562 707162 15646 707398
rect 15882 707162 51326 707398
rect 51562 707162 51646 707398
rect 51882 707162 87326 707398
rect 87562 707162 87646 707398
rect 87882 707162 123326 707398
rect 123562 707162 123646 707398
rect 123882 707162 159326 707398
rect 159562 707162 159646 707398
rect 159882 707162 195326 707398
rect 195562 707162 195646 707398
rect 195882 707162 231326 707398
rect 231562 707162 231646 707398
rect 231882 707162 267326 707398
rect 267562 707162 267646 707398
rect 267882 707162 303326 707398
rect 303562 707162 303646 707398
rect 303882 707162 339326 707398
rect 339562 707162 339646 707398
rect 339882 707162 375326 707398
rect 375562 707162 375646 707398
rect 375882 707162 411326 707398
rect 411562 707162 411646 707398
rect 411882 707162 447326 707398
rect 447562 707162 447646 707398
rect 447882 707162 483326 707398
rect 483562 707162 483646 707398
rect 483882 707162 519326 707398
rect 519562 707162 519646 707398
rect 519882 707162 555326 707398
rect 555562 707162 555646 707398
rect 555882 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect -4886 707130 588810 707162
rect -3926 706758 587850 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 10826 706758
rect 11062 706522 11146 706758
rect 11382 706522 46826 706758
rect 47062 706522 47146 706758
rect 47382 706522 82826 706758
rect 83062 706522 83146 706758
rect 83382 706522 118826 706758
rect 119062 706522 119146 706758
rect 119382 706522 154826 706758
rect 155062 706522 155146 706758
rect 155382 706522 190826 706758
rect 191062 706522 191146 706758
rect 191382 706522 226826 706758
rect 227062 706522 227146 706758
rect 227382 706522 262826 706758
rect 263062 706522 263146 706758
rect 263382 706522 298826 706758
rect 299062 706522 299146 706758
rect 299382 706522 334826 706758
rect 335062 706522 335146 706758
rect 335382 706522 370826 706758
rect 371062 706522 371146 706758
rect 371382 706522 406826 706758
rect 407062 706522 407146 706758
rect 407382 706522 442826 706758
rect 443062 706522 443146 706758
rect 443382 706522 478826 706758
rect 479062 706522 479146 706758
rect 479382 706522 514826 706758
rect 515062 706522 515146 706758
rect 515382 706522 550826 706758
rect 551062 706522 551146 706758
rect 551382 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect -3926 706438 587850 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 10826 706438
rect 11062 706202 11146 706438
rect 11382 706202 46826 706438
rect 47062 706202 47146 706438
rect 47382 706202 82826 706438
rect 83062 706202 83146 706438
rect 83382 706202 118826 706438
rect 119062 706202 119146 706438
rect 119382 706202 154826 706438
rect 155062 706202 155146 706438
rect 155382 706202 190826 706438
rect 191062 706202 191146 706438
rect 191382 706202 226826 706438
rect 227062 706202 227146 706438
rect 227382 706202 262826 706438
rect 263062 706202 263146 706438
rect 263382 706202 298826 706438
rect 299062 706202 299146 706438
rect 299382 706202 334826 706438
rect 335062 706202 335146 706438
rect 335382 706202 370826 706438
rect 371062 706202 371146 706438
rect 371382 706202 406826 706438
rect 407062 706202 407146 706438
rect 407382 706202 442826 706438
rect 443062 706202 443146 706438
rect 443382 706202 478826 706438
rect 479062 706202 479146 706438
rect 479382 706202 514826 706438
rect 515062 706202 515146 706438
rect 515382 706202 550826 706438
rect 551062 706202 551146 706438
rect 551382 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect -3926 706170 587850 706202
rect -2966 705798 586890 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 6326 705798
rect 6562 705562 6646 705798
rect 6882 705562 42326 705798
rect 42562 705562 42646 705798
rect 42882 705562 78326 705798
rect 78562 705562 78646 705798
rect 78882 705562 114326 705798
rect 114562 705562 114646 705798
rect 114882 705562 150326 705798
rect 150562 705562 150646 705798
rect 150882 705562 186326 705798
rect 186562 705562 186646 705798
rect 186882 705562 222326 705798
rect 222562 705562 222646 705798
rect 222882 705562 258326 705798
rect 258562 705562 258646 705798
rect 258882 705562 294326 705798
rect 294562 705562 294646 705798
rect 294882 705562 330326 705798
rect 330562 705562 330646 705798
rect 330882 705562 366326 705798
rect 366562 705562 366646 705798
rect 366882 705562 402326 705798
rect 402562 705562 402646 705798
rect 402882 705562 438326 705798
rect 438562 705562 438646 705798
rect 438882 705562 474326 705798
rect 474562 705562 474646 705798
rect 474882 705562 510326 705798
rect 510562 705562 510646 705798
rect 510882 705562 546326 705798
rect 546562 705562 546646 705798
rect 546882 705562 582326 705798
rect 582562 705562 582646 705798
rect 582882 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect -2966 705478 586890 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 6326 705478
rect 6562 705242 6646 705478
rect 6882 705242 42326 705478
rect 42562 705242 42646 705478
rect 42882 705242 78326 705478
rect 78562 705242 78646 705478
rect 78882 705242 114326 705478
rect 114562 705242 114646 705478
rect 114882 705242 150326 705478
rect 150562 705242 150646 705478
rect 150882 705242 186326 705478
rect 186562 705242 186646 705478
rect 186882 705242 222326 705478
rect 222562 705242 222646 705478
rect 222882 705242 258326 705478
rect 258562 705242 258646 705478
rect 258882 705242 294326 705478
rect 294562 705242 294646 705478
rect 294882 705242 330326 705478
rect 330562 705242 330646 705478
rect 330882 705242 366326 705478
rect 366562 705242 366646 705478
rect 366882 705242 402326 705478
rect 402562 705242 402646 705478
rect 402882 705242 438326 705478
rect 438562 705242 438646 705478
rect 438882 705242 474326 705478
rect 474562 705242 474646 705478
rect 474882 705242 510326 705478
rect 510562 705242 510646 705478
rect 510882 705242 546326 705478
rect 546562 705242 546646 705478
rect 546882 705242 582326 705478
rect 582562 705242 582646 705478
rect 582882 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect -2966 705210 586890 705242
rect -2006 704838 585930 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect -2006 704518 585930 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect -2006 704250 585930 704282
rect -8726 700954 592650 700986
rect -8726 700718 -4854 700954
rect -4618 700718 -4534 700954
rect -4298 700718 15326 700954
rect 15562 700718 15646 700954
rect 15882 700718 51326 700954
rect 51562 700718 51646 700954
rect 51882 700718 87326 700954
rect 87562 700718 87646 700954
rect 87882 700718 123326 700954
rect 123562 700718 123646 700954
rect 123882 700718 159326 700954
rect 159562 700718 159646 700954
rect 159882 700718 195326 700954
rect 195562 700718 195646 700954
rect 195882 700718 231326 700954
rect 231562 700718 231646 700954
rect 231882 700718 267326 700954
rect 267562 700718 267646 700954
rect 267882 700718 303326 700954
rect 303562 700718 303646 700954
rect 303882 700718 339326 700954
rect 339562 700718 339646 700954
rect 339882 700718 375326 700954
rect 375562 700718 375646 700954
rect 375882 700718 411326 700954
rect 411562 700718 411646 700954
rect 411882 700718 447326 700954
rect 447562 700718 447646 700954
rect 447882 700718 483326 700954
rect 483562 700718 483646 700954
rect 483882 700718 519326 700954
rect 519562 700718 519646 700954
rect 519882 700718 555326 700954
rect 555562 700718 555646 700954
rect 555882 700718 588222 700954
rect 588458 700718 588542 700954
rect 588778 700718 592650 700954
rect -8726 700634 592650 700718
rect -8726 700398 -4854 700634
rect -4618 700398 -4534 700634
rect -4298 700398 15326 700634
rect 15562 700398 15646 700634
rect 15882 700398 51326 700634
rect 51562 700398 51646 700634
rect 51882 700398 87326 700634
rect 87562 700398 87646 700634
rect 87882 700398 123326 700634
rect 123562 700398 123646 700634
rect 123882 700398 159326 700634
rect 159562 700398 159646 700634
rect 159882 700398 195326 700634
rect 195562 700398 195646 700634
rect 195882 700398 231326 700634
rect 231562 700398 231646 700634
rect 231882 700398 267326 700634
rect 267562 700398 267646 700634
rect 267882 700398 303326 700634
rect 303562 700398 303646 700634
rect 303882 700398 339326 700634
rect 339562 700398 339646 700634
rect 339882 700398 375326 700634
rect 375562 700398 375646 700634
rect 375882 700398 411326 700634
rect 411562 700398 411646 700634
rect 411882 700398 447326 700634
rect 447562 700398 447646 700634
rect 447882 700398 483326 700634
rect 483562 700398 483646 700634
rect 483882 700398 519326 700634
rect 519562 700398 519646 700634
rect 519882 700398 555326 700634
rect 555562 700398 555646 700634
rect 555882 700398 588222 700634
rect 588458 700398 588542 700634
rect 588778 700398 592650 700634
rect -8726 700366 592650 700398
rect -8726 696454 592650 696486
rect -8726 696218 -3894 696454
rect -3658 696218 -3574 696454
rect -3338 696218 10826 696454
rect 11062 696218 11146 696454
rect 11382 696218 46826 696454
rect 47062 696218 47146 696454
rect 47382 696218 82826 696454
rect 83062 696218 83146 696454
rect 83382 696218 118826 696454
rect 119062 696218 119146 696454
rect 119382 696218 154826 696454
rect 155062 696218 155146 696454
rect 155382 696218 190826 696454
rect 191062 696218 191146 696454
rect 191382 696218 226826 696454
rect 227062 696218 227146 696454
rect 227382 696218 262826 696454
rect 263062 696218 263146 696454
rect 263382 696218 298826 696454
rect 299062 696218 299146 696454
rect 299382 696218 334826 696454
rect 335062 696218 335146 696454
rect 335382 696218 370826 696454
rect 371062 696218 371146 696454
rect 371382 696218 406826 696454
rect 407062 696218 407146 696454
rect 407382 696218 442826 696454
rect 443062 696218 443146 696454
rect 443382 696218 478826 696454
rect 479062 696218 479146 696454
rect 479382 696218 514826 696454
rect 515062 696218 515146 696454
rect 515382 696218 550826 696454
rect 551062 696218 551146 696454
rect 551382 696218 587262 696454
rect 587498 696218 587582 696454
rect 587818 696218 592650 696454
rect -8726 696134 592650 696218
rect -8726 695898 -3894 696134
rect -3658 695898 -3574 696134
rect -3338 695898 10826 696134
rect 11062 695898 11146 696134
rect 11382 695898 46826 696134
rect 47062 695898 47146 696134
rect 47382 695898 82826 696134
rect 83062 695898 83146 696134
rect 83382 695898 118826 696134
rect 119062 695898 119146 696134
rect 119382 695898 154826 696134
rect 155062 695898 155146 696134
rect 155382 695898 190826 696134
rect 191062 695898 191146 696134
rect 191382 695898 226826 696134
rect 227062 695898 227146 696134
rect 227382 695898 262826 696134
rect 263062 695898 263146 696134
rect 263382 695898 298826 696134
rect 299062 695898 299146 696134
rect 299382 695898 334826 696134
rect 335062 695898 335146 696134
rect 335382 695898 370826 696134
rect 371062 695898 371146 696134
rect 371382 695898 406826 696134
rect 407062 695898 407146 696134
rect 407382 695898 442826 696134
rect 443062 695898 443146 696134
rect 443382 695898 478826 696134
rect 479062 695898 479146 696134
rect 479382 695898 514826 696134
rect 515062 695898 515146 696134
rect 515382 695898 550826 696134
rect 551062 695898 551146 696134
rect 551382 695898 587262 696134
rect 587498 695898 587582 696134
rect 587818 695898 592650 696134
rect -8726 695866 592650 695898
rect -8726 691954 592650 691986
rect -8726 691718 -2934 691954
rect -2698 691718 -2614 691954
rect -2378 691718 6326 691954
rect 6562 691718 6646 691954
rect 6882 691718 42326 691954
rect 42562 691718 42646 691954
rect 42882 691718 78326 691954
rect 78562 691718 78646 691954
rect 78882 691718 114326 691954
rect 114562 691718 114646 691954
rect 114882 691718 150326 691954
rect 150562 691718 150646 691954
rect 150882 691718 186326 691954
rect 186562 691718 186646 691954
rect 186882 691718 222326 691954
rect 222562 691718 222646 691954
rect 222882 691718 258326 691954
rect 258562 691718 258646 691954
rect 258882 691718 294326 691954
rect 294562 691718 294646 691954
rect 294882 691718 330326 691954
rect 330562 691718 330646 691954
rect 330882 691718 366326 691954
rect 366562 691718 366646 691954
rect 366882 691718 402326 691954
rect 402562 691718 402646 691954
rect 402882 691718 438326 691954
rect 438562 691718 438646 691954
rect 438882 691718 474326 691954
rect 474562 691718 474646 691954
rect 474882 691718 510326 691954
rect 510562 691718 510646 691954
rect 510882 691718 546326 691954
rect 546562 691718 546646 691954
rect 546882 691718 582326 691954
rect 582562 691718 582646 691954
rect 582882 691718 586302 691954
rect 586538 691718 586622 691954
rect 586858 691718 592650 691954
rect -8726 691634 592650 691718
rect -8726 691398 -2934 691634
rect -2698 691398 -2614 691634
rect -2378 691398 6326 691634
rect 6562 691398 6646 691634
rect 6882 691398 42326 691634
rect 42562 691398 42646 691634
rect 42882 691398 78326 691634
rect 78562 691398 78646 691634
rect 78882 691398 114326 691634
rect 114562 691398 114646 691634
rect 114882 691398 150326 691634
rect 150562 691398 150646 691634
rect 150882 691398 186326 691634
rect 186562 691398 186646 691634
rect 186882 691398 222326 691634
rect 222562 691398 222646 691634
rect 222882 691398 258326 691634
rect 258562 691398 258646 691634
rect 258882 691398 294326 691634
rect 294562 691398 294646 691634
rect 294882 691398 330326 691634
rect 330562 691398 330646 691634
rect 330882 691398 366326 691634
rect 366562 691398 366646 691634
rect 366882 691398 402326 691634
rect 402562 691398 402646 691634
rect 402882 691398 438326 691634
rect 438562 691398 438646 691634
rect 438882 691398 474326 691634
rect 474562 691398 474646 691634
rect 474882 691398 510326 691634
rect 510562 691398 510646 691634
rect 510882 691398 546326 691634
rect 546562 691398 546646 691634
rect 546882 691398 582326 691634
rect 582562 691398 582646 691634
rect 582882 691398 586302 691634
rect 586538 691398 586622 691634
rect 586858 691398 592650 691634
rect -8726 691366 592650 691398
rect -8726 687454 592650 687486
rect -8726 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 592650 687454
rect -8726 687134 592650 687218
rect -8726 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 592650 687134
rect -8726 686866 592650 686898
rect -8726 682954 592650 682986
rect -8726 682718 -8694 682954
rect -8458 682718 -8374 682954
rect -8138 682718 33326 682954
rect 33562 682718 33646 682954
rect 33882 682718 69326 682954
rect 69562 682718 69646 682954
rect 69882 682718 105326 682954
rect 105562 682718 105646 682954
rect 105882 682718 141326 682954
rect 141562 682718 141646 682954
rect 141882 682718 177326 682954
rect 177562 682718 177646 682954
rect 177882 682718 213326 682954
rect 213562 682718 213646 682954
rect 213882 682718 249326 682954
rect 249562 682718 249646 682954
rect 249882 682718 285326 682954
rect 285562 682718 285646 682954
rect 285882 682718 321326 682954
rect 321562 682718 321646 682954
rect 321882 682718 357326 682954
rect 357562 682718 357646 682954
rect 357882 682718 393326 682954
rect 393562 682718 393646 682954
rect 393882 682718 429326 682954
rect 429562 682718 429646 682954
rect 429882 682718 465326 682954
rect 465562 682718 465646 682954
rect 465882 682718 501326 682954
rect 501562 682718 501646 682954
rect 501882 682718 537326 682954
rect 537562 682718 537646 682954
rect 537882 682718 573326 682954
rect 573562 682718 573646 682954
rect 573882 682718 592062 682954
rect 592298 682718 592382 682954
rect 592618 682718 592650 682954
rect -8726 682634 592650 682718
rect -8726 682398 -8694 682634
rect -8458 682398 -8374 682634
rect -8138 682398 33326 682634
rect 33562 682398 33646 682634
rect 33882 682398 69326 682634
rect 69562 682398 69646 682634
rect 69882 682398 105326 682634
rect 105562 682398 105646 682634
rect 105882 682398 141326 682634
rect 141562 682398 141646 682634
rect 141882 682398 177326 682634
rect 177562 682398 177646 682634
rect 177882 682398 213326 682634
rect 213562 682398 213646 682634
rect 213882 682398 249326 682634
rect 249562 682398 249646 682634
rect 249882 682398 285326 682634
rect 285562 682398 285646 682634
rect 285882 682398 321326 682634
rect 321562 682398 321646 682634
rect 321882 682398 357326 682634
rect 357562 682398 357646 682634
rect 357882 682398 393326 682634
rect 393562 682398 393646 682634
rect 393882 682398 429326 682634
rect 429562 682398 429646 682634
rect 429882 682398 465326 682634
rect 465562 682398 465646 682634
rect 465882 682398 501326 682634
rect 501562 682398 501646 682634
rect 501882 682398 537326 682634
rect 537562 682398 537646 682634
rect 537882 682398 573326 682634
rect 573562 682398 573646 682634
rect 573882 682398 592062 682634
rect 592298 682398 592382 682634
rect 592618 682398 592650 682634
rect -8726 682366 592650 682398
rect -8726 678454 592650 678486
rect -8726 678218 -7734 678454
rect -7498 678218 -7414 678454
rect -7178 678218 28826 678454
rect 29062 678218 29146 678454
rect 29382 678218 64826 678454
rect 65062 678218 65146 678454
rect 65382 678218 100826 678454
rect 101062 678218 101146 678454
rect 101382 678218 136826 678454
rect 137062 678218 137146 678454
rect 137382 678218 172826 678454
rect 173062 678218 173146 678454
rect 173382 678218 208826 678454
rect 209062 678218 209146 678454
rect 209382 678218 244826 678454
rect 245062 678218 245146 678454
rect 245382 678218 280826 678454
rect 281062 678218 281146 678454
rect 281382 678218 316826 678454
rect 317062 678218 317146 678454
rect 317382 678218 352826 678454
rect 353062 678218 353146 678454
rect 353382 678218 388826 678454
rect 389062 678218 389146 678454
rect 389382 678218 424826 678454
rect 425062 678218 425146 678454
rect 425382 678218 460826 678454
rect 461062 678218 461146 678454
rect 461382 678218 496826 678454
rect 497062 678218 497146 678454
rect 497382 678218 532826 678454
rect 533062 678218 533146 678454
rect 533382 678218 568826 678454
rect 569062 678218 569146 678454
rect 569382 678218 591102 678454
rect 591338 678218 591422 678454
rect 591658 678218 592650 678454
rect -8726 678134 592650 678218
rect -8726 677898 -7734 678134
rect -7498 677898 -7414 678134
rect -7178 677898 28826 678134
rect 29062 677898 29146 678134
rect 29382 677898 64826 678134
rect 65062 677898 65146 678134
rect 65382 677898 100826 678134
rect 101062 677898 101146 678134
rect 101382 677898 136826 678134
rect 137062 677898 137146 678134
rect 137382 677898 172826 678134
rect 173062 677898 173146 678134
rect 173382 677898 208826 678134
rect 209062 677898 209146 678134
rect 209382 677898 244826 678134
rect 245062 677898 245146 678134
rect 245382 677898 280826 678134
rect 281062 677898 281146 678134
rect 281382 677898 316826 678134
rect 317062 677898 317146 678134
rect 317382 677898 352826 678134
rect 353062 677898 353146 678134
rect 353382 677898 388826 678134
rect 389062 677898 389146 678134
rect 389382 677898 424826 678134
rect 425062 677898 425146 678134
rect 425382 677898 460826 678134
rect 461062 677898 461146 678134
rect 461382 677898 496826 678134
rect 497062 677898 497146 678134
rect 497382 677898 532826 678134
rect 533062 677898 533146 678134
rect 533382 677898 568826 678134
rect 569062 677898 569146 678134
rect 569382 677898 591102 678134
rect 591338 677898 591422 678134
rect 591658 677898 592650 678134
rect -8726 677866 592650 677898
rect -8726 673954 592650 673986
rect -8726 673718 -6774 673954
rect -6538 673718 -6454 673954
rect -6218 673718 24326 673954
rect 24562 673718 24646 673954
rect 24882 673718 60326 673954
rect 60562 673718 60646 673954
rect 60882 673718 96326 673954
rect 96562 673718 96646 673954
rect 96882 673718 132326 673954
rect 132562 673718 132646 673954
rect 132882 673718 168326 673954
rect 168562 673718 168646 673954
rect 168882 673718 204326 673954
rect 204562 673718 204646 673954
rect 204882 673718 240326 673954
rect 240562 673718 240646 673954
rect 240882 673718 276326 673954
rect 276562 673718 276646 673954
rect 276882 673718 312326 673954
rect 312562 673718 312646 673954
rect 312882 673718 348326 673954
rect 348562 673718 348646 673954
rect 348882 673718 384326 673954
rect 384562 673718 384646 673954
rect 384882 673718 420326 673954
rect 420562 673718 420646 673954
rect 420882 673718 456326 673954
rect 456562 673718 456646 673954
rect 456882 673718 492326 673954
rect 492562 673718 492646 673954
rect 492882 673718 528326 673954
rect 528562 673718 528646 673954
rect 528882 673718 564326 673954
rect 564562 673718 564646 673954
rect 564882 673718 590142 673954
rect 590378 673718 590462 673954
rect 590698 673718 592650 673954
rect -8726 673634 592650 673718
rect -8726 673398 -6774 673634
rect -6538 673398 -6454 673634
rect -6218 673398 24326 673634
rect 24562 673398 24646 673634
rect 24882 673398 60326 673634
rect 60562 673398 60646 673634
rect 60882 673398 96326 673634
rect 96562 673398 96646 673634
rect 96882 673398 132326 673634
rect 132562 673398 132646 673634
rect 132882 673398 168326 673634
rect 168562 673398 168646 673634
rect 168882 673398 204326 673634
rect 204562 673398 204646 673634
rect 204882 673398 240326 673634
rect 240562 673398 240646 673634
rect 240882 673398 276326 673634
rect 276562 673398 276646 673634
rect 276882 673398 312326 673634
rect 312562 673398 312646 673634
rect 312882 673398 348326 673634
rect 348562 673398 348646 673634
rect 348882 673398 384326 673634
rect 384562 673398 384646 673634
rect 384882 673398 420326 673634
rect 420562 673398 420646 673634
rect 420882 673398 456326 673634
rect 456562 673398 456646 673634
rect 456882 673398 492326 673634
rect 492562 673398 492646 673634
rect 492882 673398 528326 673634
rect 528562 673398 528646 673634
rect 528882 673398 564326 673634
rect 564562 673398 564646 673634
rect 564882 673398 590142 673634
rect 590378 673398 590462 673634
rect 590698 673398 592650 673634
rect -8726 673366 592650 673398
rect -8726 669454 592650 669486
rect -8726 669218 -5814 669454
rect -5578 669218 -5494 669454
rect -5258 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 55826 669454
rect 56062 669218 56146 669454
rect 56382 669218 91826 669454
rect 92062 669218 92146 669454
rect 92382 669218 127826 669454
rect 128062 669218 128146 669454
rect 128382 669218 163826 669454
rect 164062 669218 164146 669454
rect 164382 669218 199826 669454
rect 200062 669218 200146 669454
rect 200382 669218 235826 669454
rect 236062 669218 236146 669454
rect 236382 669218 271826 669454
rect 272062 669218 272146 669454
rect 272382 669218 307826 669454
rect 308062 669218 308146 669454
rect 308382 669218 343826 669454
rect 344062 669218 344146 669454
rect 344382 669218 379826 669454
rect 380062 669218 380146 669454
rect 380382 669218 415826 669454
rect 416062 669218 416146 669454
rect 416382 669218 451826 669454
rect 452062 669218 452146 669454
rect 452382 669218 487826 669454
rect 488062 669218 488146 669454
rect 488382 669218 523826 669454
rect 524062 669218 524146 669454
rect 524382 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 589182 669454
rect 589418 669218 589502 669454
rect 589738 669218 592650 669454
rect -8726 669134 592650 669218
rect -8726 668898 -5814 669134
rect -5578 668898 -5494 669134
rect -5258 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 55826 669134
rect 56062 668898 56146 669134
rect 56382 668898 91826 669134
rect 92062 668898 92146 669134
rect 92382 668898 127826 669134
rect 128062 668898 128146 669134
rect 128382 668898 163826 669134
rect 164062 668898 164146 669134
rect 164382 668898 199826 669134
rect 200062 668898 200146 669134
rect 200382 668898 235826 669134
rect 236062 668898 236146 669134
rect 236382 668898 271826 669134
rect 272062 668898 272146 669134
rect 272382 668898 307826 669134
rect 308062 668898 308146 669134
rect 308382 668898 343826 669134
rect 344062 668898 344146 669134
rect 344382 668898 379826 669134
rect 380062 668898 380146 669134
rect 380382 668898 415826 669134
rect 416062 668898 416146 669134
rect 416382 668898 451826 669134
rect 452062 668898 452146 669134
rect 452382 668898 487826 669134
rect 488062 668898 488146 669134
rect 488382 668898 523826 669134
rect 524062 668898 524146 669134
rect 524382 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 589182 669134
rect 589418 668898 589502 669134
rect 589738 668898 592650 669134
rect -8726 668866 592650 668898
rect -8726 664954 592650 664986
rect -8726 664718 -4854 664954
rect -4618 664718 -4534 664954
rect -4298 664718 15326 664954
rect 15562 664718 15646 664954
rect 15882 664718 51326 664954
rect 51562 664718 51646 664954
rect 51882 664718 87326 664954
rect 87562 664718 87646 664954
rect 87882 664718 123326 664954
rect 123562 664718 123646 664954
rect 123882 664718 159326 664954
rect 159562 664718 159646 664954
rect 159882 664718 195326 664954
rect 195562 664718 195646 664954
rect 195882 664718 231326 664954
rect 231562 664718 231646 664954
rect 231882 664718 267326 664954
rect 267562 664718 267646 664954
rect 267882 664718 303326 664954
rect 303562 664718 303646 664954
rect 303882 664718 339326 664954
rect 339562 664718 339646 664954
rect 339882 664718 375326 664954
rect 375562 664718 375646 664954
rect 375882 664718 411326 664954
rect 411562 664718 411646 664954
rect 411882 664718 447326 664954
rect 447562 664718 447646 664954
rect 447882 664718 483326 664954
rect 483562 664718 483646 664954
rect 483882 664718 519326 664954
rect 519562 664718 519646 664954
rect 519882 664718 555326 664954
rect 555562 664718 555646 664954
rect 555882 664718 588222 664954
rect 588458 664718 588542 664954
rect 588778 664718 592650 664954
rect -8726 664634 592650 664718
rect -8726 664398 -4854 664634
rect -4618 664398 -4534 664634
rect -4298 664398 15326 664634
rect 15562 664398 15646 664634
rect 15882 664398 51326 664634
rect 51562 664398 51646 664634
rect 51882 664398 87326 664634
rect 87562 664398 87646 664634
rect 87882 664398 123326 664634
rect 123562 664398 123646 664634
rect 123882 664398 159326 664634
rect 159562 664398 159646 664634
rect 159882 664398 195326 664634
rect 195562 664398 195646 664634
rect 195882 664398 231326 664634
rect 231562 664398 231646 664634
rect 231882 664398 267326 664634
rect 267562 664398 267646 664634
rect 267882 664398 303326 664634
rect 303562 664398 303646 664634
rect 303882 664398 339326 664634
rect 339562 664398 339646 664634
rect 339882 664398 375326 664634
rect 375562 664398 375646 664634
rect 375882 664398 411326 664634
rect 411562 664398 411646 664634
rect 411882 664398 447326 664634
rect 447562 664398 447646 664634
rect 447882 664398 483326 664634
rect 483562 664398 483646 664634
rect 483882 664398 519326 664634
rect 519562 664398 519646 664634
rect 519882 664398 555326 664634
rect 555562 664398 555646 664634
rect 555882 664398 588222 664634
rect 588458 664398 588542 664634
rect 588778 664398 592650 664634
rect -8726 664366 592650 664398
rect -8726 660454 592650 660486
rect -8726 660218 -3894 660454
rect -3658 660218 -3574 660454
rect -3338 660218 10826 660454
rect 11062 660218 11146 660454
rect 11382 660218 46826 660454
rect 47062 660218 47146 660454
rect 47382 660218 82826 660454
rect 83062 660218 83146 660454
rect 83382 660218 118826 660454
rect 119062 660218 119146 660454
rect 119382 660218 154826 660454
rect 155062 660218 155146 660454
rect 155382 660218 190826 660454
rect 191062 660218 191146 660454
rect 191382 660218 226826 660454
rect 227062 660218 227146 660454
rect 227382 660218 262826 660454
rect 263062 660218 263146 660454
rect 263382 660218 298826 660454
rect 299062 660218 299146 660454
rect 299382 660218 334826 660454
rect 335062 660218 335146 660454
rect 335382 660218 370826 660454
rect 371062 660218 371146 660454
rect 371382 660218 406826 660454
rect 407062 660218 407146 660454
rect 407382 660218 442826 660454
rect 443062 660218 443146 660454
rect 443382 660218 478826 660454
rect 479062 660218 479146 660454
rect 479382 660218 514826 660454
rect 515062 660218 515146 660454
rect 515382 660218 550826 660454
rect 551062 660218 551146 660454
rect 551382 660218 587262 660454
rect 587498 660218 587582 660454
rect 587818 660218 592650 660454
rect -8726 660134 592650 660218
rect -8726 659898 -3894 660134
rect -3658 659898 -3574 660134
rect -3338 659898 10826 660134
rect 11062 659898 11146 660134
rect 11382 659898 46826 660134
rect 47062 659898 47146 660134
rect 47382 659898 82826 660134
rect 83062 659898 83146 660134
rect 83382 659898 118826 660134
rect 119062 659898 119146 660134
rect 119382 659898 154826 660134
rect 155062 659898 155146 660134
rect 155382 659898 190826 660134
rect 191062 659898 191146 660134
rect 191382 659898 226826 660134
rect 227062 659898 227146 660134
rect 227382 659898 262826 660134
rect 263062 659898 263146 660134
rect 263382 659898 298826 660134
rect 299062 659898 299146 660134
rect 299382 659898 334826 660134
rect 335062 659898 335146 660134
rect 335382 659898 370826 660134
rect 371062 659898 371146 660134
rect 371382 659898 406826 660134
rect 407062 659898 407146 660134
rect 407382 659898 442826 660134
rect 443062 659898 443146 660134
rect 443382 659898 478826 660134
rect 479062 659898 479146 660134
rect 479382 659898 514826 660134
rect 515062 659898 515146 660134
rect 515382 659898 550826 660134
rect 551062 659898 551146 660134
rect 551382 659898 587262 660134
rect 587498 659898 587582 660134
rect 587818 659898 592650 660134
rect -8726 659866 592650 659898
rect -8726 655954 592650 655986
rect -8726 655718 -2934 655954
rect -2698 655718 -2614 655954
rect -2378 655718 6326 655954
rect 6562 655718 6646 655954
rect 6882 655718 42326 655954
rect 42562 655718 42646 655954
rect 42882 655718 78326 655954
rect 78562 655718 78646 655954
rect 78882 655718 114326 655954
rect 114562 655718 114646 655954
rect 114882 655718 150326 655954
rect 150562 655718 150646 655954
rect 150882 655718 186326 655954
rect 186562 655718 186646 655954
rect 186882 655718 222326 655954
rect 222562 655718 222646 655954
rect 222882 655718 258326 655954
rect 258562 655718 258646 655954
rect 258882 655718 294326 655954
rect 294562 655718 294646 655954
rect 294882 655718 330326 655954
rect 330562 655718 330646 655954
rect 330882 655718 366326 655954
rect 366562 655718 366646 655954
rect 366882 655718 402326 655954
rect 402562 655718 402646 655954
rect 402882 655718 438326 655954
rect 438562 655718 438646 655954
rect 438882 655718 474326 655954
rect 474562 655718 474646 655954
rect 474882 655718 510326 655954
rect 510562 655718 510646 655954
rect 510882 655718 546326 655954
rect 546562 655718 546646 655954
rect 546882 655718 582326 655954
rect 582562 655718 582646 655954
rect 582882 655718 586302 655954
rect 586538 655718 586622 655954
rect 586858 655718 592650 655954
rect -8726 655634 592650 655718
rect -8726 655398 -2934 655634
rect -2698 655398 -2614 655634
rect -2378 655398 6326 655634
rect 6562 655398 6646 655634
rect 6882 655398 42326 655634
rect 42562 655398 42646 655634
rect 42882 655398 78326 655634
rect 78562 655398 78646 655634
rect 78882 655398 114326 655634
rect 114562 655398 114646 655634
rect 114882 655398 150326 655634
rect 150562 655398 150646 655634
rect 150882 655398 186326 655634
rect 186562 655398 186646 655634
rect 186882 655398 222326 655634
rect 222562 655398 222646 655634
rect 222882 655398 258326 655634
rect 258562 655398 258646 655634
rect 258882 655398 294326 655634
rect 294562 655398 294646 655634
rect 294882 655398 330326 655634
rect 330562 655398 330646 655634
rect 330882 655398 366326 655634
rect 366562 655398 366646 655634
rect 366882 655398 402326 655634
rect 402562 655398 402646 655634
rect 402882 655398 438326 655634
rect 438562 655398 438646 655634
rect 438882 655398 474326 655634
rect 474562 655398 474646 655634
rect 474882 655398 510326 655634
rect 510562 655398 510646 655634
rect 510882 655398 546326 655634
rect 546562 655398 546646 655634
rect 546882 655398 582326 655634
rect 582562 655398 582646 655634
rect 582882 655398 586302 655634
rect 586538 655398 586622 655634
rect 586858 655398 592650 655634
rect -8726 655366 592650 655398
rect -8726 651454 592650 651486
rect -8726 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 109826 651454
rect 110062 651218 110146 651454
rect 110382 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 592650 651454
rect -8726 651134 592650 651218
rect -8726 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 109826 651134
rect 110062 650898 110146 651134
rect 110382 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 592650 651134
rect -8726 650866 592650 650898
rect -8726 646954 592650 646986
rect -8726 646718 -8694 646954
rect -8458 646718 -8374 646954
rect -8138 646718 33326 646954
rect 33562 646718 33646 646954
rect 33882 646718 69326 646954
rect 69562 646718 69646 646954
rect 69882 646718 105326 646954
rect 105562 646718 105646 646954
rect 105882 646718 141326 646954
rect 141562 646718 141646 646954
rect 141882 646718 177326 646954
rect 177562 646718 177646 646954
rect 177882 646718 213326 646954
rect 213562 646718 213646 646954
rect 213882 646718 249326 646954
rect 249562 646718 249646 646954
rect 249882 646718 285326 646954
rect 285562 646718 285646 646954
rect 285882 646718 321326 646954
rect 321562 646718 321646 646954
rect 321882 646718 357326 646954
rect 357562 646718 357646 646954
rect 357882 646718 393326 646954
rect 393562 646718 393646 646954
rect 393882 646718 429326 646954
rect 429562 646718 429646 646954
rect 429882 646718 465326 646954
rect 465562 646718 465646 646954
rect 465882 646718 501326 646954
rect 501562 646718 501646 646954
rect 501882 646718 537326 646954
rect 537562 646718 537646 646954
rect 537882 646718 573326 646954
rect 573562 646718 573646 646954
rect 573882 646718 592062 646954
rect 592298 646718 592382 646954
rect 592618 646718 592650 646954
rect -8726 646634 592650 646718
rect -8726 646398 -8694 646634
rect -8458 646398 -8374 646634
rect -8138 646398 33326 646634
rect 33562 646398 33646 646634
rect 33882 646398 69326 646634
rect 69562 646398 69646 646634
rect 69882 646398 105326 646634
rect 105562 646398 105646 646634
rect 105882 646398 141326 646634
rect 141562 646398 141646 646634
rect 141882 646398 177326 646634
rect 177562 646398 177646 646634
rect 177882 646398 213326 646634
rect 213562 646398 213646 646634
rect 213882 646398 249326 646634
rect 249562 646398 249646 646634
rect 249882 646398 285326 646634
rect 285562 646398 285646 646634
rect 285882 646398 321326 646634
rect 321562 646398 321646 646634
rect 321882 646398 357326 646634
rect 357562 646398 357646 646634
rect 357882 646398 393326 646634
rect 393562 646398 393646 646634
rect 393882 646398 429326 646634
rect 429562 646398 429646 646634
rect 429882 646398 465326 646634
rect 465562 646398 465646 646634
rect 465882 646398 501326 646634
rect 501562 646398 501646 646634
rect 501882 646398 537326 646634
rect 537562 646398 537646 646634
rect 537882 646398 573326 646634
rect 573562 646398 573646 646634
rect 573882 646398 592062 646634
rect 592298 646398 592382 646634
rect 592618 646398 592650 646634
rect -8726 646366 592650 646398
rect -8726 642454 592650 642486
rect -8726 642218 -7734 642454
rect -7498 642218 -7414 642454
rect -7178 642218 28826 642454
rect 29062 642218 29146 642454
rect 29382 642218 64826 642454
rect 65062 642218 65146 642454
rect 65382 642218 100826 642454
rect 101062 642218 101146 642454
rect 101382 642218 136826 642454
rect 137062 642218 137146 642454
rect 137382 642218 172826 642454
rect 173062 642218 173146 642454
rect 173382 642218 208826 642454
rect 209062 642218 209146 642454
rect 209382 642218 244826 642454
rect 245062 642218 245146 642454
rect 245382 642218 280826 642454
rect 281062 642218 281146 642454
rect 281382 642218 316826 642454
rect 317062 642218 317146 642454
rect 317382 642218 352826 642454
rect 353062 642218 353146 642454
rect 353382 642218 388826 642454
rect 389062 642218 389146 642454
rect 389382 642218 424826 642454
rect 425062 642218 425146 642454
rect 425382 642218 460826 642454
rect 461062 642218 461146 642454
rect 461382 642218 496826 642454
rect 497062 642218 497146 642454
rect 497382 642218 532826 642454
rect 533062 642218 533146 642454
rect 533382 642218 568826 642454
rect 569062 642218 569146 642454
rect 569382 642218 591102 642454
rect 591338 642218 591422 642454
rect 591658 642218 592650 642454
rect -8726 642134 592650 642218
rect -8726 641898 -7734 642134
rect -7498 641898 -7414 642134
rect -7178 641898 28826 642134
rect 29062 641898 29146 642134
rect 29382 641898 64826 642134
rect 65062 641898 65146 642134
rect 65382 641898 100826 642134
rect 101062 641898 101146 642134
rect 101382 641898 136826 642134
rect 137062 641898 137146 642134
rect 137382 641898 172826 642134
rect 173062 641898 173146 642134
rect 173382 641898 208826 642134
rect 209062 641898 209146 642134
rect 209382 641898 244826 642134
rect 245062 641898 245146 642134
rect 245382 641898 280826 642134
rect 281062 641898 281146 642134
rect 281382 641898 316826 642134
rect 317062 641898 317146 642134
rect 317382 641898 352826 642134
rect 353062 641898 353146 642134
rect 353382 641898 388826 642134
rect 389062 641898 389146 642134
rect 389382 641898 424826 642134
rect 425062 641898 425146 642134
rect 425382 641898 460826 642134
rect 461062 641898 461146 642134
rect 461382 641898 496826 642134
rect 497062 641898 497146 642134
rect 497382 641898 532826 642134
rect 533062 641898 533146 642134
rect 533382 641898 568826 642134
rect 569062 641898 569146 642134
rect 569382 641898 591102 642134
rect 591338 641898 591422 642134
rect 591658 641898 592650 642134
rect -8726 641866 592650 641898
rect -8726 637954 592650 637986
rect -8726 637718 -6774 637954
rect -6538 637718 -6454 637954
rect -6218 637718 24326 637954
rect 24562 637718 24646 637954
rect 24882 637718 60326 637954
rect 60562 637718 60646 637954
rect 60882 637718 96326 637954
rect 96562 637718 96646 637954
rect 96882 637718 132326 637954
rect 132562 637718 132646 637954
rect 132882 637718 168326 637954
rect 168562 637718 168646 637954
rect 168882 637718 204326 637954
rect 204562 637718 204646 637954
rect 204882 637718 240326 637954
rect 240562 637718 240646 637954
rect 240882 637718 276326 637954
rect 276562 637718 276646 637954
rect 276882 637718 312326 637954
rect 312562 637718 312646 637954
rect 312882 637718 348326 637954
rect 348562 637718 348646 637954
rect 348882 637718 384326 637954
rect 384562 637718 384646 637954
rect 384882 637718 420326 637954
rect 420562 637718 420646 637954
rect 420882 637718 456326 637954
rect 456562 637718 456646 637954
rect 456882 637718 492326 637954
rect 492562 637718 492646 637954
rect 492882 637718 528326 637954
rect 528562 637718 528646 637954
rect 528882 637718 564326 637954
rect 564562 637718 564646 637954
rect 564882 637718 590142 637954
rect 590378 637718 590462 637954
rect 590698 637718 592650 637954
rect -8726 637634 592650 637718
rect -8726 637398 -6774 637634
rect -6538 637398 -6454 637634
rect -6218 637398 24326 637634
rect 24562 637398 24646 637634
rect 24882 637398 60326 637634
rect 60562 637398 60646 637634
rect 60882 637398 96326 637634
rect 96562 637398 96646 637634
rect 96882 637398 132326 637634
rect 132562 637398 132646 637634
rect 132882 637398 168326 637634
rect 168562 637398 168646 637634
rect 168882 637398 204326 637634
rect 204562 637398 204646 637634
rect 204882 637398 240326 637634
rect 240562 637398 240646 637634
rect 240882 637398 276326 637634
rect 276562 637398 276646 637634
rect 276882 637398 312326 637634
rect 312562 637398 312646 637634
rect 312882 637398 348326 637634
rect 348562 637398 348646 637634
rect 348882 637398 384326 637634
rect 384562 637398 384646 637634
rect 384882 637398 420326 637634
rect 420562 637398 420646 637634
rect 420882 637398 456326 637634
rect 456562 637398 456646 637634
rect 456882 637398 492326 637634
rect 492562 637398 492646 637634
rect 492882 637398 528326 637634
rect 528562 637398 528646 637634
rect 528882 637398 564326 637634
rect 564562 637398 564646 637634
rect 564882 637398 590142 637634
rect 590378 637398 590462 637634
rect 590698 637398 592650 637634
rect -8726 637366 592650 637398
rect -8726 633454 592650 633486
rect -8726 633218 -5814 633454
rect -5578 633218 -5494 633454
rect -5258 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 55826 633454
rect 56062 633218 56146 633454
rect 56382 633218 91826 633454
rect 92062 633218 92146 633454
rect 92382 633218 127826 633454
rect 128062 633218 128146 633454
rect 128382 633218 163826 633454
rect 164062 633218 164146 633454
rect 164382 633218 199826 633454
rect 200062 633218 200146 633454
rect 200382 633218 235826 633454
rect 236062 633218 236146 633454
rect 236382 633218 271826 633454
rect 272062 633218 272146 633454
rect 272382 633218 307826 633454
rect 308062 633218 308146 633454
rect 308382 633218 343826 633454
rect 344062 633218 344146 633454
rect 344382 633218 379826 633454
rect 380062 633218 380146 633454
rect 380382 633218 415826 633454
rect 416062 633218 416146 633454
rect 416382 633218 451826 633454
rect 452062 633218 452146 633454
rect 452382 633218 487826 633454
rect 488062 633218 488146 633454
rect 488382 633218 523826 633454
rect 524062 633218 524146 633454
rect 524382 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 589182 633454
rect 589418 633218 589502 633454
rect 589738 633218 592650 633454
rect -8726 633134 592650 633218
rect -8726 632898 -5814 633134
rect -5578 632898 -5494 633134
rect -5258 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 55826 633134
rect 56062 632898 56146 633134
rect 56382 632898 91826 633134
rect 92062 632898 92146 633134
rect 92382 632898 127826 633134
rect 128062 632898 128146 633134
rect 128382 632898 163826 633134
rect 164062 632898 164146 633134
rect 164382 632898 199826 633134
rect 200062 632898 200146 633134
rect 200382 632898 235826 633134
rect 236062 632898 236146 633134
rect 236382 632898 271826 633134
rect 272062 632898 272146 633134
rect 272382 632898 307826 633134
rect 308062 632898 308146 633134
rect 308382 632898 343826 633134
rect 344062 632898 344146 633134
rect 344382 632898 379826 633134
rect 380062 632898 380146 633134
rect 380382 632898 415826 633134
rect 416062 632898 416146 633134
rect 416382 632898 451826 633134
rect 452062 632898 452146 633134
rect 452382 632898 487826 633134
rect 488062 632898 488146 633134
rect 488382 632898 523826 633134
rect 524062 632898 524146 633134
rect 524382 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 589182 633134
rect 589418 632898 589502 633134
rect 589738 632898 592650 633134
rect -8726 632866 592650 632898
rect -8726 628954 592650 628986
rect -8726 628718 -4854 628954
rect -4618 628718 -4534 628954
rect -4298 628718 15326 628954
rect 15562 628718 15646 628954
rect 15882 628718 51326 628954
rect 51562 628718 51646 628954
rect 51882 628718 87326 628954
rect 87562 628718 87646 628954
rect 87882 628718 123326 628954
rect 123562 628718 123646 628954
rect 123882 628718 159326 628954
rect 159562 628718 159646 628954
rect 159882 628718 195326 628954
rect 195562 628718 195646 628954
rect 195882 628718 231326 628954
rect 231562 628718 231646 628954
rect 231882 628718 267326 628954
rect 267562 628718 267646 628954
rect 267882 628718 303326 628954
rect 303562 628718 303646 628954
rect 303882 628718 339326 628954
rect 339562 628718 339646 628954
rect 339882 628718 375326 628954
rect 375562 628718 375646 628954
rect 375882 628718 411326 628954
rect 411562 628718 411646 628954
rect 411882 628718 447326 628954
rect 447562 628718 447646 628954
rect 447882 628718 483326 628954
rect 483562 628718 483646 628954
rect 483882 628718 519326 628954
rect 519562 628718 519646 628954
rect 519882 628718 555326 628954
rect 555562 628718 555646 628954
rect 555882 628718 588222 628954
rect 588458 628718 588542 628954
rect 588778 628718 592650 628954
rect -8726 628634 592650 628718
rect -8726 628398 -4854 628634
rect -4618 628398 -4534 628634
rect -4298 628398 15326 628634
rect 15562 628398 15646 628634
rect 15882 628398 51326 628634
rect 51562 628398 51646 628634
rect 51882 628398 87326 628634
rect 87562 628398 87646 628634
rect 87882 628398 123326 628634
rect 123562 628398 123646 628634
rect 123882 628398 159326 628634
rect 159562 628398 159646 628634
rect 159882 628398 195326 628634
rect 195562 628398 195646 628634
rect 195882 628398 231326 628634
rect 231562 628398 231646 628634
rect 231882 628398 267326 628634
rect 267562 628398 267646 628634
rect 267882 628398 303326 628634
rect 303562 628398 303646 628634
rect 303882 628398 339326 628634
rect 339562 628398 339646 628634
rect 339882 628398 375326 628634
rect 375562 628398 375646 628634
rect 375882 628398 411326 628634
rect 411562 628398 411646 628634
rect 411882 628398 447326 628634
rect 447562 628398 447646 628634
rect 447882 628398 483326 628634
rect 483562 628398 483646 628634
rect 483882 628398 519326 628634
rect 519562 628398 519646 628634
rect 519882 628398 555326 628634
rect 555562 628398 555646 628634
rect 555882 628398 588222 628634
rect 588458 628398 588542 628634
rect 588778 628398 592650 628634
rect -8726 628366 592650 628398
rect -8726 624454 592650 624486
rect -8726 624218 -3894 624454
rect -3658 624218 -3574 624454
rect -3338 624218 10826 624454
rect 11062 624218 11146 624454
rect 11382 624218 46826 624454
rect 47062 624218 47146 624454
rect 47382 624218 82826 624454
rect 83062 624218 83146 624454
rect 83382 624218 118826 624454
rect 119062 624218 119146 624454
rect 119382 624218 154826 624454
rect 155062 624218 155146 624454
rect 155382 624218 190826 624454
rect 191062 624218 191146 624454
rect 191382 624218 226826 624454
rect 227062 624218 227146 624454
rect 227382 624218 262826 624454
rect 263062 624218 263146 624454
rect 263382 624218 298826 624454
rect 299062 624218 299146 624454
rect 299382 624218 334826 624454
rect 335062 624218 335146 624454
rect 335382 624218 370826 624454
rect 371062 624218 371146 624454
rect 371382 624218 406826 624454
rect 407062 624218 407146 624454
rect 407382 624218 442826 624454
rect 443062 624218 443146 624454
rect 443382 624218 478826 624454
rect 479062 624218 479146 624454
rect 479382 624218 514826 624454
rect 515062 624218 515146 624454
rect 515382 624218 550826 624454
rect 551062 624218 551146 624454
rect 551382 624218 587262 624454
rect 587498 624218 587582 624454
rect 587818 624218 592650 624454
rect -8726 624134 592650 624218
rect -8726 623898 -3894 624134
rect -3658 623898 -3574 624134
rect -3338 623898 10826 624134
rect 11062 623898 11146 624134
rect 11382 623898 46826 624134
rect 47062 623898 47146 624134
rect 47382 623898 82826 624134
rect 83062 623898 83146 624134
rect 83382 623898 118826 624134
rect 119062 623898 119146 624134
rect 119382 623898 154826 624134
rect 155062 623898 155146 624134
rect 155382 623898 190826 624134
rect 191062 623898 191146 624134
rect 191382 623898 226826 624134
rect 227062 623898 227146 624134
rect 227382 623898 262826 624134
rect 263062 623898 263146 624134
rect 263382 623898 298826 624134
rect 299062 623898 299146 624134
rect 299382 623898 334826 624134
rect 335062 623898 335146 624134
rect 335382 623898 370826 624134
rect 371062 623898 371146 624134
rect 371382 623898 406826 624134
rect 407062 623898 407146 624134
rect 407382 623898 442826 624134
rect 443062 623898 443146 624134
rect 443382 623898 478826 624134
rect 479062 623898 479146 624134
rect 479382 623898 514826 624134
rect 515062 623898 515146 624134
rect 515382 623898 550826 624134
rect 551062 623898 551146 624134
rect 551382 623898 587262 624134
rect 587498 623898 587582 624134
rect 587818 623898 592650 624134
rect -8726 623866 592650 623898
rect -8726 619954 592650 619986
rect -8726 619718 -2934 619954
rect -2698 619718 -2614 619954
rect -2378 619718 6326 619954
rect 6562 619718 6646 619954
rect 6882 619718 42326 619954
rect 42562 619718 42646 619954
rect 42882 619718 78326 619954
rect 78562 619718 78646 619954
rect 78882 619718 114326 619954
rect 114562 619718 114646 619954
rect 114882 619718 150326 619954
rect 150562 619718 150646 619954
rect 150882 619718 186326 619954
rect 186562 619718 186646 619954
rect 186882 619718 222326 619954
rect 222562 619718 222646 619954
rect 222882 619718 258326 619954
rect 258562 619718 258646 619954
rect 258882 619718 294326 619954
rect 294562 619718 294646 619954
rect 294882 619718 330326 619954
rect 330562 619718 330646 619954
rect 330882 619718 366326 619954
rect 366562 619718 366646 619954
rect 366882 619718 402326 619954
rect 402562 619718 402646 619954
rect 402882 619718 438326 619954
rect 438562 619718 438646 619954
rect 438882 619718 474326 619954
rect 474562 619718 474646 619954
rect 474882 619718 510326 619954
rect 510562 619718 510646 619954
rect 510882 619718 546326 619954
rect 546562 619718 546646 619954
rect 546882 619718 582326 619954
rect 582562 619718 582646 619954
rect 582882 619718 586302 619954
rect 586538 619718 586622 619954
rect 586858 619718 592650 619954
rect -8726 619634 592650 619718
rect -8726 619398 -2934 619634
rect -2698 619398 -2614 619634
rect -2378 619398 6326 619634
rect 6562 619398 6646 619634
rect 6882 619398 42326 619634
rect 42562 619398 42646 619634
rect 42882 619398 78326 619634
rect 78562 619398 78646 619634
rect 78882 619398 114326 619634
rect 114562 619398 114646 619634
rect 114882 619398 150326 619634
rect 150562 619398 150646 619634
rect 150882 619398 186326 619634
rect 186562 619398 186646 619634
rect 186882 619398 222326 619634
rect 222562 619398 222646 619634
rect 222882 619398 258326 619634
rect 258562 619398 258646 619634
rect 258882 619398 294326 619634
rect 294562 619398 294646 619634
rect 294882 619398 330326 619634
rect 330562 619398 330646 619634
rect 330882 619398 366326 619634
rect 366562 619398 366646 619634
rect 366882 619398 402326 619634
rect 402562 619398 402646 619634
rect 402882 619398 438326 619634
rect 438562 619398 438646 619634
rect 438882 619398 474326 619634
rect 474562 619398 474646 619634
rect 474882 619398 510326 619634
rect 510562 619398 510646 619634
rect 510882 619398 546326 619634
rect 546562 619398 546646 619634
rect 546882 619398 582326 619634
rect 582562 619398 582646 619634
rect 582882 619398 586302 619634
rect 586538 619398 586622 619634
rect 586858 619398 592650 619634
rect -8726 619366 592650 619398
rect -8726 615454 592650 615486
rect -8726 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 73826 615454
rect 74062 615218 74146 615454
rect 74382 615218 109826 615454
rect 110062 615218 110146 615454
rect 110382 615218 145826 615454
rect 146062 615218 146146 615454
rect 146382 615218 181826 615454
rect 182062 615218 182146 615454
rect 182382 615218 217826 615454
rect 218062 615218 218146 615454
rect 218382 615218 253826 615454
rect 254062 615218 254146 615454
rect 254382 615218 289826 615454
rect 290062 615218 290146 615454
rect 290382 615218 325826 615454
rect 326062 615218 326146 615454
rect 326382 615218 361826 615454
rect 362062 615218 362146 615454
rect 362382 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 469826 615454
rect 470062 615218 470146 615454
rect 470382 615218 505826 615454
rect 506062 615218 506146 615454
rect 506382 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 592650 615454
rect -8726 615134 592650 615218
rect -8726 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 73826 615134
rect 74062 614898 74146 615134
rect 74382 614898 109826 615134
rect 110062 614898 110146 615134
rect 110382 614898 145826 615134
rect 146062 614898 146146 615134
rect 146382 614898 181826 615134
rect 182062 614898 182146 615134
rect 182382 614898 217826 615134
rect 218062 614898 218146 615134
rect 218382 614898 253826 615134
rect 254062 614898 254146 615134
rect 254382 614898 289826 615134
rect 290062 614898 290146 615134
rect 290382 614898 325826 615134
rect 326062 614898 326146 615134
rect 326382 614898 361826 615134
rect 362062 614898 362146 615134
rect 362382 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 469826 615134
rect 470062 614898 470146 615134
rect 470382 614898 505826 615134
rect 506062 614898 506146 615134
rect 506382 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 592650 615134
rect -8726 614866 592650 614898
rect -8726 610954 592650 610986
rect -8726 610718 -8694 610954
rect -8458 610718 -8374 610954
rect -8138 610718 33326 610954
rect 33562 610718 33646 610954
rect 33882 610718 69326 610954
rect 69562 610718 69646 610954
rect 69882 610718 105326 610954
rect 105562 610718 105646 610954
rect 105882 610718 141326 610954
rect 141562 610718 141646 610954
rect 141882 610718 177326 610954
rect 177562 610718 177646 610954
rect 177882 610718 213326 610954
rect 213562 610718 213646 610954
rect 213882 610718 249326 610954
rect 249562 610718 249646 610954
rect 249882 610718 285326 610954
rect 285562 610718 285646 610954
rect 285882 610718 321326 610954
rect 321562 610718 321646 610954
rect 321882 610718 357326 610954
rect 357562 610718 357646 610954
rect 357882 610718 393326 610954
rect 393562 610718 393646 610954
rect 393882 610718 429326 610954
rect 429562 610718 429646 610954
rect 429882 610718 465326 610954
rect 465562 610718 465646 610954
rect 465882 610718 501326 610954
rect 501562 610718 501646 610954
rect 501882 610718 537326 610954
rect 537562 610718 537646 610954
rect 537882 610718 573326 610954
rect 573562 610718 573646 610954
rect 573882 610718 592062 610954
rect 592298 610718 592382 610954
rect 592618 610718 592650 610954
rect -8726 610634 592650 610718
rect -8726 610398 -8694 610634
rect -8458 610398 -8374 610634
rect -8138 610398 33326 610634
rect 33562 610398 33646 610634
rect 33882 610398 69326 610634
rect 69562 610398 69646 610634
rect 69882 610398 105326 610634
rect 105562 610398 105646 610634
rect 105882 610398 141326 610634
rect 141562 610398 141646 610634
rect 141882 610398 177326 610634
rect 177562 610398 177646 610634
rect 177882 610398 213326 610634
rect 213562 610398 213646 610634
rect 213882 610398 249326 610634
rect 249562 610398 249646 610634
rect 249882 610398 285326 610634
rect 285562 610398 285646 610634
rect 285882 610398 321326 610634
rect 321562 610398 321646 610634
rect 321882 610398 357326 610634
rect 357562 610398 357646 610634
rect 357882 610398 393326 610634
rect 393562 610398 393646 610634
rect 393882 610398 429326 610634
rect 429562 610398 429646 610634
rect 429882 610398 465326 610634
rect 465562 610398 465646 610634
rect 465882 610398 501326 610634
rect 501562 610398 501646 610634
rect 501882 610398 537326 610634
rect 537562 610398 537646 610634
rect 537882 610398 573326 610634
rect 573562 610398 573646 610634
rect 573882 610398 592062 610634
rect 592298 610398 592382 610634
rect 592618 610398 592650 610634
rect -8726 610366 592650 610398
rect -8726 606454 592650 606486
rect -8726 606218 -7734 606454
rect -7498 606218 -7414 606454
rect -7178 606218 28826 606454
rect 29062 606218 29146 606454
rect 29382 606218 64826 606454
rect 65062 606218 65146 606454
rect 65382 606218 100826 606454
rect 101062 606218 101146 606454
rect 101382 606218 136826 606454
rect 137062 606218 137146 606454
rect 137382 606218 172826 606454
rect 173062 606218 173146 606454
rect 173382 606218 208826 606454
rect 209062 606218 209146 606454
rect 209382 606218 244826 606454
rect 245062 606218 245146 606454
rect 245382 606218 280826 606454
rect 281062 606218 281146 606454
rect 281382 606218 316826 606454
rect 317062 606218 317146 606454
rect 317382 606218 352826 606454
rect 353062 606218 353146 606454
rect 353382 606218 388826 606454
rect 389062 606218 389146 606454
rect 389382 606218 424826 606454
rect 425062 606218 425146 606454
rect 425382 606218 460826 606454
rect 461062 606218 461146 606454
rect 461382 606218 496826 606454
rect 497062 606218 497146 606454
rect 497382 606218 532826 606454
rect 533062 606218 533146 606454
rect 533382 606218 568826 606454
rect 569062 606218 569146 606454
rect 569382 606218 591102 606454
rect 591338 606218 591422 606454
rect 591658 606218 592650 606454
rect -8726 606134 592650 606218
rect -8726 605898 -7734 606134
rect -7498 605898 -7414 606134
rect -7178 605898 28826 606134
rect 29062 605898 29146 606134
rect 29382 605898 64826 606134
rect 65062 605898 65146 606134
rect 65382 605898 100826 606134
rect 101062 605898 101146 606134
rect 101382 605898 136826 606134
rect 137062 605898 137146 606134
rect 137382 605898 172826 606134
rect 173062 605898 173146 606134
rect 173382 605898 208826 606134
rect 209062 605898 209146 606134
rect 209382 605898 244826 606134
rect 245062 605898 245146 606134
rect 245382 605898 280826 606134
rect 281062 605898 281146 606134
rect 281382 605898 316826 606134
rect 317062 605898 317146 606134
rect 317382 605898 352826 606134
rect 353062 605898 353146 606134
rect 353382 605898 388826 606134
rect 389062 605898 389146 606134
rect 389382 605898 424826 606134
rect 425062 605898 425146 606134
rect 425382 605898 460826 606134
rect 461062 605898 461146 606134
rect 461382 605898 496826 606134
rect 497062 605898 497146 606134
rect 497382 605898 532826 606134
rect 533062 605898 533146 606134
rect 533382 605898 568826 606134
rect 569062 605898 569146 606134
rect 569382 605898 591102 606134
rect 591338 605898 591422 606134
rect 591658 605898 592650 606134
rect -8726 605866 592650 605898
rect -8726 601954 592650 601986
rect -8726 601718 -6774 601954
rect -6538 601718 -6454 601954
rect -6218 601718 24326 601954
rect 24562 601718 24646 601954
rect 24882 601718 60326 601954
rect 60562 601718 60646 601954
rect 60882 601718 96326 601954
rect 96562 601718 96646 601954
rect 96882 601718 132326 601954
rect 132562 601718 132646 601954
rect 132882 601718 168326 601954
rect 168562 601718 168646 601954
rect 168882 601718 204326 601954
rect 204562 601718 204646 601954
rect 204882 601718 240326 601954
rect 240562 601718 240646 601954
rect 240882 601718 276326 601954
rect 276562 601718 276646 601954
rect 276882 601718 312326 601954
rect 312562 601718 312646 601954
rect 312882 601718 348326 601954
rect 348562 601718 348646 601954
rect 348882 601718 384326 601954
rect 384562 601718 384646 601954
rect 384882 601718 420326 601954
rect 420562 601718 420646 601954
rect 420882 601718 456326 601954
rect 456562 601718 456646 601954
rect 456882 601718 492326 601954
rect 492562 601718 492646 601954
rect 492882 601718 528326 601954
rect 528562 601718 528646 601954
rect 528882 601718 564326 601954
rect 564562 601718 564646 601954
rect 564882 601718 590142 601954
rect 590378 601718 590462 601954
rect 590698 601718 592650 601954
rect -8726 601634 592650 601718
rect -8726 601398 -6774 601634
rect -6538 601398 -6454 601634
rect -6218 601398 24326 601634
rect 24562 601398 24646 601634
rect 24882 601398 60326 601634
rect 60562 601398 60646 601634
rect 60882 601398 96326 601634
rect 96562 601398 96646 601634
rect 96882 601398 132326 601634
rect 132562 601398 132646 601634
rect 132882 601398 168326 601634
rect 168562 601398 168646 601634
rect 168882 601398 204326 601634
rect 204562 601398 204646 601634
rect 204882 601398 240326 601634
rect 240562 601398 240646 601634
rect 240882 601398 276326 601634
rect 276562 601398 276646 601634
rect 276882 601398 312326 601634
rect 312562 601398 312646 601634
rect 312882 601398 348326 601634
rect 348562 601398 348646 601634
rect 348882 601398 384326 601634
rect 384562 601398 384646 601634
rect 384882 601398 420326 601634
rect 420562 601398 420646 601634
rect 420882 601398 456326 601634
rect 456562 601398 456646 601634
rect 456882 601398 492326 601634
rect 492562 601398 492646 601634
rect 492882 601398 528326 601634
rect 528562 601398 528646 601634
rect 528882 601398 564326 601634
rect 564562 601398 564646 601634
rect 564882 601398 590142 601634
rect 590378 601398 590462 601634
rect 590698 601398 592650 601634
rect -8726 601366 592650 601398
rect -8726 597454 592650 597486
rect -8726 597218 -5814 597454
rect -5578 597218 -5494 597454
rect -5258 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 55826 597454
rect 56062 597218 56146 597454
rect 56382 597218 91826 597454
rect 92062 597218 92146 597454
rect 92382 597218 127826 597454
rect 128062 597218 128146 597454
rect 128382 597218 163826 597454
rect 164062 597218 164146 597454
rect 164382 597218 199826 597454
rect 200062 597218 200146 597454
rect 200382 597218 235826 597454
rect 236062 597218 236146 597454
rect 236382 597218 271826 597454
rect 272062 597218 272146 597454
rect 272382 597218 307826 597454
rect 308062 597218 308146 597454
rect 308382 597218 343826 597454
rect 344062 597218 344146 597454
rect 344382 597218 379826 597454
rect 380062 597218 380146 597454
rect 380382 597218 415826 597454
rect 416062 597218 416146 597454
rect 416382 597218 451826 597454
rect 452062 597218 452146 597454
rect 452382 597218 487826 597454
rect 488062 597218 488146 597454
rect 488382 597218 523826 597454
rect 524062 597218 524146 597454
rect 524382 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 589182 597454
rect 589418 597218 589502 597454
rect 589738 597218 592650 597454
rect -8726 597134 592650 597218
rect -8726 596898 -5814 597134
rect -5578 596898 -5494 597134
rect -5258 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 55826 597134
rect 56062 596898 56146 597134
rect 56382 596898 91826 597134
rect 92062 596898 92146 597134
rect 92382 596898 127826 597134
rect 128062 596898 128146 597134
rect 128382 596898 163826 597134
rect 164062 596898 164146 597134
rect 164382 596898 199826 597134
rect 200062 596898 200146 597134
rect 200382 596898 235826 597134
rect 236062 596898 236146 597134
rect 236382 596898 271826 597134
rect 272062 596898 272146 597134
rect 272382 596898 307826 597134
rect 308062 596898 308146 597134
rect 308382 596898 343826 597134
rect 344062 596898 344146 597134
rect 344382 596898 379826 597134
rect 380062 596898 380146 597134
rect 380382 596898 415826 597134
rect 416062 596898 416146 597134
rect 416382 596898 451826 597134
rect 452062 596898 452146 597134
rect 452382 596898 487826 597134
rect 488062 596898 488146 597134
rect 488382 596898 523826 597134
rect 524062 596898 524146 597134
rect 524382 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 589182 597134
rect 589418 596898 589502 597134
rect 589738 596898 592650 597134
rect -8726 596866 592650 596898
rect -8726 592954 592650 592986
rect -8726 592718 -4854 592954
rect -4618 592718 -4534 592954
rect -4298 592718 15326 592954
rect 15562 592718 15646 592954
rect 15882 592718 51326 592954
rect 51562 592718 51646 592954
rect 51882 592718 87326 592954
rect 87562 592718 87646 592954
rect 87882 592718 123326 592954
rect 123562 592718 123646 592954
rect 123882 592718 159326 592954
rect 159562 592718 159646 592954
rect 159882 592718 195326 592954
rect 195562 592718 195646 592954
rect 195882 592718 231326 592954
rect 231562 592718 231646 592954
rect 231882 592718 267326 592954
rect 267562 592718 267646 592954
rect 267882 592718 303326 592954
rect 303562 592718 303646 592954
rect 303882 592718 339326 592954
rect 339562 592718 339646 592954
rect 339882 592718 375326 592954
rect 375562 592718 375646 592954
rect 375882 592718 411326 592954
rect 411562 592718 411646 592954
rect 411882 592718 447326 592954
rect 447562 592718 447646 592954
rect 447882 592718 483326 592954
rect 483562 592718 483646 592954
rect 483882 592718 519326 592954
rect 519562 592718 519646 592954
rect 519882 592718 555326 592954
rect 555562 592718 555646 592954
rect 555882 592718 588222 592954
rect 588458 592718 588542 592954
rect 588778 592718 592650 592954
rect -8726 592634 592650 592718
rect -8726 592398 -4854 592634
rect -4618 592398 -4534 592634
rect -4298 592398 15326 592634
rect 15562 592398 15646 592634
rect 15882 592398 51326 592634
rect 51562 592398 51646 592634
rect 51882 592398 87326 592634
rect 87562 592398 87646 592634
rect 87882 592398 123326 592634
rect 123562 592398 123646 592634
rect 123882 592398 159326 592634
rect 159562 592398 159646 592634
rect 159882 592398 195326 592634
rect 195562 592398 195646 592634
rect 195882 592398 231326 592634
rect 231562 592398 231646 592634
rect 231882 592398 267326 592634
rect 267562 592398 267646 592634
rect 267882 592398 303326 592634
rect 303562 592398 303646 592634
rect 303882 592398 339326 592634
rect 339562 592398 339646 592634
rect 339882 592398 375326 592634
rect 375562 592398 375646 592634
rect 375882 592398 411326 592634
rect 411562 592398 411646 592634
rect 411882 592398 447326 592634
rect 447562 592398 447646 592634
rect 447882 592398 483326 592634
rect 483562 592398 483646 592634
rect 483882 592398 519326 592634
rect 519562 592398 519646 592634
rect 519882 592398 555326 592634
rect 555562 592398 555646 592634
rect 555882 592398 588222 592634
rect 588458 592398 588542 592634
rect 588778 592398 592650 592634
rect -8726 592366 592650 592398
rect -8726 588454 592650 588486
rect -8726 588218 -3894 588454
rect -3658 588218 -3574 588454
rect -3338 588218 10826 588454
rect 11062 588218 11146 588454
rect 11382 588218 46826 588454
rect 47062 588218 47146 588454
rect 47382 588218 82826 588454
rect 83062 588218 83146 588454
rect 83382 588218 118826 588454
rect 119062 588218 119146 588454
rect 119382 588218 154826 588454
rect 155062 588218 155146 588454
rect 155382 588218 190826 588454
rect 191062 588218 191146 588454
rect 191382 588218 226826 588454
rect 227062 588218 227146 588454
rect 227382 588218 262826 588454
rect 263062 588218 263146 588454
rect 263382 588218 298826 588454
rect 299062 588218 299146 588454
rect 299382 588218 334826 588454
rect 335062 588218 335146 588454
rect 335382 588218 370826 588454
rect 371062 588218 371146 588454
rect 371382 588218 406826 588454
rect 407062 588218 407146 588454
rect 407382 588218 442826 588454
rect 443062 588218 443146 588454
rect 443382 588218 478826 588454
rect 479062 588218 479146 588454
rect 479382 588218 514826 588454
rect 515062 588218 515146 588454
rect 515382 588218 550826 588454
rect 551062 588218 551146 588454
rect 551382 588218 587262 588454
rect 587498 588218 587582 588454
rect 587818 588218 592650 588454
rect -8726 588134 592650 588218
rect -8726 587898 -3894 588134
rect -3658 587898 -3574 588134
rect -3338 587898 10826 588134
rect 11062 587898 11146 588134
rect 11382 587898 46826 588134
rect 47062 587898 47146 588134
rect 47382 587898 82826 588134
rect 83062 587898 83146 588134
rect 83382 587898 118826 588134
rect 119062 587898 119146 588134
rect 119382 587898 154826 588134
rect 155062 587898 155146 588134
rect 155382 587898 190826 588134
rect 191062 587898 191146 588134
rect 191382 587898 226826 588134
rect 227062 587898 227146 588134
rect 227382 587898 262826 588134
rect 263062 587898 263146 588134
rect 263382 587898 298826 588134
rect 299062 587898 299146 588134
rect 299382 587898 334826 588134
rect 335062 587898 335146 588134
rect 335382 587898 370826 588134
rect 371062 587898 371146 588134
rect 371382 587898 406826 588134
rect 407062 587898 407146 588134
rect 407382 587898 442826 588134
rect 443062 587898 443146 588134
rect 443382 587898 478826 588134
rect 479062 587898 479146 588134
rect 479382 587898 514826 588134
rect 515062 587898 515146 588134
rect 515382 587898 550826 588134
rect 551062 587898 551146 588134
rect 551382 587898 587262 588134
rect 587498 587898 587582 588134
rect 587818 587898 592650 588134
rect -8726 587866 592650 587898
rect -8726 583954 592650 583986
rect -8726 583718 -2934 583954
rect -2698 583718 -2614 583954
rect -2378 583718 6326 583954
rect 6562 583718 6646 583954
rect 6882 583718 42326 583954
rect 42562 583718 42646 583954
rect 42882 583718 78326 583954
rect 78562 583718 78646 583954
rect 78882 583718 114326 583954
rect 114562 583718 114646 583954
rect 114882 583718 150326 583954
rect 150562 583718 150646 583954
rect 150882 583718 186326 583954
rect 186562 583718 186646 583954
rect 186882 583718 222326 583954
rect 222562 583718 222646 583954
rect 222882 583718 258326 583954
rect 258562 583718 258646 583954
rect 258882 583718 294326 583954
rect 294562 583718 294646 583954
rect 294882 583718 330326 583954
rect 330562 583718 330646 583954
rect 330882 583718 366326 583954
rect 366562 583718 366646 583954
rect 366882 583718 402326 583954
rect 402562 583718 402646 583954
rect 402882 583718 438326 583954
rect 438562 583718 438646 583954
rect 438882 583718 474326 583954
rect 474562 583718 474646 583954
rect 474882 583718 510326 583954
rect 510562 583718 510646 583954
rect 510882 583718 546326 583954
rect 546562 583718 546646 583954
rect 546882 583718 582326 583954
rect 582562 583718 582646 583954
rect 582882 583718 586302 583954
rect 586538 583718 586622 583954
rect 586858 583718 592650 583954
rect -8726 583634 592650 583718
rect -8726 583398 -2934 583634
rect -2698 583398 -2614 583634
rect -2378 583398 6326 583634
rect 6562 583398 6646 583634
rect 6882 583398 42326 583634
rect 42562 583398 42646 583634
rect 42882 583398 78326 583634
rect 78562 583398 78646 583634
rect 78882 583398 114326 583634
rect 114562 583398 114646 583634
rect 114882 583398 150326 583634
rect 150562 583398 150646 583634
rect 150882 583398 186326 583634
rect 186562 583398 186646 583634
rect 186882 583398 222326 583634
rect 222562 583398 222646 583634
rect 222882 583398 258326 583634
rect 258562 583398 258646 583634
rect 258882 583398 294326 583634
rect 294562 583398 294646 583634
rect 294882 583398 330326 583634
rect 330562 583398 330646 583634
rect 330882 583398 366326 583634
rect 366562 583398 366646 583634
rect 366882 583398 402326 583634
rect 402562 583398 402646 583634
rect 402882 583398 438326 583634
rect 438562 583398 438646 583634
rect 438882 583398 474326 583634
rect 474562 583398 474646 583634
rect 474882 583398 510326 583634
rect 510562 583398 510646 583634
rect 510882 583398 546326 583634
rect 546562 583398 546646 583634
rect 546882 583398 582326 583634
rect 582562 583398 582646 583634
rect 582882 583398 586302 583634
rect 586538 583398 586622 583634
rect 586858 583398 592650 583634
rect -8726 583366 592650 583398
rect -8726 579454 592650 579486
rect -8726 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 73826 579454
rect 74062 579218 74146 579454
rect 74382 579218 109826 579454
rect 110062 579218 110146 579454
rect 110382 579218 145826 579454
rect 146062 579218 146146 579454
rect 146382 579218 181826 579454
rect 182062 579218 182146 579454
rect 182382 579218 217826 579454
rect 218062 579218 218146 579454
rect 218382 579218 253826 579454
rect 254062 579218 254146 579454
rect 254382 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 325826 579454
rect 326062 579218 326146 579454
rect 326382 579218 361826 579454
rect 362062 579218 362146 579454
rect 362382 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 592650 579454
rect -8726 579134 592650 579218
rect -8726 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 73826 579134
rect 74062 578898 74146 579134
rect 74382 578898 109826 579134
rect 110062 578898 110146 579134
rect 110382 578898 145826 579134
rect 146062 578898 146146 579134
rect 146382 578898 181826 579134
rect 182062 578898 182146 579134
rect 182382 578898 217826 579134
rect 218062 578898 218146 579134
rect 218382 578898 253826 579134
rect 254062 578898 254146 579134
rect 254382 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 325826 579134
rect 326062 578898 326146 579134
rect 326382 578898 361826 579134
rect 362062 578898 362146 579134
rect 362382 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 592650 579134
rect -8726 578866 592650 578898
rect -8726 574954 592650 574986
rect -8726 574718 -8694 574954
rect -8458 574718 -8374 574954
rect -8138 574718 33326 574954
rect 33562 574718 33646 574954
rect 33882 574718 69326 574954
rect 69562 574718 69646 574954
rect 69882 574718 105326 574954
rect 105562 574718 105646 574954
rect 105882 574718 141326 574954
rect 141562 574718 141646 574954
rect 141882 574718 177326 574954
rect 177562 574718 177646 574954
rect 177882 574718 213326 574954
rect 213562 574718 213646 574954
rect 213882 574718 249326 574954
rect 249562 574718 249646 574954
rect 249882 574718 285326 574954
rect 285562 574718 285646 574954
rect 285882 574718 321326 574954
rect 321562 574718 321646 574954
rect 321882 574718 357326 574954
rect 357562 574718 357646 574954
rect 357882 574718 393326 574954
rect 393562 574718 393646 574954
rect 393882 574718 429326 574954
rect 429562 574718 429646 574954
rect 429882 574718 465326 574954
rect 465562 574718 465646 574954
rect 465882 574718 501326 574954
rect 501562 574718 501646 574954
rect 501882 574718 537326 574954
rect 537562 574718 537646 574954
rect 537882 574718 573326 574954
rect 573562 574718 573646 574954
rect 573882 574718 592062 574954
rect 592298 574718 592382 574954
rect 592618 574718 592650 574954
rect -8726 574634 592650 574718
rect -8726 574398 -8694 574634
rect -8458 574398 -8374 574634
rect -8138 574398 33326 574634
rect 33562 574398 33646 574634
rect 33882 574398 69326 574634
rect 69562 574398 69646 574634
rect 69882 574398 105326 574634
rect 105562 574398 105646 574634
rect 105882 574398 141326 574634
rect 141562 574398 141646 574634
rect 141882 574398 177326 574634
rect 177562 574398 177646 574634
rect 177882 574398 213326 574634
rect 213562 574398 213646 574634
rect 213882 574398 249326 574634
rect 249562 574398 249646 574634
rect 249882 574398 285326 574634
rect 285562 574398 285646 574634
rect 285882 574398 321326 574634
rect 321562 574398 321646 574634
rect 321882 574398 357326 574634
rect 357562 574398 357646 574634
rect 357882 574398 393326 574634
rect 393562 574398 393646 574634
rect 393882 574398 429326 574634
rect 429562 574398 429646 574634
rect 429882 574398 465326 574634
rect 465562 574398 465646 574634
rect 465882 574398 501326 574634
rect 501562 574398 501646 574634
rect 501882 574398 537326 574634
rect 537562 574398 537646 574634
rect 537882 574398 573326 574634
rect 573562 574398 573646 574634
rect 573882 574398 592062 574634
rect 592298 574398 592382 574634
rect 592618 574398 592650 574634
rect -8726 574366 592650 574398
rect -8726 570454 592650 570486
rect -8726 570218 -7734 570454
rect -7498 570218 -7414 570454
rect -7178 570218 28826 570454
rect 29062 570218 29146 570454
rect 29382 570218 64826 570454
rect 65062 570218 65146 570454
rect 65382 570218 100826 570454
rect 101062 570218 101146 570454
rect 101382 570218 136826 570454
rect 137062 570218 137146 570454
rect 137382 570218 172826 570454
rect 173062 570218 173146 570454
rect 173382 570218 208826 570454
rect 209062 570218 209146 570454
rect 209382 570218 244826 570454
rect 245062 570218 245146 570454
rect 245382 570218 280826 570454
rect 281062 570218 281146 570454
rect 281382 570218 316826 570454
rect 317062 570218 317146 570454
rect 317382 570218 352826 570454
rect 353062 570218 353146 570454
rect 353382 570218 388826 570454
rect 389062 570218 389146 570454
rect 389382 570218 424826 570454
rect 425062 570218 425146 570454
rect 425382 570218 460826 570454
rect 461062 570218 461146 570454
rect 461382 570218 496826 570454
rect 497062 570218 497146 570454
rect 497382 570218 532826 570454
rect 533062 570218 533146 570454
rect 533382 570218 568826 570454
rect 569062 570218 569146 570454
rect 569382 570218 591102 570454
rect 591338 570218 591422 570454
rect 591658 570218 592650 570454
rect -8726 570134 592650 570218
rect -8726 569898 -7734 570134
rect -7498 569898 -7414 570134
rect -7178 569898 28826 570134
rect 29062 569898 29146 570134
rect 29382 569898 64826 570134
rect 65062 569898 65146 570134
rect 65382 569898 100826 570134
rect 101062 569898 101146 570134
rect 101382 569898 136826 570134
rect 137062 569898 137146 570134
rect 137382 569898 172826 570134
rect 173062 569898 173146 570134
rect 173382 569898 208826 570134
rect 209062 569898 209146 570134
rect 209382 569898 244826 570134
rect 245062 569898 245146 570134
rect 245382 569898 280826 570134
rect 281062 569898 281146 570134
rect 281382 569898 316826 570134
rect 317062 569898 317146 570134
rect 317382 569898 352826 570134
rect 353062 569898 353146 570134
rect 353382 569898 388826 570134
rect 389062 569898 389146 570134
rect 389382 569898 424826 570134
rect 425062 569898 425146 570134
rect 425382 569898 460826 570134
rect 461062 569898 461146 570134
rect 461382 569898 496826 570134
rect 497062 569898 497146 570134
rect 497382 569898 532826 570134
rect 533062 569898 533146 570134
rect 533382 569898 568826 570134
rect 569062 569898 569146 570134
rect 569382 569898 591102 570134
rect 591338 569898 591422 570134
rect 591658 569898 592650 570134
rect -8726 569866 592650 569898
rect -8726 565954 592650 565986
rect -8726 565718 -6774 565954
rect -6538 565718 -6454 565954
rect -6218 565718 24326 565954
rect 24562 565718 24646 565954
rect 24882 565718 60326 565954
rect 60562 565718 60646 565954
rect 60882 565718 96326 565954
rect 96562 565718 96646 565954
rect 96882 565718 132326 565954
rect 132562 565718 132646 565954
rect 132882 565718 168326 565954
rect 168562 565718 168646 565954
rect 168882 565718 204326 565954
rect 204562 565718 204646 565954
rect 204882 565718 240326 565954
rect 240562 565718 240646 565954
rect 240882 565718 276326 565954
rect 276562 565718 276646 565954
rect 276882 565718 312326 565954
rect 312562 565718 312646 565954
rect 312882 565718 348326 565954
rect 348562 565718 348646 565954
rect 348882 565718 384326 565954
rect 384562 565718 384646 565954
rect 384882 565718 420326 565954
rect 420562 565718 420646 565954
rect 420882 565718 456326 565954
rect 456562 565718 456646 565954
rect 456882 565718 492326 565954
rect 492562 565718 492646 565954
rect 492882 565718 528326 565954
rect 528562 565718 528646 565954
rect 528882 565718 564326 565954
rect 564562 565718 564646 565954
rect 564882 565718 590142 565954
rect 590378 565718 590462 565954
rect 590698 565718 592650 565954
rect -8726 565634 592650 565718
rect -8726 565398 -6774 565634
rect -6538 565398 -6454 565634
rect -6218 565398 24326 565634
rect 24562 565398 24646 565634
rect 24882 565398 60326 565634
rect 60562 565398 60646 565634
rect 60882 565398 96326 565634
rect 96562 565398 96646 565634
rect 96882 565398 132326 565634
rect 132562 565398 132646 565634
rect 132882 565398 168326 565634
rect 168562 565398 168646 565634
rect 168882 565398 204326 565634
rect 204562 565398 204646 565634
rect 204882 565398 240326 565634
rect 240562 565398 240646 565634
rect 240882 565398 276326 565634
rect 276562 565398 276646 565634
rect 276882 565398 312326 565634
rect 312562 565398 312646 565634
rect 312882 565398 348326 565634
rect 348562 565398 348646 565634
rect 348882 565398 384326 565634
rect 384562 565398 384646 565634
rect 384882 565398 420326 565634
rect 420562 565398 420646 565634
rect 420882 565398 456326 565634
rect 456562 565398 456646 565634
rect 456882 565398 492326 565634
rect 492562 565398 492646 565634
rect 492882 565398 528326 565634
rect 528562 565398 528646 565634
rect 528882 565398 564326 565634
rect 564562 565398 564646 565634
rect 564882 565398 590142 565634
rect 590378 565398 590462 565634
rect 590698 565398 592650 565634
rect -8726 565366 592650 565398
rect -8726 561454 592650 561486
rect -8726 561218 -5814 561454
rect -5578 561218 -5494 561454
rect -5258 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 55826 561454
rect 56062 561218 56146 561454
rect 56382 561218 91826 561454
rect 92062 561218 92146 561454
rect 92382 561218 127826 561454
rect 128062 561218 128146 561454
rect 128382 561218 163826 561454
rect 164062 561218 164146 561454
rect 164382 561218 199826 561454
rect 200062 561218 200146 561454
rect 200382 561218 235826 561454
rect 236062 561218 236146 561454
rect 236382 561218 271826 561454
rect 272062 561218 272146 561454
rect 272382 561218 307826 561454
rect 308062 561218 308146 561454
rect 308382 561218 343826 561454
rect 344062 561218 344146 561454
rect 344382 561218 379826 561454
rect 380062 561218 380146 561454
rect 380382 561218 415826 561454
rect 416062 561218 416146 561454
rect 416382 561218 451826 561454
rect 452062 561218 452146 561454
rect 452382 561218 487826 561454
rect 488062 561218 488146 561454
rect 488382 561218 523826 561454
rect 524062 561218 524146 561454
rect 524382 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 589182 561454
rect 589418 561218 589502 561454
rect 589738 561218 592650 561454
rect -8726 561134 592650 561218
rect -8726 560898 -5814 561134
rect -5578 560898 -5494 561134
rect -5258 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 55826 561134
rect 56062 560898 56146 561134
rect 56382 560898 91826 561134
rect 92062 560898 92146 561134
rect 92382 560898 127826 561134
rect 128062 560898 128146 561134
rect 128382 560898 163826 561134
rect 164062 560898 164146 561134
rect 164382 560898 199826 561134
rect 200062 560898 200146 561134
rect 200382 560898 235826 561134
rect 236062 560898 236146 561134
rect 236382 560898 271826 561134
rect 272062 560898 272146 561134
rect 272382 560898 307826 561134
rect 308062 560898 308146 561134
rect 308382 560898 343826 561134
rect 344062 560898 344146 561134
rect 344382 560898 379826 561134
rect 380062 560898 380146 561134
rect 380382 560898 415826 561134
rect 416062 560898 416146 561134
rect 416382 560898 451826 561134
rect 452062 560898 452146 561134
rect 452382 560898 487826 561134
rect 488062 560898 488146 561134
rect 488382 560898 523826 561134
rect 524062 560898 524146 561134
rect 524382 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 589182 561134
rect 589418 560898 589502 561134
rect 589738 560898 592650 561134
rect -8726 560866 592650 560898
rect -8726 556954 592650 556986
rect -8726 556718 -4854 556954
rect -4618 556718 -4534 556954
rect -4298 556718 15326 556954
rect 15562 556718 15646 556954
rect 15882 556718 51326 556954
rect 51562 556718 51646 556954
rect 51882 556718 87326 556954
rect 87562 556718 87646 556954
rect 87882 556718 123326 556954
rect 123562 556718 123646 556954
rect 123882 556718 159326 556954
rect 159562 556718 159646 556954
rect 159882 556718 195326 556954
rect 195562 556718 195646 556954
rect 195882 556718 231326 556954
rect 231562 556718 231646 556954
rect 231882 556718 267326 556954
rect 267562 556718 267646 556954
rect 267882 556718 303326 556954
rect 303562 556718 303646 556954
rect 303882 556718 339326 556954
rect 339562 556718 339646 556954
rect 339882 556718 375326 556954
rect 375562 556718 375646 556954
rect 375882 556718 411326 556954
rect 411562 556718 411646 556954
rect 411882 556718 447326 556954
rect 447562 556718 447646 556954
rect 447882 556718 483326 556954
rect 483562 556718 483646 556954
rect 483882 556718 519326 556954
rect 519562 556718 519646 556954
rect 519882 556718 555326 556954
rect 555562 556718 555646 556954
rect 555882 556718 588222 556954
rect 588458 556718 588542 556954
rect 588778 556718 592650 556954
rect -8726 556634 592650 556718
rect -8726 556398 -4854 556634
rect -4618 556398 -4534 556634
rect -4298 556398 15326 556634
rect 15562 556398 15646 556634
rect 15882 556398 51326 556634
rect 51562 556398 51646 556634
rect 51882 556398 87326 556634
rect 87562 556398 87646 556634
rect 87882 556398 123326 556634
rect 123562 556398 123646 556634
rect 123882 556398 159326 556634
rect 159562 556398 159646 556634
rect 159882 556398 195326 556634
rect 195562 556398 195646 556634
rect 195882 556398 231326 556634
rect 231562 556398 231646 556634
rect 231882 556398 267326 556634
rect 267562 556398 267646 556634
rect 267882 556398 303326 556634
rect 303562 556398 303646 556634
rect 303882 556398 339326 556634
rect 339562 556398 339646 556634
rect 339882 556398 375326 556634
rect 375562 556398 375646 556634
rect 375882 556398 411326 556634
rect 411562 556398 411646 556634
rect 411882 556398 447326 556634
rect 447562 556398 447646 556634
rect 447882 556398 483326 556634
rect 483562 556398 483646 556634
rect 483882 556398 519326 556634
rect 519562 556398 519646 556634
rect 519882 556398 555326 556634
rect 555562 556398 555646 556634
rect 555882 556398 588222 556634
rect 588458 556398 588542 556634
rect 588778 556398 592650 556634
rect -8726 556366 592650 556398
rect -8726 552454 592650 552486
rect -8726 552218 -3894 552454
rect -3658 552218 -3574 552454
rect -3338 552218 10826 552454
rect 11062 552218 11146 552454
rect 11382 552218 46826 552454
rect 47062 552218 47146 552454
rect 47382 552218 82826 552454
rect 83062 552218 83146 552454
rect 83382 552218 118826 552454
rect 119062 552218 119146 552454
rect 119382 552218 154826 552454
rect 155062 552218 155146 552454
rect 155382 552218 190826 552454
rect 191062 552218 191146 552454
rect 191382 552218 226826 552454
rect 227062 552218 227146 552454
rect 227382 552218 262826 552454
rect 263062 552218 263146 552454
rect 263382 552218 298826 552454
rect 299062 552218 299146 552454
rect 299382 552218 334826 552454
rect 335062 552218 335146 552454
rect 335382 552218 370826 552454
rect 371062 552218 371146 552454
rect 371382 552218 406826 552454
rect 407062 552218 407146 552454
rect 407382 552218 442826 552454
rect 443062 552218 443146 552454
rect 443382 552218 478826 552454
rect 479062 552218 479146 552454
rect 479382 552218 514826 552454
rect 515062 552218 515146 552454
rect 515382 552218 550826 552454
rect 551062 552218 551146 552454
rect 551382 552218 587262 552454
rect 587498 552218 587582 552454
rect 587818 552218 592650 552454
rect -8726 552134 592650 552218
rect -8726 551898 -3894 552134
rect -3658 551898 -3574 552134
rect -3338 551898 10826 552134
rect 11062 551898 11146 552134
rect 11382 551898 46826 552134
rect 47062 551898 47146 552134
rect 47382 551898 82826 552134
rect 83062 551898 83146 552134
rect 83382 551898 118826 552134
rect 119062 551898 119146 552134
rect 119382 551898 154826 552134
rect 155062 551898 155146 552134
rect 155382 551898 190826 552134
rect 191062 551898 191146 552134
rect 191382 551898 226826 552134
rect 227062 551898 227146 552134
rect 227382 551898 262826 552134
rect 263062 551898 263146 552134
rect 263382 551898 298826 552134
rect 299062 551898 299146 552134
rect 299382 551898 334826 552134
rect 335062 551898 335146 552134
rect 335382 551898 370826 552134
rect 371062 551898 371146 552134
rect 371382 551898 406826 552134
rect 407062 551898 407146 552134
rect 407382 551898 442826 552134
rect 443062 551898 443146 552134
rect 443382 551898 478826 552134
rect 479062 551898 479146 552134
rect 479382 551898 514826 552134
rect 515062 551898 515146 552134
rect 515382 551898 550826 552134
rect 551062 551898 551146 552134
rect 551382 551898 587262 552134
rect 587498 551898 587582 552134
rect 587818 551898 592650 552134
rect -8726 551866 592650 551898
rect -8726 547954 592650 547986
rect -8726 547718 -2934 547954
rect -2698 547718 -2614 547954
rect -2378 547718 6326 547954
rect 6562 547718 6646 547954
rect 6882 547718 42326 547954
rect 42562 547718 42646 547954
rect 42882 547718 78326 547954
rect 78562 547718 78646 547954
rect 78882 547718 114326 547954
rect 114562 547718 114646 547954
rect 114882 547718 150326 547954
rect 150562 547718 150646 547954
rect 150882 547718 186326 547954
rect 186562 547718 186646 547954
rect 186882 547718 222326 547954
rect 222562 547718 222646 547954
rect 222882 547718 258326 547954
rect 258562 547718 258646 547954
rect 258882 547718 294326 547954
rect 294562 547718 294646 547954
rect 294882 547718 330326 547954
rect 330562 547718 330646 547954
rect 330882 547718 366326 547954
rect 366562 547718 366646 547954
rect 366882 547718 402326 547954
rect 402562 547718 402646 547954
rect 402882 547718 438326 547954
rect 438562 547718 438646 547954
rect 438882 547718 474326 547954
rect 474562 547718 474646 547954
rect 474882 547718 510326 547954
rect 510562 547718 510646 547954
rect 510882 547718 546326 547954
rect 546562 547718 546646 547954
rect 546882 547718 582326 547954
rect 582562 547718 582646 547954
rect 582882 547718 586302 547954
rect 586538 547718 586622 547954
rect 586858 547718 592650 547954
rect -8726 547634 592650 547718
rect -8726 547398 -2934 547634
rect -2698 547398 -2614 547634
rect -2378 547398 6326 547634
rect 6562 547398 6646 547634
rect 6882 547398 42326 547634
rect 42562 547398 42646 547634
rect 42882 547398 78326 547634
rect 78562 547398 78646 547634
rect 78882 547398 114326 547634
rect 114562 547398 114646 547634
rect 114882 547398 150326 547634
rect 150562 547398 150646 547634
rect 150882 547398 186326 547634
rect 186562 547398 186646 547634
rect 186882 547398 222326 547634
rect 222562 547398 222646 547634
rect 222882 547398 258326 547634
rect 258562 547398 258646 547634
rect 258882 547398 294326 547634
rect 294562 547398 294646 547634
rect 294882 547398 330326 547634
rect 330562 547398 330646 547634
rect 330882 547398 366326 547634
rect 366562 547398 366646 547634
rect 366882 547398 402326 547634
rect 402562 547398 402646 547634
rect 402882 547398 438326 547634
rect 438562 547398 438646 547634
rect 438882 547398 474326 547634
rect 474562 547398 474646 547634
rect 474882 547398 510326 547634
rect 510562 547398 510646 547634
rect 510882 547398 546326 547634
rect 546562 547398 546646 547634
rect 546882 547398 582326 547634
rect 582562 547398 582646 547634
rect 582882 547398 586302 547634
rect 586538 547398 586622 547634
rect 586858 547398 592650 547634
rect -8726 547366 592650 547398
rect -8726 543454 592650 543486
rect -8726 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 73826 543454
rect 74062 543218 74146 543454
rect 74382 543218 109826 543454
rect 110062 543218 110146 543454
rect 110382 543218 145826 543454
rect 146062 543218 146146 543454
rect 146382 543218 181826 543454
rect 182062 543218 182146 543454
rect 182382 543218 217826 543454
rect 218062 543218 218146 543454
rect 218382 543218 253826 543454
rect 254062 543218 254146 543454
rect 254382 543218 289826 543454
rect 290062 543218 290146 543454
rect 290382 543218 325826 543454
rect 326062 543218 326146 543454
rect 326382 543218 361826 543454
rect 362062 543218 362146 543454
rect 362382 543218 397826 543454
rect 398062 543218 398146 543454
rect 398382 543218 433826 543454
rect 434062 543218 434146 543454
rect 434382 543218 469826 543454
rect 470062 543218 470146 543454
rect 470382 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 592650 543454
rect -8726 543134 592650 543218
rect -8726 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 73826 543134
rect 74062 542898 74146 543134
rect 74382 542898 109826 543134
rect 110062 542898 110146 543134
rect 110382 542898 145826 543134
rect 146062 542898 146146 543134
rect 146382 542898 181826 543134
rect 182062 542898 182146 543134
rect 182382 542898 217826 543134
rect 218062 542898 218146 543134
rect 218382 542898 253826 543134
rect 254062 542898 254146 543134
rect 254382 542898 289826 543134
rect 290062 542898 290146 543134
rect 290382 542898 325826 543134
rect 326062 542898 326146 543134
rect 326382 542898 361826 543134
rect 362062 542898 362146 543134
rect 362382 542898 397826 543134
rect 398062 542898 398146 543134
rect 398382 542898 433826 543134
rect 434062 542898 434146 543134
rect 434382 542898 469826 543134
rect 470062 542898 470146 543134
rect 470382 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 592650 543134
rect -8726 542866 592650 542898
rect -8726 538954 592650 538986
rect -8726 538718 -8694 538954
rect -8458 538718 -8374 538954
rect -8138 538718 33326 538954
rect 33562 538718 33646 538954
rect 33882 538718 69326 538954
rect 69562 538718 69646 538954
rect 69882 538718 105326 538954
rect 105562 538718 105646 538954
rect 105882 538718 141326 538954
rect 141562 538718 141646 538954
rect 141882 538718 177326 538954
rect 177562 538718 177646 538954
rect 177882 538718 213326 538954
rect 213562 538718 213646 538954
rect 213882 538718 249326 538954
rect 249562 538718 249646 538954
rect 249882 538718 285326 538954
rect 285562 538718 285646 538954
rect 285882 538718 321326 538954
rect 321562 538718 321646 538954
rect 321882 538718 357326 538954
rect 357562 538718 357646 538954
rect 357882 538718 393326 538954
rect 393562 538718 393646 538954
rect 393882 538718 429326 538954
rect 429562 538718 429646 538954
rect 429882 538718 465326 538954
rect 465562 538718 465646 538954
rect 465882 538718 501326 538954
rect 501562 538718 501646 538954
rect 501882 538718 537326 538954
rect 537562 538718 537646 538954
rect 537882 538718 573326 538954
rect 573562 538718 573646 538954
rect 573882 538718 592062 538954
rect 592298 538718 592382 538954
rect 592618 538718 592650 538954
rect -8726 538634 592650 538718
rect -8726 538398 -8694 538634
rect -8458 538398 -8374 538634
rect -8138 538398 33326 538634
rect 33562 538398 33646 538634
rect 33882 538398 69326 538634
rect 69562 538398 69646 538634
rect 69882 538398 105326 538634
rect 105562 538398 105646 538634
rect 105882 538398 141326 538634
rect 141562 538398 141646 538634
rect 141882 538398 177326 538634
rect 177562 538398 177646 538634
rect 177882 538398 213326 538634
rect 213562 538398 213646 538634
rect 213882 538398 249326 538634
rect 249562 538398 249646 538634
rect 249882 538398 285326 538634
rect 285562 538398 285646 538634
rect 285882 538398 321326 538634
rect 321562 538398 321646 538634
rect 321882 538398 357326 538634
rect 357562 538398 357646 538634
rect 357882 538398 393326 538634
rect 393562 538398 393646 538634
rect 393882 538398 429326 538634
rect 429562 538398 429646 538634
rect 429882 538398 465326 538634
rect 465562 538398 465646 538634
rect 465882 538398 501326 538634
rect 501562 538398 501646 538634
rect 501882 538398 537326 538634
rect 537562 538398 537646 538634
rect 537882 538398 573326 538634
rect 573562 538398 573646 538634
rect 573882 538398 592062 538634
rect 592298 538398 592382 538634
rect 592618 538398 592650 538634
rect -8726 538366 592650 538398
rect -8726 534454 592650 534486
rect -8726 534218 -7734 534454
rect -7498 534218 -7414 534454
rect -7178 534218 28826 534454
rect 29062 534218 29146 534454
rect 29382 534218 64826 534454
rect 65062 534218 65146 534454
rect 65382 534218 100826 534454
rect 101062 534218 101146 534454
rect 101382 534218 136826 534454
rect 137062 534218 137146 534454
rect 137382 534218 172826 534454
rect 173062 534218 173146 534454
rect 173382 534218 208826 534454
rect 209062 534218 209146 534454
rect 209382 534218 244826 534454
rect 245062 534218 245146 534454
rect 245382 534218 280826 534454
rect 281062 534218 281146 534454
rect 281382 534218 316826 534454
rect 317062 534218 317146 534454
rect 317382 534218 352826 534454
rect 353062 534218 353146 534454
rect 353382 534218 388826 534454
rect 389062 534218 389146 534454
rect 389382 534218 424826 534454
rect 425062 534218 425146 534454
rect 425382 534218 460826 534454
rect 461062 534218 461146 534454
rect 461382 534218 496826 534454
rect 497062 534218 497146 534454
rect 497382 534218 532826 534454
rect 533062 534218 533146 534454
rect 533382 534218 568826 534454
rect 569062 534218 569146 534454
rect 569382 534218 591102 534454
rect 591338 534218 591422 534454
rect 591658 534218 592650 534454
rect -8726 534134 592650 534218
rect -8726 533898 -7734 534134
rect -7498 533898 -7414 534134
rect -7178 533898 28826 534134
rect 29062 533898 29146 534134
rect 29382 533898 64826 534134
rect 65062 533898 65146 534134
rect 65382 533898 100826 534134
rect 101062 533898 101146 534134
rect 101382 533898 136826 534134
rect 137062 533898 137146 534134
rect 137382 533898 172826 534134
rect 173062 533898 173146 534134
rect 173382 533898 208826 534134
rect 209062 533898 209146 534134
rect 209382 533898 244826 534134
rect 245062 533898 245146 534134
rect 245382 533898 280826 534134
rect 281062 533898 281146 534134
rect 281382 533898 316826 534134
rect 317062 533898 317146 534134
rect 317382 533898 352826 534134
rect 353062 533898 353146 534134
rect 353382 533898 388826 534134
rect 389062 533898 389146 534134
rect 389382 533898 424826 534134
rect 425062 533898 425146 534134
rect 425382 533898 460826 534134
rect 461062 533898 461146 534134
rect 461382 533898 496826 534134
rect 497062 533898 497146 534134
rect 497382 533898 532826 534134
rect 533062 533898 533146 534134
rect 533382 533898 568826 534134
rect 569062 533898 569146 534134
rect 569382 533898 591102 534134
rect 591338 533898 591422 534134
rect 591658 533898 592650 534134
rect -8726 533866 592650 533898
rect -8726 529954 592650 529986
rect -8726 529718 -6774 529954
rect -6538 529718 -6454 529954
rect -6218 529718 24326 529954
rect 24562 529718 24646 529954
rect 24882 529718 60326 529954
rect 60562 529718 60646 529954
rect 60882 529718 96326 529954
rect 96562 529718 96646 529954
rect 96882 529718 132326 529954
rect 132562 529718 132646 529954
rect 132882 529718 168326 529954
rect 168562 529718 168646 529954
rect 168882 529718 204326 529954
rect 204562 529718 204646 529954
rect 204882 529718 240326 529954
rect 240562 529718 240646 529954
rect 240882 529718 276326 529954
rect 276562 529718 276646 529954
rect 276882 529718 312326 529954
rect 312562 529718 312646 529954
rect 312882 529718 348326 529954
rect 348562 529718 348646 529954
rect 348882 529718 384326 529954
rect 384562 529718 384646 529954
rect 384882 529718 420326 529954
rect 420562 529718 420646 529954
rect 420882 529718 456326 529954
rect 456562 529718 456646 529954
rect 456882 529718 492326 529954
rect 492562 529718 492646 529954
rect 492882 529718 528326 529954
rect 528562 529718 528646 529954
rect 528882 529718 564326 529954
rect 564562 529718 564646 529954
rect 564882 529718 590142 529954
rect 590378 529718 590462 529954
rect 590698 529718 592650 529954
rect -8726 529634 592650 529718
rect -8726 529398 -6774 529634
rect -6538 529398 -6454 529634
rect -6218 529398 24326 529634
rect 24562 529398 24646 529634
rect 24882 529398 60326 529634
rect 60562 529398 60646 529634
rect 60882 529398 96326 529634
rect 96562 529398 96646 529634
rect 96882 529398 132326 529634
rect 132562 529398 132646 529634
rect 132882 529398 168326 529634
rect 168562 529398 168646 529634
rect 168882 529398 204326 529634
rect 204562 529398 204646 529634
rect 204882 529398 240326 529634
rect 240562 529398 240646 529634
rect 240882 529398 276326 529634
rect 276562 529398 276646 529634
rect 276882 529398 312326 529634
rect 312562 529398 312646 529634
rect 312882 529398 348326 529634
rect 348562 529398 348646 529634
rect 348882 529398 384326 529634
rect 384562 529398 384646 529634
rect 384882 529398 420326 529634
rect 420562 529398 420646 529634
rect 420882 529398 456326 529634
rect 456562 529398 456646 529634
rect 456882 529398 492326 529634
rect 492562 529398 492646 529634
rect 492882 529398 528326 529634
rect 528562 529398 528646 529634
rect 528882 529398 564326 529634
rect 564562 529398 564646 529634
rect 564882 529398 590142 529634
rect 590378 529398 590462 529634
rect 590698 529398 592650 529634
rect -8726 529366 592650 529398
rect -8726 525454 592650 525486
rect -8726 525218 -5814 525454
rect -5578 525218 -5494 525454
rect -5258 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 55826 525454
rect 56062 525218 56146 525454
rect 56382 525218 91826 525454
rect 92062 525218 92146 525454
rect 92382 525218 127826 525454
rect 128062 525218 128146 525454
rect 128382 525218 163826 525454
rect 164062 525218 164146 525454
rect 164382 525218 199826 525454
rect 200062 525218 200146 525454
rect 200382 525218 235826 525454
rect 236062 525218 236146 525454
rect 236382 525218 271826 525454
rect 272062 525218 272146 525454
rect 272382 525218 307826 525454
rect 308062 525218 308146 525454
rect 308382 525218 343826 525454
rect 344062 525218 344146 525454
rect 344382 525218 379826 525454
rect 380062 525218 380146 525454
rect 380382 525218 415826 525454
rect 416062 525218 416146 525454
rect 416382 525218 451826 525454
rect 452062 525218 452146 525454
rect 452382 525218 487826 525454
rect 488062 525218 488146 525454
rect 488382 525218 523826 525454
rect 524062 525218 524146 525454
rect 524382 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 589182 525454
rect 589418 525218 589502 525454
rect 589738 525218 592650 525454
rect -8726 525134 592650 525218
rect -8726 524898 -5814 525134
rect -5578 524898 -5494 525134
rect -5258 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 55826 525134
rect 56062 524898 56146 525134
rect 56382 524898 91826 525134
rect 92062 524898 92146 525134
rect 92382 524898 127826 525134
rect 128062 524898 128146 525134
rect 128382 524898 163826 525134
rect 164062 524898 164146 525134
rect 164382 524898 199826 525134
rect 200062 524898 200146 525134
rect 200382 524898 235826 525134
rect 236062 524898 236146 525134
rect 236382 524898 271826 525134
rect 272062 524898 272146 525134
rect 272382 524898 307826 525134
rect 308062 524898 308146 525134
rect 308382 524898 343826 525134
rect 344062 524898 344146 525134
rect 344382 524898 379826 525134
rect 380062 524898 380146 525134
rect 380382 524898 415826 525134
rect 416062 524898 416146 525134
rect 416382 524898 451826 525134
rect 452062 524898 452146 525134
rect 452382 524898 487826 525134
rect 488062 524898 488146 525134
rect 488382 524898 523826 525134
rect 524062 524898 524146 525134
rect 524382 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 589182 525134
rect 589418 524898 589502 525134
rect 589738 524898 592650 525134
rect -8726 524866 592650 524898
rect -8726 520954 592650 520986
rect -8726 520718 -4854 520954
rect -4618 520718 -4534 520954
rect -4298 520718 15326 520954
rect 15562 520718 15646 520954
rect 15882 520718 51326 520954
rect 51562 520718 51646 520954
rect 51882 520718 87326 520954
rect 87562 520718 87646 520954
rect 87882 520718 123326 520954
rect 123562 520718 123646 520954
rect 123882 520718 159326 520954
rect 159562 520718 159646 520954
rect 159882 520718 195326 520954
rect 195562 520718 195646 520954
rect 195882 520718 231326 520954
rect 231562 520718 231646 520954
rect 231882 520718 267326 520954
rect 267562 520718 267646 520954
rect 267882 520718 303326 520954
rect 303562 520718 303646 520954
rect 303882 520718 339326 520954
rect 339562 520718 339646 520954
rect 339882 520718 375326 520954
rect 375562 520718 375646 520954
rect 375882 520718 411326 520954
rect 411562 520718 411646 520954
rect 411882 520718 447326 520954
rect 447562 520718 447646 520954
rect 447882 520718 483326 520954
rect 483562 520718 483646 520954
rect 483882 520718 519326 520954
rect 519562 520718 519646 520954
rect 519882 520718 555326 520954
rect 555562 520718 555646 520954
rect 555882 520718 588222 520954
rect 588458 520718 588542 520954
rect 588778 520718 592650 520954
rect -8726 520634 592650 520718
rect -8726 520398 -4854 520634
rect -4618 520398 -4534 520634
rect -4298 520398 15326 520634
rect 15562 520398 15646 520634
rect 15882 520398 51326 520634
rect 51562 520398 51646 520634
rect 51882 520398 87326 520634
rect 87562 520398 87646 520634
rect 87882 520398 123326 520634
rect 123562 520398 123646 520634
rect 123882 520398 159326 520634
rect 159562 520398 159646 520634
rect 159882 520398 195326 520634
rect 195562 520398 195646 520634
rect 195882 520398 231326 520634
rect 231562 520398 231646 520634
rect 231882 520398 267326 520634
rect 267562 520398 267646 520634
rect 267882 520398 303326 520634
rect 303562 520398 303646 520634
rect 303882 520398 339326 520634
rect 339562 520398 339646 520634
rect 339882 520398 375326 520634
rect 375562 520398 375646 520634
rect 375882 520398 411326 520634
rect 411562 520398 411646 520634
rect 411882 520398 447326 520634
rect 447562 520398 447646 520634
rect 447882 520398 483326 520634
rect 483562 520398 483646 520634
rect 483882 520398 519326 520634
rect 519562 520398 519646 520634
rect 519882 520398 555326 520634
rect 555562 520398 555646 520634
rect 555882 520398 588222 520634
rect 588458 520398 588542 520634
rect 588778 520398 592650 520634
rect -8726 520366 592650 520398
rect -8726 516454 592650 516486
rect -8726 516218 -3894 516454
rect -3658 516218 -3574 516454
rect -3338 516218 10826 516454
rect 11062 516218 11146 516454
rect 11382 516218 46826 516454
rect 47062 516218 47146 516454
rect 47382 516218 82826 516454
rect 83062 516218 83146 516454
rect 83382 516218 118826 516454
rect 119062 516218 119146 516454
rect 119382 516218 154826 516454
rect 155062 516218 155146 516454
rect 155382 516218 190826 516454
rect 191062 516218 191146 516454
rect 191382 516218 226826 516454
rect 227062 516218 227146 516454
rect 227382 516218 262826 516454
rect 263062 516218 263146 516454
rect 263382 516218 298826 516454
rect 299062 516218 299146 516454
rect 299382 516218 334826 516454
rect 335062 516218 335146 516454
rect 335382 516218 370826 516454
rect 371062 516218 371146 516454
rect 371382 516218 406826 516454
rect 407062 516218 407146 516454
rect 407382 516218 442826 516454
rect 443062 516218 443146 516454
rect 443382 516218 478826 516454
rect 479062 516218 479146 516454
rect 479382 516218 514826 516454
rect 515062 516218 515146 516454
rect 515382 516218 550826 516454
rect 551062 516218 551146 516454
rect 551382 516218 587262 516454
rect 587498 516218 587582 516454
rect 587818 516218 592650 516454
rect -8726 516134 592650 516218
rect -8726 515898 -3894 516134
rect -3658 515898 -3574 516134
rect -3338 515898 10826 516134
rect 11062 515898 11146 516134
rect 11382 515898 46826 516134
rect 47062 515898 47146 516134
rect 47382 515898 82826 516134
rect 83062 515898 83146 516134
rect 83382 515898 118826 516134
rect 119062 515898 119146 516134
rect 119382 515898 154826 516134
rect 155062 515898 155146 516134
rect 155382 515898 190826 516134
rect 191062 515898 191146 516134
rect 191382 515898 226826 516134
rect 227062 515898 227146 516134
rect 227382 515898 262826 516134
rect 263062 515898 263146 516134
rect 263382 515898 298826 516134
rect 299062 515898 299146 516134
rect 299382 515898 334826 516134
rect 335062 515898 335146 516134
rect 335382 515898 370826 516134
rect 371062 515898 371146 516134
rect 371382 515898 406826 516134
rect 407062 515898 407146 516134
rect 407382 515898 442826 516134
rect 443062 515898 443146 516134
rect 443382 515898 478826 516134
rect 479062 515898 479146 516134
rect 479382 515898 514826 516134
rect 515062 515898 515146 516134
rect 515382 515898 550826 516134
rect 551062 515898 551146 516134
rect 551382 515898 587262 516134
rect 587498 515898 587582 516134
rect 587818 515898 592650 516134
rect -8726 515866 592650 515898
rect -8726 511954 592650 511986
rect -8726 511718 -2934 511954
rect -2698 511718 -2614 511954
rect -2378 511718 6326 511954
rect 6562 511718 6646 511954
rect 6882 511718 42326 511954
rect 42562 511718 42646 511954
rect 42882 511718 78326 511954
rect 78562 511718 78646 511954
rect 78882 511718 114326 511954
rect 114562 511718 114646 511954
rect 114882 511718 150326 511954
rect 150562 511718 150646 511954
rect 150882 511718 186326 511954
rect 186562 511718 186646 511954
rect 186882 511718 222326 511954
rect 222562 511718 222646 511954
rect 222882 511718 258326 511954
rect 258562 511718 258646 511954
rect 258882 511718 294326 511954
rect 294562 511718 294646 511954
rect 294882 511718 330326 511954
rect 330562 511718 330646 511954
rect 330882 511718 366326 511954
rect 366562 511718 366646 511954
rect 366882 511718 402326 511954
rect 402562 511718 402646 511954
rect 402882 511718 438326 511954
rect 438562 511718 438646 511954
rect 438882 511718 474326 511954
rect 474562 511718 474646 511954
rect 474882 511718 510326 511954
rect 510562 511718 510646 511954
rect 510882 511718 546326 511954
rect 546562 511718 546646 511954
rect 546882 511718 582326 511954
rect 582562 511718 582646 511954
rect 582882 511718 586302 511954
rect 586538 511718 586622 511954
rect 586858 511718 592650 511954
rect -8726 511634 592650 511718
rect -8726 511398 -2934 511634
rect -2698 511398 -2614 511634
rect -2378 511398 6326 511634
rect 6562 511398 6646 511634
rect 6882 511398 42326 511634
rect 42562 511398 42646 511634
rect 42882 511398 78326 511634
rect 78562 511398 78646 511634
rect 78882 511398 114326 511634
rect 114562 511398 114646 511634
rect 114882 511398 150326 511634
rect 150562 511398 150646 511634
rect 150882 511398 186326 511634
rect 186562 511398 186646 511634
rect 186882 511398 222326 511634
rect 222562 511398 222646 511634
rect 222882 511398 258326 511634
rect 258562 511398 258646 511634
rect 258882 511398 294326 511634
rect 294562 511398 294646 511634
rect 294882 511398 330326 511634
rect 330562 511398 330646 511634
rect 330882 511398 366326 511634
rect 366562 511398 366646 511634
rect 366882 511398 402326 511634
rect 402562 511398 402646 511634
rect 402882 511398 438326 511634
rect 438562 511398 438646 511634
rect 438882 511398 474326 511634
rect 474562 511398 474646 511634
rect 474882 511398 510326 511634
rect 510562 511398 510646 511634
rect 510882 511398 546326 511634
rect 546562 511398 546646 511634
rect 546882 511398 582326 511634
rect 582562 511398 582646 511634
rect 582882 511398 586302 511634
rect 586538 511398 586622 511634
rect 586858 511398 592650 511634
rect -8726 511366 592650 511398
rect -8726 507454 592650 507486
rect -8726 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 73826 507454
rect 74062 507218 74146 507454
rect 74382 507218 109826 507454
rect 110062 507218 110146 507454
rect 110382 507218 145826 507454
rect 146062 507218 146146 507454
rect 146382 507218 181826 507454
rect 182062 507218 182146 507454
rect 182382 507218 217826 507454
rect 218062 507218 218146 507454
rect 218382 507218 253826 507454
rect 254062 507218 254146 507454
rect 254382 507218 289826 507454
rect 290062 507218 290146 507454
rect 290382 507218 325826 507454
rect 326062 507218 326146 507454
rect 326382 507218 361826 507454
rect 362062 507218 362146 507454
rect 362382 507218 397826 507454
rect 398062 507218 398146 507454
rect 398382 507218 433826 507454
rect 434062 507218 434146 507454
rect 434382 507218 469826 507454
rect 470062 507218 470146 507454
rect 470382 507218 505826 507454
rect 506062 507218 506146 507454
rect 506382 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 592650 507454
rect -8726 507134 592650 507218
rect -8726 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 73826 507134
rect 74062 506898 74146 507134
rect 74382 506898 109826 507134
rect 110062 506898 110146 507134
rect 110382 506898 145826 507134
rect 146062 506898 146146 507134
rect 146382 506898 181826 507134
rect 182062 506898 182146 507134
rect 182382 506898 217826 507134
rect 218062 506898 218146 507134
rect 218382 506898 253826 507134
rect 254062 506898 254146 507134
rect 254382 506898 289826 507134
rect 290062 506898 290146 507134
rect 290382 506898 325826 507134
rect 326062 506898 326146 507134
rect 326382 506898 361826 507134
rect 362062 506898 362146 507134
rect 362382 506898 397826 507134
rect 398062 506898 398146 507134
rect 398382 506898 433826 507134
rect 434062 506898 434146 507134
rect 434382 506898 469826 507134
rect 470062 506898 470146 507134
rect 470382 506898 505826 507134
rect 506062 506898 506146 507134
rect 506382 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 592650 507134
rect -8726 506866 592650 506898
rect -8726 502954 592650 502986
rect -8726 502718 -8694 502954
rect -8458 502718 -8374 502954
rect -8138 502718 33326 502954
rect 33562 502718 33646 502954
rect 33882 502718 69326 502954
rect 69562 502718 69646 502954
rect 69882 502718 105326 502954
rect 105562 502718 105646 502954
rect 105882 502718 141326 502954
rect 141562 502718 141646 502954
rect 141882 502718 177326 502954
rect 177562 502718 177646 502954
rect 177882 502718 213326 502954
rect 213562 502718 213646 502954
rect 213882 502718 249326 502954
rect 249562 502718 249646 502954
rect 249882 502718 285326 502954
rect 285562 502718 285646 502954
rect 285882 502718 321326 502954
rect 321562 502718 321646 502954
rect 321882 502718 357326 502954
rect 357562 502718 357646 502954
rect 357882 502718 393326 502954
rect 393562 502718 393646 502954
rect 393882 502718 429326 502954
rect 429562 502718 429646 502954
rect 429882 502718 465326 502954
rect 465562 502718 465646 502954
rect 465882 502718 501326 502954
rect 501562 502718 501646 502954
rect 501882 502718 537326 502954
rect 537562 502718 537646 502954
rect 537882 502718 573326 502954
rect 573562 502718 573646 502954
rect 573882 502718 592062 502954
rect 592298 502718 592382 502954
rect 592618 502718 592650 502954
rect -8726 502634 592650 502718
rect -8726 502398 -8694 502634
rect -8458 502398 -8374 502634
rect -8138 502398 33326 502634
rect 33562 502398 33646 502634
rect 33882 502398 69326 502634
rect 69562 502398 69646 502634
rect 69882 502398 105326 502634
rect 105562 502398 105646 502634
rect 105882 502398 141326 502634
rect 141562 502398 141646 502634
rect 141882 502398 177326 502634
rect 177562 502398 177646 502634
rect 177882 502398 213326 502634
rect 213562 502398 213646 502634
rect 213882 502398 249326 502634
rect 249562 502398 249646 502634
rect 249882 502398 285326 502634
rect 285562 502398 285646 502634
rect 285882 502398 321326 502634
rect 321562 502398 321646 502634
rect 321882 502398 357326 502634
rect 357562 502398 357646 502634
rect 357882 502398 393326 502634
rect 393562 502398 393646 502634
rect 393882 502398 429326 502634
rect 429562 502398 429646 502634
rect 429882 502398 465326 502634
rect 465562 502398 465646 502634
rect 465882 502398 501326 502634
rect 501562 502398 501646 502634
rect 501882 502398 537326 502634
rect 537562 502398 537646 502634
rect 537882 502398 573326 502634
rect 573562 502398 573646 502634
rect 573882 502398 592062 502634
rect 592298 502398 592382 502634
rect 592618 502398 592650 502634
rect -8726 502366 592650 502398
rect -8726 498454 592650 498486
rect -8726 498218 -7734 498454
rect -7498 498218 -7414 498454
rect -7178 498218 28826 498454
rect 29062 498218 29146 498454
rect 29382 498218 64826 498454
rect 65062 498218 65146 498454
rect 65382 498218 100826 498454
rect 101062 498218 101146 498454
rect 101382 498218 136826 498454
rect 137062 498218 137146 498454
rect 137382 498218 172826 498454
rect 173062 498218 173146 498454
rect 173382 498218 208826 498454
rect 209062 498218 209146 498454
rect 209382 498218 244826 498454
rect 245062 498218 245146 498454
rect 245382 498218 280826 498454
rect 281062 498218 281146 498454
rect 281382 498218 316826 498454
rect 317062 498218 317146 498454
rect 317382 498218 352826 498454
rect 353062 498218 353146 498454
rect 353382 498218 388826 498454
rect 389062 498218 389146 498454
rect 389382 498218 424826 498454
rect 425062 498218 425146 498454
rect 425382 498218 460826 498454
rect 461062 498218 461146 498454
rect 461382 498218 496826 498454
rect 497062 498218 497146 498454
rect 497382 498218 532826 498454
rect 533062 498218 533146 498454
rect 533382 498218 568826 498454
rect 569062 498218 569146 498454
rect 569382 498218 591102 498454
rect 591338 498218 591422 498454
rect 591658 498218 592650 498454
rect -8726 498134 592650 498218
rect -8726 497898 -7734 498134
rect -7498 497898 -7414 498134
rect -7178 497898 28826 498134
rect 29062 497898 29146 498134
rect 29382 497898 64826 498134
rect 65062 497898 65146 498134
rect 65382 497898 100826 498134
rect 101062 497898 101146 498134
rect 101382 497898 136826 498134
rect 137062 497898 137146 498134
rect 137382 497898 172826 498134
rect 173062 497898 173146 498134
rect 173382 497898 208826 498134
rect 209062 497898 209146 498134
rect 209382 497898 244826 498134
rect 245062 497898 245146 498134
rect 245382 497898 280826 498134
rect 281062 497898 281146 498134
rect 281382 497898 316826 498134
rect 317062 497898 317146 498134
rect 317382 497898 352826 498134
rect 353062 497898 353146 498134
rect 353382 497898 388826 498134
rect 389062 497898 389146 498134
rect 389382 497898 424826 498134
rect 425062 497898 425146 498134
rect 425382 497898 460826 498134
rect 461062 497898 461146 498134
rect 461382 497898 496826 498134
rect 497062 497898 497146 498134
rect 497382 497898 532826 498134
rect 533062 497898 533146 498134
rect 533382 497898 568826 498134
rect 569062 497898 569146 498134
rect 569382 497898 591102 498134
rect 591338 497898 591422 498134
rect 591658 497898 592650 498134
rect -8726 497866 592650 497898
rect -8726 493954 592650 493986
rect -8726 493718 -6774 493954
rect -6538 493718 -6454 493954
rect -6218 493718 24326 493954
rect 24562 493718 24646 493954
rect 24882 493718 60326 493954
rect 60562 493718 60646 493954
rect 60882 493718 96326 493954
rect 96562 493718 96646 493954
rect 96882 493718 132326 493954
rect 132562 493718 132646 493954
rect 132882 493718 168326 493954
rect 168562 493718 168646 493954
rect 168882 493718 204326 493954
rect 204562 493718 204646 493954
rect 204882 493718 240326 493954
rect 240562 493718 240646 493954
rect 240882 493718 276326 493954
rect 276562 493718 276646 493954
rect 276882 493718 312326 493954
rect 312562 493718 312646 493954
rect 312882 493718 348326 493954
rect 348562 493718 348646 493954
rect 348882 493718 384326 493954
rect 384562 493718 384646 493954
rect 384882 493718 420326 493954
rect 420562 493718 420646 493954
rect 420882 493718 456326 493954
rect 456562 493718 456646 493954
rect 456882 493718 492326 493954
rect 492562 493718 492646 493954
rect 492882 493718 528326 493954
rect 528562 493718 528646 493954
rect 528882 493718 564326 493954
rect 564562 493718 564646 493954
rect 564882 493718 590142 493954
rect 590378 493718 590462 493954
rect 590698 493718 592650 493954
rect -8726 493634 592650 493718
rect -8726 493398 -6774 493634
rect -6538 493398 -6454 493634
rect -6218 493398 24326 493634
rect 24562 493398 24646 493634
rect 24882 493398 60326 493634
rect 60562 493398 60646 493634
rect 60882 493398 96326 493634
rect 96562 493398 96646 493634
rect 96882 493398 132326 493634
rect 132562 493398 132646 493634
rect 132882 493398 168326 493634
rect 168562 493398 168646 493634
rect 168882 493398 204326 493634
rect 204562 493398 204646 493634
rect 204882 493398 240326 493634
rect 240562 493398 240646 493634
rect 240882 493398 276326 493634
rect 276562 493398 276646 493634
rect 276882 493398 312326 493634
rect 312562 493398 312646 493634
rect 312882 493398 348326 493634
rect 348562 493398 348646 493634
rect 348882 493398 384326 493634
rect 384562 493398 384646 493634
rect 384882 493398 420326 493634
rect 420562 493398 420646 493634
rect 420882 493398 456326 493634
rect 456562 493398 456646 493634
rect 456882 493398 492326 493634
rect 492562 493398 492646 493634
rect 492882 493398 528326 493634
rect 528562 493398 528646 493634
rect 528882 493398 564326 493634
rect 564562 493398 564646 493634
rect 564882 493398 590142 493634
rect 590378 493398 590462 493634
rect 590698 493398 592650 493634
rect -8726 493366 592650 493398
rect -8726 489454 592650 489486
rect -8726 489218 -5814 489454
rect -5578 489218 -5494 489454
rect -5258 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 55826 489454
rect 56062 489218 56146 489454
rect 56382 489218 91826 489454
rect 92062 489218 92146 489454
rect 92382 489218 127826 489454
rect 128062 489218 128146 489454
rect 128382 489218 163826 489454
rect 164062 489218 164146 489454
rect 164382 489218 199826 489454
rect 200062 489218 200146 489454
rect 200382 489218 235826 489454
rect 236062 489218 236146 489454
rect 236382 489218 271826 489454
rect 272062 489218 272146 489454
rect 272382 489218 307826 489454
rect 308062 489218 308146 489454
rect 308382 489218 343826 489454
rect 344062 489218 344146 489454
rect 344382 489218 379826 489454
rect 380062 489218 380146 489454
rect 380382 489218 415826 489454
rect 416062 489218 416146 489454
rect 416382 489218 451826 489454
rect 452062 489218 452146 489454
rect 452382 489218 487826 489454
rect 488062 489218 488146 489454
rect 488382 489218 523826 489454
rect 524062 489218 524146 489454
rect 524382 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 589182 489454
rect 589418 489218 589502 489454
rect 589738 489218 592650 489454
rect -8726 489134 592650 489218
rect -8726 488898 -5814 489134
rect -5578 488898 -5494 489134
rect -5258 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 55826 489134
rect 56062 488898 56146 489134
rect 56382 488898 91826 489134
rect 92062 488898 92146 489134
rect 92382 488898 127826 489134
rect 128062 488898 128146 489134
rect 128382 488898 163826 489134
rect 164062 488898 164146 489134
rect 164382 488898 199826 489134
rect 200062 488898 200146 489134
rect 200382 488898 235826 489134
rect 236062 488898 236146 489134
rect 236382 488898 271826 489134
rect 272062 488898 272146 489134
rect 272382 488898 307826 489134
rect 308062 488898 308146 489134
rect 308382 488898 343826 489134
rect 344062 488898 344146 489134
rect 344382 488898 379826 489134
rect 380062 488898 380146 489134
rect 380382 488898 415826 489134
rect 416062 488898 416146 489134
rect 416382 488898 451826 489134
rect 452062 488898 452146 489134
rect 452382 488898 487826 489134
rect 488062 488898 488146 489134
rect 488382 488898 523826 489134
rect 524062 488898 524146 489134
rect 524382 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 589182 489134
rect 589418 488898 589502 489134
rect 589738 488898 592650 489134
rect -8726 488866 592650 488898
rect -8726 484954 592650 484986
rect -8726 484718 -4854 484954
rect -4618 484718 -4534 484954
rect -4298 484718 15326 484954
rect 15562 484718 15646 484954
rect 15882 484718 51326 484954
rect 51562 484718 51646 484954
rect 51882 484718 87326 484954
rect 87562 484718 87646 484954
rect 87882 484718 123326 484954
rect 123562 484718 123646 484954
rect 123882 484718 159326 484954
rect 159562 484718 159646 484954
rect 159882 484718 195326 484954
rect 195562 484718 195646 484954
rect 195882 484718 231326 484954
rect 231562 484718 231646 484954
rect 231882 484718 267326 484954
rect 267562 484718 267646 484954
rect 267882 484718 303326 484954
rect 303562 484718 303646 484954
rect 303882 484718 339326 484954
rect 339562 484718 339646 484954
rect 339882 484718 375326 484954
rect 375562 484718 375646 484954
rect 375882 484718 411326 484954
rect 411562 484718 411646 484954
rect 411882 484718 447326 484954
rect 447562 484718 447646 484954
rect 447882 484718 483326 484954
rect 483562 484718 483646 484954
rect 483882 484718 519326 484954
rect 519562 484718 519646 484954
rect 519882 484718 555326 484954
rect 555562 484718 555646 484954
rect 555882 484718 588222 484954
rect 588458 484718 588542 484954
rect 588778 484718 592650 484954
rect -8726 484634 592650 484718
rect -8726 484398 -4854 484634
rect -4618 484398 -4534 484634
rect -4298 484398 15326 484634
rect 15562 484398 15646 484634
rect 15882 484398 51326 484634
rect 51562 484398 51646 484634
rect 51882 484398 87326 484634
rect 87562 484398 87646 484634
rect 87882 484398 123326 484634
rect 123562 484398 123646 484634
rect 123882 484398 159326 484634
rect 159562 484398 159646 484634
rect 159882 484398 195326 484634
rect 195562 484398 195646 484634
rect 195882 484398 231326 484634
rect 231562 484398 231646 484634
rect 231882 484398 267326 484634
rect 267562 484398 267646 484634
rect 267882 484398 303326 484634
rect 303562 484398 303646 484634
rect 303882 484398 339326 484634
rect 339562 484398 339646 484634
rect 339882 484398 375326 484634
rect 375562 484398 375646 484634
rect 375882 484398 411326 484634
rect 411562 484398 411646 484634
rect 411882 484398 447326 484634
rect 447562 484398 447646 484634
rect 447882 484398 483326 484634
rect 483562 484398 483646 484634
rect 483882 484398 519326 484634
rect 519562 484398 519646 484634
rect 519882 484398 555326 484634
rect 555562 484398 555646 484634
rect 555882 484398 588222 484634
rect 588458 484398 588542 484634
rect 588778 484398 592650 484634
rect -8726 484366 592650 484398
rect -8726 480454 592650 480486
rect -8726 480218 -3894 480454
rect -3658 480218 -3574 480454
rect -3338 480218 10826 480454
rect 11062 480218 11146 480454
rect 11382 480218 46826 480454
rect 47062 480218 47146 480454
rect 47382 480218 82826 480454
rect 83062 480218 83146 480454
rect 83382 480218 118826 480454
rect 119062 480218 119146 480454
rect 119382 480218 154826 480454
rect 155062 480218 155146 480454
rect 155382 480218 190826 480454
rect 191062 480218 191146 480454
rect 191382 480218 226826 480454
rect 227062 480218 227146 480454
rect 227382 480218 262826 480454
rect 263062 480218 263146 480454
rect 263382 480218 298826 480454
rect 299062 480218 299146 480454
rect 299382 480218 334826 480454
rect 335062 480218 335146 480454
rect 335382 480218 370826 480454
rect 371062 480218 371146 480454
rect 371382 480218 406826 480454
rect 407062 480218 407146 480454
rect 407382 480218 442826 480454
rect 443062 480218 443146 480454
rect 443382 480218 478826 480454
rect 479062 480218 479146 480454
rect 479382 480218 514826 480454
rect 515062 480218 515146 480454
rect 515382 480218 550826 480454
rect 551062 480218 551146 480454
rect 551382 480218 587262 480454
rect 587498 480218 587582 480454
rect 587818 480218 592650 480454
rect -8726 480134 592650 480218
rect -8726 479898 -3894 480134
rect -3658 479898 -3574 480134
rect -3338 479898 10826 480134
rect 11062 479898 11146 480134
rect 11382 479898 46826 480134
rect 47062 479898 47146 480134
rect 47382 479898 82826 480134
rect 83062 479898 83146 480134
rect 83382 479898 118826 480134
rect 119062 479898 119146 480134
rect 119382 479898 154826 480134
rect 155062 479898 155146 480134
rect 155382 479898 190826 480134
rect 191062 479898 191146 480134
rect 191382 479898 226826 480134
rect 227062 479898 227146 480134
rect 227382 479898 262826 480134
rect 263062 479898 263146 480134
rect 263382 479898 298826 480134
rect 299062 479898 299146 480134
rect 299382 479898 334826 480134
rect 335062 479898 335146 480134
rect 335382 479898 370826 480134
rect 371062 479898 371146 480134
rect 371382 479898 406826 480134
rect 407062 479898 407146 480134
rect 407382 479898 442826 480134
rect 443062 479898 443146 480134
rect 443382 479898 478826 480134
rect 479062 479898 479146 480134
rect 479382 479898 514826 480134
rect 515062 479898 515146 480134
rect 515382 479898 550826 480134
rect 551062 479898 551146 480134
rect 551382 479898 587262 480134
rect 587498 479898 587582 480134
rect 587818 479898 592650 480134
rect -8726 479866 592650 479898
rect -8726 475954 592650 475986
rect -8726 475718 -2934 475954
rect -2698 475718 -2614 475954
rect -2378 475718 6326 475954
rect 6562 475718 6646 475954
rect 6882 475718 42326 475954
rect 42562 475718 42646 475954
rect 42882 475718 78326 475954
rect 78562 475718 78646 475954
rect 78882 475718 114326 475954
rect 114562 475718 114646 475954
rect 114882 475718 150326 475954
rect 150562 475718 150646 475954
rect 150882 475718 186326 475954
rect 186562 475718 186646 475954
rect 186882 475718 222326 475954
rect 222562 475718 222646 475954
rect 222882 475718 258326 475954
rect 258562 475718 258646 475954
rect 258882 475718 294326 475954
rect 294562 475718 294646 475954
rect 294882 475718 330326 475954
rect 330562 475718 330646 475954
rect 330882 475718 366326 475954
rect 366562 475718 366646 475954
rect 366882 475718 402326 475954
rect 402562 475718 402646 475954
rect 402882 475718 438326 475954
rect 438562 475718 438646 475954
rect 438882 475718 474326 475954
rect 474562 475718 474646 475954
rect 474882 475718 510326 475954
rect 510562 475718 510646 475954
rect 510882 475718 546326 475954
rect 546562 475718 546646 475954
rect 546882 475718 582326 475954
rect 582562 475718 582646 475954
rect 582882 475718 586302 475954
rect 586538 475718 586622 475954
rect 586858 475718 592650 475954
rect -8726 475634 592650 475718
rect -8726 475398 -2934 475634
rect -2698 475398 -2614 475634
rect -2378 475398 6326 475634
rect 6562 475398 6646 475634
rect 6882 475398 42326 475634
rect 42562 475398 42646 475634
rect 42882 475398 78326 475634
rect 78562 475398 78646 475634
rect 78882 475398 114326 475634
rect 114562 475398 114646 475634
rect 114882 475398 150326 475634
rect 150562 475398 150646 475634
rect 150882 475398 186326 475634
rect 186562 475398 186646 475634
rect 186882 475398 222326 475634
rect 222562 475398 222646 475634
rect 222882 475398 258326 475634
rect 258562 475398 258646 475634
rect 258882 475398 294326 475634
rect 294562 475398 294646 475634
rect 294882 475398 330326 475634
rect 330562 475398 330646 475634
rect 330882 475398 366326 475634
rect 366562 475398 366646 475634
rect 366882 475398 402326 475634
rect 402562 475398 402646 475634
rect 402882 475398 438326 475634
rect 438562 475398 438646 475634
rect 438882 475398 474326 475634
rect 474562 475398 474646 475634
rect 474882 475398 510326 475634
rect 510562 475398 510646 475634
rect 510882 475398 546326 475634
rect 546562 475398 546646 475634
rect 546882 475398 582326 475634
rect 582562 475398 582646 475634
rect 582882 475398 586302 475634
rect 586538 475398 586622 475634
rect 586858 475398 592650 475634
rect -8726 475366 592650 475398
rect -8726 471454 592650 471486
rect -8726 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 73826 471454
rect 74062 471218 74146 471454
rect 74382 471218 109826 471454
rect 110062 471218 110146 471454
rect 110382 471218 145826 471454
rect 146062 471218 146146 471454
rect 146382 471218 181826 471454
rect 182062 471218 182146 471454
rect 182382 471218 217826 471454
rect 218062 471218 218146 471454
rect 218382 471218 253826 471454
rect 254062 471218 254146 471454
rect 254382 471218 289826 471454
rect 290062 471218 290146 471454
rect 290382 471218 325826 471454
rect 326062 471218 326146 471454
rect 326382 471218 361826 471454
rect 362062 471218 362146 471454
rect 362382 471218 397826 471454
rect 398062 471218 398146 471454
rect 398382 471218 433826 471454
rect 434062 471218 434146 471454
rect 434382 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 592650 471454
rect -8726 471134 592650 471218
rect -8726 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 73826 471134
rect 74062 470898 74146 471134
rect 74382 470898 109826 471134
rect 110062 470898 110146 471134
rect 110382 470898 145826 471134
rect 146062 470898 146146 471134
rect 146382 470898 181826 471134
rect 182062 470898 182146 471134
rect 182382 470898 217826 471134
rect 218062 470898 218146 471134
rect 218382 470898 253826 471134
rect 254062 470898 254146 471134
rect 254382 470898 289826 471134
rect 290062 470898 290146 471134
rect 290382 470898 325826 471134
rect 326062 470898 326146 471134
rect 326382 470898 361826 471134
rect 362062 470898 362146 471134
rect 362382 470898 397826 471134
rect 398062 470898 398146 471134
rect 398382 470898 433826 471134
rect 434062 470898 434146 471134
rect 434382 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 592650 471134
rect -8726 470866 592650 470898
rect -8726 466954 592650 466986
rect -8726 466718 -8694 466954
rect -8458 466718 -8374 466954
rect -8138 466718 33326 466954
rect 33562 466718 33646 466954
rect 33882 466718 69326 466954
rect 69562 466718 69646 466954
rect 69882 466718 105326 466954
rect 105562 466718 105646 466954
rect 105882 466718 141326 466954
rect 141562 466718 141646 466954
rect 141882 466718 177326 466954
rect 177562 466718 177646 466954
rect 177882 466718 213326 466954
rect 213562 466718 213646 466954
rect 213882 466718 249326 466954
rect 249562 466718 249646 466954
rect 249882 466718 285326 466954
rect 285562 466718 285646 466954
rect 285882 466718 321326 466954
rect 321562 466718 321646 466954
rect 321882 466718 357326 466954
rect 357562 466718 357646 466954
rect 357882 466718 393326 466954
rect 393562 466718 393646 466954
rect 393882 466718 429326 466954
rect 429562 466718 429646 466954
rect 429882 466718 465326 466954
rect 465562 466718 465646 466954
rect 465882 466718 501326 466954
rect 501562 466718 501646 466954
rect 501882 466718 537326 466954
rect 537562 466718 537646 466954
rect 537882 466718 573326 466954
rect 573562 466718 573646 466954
rect 573882 466718 592062 466954
rect 592298 466718 592382 466954
rect 592618 466718 592650 466954
rect -8726 466634 592650 466718
rect -8726 466398 -8694 466634
rect -8458 466398 -8374 466634
rect -8138 466398 33326 466634
rect 33562 466398 33646 466634
rect 33882 466398 69326 466634
rect 69562 466398 69646 466634
rect 69882 466398 105326 466634
rect 105562 466398 105646 466634
rect 105882 466398 141326 466634
rect 141562 466398 141646 466634
rect 141882 466398 177326 466634
rect 177562 466398 177646 466634
rect 177882 466398 213326 466634
rect 213562 466398 213646 466634
rect 213882 466398 249326 466634
rect 249562 466398 249646 466634
rect 249882 466398 285326 466634
rect 285562 466398 285646 466634
rect 285882 466398 321326 466634
rect 321562 466398 321646 466634
rect 321882 466398 357326 466634
rect 357562 466398 357646 466634
rect 357882 466398 393326 466634
rect 393562 466398 393646 466634
rect 393882 466398 429326 466634
rect 429562 466398 429646 466634
rect 429882 466398 465326 466634
rect 465562 466398 465646 466634
rect 465882 466398 501326 466634
rect 501562 466398 501646 466634
rect 501882 466398 537326 466634
rect 537562 466398 537646 466634
rect 537882 466398 573326 466634
rect 573562 466398 573646 466634
rect 573882 466398 592062 466634
rect 592298 466398 592382 466634
rect 592618 466398 592650 466634
rect -8726 466366 592650 466398
rect -8726 462454 592650 462486
rect -8726 462218 -7734 462454
rect -7498 462218 -7414 462454
rect -7178 462218 28826 462454
rect 29062 462218 29146 462454
rect 29382 462218 64826 462454
rect 65062 462218 65146 462454
rect 65382 462218 100826 462454
rect 101062 462218 101146 462454
rect 101382 462218 136826 462454
rect 137062 462218 137146 462454
rect 137382 462218 172826 462454
rect 173062 462218 173146 462454
rect 173382 462218 208826 462454
rect 209062 462218 209146 462454
rect 209382 462218 244826 462454
rect 245062 462218 245146 462454
rect 245382 462218 280826 462454
rect 281062 462218 281146 462454
rect 281382 462218 316826 462454
rect 317062 462218 317146 462454
rect 317382 462218 352826 462454
rect 353062 462218 353146 462454
rect 353382 462218 388826 462454
rect 389062 462218 389146 462454
rect 389382 462218 424826 462454
rect 425062 462218 425146 462454
rect 425382 462218 460826 462454
rect 461062 462218 461146 462454
rect 461382 462218 496826 462454
rect 497062 462218 497146 462454
rect 497382 462218 532826 462454
rect 533062 462218 533146 462454
rect 533382 462218 568826 462454
rect 569062 462218 569146 462454
rect 569382 462218 591102 462454
rect 591338 462218 591422 462454
rect 591658 462218 592650 462454
rect -8726 462134 592650 462218
rect -8726 461898 -7734 462134
rect -7498 461898 -7414 462134
rect -7178 461898 28826 462134
rect 29062 461898 29146 462134
rect 29382 461898 64826 462134
rect 65062 461898 65146 462134
rect 65382 461898 100826 462134
rect 101062 461898 101146 462134
rect 101382 461898 136826 462134
rect 137062 461898 137146 462134
rect 137382 461898 172826 462134
rect 173062 461898 173146 462134
rect 173382 461898 208826 462134
rect 209062 461898 209146 462134
rect 209382 461898 244826 462134
rect 245062 461898 245146 462134
rect 245382 461898 280826 462134
rect 281062 461898 281146 462134
rect 281382 461898 316826 462134
rect 317062 461898 317146 462134
rect 317382 461898 352826 462134
rect 353062 461898 353146 462134
rect 353382 461898 388826 462134
rect 389062 461898 389146 462134
rect 389382 461898 424826 462134
rect 425062 461898 425146 462134
rect 425382 461898 460826 462134
rect 461062 461898 461146 462134
rect 461382 461898 496826 462134
rect 497062 461898 497146 462134
rect 497382 461898 532826 462134
rect 533062 461898 533146 462134
rect 533382 461898 568826 462134
rect 569062 461898 569146 462134
rect 569382 461898 591102 462134
rect 591338 461898 591422 462134
rect 591658 461898 592650 462134
rect -8726 461866 592650 461898
rect -8726 457954 592650 457986
rect -8726 457718 -6774 457954
rect -6538 457718 -6454 457954
rect -6218 457718 24326 457954
rect 24562 457718 24646 457954
rect 24882 457718 60326 457954
rect 60562 457718 60646 457954
rect 60882 457718 96326 457954
rect 96562 457718 96646 457954
rect 96882 457718 132326 457954
rect 132562 457718 132646 457954
rect 132882 457718 168326 457954
rect 168562 457718 168646 457954
rect 168882 457718 204326 457954
rect 204562 457718 204646 457954
rect 204882 457718 240326 457954
rect 240562 457718 240646 457954
rect 240882 457718 276326 457954
rect 276562 457718 276646 457954
rect 276882 457718 312326 457954
rect 312562 457718 312646 457954
rect 312882 457718 348326 457954
rect 348562 457718 348646 457954
rect 348882 457718 384326 457954
rect 384562 457718 384646 457954
rect 384882 457718 420326 457954
rect 420562 457718 420646 457954
rect 420882 457718 456326 457954
rect 456562 457718 456646 457954
rect 456882 457718 492326 457954
rect 492562 457718 492646 457954
rect 492882 457718 528326 457954
rect 528562 457718 528646 457954
rect 528882 457718 564326 457954
rect 564562 457718 564646 457954
rect 564882 457718 590142 457954
rect 590378 457718 590462 457954
rect 590698 457718 592650 457954
rect -8726 457634 592650 457718
rect -8726 457398 -6774 457634
rect -6538 457398 -6454 457634
rect -6218 457398 24326 457634
rect 24562 457398 24646 457634
rect 24882 457398 60326 457634
rect 60562 457398 60646 457634
rect 60882 457398 96326 457634
rect 96562 457398 96646 457634
rect 96882 457398 132326 457634
rect 132562 457398 132646 457634
rect 132882 457398 168326 457634
rect 168562 457398 168646 457634
rect 168882 457398 204326 457634
rect 204562 457398 204646 457634
rect 204882 457398 240326 457634
rect 240562 457398 240646 457634
rect 240882 457398 276326 457634
rect 276562 457398 276646 457634
rect 276882 457398 312326 457634
rect 312562 457398 312646 457634
rect 312882 457398 348326 457634
rect 348562 457398 348646 457634
rect 348882 457398 384326 457634
rect 384562 457398 384646 457634
rect 384882 457398 420326 457634
rect 420562 457398 420646 457634
rect 420882 457398 456326 457634
rect 456562 457398 456646 457634
rect 456882 457398 492326 457634
rect 492562 457398 492646 457634
rect 492882 457398 528326 457634
rect 528562 457398 528646 457634
rect 528882 457398 564326 457634
rect 564562 457398 564646 457634
rect 564882 457398 590142 457634
rect 590378 457398 590462 457634
rect 590698 457398 592650 457634
rect -8726 457366 592650 457398
rect -8726 453454 592650 453486
rect -8726 453218 -5814 453454
rect -5578 453218 -5494 453454
rect -5258 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 55826 453454
rect 56062 453218 56146 453454
rect 56382 453218 91826 453454
rect 92062 453218 92146 453454
rect 92382 453218 127826 453454
rect 128062 453218 128146 453454
rect 128382 453218 163826 453454
rect 164062 453218 164146 453454
rect 164382 453218 199826 453454
rect 200062 453218 200146 453454
rect 200382 453218 235826 453454
rect 236062 453218 236146 453454
rect 236382 453218 271826 453454
rect 272062 453218 272146 453454
rect 272382 453218 307826 453454
rect 308062 453218 308146 453454
rect 308382 453218 343826 453454
rect 344062 453218 344146 453454
rect 344382 453218 379826 453454
rect 380062 453218 380146 453454
rect 380382 453218 415826 453454
rect 416062 453218 416146 453454
rect 416382 453218 451826 453454
rect 452062 453218 452146 453454
rect 452382 453218 487826 453454
rect 488062 453218 488146 453454
rect 488382 453218 523826 453454
rect 524062 453218 524146 453454
rect 524382 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 589182 453454
rect 589418 453218 589502 453454
rect 589738 453218 592650 453454
rect -8726 453134 592650 453218
rect -8726 452898 -5814 453134
rect -5578 452898 -5494 453134
rect -5258 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 55826 453134
rect 56062 452898 56146 453134
rect 56382 452898 91826 453134
rect 92062 452898 92146 453134
rect 92382 452898 127826 453134
rect 128062 452898 128146 453134
rect 128382 452898 163826 453134
rect 164062 452898 164146 453134
rect 164382 452898 199826 453134
rect 200062 452898 200146 453134
rect 200382 452898 235826 453134
rect 236062 452898 236146 453134
rect 236382 452898 271826 453134
rect 272062 452898 272146 453134
rect 272382 452898 307826 453134
rect 308062 452898 308146 453134
rect 308382 452898 343826 453134
rect 344062 452898 344146 453134
rect 344382 452898 379826 453134
rect 380062 452898 380146 453134
rect 380382 452898 415826 453134
rect 416062 452898 416146 453134
rect 416382 452898 451826 453134
rect 452062 452898 452146 453134
rect 452382 452898 487826 453134
rect 488062 452898 488146 453134
rect 488382 452898 523826 453134
rect 524062 452898 524146 453134
rect 524382 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 589182 453134
rect 589418 452898 589502 453134
rect 589738 452898 592650 453134
rect -8726 452866 592650 452898
rect -8726 448954 592650 448986
rect -8726 448718 -4854 448954
rect -4618 448718 -4534 448954
rect -4298 448718 15326 448954
rect 15562 448718 15646 448954
rect 15882 448718 51326 448954
rect 51562 448718 51646 448954
rect 51882 448718 87326 448954
rect 87562 448718 87646 448954
rect 87882 448718 123326 448954
rect 123562 448718 123646 448954
rect 123882 448718 159326 448954
rect 159562 448718 159646 448954
rect 159882 448718 195326 448954
rect 195562 448718 195646 448954
rect 195882 448718 231326 448954
rect 231562 448718 231646 448954
rect 231882 448718 267326 448954
rect 267562 448718 267646 448954
rect 267882 448718 303326 448954
rect 303562 448718 303646 448954
rect 303882 448718 339326 448954
rect 339562 448718 339646 448954
rect 339882 448718 375326 448954
rect 375562 448718 375646 448954
rect 375882 448718 411326 448954
rect 411562 448718 411646 448954
rect 411882 448718 447326 448954
rect 447562 448718 447646 448954
rect 447882 448718 483326 448954
rect 483562 448718 483646 448954
rect 483882 448718 519326 448954
rect 519562 448718 519646 448954
rect 519882 448718 555326 448954
rect 555562 448718 555646 448954
rect 555882 448718 588222 448954
rect 588458 448718 588542 448954
rect 588778 448718 592650 448954
rect -8726 448634 592650 448718
rect -8726 448398 -4854 448634
rect -4618 448398 -4534 448634
rect -4298 448398 15326 448634
rect 15562 448398 15646 448634
rect 15882 448398 51326 448634
rect 51562 448398 51646 448634
rect 51882 448398 87326 448634
rect 87562 448398 87646 448634
rect 87882 448398 123326 448634
rect 123562 448398 123646 448634
rect 123882 448398 159326 448634
rect 159562 448398 159646 448634
rect 159882 448398 195326 448634
rect 195562 448398 195646 448634
rect 195882 448398 231326 448634
rect 231562 448398 231646 448634
rect 231882 448398 267326 448634
rect 267562 448398 267646 448634
rect 267882 448398 303326 448634
rect 303562 448398 303646 448634
rect 303882 448398 339326 448634
rect 339562 448398 339646 448634
rect 339882 448398 375326 448634
rect 375562 448398 375646 448634
rect 375882 448398 411326 448634
rect 411562 448398 411646 448634
rect 411882 448398 447326 448634
rect 447562 448398 447646 448634
rect 447882 448398 483326 448634
rect 483562 448398 483646 448634
rect 483882 448398 519326 448634
rect 519562 448398 519646 448634
rect 519882 448398 555326 448634
rect 555562 448398 555646 448634
rect 555882 448398 588222 448634
rect 588458 448398 588542 448634
rect 588778 448398 592650 448634
rect -8726 448366 592650 448398
rect -8726 444454 592650 444486
rect -8726 444218 -3894 444454
rect -3658 444218 -3574 444454
rect -3338 444218 10826 444454
rect 11062 444218 11146 444454
rect 11382 444218 46826 444454
rect 47062 444218 47146 444454
rect 47382 444218 82826 444454
rect 83062 444218 83146 444454
rect 83382 444218 118826 444454
rect 119062 444218 119146 444454
rect 119382 444218 154826 444454
rect 155062 444218 155146 444454
rect 155382 444218 190826 444454
rect 191062 444218 191146 444454
rect 191382 444218 226826 444454
rect 227062 444218 227146 444454
rect 227382 444218 262826 444454
rect 263062 444218 263146 444454
rect 263382 444218 298826 444454
rect 299062 444218 299146 444454
rect 299382 444218 334826 444454
rect 335062 444218 335146 444454
rect 335382 444218 370826 444454
rect 371062 444218 371146 444454
rect 371382 444218 406826 444454
rect 407062 444218 407146 444454
rect 407382 444218 442826 444454
rect 443062 444218 443146 444454
rect 443382 444218 478826 444454
rect 479062 444218 479146 444454
rect 479382 444218 514826 444454
rect 515062 444218 515146 444454
rect 515382 444218 550826 444454
rect 551062 444218 551146 444454
rect 551382 444218 587262 444454
rect 587498 444218 587582 444454
rect 587818 444218 592650 444454
rect -8726 444134 592650 444218
rect -8726 443898 -3894 444134
rect -3658 443898 -3574 444134
rect -3338 443898 10826 444134
rect 11062 443898 11146 444134
rect 11382 443898 46826 444134
rect 47062 443898 47146 444134
rect 47382 443898 82826 444134
rect 83062 443898 83146 444134
rect 83382 443898 118826 444134
rect 119062 443898 119146 444134
rect 119382 443898 154826 444134
rect 155062 443898 155146 444134
rect 155382 443898 190826 444134
rect 191062 443898 191146 444134
rect 191382 443898 226826 444134
rect 227062 443898 227146 444134
rect 227382 443898 262826 444134
rect 263062 443898 263146 444134
rect 263382 443898 298826 444134
rect 299062 443898 299146 444134
rect 299382 443898 334826 444134
rect 335062 443898 335146 444134
rect 335382 443898 370826 444134
rect 371062 443898 371146 444134
rect 371382 443898 406826 444134
rect 407062 443898 407146 444134
rect 407382 443898 442826 444134
rect 443062 443898 443146 444134
rect 443382 443898 478826 444134
rect 479062 443898 479146 444134
rect 479382 443898 514826 444134
rect 515062 443898 515146 444134
rect 515382 443898 550826 444134
rect 551062 443898 551146 444134
rect 551382 443898 587262 444134
rect 587498 443898 587582 444134
rect 587818 443898 592650 444134
rect -8726 443866 592650 443898
rect -8726 439954 592650 439986
rect -8726 439718 -2934 439954
rect -2698 439718 -2614 439954
rect -2378 439718 6326 439954
rect 6562 439718 6646 439954
rect 6882 439718 42326 439954
rect 42562 439718 42646 439954
rect 42882 439718 78326 439954
rect 78562 439718 78646 439954
rect 78882 439718 114326 439954
rect 114562 439718 114646 439954
rect 114882 439718 150326 439954
rect 150562 439718 150646 439954
rect 150882 439718 186326 439954
rect 186562 439718 186646 439954
rect 186882 439718 222326 439954
rect 222562 439718 222646 439954
rect 222882 439718 258326 439954
rect 258562 439718 258646 439954
rect 258882 439718 294326 439954
rect 294562 439718 294646 439954
rect 294882 439718 330326 439954
rect 330562 439718 330646 439954
rect 330882 439718 366326 439954
rect 366562 439718 366646 439954
rect 366882 439718 402326 439954
rect 402562 439718 402646 439954
rect 402882 439718 438326 439954
rect 438562 439718 438646 439954
rect 438882 439718 474326 439954
rect 474562 439718 474646 439954
rect 474882 439718 510326 439954
rect 510562 439718 510646 439954
rect 510882 439718 546326 439954
rect 546562 439718 546646 439954
rect 546882 439718 582326 439954
rect 582562 439718 582646 439954
rect 582882 439718 586302 439954
rect 586538 439718 586622 439954
rect 586858 439718 592650 439954
rect -8726 439634 592650 439718
rect -8726 439398 -2934 439634
rect -2698 439398 -2614 439634
rect -2378 439398 6326 439634
rect 6562 439398 6646 439634
rect 6882 439398 42326 439634
rect 42562 439398 42646 439634
rect 42882 439398 78326 439634
rect 78562 439398 78646 439634
rect 78882 439398 114326 439634
rect 114562 439398 114646 439634
rect 114882 439398 150326 439634
rect 150562 439398 150646 439634
rect 150882 439398 186326 439634
rect 186562 439398 186646 439634
rect 186882 439398 222326 439634
rect 222562 439398 222646 439634
rect 222882 439398 258326 439634
rect 258562 439398 258646 439634
rect 258882 439398 294326 439634
rect 294562 439398 294646 439634
rect 294882 439398 330326 439634
rect 330562 439398 330646 439634
rect 330882 439398 366326 439634
rect 366562 439398 366646 439634
rect 366882 439398 402326 439634
rect 402562 439398 402646 439634
rect 402882 439398 438326 439634
rect 438562 439398 438646 439634
rect 438882 439398 474326 439634
rect 474562 439398 474646 439634
rect 474882 439398 510326 439634
rect 510562 439398 510646 439634
rect 510882 439398 546326 439634
rect 546562 439398 546646 439634
rect 546882 439398 582326 439634
rect 582562 439398 582646 439634
rect 582882 439398 586302 439634
rect 586538 439398 586622 439634
rect 586858 439398 592650 439634
rect -8726 439366 592650 439398
rect -8726 435454 592650 435486
rect -8726 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 73826 435454
rect 74062 435218 74146 435454
rect 74382 435218 109826 435454
rect 110062 435218 110146 435454
rect 110382 435218 145826 435454
rect 146062 435218 146146 435454
rect 146382 435218 181826 435454
rect 182062 435218 182146 435454
rect 182382 435218 217826 435454
rect 218062 435218 218146 435454
rect 218382 435218 253826 435454
rect 254062 435218 254146 435454
rect 254382 435218 289826 435454
rect 290062 435218 290146 435454
rect 290382 435218 325826 435454
rect 326062 435218 326146 435454
rect 326382 435218 361826 435454
rect 362062 435218 362146 435454
rect 362382 435218 397826 435454
rect 398062 435218 398146 435454
rect 398382 435218 433826 435454
rect 434062 435218 434146 435454
rect 434382 435218 469826 435454
rect 470062 435218 470146 435454
rect 470382 435218 505826 435454
rect 506062 435218 506146 435454
rect 506382 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 592650 435454
rect -8726 435134 592650 435218
rect -8726 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 73826 435134
rect 74062 434898 74146 435134
rect 74382 434898 109826 435134
rect 110062 434898 110146 435134
rect 110382 434898 145826 435134
rect 146062 434898 146146 435134
rect 146382 434898 181826 435134
rect 182062 434898 182146 435134
rect 182382 434898 217826 435134
rect 218062 434898 218146 435134
rect 218382 434898 253826 435134
rect 254062 434898 254146 435134
rect 254382 434898 289826 435134
rect 290062 434898 290146 435134
rect 290382 434898 325826 435134
rect 326062 434898 326146 435134
rect 326382 434898 361826 435134
rect 362062 434898 362146 435134
rect 362382 434898 397826 435134
rect 398062 434898 398146 435134
rect 398382 434898 433826 435134
rect 434062 434898 434146 435134
rect 434382 434898 469826 435134
rect 470062 434898 470146 435134
rect 470382 434898 505826 435134
rect 506062 434898 506146 435134
rect 506382 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 592650 435134
rect -8726 434866 592650 434898
rect -8726 430954 592650 430986
rect -8726 430718 -8694 430954
rect -8458 430718 -8374 430954
rect -8138 430718 33326 430954
rect 33562 430718 33646 430954
rect 33882 430718 69326 430954
rect 69562 430718 69646 430954
rect 69882 430718 105326 430954
rect 105562 430718 105646 430954
rect 105882 430718 141326 430954
rect 141562 430718 141646 430954
rect 141882 430718 177326 430954
rect 177562 430718 177646 430954
rect 177882 430718 213326 430954
rect 213562 430718 213646 430954
rect 213882 430718 249326 430954
rect 249562 430718 249646 430954
rect 249882 430718 285326 430954
rect 285562 430718 285646 430954
rect 285882 430718 321326 430954
rect 321562 430718 321646 430954
rect 321882 430718 357326 430954
rect 357562 430718 357646 430954
rect 357882 430718 393326 430954
rect 393562 430718 393646 430954
rect 393882 430718 429326 430954
rect 429562 430718 429646 430954
rect 429882 430718 465326 430954
rect 465562 430718 465646 430954
rect 465882 430718 501326 430954
rect 501562 430718 501646 430954
rect 501882 430718 537326 430954
rect 537562 430718 537646 430954
rect 537882 430718 573326 430954
rect 573562 430718 573646 430954
rect 573882 430718 592062 430954
rect 592298 430718 592382 430954
rect 592618 430718 592650 430954
rect -8726 430634 592650 430718
rect -8726 430398 -8694 430634
rect -8458 430398 -8374 430634
rect -8138 430398 33326 430634
rect 33562 430398 33646 430634
rect 33882 430398 69326 430634
rect 69562 430398 69646 430634
rect 69882 430398 105326 430634
rect 105562 430398 105646 430634
rect 105882 430398 141326 430634
rect 141562 430398 141646 430634
rect 141882 430398 177326 430634
rect 177562 430398 177646 430634
rect 177882 430398 213326 430634
rect 213562 430398 213646 430634
rect 213882 430398 249326 430634
rect 249562 430398 249646 430634
rect 249882 430398 285326 430634
rect 285562 430398 285646 430634
rect 285882 430398 321326 430634
rect 321562 430398 321646 430634
rect 321882 430398 357326 430634
rect 357562 430398 357646 430634
rect 357882 430398 393326 430634
rect 393562 430398 393646 430634
rect 393882 430398 429326 430634
rect 429562 430398 429646 430634
rect 429882 430398 465326 430634
rect 465562 430398 465646 430634
rect 465882 430398 501326 430634
rect 501562 430398 501646 430634
rect 501882 430398 537326 430634
rect 537562 430398 537646 430634
rect 537882 430398 573326 430634
rect 573562 430398 573646 430634
rect 573882 430398 592062 430634
rect 592298 430398 592382 430634
rect 592618 430398 592650 430634
rect -8726 430366 592650 430398
rect -8726 426454 592650 426486
rect -8726 426218 -7734 426454
rect -7498 426218 -7414 426454
rect -7178 426218 28826 426454
rect 29062 426218 29146 426454
rect 29382 426218 64826 426454
rect 65062 426218 65146 426454
rect 65382 426218 100826 426454
rect 101062 426218 101146 426454
rect 101382 426218 136826 426454
rect 137062 426218 137146 426454
rect 137382 426218 172826 426454
rect 173062 426218 173146 426454
rect 173382 426218 208826 426454
rect 209062 426218 209146 426454
rect 209382 426218 244826 426454
rect 245062 426218 245146 426454
rect 245382 426218 280826 426454
rect 281062 426218 281146 426454
rect 281382 426218 316826 426454
rect 317062 426218 317146 426454
rect 317382 426218 352826 426454
rect 353062 426218 353146 426454
rect 353382 426218 388826 426454
rect 389062 426218 389146 426454
rect 389382 426218 424826 426454
rect 425062 426218 425146 426454
rect 425382 426218 460826 426454
rect 461062 426218 461146 426454
rect 461382 426218 496826 426454
rect 497062 426218 497146 426454
rect 497382 426218 532826 426454
rect 533062 426218 533146 426454
rect 533382 426218 568826 426454
rect 569062 426218 569146 426454
rect 569382 426218 591102 426454
rect 591338 426218 591422 426454
rect 591658 426218 592650 426454
rect -8726 426134 592650 426218
rect -8726 425898 -7734 426134
rect -7498 425898 -7414 426134
rect -7178 425898 28826 426134
rect 29062 425898 29146 426134
rect 29382 425898 64826 426134
rect 65062 425898 65146 426134
rect 65382 425898 100826 426134
rect 101062 425898 101146 426134
rect 101382 425898 136826 426134
rect 137062 425898 137146 426134
rect 137382 425898 172826 426134
rect 173062 425898 173146 426134
rect 173382 425898 208826 426134
rect 209062 425898 209146 426134
rect 209382 425898 244826 426134
rect 245062 425898 245146 426134
rect 245382 425898 280826 426134
rect 281062 425898 281146 426134
rect 281382 425898 316826 426134
rect 317062 425898 317146 426134
rect 317382 425898 352826 426134
rect 353062 425898 353146 426134
rect 353382 425898 388826 426134
rect 389062 425898 389146 426134
rect 389382 425898 424826 426134
rect 425062 425898 425146 426134
rect 425382 425898 460826 426134
rect 461062 425898 461146 426134
rect 461382 425898 496826 426134
rect 497062 425898 497146 426134
rect 497382 425898 532826 426134
rect 533062 425898 533146 426134
rect 533382 425898 568826 426134
rect 569062 425898 569146 426134
rect 569382 425898 591102 426134
rect 591338 425898 591422 426134
rect 591658 425898 592650 426134
rect -8726 425866 592650 425898
rect -8726 421954 592650 421986
rect -8726 421718 -6774 421954
rect -6538 421718 -6454 421954
rect -6218 421718 24326 421954
rect 24562 421718 24646 421954
rect 24882 421718 60326 421954
rect 60562 421718 60646 421954
rect 60882 421718 96326 421954
rect 96562 421718 96646 421954
rect 96882 421718 132326 421954
rect 132562 421718 132646 421954
rect 132882 421718 168326 421954
rect 168562 421718 168646 421954
rect 168882 421718 204326 421954
rect 204562 421718 204646 421954
rect 204882 421718 240326 421954
rect 240562 421718 240646 421954
rect 240882 421718 276326 421954
rect 276562 421718 276646 421954
rect 276882 421718 312326 421954
rect 312562 421718 312646 421954
rect 312882 421718 348326 421954
rect 348562 421718 348646 421954
rect 348882 421718 384326 421954
rect 384562 421718 384646 421954
rect 384882 421718 420326 421954
rect 420562 421718 420646 421954
rect 420882 421718 456326 421954
rect 456562 421718 456646 421954
rect 456882 421718 492326 421954
rect 492562 421718 492646 421954
rect 492882 421718 528326 421954
rect 528562 421718 528646 421954
rect 528882 421718 564326 421954
rect 564562 421718 564646 421954
rect 564882 421718 590142 421954
rect 590378 421718 590462 421954
rect 590698 421718 592650 421954
rect -8726 421634 592650 421718
rect -8726 421398 -6774 421634
rect -6538 421398 -6454 421634
rect -6218 421398 24326 421634
rect 24562 421398 24646 421634
rect 24882 421398 60326 421634
rect 60562 421398 60646 421634
rect 60882 421398 96326 421634
rect 96562 421398 96646 421634
rect 96882 421398 132326 421634
rect 132562 421398 132646 421634
rect 132882 421398 168326 421634
rect 168562 421398 168646 421634
rect 168882 421398 204326 421634
rect 204562 421398 204646 421634
rect 204882 421398 240326 421634
rect 240562 421398 240646 421634
rect 240882 421398 276326 421634
rect 276562 421398 276646 421634
rect 276882 421398 312326 421634
rect 312562 421398 312646 421634
rect 312882 421398 348326 421634
rect 348562 421398 348646 421634
rect 348882 421398 384326 421634
rect 384562 421398 384646 421634
rect 384882 421398 420326 421634
rect 420562 421398 420646 421634
rect 420882 421398 456326 421634
rect 456562 421398 456646 421634
rect 456882 421398 492326 421634
rect 492562 421398 492646 421634
rect 492882 421398 528326 421634
rect 528562 421398 528646 421634
rect 528882 421398 564326 421634
rect 564562 421398 564646 421634
rect 564882 421398 590142 421634
rect 590378 421398 590462 421634
rect 590698 421398 592650 421634
rect -8726 421366 592650 421398
rect -8726 417454 592650 417486
rect -8726 417218 -5814 417454
rect -5578 417218 -5494 417454
rect -5258 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 55826 417454
rect 56062 417218 56146 417454
rect 56382 417218 91826 417454
rect 92062 417218 92146 417454
rect 92382 417218 127826 417454
rect 128062 417218 128146 417454
rect 128382 417218 163826 417454
rect 164062 417218 164146 417454
rect 164382 417218 199826 417454
rect 200062 417218 200146 417454
rect 200382 417218 235826 417454
rect 236062 417218 236146 417454
rect 236382 417218 271826 417454
rect 272062 417218 272146 417454
rect 272382 417218 307826 417454
rect 308062 417218 308146 417454
rect 308382 417218 343826 417454
rect 344062 417218 344146 417454
rect 344382 417218 379826 417454
rect 380062 417218 380146 417454
rect 380382 417218 415826 417454
rect 416062 417218 416146 417454
rect 416382 417218 451826 417454
rect 452062 417218 452146 417454
rect 452382 417218 487826 417454
rect 488062 417218 488146 417454
rect 488382 417218 523826 417454
rect 524062 417218 524146 417454
rect 524382 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 589182 417454
rect 589418 417218 589502 417454
rect 589738 417218 592650 417454
rect -8726 417134 592650 417218
rect -8726 416898 -5814 417134
rect -5578 416898 -5494 417134
rect -5258 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 55826 417134
rect 56062 416898 56146 417134
rect 56382 416898 91826 417134
rect 92062 416898 92146 417134
rect 92382 416898 127826 417134
rect 128062 416898 128146 417134
rect 128382 416898 163826 417134
rect 164062 416898 164146 417134
rect 164382 416898 199826 417134
rect 200062 416898 200146 417134
rect 200382 416898 235826 417134
rect 236062 416898 236146 417134
rect 236382 416898 271826 417134
rect 272062 416898 272146 417134
rect 272382 416898 307826 417134
rect 308062 416898 308146 417134
rect 308382 416898 343826 417134
rect 344062 416898 344146 417134
rect 344382 416898 379826 417134
rect 380062 416898 380146 417134
rect 380382 416898 415826 417134
rect 416062 416898 416146 417134
rect 416382 416898 451826 417134
rect 452062 416898 452146 417134
rect 452382 416898 487826 417134
rect 488062 416898 488146 417134
rect 488382 416898 523826 417134
rect 524062 416898 524146 417134
rect 524382 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 589182 417134
rect 589418 416898 589502 417134
rect 589738 416898 592650 417134
rect -8726 416866 592650 416898
rect -8726 412954 592650 412986
rect -8726 412718 -4854 412954
rect -4618 412718 -4534 412954
rect -4298 412718 15326 412954
rect 15562 412718 15646 412954
rect 15882 412718 51326 412954
rect 51562 412718 51646 412954
rect 51882 412718 87326 412954
rect 87562 412718 87646 412954
rect 87882 412718 123326 412954
rect 123562 412718 123646 412954
rect 123882 412718 159326 412954
rect 159562 412718 159646 412954
rect 159882 412718 195326 412954
rect 195562 412718 195646 412954
rect 195882 412718 231326 412954
rect 231562 412718 231646 412954
rect 231882 412718 267326 412954
rect 267562 412718 267646 412954
rect 267882 412718 303326 412954
rect 303562 412718 303646 412954
rect 303882 412718 339326 412954
rect 339562 412718 339646 412954
rect 339882 412718 375326 412954
rect 375562 412718 375646 412954
rect 375882 412718 411326 412954
rect 411562 412718 411646 412954
rect 411882 412718 447326 412954
rect 447562 412718 447646 412954
rect 447882 412718 483326 412954
rect 483562 412718 483646 412954
rect 483882 412718 519326 412954
rect 519562 412718 519646 412954
rect 519882 412718 555326 412954
rect 555562 412718 555646 412954
rect 555882 412718 588222 412954
rect 588458 412718 588542 412954
rect 588778 412718 592650 412954
rect -8726 412634 592650 412718
rect -8726 412398 -4854 412634
rect -4618 412398 -4534 412634
rect -4298 412398 15326 412634
rect 15562 412398 15646 412634
rect 15882 412398 51326 412634
rect 51562 412398 51646 412634
rect 51882 412398 87326 412634
rect 87562 412398 87646 412634
rect 87882 412398 123326 412634
rect 123562 412398 123646 412634
rect 123882 412398 159326 412634
rect 159562 412398 159646 412634
rect 159882 412398 195326 412634
rect 195562 412398 195646 412634
rect 195882 412398 231326 412634
rect 231562 412398 231646 412634
rect 231882 412398 267326 412634
rect 267562 412398 267646 412634
rect 267882 412398 303326 412634
rect 303562 412398 303646 412634
rect 303882 412398 339326 412634
rect 339562 412398 339646 412634
rect 339882 412398 375326 412634
rect 375562 412398 375646 412634
rect 375882 412398 411326 412634
rect 411562 412398 411646 412634
rect 411882 412398 447326 412634
rect 447562 412398 447646 412634
rect 447882 412398 483326 412634
rect 483562 412398 483646 412634
rect 483882 412398 519326 412634
rect 519562 412398 519646 412634
rect 519882 412398 555326 412634
rect 555562 412398 555646 412634
rect 555882 412398 588222 412634
rect 588458 412398 588542 412634
rect 588778 412398 592650 412634
rect -8726 412366 592650 412398
rect -8726 408454 592650 408486
rect -8726 408218 -3894 408454
rect -3658 408218 -3574 408454
rect -3338 408218 10826 408454
rect 11062 408218 11146 408454
rect 11382 408218 46826 408454
rect 47062 408218 47146 408454
rect 47382 408218 82826 408454
rect 83062 408218 83146 408454
rect 83382 408218 118826 408454
rect 119062 408218 119146 408454
rect 119382 408218 154826 408454
rect 155062 408218 155146 408454
rect 155382 408218 190826 408454
rect 191062 408218 191146 408454
rect 191382 408218 226826 408454
rect 227062 408218 227146 408454
rect 227382 408218 262826 408454
rect 263062 408218 263146 408454
rect 263382 408218 298826 408454
rect 299062 408218 299146 408454
rect 299382 408218 334826 408454
rect 335062 408218 335146 408454
rect 335382 408218 370826 408454
rect 371062 408218 371146 408454
rect 371382 408218 406826 408454
rect 407062 408218 407146 408454
rect 407382 408218 442826 408454
rect 443062 408218 443146 408454
rect 443382 408218 478826 408454
rect 479062 408218 479146 408454
rect 479382 408218 514826 408454
rect 515062 408218 515146 408454
rect 515382 408218 550826 408454
rect 551062 408218 551146 408454
rect 551382 408218 587262 408454
rect 587498 408218 587582 408454
rect 587818 408218 592650 408454
rect -8726 408134 592650 408218
rect -8726 407898 -3894 408134
rect -3658 407898 -3574 408134
rect -3338 407898 10826 408134
rect 11062 407898 11146 408134
rect 11382 407898 46826 408134
rect 47062 407898 47146 408134
rect 47382 407898 82826 408134
rect 83062 407898 83146 408134
rect 83382 407898 118826 408134
rect 119062 407898 119146 408134
rect 119382 407898 154826 408134
rect 155062 407898 155146 408134
rect 155382 407898 190826 408134
rect 191062 407898 191146 408134
rect 191382 407898 226826 408134
rect 227062 407898 227146 408134
rect 227382 407898 262826 408134
rect 263062 407898 263146 408134
rect 263382 407898 298826 408134
rect 299062 407898 299146 408134
rect 299382 407898 334826 408134
rect 335062 407898 335146 408134
rect 335382 407898 370826 408134
rect 371062 407898 371146 408134
rect 371382 407898 406826 408134
rect 407062 407898 407146 408134
rect 407382 407898 442826 408134
rect 443062 407898 443146 408134
rect 443382 407898 478826 408134
rect 479062 407898 479146 408134
rect 479382 407898 514826 408134
rect 515062 407898 515146 408134
rect 515382 407898 550826 408134
rect 551062 407898 551146 408134
rect 551382 407898 587262 408134
rect 587498 407898 587582 408134
rect 587818 407898 592650 408134
rect -8726 407866 592650 407898
rect -8726 403954 592650 403986
rect -8726 403718 -2934 403954
rect -2698 403718 -2614 403954
rect -2378 403718 6326 403954
rect 6562 403718 6646 403954
rect 6882 403718 42326 403954
rect 42562 403718 42646 403954
rect 42882 403718 78326 403954
rect 78562 403718 78646 403954
rect 78882 403718 114326 403954
rect 114562 403718 114646 403954
rect 114882 403718 150326 403954
rect 150562 403718 150646 403954
rect 150882 403718 186326 403954
rect 186562 403718 186646 403954
rect 186882 403718 222326 403954
rect 222562 403718 222646 403954
rect 222882 403718 258326 403954
rect 258562 403718 258646 403954
rect 258882 403718 294326 403954
rect 294562 403718 294646 403954
rect 294882 403718 330326 403954
rect 330562 403718 330646 403954
rect 330882 403718 366326 403954
rect 366562 403718 366646 403954
rect 366882 403718 402326 403954
rect 402562 403718 402646 403954
rect 402882 403718 438326 403954
rect 438562 403718 438646 403954
rect 438882 403718 474326 403954
rect 474562 403718 474646 403954
rect 474882 403718 510326 403954
rect 510562 403718 510646 403954
rect 510882 403718 546326 403954
rect 546562 403718 546646 403954
rect 546882 403718 582326 403954
rect 582562 403718 582646 403954
rect 582882 403718 586302 403954
rect 586538 403718 586622 403954
rect 586858 403718 592650 403954
rect -8726 403634 592650 403718
rect -8726 403398 -2934 403634
rect -2698 403398 -2614 403634
rect -2378 403398 6326 403634
rect 6562 403398 6646 403634
rect 6882 403398 42326 403634
rect 42562 403398 42646 403634
rect 42882 403398 78326 403634
rect 78562 403398 78646 403634
rect 78882 403398 114326 403634
rect 114562 403398 114646 403634
rect 114882 403398 150326 403634
rect 150562 403398 150646 403634
rect 150882 403398 186326 403634
rect 186562 403398 186646 403634
rect 186882 403398 222326 403634
rect 222562 403398 222646 403634
rect 222882 403398 258326 403634
rect 258562 403398 258646 403634
rect 258882 403398 294326 403634
rect 294562 403398 294646 403634
rect 294882 403398 330326 403634
rect 330562 403398 330646 403634
rect 330882 403398 366326 403634
rect 366562 403398 366646 403634
rect 366882 403398 402326 403634
rect 402562 403398 402646 403634
rect 402882 403398 438326 403634
rect 438562 403398 438646 403634
rect 438882 403398 474326 403634
rect 474562 403398 474646 403634
rect 474882 403398 510326 403634
rect 510562 403398 510646 403634
rect 510882 403398 546326 403634
rect 546562 403398 546646 403634
rect 546882 403398 582326 403634
rect 582562 403398 582646 403634
rect 582882 403398 586302 403634
rect 586538 403398 586622 403634
rect 586858 403398 592650 403634
rect -8726 403366 592650 403398
rect -8726 399454 592650 399486
rect -8726 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 73826 399454
rect 74062 399218 74146 399454
rect 74382 399218 109826 399454
rect 110062 399218 110146 399454
rect 110382 399218 145826 399454
rect 146062 399218 146146 399454
rect 146382 399218 181826 399454
rect 182062 399218 182146 399454
rect 182382 399218 217826 399454
rect 218062 399218 218146 399454
rect 218382 399218 253826 399454
rect 254062 399218 254146 399454
rect 254382 399218 289826 399454
rect 290062 399218 290146 399454
rect 290382 399218 325826 399454
rect 326062 399218 326146 399454
rect 326382 399218 361826 399454
rect 362062 399218 362146 399454
rect 362382 399218 397826 399454
rect 398062 399218 398146 399454
rect 398382 399218 433826 399454
rect 434062 399218 434146 399454
rect 434382 399218 469826 399454
rect 470062 399218 470146 399454
rect 470382 399218 505826 399454
rect 506062 399218 506146 399454
rect 506382 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 592650 399454
rect -8726 399134 592650 399218
rect -8726 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 73826 399134
rect 74062 398898 74146 399134
rect 74382 398898 109826 399134
rect 110062 398898 110146 399134
rect 110382 398898 145826 399134
rect 146062 398898 146146 399134
rect 146382 398898 181826 399134
rect 182062 398898 182146 399134
rect 182382 398898 217826 399134
rect 218062 398898 218146 399134
rect 218382 398898 253826 399134
rect 254062 398898 254146 399134
rect 254382 398898 289826 399134
rect 290062 398898 290146 399134
rect 290382 398898 325826 399134
rect 326062 398898 326146 399134
rect 326382 398898 361826 399134
rect 362062 398898 362146 399134
rect 362382 398898 397826 399134
rect 398062 398898 398146 399134
rect 398382 398898 433826 399134
rect 434062 398898 434146 399134
rect 434382 398898 469826 399134
rect 470062 398898 470146 399134
rect 470382 398898 505826 399134
rect 506062 398898 506146 399134
rect 506382 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 592650 399134
rect -8726 398866 592650 398898
rect -8726 394954 592650 394986
rect -8726 394718 -8694 394954
rect -8458 394718 -8374 394954
rect -8138 394718 33326 394954
rect 33562 394718 33646 394954
rect 33882 394718 69326 394954
rect 69562 394718 69646 394954
rect 69882 394718 105326 394954
rect 105562 394718 105646 394954
rect 105882 394718 141326 394954
rect 141562 394718 141646 394954
rect 141882 394718 177326 394954
rect 177562 394718 177646 394954
rect 177882 394718 213326 394954
rect 213562 394718 213646 394954
rect 213882 394718 249326 394954
rect 249562 394718 249646 394954
rect 249882 394718 285326 394954
rect 285562 394718 285646 394954
rect 285882 394718 321326 394954
rect 321562 394718 321646 394954
rect 321882 394718 357326 394954
rect 357562 394718 357646 394954
rect 357882 394718 393326 394954
rect 393562 394718 393646 394954
rect 393882 394718 429326 394954
rect 429562 394718 429646 394954
rect 429882 394718 465326 394954
rect 465562 394718 465646 394954
rect 465882 394718 501326 394954
rect 501562 394718 501646 394954
rect 501882 394718 537326 394954
rect 537562 394718 537646 394954
rect 537882 394718 573326 394954
rect 573562 394718 573646 394954
rect 573882 394718 592062 394954
rect 592298 394718 592382 394954
rect 592618 394718 592650 394954
rect -8726 394634 592650 394718
rect -8726 394398 -8694 394634
rect -8458 394398 -8374 394634
rect -8138 394398 33326 394634
rect 33562 394398 33646 394634
rect 33882 394398 69326 394634
rect 69562 394398 69646 394634
rect 69882 394398 105326 394634
rect 105562 394398 105646 394634
rect 105882 394398 141326 394634
rect 141562 394398 141646 394634
rect 141882 394398 177326 394634
rect 177562 394398 177646 394634
rect 177882 394398 213326 394634
rect 213562 394398 213646 394634
rect 213882 394398 249326 394634
rect 249562 394398 249646 394634
rect 249882 394398 285326 394634
rect 285562 394398 285646 394634
rect 285882 394398 321326 394634
rect 321562 394398 321646 394634
rect 321882 394398 357326 394634
rect 357562 394398 357646 394634
rect 357882 394398 393326 394634
rect 393562 394398 393646 394634
rect 393882 394398 429326 394634
rect 429562 394398 429646 394634
rect 429882 394398 465326 394634
rect 465562 394398 465646 394634
rect 465882 394398 501326 394634
rect 501562 394398 501646 394634
rect 501882 394398 537326 394634
rect 537562 394398 537646 394634
rect 537882 394398 573326 394634
rect 573562 394398 573646 394634
rect 573882 394398 592062 394634
rect 592298 394398 592382 394634
rect 592618 394398 592650 394634
rect -8726 394366 592650 394398
rect -8726 390454 592650 390486
rect -8726 390218 -7734 390454
rect -7498 390218 -7414 390454
rect -7178 390218 28826 390454
rect 29062 390218 29146 390454
rect 29382 390218 64826 390454
rect 65062 390218 65146 390454
rect 65382 390218 100826 390454
rect 101062 390218 101146 390454
rect 101382 390218 136826 390454
rect 137062 390218 137146 390454
rect 137382 390218 172826 390454
rect 173062 390218 173146 390454
rect 173382 390218 208826 390454
rect 209062 390218 209146 390454
rect 209382 390218 244826 390454
rect 245062 390218 245146 390454
rect 245382 390218 280826 390454
rect 281062 390218 281146 390454
rect 281382 390218 316826 390454
rect 317062 390218 317146 390454
rect 317382 390218 352826 390454
rect 353062 390218 353146 390454
rect 353382 390218 388826 390454
rect 389062 390218 389146 390454
rect 389382 390218 424826 390454
rect 425062 390218 425146 390454
rect 425382 390218 460826 390454
rect 461062 390218 461146 390454
rect 461382 390218 496826 390454
rect 497062 390218 497146 390454
rect 497382 390218 532826 390454
rect 533062 390218 533146 390454
rect 533382 390218 568826 390454
rect 569062 390218 569146 390454
rect 569382 390218 591102 390454
rect 591338 390218 591422 390454
rect 591658 390218 592650 390454
rect -8726 390134 592650 390218
rect -8726 389898 -7734 390134
rect -7498 389898 -7414 390134
rect -7178 389898 28826 390134
rect 29062 389898 29146 390134
rect 29382 389898 64826 390134
rect 65062 389898 65146 390134
rect 65382 389898 100826 390134
rect 101062 389898 101146 390134
rect 101382 389898 136826 390134
rect 137062 389898 137146 390134
rect 137382 389898 172826 390134
rect 173062 389898 173146 390134
rect 173382 389898 208826 390134
rect 209062 389898 209146 390134
rect 209382 389898 244826 390134
rect 245062 389898 245146 390134
rect 245382 389898 280826 390134
rect 281062 389898 281146 390134
rect 281382 389898 316826 390134
rect 317062 389898 317146 390134
rect 317382 389898 352826 390134
rect 353062 389898 353146 390134
rect 353382 389898 388826 390134
rect 389062 389898 389146 390134
rect 389382 389898 424826 390134
rect 425062 389898 425146 390134
rect 425382 389898 460826 390134
rect 461062 389898 461146 390134
rect 461382 389898 496826 390134
rect 497062 389898 497146 390134
rect 497382 389898 532826 390134
rect 533062 389898 533146 390134
rect 533382 389898 568826 390134
rect 569062 389898 569146 390134
rect 569382 389898 591102 390134
rect 591338 389898 591422 390134
rect 591658 389898 592650 390134
rect -8726 389866 592650 389898
rect -8726 385954 592650 385986
rect -8726 385718 -6774 385954
rect -6538 385718 -6454 385954
rect -6218 385718 24326 385954
rect 24562 385718 24646 385954
rect 24882 385718 60326 385954
rect 60562 385718 60646 385954
rect 60882 385718 96326 385954
rect 96562 385718 96646 385954
rect 96882 385718 132326 385954
rect 132562 385718 132646 385954
rect 132882 385718 168326 385954
rect 168562 385718 168646 385954
rect 168882 385718 204326 385954
rect 204562 385718 204646 385954
rect 204882 385718 240326 385954
rect 240562 385718 240646 385954
rect 240882 385718 276326 385954
rect 276562 385718 276646 385954
rect 276882 385718 312326 385954
rect 312562 385718 312646 385954
rect 312882 385718 348326 385954
rect 348562 385718 348646 385954
rect 348882 385718 384326 385954
rect 384562 385718 384646 385954
rect 384882 385718 420326 385954
rect 420562 385718 420646 385954
rect 420882 385718 456326 385954
rect 456562 385718 456646 385954
rect 456882 385718 492326 385954
rect 492562 385718 492646 385954
rect 492882 385718 528326 385954
rect 528562 385718 528646 385954
rect 528882 385718 564326 385954
rect 564562 385718 564646 385954
rect 564882 385718 590142 385954
rect 590378 385718 590462 385954
rect 590698 385718 592650 385954
rect -8726 385634 592650 385718
rect -8726 385398 -6774 385634
rect -6538 385398 -6454 385634
rect -6218 385398 24326 385634
rect 24562 385398 24646 385634
rect 24882 385398 60326 385634
rect 60562 385398 60646 385634
rect 60882 385398 96326 385634
rect 96562 385398 96646 385634
rect 96882 385398 132326 385634
rect 132562 385398 132646 385634
rect 132882 385398 168326 385634
rect 168562 385398 168646 385634
rect 168882 385398 204326 385634
rect 204562 385398 204646 385634
rect 204882 385398 240326 385634
rect 240562 385398 240646 385634
rect 240882 385398 276326 385634
rect 276562 385398 276646 385634
rect 276882 385398 312326 385634
rect 312562 385398 312646 385634
rect 312882 385398 348326 385634
rect 348562 385398 348646 385634
rect 348882 385398 384326 385634
rect 384562 385398 384646 385634
rect 384882 385398 420326 385634
rect 420562 385398 420646 385634
rect 420882 385398 456326 385634
rect 456562 385398 456646 385634
rect 456882 385398 492326 385634
rect 492562 385398 492646 385634
rect 492882 385398 528326 385634
rect 528562 385398 528646 385634
rect 528882 385398 564326 385634
rect 564562 385398 564646 385634
rect 564882 385398 590142 385634
rect 590378 385398 590462 385634
rect 590698 385398 592650 385634
rect -8726 385366 592650 385398
rect -8726 381454 592650 381486
rect -8726 381218 -5814 381454
rect -5578 381218 -5494 381454
rect -5258 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 55826 381454
rect 56062 381218 56146 381454
rect 56382 381218 91826 381454
rect 92062 381218 92146 381454
rect 92382 381218 127826 381454
rect 128062 381218 128146 381454
rect 128382 381218 163826 381454
rect 164062 381218 164146 381454
rect 164382 381218 199826 381454
rect 200062 381218 200146 381454
rect 200382 381218 235826 381454
rect 236062 381218 236146 381454
rect 236382 381218 271826 381454
rect 272062 381218 272146 381454
rect 272382 381218 307826 381454
rect 308062 381218 308146 381454
rect 308382 381218 343826 381454
rect 344062 381218 344146 381454
rect 344382 381218 379826 381454
rect 380062 381218 380146 381454
rect 380382 381218 415826 381454
rect 416062 381218 416146 381454
rect 416382 381218 451826 381454
rect 452062 381218 452146 381454
rect 452382 381218 487826 381454
rect 488062 381218 488146 381454
rect 488382 381218 523826 381454
rect 524062 381218 524146 381454
rect 524382 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 589182 381454
rect 589418 381218 589502 381454
rect 589738 381218 592650 381454
rect -8726 381134 592650 381218
rect -8726 380898 -5814 381134
rect -5578 380898 -5494 381134
rect -5258 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 55826 381134
rect 56062 380898 56146 381134
rect 56382 380898 91826 381134
rect 92062 380898 92146 381134
rect 92382 380898 127826 381134
rect 128062 380898 128146 381134
rect 128382 380898 163826 381134
rect 164062 380898 164146 381134
rect 164382 380898 199826 381134
rect 200062 380898 200146 381134
rect 200382 380898 235826 381134
rect 236062 380898 236146 381134
rect 236382 380898 271826 381134
rect 272062 380898 272146 381134
rect 272382 380898 307826 381134
rect 308062 380898 308146 381134
rect 308382 380898 343826 381134
rect 344062 380898 344146 381134
rect 344382 380898 379826 381134
rect 380062 380898 380146 381134
rect 380382 380898 415826 381134
rect 416062 380898 416146 381134
rect 416382 380898 451826 381134
rect 452062 380898 452146 381134
rect 452382 380898 487826 381134
rect 488062 380898 488146 381134
rect 488382 380898 523826 381134
rect 524062 380898 524146 381134
rect 524382 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 589182 381134
rect 589418 380898 589502 381134
rect 589738 380898 592650 381134
rect -8726 380866 592650 380898
rect -8726 376954 592650 376986
rect -8726 376718 -4854 376954
rect -4618 376718 -4534 376954
rect -4298 376718 15326 376954
rect 15562 376718 15646 376954
rect 15882 376718 51326 376954
rect 51562 376718 51646 376954
rect 51882 376718 87326 376954
rect 87562 376718 87646 376954
rect 87882 376718 123326 376954
rect 123562 376718 123646 376954
rect 123882 376718 159326 376954
rect 159562 376718 159646 376954
rect 159882 376718 195326 376954
rect 195562 376718 195646 376954
rect 195882 376718 231326 376954
rect 231562 376718 231646 376954
rect 231882 376718 267326 376954
rect 267562 376718 267646 376954
rect 267882 376718 303326 376954
rect 303562 376718 303646 376954
rect 303882 376718 339326 376954
rect 339562 376718 339646 376954
rect 339882 376718 375326 376954
rect 375562 376718 375646 376954
rect 375882 376718 411326 376954
rect 411562 376718 411646 376954
rect 411882 376718 447326 376954
rect 447562 376718 447646 376954
rect 447882 376718 483326 376954
rect 483562 376718 483646 376954
rect 483882 376718 519326 376954
rect 519562 376718 519646 376954
rect 519882 376718 555326 376954
rect 555562 376718 555646 376954
rect 555882 376718 588222 376954
rect 588458 376718 588542 376954
rect 588778 376718 592650 376954
rect -8726 376634 592650 376718
rect -8726 376398 -4854 376634
rect -4618 376398 -4534 376634
rect -4298 376398 15326 376634
rect 15562 376398 15646 376634
rect 15882 376398 51326 376634
rect 51562 376398 51646 376634
rect 51882 376398 87326 376634
rect 87562 376398 87646 376634
rect 87882 376398 123326 376634
rect 123562 376398 123646 376634
rect 123882 376398 159326 376634
rect 159562 376398 159646 376634
rect 159882 376398 195326 376634
rect 195562 376398 195646 376634
rect 195882 376398 231326 376634
rect 231562 376398 231646 376634
rect 231882 376398 267326 376634
rect 267562 376398 267646 376634
rect 267882 376398 303326 376634
rect 303562 376398 303646 376634
rect 303882 376398 339326 376634
rect 339562 376398 339646 376634
rect 339882 376398 375326 376634
rect 375562 376398 375646 376634
rect 375882 376398 411326 376634
rect 411562 376398 411646 376634
rect 411882 376398 447326 376634
rect 447562 376398 447646 376634
rect 447882 376398 483326 376634
rect 483562 376398 483646 376634
rect 483882 376398 519326 376634
rect 519562 376398 519646 376634
rect 519882 376398 555326 376634
rect 555562 376398 555646 376634
rect 555882 376398 588222 376634
rect 588458 376398 588542 376634
rect 588778 376398 592650 376634
rect -8726 376366 592650 376398
rect -8726 372454 592650 372486
rect -8726 372218 -3894 372454
rect -3658 372218 -3574 372454
rect -3338 372218 10826 372454
rect 11062 372218 11146 372454
rect 11382 372218 46826 372454
rect 47062 372218 47146 372454
rect 47382 372218 82826 372454
rect 83062 372218 83146 372454
rect 83382 372218 118826 372454
rect 119062 372218 119146 372454
rect 119382 372218 154826 372454
rect 155062 372218 155146 372454
rect 155382 372218 190826 372454
rect 191062 372218 191146 372454
rect 191382 372218 226826 372454
rect 227062 372218 227146 372454
rect 227382 372218 262826 372454
rect 263062 372218 263146 372454
rect 263382 372218 298826 372454
rect 299062 372218 299146 372454
rect 299382 372218 334826 372454
rect 335062 372218 335146 372454
rect 335382 372218 370826 372454
rect 371062 372218 371146 372454
rect 371382 372218 406826 372454
rect 407062 372218 407146 372454
rect 407382 372218 442826 372454
rect 443062 372218 443146 372454
rect 443382 372218 478826 372454
rect 479062 372218 479146 372454
rect 479382 372218 514826 372454
rect 515062 372218 515146 372454
rect 515382 372218 550826 372454
rect 551062 372218 551146 372454
rect 551382 372218 587262 372454
rect 587498 372218 587582 372454
rect 587818 372218 592650 372454
rect -8726 372134 592650 372218
rect -8726 371898 -3894 372134
rect -3658 371898 -3574 372134
rect -3338 371898 10826 372134
rect 11062 371898 11146 372134
rect 11382 371898 46826 372134
rect 47062 371898 47146 372134
rect 47382 371898 82826 372134
rect 83062 371898 83146 372134
rect 83382 371898 118826 372134
rect 119062 371898 119146 372134
rect 119382 371898 154826 372134
rect 155062 371898 155146 372134
rect 155382 371898 190826 372134
rect 191062 371898 191146 372134
rect 191382 371898 226826 372134
rect 227062 371898 227146 372134
rect 227382 371898 262826 372134
rect 263062 371898 263146 372134
rect 263382 371898 298826 372134
rect 299062 371898 299146 372134
rect 299382 371898 334826 372134
rect 335062 371898 335146 372134
rect 335382 371898 370826 372134
rect 371062 371898 371146 372134
rect 371382 371898 406826 372134
rect 407062 371898 407146 372134
rect 407382 371898 442826 372134
rect 443062 371898 443146 372134
rect 443382 371898 478826 372134
rect 479062 371898 479146 372134
rect 479382 371898 514826 372134
rect 515062 371898 515146 372134
rect 515382 371898 550826 372134
rect 551062 371898 551146 372134
rect 551382 371898 587262 372134
rect 587498 371898 587582 372134
rect 587818 371898 592650 372134
rect -8726 371866 592650 371898
rect -8726 367954 592650 367986
rect -8726 367718 -2934 367954
rect -2698 367718 -2614 367954
rect -2378 367718 6326 367954
rect 6562 367718 6646 367954
rect 6882 367718 42326 367954
rect 42562 367718 42646 367954
rect 42882 367718 78326 367954
rect 78562 367718 78646 367954
rect 78882 367718 114326 367954
rect 114562 367718 114646 367954
rect 114882 367718 150326 367954
rect 150562 367718 150646 367954
rect 150882 367718 186326 367954
rect 186562 367718 186646 367954
rect 186882 367718 222326 367954
rect 222562 367718 222646 367954
rect 222882 367718 258326 367954
rect 258562 367718 258646 367954
rect 258882 367718 294326 367954
rect 294562 367718 294646 367954
rect 294882 367718 330326 367954
rect 330562 367718 330646 367954
rect 330882 367718 366326 367954
rect 366562 367718 366646 367954
rect 366882 367718 402326 367954
rect 402562 367718 402646 367954
rect 402882 367718 438326 367954
rect 438562 367718 438646 367954
rect 438882 367718 474326 367954
rect 474562 367718 474646 367954
rect 474882 367718 510326 367954
rect 510562 367718 510646 367954
rect 510882 367718 546326 367954
rect 546562 367718 546646 367954
rect 546882 367718 582326 367954
rect 582562 367718 582646 367954
rect 582882 367718 586302 367954
rect 586538 367718 586622 367954
rect 586858 367718 592650 367954
rect -8726 367634 592650 367718
rect -8726 367398 -2934 367634
rect -2698 367398 -2614 367634
rect -2378 367398 6326 367634
rect 6562 367398 6646 367634
rect 6882 367398 42326 367634
rect 42562 367398 42646 367634
rect 42882 367398 78326 367634
rect 78562 367398 78646 367634
rect 78882 367398 114326 367634
rect 114562 367398 114646 367634
rect 114882 367398 150326 367634
rect 150562 367398 150646 367634
rect 150882 367398 186326 367634
rect 186562 367398 186646 367634
rect 186882 367398 222326 367634
rect 222562 367398 222646 367634
rect 222882 367398 258326 367634
rect 258562 367398 258646 367634
rect 258882 367398 294326 367634
rect 294562 367398 294646 367634
rect 294882 367398 330326 367634
rect 330562 367398 330646 367634
rect 330882 367398 366326 367634
rect 366562 367398 366646 367634
rect 366882 367398 402326 367634
rect 402562 367398 402646 367634
rect 402882 367398 438326 367634
rect 438562 367398 438646 367634
rect 438882 367398 474326 367634
rect 474562 367398 474646 367634
rect 474882 367398 510326 367634
rect 510562 367398 510646 367634
rect 510882 367398 546326 367634
rect 546562 367398 546646 367634
rect 546882 367398 582326 367634
rect 582562 367398 582646 367634
rect 582882 367398 586302 367634
rect 586538 367398 586622 367634
rect 586858 367398 592650 367634
rect -8726 367366 592650 367398
rect -8726 363454 592650 363486
rect -8726 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 73826 363454
rect 74062 363218 74146 363454
rect 74382 363218 109826 363454
rect 110062 363218 110146 363454
rect 110382 363218 145826 363454
rect 146062 363218 146146 363454
rect 146382 363218 181826 363454
rect 182062 363218 182146 363454
rect 182382 363218 217826 363454
rect 218062 363218 218146 363454
rect 218382 363218 253826 363454
rect 254062 363218 254146 363454
rect 254382 363218 289826 363454
rect 290062 363218 290146 363454
rect 290382 363218 325826 363454
rect 326062 363218 326146 363454
rect 326382 363218 361826 363454
rect 362062 363218 362146 363454
rect 362382 363218 397826 363454
rect 398062 363218 398146 363454
rect 398382 363218 433826 363454
rect 434062 363218 434146 363454
rect 434382 363218 469826 363454
rect 470062 363218 470146 363454
rect 470382 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 592650 363454
rect -8726 363134 592650 363218
rect -8726 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 73826 363134
rect 74062 362898 74146 363134
rect 74382 362898 109826 363134
rect 110062 362898 110146 363134
rect 110382 362898 145826 363134
rect 146062 362898 146146 363134
rect 146382 362898 181826 363134
rect 182062 362898 182146 363134
rect 182382 362898 217826 363134
rect 218062 362898 218146 363134
rect 218382 362898 253826 363134
rect 254062 362898 254146 363134
rect 254382 362898 289826 363134
rect 290062 362898 290146 363134
rect 290382 362898 325826 363134
rect 326062 362898 326146 363134
rect 326382 362898 361826 363134
rect 362062 362898 362146 363134
rect 362382 362898 397826 363134
rect 398062 362898 398146 363134
rect 398382 362898 433826 363134
rect 434062 362898 434146 363134
rect 434382 362898 469826 363134
rect 470062 362898 470146 363134
rect 470382 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 592650 363134
rect -8726 362866 592650 362898
rect -8726 358954 592650 358986
rect -8726 358718 -8694 358954
rect -8458 358718 -8374 358954
rect -8138 358718 33326 358954
rect 33562 358718 33646 358954
rect 33882 358718 69326 358954
rect 69562 358718 69646 358954
rect 69882 358718 105326 358954
rect 105562 358718 105646 358954
rect 105882 358718 141326 358954
rect 141562 358718 141646 358954
rect 141882 358718 177326 358954
rect 177562 358718 177646 358954
rect 177882 358718 213326 358954
rect 213562 358718 213646 358954
rect 213882 358718 249326 358954
rect 249562 358718 249646 358954
rect 249882 358718 285326 358954
rect 285562 358718 285646 358954
rect 285882 358718 321326 358954
rect 321562 358718 321646 358954
rect 321882 358718 357326 358954
rect 357562 358718 357646 358954
rect 357882 358718 393326 358954
rect 393562 358718 393646 358954
rect 393882 358718 429326 358954
rect 429562 358718 429646 358954
rect 429882 358718 465326 358954
rect 465562 358718 465646 358954
rect 465882 358718 501326 358954
rect 501562 358718 501646 358954
rect 501882 358718 537326 358954
rect 537562 358718 537646 358954
rect 537882 358718 573326 358954
rect 573562 358718 573646 358954
rect 573882 358718 592062 358954
rect 592298 358718 592382 358954
rect 592618 358718 592650 358954
rect -8726 358634 592650 358718
rect -8726 358398 -8694 358634
rect -8458 358398 -8374 358634
rect -8138 358398 33326 358634
rect 33562 358398 33646 358634
rect 33882 358398 69326 358634
rect 69562 358398 69646 358634
rect 69882 358398 105326 358634
rect 105562 358398 105646 358634
rect 105882 358398 141326 358634
rect 141562 358398 141646 358634
rect 141882 358398 177326 358634
rect 177562 358398 177646 358634
rect 177882 358398 213326 358634
rect 213562 358398 213646 358634
rect 213882 358398 249326 358634
rect 249562 358398 249646 358634
rect 249882 358398 285326 358634
rect 285562 358398 285646 358634
rect 285882 358398 321326 358634
rect 321562 358398 321646 358634
rect 321882 358398 357326 358634
rect 357562 358398 357646 358634
rect 357882 358398 393326 358634
rect 393562 358398 393646 358634
rect 393882 358398 429326 358634
rect 429562 358398 429646 358634
rect 429882 358398 465326 358634
rect 465562 358398 465646 358634
rect 465882 358398 501326 358634
rect 501562 358398 501646 358634
rect 501882 358398 537326 358634
rect 537562 358398 537646 358634
rect 537882 358398 573326 358634
rect 573562 358398 573646 358634
rect 573882 358398 592062 358634
rect 592298 358398 592382 358634
rect 592618 358398 592650 358634
rect -8726 358366 592650 358398
rect -8726 354454 592650 354486
rect -8726 354218 -7734 354454
rect -7498 354218 -7414 354454
rect -7178 354218 28826 354454
rect 29062 354218 29146 354454
rect 29382 354218 64826 354454
rect 65062 354218 65146 354454
rect 65382 354218 100826 354454
rect 101062 354218 101146 354454
rect 101382 354218 136826 354454
rect 137062 354218 137146 354454
rect 137382 354218 172826 354454
rect 173062 354218 173146 354454
rect 173382 354218 208826 354454
rect 209062 354218 209146 354454
rect 209382 354218 244826 354454
rect 245062 354218 245146 354454
rect 245382 354218 280826 354454
rect 281062 354218 281146 354454
rect 281382 354218 316826 354454
rect 317062 354218 317146 354454
rect 317382 354218 352826 354454
rect 353062 354218 353146 354454
rect 353382 354218 388826 354454
rect 389062 354218 389146 354454
rect 389382 354218 424826 354454
rect 425062 354218 425146 354454
rect 425382 354218 460826 354454
rect 461062 354218 461146 354454
rect 461382 354218 496826 354454
rect 497062 354218 497146 354454
rect 497382 354218 532826 354454
rect 533062 354218 533146 354454
rect 533382 354218 568826 354454
rect 569062 354218 569146 354454
rect 569382 354218 591102 354454
rect 591338 354218 591422 354454
rect 591658 354218 592650 354454
rect -8726 354134 592650 354218
rect -8726 353898 -7734 354134
rect -7498 353898 -7414 354134
rect -7178 353898 28826 354134
rect 29062 353898 29146 354134
rect 29382 353898 64826 354134
rect 65062 353898 65146 354134
rect 65382 353898 100826 354134
rect 101062 353898 101146 354134
rect 101382 353898 136826 354134
rect 137062 353898 137146 354134
rect 137382 353898 172826 354134
rect 173062 353898 173146 354134
rect 173382 353898 208826 354134
rect 209062 353898 209146 354134
rect 209382 353898 244826 354134
rect 245062 353898 245146 354134
rect 245382 353898 280826 354134
rect 281062 353898 281146 354134
rect 281382 353898 316826 354134
rect 317062 353898 317146 354134
rect 317382 353898 352826 354134
rect 353062 353898 353146 354134
rect 353382 353898 388826 354134
rect 389062 353898 389146 354134
rect 389382 353898 424826 354134
rect 425062 353898 425146 354134
rect 425382 353898 460826 354134
rect 461062 353898 461146 354134
rect 461382 353898 496826 354134
rect 497062 353898 497146 354134
rect 497382 353898 532826 354134
rect 533062 353898 533146 354134
rect 533382 353898 568826 354134
rect 569062 353898 569146 354134
rect 569382 353898 591102 354134
rect 591338 353898 591422 354134
rect 591658 353898 592650 354134
rect -8726 353866 592650 353898
rect -8726 349954 592650 349986
rect -8726 349718 -6774 349954
rect -6538 349718 -6454 349954
rect -6218 349718 24326 349954
rect 24562 349718 24646 349954
rect 24882 349718 60326 349954
rect 60562 349718 60646 349954
rect 60882 349718 96326 349954
rect 96562 349718 96646 349954
rect 96882 349718 132326 349954
rect 132562 349718 132646 349954
rect 132882 349718 168326 349954
rect 168562 349718 168646 349954
rect 168882 349718 204326 349954
rect 204562 349718 204646 349954
rect 204882 349718 240326 349954
rect 240562 349718 240646 349954
rect 240882 349718 276326 349954
rect 276562 349718 276646 349954
rect 276882 349718 312326 349954
rect 312562 349718 312646 349954
rect 312882 349718 348326 349954
rect 348562 349718 348646 349954
rect 348882 349718 384326 349954
rect 384562 349718 384646 349954
rect 384882 349718 420326 349954
rect 420562 349718 420646 349954
rect 420882 349718 456326 349954
rect 456562 349718 456646 349954
rect 456882 349718 492326 349954
rect 492562 349718 492646 349954
rect 492882 349718 528326 349954
rect 528562 349718 528646 349954
rect 528882 349718 564326 349954
rect 564562 349718 564646 349954
rect 564882 349718 590142 349954
rect 590378 349718 590462 349954
rect 590698 349718 592650 349954
rect -8726 349634 592650 349718
rect -8726 349398 -6774 349634
rect -6538 349398 -6454 349634
rect -6218 349398 24326 349634
rect 24562 349398 24646 349634
rect 24882 349398 60326 349634
rect 60562 349398 60646 349634
rect 60882 349398 96326 349634
rect 96562 349398 96646 349634
rect 96882 349398 132326 349634
rect 132562 349398 132646 349634
rect 132882 349398 168326 349634
rect 168562 349398 168646 349634
rect 168882 349398 204326 349634
rect 204562 349398 204646 349634
rect 204882 349398 240326 349634
rect 240562 349398 240646 349634
rect 240882 349398 276326 349634
rect 276562 349398 276646 349634
rect 276882 349398 312326 349634
rect 312562 349398 312646 349634
rect 312882 349398 348326 349634
rect 348562 349398 348646 349634
rect 348882 349398 384326 349634
rect 384562 349398 384646 349634
rect 384882 349398 420326 349634
rect 420562 349398 420646 349634
rect 420882 349398 456326 349634
rect 456562 349398 456646 349634
rect 456882 349398 492326 349634
rect 492562 349398 492646 349634
rect 492882 349398 528326 349634
rect 528562 349398 528646 349634
rect 528882 349398 564326 349634
rect 564562 349398 564646 349634
rect 564882 349398 590142 349634
rect 590378 349398 590462 349634
rect 590698 349398 592650 349634
rect -8726 349366 592650 349398
rect -8726 345454 592650 345486
rect -8726 345218 -5814 345454
rect -5578 345218 -5494 345454
rect -5258 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 55826 345454
rect 56062 345218 56146 345454
rect 56382 345218 91826 345454
rect 92062 345218 92146 345454
rect 92382 345218 127826 345454
rect 128062 345218 128146 345454
rect 128382 345218 163826 345454
rect 164062 345218 164146 345454
rect 164382 345218 199826 345454
rect 200062 345218 200146 345454
rect 200382 345218 235826 345454
rect 236062 345218 236146 345454
rect 236382 345218 271826 345454
rect 272062 345218 272146 345454
rect 272382 345218 307826 345454
rect 308062 345218 308146 345454
rect 308382 345218 343826 345454
rect 344062 345218 344146 345454
rect 344382 345218 379826 345454
rect 380062 345218 380146 345454
rect 380382 345218 415826 345454
rect 416062 345218 416146 345454
rect 416382 345218 451826 345454
rect 452062 345218 452146 345454
rect 452382 345218 487826 345454
rect 488062 345218 488146 345454
rect 488382 345218 523826 345454
rect 524062 345218 524146 345454
rect 524382 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 589182 345454
rect 589418 345218 589502 345454
rect 589738 345218 592650 345454
rect -8726 345134 592650 345218
rect -8726 344898 -5814 345134
rect -5578 344898 -5494 345134
rect -5258 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 55826 345134
rect 56062 344898 56146 345134
rect 56382 344898 91826 345134
rect 92062 344898 92146 345134
rect 92382 344898 127826 345134
rect 128062 344898 128146 345134
rect 128382 344898 163826 345134
rect 164062 344898 164146 345134
rect 164382 344898 199826 345134
rect 200062 344898 200146 345134
rect 200382 344898 235826 345134
rect 236062 344898 236146 345134
rect 236382 344898 271826 345134
rect 272062 344898 272146 345134
rect 272382 344898 307826 345134
rect 308062 344898 308146 345134
rect 308382 344898 343826 345134
rect 344062 344898 344146 345134
rect 344382 344898 379826 345134
rect 380062 344898 380146 345134
rect 380382 344898 415826 345134
rect 416062 344898 416146 345134
rect 416382 344898 451826 345134
rect 452062 344898 452146 345134
rect 452382 344898 487826 345134
rect 488062 344898 488146 345134
rect 488382 344898 523826 345134
rect 524062 344898 524146 345134
rect 524382 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 589182 345134
rect 589418 344898 589502 345134
rect 589738 344898 592650 345134
rect -8726 344866 592650 344898
rect -8726 340954 592650 340986
rect -8726 340718 -4854 340954
rect -4618 340718 -4534 340954
rect -4298 340718 15326 340954
rect 15562 340718 15646 340954
rect 15882 340718 51326 340954
rect 51562 340718 51646 340954
rect 51882 340718 87326 340954
rect 87562 340718 87646 340954
rect 87882 340718 123326 340954
rect 123562 340718 123646 340954
rect 123882 340718 159326 340954
rect 159562 340718 159646 340954
rect 159882 340718 195326 340954
rect 195562 340718 195646 340954
rect 195882 340718 231326 340954
rect 231562 340718 231646 340954
rect 231882 340718 267326 340954
rect 267562 340718 267646 340954
rect 267882 340718 303326 340954
rect 303562 340718 303646 340954
rect 303882 340718 339326 340954
rect 339562 340718 339646 340954
rect 339882 340718 375326 340954
rect 375562 340718 375646 340954
rect 375882 340718 411326 340954
rect 411562 340718 411646 340954
rect 411882 340718 447326 340954
rect 447562 340718 447646 340954
rect 447882 340718 483326 340954
rect 483562 340718 483646 340954
rect 483882 340718 519326 340954
rect 519562 340718 519646 340954
rect 519882 340718 555326 340954
rect 555562 340718 555646 340954
rect 555882 340718 588222 340954
rect 588458 340718 588542 340954
rect 588778 340718 592650 340954
rect -8726 340634 592650 340718
rect -8726 340398 -4854 340634
rect -4618 340398 -4534 340634
rect -4298 340398 15326 340634
rect 15562 340398 15646 340634
rect 15882 340398 51326 340634
rect 51562 340398 51646 340634
rect 51882 340398 87326 340634
rect 87562 340398 87646 340634
rect 87882 340398 123326 340634
rect 123562 340398 123646 340634
rect 123882 340398 159326 340634
rect 159562 340398 159646 340634
rect 159882 340398 195326 340634
rect 195562 340398 195646 340634
rect 195882 340398 231326 340634
rect 231562 340398 231646 340634
rect 231882 340398 267326 340634
rect 267562 340398 267646 340634
rect 267882 340398 303326 340634
rect 303562 340398 303646 340634
rect 303882 340398 339326 340634
rect 339562 340398 339646 340634
rect 339882 340398 375326 340634
rect 375562 340398 375646 340634
rect 375882 340398 411326 340634
rect 411562 340398 411646 340634
rect 411882 340398 447326 340634
rect 447562 340398 447646 340634
rect 447882 340398 483326 340634
rect 483562 340398 483646 340634
rect 483882 340398 519326 340634
rect 519562 340398 519646 340634
rect 519882 340398 555326 340634
rect 555562 340398 555646 340634
rect 555882 340398 588222 340634
rect 588458 340398 588542 340634
rect 588778 340398 592650 340634
rect -8726 340366 592650 340398
rect -8726 336454 592650 336486
rect -8726 336218 -3894 336454
rect -3658 336218 -3574 336454
rect -3338 336218 10826 336454
rect 11062 336218 11146 336454
rect 11382 336218 46826 336454
rect 47062 336218 47146 336454
rect 47382 336218 82826 336454
rect 83062 336218 83146 336454
rect 83382 336218 118826 336454
rect 119062 336218 119146 336454
rect 119382 336218 154826 336454
rect 155062 336218 155146 336454
rect 155382 336218 190826 336454
rect 191062 336218 191146 336454
rect 191382 336218 226826 336454
rect 227062 336218 227146 336454
rect 227382 336218 262826 336454
rect 263062 336218 263146 336454
rect 263382 336218 298826 336454
rect 299062 336218 299146 336454
rect 299382 336218 334826 336454
rect 335062 336218 335146 336454
rect 335382 336218 370826 336454
rect 371062 336218 371146 336454
rect 371382 336218 406826 336454
rect 407062 336218 407146 336454
rect 407382 336218 442826 336454
rect 443062 336218 443146 336454
rect 443382 336218 478826 336454
rect 479062 336218 479146 336454
rect 479382 336218 514826 336454
rect 515062 336218 515146 336454
rect 515382 336218 550826 336454
rect 551062 336218 551146 336454
rect 551382 336218 587262 336454
rect 587498 336218 587582 336454
rect 587818 336218 592650 336454
rect -8726 336134 592650 336218
rect -8726 335898 -3894 336134
rect -3658 335898 -3574 336134
rect -3338 335898 10826 336134
rect 11062 335898 11146 336134
rect 11382 335898 46826 336134
rect 47062 335898 47146 336134
rect 47382 335898 82826 336134
rect 83062 335898 83146 336134
rect 83382 335898 118826 336134
rect 119062 335898 119146 336134
rect 119382 335898 154826 336134
rect 155062 335898 155146 336134
rect 155382 335898 190826 336134
rect 191062 335898 191146 336134
rect 191382 335898 226826 336134
rect 227062 335898 227146 336134
rect 227382 335898 262826 336134
rect 263062 335898 263146 336134
rect 263382 335898 298826 336134
rect 299062 335898 299146 336134
rect 299382 335898 334826 336134
rect 335062 335898 335146 336134
rect 335382 335898 370826 336134
rect 371062 335898 371146 336134
rect 371382 335898 406826 336134
rect 407062 335898 407146 336134
rect 407382 335898 442826 336134
rect 443062 335898 443146 336134
rect 443382 335898 478826 336134
rect 479062 335898 479146 336134
rect 479382 335898 514826 336134
rect 515062 335898 515146 336134
rect 515382 335898 550826 336134
rect 551062 335898 551146 336134
rect 551382 335898 587262 336134
rect 587498 335898 587582 336134
rect 587818 335898 592650 336134
rect -8726 335866 592650 335898
rect -8726 331954 592650 331986
rect -8726 331718 -2934 331954
rect -2698 331718 -2614 331954
rect -2378 331718 6326 331954
rect 6562 331718 6646 331954
rect 6882 331718 42326 331954
rect 42562 331718 42646 331954
rect 42882 331718 78326 331954
rect 78562 331718 78646 331954
rect 78882 331718 114326 331954
rect 114562 331718 114646 331954
rect 114882 331718 150326 331954
rect 150562 331718 150646 331954
rect 150882 331718 186326 331954
rect 186562 331718 186646 331954
rect 186882 331718 222326 331954
rect 222562 331718 222646 331954
rect 222882 331718 258326 331954
rect 258562 331718 258646 331954
rect 258882 331718 294326 331954
rect 294562 331718 294646 331954
rect 294882 331718 330326 331954
rect 330562 331718 330646 331954
rect 330882 331718 366326 331954
rect 366562 331718 366646 331954
rect 366882 331718 402326 331954
rect 402562 331718 402646 331954
rect 402882 331718 438326 331954
rect 438562 331718 438646 331954
rect 438882 331718 474326 331954
rect 474562 331718 474646 331954
rect 474882 331718 510326 331954
rect 510562 331718 510646 331954
rect 510882 331718 546326 331954
rect 546562 331718 546646 331954
rect 546882 331718 582326 331954
rect 582562 331718 582646 331954
rect 582882 331718 586302 331954
rect 586538 331718 586622 331954
rect 586858 331718 592650 331954
rect -8726 331634 592650 331718
rect -8726 331398 -2934 331634
rect -2698 331398 -2614 331634
rect -2378 331398 6326 331634
rect 6562 331398 6646 331634
rect 6882 331398 42326 331634
rect 42562 331398 42646 331634
rect 42882 331398 78326 331634
rect 78562 331398 78646 331634
rect 78882 331398 114326 331634
rect 114562 331398 114646 331634
rect 114882 331398 150326 331634
rect 150562 331398 150646 331634
rect 150882 331398 186326 331634
rect 186562 331398 186646 331634
rect 186882 331398 222326 331634
rect 222562 331398 222646 331634
rect 222882 331398 258326 331634
rect 258562 331398 258646 331634
rect 258882 331398 294326 331634
rect 294562 331398 294646 331634
rect 294882 331398 330326 331634
rect 330562 331398 330646 331634
rect 330882 331398 366326 331634
rect 366562 331398 366646 331634
rect 366882 331398 402326 331634
rect 402562 331398 402646 331634
rect 402882 331398 438326 331634
rect 438562 331398 438646 331634
rect 438882 331398 474326 331634
rect 474562 331398 474646 331634
rect 474882 331398 510326 331634
rect 510562 331398 510646 331634
rect 510882 331398 546326 331634
rect 546562 331398 546646 331634
rect 546882 331398 582326 331634
rect 582562 331398 582646 331634
rect 582882 331398 586302 331634
rect 586538 331398 586622 331634
rect 586858 331398 592650 331634
rect -8726 331366 592650 331398
rect -8726 327454 592650 327486
rect -8726 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 73826 327454
rect 74062 327218 74146 327454
rect 74382 327218 109826 327454
rect 110062 327218 110146 327454
rect 110382 327218 145826 327454
rect 146062 327218 146146 327454
rect 146382 327218 181826 327454
rect 182062 327218 182146 327454
rect 182382 327218 217826 327454
rect 218062 327218 218146 327454
rect 218382 327218 253826 327454
rect 254062 327218 254146 327454
rect 254382 327218 289826 327454
rect 290062 327218 290146 327454
rect 290382 327218 325826 327454
rect 326062 327218 326146 327454
rect 326382 327218 361826 327454
rect 362062 327218 362146 327454
rect 362382 327218 397826 327454
rect 398062 327218 398146 327454
rect 398382 327218 433826 327454
rect 434062 327218 434146 327454
rect 434382 327218 469826 327454
rect 470062 327218 470146 327454
rect 470382 327218 505826 327454
rect 506062 327218 506146 327454
rect 506382 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 592650 327454
rect -8726 327134 592650 327218
rect -8726 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 73826 327134
rect 74062 326898 74146 327134
rect 74382 326898 109826 327134
rect 110062 326898 110146 327134
rect 110382 326898 145826 327134
rect 146062 326898 146146 327134
rect 146382 326898 181826 327134
rect 182062 326898 182146 327134
rect 182382 326898 217826 327134
rect 218062 326898 218146 327134
rect 218382 326898 253826 327134
rect 254062 326898 254146 327134
rect 254382 326898 289826 327134
rect 290062 326898 290146 327134
rect 290382 326898 325826 327134
rect 326062 326898 326146 327134
rect 326382 326898 361826 327134
rect 362062 326898 362146 327134
rect 362382 326898 397826 327134
rect 398062 326898 398146 327134
rect 398382 326898 433826 327134
rect 434062 326898 434146 327134
rect 434382 326898 469826 327134
rect 470062 326898 470146 327134
rect 470382 326898 505826 327134
rect 506062 326898 506146 327134
rect 506382 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 592650 327134
rect -8726 326866 592650 326898
rect -8726 322954 592650 322986
rect -8726 322718 -8694 322954
rect -8458 322718 -8374 322954
rect -8138 322718 33326 322954
rect 33562 322718 33646 322954
rect 33882 322718 69326 322954
rect 69562 322718 69646 322954
rect 69882 322718 105326 322954
rect 105562 322718 105646 322954
rect 105882 322718 141326 322954
rect 141562 322718 141646 322954
rect 141882 322718 177326 322954
rect 177562 322718 177646 322954
rect 177882 322718 213326 322954
rect 213562 322718 213646 322954
rect 213882 322718 249326 322954
rect 249562 322718 249646 322954
rect 249882 322718 285326 322954
rect 285562 322718 285646 322954
rect 285882 322718 321326 322954
rect 321562 322718 321646 322954
rect 321882 322718 357326 322954
rect 357562 322718 357646 322954
rect 357882 322718 393326 322954
rect 393562 322718 393646 322954
rect 393882 322718 429326 322954
rect 429562 322718 429646 322954
rect 429882 322718 465326 322954
rect 465562 322718 465646 322954
rect 465882 322718 501326 322954
rect 501562 322718 501646 322954
rect 501882 322718 537326 322954
rect 537562 322718 537646 322954
rect 537882 322718 573326 322954
rect 573562 322718 573646 322954
rect 573882 322718 592062 322954
rect 592298 322718 592382 322954
rect 592618 322718 592650 322954
rect -8726 322634 592650 322718
rect -8726 322398 -8694 322634
rect -8458 322398 -8374 322634
rect -8138 322398 33326 322634
rect 33562 322398 33646 322634
rect 33882 322398 69326 322634
rect 69562 322398 69646 322634
rect 69882 322398 105326 322634
rect 105562 322398 105646 322634
rect 105882 322398 141326 322634
rect 141562 322398 141646 322634
rect 141882 322398 177326 322634
rect 177562 322398 177646 322634
rect 177882 322398 213326 322634
rect 213562 322398 213646 322634
rect 213882 322398 249326 322634
rect 249562 322398 249646 322634
rect 249882 322398 285326 322634
rect 285562 322398 285646 322634
rect 285882 322398 321326 322634
rect 321562 322398 321646 322634
rect 321882 322398 357326 322634
rect 357562 322398 357646 322634
rect 357882 322398 393326 322634
rect 393562 322398 393646 322634
rect 393882 322398 429326 322634
rect 429562 322398 429646 322634
rect 429882 322398 465326 322634
rect 465562 322398 465646 322634
rect 465882 322398 501326 322634
rect 501562 322398 501646 322634
rect 501882 322398 537326 322634
rect 537562 322398 537646 322634
rect 537882 322398 573326 322634
rect 573562 322398 573646 322634
rect 573882 322398 592062 322634
rect 592298 322398 592382 322634
rect 592618 322398 592650 322634
rect -8726 322366 592650 322398
rect -8726 318454 592650 318486
rect -8726 318218 -7734 318454
rect -7498 318218 -7414 318454
rect -7178 318218 28826 318454
rect 29062 318218 29146 318454
rect 29382 318218 64826 318454
rect 65062 318218 65146 318454
rect 65382 318218 100826 318454
rect 101062 318218 101146 318454
rect 101382 318218 136826 318454
rect 137062 318218 137146 318454
rect 137382 318218 172826 318454
rect 173062 318218 173146 318454
rect 173382 318218 208826 318454
rect 209062 318218 209146 318454
rect 209382 318218 244826 318454
rect 245062 318218 245146 318454
rect 245382 318218 280826 318454
rect 281062 318218 281146 318454
rect 281382 318218 316826 318454
rect 317062 318218 317146 318454
rect 317382 318218 352826 318454
rect 353062 318218 353146 318454
rect 353382 318218 388826 318454
rect 389062 318218 389146 318454
rect 389382 318218 424826 318454
rect 425062 318218 425146 318454
rect 425382 318218 460826 318454
rect 461062 318218 461146 318454
rect 461382 318218 496826 318454
rect 497062 318218 497146 318454
rect 497382 318218 532826 318454
rect 533062 318218 533146 318454
rect 533382 318218 568826 318454
rect 569062 318218 569146 318454
rect 569382 318218 591102 318454
rect 591338 318218 591422 318454
rect 591658 318218 592650 318454
rect -8726 318134 592650 318218
rect -8726 317898 -7734 318134
rect -7498 317898 -7414 318134
rect -7178 317898 28826 318134
rect 29062 317898 29146 318134
rect 29382 317898 64826 318134
rect 65062 317898 65146 318134
rect 65382 317898 100826 318134
rect 101062 317898 101146 318134
rect 101382 317898 136826 318134
rect 137062 317898 137146 318134
rect 137382 317898 172826 318134
rect 173062 317898 173146 318134
rect 173382 317898 208826 318134
rect 209062 317898 209146 318134
rect 209382 317898 244826 318134
rect 245062 317898 245146 318134
rect 245382 317898 280826 318134
rect 281062 317898 281146 318134
rect 281382 317898 316826 318134
rect 317062 317898 317146 318134
rect 317382 317898 352826 318134
rect 353062 317898 353146 318134
rect 353382 317898 388826 318134
rect 389062 317898 389146 318134
rect 389382 317898 424826 318134
rect 425062 317898 425146 318134
rect 425382 317898 460826 318134
rect 461062 317898 461146 318134
rect 461382 317898 496826 318134
rect 497062 317898 497146 318134
rect 497382 317898 532826 318134
rect 533062 317898 533146 318134
rect 533382 317898 568826 318134
rect 569062 317898 569146 318134
rect 569382 317898 591102 318134
rect 591338 317898 591422 318134
rect 591658 317898 592650 318134
rect -8726 317866 592650 317898
rect -8726 313954 592650 313986
rect -8726 313718 -6774 313954
rect -6538 313718 -6454 313954
rect -6218 313718 24326 313954
rect 24562 313718 24646 313954
rect 24882 313718 60326 313954
rect 60562 313718 60646 313954
rect 60882 313718 96326 313954
rect 96562 313718 96646 313954
rect 96882 313718 132326 313954
rect 132562 313718 132646 313954
rect 132882 313718 168326 313954
rect 168562 313718 168646 313954
rect 168882 313718 204326 313954
rect 204562 313718 204646 313954
rect 204882 313718 240326 313954
rect 240562 313718 240646 313954
rect 240882 313718 276326 313954
rect 276562 313718 276646 313954
rect 276882 313718 312326 313954
rect 312562 313718 312646 313954
rect 312882 313718 348326 313954
rect 348562 313718 348646 313954
rect 348882 313718 384326 313954
rect 384562 313718 384646 313954
rect 384882 313718 420326 313954
rect 420562 313718 420646 313954
rect 420882 313718 456326 313954
rect 456562 313718 456646 313954
rect 456882 313718 492326 313954
rect 492562 313718 492646 313954
rect 492882 313718 528326 313954
rect 528562 313718 528646 313954
rect 528882 313718 564326 313954
rect 564562 313718 564646 313954
rect 564882 313718 590142 313954
rect 590378 313718 590462 313954
rect 590698 313718 592650 313954
rect -8726 313634 592650 313718
rect -8726 313398 -6774 313634
rect -6538 313398 -6454 313634
rect -6218 313398 24326 313634
rect 24562 313398 24646 313634
rect 24882 313398 60326 313634
rect 60562 313398 60646 313634
rect 60882 313398 96326 313634
rect 96562 313398 96646 313634
rect 96882 313398 132326 313634
rect 132562 313398 132646 313634
rect 132882 313398 168326 313634
rect 168562 313398 168646 313634
rect 168882 313398 204326 313634
rect 204562 313398 204646 313634
rect 204882 313398 240326 313634
rect 240562 313398 240646 313634
rect 240882 313398 276326 313634
rect 276562 313398 276646 313634
rect 276882 313398 312326 313634
rect 312562 313398 312646 313634
rect 312882 313398 348326 313634
rect 348562 313398 348646 313634
rect 348882 313398 384326 313634
rect 384562 313398 384646 313634
rect 384882 313398 420326 313634
rect 420562 313398 420646 313634
rect 420882 313398 456326 313634
rect 456562 313398 456646 313634
rect 456882 313398 492326 313634
rect 492562 313398 492646 313634
rect 492882 313398 528326 313634
rect 528562 313398 528646 313634
rect 528882 313398 564326 313634
rect 564562 313398 564646 313634
rect 564882 313398 590142 313634
rect 590378 313398 590462 313634
rect 590698 313398 592650 313634
rect -8726 313366 592650 313398
rect -8726 309454 592650 309486
rect -8726 309218 -5814 309454
rect -5578 309218 -5494 309454
rect -5258 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 55826 309454
rect 56062 309218 56146 309454
rect 56382 309218 91826 309454
rect 92062 309218 92146 309454
rect 92382 309218 127826 309454
rect 128062 309218 128146 309454
rect 128382 309218 163826 309454
rect 164062 309218 164146 309454
rect 164382 309218 199826 309454
rect 200062 309218 200146 309454
rect 200382 309218 235826 309454
rect 236062 309218 236146 309454
rect 236382 309218 271826 309454
rect 272062 309218 272146 309454
rect 272382 309218 307826 309454
rect 308062 309218 308146 309454
rect 308382 309218 343826 309454
rect 344062 309218 344146 309454
rect 344382 309218 379826 309454
rect 380062 309218 380146 309454
rect 380382 309218 415826 309454
rect 416062 309218 416146 309454
rect 416382 309218 451826 309454
rect 452062 309218 452146 309454
rect 452382 309218 487826 309454
rect 488062 309218 488146 309454
rect 488382 309218 523826 309454
rect 524062 309218 524146 309454
rect 524382 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 589182 309454
rect 589418 309218 589502 309454
rect 589738 309218 592650 309454
rect -8726 309134 592650 309218
rect -8726 308898 -5814 309134
rect -5578 308898 -5494 309134
rect -5258 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 55826 309134
rect 56062 308898 56146 309134
rect 56382 308898 91826 309134
rect 92062 308898 92146 309134
rect 92382 308898 127826 309134
rect 128062 308898 128146 309134
rect 128382 308898 163826 309134
rect 164062 308898 164146 309134
rect 164382 308898 199826 309134
rect 200062 308898 200146 309134
rect 200382 308898 235826 309134
rect 236062 308898 236146 309134
rect 236382 308898 271826 309134
rect 272062 308898 272146 309134
rect 272382 308898 307826 309134
rect 308062 308898 308146 309134
rect 308382 308898 343826 309134
rect 344062 308898 344146 309134
rect 344382 308898 379826 309134
rect 380062 308898 380146 309134
rect 380382 308898 415826 309134
rect 416062 308898 416146 309134
rect 416382 308898 451826 309134
rect 452062 308898 452146 309134
rect 452382 308898 487826 309134
rect 488062 308898 488146 309134
rect 488382 308898 523826 309134
rect 524062 308898 524146 309134
rect 524382 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 589182 309134
rect 589418 308898 589502 309134
rect 589738 308898 592650 309134
rect -8726 308866 592650 308898
rect -8726 304954 592650 304986
rect -8726 304718 -4854 304954
rect -4618 304718 -4534 304954
rect -4298 304718 15326 304954
rect 15562 304718 15646 304954
rect 15882 304718 51326 304954
rect 51562 304718 51646 304954
rect 51882 304718 87326 304954
rect 87562 304718 87646 304954
rect 87882 304718 123326 304954
rect 123562 304718 123646 304954
rect 123882 304718 159326 304954
rect 159562 304718 159646 304954
rect 159882 304718 195326 304954
rect 195562 304718 195646 304954
rect 195882 304718 231326 304954
rect 231562 304718 231646 304954
rect 231882 304718 267326 304954
rect 267562 304718 267646 304954
rect 267882 304718 303326 304954
rect 303562 304718 303646 304954
rect 303882 304718 339326 304954
rect 339562 304718 339646 304954
rect 339882 304718 375326 304954
rect 375562 304718 375646 304954
rect 375882 304718 411326 304954
rect 411562 304718 411646 304954
rect 411882 304718 447326 304954
rect 447562 304718 447646 304954
rect 447882 304718 483326 304954
rect 483562 304718 483646 304954
rect 483882 304718 519326 304954
rect 519562 304718 519646 304954
rect 519882 304718 555326 304954
rect 555562 304718 555646 304954
rect 555882 304718 588222 304954
rect 588458 304718 588542 304954
rect 588778 304718 592650 304954
rect -8726 304634 592650 304718
rect -8726 304398 -4854 304634
rect -4618 304398 -4534 304634
rect -4298 304398 15326 304634
rect 15562 304398 15646 304634
rect 15882 304398 51326 304634
rect 51562 304398 51646 304634
rect 51882 304398 87326 304634
rect 87562 304398 87646 304634
rect 87882 304398 123326 304634
rect 123562 304398 123646 304634
rect 123882 304398 159326 304634
rect 159562 304398 159646 304634
rect 159882 304398 195326 304634
rect 195562 304398 195646 304634
rect 195882 304398 231326 304634
rect 231562 304398 231646 304634
rect 231882 304398 267326 304634
rect 267562 304398 267646 304634
rect 267882 304398 303326 304634
rect 303562 304398 303646 304634
rect 303882 304398 339326 304634
rect 339562 304398 339646 304634
rect 339882 304398 375326 304634
rect 375562 304398 375646 304634
rect 375882 304398 411326 304634
rect 411562 304398 411646 304634
rect 411882 304398 447326 304634
rect 447562 304398 447646 304634
rect 447882 304398 483326 304634
rect 483562 304398 483646 304634
rect 483882 304398 519326 304634
rect 519562 304398 519646 304634
rect 519882 304398 555326 304634
rect 555562 304398 555646 304634
rect 555882 304398 588222 304634
rect 588458 304398 588542 304634
rect 588778 304398 592650 304634
rect -8726 304366 592650 304398
rect -8726 300454 592650 300486
rect -8726 300218 -3894 300454
rect -3658 300218 -3574 300454
rect -3338 300218 10826 300454
rect 11062 300218 11146 300454
rect 11382 300218 46826 300454
rect 47062 300218 47146 300454
rect 47382 300218 82826 300454
rect 83062 300218 83146 300454
rect 83382 300218 118826 300454
rect 119062 300218 119146 300454
rect 119382 300218 154826 300454
rect 155062 300218 155146 300454
rect 155382 300218 190826 300454
rect 191062 300218 191146 300454
rect 191382 300218 226826 300454
rect 227062 300218 227146 300454
rect 227382 300218 262826 300454
rect 263062 300218 263146 300454
rect 263382 300218 298826 300454
rect 299062 300218 299146 300454
rect 299382 300218 334826 300454
rect 335062 300218 335146 300454
rect 335382 300218 370826 300454
rect 371062 300218 371146 300454
rect 371382 300218 406826 300454
rect 407062 300218 407146 300454
rect 407382 300218 442826 300454
rect 443062 300218 443146 300454
rect 443382 300218 478826 300454
rect 479062 300218 479146 300454
rect 479382 300218 514826 300454
rect 515062 300218 515146 300454
rect 515382 300218 550826 300454
rect 551062 300218 551146 300454
rect 551382 300218 587262 300454
rect 587498 300218 587582 300454
rect 587818 300218 592650 300454
rect -8726 300134 592650 300218
rect -8726 299898 -3894 300134
rect -3658 299898 -3574 300134
rect -3338 299898 10826 300134
rect 11062 299898 11146 300134
rect 11382 299898 46826 300134
rect 47062 299898 47146 300134
rect 47382 299898 82826 300134
rect 83062 299898 83146 300134
rect 83382 299898 118826 300134
rect 119062 299898 119146 300134
rect 119382 299898 154826 300134
rect 155062 299898 155146 300134
rect 155382 299898 190826 300134
rect 191062 299898 191146 300134
rect 191382 299898 226826 300134
rect 227062 299898 227146 300134
rect 227382 299898 262826 300134
rect 263062 299898 263146 300134
rect 263382 299898 298826 300134
rect 299062 299898 299146 300134
rect 299382 299898 334826 300134
rect 335062 299898 335146 300134
rect 335382 299898 370826 300134
rect 371062 299898 371146 300134
rect 371382 299898 406826 300134
rect 407062 299898 407146 300134
rect 407382 299898 442826 300134
rect 443062 299898 443146 300134
rect 443382 299898 478826 300134
rect 479062 299898 479146 300134
rect 479382 299898 514826 300134
rect 515062 299898 515146 300134
rect 515382 299898 550826 300134
rect 551062 299898 551146 300134
rect 551382 299898 587262 300134
rect 587498 299898 587582 300134
rect 587818 299898 592650 300134
rect -8726 299866 592650 299898
rect -8726 295954 592650 295986
rect -8726 295718 -2934 295954
rect -2698 295718 -2614 295954
rect -2378 295718 6326 295954
rect 6562 295718 6646 295954
rect 6882 295718 42326 295954
rect 42562 295718 42646 295954
rect 42882 295718 78326 295954
rect 78562 295718 78646 295954
rect 78882 295718 114326 295954
rect 114562 295718 114646 295954
rect 114882 295718 150326 295954
rect 150562 295718 150646 295954
rect 150882 295718 186326 295954
rect 186562 295718 186646 295954
rect 186882 295718 222326 295954
rect 222562 295718 222646 295954
rect 222882 295718 258326 295954
rect 258562 295718 258646 295954
rect 258882 295718 294326 295954
rect 294562 295718 294646 295954
rect 294882 295718 330326 295954
rect 330562 295718 330646 295954
rect 330882 295718 366326 295954
rect 366562 295718 366646 295954
rect 366882 295718 402326 295954
rect 402562 295718 402646 295954
rect 402882 295718 438326 295954
rect 438562 295718 438646 295954
rect 438882 295718 474326 295954
rect 474562 295718 474646 295954
rect 474882 295718 510326 295954
rect 510562 295718 510646 295954
rect 510882 295718 546326 295954
rect 546562 295718 546646 295954
rect 546882 295718 582326 295954
rect 582562 295718 582646 295954
rect 582882 295718 586302 295954
rect 586538 295718 586622 295954
rect 586858 295718 592650 295954
rect -8726 295634 592650 295718
rect -8726 295398 -2934 295634
rect -2698 295398 -2614 295634
rect -2378 295398 6326 295634
rect 6562 295398 6646 295634
rect 6882 295398 42326 295634
rect 42562 295398 42646 295634
rect 42882 295398 78326 295634
rect 78562 295398 78646 295634
rect 78882 295398 114326 295634
rect 114562 295398 114646 295634
rect 114882 295398 150326 295634
rect 150562 295398 150646 295634
rect 150882 295398 186326 295634
rect 186562 295398 186646 295634
rect 186882 295398 222326 295634
rect 222562 295398 222646 295634
rect 222882 295398 258326 295634
rect 258562 295398 258646 295634
rect 258882 295398 294326 295634
rect 294562 295398 294646 295634
rect 294882 295398 330326 295634
rect 330562 295398 330646 295634
rect 330882 295398 366326 295634
rect 366562 295398 366646 295634
rect 366882 295398 402326 295634
rect 402562 295398 402646 295634
rect 402882 295398 438326 295634
rect 438562 295398 438646 295634
rect 438882 295398 474326 295634
rect 474562 295398 474646 295634
rect 474882 295398 510326 295634
rect 510562 295398 510646 295634
rect 510882 295398 546326 295634
rect 546562 295398 546646 295634
rect 546882 295398 582326 295634
rect 582562 295398 582646 295634
rect 582882 295398 586302 295634
rect 586538 295398 586622 295634
rect 586858 295398 592650 295634
rect -8726 295366 592650 295398
rect -8726 291454 592650 291486
rect -8726 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 73826 291454
rect 74062 291218 74146 291454
rect 74382 291218 109826 291454
rect 110062 291218 110146 291454
rect 110382 291218 145826 291454
rect 146062 291218 146146 291454
rect 146382 291218 181826 291454
rect 182062 291218 182146 291454
rect 182382 291218 217826 291454
rect 218062 291218 218146 291454
rect 218382 291218 253826 291454
rect 254062 291218 254146 291454
rect 254382 291218 289826 291454
rect 290062 291218 290146 291454
rect 290382 291218 325826 291454
rect 326062 291218 326146 291454
rect 326382 291218 361826 291454
rect 362062 291218 362146 291454
rect 362382 291218 397826 291454
rect 398062 291218 398146 291454
rect 398382 291218 433826 291454
rect 434062 291218 434146 291454
rect 434382 291218 469826 291454
rect 470062 291218 470146 291454
rect 470382 291218 505826 291454
rect 506062 291218 506146 291454
rect 506382 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 592650 291454
rect -8726 291134 592650 291218
rect -8726 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 73826 291134
rect 74062 290898 74146 291134
rect 74382 290898 109826 291134
rect 110062 290898 110146 291134
rect 110382 290898 145826 291134
rect 146062 290898 146146 291134
rect 146382 290898 181826 291134
rect 182062 290898 182146 291134
rect 182382 290898 217826 291134
rect 218062 290898 218146 291134
rect 218382 290898 253826 291134
rect 254062 290898 254146 291134
rect 254382 290898 289826 291134
rect 290062 290898 290146 291134
rect 290382 290898 325826 291134
rect 326062 290898 326146 291134
rect 326382 290898 361826 291134
rect 362062 290898 362146 291134
rect 362382 290898 397826 291134
rect 398062 290898 398146 291134
rect 398382 290898 433826 291134
rect 434062 290898 434146 291134
rect 434382 290898 469826 291134
rect 470062 290898 470146 291134
rect 470382 290898 505826 291134
rect 506062 290898 506146 291134
rect 506382 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 592650 291134
rect -8726 290866 592650 290898
rect -8726 286954 592650 286986
rect -8726 286718 -8694 286954
rect -8458 286718 -8374 286954
rect -8138 286718 33326 286954
rect 33562 286718 33646 286954
rect 33882 286718 69326 286954
rect 69562 286718 69646 286954
rect 69882 286718 105326 286954
rect 105562 286718 105646 286954
rect 105882 286718 141326 286954
rect 141562 286718 141646 286954
rect 141882 286718 177326 286954
rect 177562 286718 177646 286954
rect 177882 286718 213326 286954
rect 213562 286718 213646 286954
rect 213882 286718 249326 286954
rect 249562 286718 249646 286954
rect 249882 286718 285326 286954
rect 285562 286718 285646 286954
rect 285882 286718 321326 286954
rect 321562 286718 321646 286954
rect 321882 286718 357326 286954
rect 357562 286718 357646 286954
rect 357882 286718 393326 286954
rect 393562 286718 393646 286954
rect 393882 286718 429326 286954
rect 429562 286718 429646 286954
rect 429882 286718 465326 286954
rect 465562 286718 465646 286954
rect 465882 286718 501326 286954
rect 501562 286718 501646 286954
rect 501882 286718 537326 286954
rect 537562 286718 537646 286954
rect 537882 286718 573326 286954
rect 573562 286718 573646 286954
rect 573882 286718 592062 286954
rect 592298 286718 592382 286954
rect 592618 286718 592650 286954
rect -8726 286634 592650 286718
rect -8726 286398 -8694 286634
rect -8458 286398 -8374 286634
rect -8138 286398 33326 286634
rect 33562 286398 33646 286634
rect 33882 286398 69326 286634
rect 69562 286398 69646 286634
rect 69882 286398 105326 286634
rect 105562 286398 105646 286634
rect 105882 286398 141326 286634
rect 141562 286398 141646 286634
rect 141882 286398 177326 286634
rect 177562 286398 177646 286634
rect 177882 286398 213326 286634
rect 213562 286398 213646 286634
rect 213882 286398 249326 286634
rect 249562 286398 249646 286634
rect 249882 286398 285326 286634
rect 285562 286398 285646 286634
rect 285882 286398 321326 286634
rect 321562 286398 321646 286634
rect 321882 286398 357326 286634
rect 357562 286398 357646 286634
rect 357882 286398 393326 286634
rect 393562 286398 393646 286634
rect 393882 286398 429326 286634
rect 429562 286398 429646 286634
rect 429882 286398 465326 286634
rect 465562 286398 465646 286634
rect 465882 286398 501326 286634
rect 501562 286398 501646 286634
rect 501882 286398 537326 286634
rect 537562 286398 537646 286634
rect 537882 286398 573326 286634
rect 573562 286398 573646 286634
rect 573882 286398 592062 286634
rect 592298 286398 592382 286634
rect 592618 286398 592650 286634
rect -8726 286366 592650 286398
rect -8726 282454 592650 282486
rect -8726 282218 -7734 282454
rect -7498 282218 -7414 282454
rect -7178 282218 28826 282454
rect 29062 282218 29146 282454
rect 29382 282218 64826 282454
rect 65062 282218 65146 282454
rect 65382 282218 100826 282454
rect 101062 282218 101146 282454
rect 101382 282218 136826 282454
rect 137062 282218 137146 282454
rect 137382 282218 172826 282454
rect 173062 282218 173146 282454
rect 173382 282218 208826 282454
rect 209062 282218 209146 282454
rect 209382 282218 244826 282454
rect 245062 282218 245146 282454
rect 245382 282218 280826 282454
rect 281062 282218 281146 282454
rect 281382 282218 316826 282454
rect 317062 282218 317146 282454
rect 317382 282218 352826 282454
rect 353062 282218 353146 282454
rect 353382 282218 388826 282454
rect 389062 282218 389146 282454
rect 389382 282218 424826 282454
rect 425062 282218 425146 282454
rect 425382 282218 460826 282454
rect 461062 282218 461146 282454
rect 461382 282218 496826 282454
rect 497062 282218 497146 282454
rect 497382 282218 532826 282454
rect 533062 282218 533146 282454
rect 533382 282218 568826 282454
rect 569062 282218 569146 282454
rect 569382 282218 591102 282454
rect 591338 282218 591422 282454
rect 591658 282218 592650 282454
rect -8726 282134 592650 282218
rect -8726 281898 -7734 282134
rect -7498 281898 -7414 282134
rect -7178 281898 28826 282134
rect 29062 281898 29146 282134
rect 29382 281898 64826 282134
rect 65062 281898 65146 282134
rect 65382 281898 100826 282134
rect 101062 281898 101146 282134
rect 101382 281898 136826 282134
rect 137062 281898 137146 282134
rect 137382 281898 172826 282134
rect 173062 281898 173146 282134
rect 173382 281898 208826 282134
rect 209062 281898 209146 282134
rect 209382 281898 244826 282134
rect 245062 281898 245146 282134
rect 245382 281898 280826 282134
rect 281062 281898 281146 282134
rect 281382 281898 316826 282134
rect 317062 281898 317146 282134
rect 317382 281898 352826 282134
rect 353062 281898 353146 282134
rect 353382 281898 388826 282134
rect 389062 281898 389146 282134
rect 389382 281898 424826 282134
rect 425062 281898 425146 282134
rect 425382 281898 460826 282134
rect 461062 281898 461146 282134
rect 461382 281898 496826 282134
rect 497062 281898 497146 282134
rect 497382 281898 532826 282134
rect 533062 281898 533146 282134
rect 533382 281898 568826 282134
rect 569062 281898 569146 282134
rect 569382 281898 591102 282134
rect 591338 281898 591422 282134
rect 591658 281898 592650 282134
rect -8726 281866 592650 281898
rect -8726 277954 592650 277986
rect -8726 277718 -6774 277954
rect -6538 277718 -6454 277954
rect -6218 277718 24326 277954
rect 24562 277718 24646 277954
rect 24882 277718 60326 277954
rect 60562 277718 60646 277954
rect 60882 277718 96326 277954
rect 96562 277718 96646 277954
rect 96882 277718 132326 277954
rect 132562 277718 132646 277954
rect 132882 277718 168326 277954
rect 168562 277718 168646 277954
rect 168882 277718 204326 277954
rect 204562 277718 204646 277954
rect 204882 277718 240326 277954
rect 240562 277718 240646 277954
rect 240882 277718 276326 277954
rect 276562 277718 276646 277954
rect 276882 277718 312326 277954
rect 312562 277718 312646 277954
rect 312882 277718 348326 277954
rect 348562 277718 348646 277954
rect 348882 277718 384326 277954
rect 384562 277718 384646 277954
rect 384882 277718 420326 277954
rect 420562 277718 420646 277954
rect 420882 277718 456326 277954
rect 456562 277718 456646 277954
rect 456882 277718 492326 277954
rect 492562 277718 492646 277954
rect 492882 277718 528326 277954
rect 528562 277718 528646 277954
rect 528882 277718 564326 277954
rect 564562 277718 564646 277954
rect 564882 277718 590142 277954
rect 590378 277718 590462 277954
rect 590698 277718 592650 277954
rect -8726 277634 592650 277718
rect -8726 277398 -6774 277634
rect -6538 277398 -6454 277634
rect -6218 277398 24326 277634
rect 24562 277398 24646 277634
rect 24882 277398 60326 277634
rect 60562 277398 60646 277634
rect 60882 277398 96326 277634
rect 96562 277398 96646 277634
rect 96882 277398 132326 277634
rect 132562 277398 132646 277634
rect 132882 277398 168326 277634
rect 168562 277398 168646 277634
rect 168882 277398 204326 277634
rect 204562 277398 204646 277634
rect 204882 277398 240326 277634
rect 240562 277398 240646 277634
rect 240882 277398 276326 277634
rect 276562 277398 276646 277634
rect 276882 277398 312326 277634
rect 312562 277398 312646 277634
rect 312882 277398 348326 277634
rect 348562 277398 348646 277634
rect 348882 277398 384326 277634
rect 384562 277398 384646 277634
rect 384882 277398 420326 277634
rect 420562 277398 420646 277634
rect 420882 277398 456326 277634
rect 456562 277398 456646 277634
rect 456882 277398 492326 277634
rect 492562 277398 492646 277634
rect 492882 277398 528326 277634
rect 528562 277398 528646 277634
rect 528882 277398 564326 277634
rect 564562 277398 564646 277634
rect 564882 277398 590142 277634
rect 590378 277398 590462 277634
rect 590698 277398 592650 277634
rect -8726 277366 592650 277398
rect -8726 273454 592650 273486
rect -8726 273218 -5814 273454
rect -5578 273218 -5494 273454
rect -5258 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 55826 273454
rect 56062 273218 56146 273454
rect 56382 273218 91826 273454
rect 92062 273218 92146 273454
rect 92382 273218 127826 273454
rect 128062 273218 128146 273454
rect 128382 273218 163826 273454
rect 164062 273218 164146 273454
rect 164382 273218 199826 273454
rect 200062 273218 200146 273454
rect 200382 273218 235826 273454
rect 236062 273218 236146 273454
rect 236382 273218 271826 273454
rect 272062 273218 272146 273454
rect 272382 273218 307826 273454
rect 308062 273218 308146 273454
rect 308382 273218 343826 273454
rect 344062 273218 344146 273454
rect 344382 273218 379826 273454
rect 380062 273218 380146 273454
rect 380382 273218 415826 273454
rect 416062 273218 416146 273454
rect 416382 273218 451826 273454
rect 452062 273218 452146 273454
rect 452382 273218 487826 273454
rect 488062 273218 488146 273454
rect 488382 273218 523826 273454
rect 524062 273218 524146 273454
rect 524382 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 589182 273454
rect 589418 273218 589502 273454
rect 589738 273218 592650 273454
rect -8726 273134 592650 273218
rect -8726 272898 -5814 273134
rect -5578 272898 -5494 273134
rect -5258 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 55826 273134
rect 56062 272898 56146 273134
rect 56382 272898 91826 273134
rect 92062 272898 92146 273134
rect 92382 272898 127826 273134
rect 128062 272898 128146 273134
rect 128382 272898 163826 273134
rect 164062 272898 164146 273134
rect 164382 272898 199826 273134
rect 200062 272898 200146 273134
rect 200382 272898 235826 273134
rect 236062 272898 236146 273134
rect 236382 272898 271826 273134
rect 272062 272898 272146 273134
rect 272382 272898 307826 273134
rect 308062 272898 308146 273134
rect 308382 272898 343826 273134
rect 344062 272898 344146 273134
rect 344382 272898 379826 273134
rect 380062 272898 380146 273134
rect 380382 272898 415826 273134
rect 416062 272898 416146 273134
rect 416382 272898 451826 273134
rect 452062 272898 452146 273134
rect 452382 272898 487826 273134
rect 488062 272898 488146 273134
rect 488382 272898 523826 273134
rect 524062 272898 524146 273134
rect 524382 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 589182 273134
rect 589418 272898 589502 273134
rect 589738 272898 592650 273134
rect -8726 272866 592650 272898
rect -8726 268954 592650 268986
rect -8726 268718 -4854 268954
rect -4618 268718 -4534 268954
rect -4298 268718 15326 268954
rect 15562 268718 15646 268954
rect 15882 268718 51326 268954
rect 51562 268718 51646 268954
rect 51882 268718 87326 268954
rect 87562 268718 87646 268954
rect 87882 268718 123326 268954
rect 123562 268718 123646 268954
rect 123882 268718 159326 268954
rect 159562 268718 159646 268954
rect 159882 268718 195326 268954
rect 195562 268718 195646 268954
rect 195882 268718 231326 268954
rect 231562 268718 231646 268954
rect 231882 268718 267326 268954
rect 267562 268718 267646 268954
rect 267882 268718 303326 268954
rect 303562 268718 303646 268954
rect 303882 268718 339326 268954
rect 339562 268718 339646 268954
rect 339882 268718 375326 268954
rect 375562 268718 375646 268954
rect 375882 268718 411326 268954
rect 411562 268718 411646 268954
rect 411882 268718 447326 268954
rect 447562 268718 447646 268954
rect 447882 268718 483326 268954
rect 483562 268718 483646 268954
rect 483882 268718 519326 268954
rect 519562 268718 519646 268954
rect 519882 268718 555326 268954
rect 555562 268718 555646 268954
rect 555882 268718 588222 268954
rect 588458 268718 588542 268954
rect 588778 268718 592650 268954
rect -8726 268634 592650 268718
rect -8726 268398 -4854 268634
rect -4618 268398 -4534 268634
rect -4298 268398 15326 268634
rect 15562 268398 15646 268634
rect 15882 268398 51326 268634
rect 51562 268398 51646 268634
rect 51882 268398 87326 268634
rect 87562 268398 87646 268634
rect 87882 268398 123326 268634
rect 123562 268398 123646 268634
rect 123882 268398 159326 268634
rect 159562 268398 159646 268634
rect 159882 268398 195326 268634
rect 195562 268398 195646 268634
rect 195882 268398 231326 268634
rect 231562 268398 231646 268634
rect 231882 268398 267326 268634
rect 267562 268398 267646 268634
rect 267882 268398 303326 268634
rect 303562 268398 303646 268634
rect 303882 268398 339326 268634
rect 339562 268398 339646 268634
rect 339882 268398 375326 268634
rect 375562 268398 375646 268634
rect 375882 268398 411326 268634
rect 411562 268398 411646 268634
rect 411882 268398 447326 268634
rect 447562 268398 447646 268634
rect 447882 268398 483326 268634
rect 483562 268398 483646 268634
rect 483882 268398 519326 268634
rect 519562 268398 519646 268634
rect 519882 268398 555326 268634
rect 555562 268398 555646 268634
rect 555882 268398 588222 268634
rect 588458 268398 588542 268634
rect 588778 268398 592650 268634
rect -8726 268366 592650 268398
rect -8726 264454 592650 264486
rect -8726 264218 -3894 264454
rect -3658 264218 -3574 264454
rect -3338 264218 10826 264454
rect 11062 264218 11146 264454
rect 11382 264218 46826 264454
rect 47062 264218 47146 264454
rect 47382 264218 82826 264454
rect 83062 264218 83146 264454
rect 83382 264218 118826 264454
rect 119062 264218 119146 264454
rect 119382 264218 154826 264454
rect 155062 264218 155146 264454
rect 155382 264218 190826 264454
rect 191062 264218 191146 264454
rect 191382 264218 226826 264454
rect 227062 264218 227146 264454
rect 227382 264218 262826 264454
rect 263062 264218 263146 264454
rect 263382 264218 298826 264454
rect 299062 264218 299146 264454
rect 299382 264218 334826 264454
rect 335062 264218 335146 264454
rect 335382 264218 370826 264454
rect 371062 264218 371146 264454
rect 371382 264218 406826 264454
rect 407062 264218 407146 264454
rect 407382 264218 442826 264454
rect 443062 264218 443146 264454
rect 443382 264218 478826 264454
rect 479062 264218 479146 264454
rect 479382 264218 514826 264454
rect 515062 264218 515146 264454
rect 515382 264218 550826 264454
rect 551062 264218 551146 264454
rect 551382 264218 587262 264454
rect 587498 264218 587582 264454
rect 587818 264218 592650 264454
rect -8726 264134 592650 264218
rect -8726 263898 -3894 264134
rect -3658 263898 -3574 264134
rect -3338 263898 10826 264134
rect 11062 263898 11146 264134
rect 11382 263898 46826 264134
rect 47062 263898 47146 264134
rect 47382 263898 82826 264134
rect 83062 263898 83146 264134
rect 83382 263898 118826 264134
rect 119062 263898 119146 264134
rect 119382 263898 154826 264134
rect 155062 263898 155146 264134
rect 155382 263898 190826 264134
rect 191062 263898 191146 264134
rect 191382 263898 226826 264134
rect 227062 263898 227146 264134
rect 227382 263898 262826 264134
rect 263062 263898 263146 264134
rect 263382 263898 298826 264134
rect 299062 263898 299146 264134
rect 299382 263898 334826 264134
rect 335062 263898 335146 264134
rect 335382 263898 370826 264134
rect 371062 263898 371146 264134
rect 371382 263898 406826 264134
rect 407062 263898 407146 264134
rect 407382 263898 442826 264134
rect 443062 263898 443146 264134
rect 443382 263898 478826 264134
rect 479062 263898 479146 264134
rect 479382 263898 514826 264134
rect 515062 263898 515146 264134
rect 515382 263898 550826 264134
rect 551062 263898 551146 264134
rect 551382 263898 587262 264134
rect 587498 263898 587582 264134
rect 587818 263898 592650 264134
rect -8726 263866 592650 263898
rect -8726 259954 592650 259986
rect -8726 259718 -2934 259954
rect -2698 259718 -2614 259954
rect -2378 259718 6326 259954
rect 6562 259718 6646 259954
rect 6882 259718 42326 259954
rect 42562 259718 42646 259954
rect 42882 259718 78326 259954
rect 78562 259718 78646 259954
rect 78882 259718 114326 259954
rect 114562 259718 114646 259954
rect 114882 259718 222326 259954
rect 222562 259718 222646 259954
rect 222882 259718 258326 259954
rect 258562 259718 258646 259954
rect 258882 259718 294326 259954
rect 294562 259718 294646 259954
rect 294882 259718 330326 259954
rect 330562 259718 330646 259954
rect 330882 259718 366326 259954
rect 366562 259718 366646 259954
rect 366882 259718 402326 259954
rect 402562 259718 402646 259954
rect 402882 259718 438326 259954
rect 438562 259718 438646 259954
rect 438882 259718 474326 259954
rect 474562 259718 474646 259954
rect 474882 259718 510326 259954
rect 510562 259718 510646 259954
rect 510882 259718 546326 259954
rect 546562 259718 546646 259954
rect 546882 259718 582326 259954
rect 582562 259718 582646 259954
rect 582882 259718 586302 259954
rect 586538 259718 586622 259954
rect 586858 259718 592650 259954
rect -8726 259634 592650 259718
rect -8726 259398 -2934 259634
rect -2698 259398 -2614 259634
rect -2378 259398 6326 259634
rect 6562 259398 6646 259634
rect 6882 259398 42326 259634
rect 42562 259398 42646 259634
rect 42882 259398 78326 259634
rect 78562 259398 78646 259634
rect 78882 259398 114326 259634
rect 114562 259398 114646 259634
rect 114882 259398 222326 259634
rect 222562 259398 222646 259634
rect 222882 259398 258326 259634
rect 258562 259398 258646 259634
rect 258882 259398 294326 259634
rect 294562 259398 294646 259634
rect 294882 259398 330326 259634
rect 330562 259398 330646 259634
rect 330882 259398 366326 259634
rect 366562 259398 366646 259634
rect 366882 259398 402326 259634
rect 402562 259398 402646 259634
rect 402882 259398 438326 259634
rect 438562 259398 438646 259634
rect 438882 259398 474326 259634
rect 474562 259398 474646 259634
rect 474882 259398 510326 259634
rect 510562 259398 510646 259634
rect 510882 259398 546326 259634
rect 546562 259398 546646 259634
rect 546882 259398 582326 259634
rect 582562 259398 582646 259634
rect 582882 259398 586302 259634
rect 586538 259398 586622 259634
rect 586858 259398 592650 259634
rect -8726 259366 592650 259398
rect -8726 255454 592650 255486
rect -8726 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 73826 255454
rect 74062 255218 74146 255454
rect 74382 255218 109826 255454
rect 110062 255218 110146 255454
rect 110382 255218 124250 255454
rect 124486 255218 154970 255454
rect 155206 255218 185690 255454
rect 185926 255218 217826 255454
rect 218062 255218 218146 255454
rect 218382 255218 253826 255454
rect 254062 255218 254146 255454
rect 254382 255218 289826 255454
rect 290062 255218 290146 255454
rect 290382 255218 325826 255454
rect 326062 255218 326146 255454
rect 326382 255218 361826 255454
rect 362062 255218 362146 255454
rect 362382 255218 397826 255454
rect 398062 255218 398146 255454
rect 398382 255218 433826 255454
rect 434062 255218 434146 255454
rect 434382 255218 469826 255454
rect 470062 255218 470146 255454
rect 470382 255218 505826 255454
rect 506062 255218 506146 255454
rect 506382 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 592650 255454
rect -8726 255134 592650 255218
rect -8726 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 73826 255134
rect 74062 254898 74146 255134
rect 74382 254898 109826 255134
rect 110062 254898 110146 255134
rect 110382 254898 124250 255134
rect 124486 254898 154970 255134
rect 155206 254898 185690 255134
rect 185926 254898 217826 255134
rect 218062 254898 218146 255134
rect 218382 254898 253826 255134
rect 254062 254898 254146 255134
rect 254382 254898 289826 255134
rect 290062 254898 290146 255134
rect 290382 254898 325826 255134
rect 326062 254898 326146 255134
rect 326382 254898 361826 255134
rect 362062 254898 362146 255134
rect 362382 254898 397826 255134
rect 398062 254898 398146 255134
rect 398382 254898 433826 255134
rect 434062 254898 434146 255134
rect 434382 254898 469826 255134
rect 470062 254898 470146 255134
rect 470382 254898 505826 255134
rect 506062 254898 506146 255134
rect 506382 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 592650 255134
rect -8726 254866 592650 254898
rect -8726 250954 592650 250986
rect -8726 250718 -8694 250954
rect -8458 250718 -8374 250954
rect -8138 250718 33326 250954
rect 33562 250718 33646 250954
rect 33882 250718 69326 250954
rect 69562 250718 69646 250954
rect 69882 250718 105326 250954
rect 105562 250718 105646 250954
rect 105882 250718 213326 250954
rect 213562 250718 213646 250954
rect 213882 250718 249326 250954
rect 249562 250718 249646 250954
rect 249882 250718 285326 250954
rect 285562 250718 285646 250954
rect 285882 250718 321326 250954
rect 321562 250718 321646 250954
rect 321882 250718 357326 250954
rect 357562 250718 357646 250954
rect 357882 250718 393326 250954
rect 393562 250718 393646 250954
rect 393882 250718 429326 250954
rect 429562 250718 429646 250954
rect 429882 250718 465326 250954
rect 465562 250718 465646 250954
rect 465882 250718 501326 250954
rect 501562 250718 501646 250954
rect 501882 250718 537326 250954
rect 537562 250718 537646 250954
rect 537882 250718 573326 250954
rect 573562 250718 573646 250954
rect 573882 250718 592062 250954
rect 592298 250718 592382 250954
rect 592618 250718 592650 250954
rect -8726 250634 592650 250718
rect -8726 250398 -8694 250634
rect -8458 250398 -8374 250634
rect -8138 250398 33326 250634
rect 33562 250398 33646 250634
rect 33882 250398 69326 250634
rect 69562 250398 69646 250634
rect 69882 250398 105326 250634
rect 105562 250398 105646 250634
rect 105882 250398 213326 250634
rect 213562 250398 213646 250634
rect 213882 250398 249326 250634
rect 249562 250398 249646 250634
rect 249882 250398 285326 250634
rect 285562 250398 285646 250634
rect 285882 250398 321326 250634
rect 321562 250398 321646 250634
rect 321882 250398 357326 250634
rect 357562 250398 357646 250634
rect 357882 250398 393326 250634
rect 393562 250398 393646 250634
rect 393882 250398 429326 250634
rect 429562 250398 429646 250634
rect 429882 250398 465326 250634
rect 465562 250398 465646 250634
rect 465882 250398 501326 250634
rect 501562 250398 501646 250634
rect 501882 250398 537326 250634
rect 537562 250398 537646 250634
rect 537882 250398 573326 250634
rect 573562 250398 573646 250634
rect 573882 250398 592062 250634
rect 592298 250398 592382 250634
rect 592618 250398 592650 250634
rect -8726 250366 592650 250398
rect -8726 246454 592650 246486
rect -8726 246218 -7734 246454
rect -7498 246218 -7414 246454
rect -7178 246218 28826 246454
rect 29062 246218 29146 246454
rect 29382 246218 64826 246454
rect 65062 246218 65146 246454
rect 65382 246218 100826 246454
rect 101062 246218 101146 246454
rect 101382 246218 208826 246454
rect 209062 246218 209146 246454
rect 209382 246218 244826 246454
rect 245062 246218 245146 246454
rect 245382 246218 280826 246454
rect 281062 246218 281146 246454
rect 281382 246218 316826 246454
rect 317062 246218 317146 246454
rect 317382 246218 352826 246454
rect 353062 246218 353146 246454
rect 353382 246218 388826 246454
rect 389062 246218 389146 246454
rect 389382 246218 424826 246454
rect 425062 246218 425146 246454
rect 425382 246218 460826 246454
rect 461062 246218 461146 246454
rect 461382 246218 496826 246454
rect 497062 246218 497146 246454
rect 497382 246218 532826 246454
rect 533062 246218 533146 246454
rect 533382 246218 568826 246454
rect 569062 246218 569146 246454
rect 569382 246218 591102 246454
rect 591338 246218 591422 246454
rect 591658 246218 592650 246454
rect -8726 246134 592650 246218
rect -8726 245898 -7734 246134
rect -7498 245898 -7414 246134
rect -7178 245898 28826 246134
rect 29062 245898 29146 246134
rect 29382 245898 64826 246134
rect 65062 245898 65146 246134
rect 65382 245898 100826 246134
rect 101062 245898 101146 246134
rect 101382 245898 208826 246134
rect 209062 245898 209146 246134
rect 209382 245898 244826 246134
rect 245062 245898 245146 246134
rect 245382 245898 280826 246134
rect 281062 245898 281146 246134
rect 281382 245898 316826 246134
rect 317062 245898 317146 246134
rect 317382 245898 352826 246134
rect 353062 245898 353146 246134
rect 353382 245898 388826 246134
rect 389062 245898 389146 246134
rect 389382 245898 424826 246134
rect 425062 245898 425146 246134
rect 425382 245898 460826 246134
rect 461062 245898 461146 246134
rect 461382 245898 496826 246134
rect 497062 245898 497146 246134
rect 497382 245898 532826 246134
rect 533062 245898 533146 246134
rect 533382 245898 568826 246134
rect 569062 245898 569146 246134
rect 569382 245898 591102 246134
rect 591338 245898 591422 246134
rect 591658 245898 592650 246134
rect -8726 245866 592650 245898
rect -8726 241954 592650 241986
rect -8726 241718 -6774 241954
rect -6538 241718 -6454 241954
rect -6218 241718 24326 241954
rect 24562 241718 24646 241954
rect 24882 241718 60326 241954
rect 60562 241718 60646 241954
rect 60882 241718 96326 241954
rect 96562 241718 96646 241954
rect 96882 241718 204326 241954
rect 204562 241718 204646 241954
rect 204882 241718 240326 241954
rect 240562 241718 240646 241954
rect 240882 241718 276326 241954
rect 276562 241718 276646 241954
rect 276882 241718 312326 241954
rect 312562 241718 312646 241954
rect 312882 241718 348326 241954
rect 348562 241718 348646 241954
rect 348882 241718 384326 241954
rect 384562 241718 384646 241954
rect 384882 241718 420326 241954
rect 420562 241718 420646 241954
rect 420882 241718 456326 241954
rect 456562 241718 456646 241954
rect 456882 241718 492326 241954
rect 492562 241718 492646 241954
rect 492882 241718 528326 241954
rect 528562 241718 528646 241954
rect 528882 241718 564326 241954
rect 564562 241718 564646 241954
rect 564882 241718 590142 241954
rect 590378 241718 590462 241954
rect 590698 241718 592650 241954
rect -8726 241634 592650 241718
rect -8726 241398 -6774 241634
rect -6538 241398 -6454 241634
rect -6218 241398 24326 241634
rect 24562 241398 24646 241634
rect 24882 241398 60326 241634
rect 60562 241398 60646 241634
rect 60882 241398 96326 241634
rect 96562 241398 96646 241634
rect 96882 241398 204326 241634
rect 204562 241398 204646 241634
rect 204882 241398 240326 241634
rect 240562 241398 240646 241634
rect 240882 241398 276326 241634
rect 276562 241398 276646 241634
rect 276882 241398 312326 241634
rect 312562 241398 312646 241634
rect 312882 241398 348326 241634
rect 348562 241398 348646 241634
rect 348882 241398 384326 241634
rect 384562 241398 384646 241634
rect 384882 241398 420326 241634
rect 420562 241398 420646 241634
rect 420882 241398 456326 241634
rect 456562 241398 456646 241634
rect 456882 241398 492326 241634
rect 492562 241398 492646 241634
rect 492882 241398 528326 241634
rect 528562 241398 528646 241634
rect 528882 241398 564326 241634
rect 564562 241398 564646 241634
rect 564882 241398 590142 241634
rect 590378 241398 590462 241634
rect 590698 241398 592650 241634
rect -8726 241366 592650 241398
rect -8726 237454 592650 237486
rect -8726 237218 -5814 237454
rect -5578 237218 -5494 237454
rect -5258 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 55826 237454
rect 56062 237218 56146 237454
rect 56382 237218 91826 237454
rect 92062 237218 92146 237454
rect 92382 237218 199826 237454
rect 200062 237218 200146 237454
rect 200382 237218 235826 237454
rect 236062 237218 236146 237454
rect 236382 237218 271826 237454
rect 272062 237218 272146 237454
rect 272382 237218 307826 237454
rect 308062 237218 308146 237454
rect 308382 237218 343826 237454
rect 344062 237218 344146 237454
rect 344382 237218 379826 237454
rect 380062 237218 380146 237454
rect 380382 237218 415826 237454
rect 416062 237218 416146 237454
rect 416382 237218 451826 237454
rect 452062 237218 452146 237454
rect 452382 237218 487826 237454
rect 488062 237218 488146 237454
rect 488382 237218 523826 237454
rect 524062 237218 524146 237454
rect 524382 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 589182 237454
rect 589418 237218 589502 237454
rect 589738 237218 592650 237454
rect -8726 237134 592650 237218
rect -8726 236898 -5814 237134
rect -5578 236898 -5494 237134
rect -5258 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 55826 237134
rect 56062 236898 56146 237134
rect 56382 236898 91826 237134
rect 92062 236898 92146 237134
rect 92382 236898 199826 237134
rect 200062 236898 200146 237134
rect 200382 236898 235826 237134
rect 236062 236898 236146 237134
rect 236382 236898 271826 237134
rect 272062 236898 272146 237134
rect 272382 236898 307826 237134
rect 308062 236898 308146 237134
rect 308382 236898 343826 237134
rect 344062 236898 344146 237134
rect 344382 236898 379826 237134
rect 380062 236898 380146 237134
rect 380382 236898 415826 237134
rect 416062 236898 416146 237134
rect 416382 236898 451826 237134
rect 452062 236898 452146 237134
rect 452382 236898 487826 237134
rect 488062 236898 488146 237134
rect 488382 236898 523826 237134
rect 524062 236898 524146 237134
rect 524382 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 589182 237134
rect 589418 236898 589502 237134
rect 589738 236898 592650 237134
rect -8726 236866 592650 236898
rect -8726 232954 592650 232986
rect -8726 232718 -4854 232954
rect -4618 232718 -4534 232954
rect -4298 232718 15326 232954
rect 15562 232718 15646 232954
rect 15882 232718 51326 232954
rect 51562 232718 51646 232954
rect 51882 232718 87326 232954
rect 87562 232718 87646 232954
rect 87882 232718 195326 232954
rect 195562 232718 195646 232954
rect 195882 232718 231326 232954
rect 231562 232718 231646 232954
rect 231882 232718 267326 232954
rect 267562 232718 267646 232954
rect 267882 232718 303326 232954
rect 303562 232718 303646 232954
rect 303882 232718 339326 232954
rect 339562 232718 339646 232954
rect 339882 232718 375326 232954
rect 375562 232718 375646 232954
rect 375882 232718 411326 232954
rect 411562 232718 411646 232954
rect 411882 232718 447326 232954
rect 447562 232718 447646 232954
rect 447882 232718 483326 232954
rect 483562 232718 483646 232954
rect 483882 232718 519326 232954
rect 519562 232718 519646 232954
rect 519882 232718 555326 232954
rect 555562 232718 555646 232954
rect 555882 232718 588222 232954
rect 588458 232718 588542 232954
rect 588778 232718 592650 232954
rect -8726 232634 592650 232718
rect -8726 232398 -4854 232634
rect -4618 232398 -4534 232634
rect -4298 232398 15326 232634
rect 15562 232398 15646 232634
rect 15882 232398 51326 232634
rect 51562 232398 51646 232634
rect 51882 232398 87326 232634
rect 87562 232398 87646 232634
rect 87882 232398 195326 232634
rect 195562 232398 195646 232634
rect 195882 232398 231326 232634
rect 231562 232398 231646 232634
rect 231882 232398 267326 232634
rect 267562 232398 267646 232634
rect 267882 232398 303326 232634
rect 303562 232398 303646 232634
rect 303882 232398 339326 232634
rect 339562 232398 339646 232634
rect 339882 232398 375326 232634
rect 375562 232398 375646 232634
rect 375882 232398 411326 232634
rect 411562 232398 411646 232634
rect 411882 232398 447326 232634
rect 447562 232398 447646 232634
rect 447882 232398 483326 232634
rect 483562 232398 483646 232634
rect 483882 232398 519326 232634
rect 519562 232398 519646 232634
rect 519882 232398 555326 232634
rect 555562 232398 555646 232634
rect 555882 232398 588222 232634
rect 588458 232398 588542 232634
rect 588778 232398 592650 232634
rect -8726 232366 592650 232398
rect -8726 228454 592650 228486
rect -8726 228218 -3894 228454
rect -3658 228218 -3574 228454
rect -3338 228218 10826 228454
rect 11062 228218 11146 228454
rect 11382 228218 46826 228454
rect 47062 228218 47146 228454
rect 47382 228218 82826 228454
rect 83062 228218 83146 228454
rect 83382 228218 226826 228454
rect 227062 228218 227146 228454
rect 227382 228218 262826 228454
rect 263062 228218 263146 228454
rect 263382 228218 298826 228454
rect 299062 228218 299146 228454
rect 299382 228218 334826 228454
rect 335062 228218 335146 228454
rect 335382 228218 370826 228454
rect 371062 228218 371146 228454
rect 371382 228218 406826 228454
rect 407062 228218 407146 228454
rect 407382 228218 442826 228454
rect 443062 228218 443146 228454
rect 443382 228218 478826 228454
rect 479062 228218 479146 228454
rect 479382 228218 514826 228454
rect 515062 228218 515146 228454
rect 515382 228218 550826 228454
rect 551062 228218 551146 228454
rect 551382 228218 587262 228454
rect 587498 228218 587582 228454
rect 587818 228218 592650 228454
rect -8726 228134 592650 228218
rect -8726 227898 -3894 228134
rect -3658 227898 -3574 228134
rect -3338 227898 10826 228134
rect 11062 227898 11146 228134
rect 11382 227898 46826 228134
rect 47062 227898 47146 228134
rect 47382 227898 82826 228134
rect 83062 227898 83146 228134
rect 83382 227898 226826 228134
rect 227062 227898 227146 228134
rect 227382 227898 262826 228134
rect 263062 227898 263146 228134
rect 263382 227898 298826 228134
rect 299062 227898 299146 228134
rect 299382 227898 334826 228134
rect 335062 227898 335146 228134
rect 335382 227898 370826 228134
rect 371062 227898 371146 228134
rect 371382 227898 406826 228134
rect 407062 227898 407146 228134
rect 407382 227898 442826 228134
rect 443062 227898 443146 228134
rect 443382 227898 478826 228134
rect 479062 227898 479146 228134
rect 479382 227898 514826 228134
rect 515062 227898 515146 228134
rect 515382 227898 550826 228134
rect 551062 227898 551146 228134
rect 551382 227898 587262 228134
rect 587498 227898 587582 228134
rect 587818 227898 592650 228134
rect -8726 227866 592650 227898
rect -8726 223954 592650 223986
rect -8726 223718 -2934 223954
rect -2698 223718 -2614 223954
rect -2378 223718 6326 223954
rect 6562 223718 6646 223954
rect 6882 223718 42326 223954
rect 42562 223718 42646 223954
rect 42882 223718 78326 223954
rect 78562 223718 78646 223954
rect 78882 223718 114326 223954
rect 114562 223718 114646 223954
rect 114882 223718 139610 223954
rect 139846 223718 170330 223954
rect 170566 223718 222326 223954
rect 222562 223718 222646 223954
rect 222882 223718 258326 223954
rect 258562 223718 258646 223954
rect 258882 223718 294326 223954
rect 294562 223718 294646 223954
rect 294882 223718 330326 223954
rect 330562 223718 330646 223954
rect 330882 223718 366326 223954
rect 366562 223718 366646 223954
rect 366882 223718 402326 223954
rect 402562 223718 402646 223954
rect 402882 223718 438326 223954
rect 438562 223718 438646 223954
rect 438882 223718 474326 223954
rect 474562 223718 474646 223954
rect 474882 223718 510326 223954
rect 510562 223718 510646 223954
rect 510882 223718 546326 223954
rect 546562 223718 546646 223954
rect 546882 223718 582326 223954
rect 582562 223718 582646 223954
rect 582882 223718 586302 223954
rect 586538 223718 586622 223954
rect 586858 223718 592650 223954
rect -8726 223634 592650 223718
rect -8726 223398 -2934 223634
rect -2698 223398 -2614 223634
rect -2378 223398 6326 223634
rect 6562 223398 6646 223634
rect 6882 223398 42326 223634
rect 42562 223398 42646 223634
rect 42882 223398 78326 223634
rect 78562 223398 78646 223634
rect 78882 223398 114326 223634
rect 114562 223398 114646 223634
rect 114882 223398 139610 223634
rect 139846 223398 170330 223634
rect 170566 223398 222326 223634
rect 222562 223398 222646 223634
rect 222882 223398 258326 223634
rect 258562 223398 258646 223634
rect 258882 223398 294326 223634
rect 294562 223398 294646 223634
rect 294882 223398 330326 223634
rect 330562 223398 330646 223634
rect 330882 223398 366326 223634
rect 366562 223398 366646 223634
rect 366882 223398 402326 223634
rect 402562 223398 402646 223634
rect 402882 223398 438326 223634
rect 438562 223398 438646 223634
rect 438882 223398 474326 223634
rect 474562 223398 474646 223634
rect 474882 223398 510326 223634
rect 510562 223398 510646 223634
rect 510882 223398 546326 223634
rect 546562 223398 546646 223634
rect 546882 223398 582326 223634
rect 582562 223398 582646 223634
rect 582882 223398 586302 223634
rect 586538 223398 586622 223634
rect 586858 223398 592650 223634
rect -8726 223366 592650 223398
rect -8726 219454 592650 219486
rect -8726 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 73826 219454
rect 74062 219218 74146 219454
rect 74382 219218 109826 219454
rect 110062 219218 110146 219454
rect 110382 219218 124250 219454
rect 124486 219218 154970 219454
rect 155206 219218 185690 219454
rect 185926 219218 217826 219454
rect 218062 219218 218146 219454
rect 218382 219218 253826 219454
rect 254062 219218 254146 219454
rect 254382 219218 289826 219454
rect 290062 219218 290146 219454
rect 290382 219218 325826 219454
rect 326062 219218 326146 219454
rect 326382 219218 361826 219454
rect 362062 219218 362146 219454
rect 362382 219218 397826 219454
rect 398062 219218 398146 219454
rect 398382 219218 433826 219454
rect 434062 219218 434146 219454
rect 434382 219218 469826 219454
rect 470062 219218 470146 219454
rect 470382 219218 505826 219454
rect 506062 219218 506146 219454
rect 506382 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 592650 219454
rect -8726 219134 592650 219218
rect -8726 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 73826 219134
rect 74062 218898 74146 219134
rect 74382 218898 109826 219134
rect 110062 218898 110146 219134
rect 110382 218898 124250 219134
rect 124486 218898 154970 219134
rect 155206 218898 185690 219134
rect 185926 218898 217826 219134
rect 218062 218898 218146 219134
rect 218382 218898 253826 219134
rect 254062 218898 254146 219134
rect 254382 218898 289826 219134
rect 290062 218898 290146 219134
rect 290382 218898 325826 219134
rect 326062 218898 326146 219134
rect 326382 218898 361826 219134
rect 362062 218898 362146 219134
rect 362382 218898 397826 219134
rect 398062 218898 398146 219134
rect 398382 218898 433826 219134
rect 434062 218898 434146 219134
rect 434382 218898 469826 219134
rect 470062 218898 470146 219134
rect 470382 218898 505826 219134
rect 506062 218898 506146 219134
rect 506382 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 592650 219134
rect -8726 218866 592650 218898
rect -8726 214954 592650 214986
rect -8726 214718 -8694 214954
rect -8458 214718 -8374 214954
rect -8138 214718 33326 214954
rect 33562 214718 33646 214954
rect 33882 214718 69326 214954
rect 69562 214718 69646 214954
rect 69882 214718 105326 214954
rect 105562 214718 105646 214954
rect 105882 214718 213326 214954
rect 213562 214718 213646 214954
rect 213882 214718 249326 214954
rect 249562 214718 249646 214954
rect 249882 214718 285326 214954
rect 285562 214718 285646 214954
rect 285882 214718 321326 214954
rect 321562 214718 321646 214954
rect 321882 214718 357326 214954
rect 357562 214718 357646 214954
rect 357882 214718 393326 214954
rect 393562 214718 393646 214954
rect 393882 214718 429326 214954
rect 429562 214718 429646 214954
rect 429882 214718 465326 214954
rect 465562 214718 465646 214954
rect 465882 214718 501326 214954
rect 501562 214718 501646 214954
rect 501882 214718 537326 214954
rect 537562 214718 537646 214954
rect 537882 214718 573326 214954
rect 573562 214718 573646 214954
rect 573882 214718 592062 214954
rect 592298 214718 592382 214954
rect 592618 214718 592650 214954
rect -8726 214634 592650 214718
rect -8726 214398 -8694 214634
rect -8458 214398 -8374 214634
rect -8138 214398 33326 214634
rect 33562 214398 33646 214634
rect 33882 214398 69326 214634
rect 69562 214398 69646 214634
rect 69882 214398 105326 214634
rect 105562 214398 105646 214634
rect 105882 214398 213326 214634
rect 213562 214398 213646 214634
rect 213882 214398 249326 214634
rect 249562 214398 249646 214634
rect 249882 214398 285326 214634
rect 285562 214398 285646 214634
rect 285882 214398 321326 214634
rect 321562 214398 321646 214634
rect 321882 214398 357326 214634
rect 357562 214398 357646 214634
rect 357882 214398 393326 214634
rect 393562 214398 393646 214634
rect 393882 214398 429326 214634
rect 429562 214398 429646 214634
rect 429882 214398 465326 214634
rect 465562 214398 465646 214634
rect 465882 214398 501326 214634
rect 501562 214398 501646 214634
rect 501882 214398 537326 214634
rect 537562 214398 537646 214634
rect 537882 214398 573326 214634
rect 573562 214398 573646 214634
rect 573882 214398 592062 214634
rect 592298 214398 592382 214634
rect 592618 214398 592650 214634
rect -8726 214366 592650 214398
rect -8726 210454 592650 210486
rect -8726 210218 -7734 210454
rect -7498 210218 -7414 210454
rect -7178 210218 28826 210454
rect 29062 210218 29146 210454
rect 29382 210218 64826 210454
rect 65062 210218 65146 210454
rect 65382 210218 100826 210454
rect 101062 210218 101146 210454
rect 101382 210218 208826 210454
rect 209062 210218 209146 210454
rect 209382 210218 244826 210454
rect 245062 210218 245146 210454
rect 245382 210218 280826 210454
rect 281062 210218 281146 210454
rect 281382 210218 316826 210454
rect 317062 210218 317146 210454
rect 317382 210218 352826 210454
rect 353062 210218 353146 210454
rect 353382 210218 388826 210454
rect 389062 210218 389146 210454
rect 389382 210218 424826 210454
rect 425062 210218 425146 210454
rect 425382 210218 460826 210454
rect 461062 210218 461146 210454
rect 461382 210218 496826 210454
rect 497062 210218 497146 210454
rect 497382 210218 532826 210454
rect 533062 210218 533146 210454
rect 533382 210218 568826 210454
rect 569062 210218 569146 210454
rect 569382 210218 591102 210454
rect 591338 210218 591422 210454
rect 591658 210218 592650 210454
rect -8726 210134 592650 210218
rect -8726 209898 -7734 210134
rect -7498 209898 -7414 210134
rect -7178 209898 28826 210134
rect 29062 209898 29146 210134
rect 29382 209898 64826 210134
rect 65062 209898 65146 210134
rect 65382 209898 100826 210134
rect 101062 209898 101146 210134
rect 101382 209898 208826 210134
rect 209062 209898 209146 210134
rect 209382 209898 244826 210134
rect 245062 209898 245146 210134
rect 245382 209898 280826 210134
rect 281062 209898 281146 210134
rect 281382 209898 316826 210134
rect 317062 209898 317146 210134
rect 317382 209898 352826 210134
rect 353062 209898 353146 210134
rect 353382 209898 388826 210134
rect 389062 209898 389146 210134
rect 389382 209898 424826 210134
rect 425062 209898 425146 210134
rect 425382 209898 460826 210134
rect 461062 209898 461146 210134
rect 461382 209898 496826 210134
rect 497062 209898 497146 210134
rect 497382 209898 532826 210134
rect 533062 209898 533146 210134
rect 533382 209898 568826 210134
rect 569062 209898 569146 210134
rect 569382 209898 591102 210134
rect 591338 209898 591422 210134
rect 591658 209898 592650 210134
rect -8726 209866 592650 209898
rect -8726 205954 592650 205986
rect -8726 205718 -6774 205954
rect -6538 205718 -6454 205954
rect -6218 205718 24326 205954
rect 24562 205718 24646 205954
rect 24882 205718 60326 205954
rect 60562 205718 60646 205954
rect 60882 205718 96326 205954
rect 96562 205718 96646 205954
rect 96882 205718 204326 205954
rect 204562 205718 204646 205954
rect 204882 205718 240326 205954
rect 240562 205718 240646 205954
rect 240882 205718 276326 205954
rect 276562 205718 276646 205954
rect 276882 205718 312326 205954
rect 312562 205718 312646 205954
rect 312882 205718 348326 205954
rect 348562 205718 348646 205954
rect 348882 205718 384326 205954
rect 384562 205718 384646 205954
rect 384882 205718 420326 205954
rect 420562 205718 420646 205954
rect 420882 205718 456326 205954
rect 456562 205718 456646 205954
rect 456882 205718 492326 205954
rect 492562 205718 492646 205954
rect 492882 205718 528326 205954
rect 528562 205718 528646 205954
rect 528882 205718 564326 205954
rect 564562 205718 564646 205954
rect 564882 205718 590142 205954
rect 590378 205718 590462 205954
rect 590698 205718 592650 205954
rect -8726 205634 592650 205718
rect -8726 205398 -6774 205634
rect -6538 205398 -6454 205634
rect -6218 205398 24326 205634
rect 24562 205398 24646 205634
rect 24882 205398 60326 205634
rect 60562 205398 60646 205634
rect 60882 205398 96326 205634
rect 96562 205398 96646 205634
rect 96882 205398 204326 205634
rect 204562 205398 204646 205634
rect 204882 205398 240326 205634
rect 240562 205398 240646 205634
rect 240882 205398 276326 205634
rect 276562 205398 276646 205634
rect 276882 205398 312326 205634
rect 312562 205398 312646 205634
rect 312882 205398 348326 205634
rect 348562 205398 348646 205634
rect 348882 205398 384326 205634
rect 384562 205398 384646 205634
rect 384882 205398 420326 205634
rect 420562 205398 420646 205634
rect 420882 205398 456326 205634
rect 456562 205398 456646 205634
rect 456882 205398 492326 205634
rect 492562 205398 492646 205634
rect 492882 205398 528326 205634
rect 528562 205398 528646 205634
rect 528882 205398 564326 205634
rect 564562 205398 564646 205634
rect 564882 205398 590142 205634
rect 590378 205398 590462 205634
rect 590698 205398 592650 205634
rect -8726 205366 592650 205398
rect -8726 201454 592650 201486
rect -8726 201218 -5814 201454
rect -5578 201218 -5494 201454
rect -5258 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 55826 201454
rect 56062 201218 56146 201454
rect 56382 201218 91826 201454
rect 92062 201218 92146 201454
rect 92382 201218 199826 201454
rect 200062 201218 200146 201454
rect 200382 201218 235826 201454
rect 236062 201218 236146 201454
rect 236382 201218 271826 201454
rect 272062 201218 272146 201454
rect 272382 201218 307826 201454
rect 308062 201218 308146 201454
rect 308382 201218 343826 201454
rect 344062 201218 344146 201454
rect 344382 201218 379826 201454
rect 380062 201218 380146 201454
rect 380382 201218 415826 201454
rect 416062 201218 416146 201454
rect 416382 201218 451826 201454
rect 452062 201218 452146 201454
rect 452382 201218 487826 201454
rect 488062 201218 488146 201454
rect 488382 201218 523826 201454
rect 524062 201218 524146 201454
rect 524382 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 589182 201454
rect 589418 201218 589502 201454
rect 589738 201218 592650 201454
rect -8726 201134 592650 201218
rect -8726 200898 -5814 201134
rect -5578 200898 -5494 201134
rect -5258 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 55826 201134
rect 56062 200898 56146 201134
rect 56382 200898 91826 201134
rect 92062 200898 92146 201134
rect 92382 200898 199826 201134
rect 200062 200898 200146 201134
rect 200382 200898 235826 201134
rect 236062 200898 236146 201134
rect 236382 200898 271826 201134
rect 272062 200898 272146 201134
rect 272382 200898 307826 201134
rect 308062 200898 308146 201134
rect 308382 200898 343826 201134
rect 344062 200898 344146 201134
rect 344382 200898 379826 201134
rect 380062 200898 380146 201134
rect 380382 200898 415826 201134
rect 416062 200898 416146 201134
rect 416382 200898 451826 201134
rect 452062 200898 452146 201134
rect 452382 200898 487826 201134
rect 488062 200898 488146 201134
rect 488382 200898 523826 201134
rect 524062 200898 524146 201134
rect 524382 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 589182 201134
rect 589418 200898 589502 201134
rect 589738 200898 592650 201134
rect -8726 200866 592650 200898
rect -8726 196954 592650 196986
rect -8726 196718 -4854 196954
rect -4618 196718 -4534 196954
rect -4298 196718 15326 196954
rect 15562 196718 15646 196954
rect 15882 196718 51326 196954
rect 51562 196718 51646 196954
rect 51882 196718 87326 196954
rect 87562 196718 87646 196954
rect 87882 196718 123326 196954
rect 123562 196718 123646 196954
rect 123882 196718 159326 196954
rect 159562 196718 159646 196954
rect 159882 196718 195326 196954
rect 195562 196718 195646 196954
rect 195882 196718 231326 196954
rect 231562 196718 231646 196954
rect 231882 196718 267326 196954
rect 267562 196718 267646 196954
rect 267882 196718 303326 196954
rect 303562 196718 303646 196954
rect 303882 196718 339326 196954
rect 339562 196718 339646 196954
rect 339882 196718 375326 196954
rect 375562 196718 375646 196954
rect 375882 196718 411326 196954
rect 411562 196718 411646 196954
rect 411882 196718 447326 196954
rect 447562 196718 447646 196954
rect 447882 196718 483326 196954
rect 483562 196718 483646 196954
rect 483882 196718 519326 196954
rect 519562 196718 519646 196954
rect 519882 196718 555326 196954
rect 555562 196718 555646 196954
rect 555882 196718 588222 196954
rect 588458 196718 588542 196954
rect 588778 196718 592650 196954
rect -8726 196634 592650 196718
rect -8726 196398 -4854 196634
rect -4618 196398 -4534 196634
rect -4298 196398 15326 196634
rect 15562 196398 15646 196634
rect 15882 196398 51326 196634
rect 51562 196398 51646 196634
rect 51882 196398 87326 196634
rect 87562 196398 87646 196634
rect 87882 196398 123326 196634
rect 123562 196398 123646 196634
rect 123882 196398 159326 196634
rect 159562 196398 159646 196634
rect 159882 196398 195326 196634
rect 195562 196398 195646 196634
rect 195882 196398 231326 196634
rect 231562 196398 231646 196634
rect 231882 196398 267326 196634
rect 267562 196398 267646 196634
rect 267882 196398 303326 196634
rect 303562 196398 303646 196634
rect 303882 196398 339326 196634
rect 339562 196398 339646 196634
rect 339882 196398 375326 196634
rect 375562 196398 375646 196634
rect 375882 196398 411326 196634
rect 411562 196398 411646 196634
rect 411882 196398 447326 196634
rect 447562 196398 447646 196634
rect 447882 196398 483326 196634
rect 483562 196398 483646 196634
rect 483882 196398 519326 196634
rect 519562 196398 519646 196634
rect 519882 196398 555326 196634
rect 555562 196398 555646 196634
rect 555882 196398 588222 196634
rect 588458 196398 588542 196634
rect 588778 196398 592650 196634
rect -8726 196366 592650 196398
rect -8726 192454 592650 192486
rect -8726 192218 -3894 192454
rect -3658 192218 -3574 192454
rect -3338 192218 10826 192454
rect 11062 192218 11146 192454
rect 11382 192218 46826 192454
rect 47062 192218 47146 192454
rect 47382 192218 82826 192454
rect 83062 192218 83146 192454
rect 83382 192218 118826 192454
rect 119062 192218 119146 192454
rect 119382 192218 154826 192454
rect 155062 192218 155146 192454
rect 155382 192218 190826 192454
rect 191062 192218 191146 192454
rect 191382 192218 226826 192454
rect 227062 192218 227146 192454
rect 227382 192218 262826 192454
rect 263062 192218 263146 192454
rect 263382 192218 298826 192454
rect 299062 192218 299146 192454
rect 299382 192218 334826 192454
rect 335062 192218 335146 192454
rect 335382 192218 370826 192454
rect 371062 192218 371146 192454
rect 371382 192218 406826 192454
rect 407062 192218 407146 192454
rect 407382 192218 442826 192454
rect 443062 192218 443146 192454
rect 443382 192218 478826 192454
rect 479062 192218 479146 192454
rect 479382 192218 514826 192454
rect 515062 192218 515146 192454
rect 515382 192218 550826 192454
rect 551062 192218 551146 192454
rect 551382 192218 587262 192454
rect 587498 192218 587582 192454
rect 587818 192218 592650 192454
rect -8726 192134 592650 192218
rect -8726 191898 -3894 192134
rect -3658 191898 -3574 192134
rect -3338 191898 10826 192134
rect 11062 191898 11146 192134
rect 11382 191898 46826 192134
rect 47062 191898 47146 192134
rect 47382 191898 82826 192134
rect 83062 191898 83146 192134
rect 83382 191898 118826 192134
rect 119062 191898 119146 192134
rect 119382 191898 154826 192134
rect 155062 191898 155146 192134
rect 155382 191898 190826 192134
rect 191062 191898 191146 192134
rect 191382 191898 226826 192134
rect 227062 191898 227146 192134
rect 227382 191898 262826 192134
rect 263062 191898 263146 192134
rect 263382 191898 298826 192134
rect 299062 191898 299146 192134
rect 299382 191898 334826 192134
rect 335062 191898 335146 192134
rect 335382 191898 370826 192134
rect 371062 191898 371146 192134
rect 371382 191898 406826 192134
rect 407062 191898 407146 192134
rect 407382 191898 442826 192134
rect 443062 191898 443146 192134
rect 443382 191898 478826 192134
rect 479062 191898 479146 192134
rect 479382 191898 514826 192134
rect 515062 191898 515146 192134
rect 515382 191898 550826 192134
rect 551062 191898 551146 192134
rect 551382 191898 587262 192134
rect 587498 191898 587582 192134
rect 587818 191898 592650 192134
rect -8726 191866 592650 191898
rect -8726 187954 592650 187986
rect -8726 187718 -2934 187954
rect -2698 187718 -2614 187954
rect -2378 187718 6326 187954
rect 6562 187718 6646 187954
rect 6882 187718 42326 187954
rect 42562 187718 42646 187954
rect 42882 187718 78326 187954
rect 78562 187718 78646 187954
rect 78882 187718 114326 187954
rect 114562 187718 114646 187954
rect 114882 187718 150326 187954
rect 150562 187718 150646 187954
rect 150882 187718 186326 187954
rect 186562 187718 186646 187954
rect 186882 187718 222326 187954
rect 222562 187718 222646 187954
rect 222882 187718 258326 187954
rect 258562 187718 258646 187954
rect 258882 187718 294326 187954
rect 294562 187718 294646 187954
rect 294882 187718 330326 187954
rect 330562 187718 330646 187954
rect 330882 187718 366326 187954
rect 366562 187718 366646 187954
rect 366882 187718 402326 187954
rect 402562 187718 402646 187954
rect 402882 187718 438326 187954
rect 438562 187718 438646 187954
rect 438882 187718 474326 187954
rect 474562 187718 474646 187954
rect 474882 187718 510326 187954
rect 510562 187718 510646 187954
rect 510882 187718 546326 187954
rect 546562 187718 546646 187954
rect 546882 187718 582326 187954
rect 582562 187718 582646 187954
rect 582882 187718 586302 187954
rect 586538 187718 586622 187954
rect 586858 187718 592650 187954
rect -8726 187634 592650 187718
rect -8726 187398 -2934 187634
rect -2698 187398 -2614 187634
rect -2378 187398 6326 187634
rect 6562 187398 6646 187634
rect 6882 187398 42326 187634
rect 42562 187398 42646 187634
rect 42882 187398 78326 187634
rect 78562 187398 78646 187634
rect 78882 187398 114326 187634
rect 114562 187398 114646 187634
rect 114882 187398 150326 187634
rect 150562 187398 150646 187634
rect 150882 187398 186326 187634
rect 186562 187398 186646 187634
rect 186882 187398 222326 187634
rect 222562 187398 222646 187634
rect 222882 187398 258326 187634
rect 258562 187398 258646 187634
rect 258882 187398 294326 187634
rect 294562 187398 294646 187634
rect 294882 187398 330326 187634
rect 330562 187398 330646 187634
rect 330882 187398 366326 187634
rect 366562 187398 366646 187634
rect 366882 187398 402326 187634
rect 402562 187398 402646 187634
rect 402882 187398 438326 187634
rect 438562 187398 438646 187634
rect 438882 187398 474326 187634
rect 474562 187398 474646 187634
rect 474882 187398 510326 187634
rect 510562 187398 510646 187634
rect 510882 187398 546326 187634
rect 546562 187398 546646 187634
rect 546882 187398 582326 187634
rect 582562 187398 582646 187634
rect 582882 187398 586302 187634
rect 586538 187398 586622 187634
rect 586858 187398 592650 187634
rect -8726 187366 592650 187398
rect -8726 183454 592650 183486
rect -8726 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 73826 183454
rect 74062 183218 74146 183454
rect 74382 183218 109826 183454
rect 110062 183218 110146 183454
rect 110382 183218 145826 183454
rect 146062 183218 146146 183454
rect 146382 183218 181826 183454
rect 182062 183218 182146 183454
rect 182382 183218 217826 183454
rect 218062 183218 218146 183454
rect 218382 183218 253826 183454
rect 254062 183218 254146 183454
rect 254382 183218 289826 183454
rect 290062 183218 290146 183454
rect 290382 183218 325826 183454
rect 326062 183218 326146 183454
rect 326382 183218 361826 183454
rect 362062 183218 362146 183454
rect 362382 183218 397826 183454
rect 398062 183218 398146 183454
rect 398382 183218 433826 183454
rect 434062 183218 434146 183454
rect 434382 183218 469826 183454
rect 470062 183218 470146 183454
rect 470382 183218 505826 183454
rect 506062 183218 506146 183454
rect 506382 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 592650 183454
rect -8726 183134 592650 183218
rect -8726 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 73826 183134
rect 74062 182898 74146 183134
rect 74382 182898 109826 183134
rect 110062 182898 110146 183134
rect 110382 182898 145826 183134
rect 146062 182898 146146 183134
rect 146382 182898 181826 183134
rect 182062 182898 182146 183134
rect 182382 182898 217826 183134
rect 218062 182898 218146 183134
rect 218382 182898 253826 183134
rect 254062 182898 254146 183134
rect 254382 182898 289826 183134
rect 290062 182898 290146 183134
rect 290382 182898 325826 183134
rect 326062 182898 326146 183134
rect 326382 182898 361826 183134
rect 362062 182898 362146 183134
rect 362382 182898 397826 183134
rect 398062 182898 398146 183134
rect 398382 182898 433826 183134
rect 434062 182898 434146 183134
rect 434382 182898 469826 183134
rect 470062 182898 470146 183134
rect 470382 182898 505826 183134
rect 506062 182898 506146 183134
rect 506382 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 592650 183134
rect -8726 182866 592650 182898
rect -8726 178954 592650 178986
rect -8726 178718 -8694 178954
rect -8458 178718 -8374 178954
rect -8138 178718 33326 178954
rect 33562 178718 33646 178954
rect 33882 178718 69326 178954
rect 69562 178718 69646 178954
rect 69882 178718 105326 178954
rect 105562 178718 105646 178954
rect 105882 178718 141326 178954
rect 141562 178718 141646 178954
rect 141882 178718 177326 178954
rect 177562 178718 177646 178954
rect 177882 178718 213326 178954
rect 213562 178718 213646 178954
rect 213882 178718 249326 178954
rect 249562 178718 249646 178954
rect 249882 178718 285326 178954
rect 285562 178718 285646 178954
rect 285882 178718 321326 178954
rect 321562 178718 321646 178954
rect 321882 178718 357326 178954
rect 357562 178718 357646 178954
rect 357882 178718 393326 178954
rect 393562 178718 393646 178954
rect 393882 178718 429326 178954
rect 429562 178718 429646 178954
rect 429882 178718 465326 178954
rect 465562 178718 465646 178954
rect 465882 178718 501326 178954
rect 501562 178718 501646 178954
rect 501882 178718 537326 178954
rect 537562 178718 537646 178954
rect 537882 178718 573326 178954
rect 573562 178718 573646 178954
rect 573882 178718 592062 178954
rect 592298 178718 592382 178954
rect 592618 178718 592650 178954
rect -8726 178634 592650 178718
rect -8726 178398 -8694 178634
rect -8458 178398 -8374 178634
rect -8138 178398 33326 178634
rect 33562 178398 33646 178634
rect 33882 178398 69326 178634
rect 69562 178398 69646 178634
rect 69882 178398 105326 178634
rect 105562 178398 105646 178634
rect 105882 178398 141326 178634
rect 141562 178398 141646 178634
rect 141882 178398 177326 178634
rect 177562 178398 177646 178634
rect 177882 178398 213326 178634
rect 213562 178398 213646 178634
rect 213882 178398 249326 178634
rect 249562 178398 249646 178634
rect 249882 178398 285326 178634
rect 285562 178398 285646 178634
rect 285882 178398 321326 178634
rect 321562 178398 321646 178634
rect 321882 178398 357326 178634
rect 357562 178398 357646 178634
rect 357882 178398 393326 178634
rect 393562 178398 393646 178634
rect 393882 178398 429326 178634
rect 429562 178398 429646 178634
rect 429882 178398 465326 178634
rect 465562 178398 465646 178634
rect 465882 178398 501326 178634
rect 501562 178398 501646 178634
rect 501882 178398 537326 178634
rect 537562 178398 537646 178634
rect 537882 178398 573326 178634
rect 573562 178398 573646 178634
rect 573882 178398 592062 178634
rect 592298 178398 592382 178634
rect 592618 178398 592650 178634
rect -8726 178366 592650 178398
rect -8726 174454 592650 174486
rect -8726 174218 -7734 174454
rect -7498 174218 -7414 174454
rect -7178 174218 28826 174454
rect 29062 174218 29146 174454
rect 29382 174218 64826 174454
rect 65062 174218 65146 174454
rect 65382 174218 100826 174454
rect 101062 174218 101146 174454
rect 101382 174218 208826 174454
rect 209062 174218 209146 174454
rect 209382 174218 244826 174454
rect 245062 174218 245146 174454
rect 245382 174218 280826 174454
rect 281062 174218 281146 174454
rect 281382 174218 316826 174454
rect 317062 174218 317146 174454
rect 317382 174218 352826 174454
rect 353062 174218 353146 174454
rect 353382 174218 388826 174454
rect 389062 174218 389146 174454
rect 389382 174218 424826 174454
rect 425062 174218 425146 174454
rect 425382 174218 460826 174454
rect 461062 174218 461146 174454
rect 461382 174218 496826 174454
rect 497062 174218 497146 174454
rect 497382 174218 532826 174454
rect 533062 174218 533146 174454
rect 533382 174218 568826 174454
rect 569062 174218 569146 174454
rect 569382 174218 591102 174454
rect 591338 174218 591422 174454
rect 591658 174218 592650 174454
rect -8726 174134 592650 174218
rect -8726 173898 -7734 174134
rect -7498 173898 -7414 174134
rect -7178 173898 28826 174134
rect 29062 173898 29146 174134
rect 29382 173898 64826 174134
rect 65062 173898 65146 174134
rect 65382 173898 100826 174134
rect 101062 173898 101146 174134
rect 101382 173898 208826 174134
rect 209062 173898 209146 174134
rect 209382 173898 244826 174134
rect 245062 173898 245146 174134
rect 245382 173898 280826 174134
rect 281062 173898 281146 174134
rect 281382 173898 316826 174134
rect 317062 173898 317146 174134
rect 317382 173898 352826 174134
rect 353062 173898 353146 174134
rect 353382 173898 388826 174134
rect 389062 173898 389146 174134
rect 389382 173898 424826 174134
rect 425062 173898 425146 174134
rect 425382 173898 460826 174134
rect 461062 173898 461146 174134
rect 461382 173898 496826 174134
rect 497062 173898 497146 174134
rect 497382 173898 532826 174134
rect 533062 173898 533146 174134
rect 533382 173898 568826 174134
rect 569062 173898 569146 174134
rect 569382 173898 591102 174134
rect 591338 173898 591422 174134
rect 591658 173898 592650 174134
rect -8726 173866 592650 173898
rect -8726 169954 592650 169986
rect -8726 169718 -6774 169954
rect -6538 169718 -6454 169954
rect -6218 169718 24326 169954
rect 24562 169718 24646 169954
rect 24882 169718 60326 169954
rect 60562 169718 60646 169954
rect 60882 169718 96326 169954
rect 96562 169718 96646 169954
rect 96882 169718 204326 169954
rect 204562 169718 204646 169954
rect 204882 169718 240326 169954
rect 240562 169718 240646 169954
rect 240882 169718 276326 169954
rect 276562 169718 276646 169954
rect 276882 169718 312326 169954
rect 312562 169718 312646 169954
rect 312882 169718 348326 169954
rect 348562 169718 348646 169954
rect 348882 169718 384326 169954
rect 384562 169718 384646 169954
rect 384882 169718 420326 169954
rect 420562 169718 420646 169954
rect 420882 169718 456326 169954
rect 456562 169718 456646 169954
rect 456882 169718 492326 169954
rect 492562 169718 492646 169954
rect 492882 169718 528326 169954
rect 528562 169718 528646 169954
rect 528882 169718 564326 169954
rect 564562 169718 564646 169954
rect 564882 169718 590142 169954
rect 590378 169718 590462 169954
rect 590698 169718 592650 169954
rect -8726 169634 592650 169718
rect -8726 169398 -6774 169634
rect -6538 169398 -6454 169634
rect -6218 169398 24326 169634
rect 24562 169398 24646 169634
rect 24882 169398 60326 169634
rect 60562 169398 60646 169634
rect 60882 169398 96326 169634
rect 96562 169398 96646 169634
rect 96882 169398 204326 169634
rect 204562 169398 204646 169634
rect 204882 169398 240326 169634
rect 240562 169398 240646 169634
rect 240882 169398 276326 169634
rect 276562 169398 276646 169634
rect 276882 169398 312326 169634
rect 312562 169398 312646 169634
rect 312882 169398 348326 169634
rect 348562 169398 348646 169634
rect 348882 169398 384326 169634
rect 384562 169398 384646 169634
rect 384882 169398 420326 169634
rect 420562 169398 420646 169634
rect 420882 169398 456326 169634
rect 456562 169398 456646 169634
rect 456882 169398 492326 169634
rect 492562 169398 492646 169634
rect 492882 169398 528326 169634
rect 528562 169398 528646 169634
rect 528882 169398 564326 169634
rect 564562 169398 564646 169634
rect 564882 169398 590142 169634
rect 590378 169398 590462 169634
rect 590698 169398 592650 169634
rect -8726 169366 592650 169398
rect -8726 165454 592650 165486
rect -8726 165218 -5814 165454
rect -5578 165218 -5494 165454
rect -5258 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 55826 165454
rect 56062 165218 56146 165454
rect 56382 165218 91826 165454
rect 92062 165218 92146 165454
rect 92382 165218 199826 165454
rect 200062 165218 200146 165454
rect 200382 165218 235826 165454
rect 236062 165218 236146 165454
rect 236382 165218 271826 165454
rect 272062 165218 272146 165454
rect 272382 165218 307826 165454
rect 308062 165218 308146 165454
rect 308382 165218 343826 165454
rect 344062 165218 344146 165454
rect 344382 165218 379826 165454
rect 380062 165218 380146 165454
rect 380382 165218 415826 165454
rect 416062 165218 416146 165454
rect 416382 165218 451826 165454
rect 452062 165218 452146 165454
rect 452382 165218 487826 165454
rect 488062 165218 488146 165454
rect 488382 165218 523826 165454
rect 524062 165218 524146 165454
rect 524382 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 589182 165454
rect 589418 165218 589502 165454
rect 589738 165218 592650 165454
rect -8726 165134 592650 165218
rect -8726 164898 -5814 165134
rect -5578 164898 -5494 165134
rect -5258 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 55826 165134
rect 56062 164898 56146 165134
rect 56382 164898 91826 165134
rect 92062 164898 92146 165134
rect 92382 164898 199826 165134
rect 200062 164898 200146 165134
rect 200382 164898 235826 165134
rect 236062 164898 236146 165134
rect 236382 164898 271826 165134
rect 272062 164898 272146 165134
rect 272382 164898 307826 165134
rect 308062 164898 308146 165134
rect 308382 164898 343826 165134
rect 344062 164898 344146 165134
rect 344382 164898 379826 165134
rect 380062 164898 380146 165134
rect 380382 164898 415826 165134
rect 416062 164898 416146 165134
rect 416382 164898 451826 165134
rect 452062 164898 452146 165134
rect 452382 164898 487826 165134
rect 488062 164898 488146 165134
rect 488382 164898 523826 165134
rect 524062 164898 524146 165134
rect 524382 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 589182 165134
rect 589418 164898 589502 165134
rect 589738 164898 592650 165134
rect -8726 164866 592650 164898
rect -8726 160954 592650 160986
rect -8726 160718 -4854 160954
rect -4618 160718 -4534 160954
rect -4298 160718 15326 160954
rect 15562 160718 15646 160954
rect 15882 160718 51326 160954
rect 51562 160718 51646 160954
rect 51882 160718 87326 160954
rect 87562 160718 87646 160954
rect 87882 160718 123326 160954
rect 123562 160718 123646 160954
rect 123882 160718 159326 160954
rect 159562 160718 159646 160954
rect 159882 160718 195326 160954
rect 195562 160718 195646 160954
rect 195882 160718 231326 160954
rect 231562 160718 231646 160954
rect 231882 160718 267326 160954
rect 267562 160718 267646 160954
rect 267882 160718 303326 160954
rect 303562 160718 303646 160954
rect 303882 160718 339326 160954
rect 339562 160718 339646 160954
rect 339882 160718 375326 160954
rect 375562 160718 375646 160954
rect 375882 160718 411326 160954
rect 411562 160718 411646 160954
rect 411882 160718 447326 160954
rect 447562 160718 447646 160954
rect 447882 160718 483326 160954
rect 483562 160718 483646 160954
rect 483882 160718 519326 160954
rect 519562 160718 519646 160954
rect 519882 160718 555326 160954
rect 555562 160718 555646 160954
rect 555882 160718 588222 160954
rect 588458 160718 588542 160954
rect 588778 160718 592650 160954
rect -8726 160634 592650 160718
rect -8726 160398 -4854 160634
rect -4618 160398 -4534 160634
rect -4298 160398 15326 160634
rect 15562 160398 15646 160634
rect 15882 160398 51326 160634
rect 51562 160398 51646 160634
rect 51882 160398 87326 160634
rect 87562 160398 87646 160634
rect 87882 160398 123326 160634
rect 123562 160398 123646 160634
rect 123882 160398 159326 160634
rect 159562 160398 159646 160634
rect 159882 160398 195326 160634
rect 195562 160398 195646 160634
rect 195882 160398 231326 160634
rect 231562 160398 231646 160634
rect 231882 160398 267326 160634
rect 267562 160398 267646 160634
rect 267882 160398 303326 160634
rect 303562 160398 303646 160634
rect 303882 160398 339326 160634
rect 339562 160398 339646 160634
rect 339882 160398 375326 160634
rect 375562 160398 375646 160634
rect 375882 160398 411326 160634
rect 411562 160398 411646 160634
rect 411882 160398 447326 160634
rect 447562 160398 447646 160634
rect 447882 160398 483326 160634
rect 483562 160398 483646 160634
rect 483882 160398 519326 160634
rect 519562 160398 519646 160634
rect 519882 160398 555326 160634
rect 555562 160398 555646 160634
rect 555882 160398 588222 160634
rect 588458 160398 588542 160634
rect 588778 160398 592650 160634
rect -8726 160366 592650 160398
rect -8726 156454 592650 156486
rect -8726 156218 -3894 156454
rect -3658 156218 -3574 156454
rect -3338 156218 10826 156454
rect 11062 156218 11146 156454
rect 11382 156218 46826 156454
rect 47062 156218 47146 156454
rect 47382 156218 82826 156454
rect 83062 156218 83146 156454
rect 83382 156218 118826 156454
rect 119062 156218 119146 156454
rect 119382 156218 154826 156454
rect 155062 156218 155146 156454
rect 155382 156218 190826 156454
rect 191062 156218 191146 156454
rect 191382 156218 226826 156454
rect 227062 156218 227146 156454
rect 227382 156218 262826 156454
rect 263062 156218 263146 156454
rect 263382 156218 298826 156454
rect 299062 156218 299146 156454
rect 299382 156218 334826 156454
rect 335062 156218 335146 156454
rect 335382 156218 370826 156454
rect 371062 156218 371146 156454
rect 371382 156218 406826 156454
rect 407062 156218 407146 156454
rect 407382 156218 442826 156454
rect 443062 156218 443146 156454
rect 443382 156218 478826 156454
rect 479062 156218 479146 156454
rect 479382 156218 514826 156454
rect 515062 156218 515146 156454
rect 515382 156218 550826 156454
rect 551062 156218 551146 156454
rect 551382 156218 587262 156454
rect 587498 156218 587582 156454
rect 587818 156218 592650 156454
rect -8726 156134 592650 156218
rect -8726 155898 -3894 156134
rect -3658 155898 -3574 156134
rect -3338 155898 10826 156134
rect 11062 155898 11146 156134
rect 11382 155898 46826 156134
rect 47062 155898 47146 156134
rect 47382 155898 82826 156134
rect 83062 155898 83146 156134
rect 83382 155898 118826 156134
rect 119062 155898 119146 156134
rect 119382 155898 154826 156134
rect 155062 155898 155146 156134
rect 155382 155898 190826 156134
rect 191062 155898 191146 156134
rect 191382 155898 226826 156134
rect 227062 155898 227146 156134
rect 227382 155898 262826 156134
rect 263062 155898 263146 156134
rect 263382 155898 298826 156134
rect 299062 155898 299146 156134
rect 299382 155898 334826 156134
rect 335062 155898 335146 156134
rect 335382 155898 370826 156134
rect 371062 155898 371146 156134
rect 371382 155898 406826 156134
rect 407062 155898 407146 156134
rect 407382 155898 442826 156134
rect 443062 155898 443146 156134
rect 443382 155898 478826 156134
rect 479062 155898 479146 156134
rect 479382 155898 514826 156134
rect 515062 155898 515146 156134
rect 515382 155898 550826 156134
rect 551062 155898 551146 156134
rect 551382 155898 587262 156134
rect 587498 155898 587582 156134
rect 587818 155898 592650 156134
rect -8726 155866 592650 155898
rect -8726 151954 592650 151986
rect -8726 151718 -2934 151954
rect -2698 151718 -2614 151954
rect -2378 151718 6326 151954
rect 6562 151718 6646 151954
rect 6882 151718 42326 151954
rect 42562 151718 42646 151954
rect 42882 151718 78326 151954
rect 78562 151718 78646 151954
rect 78882 151718 114326 151954
rect 114562 151718 114646 151954
rect 114882 151718 150326 151954
rect 150562 151718 150646 151954
rect 150882 151718 186326 151954
rect 186562 151718 186646 151954
rect 186882 151718 222326 151954
rect 222562 151718 222646 151954
rect 222882 151718 258326 151954
rect 258562 151718 258646 151954
rect 258882 151718 294326 151954
rect 294562 151718 294646 151954
rect 294882 151718 330326 151954
rect 330562 151718 330646 151954
rect 330882 151718 366326 151954
rect 366562 151718 366646 151954
rect 366882 151718 402326 151954
rect 402562 151718 402646 151954
rect 402882 151718 438326 151954
rect 438562 151718 438646 151954
rect 438882 151718 474326 151954
rect 474562 151718 474646 151954
rect 474882 151718 510326 151954
rect 510562 151718 510646 151954
rect 510882 151718 546326 151954
rect 546562 151718 546646 151954
rect 546882 151718 582326 151954
rect 582562 151718 582646 151954
rect 582882 151718 586302 151954
rect 586538 151718 586622 151954
rect 586858 151718 592650 151954
rect -8726 151634 592650 151718
rect -8726 151398 -2934 151634
rect -2698 151398 -2614 151634
rect -2378 151398 6326 151634
rect 6562 151398 6646 151634
rect 6882 151398 42326 151634
rect 42562 151398 42646 151634
rect 42882 151398 78326 151634
rect 78562 151398 78646 151634
rect 78882 151398 114326 151634
rect 114562 151398 114646 151634
rect 114882 151398 150326 151634
rect 150562 151398 150646 151634
rect 150882 151398 186326 151634
rect 186562 151398 186646 151634
rect 186882 151398 222326 151634
rect 222562 151398 222646 151634
rect 222882 151398 258326 151634
rect 258562 151398 258646 151634
rect 258882 151398 294326 151634
rect 294562 151398 294646 151634
rect 294882 151398 330326 151634
rect 330562 151398 330646 151634
rect 330882 151398 366326 151634
rect 366562 151398 366646 151634
rect 366882 151398 402326 151634
rect 402562 151398 402646 151634
rect 402882 151398 438326 151634
rect 438562 151398 438646 151634
rect 438882 151398 474326 151634
rect 474562 151398 474646 151634
rect 474882 151398 510326 151634
rect 510562 151398 510646 151634
rect 510882 151398 546326 151634
rect 546562 151398 546646 151634
rect 546882 151398 582326 151634
rect 582562 151398 582646 151634
rect 582882 151398 586302 151634
rect 586538 151398 586622 151634
rect 586858 151398 592650 151634
rect -8726 151366 592650 151398
rect -8726 147454 592650 147486
rect -8726 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 73826 147454
rect 74062 147218 74146 147454
rect 74382 147218 109826 147454
rect 110062 147218 110146 147454
rect 110382 147218 145826 147454
rect 146062 147218 146146 147454
rect 146382 147218 181826 147454
rect 182062 147218 182146 147454
rect 182382 147218 217826 147454
rect 218062 147218 218146 147454
rect 218382 147218 253826 147454
rect 254062 147218 254146 147454
rect 254382 147218 289826 147454
rect 290062 147218 290146 147454
rect 290382 147218 325826 147454
rect 326062 147218 326146 147454
rect 326382 147218 361826 147454
rect 362062 147218 362146 147454
rect 362382 147218 397826 147454
rect 398062 147218 398146 147454
rect 398382 147218 433826 147454
rect 434062 147218 434146 147454
rect 434382 147218 469826 147454
rect 470062 147218 470146 147454
rect 470382 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 592650 147454
rect -8726 147134 592650 147218
rect -8726 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 73826 147134
rect 74062 146898 74146 147134
rect 74382 146898 109826 147134
rect 110062 146898 110146 147134
rect 110382 146898 145826 147134
rect 146062 146898 146146 147134
rect 146382 146898 181826 147134
rect 182062 146898 182146 147134
rect 182382 146898 217826 147134
rect 218062 146898 218146 147134
rect 218382 146898 253826 147134
rect 254062 146898 254146 147134
rect 254382 146898 289826 147134
rect 290062 146898 290146 147134
rect 290382 146898 325826 147134
rect 326062 146898 326146 147134
rect 326382 146898 361826 147134
rect 362062 146898 362146 147134
rect 362382 146898 397826 147134
rect 398062 146898 398146 147134
rect 398382 146898 433826 147134
rect 434062 146898 434146 147134
rect 434382 146898 469826 147134
rect 470062 146898 470146 147134
rect 470382 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 592650 147134
rect -8726 146866 592650 146898
rect -8726 142954 592650 142986
rect -8726 142718 -8694 142954
rect -8458 142718 -8374 142954
rect -8138 142718 33326 142954
rect 33562 142718 33646 142954
rect 33882 142718 69326 142954
rect 69562 142718 69646 142954
rect 69882 142718 105326 142954
rect 105562 142718 105646 142954
rect 105882 142718 141326 142954
rect 141562 142718 141646 142954
rect 141882 142718 177326 142954
rect 177562 142718 177646 142954
rect 177882 142718 213326 142954
rect 213562 142718 213646 142954
rect 213882 142718 249326 142954
rect 249562 142718 249646 142954
rect 249882 142718 285326 142954
rect 285562 142718 285646 142954
rect 285882 142718 321326 142954
rect 321562 142718 321646 142954
rect 321882 142718 357326 142954
rect 357562 142718 357646 142954
rect 357882 142718 393326 142954
rect 393562 142718 393646 142954
rect 393882 142718 429326 142954
rect 429562 142718 429646 142954
rect 429882 142718 465326 142954
rect 465562 142718 465646 142954
rect 465882 142718 501326 142954
rect 501562 142718 501646 142954
rect 501882 142718 537326 142954
rect 537562 142718 537646 142954
rect 537882 142718 573326 142954
rect 573562 142718 573646 142954
rect 573882 142718 592062 142954
rect 592298 142718 592382 142954
rect 592618 142718 592650 142954
rect -8726 142634 592650 142718
rect -8726 142398 -8694 142634
rect -8458 142398 -8374 142634
rect -8138 142398 33326 142634
rect 33562 142398 33646 142634
rect 33882 142398 69326 142634
rect 69562 142398 69646 142634
rect 69882 142398 105326 142634
rect 105562 142398 105646 142634
rect 105882 142398 141326 142634
rect 141562 142398 141646 142634
rect 141882 142398 177326 142634
rect 177562 142398 177646 142634
rect 177882 142398 213326 142634
rect 213562 142398 213646 142634
rect 213882 142398 249326 142634
rect 249562 142398 249646 142634
rect 249882 142398 285326 142634
rect 285562 142398 285646 142634
rect 285882 142398 321326 142634
rect 321562 142398 321646 142634
rect 321882 142398 357326 142634
rect 357562 142398 357646 142634
rect 357882 142398 393326 142634
rect 393562 142398 393646 142634
rect 393882 142398 429326 142634
rect 429562 142398 429646 142634
rect 429882 142398 465326 142634
rect 465562 142398 465646 142634
rect 465882 142398 501326 142634
rect 501562 142398 501646 142634
rect 501882 142398 537326 142634
rect 537562 142398 537646 142634
rect 537882 142398 573326 142634
rect 573562 142398 573646 142634
rect 573882 142398 592062 142634
rect 592298 142398 592382 142634
rect 592618 142398 592650 142634
rect -8726 142366 592650 142398
rect -8726 138454 592650 138486
rect -8726 138218 -7734 138454
rect -7498 138218 -7414 138454
rect -7178 138218 28826 138454
rect 29062 138218 29146 138454
rect 29382 138218 64826 138454
rect 65062 138218 65146 138454
rect 65382 138218 100826 138454
rect 101062 138218 101146 138454
rect 101382 138218 208826 138454
rect 209062 138218 209146 138454
rect 209382 138218 244826 138454
rect 245062 138218 245146 138454
rect 245382 138218 280826 138454
rect 281062 138218 281146 138454
rect 281382 138218 316826 138454
rect 317062 138218 317146 138454
rect 317382 138218 352826 138454
rect 353062 138218 353146 138454
rect 353382 138218 388826 138454
rect 389062 138218 389146 138454
rect 389382 138218 424826 138454
rect 425062 138218 425146 138454
rect 425382 138218 460826 138454
rect 461062 138218 461146 138454
rect 461382 138218 496826 138454
rect 497062 138218 497146 138454
rect 497382 138218 532826 138454
rect 533062 138218 533146 138454
rect 533382 138218 568826 138454
rect 569062 138218 569146 138454
rect 569382 138218 591102 138454
rect 591338 138218 591422 138454
rect 591658 138218 592650 138454
rect -8726 138134 592650 138218
rect -8726 137898 -7734 138134
rect -7498 137898 -7414 138134
rect -7178 137898 28826 138134
rect 29062 137898 29146 138134
rect 29382 137898 64826 138134
rect 65062 137898 65146 138134
rect 65382 137898 100826 138134
rect 101062 137898 101146 138134
rect 101382 137898 208826 138134
rect 209062 137898 209146 138134
rect 209382 137898 244826 138134
rect 245062 137898 245146 138134
rect 245382 137898 280826 138134
rect 281062 137898 281146 138134
rect 281382 137898 316826 138134
rect 317062 137898 317146 138134
rect 317382 137898 352826 138134
rect 353062 137898 353146 138134
rect 353382 137898 388826 138134
rect 389062 137898 389146 138134
rect 389382 137898 424826 138134
rect 425062 137898 425146 138134
rect 425382 137898 460826 138134
rect 461062 137898 461146 138134
rect 461382 137898 496826 138134
rect 497062 137898 497146 138134
rect 497382 137898 532826 138134
rect 533062 137898 533146 138134
rect 533382 137898 568826 138134
rect 569062 137898 569146 138134
rect 569382 137898 591102 138134
rect 591338 137898 591422 138134
rect 591658 137898 592650 138134
rect -8726 137866 592650 137898
rect -8726 133954 592650 133986
rect -8726 133718 -6774 133954
rect -6538 133718 -6454 133954
rect -6218 133718 24326 133954
rect 24562 133718 24646 133954
rect 24882 133718 60326 133954
rect 60562 133718 60646 133954
rect 60882 133718 96326 133954
rect 96562 133718 96646 133954
rect 96882 133718 204326 133954
rect 204562 133718 204646 133954
rect 204882 133718 240326 133954
rect 240562 133718 240646 133954
rect 240882 133718 276326 133954
rect 276562 133718 276646 133954
rect 276882 133718 312326 133954
rect 312562 133718 312646 133954
rect 312882 133718 348326 133954
rect 348562 133718 348646 133954
rect 348882 133718 384326 133954
rect 384562 133718 384646 133954
rect 384882 133718 420326 133954
rect 420562 133718 420646 133954
rect 420882 133718 456326 133954
rect 456562 133718 456646 133954
rect 456882 133718 492326 133954
rect 492562 133718 492646 133954
rect 492882 133718 528326 133954
rect 528562 133718 528646 133954
rect 528882 133718 564326 133954
rect 564562 133718 564646 133954
rect 564882 133718 590142 133954
rect 590378 133718 590462 133954
rect 590698 133718 592650 133954
rect -8726 133634 592650 133718
rect -8726 133398 -6774 133634
rect -6538 133398 -6454 133634
rect -6218 133398 24326 133634
rect 24562 133398 24646 133634
rect 24882 133398 60326 133634
rect 60562 133398 60646 133634
rect 60882 133398 96326 133634
rect 96562 133398 96646 133634
rect 96882 133398 204326 133634
rect 204562 133398 204646 133634
rect 204882 133398 240326 133634
rect 240562 133398 240646 133634
rect 240882 133398 276326 133634
rect 276562 133398 276646 133634
rect 276882 133398 312326 133634
rect 312562 133398 312646 133634
rect 312882 133398 348326 133634
rect 348562 133398 348646 133634
rect 348882 133398 384326 133634
rect 384562 133398 384646 133634
rect 384882 133398 420326 133634
rect 420562 133398 420646 133634
rect 420882 133398 456326 133634
rect 456562 133398 456646 133634
rect 456882 133398 492326 133634
rect 492562 133398 492646 133634
rect 492882 133398 528326 133634
rect 528562 133398 528646 133634
rect 528882 133398 564326 133634
rect 564562 133398 564646 133634
rect 564882 133398 590142 133634
rect 590378 133398 590462 133634
rect 590698 133398 592650 133634
rect -8726 133366 592650 133398
rect -8726 129454 592650 129486
rect -8726 129218 -5814 129454
rect -5578 129218 -5494 129454
rect -5258 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 55826 129454
rect 56062 129218 56146 129454
rect 56382 129218 91826 129454
rect 92062 129218 92146 129454
rect 92382 129218 199826 129454
rect 200062 129218 200146 129454
rect 200382 129218 235826 129454
rect 236062 129218 236146 129454
rect 236382 129218 271826 129454
rect 272062 129218 272146 129454
rect 272382 129218 307826 129454
rect 308062 129218 308146 129454
rect 308382 129218 343826 129454
rect 344062 129218 344146 129454
rect 344382 129218 379826 129454
rect 380062 129218 380146 129454
rect 380382 129218 415826 129454
rect 416062 129218 416146 129454
rect 416382 129218 451826 129454
rect 452062 129218 452146 129454
rect 452382 129218 487826 129454
rect 488062 129218 488146 129454
rect 488382 129218 523826 129454
rect 524062 129218 524146 129454
rect 524382 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 589182 129454
rect 589418 129218 589502 129454
rect 589738 129218 592650 129454
rect -8726 129134 592650 129218
rect -8726 128898 -5814 129134
rect -5578 128898 -5494 129134
rect -5258 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 55826 129134
rect 56062 128898 56146 129134
rect 56382 128898 91826 129134
rect 92062 128898 92146 129134
rect 92382 128898 199826 129134
rect 200062 128898 200146 129134
rect 200382 128898 235826 129134
rect 236062 128898 236146 129134
rect 236382 128898 271826 129134
rect 272062 128898 272146 129134
rect 272382 128898 307826 129134
rect 308062 128898 308146 129134
rect 308382 128898 343826 129134
rect 344062 128898 344146 129134
rect 344382 128898 379826 129134
rect 380062 128898 380146 129134
rect 380382 128898 415826 129134
rect 416062 128898 416146 129134
rect 416382 128898 451826 129134
rect 452062 128898 452146 129134
rect 452382 128898 487826 129134
rect 488062 128898 488146 129134
rect 488382 128898 523826 129134
rect 524062 128898 524146 129134
rect 524382 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 589182 129134
rect 589418 128898 589502 129134
rect 589738 128898 592650 129134
rect -8726 128866 592650 128898
rect -8726 124954 592650 124986
rect -8726 124718 -4854 124954
rect -4618 124718 -4534 124954
rect -4298 124718 15326 124954
rect 15562 124718 15646 124954
rect 15882 124718 51326 124954
rect 51562 124718 51646 124954
rect 51882 124718 87326 124954
rect 87562 124718 87646 124954
rect 87882 124718 195326 124954
rect 195562 124718 195646 124954
rect 195882 124718 231326 124954
rect 231562 124718 231646 124954
rect 231882 124718 267326 124954
rect 267562 124718 267646 124954
rect 267882 124718 303326 124954
rect 303562 124718 303646 124954
rect 303882 124718 339326 124954
rect 339562 124718 339646 124954
rect 339882 124718 375326 124954
rect 375562 124718 375646 124954
rect 375882 124718 411326 124954
rect 411562 124718 411646 124954
rect 411882 124718 447326 124954
rect 447562 124718 447646 124954
rect 447882 124718 483326 124954
rect 483562 124718 483646 124954
rect 483882 124718 519326 124954
rect 519562 124718 519646 124954
rect 519882 124718 555326 124954
rect 555562 124718 555646 124954
rect 555882 124718 588222 124954
rect 588458 124718 588542 124954
rect 588778 124718 592650 124954
rect -8726 124634 592650 124718
rect -8726 124398 -4854 124634
rect -4618 124398 -4534 124634
rect -4298 124398 15326 124634
rect 15562 124398 15646 124634
rect 15882 124398 51326 124634
rect 51562 124398 51646 124634
rect 51882 124398 87326 124634
rect 87562 124398 87646 124634
rect 87882 124398 195326 124634
rect 195562 124398 195646 124634
rect 195882 124398 231326 124634
rect 231562 124398 231646 124634
rect 231882 124398 267326 124634
rect 267562 124398 267646 124634
rect 267882 124398 303326 124634
rect 303562 124398 303646 124634
rect 303882 124398 339326 124634
rect 339562 124398 339646 124634
rect 339882 124398 375326 124634
rect 375562 124398 375646 124634
rect 375882 124398 411326 124634
rect 411562 124398 411646 124634
rect 411882 124398 447326 124634
rect 447562 124398 447646 124634
rect 447882 124398 483326 124634
rect 483562 124398 483646 124634
rect 483882 124398 519326 124634
rect 519562 124398 519646 124634
rect 519882 124398 555326 124634
rect 555562 124398 555646 124634
rect 555882 124398 588222 124634
rect 588458 124398 588542 124634
rect 588778 124398 592650 124634
rect -8726 124366 592650 124398
rect -8726 120454 592650 120486
rect -8726 120218 -3894 120454
rect -3658 120218 -3574 120454
rect -3338 120218 10826 120454
rect 11062 120218 11146 120454
rect 11382 120218 46826 120454
rect 47062 120218 47146 120454
rect 47382 120218 82826 120454
rect 83062 120218 83146 120454
rect 83382 120218 226826 120454
rect 227062 120218 227146 120454
rect 227382 120218 262826 120454
rect 263062 120218 263146 120454
rect 263382 120218 298826 120454
rect 299062 120218 299146 120454
rect 299382 120218 334826 120454
rect 335062 120218 335146 120454
rect 335382 120218 370826 120454
rect 371062 120218 371146 120454
rect 371382 120218 406826 120454
rect 407062 120218 407146 120454
rect 407382 120218 442826 120454
rect 443062 120218 443146 120454
rect 443382 120218 478826 120454
rect 479062 120218 479146 120454
rect 479382 120218 514826 120454
rect 515062 120218 515146 120454
rect 515382 120218 550826 120454
rect 551062 120218 551146 120454
rect 551382 120218 587262 120454
rect 587498 120218 587582 120454
rect 587818 120218 592650 120454
rect -8726 120134 592650 120218
rect -8726 119898 -3894 120134
rect -3658 119898 -3574 120134
rect -3338 119898 10826 120134
rect 11062 119898 11146 120134
rect 11382 119898 46826 120134
rect 47062 119898 47146 120134
rect 47382 119898 82826 120134
rect 83062 119898 83146 120134
rect 83382 119898 226826 120134
rect 227062 119898 227146 120134
rect 227382 119898 262826 120134
rect 263062 119898 263146 120134
rect 263382 119898 298826 120134
rect 299062 119898 299146 120134
rect 299382 119898 334826 120134
rect 335062 119898 335146 120134
rect 335382 119898 370826 120134
rect 371062 119898 371146 120134
rect 371382 119898 406826 120134
rect 407062 119898 407146 120134
rect 407382 119898 442826 120134
rect 443062 119898 443146 120134
rect 443382 119898 478826 120134
rect 479062 119898 479146 120134
rect 479382 119898 514826 120134
rect 515062 119898 515146 120134
rect 515382 119898 550826 120134
rect 551062 119898 551146 120134
rect 551382 119898 587262 120134
rect 587498 119898 587582 120134
rect 587818 119898 592650 120134
rect -8726 119866 592650 119898
rect -8726 115954 592650 115986
rect -8726 115718 -2934 115954
rect -2698 115718 -2614 115954
rect -2378 115718 6326 115954
rect 6562 115718 6646 115954
rect 6882 115718 42326 115954
rect 42562 115718 42646 115954
rect 42882 115718 78326 115954
rect 78562 115718 78646 115954
rect 78882 115718 114326 115954
rect 114562 115718 114646 115954
rect 114882 115718 139610 115954
rect 139846 115718 170330 115954
rect 170566 115718 222326 115954
rect 222562 115718 222646 115954
rect 222882 115718 258326 115954
rect 258562 115718 258646 115954
rect 258882 115718 294326 115954
rect 294562 115718 294646 115954
rect 294882 115718 330326 115954
rect 330562 115718 330646 115954
rect 330882 115718 366326 115954
rect 366562 115718 366646 115954
rect 366882 115718 402326 115954
rect 402562 115718 402646 115954
rect 402882 115718 438326 115954
rect 438562 115718 438646 115954
rect 438882 115718 474326 115954
rect 474562 115718 474646 115954
rect 474882 115718 510326 115954
rect 510562 115718 510646 115954
rect 510882 115718 546326 115954
rect 546562 115718 546646 115954
rect 546882 115718 582326 115954
rect 582562 115718 582646 115954
rect 582882 115718 586302 115954
rect 586538 115718 586622 115954
rect 586858 115718 592650 115954
rect -8726 115634 592650 115718
rect -8726 115398 -2934 115634
rect -2698 115398 -2614 115634
rect -2378 115398 6326 115634
rect 6562 115398 6646 115634
rect 6882 115398 42326 115634
rect 42562 115398 42646 115634
rect 42882 115398 78326 115634
rect 78562 115398 78646 115634
rect 78882 115398 114326 115634
rect 114562 115398 114646 115634
rect 114882 115398 139610 115634
rect 139846 115398 170330 115634
rect 170566 115398 222326 115634
rect 222562 115398 222646 115634
rect 222882 115398 258326 115634
rect 258562 115398 258646 115634
rect 258882 115398 294326 115634
rect 294562 115398 294646 115634
rect 294882 115398 330326 115634
rect 330562 115398 330646 115634
rect 330882 115398 366326 115634
rect 366562 115398 366646 115634
rect 366882 115398 402326 115634
rect 402562 115398 402646 115634
rect 402882 115398 438326 115634
rect 438562 115398 438646 115634
rect 438882 115398 474326 115634
rect 474562 115398 474646 115634
rect 474882 115398 510326 115634
rect 510562 115398 510646 115634
rect 510882 115398 546326 115634
rect 546562 115398 546646 115634
rect 546882 115398 582326 115634
rect 582562 115398 582646 115634
rect 582882 115398 586302 115634
rect 586538 115398 586622 115634
rect 586858 115398 592650 115634
rect -8726 115366 592650 115398
rect -8726 111454 592650 111486
rect -8726 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 73826 111454
rect 74062 111218 74146 111454
rect 74382 111218 109826 111454
rect 110062 111218 110146 111454
rect 110382 111218 124250 111454
rect 124486 111218 154970 111454
rect 155206 111218 185690 111454
rect 185926 111218 217826 111454
rect 218062 111218 218146 111454
rect 218382 111218 253826 111454
rect 254062 111218 254146 111454
rect 254382 111218 289826 111454
rect 290062 111218 290146 111454
rect 290382 111218 325826 111454
rect 326062 111218 326146 111454
rect 326382 111218 361826 111454
rect 362062 111218 362146 111454
rect 362382 111218 397826 111454
rect 398062 111218 398146 111454
rect 398382 111218 433826 111454
rect 434062 111218 434146 111454
rect 434382 111218 469826 111454
rect 470062 111218 470146 111454
rect 470382 111218 505826 111454
rect 506062 111218 506146 111454
rect 506382 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 592650 111454
rect -8726 111134 592650 111218
rect -8726 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 73826 111134
rect 74062 110898 74146 111134
rect 74382 110898 109826 111134
rect 110062 110898 110146 111134
rect 110382 110898 124250 111134
rect 124486 110898 154970 111134
rect 155206 110898 185690 111134
rect 185926 110898 217826 111134
rect 218062 110898 218146 111134
rect 218382 110898 253826 111134
rect 254062 110898 254146 111134
rect 254382 110898 289826 111134
rect 290062 110898 290146 111134
rect 290382 110898 325826 111134
rect 326062 110898 326146 111134
rect 326382 110898 361826 111134
rect 362062 110898 362146 111134
rect 362382 110898 397826 111134
rect 398062 110898 398146 111134
rect 398382 110898 433826 111134
rect 434062 110898 434146 111134
rect 434382 110898 469826 111134
rect 470062 110898 470146 111134
rect 470382 110898 505826 111134
rect 506062 110898 506146 111134
rect 506382 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 592650 111134
rect -8726 110866 592650 110898
rect -8726 106954 592650 106986
rect -8726 106718 -8694 106954
rect -8458 106718 -8374 106954
rect -8138 106718 33326 106954
rect 33562 106718 33646 106954
rect 33882 106718 69326 106954
rect 69562 106718 69646 106954
rect 69882 106718 105326 106954
rect 105562 106718 105646 106954
rect 105882 106718 213326 106954
rect 213562 106718 213646 106954
rect 213882 106718 249326 106954
rect 249562 106718 249646 106954
rect 249882 106718 285326 106954
rect 285562 106718 285646 106954
rect 285882 106718 321326 106954
rect 321562 106718 321646 106954
rect 321882 106718 357326 106954
rect 357562 106718 357646 106954
rect 357882 106718 393326 106954
rect 393562 106718 393646 106954
rect 393882 106718 429326 106954
rect 429562 106718 429646 106954
rect 429882 106718 465326 106954
rect 465562 106718 465646 106954
rect 465882 106718 501326 106954
rect 501562 106718 501646 106954
rect 501882 106718 537326 106954
rect 537562 106718 537646 106954
rect 537882 106718 573326 106954
rect 573562 106718 573646 106954
rect 573882 106718 592062 106954
rect 592298 106718 592382 106954
rect 592618 106718 592650 106954
rect -8726 106634 592650 106718
rect -8726 106398 -8694 106634
rect -8458 106398 -8374 106634
rect -8138 106398 33326 106634
rect 33562 106398 33646 106634
rect 33882 106398 69326 106634
rect 69562 106398 69646 106634
rect 69882 106398 105326 106634
rect 105562 106398 105646 106634
rect 105882 106398 213326 106634
rect 213562 106398 213646 106634
rect 213882 106398 249326 106634
rect 249562 106398 249646 106634
rect 249882 106398 285326 106634
rect 285562 106398 285646 106634
rect 285882 106398 321326 106634
rect 321562 106398 321646 106634
rect 321882 106398 357326 106634
rect 357562 106398 357646 106634
rect 357882 106398 393326 106634
rect 393562 106398 393646 106634
rect 393882 106398 429326 106634
rect 429562 106398 429646 106634
rect 429882 106398 465326 106634
rect 465562 106398 465646 106634
rect 465882 106398 501326 106634
rect 501562 106398 501646 106634
rect 501882 106398 537326 106634
rect 537562 106398 537646 106634
rect 537882 106398 573326 106634
rect 573562 106398 573646 106634
rect 573882 106398 592062 106634
rect 592298 106398 592382 106634
rect 592618 106398 592650 106634
rect -8726 106366 592650 106398
rect -8726 102454 592650 102486
rect -8726 102218 -7734 102454
rect -7498 102218 -7414 102454
rect -7178 102218 28826 102454
rect 29062 102218 29146 102454
rect 29382 102218 64826 102454
rect 65062 102218 65146 102454
rect 65382 102218 100826 102454
rect 101062 102218 101146 102454
rect 101382 102218 208826 102454
rect 209062 102218 209146 102454
rect 209382 102218 244826 102454
rect 245062 102218 245146 102454
rect 245382 102218 280826 102454
rect 281062 102218 281146 102454
rect 281382 102218 316826 102454
rect 317062 102218 317146 102454
rect 317382 102218 352826 102454
rect 353062 102218 353146 102454
rect 353382 102218 388826 102454
rect 389062 102218 389146 102454
rect 389382 102218 424826 102454
rect 425062 102218 425146 102454
rect 425382 102218 460826 102454
rect 461062 102218 461146 102454
rect 461382 102218 496826 102454
rect 497062 102218 497146 102454
rect 497382 102218 532826 102454
rect 533062 102218 533146 102454
rect 533382 102218 568826 102454
rect 569062 102218 569146 102454
rect 569382 102218 591102 102454
rect 591338 102218 591422 102454
rect 591658 102218 592650 102454
rect -8726 102134 592650 102218
rect -8726 101898 -7734 102134
rect -7498 101898 -7414 102134
rect -7178 101898 28826 102134
rect 29062 101898 29146 102134
rect 29382 101898 64826 102134
rect 65062 101898 65146 102134
rect 65382 101898 100826 102134
rect 101062 101898 101146 102134
rect 101382 101898 208826 102134
rect 209062 101898 209146 102134
rect 209382 101898 244826 102134
rect 245062 101898 245146 102134
rect 245382 101898 280826 102134
rect 281062 101898 281146 102134
rect 281382 101898 316826 102134
rect 317062 101898 317146 102134
rect 317382 101898 352826 102134
rect 353062 101898 353146 102134
rect 353382 101898 388826 102134
rect 389062 101898 389146 102134
rect 389382 101898 424826 102134
rect 425062 101898 425146 102134
rect 425382 101898 460826 102134
rect 461062 101898 461146 102134
rect 461382 101898 496826 102134
rect 497062 101898 497146 102134
rect 497382 101898 532826 102134
rect 533062 101898 533146 102134
rect 533382 101898 568826 102134
rect 569062 101898 569146 102134
rect 569382 101898 591102 102134
rect 591338 101898 591422 102134
rect 591658 101898 592650 102134
rect -8726 101866 592650 101898
rect -8726 97954 592650 97986
rect -8726 97718 -6774 97954
rect -6538 97718 -6454 97954
rect -6218 97718 24326 97954
rect 24562 97718 24646 97954
rect 24882 97718 60326 97954
rect 60562 97718 60646 97954
rect 60882 97718 96326 97954
rect 96562 97718 96646 97954
rect 96882 97718 204326 97954
rect 204562 97718 204646 97954
rect 204882 97718 240326 97954
rect 240562 97718 240646 97954
rect 240882 97718 276326 97954
rect 276562 97718 276646 97954
rect 276882 97718 312326 97954
rect 312562 97718 312646 97954
rect 312882 97718 348326 97954
rect 348562 97718 348646 97954
rect 348882 97718 384326 97954
rect 384562 97718 384646 97954
rect 384882 97718 420326 97954
rect 420562 97718 420646 97954
rect 420882 97718 456326 97954
rect 456562 97718 456646 97954
rect 456882 97718 492326 97954
rect 492562 97718 492646 97954
rect 492882 97718 528326 97954
rect 528562 97718 528646 97954
rect 528882 97718 564326 97954
rect 564562 97718 564646 97954
rect 564882 97718 590142 97954
rect 590378 97718 590462 97954
rect 590698 97718 592650 97954
rect -8726 97634 592650 97718
rect -8726 97398 -6774 97634
rect -6538 97398 -6454 97634
rect -6218 97398 24326 97634
rect 24562 97398 24646 97634
rect 24882 97398 60326 97634
rect 60562 97398 60646 97634
rect 60882 97398 96326 97634
rect 96562 97398 96646 97634
rect 96882 97398 204326 97634
rect 204562 97398 204646 97634
rect 204882 97398 240326 97634
rect 240562 97398 240646 97634
rect 240882 97398 276326 97634
rect 276562 97398 276646 97634
rect 276882 97398 312326 97634
rect 312562 97398 312646 97634
rect 312882 97398 348326 97634
rect 348562 97398 348646 97634
rect 348882 97398 384326 97634
rect 384562 97398 384646 97634
rect 384882 97398 420326 97634
rect 420562 97398 420646 97634
rect 420882 97398 456326 97634
rect 456562 97398 456646 97634
rect 456882 97398 492326 97634
rect 492562 97398 492646 97634
rect 492882 97398 528326 97634
rect 528562 97398 528646 97634
rect 528882 97398 564326 97634
rect 564562 97398 564646 97634
rect 564882 97398 590142 97634
rect 590378 97398 590462 97634
rect 590698 97398 592650 97634
rect -8726 97366 592650 97398
rect -8726 93454 592650 93486
rect -8726 93218 -5814 93454
rect -5578 93218 -5494 93454
rect -5258 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 55826 93454
rect 56062 93218 56146 93454
rect 56382 93218 91826 93454
rect 92062 93218 92146 93454
rect 92382 93218 199826 93454
rect 200062 93218 200146 93454
rect 200382 93218 235826 93454
rect 236062 93218 236146 93454
rect 236382 93218 271826 93454
rect 272062 93218 272146 93454
rect 272382 93218 307826 93454
rect 308062 93218 308146 93454
rect 308382 93218 343826 93454
rect 344062 93218 344146 93454
rect 344382 93218 379826 93454
rect 380062 93218 380146 93454
rect 380382 93218 415826 93454
rect 416062 93218 416146 93454
rect 416382 93218 451826 93454
rect 452062 93218 452146 93454
rect 452382 93218 487826 93454
rect 488062 93218 488146 93454
rect 488382 93218 523826 93454
rect 524062 93218 524146 93454
rect 524382 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 589182 93454
rect 589418 93218 589502 93454
rect 589738 93218 592650 93454
rect -8726 93134 592650 93218
rect -8726 92898 -5814 93134
rect -5578 92898 -5494 93134
rect -5258 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 55826 93134
rect 56062 92898 56146 93134
rect 56382 92898 91826 93134
rect 92062 92898 92146 93134
rect 92382 92898 199826 93134
rect 200062 92898 200146 93134
rect 200382 92898 235826 93134
rect 236062 92898 236146 93134
rect 236382 92898 271826 93134
rect 272062 92898 272146 93134
rect 272382 92898 307826 93134
rect 308062 92898 308146 93134
rect 308382 92898 343826 93134
rect 344062 92898 344146 93134
rect 344382 92898 379826 93134
rect 380062 92898 380146 93134
rect 380382 92898 415826 93134
rect 416062 92898 416146 93134
rect 416382 92898 451826 93134
rect 452062 92898 452146 93134
rect 452382 92898 487826 93134
rect 488062 92898 488146 93134
rect 488382 92898 523826 93134
rect 524062 92898 524146 93134
rect 524382 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 589182 93134
rect 589418 92898 589502 93134
rect 589738 92898 592650 93134
rect -8726 92866 592650 92898
rect -8726 88954 592650 88986
rect -8726 88718 -4854 88954
rect -4618 88718 -4534 88954
rect -4298 88718 15326 88954
rect 15562 88718 15646 88954
rect 15882 88718 51326 88954
rect 51562 88718 51646 88954
rect 51882 88718 87326 88954
rect 87562 88718 87646 88954
rect 87882 88718 195326 88954
rect 195562 88718 195646 88954
rect 195882 88718 231326 88954
rect 231562 88718 231646 88954
rect 231882 88718 267326 88954
rect 267562 88718 267646 88954
rect 267882 88718 303326 88954
rect 303562 88718 303646 88954
rect 303882 88718 339326 88954
rect 339562 88718 339646 88954
rect 339882 88718 375326 88954
rect 375562 88718 375646 88954
rect 375882 88718 411326 88954
rect 411562 88718 411646 88954
rect 411882 88718 447326 88954
rect 447562 88718 447646 88954
rect 447882 88718 483326 88954
rect 483562 88718 483646 88954
rect 483882 88718 519326 88954
rect 519562 88718 519646 88954
rect 519882 88718 555326 88954
rect 555562 88718 555646 88954
rect 555882 88718 588222 88954
rect 588458 88718 588542 88954
rect 588778 88718 592650 88954
rect -8726 88634 592650 88718
rect -8726 88398 -4854 88634
rect -4618 88398 -4534 88634
rect -4298 88398 15326 88634
rect 15562 88398 15646 88634
rect 15882 88398 51326 88634
rect 51562 88398 51646 88634
rect 51882 88398 87326 88634
rect 87562 88398 87646 88634
rect 87882 88398 195326 88634
rect 195562 88398 195646 88634
rect 195882 88398 231326 88634
rect 231562 88398 231646 88634
rect 231882 88398 267326 88634
rect 267562 88398 267646 88634
rect 267882 88398 303326 88634
rect 303562 88398 303646 88634
rect 303882 88398 339326 88634
rect 339562 88398 339646 88634
rect 339882 88398 375326 88634
rect 375562 88398 375646 88634
rect 375882 88398 411326 88634
rect 411562 88398 411646 88634
rect 411882 88398 447326 88634
rect 447562 88398 447646 88634
rect 447882 88398 483326 88634
rect 483562 88398 483646 88634
rect 483882 88398 519326 88634
rect 519562 88398 519646 88634
rect 519882 88398 555326 88634
rect 555562 88398 555646 88634
rect 555882 88398 588222 88634
rect 588458 88398 588542 88634
rect 588778 88398 592650 88634
rect -8726 88366 592650 88398
rect -8726 84454 592650 84486
rect -8726 84218 -3894 84454
rect -3658 84218 -3574 84454
rect -3338 84218 10826 84454
rect 11062 84218 11146 84454
rect 11382 84218 46826 84454
rect 47062 84218 47146 84454
rect 47382 84218 82826 84454
rect 83062 84218 83146 84454
rect 83382 84218 226826 84454
rect 227062 84218 227146 84454
rect 227382 84218 262826 84454
rect 263062 84218 263146 84454
rect 263382 84218 298826 84454
rect 299062 84218 299146 84454
rect 299382 84218 334826 84454
rect 335062 84218 335146 84454
rect 335382 84218 370826 84454
rect 371062 84218 371146 84454
rect 371382 84218 406826 84454
rect 407062 84218 407146 84454
rect 407382 84218 442826 84454
rect 443062 84218 443146 84454
rect 443382 84218 478826 84454
rect 479062 84218 479146 84454
rect 479382 84218 514826 84454
rect 515062 84218 515146 84454
rect 515382 84218 550826 84454
rect 551062 84218 551146 84454
rect 551382 84218 587262 84454
rect 587498 84218 587582 84454
rect 587818 84218 592650 84454
rect -8726 84134 592650 84218
rect -8726 83898 -3894 84134
rect -3658 83898 -3574 84134
rect -3338 83898 10826 84134
rect 11062 83898 11146 84134
rect 11382 83898 46826 84134
rect 47062 83898 47146 84134
rect 47382 83898 82826 84134
rect 83062 83898 83146 84134
rect 83382 83898 226826 84134
rect 227062 83898 227146 84134
rect 227382 83898 262826 84134
rect 263062 83898 263146 84134
rect 263382 83898 298826 84134
rect 299062 83898 299146 84134
rect 299382 83898 334826 84134
rect 335062 83898 335146 84134
rect 335382 83898 370826 84134
rect 371062 83898 371146 84134
rect 371382 83898 406826 84134
rect 407062 83898 407146 84134
rect 407382 83898 442826 84134
rect 443062 83898 443146 84134
rect 443382 83898 478826 84134
rect 479062 83898 479146 84134
rect 479382 83898 514826 84134
rect 515062 83898 515146 84134
rect 515382 83898 550826 84134
rect 551062 83898 551146 84134
rect 551382 83898 587262 84134
rect 587498 83898 587582 84134
rect 587818 83898 592650 84134
rect -8726 83866 592650 83898
rect -8726 79954 592650 79986
rect -8726 79718 -2934 79954
rect -2698 79718 -2614 79954
rect -2378 79718 6326 79954
rect 6562 79718 6646 79954
rect 6882 79718 42326 79954
rect 42562 79718 42646 79954
rect 42882 79718 78326 79954
rect 78562 79718 78646 79954
rect 78882 79718 114326 79954
rect 114562 79718 114646 79954
rect 114882 79718 222326 79954
rect 222562 79718 222646 79954
rect 222882 79718 258326 79954
rect 258562 79718 258646 79954
rect 258882 79718 294326 79954
rect 294562 79718 294646 79954
rect 294882 79718 330326 79954
rect 330562 79718 330646 79954
rect 330882 79718 366326 79954
rect 366562 79718 366646 79954
rect 366882 79718 402326 79954
rect 402562 79718 402646 79954
rect 402882 79718 438326 79954
rect 438562 79718 438646 79954
rect 438882 79718 474326 79954
rect 474562 79718 474646 79954
rect 474882 79718 510326 79954
rect 510562 79718 510646 79954
rect 510882 79718 546326 79954
rect 546562 79718 546646 79954
rect 546882 79718 582326 79954
rect 582562 79718 582646 79954
rect 582882 79718 586302 79954
rect 586538 79718 586622 79954
rect 586858 79718 592650 79954
rect -8726 79634 592650 79718
rect -8726 79398 -2934 79634
rect -2698 79398 -2614 79634
rect -2378 79398 6326 79634
rect 6562 79398 6646 79634
rect 6882 79398 42326 79634
rect 42562 79398 42646 79634
rect 42882 79398 78326 79634
rect 78562 79398 78646 79634
rect 78882 79398 114326 79634
rect 114562 79398 114646 79634
rect 114882 79398 222326 79634
rect 222562 79398 222646 79634
rect 222882 79398 258326 79634
rect 258562 79398 258646 79634
rect 258882 79398 294326 79634
rect 294562 79398 294646 79634
rect 294882 79398 330326 79634
rect 330562 79398 330646 79634
rect 330882 79398 366326 79634
rect 366562 79398 366646 79634
rect 366882 79398 402326 79634
rect 402562 79398 402646 79634
rect 402882 79398 438326 79634
rect 438562 79398 438646 79634
rect 438882 79398 474326 79634
rect 474562 79398 474646 79634
rect 474882 79398 510326 79634
rect 510562 79398 510646 79634
rect 510882 79398 546326 79634
rect 546562 79398 546646 79634
rect 546882 79398 582326 79634
rect 582562 79398 582646 79634
rect 582882 79398 586302 79634
rect 586538 79398 586622 79634
rect 586858 79398 592650 79634
rect -8726 79366 592650 79398
rect -8726 75454 592650 75486
rect -8726 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 73826 75454
rect 74062 75218 74146 75454
rect 74382 75218 109826 75454
rect 110062 75218 110146 75454
rect 110382 75218 145826 75454
rect 146062 75218 146146 75454
rect 146382 75218 181826 75454
rect 182062 75218 182146 75454
rect 182382 75218 217826 75454
rect 218062 75218 218146 75454
rect 218382 75218 253826 75454
rect 254062 75218 254146 75454
rect 254382 75218 289826 75454
rect 290062 75218 290146 75454
rect 290382 75218 325826 75454
rect 326062 75218 326146 75454
rect 326382 75218 361826 75454
rect 362062 75218 362146 75454
rect 362382 75218 397826 75454
rect 398062 75218 398146 75454
rect 398382 75218 433826 75454
rect 434062 75218 434146 75454
rect 434382 75218 469826 75454
rect 470062 75218 470146 75454
rect 470382 75218 505826 75454
rect 506062 75218 506146 75454
rect 506382 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 592650 75454
rect -8726 75134 592650 75218
rect -8726 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 73826 75134
rect 74062 74898 74146 75134
rect 74382 74898 109826 75134
rect 110062 74898 110146 75134
rect 110382 74898 145826 75134
rect 146062 74898 146146 75134
rect 146382 74898 181826 75134
rect 182062 74898 182146 75134
rect 182382 74898 217826 75134
rect 218062 74898 218146 75134
rect 218382 74898 253826 75134
rect 254062 74898 254146 75134
rect 254382 74898 289826 75134
rect 290062 74898 290146 75134
rect 290382 74898 325826 75134
rect 326062 74898 326146 75134
rect 326382 74898 361826 75134
rect 362062 74898 362146 75134
rect 362382 74898 397826 75134
rect 398062 74898 398146 75134
rect 398382 74898 433826 75134
rect 434062 74898 434146 75134
rect 434382 74898 469826 75134
rect 470062 74898 470146 75134
rect 470382 74898 505826 75134
rect 506062 74898 506146 75134
rect 506382 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 592650 75134
rect -8726 74866 592650 74898
rect -8726 70954 592650 70986
rect -8726 70718 -8694 70954
rect -8458 70718 -8374 70954
rect -8138 70718 33326 70954
rect 33562 70718 33646 70954
rect 33882 70718 69326 70954
rect 69562 70718 69646 70954
rect 69882 70718 105326 70954
rect 105562 70718 105646 70954
rect 105882 70718 141326 70954
rect 141562 70718 141646 70954
rect 141882 70718 177326 70954
rect 177562 70718 177646 70954
rect 177882 70718 213326 70954
rect 213562 70718 213646 70954
rect 213882 70718 249326 70954
rect 249562 70718 249646 70954
rect 249882 70718 285326 70954
rect 285562 70718 285646 70954
rect 285882 70718 321326 70954
rect 321562 70718 321646 70954
rect 321882 70718 357326 70954
rect 357562 70718 357646 70954
rect 357882 70718 393326 70954
rect 393562 70718 393646 70954
rect 393882 70718 429326 70954
rect 429562 70718 429646 70954
rect 429882 70718 465326 70954
rect 465562 70718 465646 70954
rect 465882 70718 501326 70954
rect 501562 70718 501646 70954
rect 501882 70718 537326 70954
rect 537562 70718 537646 70954
rect 537882 70718 573326 70954
rect 573562 70718 573646 70954
rect 573882 70718 592062 70954
rect 592298 70718 592382 70954
rect 592618 70718 592650 70954
rect -8726 70634 592650 70718
rect -8726 70398 -8694 70634
rect -8458 70398 -8374 70634
rect -8138 70398 33326 70634
rect 33562 70398 33646 70634
rect 33882 70398 69326 70634
rect 69562 70398 69646 70634
rect 69882 70398 105326 70634
rect 105562 70398 105646 70634
rect 105882 70398 141326 70634
rect 141562 70398 141646 70634
rect 141882 70398 177326 70634
rect 177562 70398 177646 70634
rect 177882 70398 213326 70634
rect 213562 70398 213646 70634
rect 213882 70398 249326 70634
rect 249562 70398 249646 70634
rect 249882 70398 285326 70634
rect 285562 70398 285646 70634
rect 285882 70398 321326 70634
rect 321562 70398 321646 70634
rect 321882 70398 357326 70634
rect 357562 70398 357646 70634
rect 357882 70398 393326 70634
rect 393562 70398 393646 70634
rect 393882 70398 429326 70634
rect 429562 70398 429646 70634
rect 429882 70398 465326 70634
rect 465562 70398 465646 70634
rect 465882 70398 501326 70634
rect 501562 70398 501646 70634
rect 501882 70398 537326 70634
rect 537562 70398 537646 70634
rect 537882 70398 573326 70634
rect 573562 70398 573646 70634
rect 573882 70398 592062 70634
rect 592298 70398 592382 70634
rect 592618 70398 592650 70634
rect -8726 70366 592650 70398
rect -8726 66454 592650 66486
rect -8726 66218 -7734 66454
rect -7498 66218 -7414 66454
rect -7178 66218 28826 66454
rect 29062 66218 29146 66454
rect 29382 66218 64826 66454
rect 65062 66218 65146 66454
rect 65382 66218 100826 66454
rect 101062 66218 101146 66454
rect 101382 66218 136826 66454
rect 137062 66218 137146 66454
rect 137382 66218 172826 66454
rect 173062 66218 173146 66454
rect 173382 66218 208826 66454
rect 209062 66218 209146 66454
rect 209382 66218 244826 66454
rect 245062 66218 245146 66454
rect 245382 66218 280826 66454
rect 281062 66218 281146 66454
rect 281382 66218 316826 66454
rect 317062 66218 317146 66454
rect 317382 66218 352826 66454
rect 353062 66218 353146 66454
rect 353382 66218 388826 66454
rect 389062 66218 389146 66454
rect 389382 66218 424826 66454
rect 425062 66218 425146 66454
rect 425382 66218 460826 66454
rect 461062 66218 461146 66454
rect 461382 66218 496826 66454
rect 497062 66218 497146 66454
rect 497382 66218 532826 66454
rect 533062 66218 533146 66454
rect 533382 66218 568826 66454
rect 569062 66218 569146 66454
rect 569382 66218 591102 66454
rect 591338 66218 591422 66454
rect 591658 66218 592650 66454
rect -8726 66134 592650 66218
rect -8726 65898 -7734 66134
rect -7498 65898 -7414 66134
rect -7178 65898 28826 66134
rect 29062 65898 29146 66134
rect 29382 65898 64826 66134
rect 65062 65898 65146 66134
rect 65382 65898 100826 66134
rect 101062 65898 101146 66134
rect 101382 65898 136826 66134
rect 137062 65898 137146 66134
rect 137382 65898 172826 66134
rect 173062 65898 173146 66134
rect 173382 65898 208826 66134
rect 209062 65898 209146 66134
rect 209382 65898 244826 66134
rect 245062 65898 245146 66134
rect 245382 65898 280826 66134
rect 281062 65898 281146 66134
rect 281382 65898 316826 66134
rect 317062 65898 317146 66134
rect 317382 65898 352826 66134
rect 353062 65898 353146 66134
rect 353382 65898 388826 66134
rect 389062 65898 389146 66134
rect 389382 65898 424826 66134
rect 425062 65898 425146 66134
rect 425382 65898 460826 66134
rect 461062 65898 461146 66134
rect 461382 65898 496826 66134
rect 497062 65898 497146 66134
rect 497382 65898 532826 66134
rect 533062 65898 533146 66134
rect 533382 65898 568826 66134
rect 569062 65898 569146 66134
rect 569382 65898 591102 66134
rect 591338 65898 591422 66134
rect 591658 65898 592650 66134
rect -8726 65866 592650 65898
rect -8726 61954 592650 61986
rect -8726 61718 -6774 61954
rect -6538 61718 -6454 61954
rect -6218 61718 24326 61954
rect 24562 61718 24646 61954
rect 24882 61718 60326 61954
rect 60562 61718 60646 61954
rect 60882 61718 96326 61954
rect 96562 61718 96646 61954
rect 96882 61718 132326 61954
rect 132562 61718 132646 61954
rect 132882 61718 168326 61954
rect 168562 61718 168646 61954
rect 168882 61718 204326 61954
rect 204562 61718 204646 61954
rect 204882 61718 240326 61954
rect 240562 61718 240646 61954
rect 240882 61718 276326 61954
rect 276562 61718 276646 61954
rect 276882 61718 312326 61954
rect 312562 61718 312646 61954
rect 312882 61718 348326 61954
rect 348562 61718 348646 61954
rect 348882 61718 384326 61954
rect 384562 61718 384646 61954
rect 384882 61718 420326 61954
rect 420562 61718 420646 61954
rect 420882 61718 456326 61954
rect 456562 61718 456646 61954
rect 456882 61718 492326 61954
rect 492562 61718 492646 61954
rect 492882 61718 528326 61954
rect 528562 61718 528646 61954
rect 528882 61718 564326 61954
rect 564562 61718 564646 61954
rect 564882 61718 590142 61954
rect 590378 61718 590462 61954
rect 590698 61718 592650 61954
rect -8726 61634 592650 61718
rect -8726 61398 -6774 61634
rect -6538 61398 -6454 61634
rect -6218 61398 24326 61634
rect 24562 61398 24646 61634
rect 24882 61398 60326 61634
rect 60562 61398 60646 61634
rect 60882 61398 96326 61634
rect 96562 61398 96646 61634
rect 96882 61398 132326 61634
rect 132562 61398 132646 61634
rect 132882 61398 168326 61634
rect 168562 61398 168646 61634
rect 168882 61398 204326 61634
rect 204562 61398 204646 61634
rect 204882 61398 240326 61634
rect 240562 61398 240646 61634
rect 240882 61398 276326 61634
rect 276562 61398 276646 61634
rect 276882 61398 312326 61634
rect 312562 61398 312646 61634
rect 312882 61398 348326 61634
rect 348562 61398 348646 61634
rect 348882 61398 384326 61634
rect 384562 61398 384646 61634
rect 384882 61398 420326 61634
rect 420562 61398 420646 61634
rect 420882 61398 456326 61634
rect 456562 61398 456646 61634
rect 456882 61398 492326 61634
rect 492562 61398 492646 61634
rect 492882 61398 528326 61634
rect 528562 61398 528646 61634
rect 528882 61398 564326 61634
rect 564562 61398 564646 61634
rect 564882 61398 590142 61634
rect 590378 61398 590462 61634
rect 590698 61398 592650 61634
rect -8726 61366 592650 61398
rect -8726 57454 592650 57486
rect -8726 57218 -5814 57454
rect -5578 57218 -5494 57454
rect -5258 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 55826 57454
rect 56062 57218 56146 57454
rect 56382 57218 91826 57454
rect 92062 57218 92146 57454
rect 92382 57218 127826 57454
rect 128062 57218 128146 57454
rect 128382 57218 163826 57454
rect 164062 57218 164146 57454
rect 164382 57218 199826 57454
rect 200062 57218 200146 57454
rect 200382 57218 235826 57454
rect 236062 57218 236146 57454
rect 236382 57218 271826 57454
rect 272062 57218 272146 57454
rect 272382 57218 307826 57454
rect 308062 57218 308146 57454
rect 308382 57218 343826 57454
rect 344062 57218 344146 57454
rect 344382 57218 379826 57454
rect 380062 57218 380146 57454
rect 380382 57218 415826 57454
rect 416062 57218 416146 57454
rect 416382 57218 451826 57454
rect 452062 57218 452146 57454
rect 452382 57218 487826 57454
rect 488062 57218 488146 57454
rect 488382 57218 523826 57454
rect 524062 57218 524146 57454
rect 524382 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 589182 57454
rect 589418 57218 589502 57454
rect 589738 57218 592650 57454
rect -8726 57134 592650 57218
rect -8726 56898 -5814 57134
rect -5578 56898 -5494 57134
rect -5258 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 55826 57134
rect 56062 56898 56146 57134
rect 56382 56898 91826 57134
rect 92062 56898 92146 57134
rect 92382 56898 127826 57134
rect 128062 56898 128146 57134
rect 128382 56898 163826 57134
rect 164062 56898 164146 57134
rect 164382 56898 199826 57134
rect 200062 56898 200146 57134
rect 200382 56898 235826 57134
rect 236062 56898 236146 57134
rect 236382 56898 271826 57134
rect 272062 56898 272146 57134
rect 272382 56898 307826 57134
rect 308062 56898 308146 57134
rect 308382 56898 343826 57134
rect 344062 56898 344146 57134
rect 344382 56898 379826 57134
rect 380062 56898 380146 57134
rect 380382 56898 415826 57134
rect 416062 56898 416146 57134
rect 416382 56898 451826 57134
rect 452062 56898 452146 57134
rect 452382 56898 487826 57134
rect 488062 56898 488146 57134
rect 488382 56898 523826 57134
rect 524062 56898 524146 57134
rect 524382 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 589182 57134
rect 589418 56898 589502 57134
rect 589738 56898 592650 57134
rect -8726 56866 592650 56898
rect -8726 52954 592650 52986
rect -8726 52718 -4854 52954
rect -4618 52718 -4534 52954
rect -4298 52718 15326 52954
rect 15562 52718 15646 52954
rect 15882 52718 51326 52954
rect 51562 52718 51646 52954
rect 51882 52718 87326 52954
rect 87562 52718 87646 52954
rect 87882 52718 123326 52954
rect 123562 52718 123646 52954
rect 123882 52718 159326 52954
rect 159562 52718 159646 52954
rect 159882 52718 195326 52954
rect 195562 52718 195646 52954
rect 195882 52718 231326 52954
rect 231562 52718 231646 52954
rect 231882 52718 267326 52954
rect 267562 52718 267646 52954
rect 267882 52718 303326 52954
rect 303562 52718 303646 52954
rect 303882 52718 339326 52954
rect 339562 52718 339646 52954
rect 339882 52718 375326 52954
rect 375562 52718 375646 52954
rect 375882 52718 411326 52954
rect 411562 52718 411646 52954
rect 411882 52718 447326 52954
rect 447562 52718 447646 52954
rect 447882 52718 483326 52954
rect 483562 52718 483646 52954
rect 483882 52718 519326 52954
rect 519562 52718 519646 52954
rect 519882 52718 555326 52954
rect 555562 52718 555646 52954
rect 555882 52718 588222 52954
rect 588458 52718 588542 52954
rect 588778 52718 592650 52954
rect -8726 52634 592650 52718
rect -8726 52398 -4854 52634
rect -4618 52398 -4534 52634
rect -4298 52398 15326 52634
rect 15562 52398 15646 52634
rect 15882 52398 51326 52634
rect 51562 52398 51646 52634
rect 51882 52398 87326 52634
rect 87562 52398 87646 52634
rect 87882 52398 123326 52634
rect 123562 52398 123646 52634
rect 123882 52398 159326 52634
rect 159562 52398 159646 52634
rect 159882 52398 195326 52634
rect 195562 52398 195646 52634
rect 195882 52398 231326 52634
rect 231562 52398 231646 52634
rect 231882 52398 267326 52634
rect 267562 52398 267646 52634
rect 267882 52398 303326 52634
rect 303562 52398 303646 52634
rect 303882 52398 339326 52634
rect 339562 52398 339646 52634
rect 339882 52398 375326 52634
rect 375562 52398 375646 52634
rect 375882 52398 411326 52634
rect 411562 52398 411646 52634
rect 411882 52398 447326 52634
rect 447562 52398 447646 52634
rect 447882 52398 483326 52634
rect 483562 52398 483646 52634
rect 483882 52398 519326 52634
rect 519562 52398 519646 52634
rect 519882 52398 555326 52634
rect 555562 52398 555646 52634
rect 555882 52398 588222 52634
rect 588458 52398 588542 52634
rect 588778 52398 592650 52634
rect -8726 52366 592650 52398
rect -8726 48454 592650 48486
rect -8726 48218 -3894 48454
rect -3658 48218 -3574 48454
rect -3338 48218 10826 48454
rect 11062 48218 11146 48454
rect 11382 48218 46826 48454
rect 47062 48218 47146 48454
rect 47382 48218 82826 48454
rect 83062 48218 83146 48454
rect 83382 48218 118826 48454
rect 119062 48218 119146 48454
rect 119382 48218 154826 48454
rect 155062 48218 155146 48454
rect 155382 48218 190826 48454
rect 191062 48218 191146 48454
rect 191382 48218 226826 48454
rect 227062 48218 227146 48454
rect 227382 48218 262826 48454
rect 263062 48218 263146 48454
rect 263382 48218 298826 48454
rect 299062 48218 299146 48454
rect 299382 48218 334826 48454
rect 335062 48218 335146 48454
rect 335382 48218 370826 48454
rect 371062 48218 371146 48454
rect 371382 48218 406826 48454
rect 407062 48218 407146 48454
rect 407382 48218 442826 48454
rect 443062 48218 443146 48454
rect 443382 48218 478826 48454
rect 479062 48218 479146 48454
rect 479382 48218 514826 48454
rect 515062 48218 515146 48454
rect 515382 48218 550826 48454
rect 551062 48218 551146 48454
rect 551382 48218 587262 48454
rect 587498 48218 587582 48454
rect 587818 48218 592650 48454
rect -8726 48134 592650 48218
rect -8726 47898 -3894 48134
rect -3658 47898 -3574 48134
rect -3338 47898 10826 48134
rect 11062 47898 11146 48134
rect 11382 47898 46826 48134
rect 47062 47898 47146 48134
rect 47382 47898 82826 48134
rect 83062 47898 83146 48134
rect 83382 47898 118826 48134
rect 119062 47898 119146 48134
rect 119382 47898 154826 48134
rect 155062 47898 155146 48134
rect 155382 47898 190826 48134
rect 191062 47898 191146 48134
rect 191382 47898 226826 48134
rect 227062 47898 227146 48134
rect 227382 47898 262826 48134
rect 263062 47898 263146 48134
rect 263382 47898 298826 48134
rect 299062 47898 299146 48134
rect 299382 47898 334826 48134
rect 335062 47898 335146 48134
rect 335382 47898 370826 48134
rect 371062 47898 371146 48134
rect 371382 47898 406826 48134
rect 407062 47898 407146 48134
rect 407382 47898 442826 48134
rect 443062 47898 443146 48134
rect 443382 47898 478826 48134
rect 479062 47898 479146 48134
rect 479382 47898 514826 48134
rect 515062 47898 515146 48134
rect 515382 47898 550826 48134
rect 551062 47898 551146 48134
rect 551382 47898 587262 48134
rect 587498 47898 587582 48134
rect 587818 47898 592650 48134
rect -8726 47866 592650 47898
rect -8726 43954 592650 43986
rect -8726 43718 -2934 43954
rect -2698 43718 -2614 43954
rect -2378 43718 6326 43954
rect 6562 43718 6646 43954
rect 6882 43718 42326 43954
rect 42562 43718 42646 43954
rect 42882 43718 78326 43954
rect 78562 43718 78646 43954
rect 78882 43718 114326 43954
rect 114562 43718 114646 43954
rect 114882 43718 150326 43954
rect 150562 43718 150646 43954
rect 150882 43718 186326 43954
rect 186562 43718 186646 43954
rect 186882 43718 222326 43954
rect 222562 43718 222646 43954
rect 222882 43718 258326 43954
rect 258562 43718 258646 43954
rect 258882 43718 294326 43954
rect 294562 43718 294646 43954
rect 294882 43718 330326 43954
rect 330562 43718 330646 43954
rect 330882 43718 366326 43954
rect 366562 43718 366646 43954
rect 366882 43718 402326 43954
rect 402562 43718 402646 43954
rect 402882 43718 438326 43954
rect 438562 43718 438646 43954
rect 438882 43718 474326 43954
rect 474562 43718 474646 43954
rect 474882 43718 510326 43954
rect 510562 43718 510646 43954
rect 510882 43718 546326 43954
rect 546562 43718 546646 43954
rect 546882 43718 582326 43954
rect 582562 43718 582646 43954
rect 582882 43718 586302 43954
rect 586538 43718 586622 43954
rect 586858 43718 592650 43954
rect -8726 43634 592650 43718
rect -8726 43398 -2934 43634
rect -2698 43398 -2614 43634
rect -2378 43398 6326 43634
rect 6562 43398 6646 43634
rect 6882 43398 42326 43634
rect 42562 43398 42646 43634
rect 42882 43398 78326 43634
rect 78562 43398 78646 43634
rect 78882 43398 114326 43634
rect 114562 43398 114646 43634
rect 114882 43398 150326 43634
rect 150562 43398 150646 43634
rect 150882 43398 186326 43634
rect 186562 43398 186646 43634
rect 186882 43398 222326 43634
rect 222562 43398 222646 43634
rect 222882 43398 258326 43634
rect 258562 43398 258646 43634
rect 258882 43398 294326 43634
rect 294562 43398 294646 43634
rect 294882 43398 330326 43634
rect 330562 43398 330646 43634
rect 330882 43398 366326 43634
rect 366562 43398 366646 43634
rect 366882 43398 402326 43634
rect 402562 43398 402646 43634
rect 402882 43398 438326 43634
rect 438562 43398 438646 43634
rect 438882 43398 474326 43634
rect 474562 43398 474646 43634
rect 474882 43398 510326 43634
rect 510562 43398 510646 43634
rect 510882 43398 546326 43634
rect 546562 43398 546646 43634
rect 546882 43398 582326 43634
rect 582562 43398 582646 43634
rect 582882 43398 586302 43634
rect 586538 43398 586622 43634
rect 586858 43398 592650 43634
rect -8726 43366 592650 43398
rect -8726 39454 592650 39486
rect -8726 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 592650 39454
rect -8726 39134 592650 39218
rect -8726 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 592650 39134
rect -8726 38866 592650 38898
rect -8726 34954 592650 34986
rect -8726 34718 -8694 34954
rect -8458 34718 -8374 34954
rect -8138 34718 33326 34954
rect 33562 34718 33646 34954
rect 33882 34718 69326 34954
rect 69562 34718 69646 34954
rect 69882 34718 105326 34954
rect 105562 34718 105646 34954
rect 105882 34718 141326 34954
rect 141562 34718 141646 34954
rect 141882 34718 177326 34954
rect 177562 34718 177646 34954
rect 177882 34718 213326 34954
rect 213562 34718 213646 34954
rect 213882 34718 249326 34954
rect 249562 34718 249646 34954
rect 249882 34718 285326 34954
rect 285562 34718 285646 34954
rect 285882 34718 321326 34954
rect 321562 34718 321646 34954
rect 321882 34718 357326 34954
rect 357562 34718 357646 34954
rect 357882 34718 393326 34954
rect 393562 34718 393646 34954
rect 393882 34718 429326 34954
rect 429562 34718 429646 34954
rect 429882 34718 465326 34954
rect 465562 34718 465646 34954
rect 465882 34718 501326 34954
rect 501562 34718 501646 34954
rect 501882 34718 537326 34954
rect 537562 34718 537646 34954
rect 537882 34718 573326 34954
rect 573562 34718 573646 34954
rect 573882 34718 592062 34954
rect 592298 34718 592382 34954
rect 592618 34718 592650 34954
rect -8726 34634 592650 34718
rect -8726 34398 -8694 34634
rect -8458 34398 -8374 34634
rect -8138 34398 33326 34634
rect 33562 34398 33646 34634
rect 33882 34398 69326 34634
rect 69562 34398 69646 34634
rect 69882 34398 105326 34634
rect 105562 34398 105646 34634
rect 105882 34398 141326 34634
rect 141562 34398 141646 34634
rect 141882 34398 177326 34634
rect 177562 34398 177646 34634
rect 177882 34398 213326 34634
rect 213562 34398 213646 34634
rect 213882 34398 249326 34634
rect 249562 34398 249646 34634
rect 249882 34398 285326 34634
rect 285562 34398 285646 34634
rect 285882 34398 321326 34634
rect 321562 34398 321646 34634
rect 321882 34398 357326 34634
rect 357562 34398 357646 34634
rect 357882 34398 393326 34634
rect 393562 34398 393646 34634
rect 393882 34398 429326 34634
rect 429562 34398 429646 34634
rect 429882 34398 465326 34634
rect 465562 34398 465646 34634
rect 465882 34398 501326 34634
rect 501562 34398 501646 34634
rect 501882 34398 537326 34634
rect 537562 34398 537646 34634
rect 537882 34398 573326 34634
rect 573562 34398 573646 34634
rect 573882 34398 592062 34634
rect 592298 34398 592382 34634
rect 592618 34398 592650 34634
rect -8726 34366 592650 34398
rect -8726 30454 592650 30486
rect -8726 30218 -7734 30454
rect -7498 30218 -7414 30454
rect -7178 30218 28826 30454
rect 29062 30218 29146 30454
rect 29382 30218 64826 30454
rect 65062 30218 65146 30454
rect 65382 30218 100826 30454
rect 101062 30218 101146 30454
rect 101382 30218 136826 30454
rect 137062 30218 137146 30454
rect 137382 30218 172826 30454
rect 173062 30218 173146 30454
rect 173382 30218 208826 30454
rect 209062 30218 209146 30454
rect 209382 30218 244826 30454
rect 245062 30218 245146 30454
rect 245382 30218 280826 30454
rect 281062 30218 281146 30454
rect 281382 30218 316826 30454
rect 317062 30218 317146 30454
rect 317382 30218 352826 30454
rect 353062 30218 353146 30454
rect 353382 30218 388826 30454
rect 389062 30218 389146 30454
rect 389382 30218 424826 30454
rect 425062 30218 425146 30454
rect 425382 30218 460826 30454
rect 461062 30218 461146 30454
rect 461382 30218 496826 30454
rect 497062 30218 497146 30454
rect 497382 30218 532826 30454
rect 533062 30218 533146 30454
rect 533382 30218 568826 30454
rect 569062 30218 569146 30454
rect 569382 30218 591102 30454
rect 591338 30218 591422 30454
rect 591658 30218 592650 30454
rect -8726 30134 592650 30218
rect -8726 29898 -7734 30134
rect -7498 29898 -7414 30134
rect -7178 29898 28826 30134
rect 29062 29898 29146 30134
rect 29382 29898 64826 30134
rect 65062 29898 65146 30134
rect 65382 29898 100826 30134
rect 101062 29898 101146 30134
rect 101382 29898 136826 30134
rect 137062 29898 137146 30134
rect 137382 29898 172826 30134
rect 173062 29898 173146 30134
rect 173382 29898 208826 30134
rect 209062 29898 209146 30134
rect 209382 29898 244826 30134
rect 245062 29898 245146 30134
rect 245382 29898 280826 30134
rect 281062 29898 281146 30134
rect 281382 29898 316826 30134
rect 317062 29898 317146 30134
rect 317382 29898 352826 30134
rect 353062 29898 353146 30134
rect 353382 29898 388826 30134
rect 389062 29898 389146 30134
rect 389382 29898 424826 30134
rect 425062 29898 425146 30134
rect 425382 29898 460826 30134
rect 461062 29898 461146 30134
rect 461382 29898 496826 30134
rect 497062 29898 497146 30134
rect 497382 29898 532826 30134
rect 533062 29898 533146 30134
rect 533382 29898 568826 30134
rect 569062 29898 569146 30134
rect 569382 29898 591102 30134
rect 591338 29898 591422 30134
rect 591658 29898 592650 30134
rect -8726 29866 592650 29898
rect -8726 25954 592650 25986
rect -8726 25718 -6774 25954
rect -6538 25718 -6454 25954
rect -6218 25718 24326 25954
rect 24562 25718 24646 25954
rect 24882 25718 60326 25954
rect 60562 25718 60646 25954
rect 60882 25718 96326 25954
rect 96562 25718 96646 25954
rect 96882 25718 132326 25954
rect 132562 25718 132646 25954
rect 132882 25718 168326 25954
rect 168562 25718 168646 25954
rect 168882 25718 204326 25954
rect 204562 25718 204646 25954
rect 204882 25718 240326 25954
rect 240562 25718 240646 25954
rect 240882 25718 276326 25954
rect 276562 25718 276646 25954
rect 276882 25718 312326 25954
rect 312562 25718 312646 25954
rect 312882 25718 348326 25954
rect 348562 25718 348646 25954
rect 348882 25718 384326 25954
rect 384562 25718 384646 25954
rect 384882 25718 420326 25954
rect 420562 25718 420646 25954
rect 420882 25718 456326 25954
rect 456562 25718 456646 25954
rect 456882 25718 492326 25954
rect 492562 25718 492646 25954
rect 492882 25718 528326 25954
rect 528562 25718 528646 25954
rect 528882 25718 564326 25954
rect 564562 25718 564646 25954
rect 564882 25718 590142 25954
rect 590378 25718 590462 25954
rect 590698 25718 592650 25954
rect -8726 25634 592650 25718
rect -8726 25398 -6774 25634
rect -6538 25398 -6454 25634
rect -6218 25398 24326 25634
rect 24562 25398 24646 25634
rect 24882 25398 60326 25634
rect 60562 25398 60646 25634
rect 60882 25398 96326 25634
rect 96562 25398 96646 25634
rect 96882 25398 132326 25634
rect 132562 25398 132646 25634
rect 132882 25398 168326 25634
rect 168562 25398 168646 25634
rect 168882 25398 204326 25634
rect 204562 25398 204646 25634
rect 204882 25398 240326 25634
rect 240562 25398 240646 25634
rect 240882 25398 276326 25634
rect 276562 25398 276646 25634
rect 276882 25398 312326 25634
rect 312562 25398 312646 25634
rect 312882 25398 348326 25634
rect 348562 25398 348646 25634
rect 348882 25398 384326 25634
rect 384562 25398 384646 25634
rect 384882 25398 420326 25634
rect 420562 25398 420646 25634
rect 420882 25398 456326 25634
rect 456562 25398 456646 25634
rect 456882 25398 492326 25634
rect 492562 25398 492646 25634
rect 492882 25398 528326 25634
rect 528562 25398 528646 25634
rect 528882 25398 564326 25634
rect 564562 25398 564646 25634
rect 564882 25398 590142 25634
rect 590378 25398 590462 25634
rect 590698 25398 592650 25634
rect -8726 25366 592650 25398
rect -8726 21454 592650 21486
rect -8726 21218 -5814 21454
rect -5578 21218 -5494 21454
rect -5258 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 589182 21454
rect 589418 21218 589502 21454
rect 589738 21218 592650 21454
rect -8726 21134 592650 21218
rect -8726 20898 -5814 21134
rect -5578 20898 -5494 21134
rect -5258 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 589182 21134
rect 589418 20898 589502 21134
rect 589738 20898 592650 21134
rect -8726 20866 592650 20898
rect -8726 16954 592650 16986
rect -8726 16718 -4854 16954
rect -4618 16718 -4534 16954
rect -4298 16718 15326 16954
rect 15562 16718 15646 16954
rect 15882 16718 51326 16954
rect 51562 16718 51646 16954
rect 51882 16718 87326 16954
rect 87562 16718 87646 16954
rect 87882 16718 123326 16954
rect 123562 16718 123646 16954
rect 123882 16718 159326 16954
rect 159562 16718 159646 16954
rect 159882 16718 195326 16954
rect 195562 16718 195646 16954
rect 195882 16718 231326 16954
rect 231562 16718 231646 16954
rect 231882 16718 267326 16954
rect 267562 16718 267646 16954
rect 267882 16718 303326 16954
rect 303562 16718 303646 16954
rect 303882 16718 339326 16954
rect 339562 16718 339646 16954
rect 339882 16718 375326 16954
rect 375562 16718 375646 16954
rect 375882 16718 411326 16954
rect 411562 16718 411646 16954
rect 411882 16718 447326 16954
rect 447562 16718 447646 16954
rect 447882 16718 483326 16954
rect 483562 16718 483646 16954
rect 483882 16718 519326 16954
rect 519562 16718 519646 16954
rect 519882 16718 555326 16954
rect 555562 16718 555646 16954
rect 555882 16718 588222 16954
rect 588458 16718 588542 16954
rect 588778 16718 592650 16954
rect -8726 16634 592650 16718
rect -8726 16398 -4854 16634
rect -4618 16398 -4534 16634
rect -4298 16398 15326 16634
rect 15562 16398 15646 16634
rect 15882 16398 51326 16634
rect 51562 16398 51646 16634
rect 51882 16398 87326 16634
rect 87562 16398 87646 16634
rect 87882 16398 123326 16634
rect 123562 16398 123646 16634
rect 123882 16398 159326 16634
rect 159562 16398 159646 16634
rect 159882 16398 195326 16634
rect 195562 16398 195646 16634
rect 195882 16398 231326 16634
rect 231562 16398 231646 16634
rect 231882 16398 267326 16634
rect 267562 16398 267646 16634
rect 267882 16398 303326 16634
rect 303562 16398 303646 16634
rect 303882 16398 339326 16634
rect 339562 16398 339646 16634
rect 339882 16398 375326 16634
rect 375562 16398 375646 16634
rect 375882 16398 411326 16634
rect 411562 16398 411646 16634
rect 411882 16398 447326 16634
rect 447562 16398 447646 16634
rect 447882 16398 483326 16634
rect 483562 16398 483646 16634
rect 483882 16398 519326 16634
rect 519562 16398 519646 16634
rect 519882 16398 555326 16634
rect 555562 16398 555646 16634
rect 555882 16398 588222 16634
rect 588458 16398 588542 16634
rect 588778 16398 592650 16634
rect -8726 16366 592650 16398
rect -8726 12454 592650 12486
rect -8726 12218 -3894 12454
rect -3658 12218 -3574 12454
rect -3338 12218 10826 12454
rect 11062 12218 11146 12454
rect 11382 12218 46826 12454
rect 47062 12218 47146 12454
rect 47382 12218 82826 12454
rect 83062 12218 83146 12454
rect 83382 12218 118826 12454
rect 119062 12218 119146 12454
rect 119382 12218 154826 12454
rect 155062 12218 155146 12454
rect 155382 12218 190826 12454
rect 191062 12218 191146 12454
rect 191382 12218 226826 12454
rect 227062 12218 227146 12454
rect 227382 12218 262826 12454
rect 263062 12218 263146 12454
rect 263382 12218 298826 12454
rect 299062 12218 299146 12454
rect 299382 12218 334826 12454
rect 335062 12218 335146 12454
rect 335382 12218 370826 12454
rect 371062 12218 371146 12454
rect 371382 12218 406826 12454
rect 407062 12218 407146 12454
rect 407382 12218 442826 12454
rect 443062 12218 443146 12454
rect 443382 12218 478826 12454
rect 479062 12218 479146 12454
rect 479382 12218 514826 12454
rect 515062 12218 515146 12454
rect 515382 12218 550826 12454
rect 551062 12218 551146 12454
rect 551382 12218 587262 12454
rect 587498 12218 587582 12454
rect 587818 12218 592650 12454
rect -8726 12134 592650 12218
rect -8726 11898 -3894 12134
rect -3658 11898 -3574 12134
rect -3338 11898 10826 12134
rect 11062 11898 11146 12134
rect 11382 11898 46826 12134
rect 47062 11898 47146 12134
rect 47382 11898 82826 12134
rect 83062 11898 83146 12134
rect 83382 11898 118826 12134
rect 119062 11898 119146 12134
rect 119382 11898 154826 12134
rect 155062 11898 155146 12134
rect 155382 11898 190826 12134
rect 191062 11898 191146 12134
rect 191382 11898 226826 12134
rect 227062 11898 227146 12134
rect 227382 11898 262826 12134
rect 263062 11898 263146 12134
rect 263382 11898 298826 12134
rect 299062 11898 299146 12134
rect 299382 11898 334826 12134
rect 335062 11898 335146 12134
rect 335382 11898 370826 12134
rect 371062 11898 371146 12134
rect 371382 11898 406826 12134
rect 407062 11898 407146 12134
rect 407382 11898 442826 12134
rect 443062 11898 443146 12134
rect 443382 11898 478826 12134
rect 479062 11898 479146 12134
rect 479382 11898 514826 12134
rect 515062 11898 515146 12134
rect 515382 11898 550826 12134
rect 551062 11898 551146 12134
rect 551382 11898 587262 12134
rect 587498 11898 587582 12134
rect 587818 11898 592650 12134
rect -8726 11866 592650 11898
rect -8726 7954 592650 7986
rect -8726 7718 -2934 7954
rect -2698 7718 -2614 7954
rect -2378 7718 6326 7954
rect 6562 7718 6646 7954
rect 6882 7718 42326 7954
rect 42562 7718 42646 7954
rect 42882 7718 78326 7954
rect 78562 7718 78646 7954
rect 78882 7718 114326 7954
rect 114562 7718 114646 7954
rect 114882 7718 150326 7954
rect 150562 7718 150646 7954
rect 150882 7718 186326 7954
rect 186562 7718 186646 7954
rect 186882 7718 222326 7954
rect 222562 7718 222646 7954
rect 222882 7718 258326 7954
rect 258562 7718 258646 7954
rect 258882 7718 294326 7954
rect 294562 7718 294646 7954
rect 294882 7718 330326 7954
rect 330562 7718 330646 7954
rect 330882 7718 366326 7954
rect 366562 7718 366646 7954
rect 366882 7718 402326 7954
rect 402562 7718 402646 7954
rect 402882 7718 438326 7954
rect 438562 7718 438646 7954
rect 438882 7718 474326 7954
rect 474562 7718 474646 7954
rect 474882 7718 510326 7954
rect 510562 7718 510646 7954
rect 510882 7718 546326 7954
rect 546562 7718 546646 7954
rect 546882 7718 582326 7954
rect 582562 7718 582646 7954
rect 582882 7718 586302 7954
rect 586538 7718 586622 7954
rect 586858 7718 592650 7954
rect -8726 7634 592650 7718
rect -8726 7398 -2934 7634
rect -2698 7398 -2614 7634
rect -2378 7398 6326 7634
rect 6562 7398 6646 7634
rect 6882 7398 42326 7634
rect 42562 7398 42646 7634
rect 42882 7398 78326 7634
rect 78562 7398 78646 7634
rect 78882 7398 114326 7634
rect 114562 7398 114646 7634
rect 114882 7398 150326 7634
rect 150562 7398 150646 7634
rect 150882 7398 186326 7634
rect 186562 7398 186646 7634
rect 186882 7398 222326 7634
rect 222562 7398 222646 7634
rect 222882 7398 258326 7634
rect 258562 7398 258646 7634
rect 258882 7398 294326 7634
rect 294562 7398 294646 7634
rect 294882 7398 330326 7634
rect 330562 7398 330646 7634
rect 330882 7398 366326 7634
rect 366562 7398 366646 7634
rect 366882 7398 402326 7634
rect 402562 7398 402646 7634
rect 402882 7398 438326 7634
rect 438562 7398 438646 7634
rect 438882 7398 474326 7634
rect 474562 7398 474646 7634
rect 474882 7398 510326 7634
rect 510562 7398 510646 7634
rect 510882 7398 546326 7634
rect 546562 7398 546646 7634
rect 546882 7398 582326 7634
rect 582562 7398 582646 7634
rect 582882 7398 586302 7634
rect 586538 7398 586622 7634
rect 586858 7398 592650 7634
rect -8726 7366 592650 7398
rect -8726 3454 592650 3486
rect -8726 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 592650 3454
rect -8726 3134 592650 3218
rect -8726 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 592650 3134
rect -8726 2866 592650 2898
rect -2006 -346 585930 -314
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect -2006 -666 585930 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect -2006 -934 585930 -902
rect -2966 -1306 586890 -1274
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 6326 -1306
rect 6562 -1542 6646 -1306
rect 6882 -1542 42326 -1306
rect 42562 -1542 42646 -1306
rect 42882 -1542 78326 -1306
rect 78562 -1542 78646 -1306
rect 78882 -1542 114326 -1306
rect 114562 -1542 114646 -1306
rect 114882 -1542 150326 -1306
rect 150562 -1542 150646 -1306
rect 150882 -1542 186326 -1306
rect 186562 -1542 186646 -1306
rect 186882 -1542 222326 -1306
rect 222562 -1542 222646 -1306
rect 222882 -1542 258326 -1306
rect 258562 -1542 258646 -1306
rect 258882 -1542 294326 -1306
rect 294562 -1542 294646 -1306
rect 294882 -1542 330326 -1306
rect 330562 -1542 330646 -1306
rect 330882 -1542 366326 -1306
rect 366562 -1542 366646 -1306
rect 366882 -1542 402326 -1306
rect 402562 -1542 402646 -1306
rect 402882 -1542 438326 -1306
rect 438562 -1542 438646 -1306
rect 438882 -1542 474326 -1306
rect 474562 -1542 474646 -1306
rect 474882 -1542 510326 -1306
rect 510562 -1542 510646 -1306
rect 510882 -1542 546326 -1306
rect 546562 -1542 546646 -1306
rect 546882 -1542 582326 -1306
rect 582562 -1542 582646 -1306
rect 582882 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect -2966 -1626 586890 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 6326 -1626
rect 6562 -1862 6646 -1626
rect 6882 -1862 42326 -1626
rect 42562 -1862 42646 -1626
rect 42882 -1862 78326 -1626
rect 78562 -1862 78646 -1626
rect 78882 -1862 114326 -1626
rect 114562 -1862 114646 -1626
rect 114882 -1862 150326 -1626
rect 150562 -1862 150646 -1626
rect 150882 -1862 186326 -1626
rect 186562 -1862 186646 -1626
rect 186882 -1862 222326 -1626
rect 222562 -1862 222646 -1626
rect 222882 -1862 258326 -1626
rect 258562 -1862 258646 -1626
rect 258882 -1862 294326 -1626
rect 294562 -1862 294646 -1626
rect 294882 -1862 330326 -1626
rect 330562 -1862 330646 -1626
rect 330882 -1862 366326 -1626
rect 366562 -1862 366646 -1626
rect 366882 -1862 402326 -1626
rect 402562 -1862 402646 -1626
rect 402882 -1862 438326 -1626
rect 438562 -1862 438646 -1626
rect 438882 -1862 474326 -1626
rect 474562 -1862 474646 -1626
rect 474882 -1862 510326 -1626
rect 510562 -1862 510646 -1626
rect 510882 -1862 546326 -1626
rect 546562 -1862 546646 -1626
rect 546882 -1862 582326 -1626
rect 582562 -1862 582646 -1626
rect 582882 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect -2966 -1894 586890 -1862
rect -3926 -2266 587850 -2234
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 10826 -2266
rect 11062 -2502 11146 -2266
rect 11382 -2502 46826 -2266
rect 47062 -2502 47146 -2266
rect 47382 -2502 82826 -2266
rect 83062 -2502 83146 -2266
rect 83382 -2502 118826 -2266
rect 119062 -2502 119146 -2266
rect 119382 -2502 154826 -2266
rect 155062 -2502 155146 -2266
rect 155382 -2502 190826 -2266
rect 191062 -2502 191146 -2266
rect 191382 -2502 226826 -2266
rect 227062 -2502 227146 -2266
rect 227382 -2502 262826 -2266
rect 263062 -2502 263146 -2266
rect 263382 -2502 298826 -2266
rect 299062 -2502 299146 -2266
rect 299382 -2502 334826 -2266
rect 335062 -2502 335146 -2266
rect 335382 -2502 370826 -2266
rect 371062 -2502 371146 -2266
rect 371382 -2502 406826 -2266
rect 407062 -2502 407146 -2266
rect 407382 -2502 442826 -2266
rect 443062 -2502 443146 -2266
rect 443382 -2502 478826 -2266
rect 479062 -2502 479146 -2266
rect 479382 -2502 514826 -2266
rect 515062 -2502 515146 -2266
rect 515382 -2502 550826 -2266
rect 551062 -2502 551146 -2266
rect 551382 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect -3926 -2586 587850 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 10826 -2586
rect 11062 -2822 11146 -2586
rect 11382 -2822 46826 -2586
rect 47062 -2822 47146 -2586
rect 47382 -2822 82826 -2586
rect 83062 -2822 83146 -2586
rect 83382 -2822 118826 -2586
rect 119062 -2822 119146 -2586
rect 119382 -2822 154826 -2586
rect 155062 -2822 155146 -2586
rect 155382 -2822 190826 -2586
rect 191062 -2822 191146 -2586
rect 191382 -2822 226826 -2586
rect 227062 -2822 227146 -2586
rect 227382 -2822 262826 -2586
rect 263062 -2822 263146 -2586
rect 263382 -2822 298826 -2586
rect 299062 -2822 299146 -2586
rect 299382 -2822 334826 -2586
rect 335062 -2822 335146 -2586
rect 335382 -2822 370826 -2586
rect 371062 -2822 371146 -2586
rect 371382 -2822 406826 -2586
rect 407062 -2822 407146 -2586
rect 407382 -2822 442826 -2586
rect 443062 -2822 443146 -2586
rect 443382 -2822 478826 -2586
rect 479062 -2822 479146 -2586
rect 479382 -2822 514826 -2586
rect 515062 -2822 515146 -2586
rect 515382 -2822 550826 -2586
rect 551062 -2822 551146 -2586
rect 551382 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect -3926 -2854 587850 -2822
rect -4886 -3226 588810 -3194
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 15326 -3226
rect 15562 -3462 15646 -3226
rect 15882 -3462 51326 -3226
rect 51562 -3462 51646 -3226
rect 51882 -3462 87326 -3226
rect 87562 -3462 87646 -3226
rect 87882 -3462 123326 -3226
rect 123562 -3462 123646 -3226
rect 123882 -3462 159326 -3226
rect 159562 -3462 159646 -3226
rect 159882 -3462 195326 -3226
rect 195562 -3462 195646 -3226
rect 195882 -3462 231326 -3226
rect 231562 -3462 231646 -3226
rect 231882 -3462 267326 -3226
rect 267562 -3462 267646 -3226
rect 267882 -3462 303326 -3226
rect 303562 -3462 303646 -3226
rect 303882 -3462 339326 -3226
rect 339562 -3462 339646 -3226
rect 339882 -3462 375326 -3226
rect 375562 -3462 375646 -3226
rect 375882 -3462 411326 -3226
rect 411562 -3462 411646 -3226
rect 411882 -3462 447326 -3226
rect 447562 -3462 447646 -3226
rect 447882 -3462 483326 -3226
rect 483562 -3462 483646 -3226
rect 483882 -3462 519326 -3226
rect 519562 -3462 519646 -3226
rect 519882 -3462 555326 -3226
rect 555562 -3462 555646 -3226
rect 555882 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect -4886 -3546 588810 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 15326 -3546
rect 15562 -3782 15646 -3546
rect 15882 -3782 51326 -3546
rect 51562 -3782 51646 -3546
rect 51882 -3782 87326 -3546
rect 87562 -3782 87646 -3546
rect 87882 -3782 123326 -3546
rect 123562 -3782 123646 -3546
rect 123882 -3782 159326 -3546
rect 159562 -3782 159646 -3546
rect 159882 -3782 195326 -3546
rect 195562 -3782 195646 -3546
rect 195882 -3782 231326 -3546
rect 231562 -3782 231646 -3546
rect 231882 -3782 267326 -3546
rect 267562 -3782 267646 -3546
rect 267882 -3782 303326 -3546
rect 303562 -3782 303646 -3546
rect 303882 -3782 339326 -3546
rect 339562 -3782 339646 -3546
rect 339882 -3782 375326 -3546
rect 375562 -3782 375646 -3546
rect 375882 -3782 411326 -3546
rect 411562 -3782 411646 -3546
rect 411882 -3782 447326 -3546
rect 447562 -3782 447646 -3546
rect 447882 -3782 483326 -3546
rect 483562 -3782 483646 -3546
rect 483882 -3782 519326 -3546
rect 519562 -3782 519646 -3546
rect 519882 -3782 555326 -3546
rect 555562 -3782 555646 -3546
rect 555882 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect -4886 -3814 588810 -3782
rect -5846 -4186 589770 -4154
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 19826 -4186
rect 20062 -4422 20146 -4186
rect 20382 -4422 55826 -4186
rect 56062 -4422 56146 -4186
rect 56382 -4422 91826 -4186
rect 92062 -4422 92146 -4186
rect 92382 -4422 127826 -4186
rect 128062 -4422 128146 -4186
rect 128382 -4422 163826 -4186
rect 164062 -4422 164146 -4186
rect 164382 -4422 199826 -4186
rect 200062 -4422 200146 -4186
rect 200382 -4422 235826 -4186
rect 236062 -4422 236146 -4186
rect 236382 -4422 271826 -4186
rect 272062 -4422 272146 -4186
rect 272382 -4422 307826 -4186
rect 308062 -4422 308146 -4186
rect 308382 -4422 343826 -4186
rect 344062 -4422 344146 -4186
rect 344382 -4422 379826 -4186
rect 380062 -4422 380146 -4186
rect 380382 -4422 415826 -4186
rect 416062 -4422 416146 -4186
rect 416382 -4422 451826 -4186
rect 452062 -4422 452146 -4186
rect 452382 -4422 487826 -4186
rect 488062 -4422 488146 -4186
rect 488382 -4422 523826 -4186
rect 524062 -4422 524146 -4186
rect 524382 -4422 559826 -4186
rect 560062 -4422 560146 -4186
rect 560382 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect -5846 -4506 589770 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 19826 -4506
rect 20062 -4742 20146 -4506
rect 20382 -4742 55826 -4506
rect 56062 -4742 56146 -4506
rect 56382 -4742 91826 -4506
rect 92062 -4742 92146 -4506
rect 92382 -4742 127826 -4506
rect 128062 -4742 128146 -4506
rect 128382 -4742 163826 -4506
rect 164062 -4742 164146 -4506
rect 164382 -4742 199826 -4506
rect 200062 -4742 200146 -4506
rect 200382 -4742 235826 -4506
rect 236062 -4742 236146 -4506
rect 236382 -4742 271826 -4506
rect 272062 -4742 272146 -4506
rect 272382 -4742 307826 -4506
rect 308062 -4742 308146 -4506
rect 308382 -4742 343826 -4506
rect 344062 -4742 344146 -4506
rect 344382 -4742 379826 -4506
rect 380062 -4742 380146 -4506
rect 380382 -4742 415826 -4506
rect 416062 -4742 416146 -4506
rect 416382 -4742 451826 -4506
rect 452062 -4742 452146 -4506
rect 452382 -4742 487826 -4506
rect 488062 -4742 488146 -4506
rect 488382 -4742 523826 -4506
rect 524062 -4742 524146 -4506
rect 524382 -4742 559826 -4506
rect 560062 -4742 560146 -4506
rect 560382 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect -5846 -4774 589770 -4742
rect -6806 -5146 590730 -5114
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 24326 -5146
rect 24562 -5382 24646 -5146
rect 24882 -5382 60326 -5146
rect 60562 -5382 60646 -5146
rect 60882 -5382 96326 -5146
rect 96562 -5382 96646 -5146
rect 96882 -5382 132326 -5146
rect 132562 -5382 132646 -5146
rect 132882 -5382 168326 -5146
rect 168562 -5382 168646 -5146
rect 168882 -5382 204326 -5146
rect 204562 -5382 204646 -5146
rect 204882 -5382 240326 -5146
rect 240562 -5382 240646 -5146
rect 240882 -5382 276326 -5146
rect 276562 -5382 276646 -5146
rect 276882 -5382 312326 -5146
rect 312562 -5382 312646 -5146
rect 312882 -5382 348326 -5146
rect 348562 -5382 348646 -5146
rect 348882 -5382 384326 -5146
rect 384562 -5382 384646 -5146
rect 384882 -5382 420326 -5146
rect 420562 -5382 420646 -5146
rect 420882 -5382 456326 -5146
rect 456562 -5382 456646 -5146
rect 456882 -5382 492326 -5146
rect 492562 -5382 492646 -5146
rect 492882 -5382 528326 -5146
rect 528562 -5382 528646 -5146
rect 528882 -5382 564326 -5146
rect 564562 -5382 564646 -5146
rect 564882 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect -6806 -5466 590730 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 24326 -5466
rect 24562 -5702 24646 -5466
rect 24882 -5702 60326 -5466
rect 60562 -5702 60646 -5466
rect 60882 -5702 96326 -5466
rect 96562 -5702 96646 -5466
rect 96882 -5702 132326 -5466
rect 132562 -5702 132646 -5466
rect 132882 -5702 168326 -5466
rect 168562 -5702 168646 -5466
rect 168882 -5702 204326 -5466
rect 204562 -5702 204646 -5466
rect 204882 -5702 240326 -5466
rect 240562 -5702 240646 -5466
rect 240882 -5702 276326 -5466
rect 276562 -5702 276646 -5466
rect 276882 -5702 312326 -5466
rect 312562 -5702 312646 -5466
rect 312882 -5702 348326 -5466
rect 348562 -5702 348646 -5466
rect 348882 -5702 384326 -5466
rect 384562 -5702 384646 -5466
rect 384882 -5702 420326 -5466
rect 420562 -5702 420646 -5466
rect 420882 -5702 456326 -5466
rect 456562 -5702 456646 -5466
rect 456882 -5702 492326 -5466
rect 492562 -5702 492646 -5466
rect 492882 -5702 528326 -5466
rect 528562 -5702 528646 -5466
rect 528882 -5702 564326 -5466
rect 564562 -5702 564646 -5466
rect 564882 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect -6806 -5734 590730 -5702
rect -7766 -6106 591690 -6074
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 28826 -6106
rect 29062 -6342 29146 -6106
rect 29382 -6342 64826 -6106
rect 65062 -6342 65146 -6106
rect 65382 -6342 100826 -6106
rect 101062 -6342 101146 -6106
rect 101382 -6342 136826 -6106
rect 137062 -6342 137146 -6106
rect 137382 -6342 172826 -6106
rect 173062 -6342 173146 -6106
rect 173382 -6342 208826 -6106
rect 209062 -6342 209146 -6106
rect 209382 -6342 244826 -6106
rect 245062 -6342 245146 -6106
rect 245382 -6342 280826 -6106
rect 281062 -6342 281146 -6106
rect 281382 -6342 316826 -6106
rect 317062 -6342 317146 -6106
rect 317382 -6342 352826 -6106
rect 353062 -6342 353146 -6106
rect 353382 -6342 388826 -6106
rect 389062 -6342 389146 -6106
rect 389382 -6342 424826 -6106
rect 425062 -6342 425146 -6106
rect 425382 -6342 460826 -6106
rect 461062 -6342 461146 -6106
rect 461382 -6342 496826 -6106
rect 497062 -6342 497146 -6106
rect 497382 -6342 532826 -6106
rect 533062 -6342 533146 -6106
rect 533382 -6342 568826 -6106
rect 569062 -6342 569146 -6106
rect 569382 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect -7766 -6426 591690 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 28826 -6426
rect 29062 -6662 29146 -6426
rect 29382 -6662 64826 -6426
rect 65062 -6662 65146 -6426
rect 65382 -6662 100826 -6426
rect 101062 -6662 101146 -6426
rect 101382 -6662 136826 -6426
rect 137062 -6662 137146 -6426
rect 137382 -6662 172826 -6426
rect 173062 -6662 173146 -6426
rect 173382 -6662 208826 -6426
rect 209062 -6662 209146 -6426
rect 209382 -6662 244826 -6426
rect 245062 -6662 245146 -6426
rect 245382 -6662 280826 -6426
rect 281062 -6662 281146 -6426
rect 281382 -6662 316826 -6426
rect 317062 -6662 317146 -6426
rect 317382 -6662 352826 -6426
rect 353062 -6662 353146 -6426
rect 353382 -6662 388826 -6426
rect 389062 -6662 389146 -6426
rect 389382 -6662 424826 -6426
rect 425062 -6662 425146 -6426
rect 425382 -6662 460826 -6426
rect 461062 -6662 461146 -6426
rect 461382 -6662 496826 -6426
rect 497062 -6662 497146 -6426
rect 497382 -6662 532826 -6426
rect 533062 -6662 533146 -6426
rect 533382 -6662 568826 -6426
rect 569062 -6662 569146 -6426
rect 569382 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect -7766 -6694 591690 -6662
rect -8726 -7066 592650 -7034
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 33326 -7066
rect 33562 -7302 33646 -7066
rect 33882 -7302 69326 -7066
rect 69562 -7302 69646 -7066
rect 69882 -7302 105326 -7066
rect 105562 -7302 105646 -7066
rect 105882 -7302 141326 -7066
rect 141562 -7302 141646 -7066
rect 141882 -7302 177326 -7066
rect 177562 -7302 177646 -7066
rect 177882 -7302 213326 -7066
rect 213562 -7302 213646 -7066
rect 213882 -7302 249326 -7066
rect 249562 -7302 249646 -7066
rect 249882 -7302 285326 -7066
rect 285562 -7302 285646 -7066
rect 285882 -7302 321326 -7066
rect 321562 -7302 321646 -7066
rect 321882 -7302 357326 -7066
rect 357562 -7302 357646 -7066
rect 357882 -7302 393326 -7066
rect 393562 -7302 393646 -7066
rect 393882 -7302 429326 -7066
rect 429562 -7302 429646 -7066
rect 429882 -7302 465326 -7066
rect 465562 -7302 465646 -7066
rect 465882 -7302 501326 -7066
rect 501562 -7302 501646 -7066
rect 501882 -7302 537326 -7066
rect 537562 -7302 537646 -7066
rect 537882 -7302 573326 -7066
rect 573562 -7302 573646 -7066
rect 573882 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect -8726 -7386 592650 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 33326 -7386
rect 33562 -7622 33646 -7386
rect 33882 -7622 69326 -7386
rect 69562 -7622 69646 -7386
rect 69882 -7622 105326 -7386
rect 105562 -7622 105646 -7386
rect 105882 -7622 141326 -7386
rect 141562 -7622 141646 -7386
rect 141882 -7622 177326 -7386
rect 177562 -7622 177646 -7386
rect 177882 -7622 213326 -7386
rect 213562 -7622 213646 -7386
rect 213882 -7622 249326 -7386
rect 249562 -7622 249646 -7386
rect 249882 -7622 285326 -7386
rect 285562 -7622 285646 -7386
rect 285882 -7622 321326 -7386
rect 321562 -7622 321646 -7386
rect 321882 -7622 357326 -7386
rect 357562 -7622 357646 -7386
rect 357882 -7622 393326 -7386
rect 393562 -7622 393646 -7386
rect 393882 -7622 429326 -7386
rect 429562 -7622 429646 -7386
rect 429882 -7622 465326 -7386
rect 465562 -7622 465646 -7386
rect 465882 -7622 501326 -7386
rect 501562 -7622 501646 -7386
rect 501882 -7622 537326 -7386
rect 537562 -7622 537646 -7386
rect 537882 -7622 573326 -7386
rect 573562 -7622 573646 -7386
rect 573882 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect -8726 -7654 592650 -7622
use pixel_macro  pixel_macro0
timestamp 0
transform 1 0 120000 0 1 200000
box 570 0 69354 60000
use rlbp_macro  rlbp_macro0
timestamp 0
transform 1 0 120000 0 1 80000
box 1066 0 68854 60000
<< labels >>
flabel metal2 s 506174 703520 506286 704960 0 FreeSans 448 90 0 0 gpio_analog[0]
port 0 nsew signal bidirectional
flabel metal2 s 159058 -960 159170 480 0 FreeSans 448 90 0 0 gpio_analog[10]
port 1 nsew signal bidirectional
flabel metal3 s 583520 417468 584960 417708 0 FreeSans 960 0 0 0 gpio_analog[11]
port 2 nsew signal bidirectional
flabel metal3 s -960 573188 480 573428 0 FreeSans 960 0 0 0 gpio_analog[12]
port 3 nsew signal bidirectional
flabel metal3 s 583520 593588 584960 593828 0 FreeSans 960 0 0 0 gpio_analog[13]
port 4 nsew signal bidirectional
flabel metal2 s 56662 -960 56774 480 0 FreeSans 448 90 0 0 gpio_analog[14]
port 5 nsew signal bidirectional
flabel metal2 s 160346 703520 160458 704960 0 FreeSans 448 90 0 0 gpio_analog[15]
port 6 nsew signal bidirectional
flabel metal3 s 583520 212788 584960 213028 0 FreeSans 960 0 0 0 gpio_analog[16]
port 7 nsew signal bidirectional
flabel metal3 s -960 501108 480 501348 0 FreeSans 960 0 0 0 gpio_analog[17]
port 8 nsew signal bidirectional
flabel metal2 s 223458 -960 223570 480 0 FreeSans 448 90 0 0 gpio_analog[1]
port 9 nsew signal bidirectional
flabel metal3 s 583520 229108 584960 229348 0 FreeSans 960 0 0 0 gpio_analog[2]
port 10 nsew signal bidirectional
flabel metal3 s -960 268548 480 268788 0 FreeSans 960 0 0 0 gpio_analog[3]
port 11 nsew signal bidirectional
flabel metal2 s 428894 -960 429006 480 0 FreeSans 448 90 0 0 gpio_analog[4]
port 12 nsew signal bidirectional
flabel metal3 s 583520 124388 584960 124628 0 FreeSans 960 0 0 0 gpio_analog[5]
port 13 nsew signal bidirectional
flabel metal3 s 583520 513348 584960 513588 0 FreeSans 960 0 0 0 gpio_analog[6]
port 14 nsew signal bidirectional
flabel metal2 s 270470 703520 270582 704960 0 FreeSans 448 90 0 0 gpio_analog[7]
port 15 nsew signal bidirectional
flabel metal3 s 583520 329068 584960 329308 0 FreeSans 960 0 0 0 gpio_analog[8]
port 16 nsew signal bidirectional
flabel metal2 s 405710 -960 405822 480 0 FreeSans 448 90 0 0 gpio_analog[9]
port 17 nsew signal bidirectional
flabel metal2 s 37342 -960 37454 480 0 FreeSans 448 90 0 0 gpio_noesd[0]
port 18 nsew signal bidirectional
flabel metal3 s 583520 136628 584960 136868 0 FreeSans 960 0 0 0 gpio_noesd[10]
port 19 nsew signal bidirectional
flabel metal2 s 337446 -960 337558 480 0 FreeSans 448 90 0 0 gpio_noesd[11]
port 20 nsew signal bidirectional
flabel metal2 s 440486 -960 440598 480 0 FreeSans 448 90 0 0 gpio_noesd[12]
port 21 nsew signal bidirectional
flabel metal3 s -960 276028 480 276268 0 FreeSans 960 0 0 0 gpio_noesd[13]
port 22 nsew signal bidirectional
flabel metal3 s 583520 409308 584960 409548 0 FreeSans 960 0 0 0 gpio_noesd[14]
port 23 nsew signal bidirectional
flabel metal3 s 583520 120988 584960 121228 0 FreeSans 960 0 0 0 gpio_noesd[15]
port 24 nsew signal bidirectional
flabel metal3 s 583520 665668 584960 665908 0 FreeSans 960 0 0 0 gpio_noesd[16]
port 25 nsew signal bidirectional
flabel metal2 s 367714 -960 367826 480 0 FreeSans 448 90 0 0 gpio_noesd[17]
port 26 nsew signal bidirectional
flabel metal2 s 292366 -960 292478 480 0 FreeSans 448 90 0 0 gpio_noesd[1]
port 27 nsew signal bidirectional
flabel metal3 s 583520 324988 584960 325228 0 FreeSans 960 0 0 0 gpio_noesd[2]
port 28 nsew signal bidirectional
flabel metal3 s 583520 421548 584960 421788 0 FreeSans 960 0 0 0 gpio_noesd[3]
port 29 nsew signal bidirectional
flabel metal2 s 569286 -960 569398 480 0 FreeSans 448 90 0 0 gpio_noesd[4]
port 30 nsew signal bidirectional
flabel metal2 s 224746 703520 224858 704960 0 FreeSans 448 90 0 0 gpio_noesd[5]
port 31 nsew signal bidirectional
flabel metal3 s -960 669068 480 669308 0 FreeSans 960 0 0 0 gpio_noesd[6]
port 32 nsew signal bidirectional
flabel metal2 s 372866 703520 372978 704960 0 FreeSans 448 90 0 0 gpio_noesd[7]
port 33 nsew signal bidirectional
flabel metal2 s 413438 -960 413550 480 0 FreeSans 448 90 0 0 gpio_noesd[8]
port 34 nsew signal bidirectional
flabel metal3 s 583520 633708 584960 633948 0 FreeSans 960 0 0 0 gpio_noesd[9]
port 35 nsew signal bidirectional
flabel metal3 s -960 148188 480 148428 0 FreeSans 960 0 0 0 io_analog[0]
port 36 nsew signal bidirectional
flabel metal2 s 238914 -960 239026 480 0 FreeSans 448 90 0 0 io_analog[10]
port 37 nsew signal bidirectional
flabel metal2 s 130078 703520 130190 704960 0 FreeSans 448 90 0 0 io_analog[1]
port 38 nsew signal bidirectional
flabel metal3 s -960 31908 480 32148 0 FreeSans 960 0 0 0 io_analog[2]
port 39 nsew signal bidirectional
flabel metal3 s -960 203948 480 204188 0 FreeSans 960 0 0 0 io_analog[3]
port 40 nsew signal bidirectional
flabel metal2 s 60526 -960 60638 480 0 FreeSans 448 90 0 0 io_analog[4]
port 41 nsew signal bidirectional
flabel metal2 s 296874 703520 296986 704960 0 FreeSans 448 90 0 0 io_analog[5]
port 42 nsew signal bidirectional
flabel metal3 s -960 693548 480 693788 0 FreeSans 960 0 0 0 io_analog[6]
port 43 nsew signal bidirectional
flabel metal3 s 583520 561628 584960 561868 0 FreeSans 960 0 0 0 io_analog[7]
port 44 nsew signal bidirectional
flabel metal3 s -960 673148 480 673388 0 FreeSans 960 0 0 0 io_analog[8]
port 45 nsew signal bidirectional
flabel metal2 s 388322 703520 388434 704960 0 FreeSans 448 90 0 0 io_analog[9]
port 46 nsew signal bidirectional
flabel metal2 s 186750 703520 186862 704960 0 FreeSans 448 90 0 0 io_clamp_high[0]
port 47 nsew signal bidirectional
flabel metal3 s -960 424948 480 425188 0 FreeSans 960 0 0 0 io_clamp_high[1]
port 48 nsew signal bidirectional
flabel metal2 s 22530 -960 22642 480 0 FreeSans 448 90 0 0 io_clamp_high[2]
port 49 nsew signal bidirectional
flabel metal3 s 583520 618068 584960 618308 0 FreeSans 960 0 0 0 io_clamp_low[0]
port 50 nsew signal bidirectional
flabel metal3 s 583520 160428 584960 160668 0 FreeSans 960 0 0 0 io_clamp_low[1]
port 51 nsew signal bidirectional
flabel metal3 s -960 55708 480 55948 0 FreeSans 960 0 0 0 io_clamp_low[2]
port 52 nsew signal bidirectional
flabel metal3 s 583520 537828 584960 538068 0 FreeSans 960 0 0 0 io_in[0]
port 53 nsew signal input
flabel metal3 s 583520 356948 584960 357188 0 FreeSans 960 0 0 0 io_in[10]
port 54 nsew signal input
flabel metal3 s 583520 92428 584960 92668 0 FreeSans 960 0 0 0 io_in[11]
port 55 nsew signal input
flabel metal2 s 113334 -960 113446 480 0 FreeSans 448 90 0 0 io_in[12]
port 56 nsew signal input
flabel metal2 s 34766 703520 34878 704960 0 FreeSans 448 90 0 0 io_in[13]
port 57 nsew signal input
flabel metal2 s 441130 703520 441242 704960 0 FreeSans 448 90 0 0 io_in[14]
port 58 nsew signal input
flabel metal3 s 583520 216868 584960 217108 0 FreeSans 960 0 0 0 io_in[15]
port 59 nsew signal input
flabel metal2 s 493294 -960 493406 480 0 FreeSans 448 90 0 0 io_in[16]
port 60 nsew signal input
flabel metal3 s 583520 381428 584960 381668 0 FreeSans 960 0 0 0 io_in[17]
port 61 nsew signal input
flabel metal2 s 147466 -960 147578 480 0 FreeSans 448 90 0 0 io_in[18]
port 62 nsew signal input
flabel metal3 s -960 533068 480 533308 0 FreeSans 960 0 0 0 io_in[19]
port 63 nsew signal input
flabel metal2 s 95946 703520 96058 704960 0 FreeSans 448 90 0 0 io_in[1]
port 64 nsew signal input
flabel metal2 s 361918 703520 362030 704960 0 FreeSans 448 90 0 0 io_in[20]
port 65 nsew signal input
flabel metal2 s 68898 703520 69010 704960 0 FreeSans 448 90 0 0 io_in[21]
port 66 nsew signal input
flabel metal2 s 417302 -960 417414 480 0 FreeSans 448 90 0 0 io_in[22]
port 67 nsew signal input
flabel metal2 s 136518 -960 136630 480 0 FreeSans 448 90 0 0 io_in[23]
port 68 nsew signal input
flabel metal3 s -960 239988 480 240228 0 FreeSans 960 0 0 0 io_in[24]
port 69 nsew signal input
flabel metal2 s 133942 703520 134054 704960 0 FreeSans 448 90 0 0 io_in[25]
port 70 nsew signal input
flabel metal3 s 583520 485468 584960 485708 0 FreeSans 960 0 0 0 io_in[26]
port 71 nsew signal input
flabel metal2 s 98522 -960 98634 480 0 FreeSans 448 90 0 0 io_in[2]
port 72 nsew signal input
flabel metal2 s 83066 -960 83178 480 0 FreeSans 448 90 0 0 io_in[3]
port 73 nsew signal input
flabel metal3 s 583520 565708 584960 565948 0 FreeSans 960 0 0 0 io_in[4]
port 74 nsew signal input
flabel metal2 s 288502 -960 288614 480 0 FreeSans 448 90 0 0 io_in[5]
port 75 nsew signal input
flabel metal3 s -960 617388 480 617628 0 FreeSans 960 0 0 0 io_in[6]
port 76 nsew signal input
flabel metal3 s -960 340628 480 340868 0 FreeSans 960 0 0 0 io_in[7]
port 77 nsew signal input
flabel metal3 s 583520 68628 584960 68868 0 FreeSans 960 0 0 0 io_in[8]
port 78 nsew signal input
flabel metal3 s -960 192388 480 192628 0 FreeSans 960 0 0 0 io_in[9]
port 79 nsew signal input
flabel metal2 s 338734 703520 338846 704960 0 FreeSans 448 90 0 0 io_in_3v3[0]
port 80 nsew signal input
flabel metal3 s -960 392308 480 392548 0 FreeSans 960 0 0 0 io_in_3v3[10]
port 81 nsew signal input
flabel metal2 s 86930 -960 87042 480 0 FreeSans 448 90 0 0 io_in_3v3[11]
port 82 nsew signal input
flabel metal2 s 258878 703520 258990 704960 0 FreeSans 448 90 0 0 io_in_3v3[12]
port 83 nsew signal input
flabel metal2 s 122350 703520 122462 704960 0 FreeSans 448 90 0 0 io_in_3v3[13]
port 84 nsew signal input
flabel metal3 s -960 312068 480 312308 0 FreeSans 960 0 0 0 io_in_3v3[14]
port 85 nsew signal input
flabel metal3 s 583520 148868 584960 149108 0 FreeSans 960 0 0 0 io_in_3v3[15]
port 86 nsew signal input
flabel metal3 s -960 176068 480 176308 0 FreeSans 960 0 0 0 io_in_3v3[16]
port 87 nsew signal input
flabel metal2 s 10938 -960 11050 480 0 FreeSans 448 90 0 0 io_in_3v3[17]
port 88 nsew signal input
flabel metal3 s -960 649348 480 649588 0 FreeSans 960 0 0 0 io_in_3v3[18]
port 89 nsew signal input
flabel metal2 s 414726 703520 414838 704960 0 FreeSans 448 90 0 0 io_in_3v3[19]
port 90 nsew signal input
flabel metal3 s 583520 577948 584960 578188 0 FreeSans 960 0 0 0 io_in_3v3[1]
port 91 nsew signal input
flabel metal3 s -960 420868 480 421108 0 FreeSans 960 0 0 0 io_in_3v3[20]
port 92 nsew signal input
flabel metal2 s 217018 703520 217130 704960 0 FreeSans 448 90 0 0 io_in_3v3[21]
port 93 nsew signal input
flabel metal2 s 451434 -960 451546 480 0 FreeSans 448 90 0 0 io_in_3v3[22]
port 94 nsew signal input
flabel metal3 s 583520 64548 584960 64788 0 FreeSans 960 0 0 0 io_in_3v3[23]
port 95 nsew signal input
flabel metal3 s -960 628948 480 629188 0 FreeSans 960 0 0 0 io_in_3v3[24]
port 96 nsew signal input
flabel metal3 s 583520 397068 584960 397308 0 FreeSans 960 0 0 0 io_in_3v3[25]
port 97 nsew signal input
flabel metal2 s 213798 703520 213910 704960 0 FreeSans 448 90 0 0 io_in_3v3[26]
port 98 nsew signal input
flabel metal3 s 583520 650028 584960 650268 0 FreeSans 960 0 0 0 io_in_3v3[2]
port 99 nsew signal input
flabel metal3 s -960 565028 480 565268 0 FreeSans 960 0 0 0 io_in_3v3[3]
port 100 nsew signal input
flabel metal2 s 126214 703520 126326 704960 0 FreeSans 448 90 0 0 io_in_3v3[4]
port 101 nsew signal input
flabel metal2 s 273046 -960 273158 480 0 FreeSans 448 90 0 0 io_in_3v3[5]
port 102 nsew signal input
flabel metal3 s 583520 582028 584960 582268 0 FreeSans 960 0 0 0 io_in_3v3[6]
port 103 nsew signal input
flabel metal2 s 346462 703520 346574 704960 0 FreeSans 448 90 0 0 io_in_3v3[7]
port 104 nsew signal input
flabel metal3 s -960 63868 480 64108 0 FreeSans 960 0 0 0 io_in_3v3[8]
port 105 nsew signal input
flabel metal2 s 523562 -960 523674 480 0 FreeSans 448 90 0 0 io_in_3v3[9]
port 106 nsew signal input
flabel metal3 s 583520 605828 584960 606068 0 FreeSans 960 0 0 0 io_oeb[0]
port 107 nsew signal tristate
flabel metal3 s 583520 297108 584960 297348 0 FreeSans 960 0 0 0 io_oeb[10]
port 108 nsew signal tristate
flabel metal2 s 289146 703520 289258 704960 0 FreeSans 448 90 0 0 io_oeb[11]
port 109 nsew signal tristate
flabel metal2 s 212510 -960 212622 480 0 FreeSans 448 90 0 0 io_oeb[12]
port 110 nsew signal tristate
flabel metal3 s 583520 204628 584960 204868 0 FreeSans 960 0 0 0 io_oeb[13]
port 111 nsew signal tristate
flabel metal3 s -960 396388 480 396628 0 FreeSans 960 0 0 0 io_oeb[14]
port 112 nsew signal tristate
flabel metal3 s 583520 172668 584960 172908 0 FreeSans 960 0 0 0 io_oeb[15]
port 113 nsew signal tristate
flabel metal3 s 583520 168588 584960 168828 0 FreeSans 960 0 0 0 io_oeb[16]
port 114 nsew signal tristate
flabel metal3 s -960 119628 480 119868 0 FreeSans 960 0 0 0 io_oeb[17]
port 115 nsew signal tristate
flabel metal3 s -960 364428 480 364668 0 FreeSans 960 0 0 0 io_oeb[18]
port 116 nsew signal tristate
flabel metal3 s 583520 84268 584960 84508 0 FreeSans 960 0 0 0 io_oeb[19]
port 117 nsew signal tristate
flabel metal2 s 396050 703520 396162 704960 0 FreeSans 448 90 0 0 io_oeb[1]
port 118 nsew signal tristate
flabel metal3 s -960 271948 480 272188 0 FreeSans 960 0 0 0 io_oeb[20]
port 119 nsew signal tristate
flabel metal3 s -960 87668 480 87908 0 FreeSans 960 0 0 0 io_oeb[21]
port 120 nsew signal tristate
flabel metal3 s 583520 252908 584960 253148 0 FreeSans 960 0 0 0 io_oeb[22]
port 121 nsew signal tristate
flabel metal2 s 166786 -960 166898 480 0 FreeSans 448 90 0 0 io_oeb[23]
port 122 nsew signal tristate
flabel metal3 s -960 588828 480 589068 0 FreeSans 960 0 0 0 io_oeb[24]
port 123 nsew signal tristate
flabel metal2 s 330362 -960 330474 480 0 FreeSans 448 90 0 0 io_oeb[25]
port 124 nsew signal tristate
flabel metal3 s -960 400468 480 400708 0 FreeSans 960 0 0 0 io_oeb[26]
port 125 nsew signal tristate
flabel metal3 s -960 320228 480 320468 0 FreeSans 960 0 0 0 io_oeb[2]
port 126 nsew signal tristate
flabel metal2 s 148754 703520 148866 704960 0 FreeSans 448 90 0 0 io_oeb[3]
port 127 nsew signal tristate
flabel metal2 s 327142 703520 327254 704960 0 FreeSans 448 90 0 0 io_oeb[4]
port 128 nsew signal tristate
flabel metal3 s 583520 76788 584960 77028 0 FreeSans 960 0 0 0 io_oeb[5]
port 129 nsew signal tristate
flabel metal3 s -960 116228 480 116468 0 FreeSans 960 0 0 0 io_oeb[6]
port 130 nsew signal tristate
flabel metal2 s 144890 703520 145002 704960 0 FreeSans 448 90 0 0 io_oeb[7]
port 131 nsew signal tristate
flabel metal2 s 547390 703520 547502 704960 0 FreeSans 448 90 0 0 io_oeb[8]
port 132 nsew signal tristate
flabel metal2 s 128790 -960 128902 480 0 FreeSans 448 90 0 0 io_oeb[9]
port 133 nsew signal tristate
flabel metal3 s -960 23748 480 23988 0 FreeSans 960 0 0 0 io_out[0]
port 134 nsew signal tristate
flabel metal3 s -960 416788 480 417028 0 FreeSans 960 0 0 0 io_out[10]
port 135 nsew signal tristate
flabel metal2 s 512614 -960 512726 480 0 FreeSans 448 90 0 0 io_out[11]
port 136 nsew signal tristate
flabel metal3 s 583520 698308 584960 698548 0 FreeSans 960 0 0 0 io_out[12]
port 137 nsew signal tristate
flabel metal2 s 482990 703520 483102 704960 0 FreeSans 448 90 0 0 io_out[13]
port 138 nsew signal tristate
flabel metal2 s 182886 703520 182998 704960 0 FreeSans 448 90 0 0 io_out[14]
port 139 nsew signal tristate
flabel metal3 s 583520 673828 584960 674068 0 FreeSans 960 0 0 0 io_out[15]
port 140 nsew signal tristate
flabel metal3 s -960 296428 480 296668 0 FreeSans 960 0 0 0 io_out[16]
port 141 nsew signal tristate
flabel metal2 s 38630 703520 38742 704960 0 FreeSans 448 90 0 0 io_out[17]
port 142 nsew signal tristate
flabel metal2 s 570574 703520 570686 704960 0 FreeSans 448 90 0 0 io_out[18]
port 143 nsew signal tristate
flabel metal2 s 468178 703520 468290 704960 0 FreeSans 448 90 0 0 io_out[19]
port 144 nsew signal tristate
flabel metal3 s 583520 658188 584960 658428 0 FreeSans 960 0 0 0 io_out[1]
port 145 nsew signal tristate
flabel metal2 s 285926 703520 286038 704960 0 FreeSans 448 90 0 0 io_out[20]
port 146 nsew signal tristate
flabel metal3 s -960 637108 480 637348 0 FreeSans 960 0 0 0 io_out[21]
port 147 nsew signal tristate
flabel metal2 s 444994 703520 445106 704960 0 FreeSans 448 90 0 0 io_out[22]
port 148 nsew signal tristate
flabel metal3 s 583520 645948 584960 646188 0 FreeSans 960 0 0 0 io_out[23]
port 149 nsew signal tristate
flabel metal3 s -960 3348 480 3588 0 FreeSans 960 0 0 0 io_out[24]
port 150 nsew signal tristate
flabel metal3 s -960 436508 480 436748 0 FreeSans 960 0 0 0 io_out[25]
port 151 nsew signal tristate
flabel metal3 s 583520 60468 584960 60708 0 FreeSans 960 0 0 0 io_out[26]
port 152 nsew signal tristate
flabel metal3 s -960 504508 480 504748 0 FreeSans 960 0 0 0 io_out[2]
port 153 nsew signal tristate
flabel metal3 s 583520 337228 584960 337468 0 FreeSans 960 0 0 0 io_out[3]
port 154 nsew signal tristate
flabel metal3 s -960 701028 480 701268 0 FreeSans 960 0 0 0 io_out[4]
port 155 nsew signal tristate
flabel metal3 s -960 689468 480 689708 0 FreeSans 960 0 0 0 io_out[5]
port 156 nsew signal tristate
flabel metal3 s -960 452828 480 453068 0 FreeSans 960 0 0 0 io_out[6]
port 157 nsew signal tristate
flabel metal2 s 174514 -960 174626 480 0 FreeSans 448 90 0 0 io_out[7]
port 158 nsew signal tristate
flabel metal2 s 45070 -960 45182 480 0 FreeSans 448 90 0 0 io_out[8]
port 159 nsew signal tristate
flabel metal2 s 519698 -960 519810 480 0 FreeSans 448 90 0 0 io_out[9]
port 160 nsew signal tristate
flabel metal2 s 23818 703520 23930 704960 0 FreeSans 448 90 0 0 la_data_in[0]
port 161 nsew signal input
flabel metal3 s 583520 597668 584960 597908 0 FreeSans 960 0 0 0 la_data_in[100]
port 162 nsew signal input
flabel metal3 s -960 560948 480 561188 0 FreeSans 960 0 0 0 la_data_in[101]
port 163 nsew signal input
flabel metal3 s -960 380748 480 380988 0 FreeSans 960 0 0 0 la_data_in[102]
port 164 nsew signal input
flabel metal2 s 376730 703520 376842 704960 0 FreeSans 448 90 0 0 la_data_in[103]
port 165 nsew signal input
flabel metal2 s 269182 -960 269294 480 0 FreeSans 448 90 0 0 la_data_in[104]
port 166 nsew signal input
flabel metal3 s 583520 225028 584960 225268 0 FreeSans 960 0 0 0 la_data_in[105]
port 167 nsew signal input
flabel metal3 s 583520 8108 584960 8348 0 FreeSans 960 0 0 0 la_data_in[106]
port 168 nsew signal input
flabel metal3 s -960 624868 480 625108 0 FreeSans 960 0 0 0 la_data_in[107]
port 169 nsew signal input
flabel metal3 s -960 520828 480 521068 0 FreeSans 960 0 0 0 la_data_in[108]
port 170 nsew signal input
flabel metal2 s 485566 -960 485678 480 0 FreeSans 448 90 0 0 la_data_in[109]
port 171 nsew signal input
flabel metal3 s -960 47548 480 47788 0 FreeSans 960 0 0 0 la_data_in[10]
port 172 nsew signal input
flabel metal3 s 583520 529668 584960 529908 0 FreeSans 960 0 0 0 la_data_in[110]
port 173 nsew signal input
flabel metal3 s 583520 24428 584960 24668 0 FreeSans 960 0 0 0 la_data_in[111]
port 174 nsew signal input
flabel metal3 s -960 681308 480 681548 0 FreeSans 960 0 0 0 la_data_in[112]
port 175 nsew signal input
flabel metal3 s -960 184228 480 184468 0 FreeSans 960 0 0 0 la_data_in[113]
port 176 nsew signal input
flabel metal2 s 314906 -960 315018 480 0 FreeSans 448 90 0 0 la_data_in[114]
port 177 nsew signal input
flabel metal3 s 583520 389588 584960 389828 0 FreeSans 960 0 0 0 la_data_in[115]
port 178 nsew signal input
flabel metal3 s -960 180148 480 180388 0 FreeSans 960 0 0 0 la_data_in[116]
port 179 nsew signal input
flabel metal2 s 121062 -960 121174 480 0 FreeSans 448 90 0 0 la_data_in[117]
port 180 nsew signal input
flabel metal3 s -960 512668 480 512908 0 FreeSans 960 0 0 0 la_data_in[118]
port 181 nsew signal input
flabel metal2 s 447570 -960 447682 480 0 FreeSans 448 90 0 0 la_data_in[119]
port 182 nsew signal input
flabel metal2 s 535154 -960 535266 480 0 FreeSans 448 90 0 0 la_data_in[11]
port 183 nsew signal input
flabel metal3 s 583520 301188 584960 301428 0 FreeSans 960 0 0 0 la_data_in[120]
port 184 nsew signal input
flabel metal2 s 342598 703520 342710 704960 0 FreeSans 448 90 0 0 la_data_in[121]
port 185 nsew signal input
flabel metal3 s -960 484788 480 485028 0 FreeSans 960 0 0 0 la_data_in[122]
port 186 nsew signal input
flabel metal3 s 583520 493628 584960 493868 0 FreeSans 960 0 0 0 la_data_in[123]
port 187 nsew signal input
flabel metal2 s 244066 703520 244178 704960 0 FreeSans 448 90 0 0 la_data_in[124]
port 188 nsew signal input
flabel metal2 s 162922 -960 163034 480 0 FreeSans 448 90 0 0 la_data_in[125]
port 189 nsew signal input
flabel metal3 s -960 621468 480 621708 0 FreeSans 960 0 0 0 la_data_in[126]
port 190 nsew signal input
flabel metal3 s 583520 269228 584960 269468 0 FreeSans 960 0 0 0 la_data_in[127]
port 191 nsew signal input
flabel metal3 s -960 444668 480 444908 0 FreeSans 960 0 0 0 la_data_in[12]
port 192 nsew signal input
flabel metal2 s 489430 -960 489542 480 0 FreeSans 448 90 0 0 la_data_in[13]
port 193 nsew signal input
flabel metal3 s 583520 589508 584960 589748 0 FreeSans 960 0 0 0 la_data_in[14]
port 194 nsew signal input
flabel metal3 s 583520 626228 584960 626468 0 FreeSans 960 0 0 0 la_data_in[15]
port 195 nsew signal input
flabel metal3 s 583520 425628 584960 425868 0 FreeSans 960 0 0 0 la_data_in[16]
port 196 nsew signal input
flabel metal2 s 261454 -960 261566 480 0 FreeSans 448 90 0 0 la_data_in[17]
port 197 nsew signal input
flabel metal3 s 583520 553468 584960 553708 0 FreeSans 960 0 0 0 la_data_in[18]
port 198 nsew signal input
flabel metal3 s -960 544628 480 544868 0 FreeSans 960 0 0 0 la_data_in[19]
port 199 nsew signal input
flabel metal2 s 477838 -960 477950 480 0 FreeSans 448 90 0 0 la_data_in[1]
port 200 nsew signal input
flabel metal3 s -960 163828 480 164068 0 FreeSans 960 0 0 0 la_data_in[20]
port 201 nsew signal input
flabel metal3 s 583520 108748 584960 108988 0 FreeSans 960 0 0 0 la_data_in[21]
port 202 nsew signal input
flabel metal3 s -960 344708 480 344948 0 FreeSans 960 0 0 0 la_data_in[22]
port 203 nsew signal input
flabel metal2 s 303314 -960 303426 480 0 FreeSans 448 90 0 0 la_data_in[23]
port 204 nsew signal input
flabel metal2 s 517122 703520 517234 704960 0 FreeSans 448 90 0 0 la_data_in[24]
port 205 nsew signal input
flabel metal3 s 583520 188988 584960 189228 0 FreeSans 960 0 0 0 la_data_in[25]
port 206 nsew signal input
flabel metal2 s 463026 -960 463138 480 0 FreeSans 448 90 0 0 la_data_in[26]
port 207 nsew signal input
flabel metal3 s -960 697628 480 697868 0 FreeSans 960 0 0 0 la_data_in[27]
port 208 nsew signal input
flabel metal2 s 528714 703520 528826 704960 0 FreeSans 448 90 0 0 la_data_in[28]
port 209 nsew signal input
flabel metal3 s -960 605148 480 605388 0 FreeSans 960 0 0 0 la_data_in[29]
port 210 nsew signal input
flabel metal3 s -960 304588 480 304828 0 FreeSans 960 0 0 0 la_data_in[2]
port 211 nsew signal input
flabel metal2 s 295586 -960 295698 480 0 FreeSans 448 90 0 0 la_data_in[30]
port 212 nsew signal input
flabel metal3 s -960 456908 480 457148 0 FreeSans 960 0 0 0 la_data_in[31]
port 213 nsew signal input
flabel metal2 s 75338 -960 75450 480 0 FreeSans 448 90 0 0 la_data_in[32]
port 214 nsew signal input
flabel metal2 s 175802 703520 175914 704960 0 FreeSans 448 90 0 0 la_data_in[33]
port 215 nsew signal input
flabel metal2 s 304602 703520 304714 704960 0 FreeSans 448 90 0 0 la_data_in[34]
port 216 nsew signal input
flabel metal3 s -960 332468 480 332708 0 FreeSans 960 0 0 0 la_data_in[35]
port 217 nsew signal input
flabel metal3 s -960 657508 480 657748 0 FreeSans 960 0 0 0 la_data_in[36]
port 218 nsew signal input
flabel metal3 s 583520 521508 584960 521748 0 FreeSans 960 0 0 0 la_data_in[37]
port 219 nsew signal input
flabel metal3 s 583520 453508 584960 453748 0 FreeSans 960 0 0 0 la_data_in[38]
port 220 nsew signal input
flabel metal3 s -960 159748 480 159988 0 FreeSans 960 0 0 0 la_data_in[39]
port 221 nsew signal input
flabel metal2 s 546746 -960 546858 480 0 FreeSans 448 90 0 0 la_data_in[3]
port 222 nsew signal input
flabel metal2 s 540306 703520 540418 704960 0 FreeSans 448 90 0 0 la_data_in[40]
port 223 nsew signal input
flabel metal3 s 583520 52308 584960 52548 0 FreeSans 960 0 0 0 la_data_in[41]
port 224 nsew signal input
flabel metal3 s 583520 365108 584960 365348 0 FreeSans 960 0 0 0 la_data_in[42]
port 225 nsew signal input
flabel metal3 s -960 76108 480 76348 0 FreeSans 960 0 0 0 la_data_in[43]
port 226 nsew signal input
flabel metal3 s -960 7428 480 7668 0 FreeSans 960 0 0 0 la_data_in[44]
port 227 nsew signal input
flabel metal2 s 204782 -960 204894 480 0 FreeSans 448 90 0 0 la_data_in[45]
port 228 nsew signal input
flabel metal3 s -960 144108 480 144348 0 FreeSans 960 0 0 0 la_data_in[46]
port 229 nsew signal input
flabel metal3 s 583520 40748 584960 40988 0 FreeSans 960 0 0 0 la_data_in[47]
port 230 nsew signal input
flabel metal2 s 151330 -960 151442 480 0 FreeSans 448 90 0 0 la_data_in[48]
port 231 nsew signal input
flabel metal2 s 197054 -960 197166 480 0 FreeSans 448 90 0 0 la_data_in[49]
port 232 nsew signal input
flabel metal3 s 583520 313428 584960 313668 0 FreeSans 960 0 0 0 la_data_in[4]
port 233 nsew signal input
flabel metal2 s 580878 -960 580990 480 0 FreeSans 448 90 0 0 la_data_in[50]
port 234 nsew signal input
flabel metal2 s 266606 703520 266718 704960 0 FreeSans 448 90 0 0 la_data_in[51]
port 235 nsew signal input
flabel metal3 s -960 428348 480 428588 0 FreeSans 960 0 0 0 la_data_in[52]
port 236 nsew signal input
flabel metal3 s -960 123708 480 123948 0 FreeSans 960 0 0 0 la_data_in[53]
port 237 nsew signal input
flabel metal2 s 262742 703520 262854 704960 0 FreeSans 448 90 0 0 la_data_in[54]
port 238 nsew signal input
flabel metal3 s 583520 509948 584960 510188 0 FreeSans 960 0 0 0 la_data_in[55]
port 239 nsew signal input
flabel metal3 s -960 548708 480 548948 0 FreeSans 960 0 0 0 la_data_in[56]
port 240 nsew signal input
flabel metal2 s 257590 -960 257702 480 0 FreeSans 448 90 0 0 la_data_in[57]
port 241 nsew signal input
flabel metal2 s 3210 -960 3322 480 0 FreeSans 448 90 0 0 la_data_in[58]
port 242 nsew signal input
flabel metal3 s 583520 441268 584960 441508 0 FreeSans 960 0 0 0 la_data_in[59]
port 243 nsew signal input
flabel metal3 s 583520 32588 584960 32828 0 FreeSans 960 0 0 0 la_data_in[5]
port 244 nsew signal input
flabel metal2 s 57950 703520 58062 704960 0 FreeSans 448 90 0 0 la_data_in[60]
port 245 nsew signal input
flabel metal3 s 583520 501788 584960 502028 0 FreeSans 960 0 0 0 la_data_in[61]
port 246 nsew signal input
flabel metal3 s -960 95828 480 96068 0 FreeSans 960 0 0 0 la_data_in[62]
port 247 nsew signal input
flabel metal3 s -960 488868 480 489108 0 FreeSans 960 0 0 0 la_data_in[63]
port 248 nsew signal input
flabel metal3 s -960 528988 480 529228 0 FreeSans 960 0 0 0 la_data_in[64]
port 249 nsew signal input
flabel metal3 s -960 677228 480 677468 0 FreeSans 960 0 0 0 la_data_in[65]
port 250 nsew signal input
flabel metal3 s 583520 56388 584960 56628 0 FreeSans 960 0 0 0 la_data_in[66]
port 251 nsew signal input
flabel metal2 s 448858 703520 448970 704960 0 FreeSans 448 90 0 0 la_data_in[67]
port 252 nsew signal input
flabel metal3 s 583520 180828 584960 181068 0 FreeSans 960 0 0 0 la_data_in[68]
port 253 nsew signal input
flabel metal3 s 583520 586108 584960 586348 0 FreeSans 960 0 0 0 la_data_in[69]
port 254 nsew signal input
flabel metal3 s 583520 341308 584960 341548 0 FreeSans 960 0 0 0 la_data_in[6]
port 255 nsew signal input
flabel metal2 s 79202 -960 79314 480 0 FreeSans 448 90 0 0 la_data_in[70]
port 256 nsew signal input
flabel metal3 s 583520 573868 584960 574108 0 FreeSans 960 0 0 0 la_data_in[71]
port 257 nsew signal input
flabel metal3 s -960 308668 480 308908 0 FreeSans 960 0 0 0 la_data_in[72]
port 258 nsew signal input
flabel metal2 s 118486 703520 118598 704960 0 FreeSans 448 90 0 0 la_data_in[73]
port 259 nsew signal input
flabel metal3 s 583520 549388 584960 549628 0 FreeSans 960 0 0 0 la_data_in[74]
port 260 nsew signal input
flabel metal2 s 392186 703520 392298 704960 0 FreeSans 448 90 0 0 la_data_in[75]
port 261 nsew signal input
flabel metal2 s 520986 703520 521098 704960 0 FreeSans 448 90 0 0 la_data_in[76]
port 262 nsew signal input
flabel metal3 s -960 288268 480 288508 0 FreeSans 960 0 0 0 la_data_in[77]
port 263 nsew signal input
flabel metal3 s 583520 333148 584960 333388 0 FreeSans 960 0 0 0 la_data_in[78]
port 264 nsew signal input
flabel metal3 s 583520 677908 584960 678148 0 FreeSans 960 0 0 0 la_data_in[79]
port 265 nsew signal input
flabel metal2 s 194478 703520 194590 704960 0 FreeSans 448 90 0 0 la_data_in[7]
port 266 nsew signal input
flabel metal2 s 494582 703520 494694 704960 0 FreeSans 448 90 0 0 la_data_in[80]
port 267 nsew signal input
flabel metal2 s 232474 703520 232586 704960 0 FreeSans 448 90 0 0 la_data_in[81]
port 268 nsew signal input
flabel metal3 s -960 480708 480 480948 0 FreeSans 960 0 0 0 la_data_in[82]
port 269 nsew signal input
flabel metal3 s -960 72028 480 72268 0 FreeSans 960 0 0 0 la_data_in[83]
port 270 nsew signal input
flabel metal2 s 490718 703520 490830 704960 0 FreeSans 448 90 0 0 la_data_in[84]
port 271 nsew signal input
flabel metal3 s -960 328388 480 328628 0 FreeSans 960 0 0 0 la_data_in[85]
port 272 nsew signal input
flabel metal3 s 583520 349468 584960 349708 0 FreeSans 960 0 0 0 la_data_in[86]
port 273 nsew signal input
flabel metal3 s -960 91748 480 91988 0 FreeSans 960 0 0 0 la_data_in[87]
port 274 nsew signal input
flabel metal3 s 583520 628 584960 868 0 FreeSans 960 0 0 0 la_data_in[88]
port 275 nsew signal input
flabel metal3 s -960 284188 480 284428 0 FreeSans 960 0 0 0 la_data_in[89]
port 276 nsew signal input
flabel metal3 s -960 103988 480 104228 0 FreeSans 960 0 0 0 la_data_in[8]
port 277 nsew signal input
flabel metal2 s 94658 -960 94770 480 0 FreeSans 448 90 0 0 la_data_in[90]
port 278 nsew signal input
flabel metal3 s -960 195788 480 196028 0 FreeSans 960 0 0 0 la_data_in[91]
port 279 nsew signal input
flabel metal2 s 254370 -960 254482 480 0 FreeSans 448 90 0 0 la_data_in[92]
port 280 nsew signal input
flabel metal2 s 276910 -960 277022 480 0 FreeSans 448 90 0 0 la_data_in[93]
port 281 nsew signal input
flabel metal2 s 50222 703520 50334 704960 0 FreeSans 448 90 0 0 la_data_in[94]
port 282 nsew signal input
flabel metal2 s 553830 -960 553942 480 0 FreeSans 448 90 0 0 la_data_in[95]
port 283 nsew signal input
flabel metal2 s 555118 703520 555230 704960 0 FreeSans 448 90 0 0 la_data_in[96]
port 284 nsew signal input
flabel metal3 s -960 232508 480 232748 0 FreeSans 960 0 0 0 la_data_in[97]
port 285 nsew signal input
flabel metal3 s 583520 320908 584960 321148 0 FreeSans 960 0 0 0 la_data_in[98]
port 286 nsew signal input
flabel metal2 s 189326 -960 189438 480 0 FreeSans 448 90 0 0 la_data_in[99]
port 287 nsew signal input
flabel metal3 s -960 508588 480 508828 0 FreeSans 960 0 0 0 la_data_in[9]
port 288 nsew signal input
flabel metal3 s -960 609228 480 609468 0 FreeSans 960 0 0 0 la_data_out[0]
port 289 nsew signal tristate
flabel metal2 s 284638 -960 284750 480 0 FreeSans 448 90 0 0 la_data_out[100]
port 290 nsew signal tristate
flabel metal3 s 583520 197148 584960 197388 0 FreeSans 960 0 0 0 la_data_out[101]
port 291 nsew signal tristate
flabel metal3 s 583520 413388 584960 413628 0 FreeSans 960 0 0 0 la_data_out[102]
port 292 nsew signal tristate
flabel metal3 s -960 685388 480 685628 0 FreeSans 960 0 0 0 la_data_out[103]
port 293 nsew signal tristate
flabel metal3 s -960 645268 480 645508 0 FreeSans 960 0 0 0 la_data_out[104]
port 294 nsew signal tristate
flabel metal2 s 231186 -960 231298 480 0 FreeSans 448 90 0 0 la_data_out[105]
port 295 nsew signal tristate
flabel metal2 s 164210 703520 164322 704960 0 FreeSans 448 90 0 0 la_data_out[106]
port 296 nsew signal tristate
flabel metal3 s 583520 261068 584960 261308 0 FreeSans 960 0 0 0 la_data_out[107]
port 297 nsew signal tristate
flabel metal2 s 156482 703520 156594 704960 0 FreeSans 448 90 0 0 la_data_out[108]
port 298 nsew signal tristate
flabel metal2 s 84354 703520 84466 704960 0 FreeSans 448 90 0 0 la_data_out[109]
port 299 nsew signal tristate
flabel metal2 s 155194 -960 155306 480 0 FreeSans 448 90 0 0 la_data_out[10]
port 300 nsew signal tristate
flabel metal3 s 583520 392988 584960 393228 0 FreeSans 960 0 0 0 la_data_out[110]
port 301 nsew signal tristate
flabel metal3 s -960 465068 480 465308 0 FreeSans 960 0 0 0 la_data_out[111]
port 302 nsew signal tristate
flabel metal2 s 502310 703520 502422 704960 0 FreeSans 448 90 0 0 la_data_out[112]
port 303 nsew signal tristate
flabel metal3 s -960 384828 480 385068 0 FreeSans 960 0 0 0 la_data_out[113]
port 304 nsew signal tristate
flabel metal3 s -960 212108 480 212348 0 FreeSans 960 0 0 0 la_data_out[114]
port 305 nsew signal tristate
flabel metal2 s 566710 703520 566822 704960 0 FreeSans 448 90 0 0 la_data_out[115]
port 306 nsew signal tristate
flabel metal3 s -960 497028 480 497268 0 FreeSans 960 0 0 0 la_data_out[116]
port 307 nsew signal tristate
flabel metal2 s 200918 -960 201030 480 0 FreeSans 448 90 0 0 la_data_out[117]
port 308 nsew signal tristate
flabel metal2 s 562846 703520 562958 704960 0 FreeSans 448 90 0 0 la_data_out[118]
port 309 nsew signal tristate
flabel metal3 s -960 67948 480 68188 0 FreeSans 960 0 0 0 la_data_out[119]
port 310 nsew signal tristate
flabel metal2 s 409574 -960 409686 480 0 FreeSans 448 90 0 0 la_data_out[11]
port 311 nsew signal tristate
flabel metal3 s 583520 654108 584960 654348 0 FreeSans 960 0 0 0 la_data_out[120]
port 312 nsew signal tristate
flabel metal3 s 583520 401148 584960 401388 0 FreeSans 960 0 0 0 la_data_out[121]
port 313 nsew signal tristate
flabel metal3 s 583520 28508 584960 28748 0 FreeSans 960 0 0 0 la_data_out[122]
port 314 nsew signal tristate
flabel metal3 s -960 188308 480 188548 0 FreeSans 960 0 0 0 la_data_out[123]
port 315 nsew signal tristate
flabel metal2 s 18666 -960 18778 480 0 FreeSans 448 90 0 0 la_data_out[124]
port 316 nsew signal tristate
flabel metal2 s 179022 703520 179134 704960 0 FreeSans 448 90 0 0 la_data_out[125]
port 317 nsew signal tristate
flabel metal2 s 106894 703520 107006 704960 0 FreeSans 448 90 0 0 la_data_out[126]
port 318 nsew signal tristate
flabel metal2 s 475262 703520 475374 704960 0 FreeSans 448 90 0 0 la_data_out[127]
port 319 nsew signal tristate
flabel metal3 s 583520 140708 584960 140948 0 FreeSans 960 0 0 0 la_data_out[12]
port 320 nsew signal tristate
flabel metal3 s 583520 489548 584960 489788 0 FreeSans 960 0 0 0 la_data_out[13]
port 321 nsew signal tristate
flabel metal3 s -960 27828 480 28068 0 FreeSans 960 0 0 0 la_data_out[14]
port 322 nsew signal tristate
flabel metal3 s 583520 284868 584960 285108 0 FreeSans 960 0 0 0 la_data_out[15]
port 323 nsew signal tristate
flabel metal2 s 227322 -960 227434 480 0 FreeSans 448 90 0 0 la_data_out[16]
port 324 nsew signal tristate
flabel metal3 s 583520 44148 584960 44388 0 FreeSans 960 0 0 0 la_data_out[17]
port 325 nsew signal tristate
flabel metal2 s 394762 -960 394874 480 0 FreeSans 448 90 0 0 la_data_out[18]
port 326 nsew signal tristate
flabel metal2 s 88218 703520 88330 704960 0 FreeSans 448 90 0 0 la_data_out[19]
port 327 nsew signal tristate
flabel metal2 s 334870 703520 334982 704960 0 FreeSans 448 90 0 0 la_data_out[1]
port 328 nsew signal tristate
flabel metal2 s 168074 703520 168186 704960 0 FreeSans 448 90 0 0 la_data_out[20]
port 329 nsew signal tristate
flabel metal2 s 110114 -960 110226 480 0 FreeSans 448 90 0 0 la_data_out[21]
port 330 nsew signal tristate
flabel metal3 s 583520 469828 584960 470068 0 FreeSans 960 0 0 0 la_data_out[22]
port 331 nsew signal tristate
flabel metal3 s -960 448748 480 448988 0 FreeSans 960 0 0 0 la_data_out[23]
port 332 nsew signal tristate
flabel metal2 s 504886 -960 504998 480 0 FreeSans 448 90 0 0 la_data_out[24]
port 333 nsew signal tristate
flabel metal3 s 583520 233188 584960 233428 0 FreeSans 960 0 0 0 la_data_out[25]
port 334 nsew signal tristate
flabel metal2 s 582166 703520 582278 704960 0 FreeSans 448 90 0 0 la_data_out[26]
port 335 nsew signal tristate
flabel metal3 s -960 440588 480 440828 0 FreeSans 960 0 0 0 la_data_out[27]
port 336 nsew signal tristate
flabel metal3 s 583520 16268 584960 16508 0 FreeSans 960 0 0 0 la_data_out[28]
port 337 nsew signal tristate
flabel metal2 s 472042 703520 472154 704960 0 FreeSans 448 90 0 0 la_data_out[29]
port 338 nsew signal tristate
flabel metal3 s 583520 477308 584960 477548 0 FreeSans 960 0 0 0 la_data_out[2]
port 339 nsew signal tristate
flabel metal3 s 583520 377348 584960 377588 0 FreeSans 960 0 0 0 la_data_out[30]
port 340 nsew signal tristate
flabel metal2 s 311042 -960 311154 480 0 FreeSans 448 90 0 0 la_data_out[31]
port 341 nsew signal tristate
flabel metal2 s 307178 -960 307290 480 0 FreeSans 448 90 0 0 la_data_out[32]
port 342 nsew signal tristate
flabel metal3 s -960 412708 480 412948 0 FreeSans 960 0 0 0 la_data_out[33]
port 343 nsew signal tristate
flabel metal3 s 583520 433108 584960 433348 0 FreeSans 960 0 0 0 la_data_out[34]
port 344 nsew signal tristate
flabel metal3 s -960 235908 480 236148 0 FreeSans 960 0 0 0 la_data_out[35]
port 345 nsew signal tristate
flabel metal3 s 583520 316828 584960 317068 0 FreeSans 960 0 0 0 la_data_out[36]
port 346 nsew signal tristate
flabel metal3 s 583520 208708 584960 208948 0 FreeSans 960 0 0 0 la_data_out[37]
port 347 nsew signal tristate
flabel metal3 s -960 127788 480 128028 0 FreeSans 960 0 0 0 la_data_out[38]
port 348 nsew signal tristate
flabel metal3 s 583520 157028 584960 157268 0 FreeSans 960 0 0 0 la_data_out[39]
port 349 nsew signal tristate
flabel metal2 s 524850 703520 524962 704960 0 FreeSans 448 90 0 0 la_data_out[3]
port 350 nsew signal tristate
flabel metal3 s 583520 12188 584960 12428 0 FreeSans 960 0 0 0 la_data_out[40]
port 351 nsew signal tristate
flabel metal3 s 583520 72708 584960 72948 0 FreeSans 960 0 0 0 la_data_out[41]
port 352 nsew signal tristate
flabel metal3 s 583520 132548 584960 132788 0 FreeSans 960 0 0 0 la_data_out[42]
port 353 nsew signal tristate
flabel metal2 s 251794 703520 251906 704960 0 FreeSans 448 90 0 0 la_data_out[43]
port 354 nsew signal tristate
flabel metal3 s 583520 353548 584960 353788 0 FreeSans 960 0 0 0 la_data_out[44]
port 355 nsew signal tristate
flabel metal2 s 322634 -960 322746 480 0 FreeSans 448 90 0 0 la_data_out[45]
port 356 nsew signal tristate
flabel metal2 s 240202 703520 240314 704960 0 FreeSans 448 90 0 0 la_data_out[46]
port 357 nsew signal tristate
flabel metal3 s -960 633028 480 633268 0 FreeSans 960 0 0 0 la_data_out[47]
port 358 nsew signal tristate
flabel metal2 s 470754 -960 470866 480 0 FreeSans 448 90 0 0 la_data_out[48]
port 359 nsew signal tristate
flabel metal2 s 379306 -960 379418 480 0 FreeSans 448 90 0 0 la_data_out[49]
port 360 nsew signal tristate
flabel metal2 s 80490 703520 80602 704960 0 FreeSans 448 90 0 0 la_data_out[4]
port 361 nsew signal tristate
flabel metal2 s 61814 703520 61926 704960 0 FreeSans 448 90 0 0 la_data_out[50]
port 362 nsew signal tristate
flabel metal3 s -960 516748 480 516988 0 FreeSans 960 0 0 0 la_data_out[51]
port 363 nsew signal tristate
flabel metal2 s 141670 703520 141782 704960 0 FreeSans 448 90 0 0 la_data_out[52]
port 364 nsew signal tristate
flabel metal3 s -960 228428 480 228668 0 FreeSans 960 0 0 0 la_data_out[53]
port 365 nsew signal tristate
flabel metal3 s -960 352188 480 352428 0 FreeSans 960 0 0 0 la_data_out[54]
port 366 nsew signal tristate
flabel metal2 s 371578 -960 371690 480 0 FreeSans 448 90 0 0 la_data_out[55]
port 367 nsew signal tristate
flabel metal3 s -960 83588 480 83828 0 FreeSans 960 0 0 0 la_data_out[56]
port 368 nsew signal tristate
flabel metal2 s 434046 703520 434158 704960 0 FreeSans 448 90 0 0 la_data_out[57]
port 369 nsew signal tristate
flabel metal2 s 398626 -960 398738 480 0 FreeSans 448 90 0 0 la_data_out[58]
port 370 nsew signal tristate
flabel metal3 s -960 199868 480 200108 0 FreeSans 960 0 0 0 la_data_out[59]
port 371 nsew signal tristate
flabel metal2 s 274334 703520 274446 704960 0 FreeSans 448 90 0 0 la_data_out[5]
port 372 nsew signal tristate
flabel metal3 s 583520 449428 584960 449668 0 FreeSans 960 0 0 0 la_data_out[60]
port 373 nsew signal tristate
flabel metal3 s 583520 128468 584960 128708 0 FreeSans 960 0 0 0 la_data_out[61]
port 374 nsew signal tristate
flabel metal3 s 583520 429708 584960 429948 0 FreeSans 960 0 0 0 la_data_out[62]
port 375 nsew signal tristate
flabel metal2 s 356766 -960 356878 480 0 FreeSans 448 90 0 0 la_data_out[63]
port 376 nsew signal tristate
flabel metal3 s -960 641188 480 641428 0 FreeSans 960 0 0 0 la_data_out[64]
port 377 nsew signal tristate
flabel metal2 s 452722 703520 452834 704960 0 FreeSans 448 90 0 0 la_data_out[65]
port 378 nsew signal tristate
flabel metal2 s 364494 -960 364606 480 0 FreeSans 448 90 0 0 la_data_out[66]
port 379 nsew signal tristate
flabel metal2 s 430182 703520 430294 704960 0 FreeSans 448 90 0 0 la_data_out[67]
port 380 nsew signal tristate
flabel metal3 s -960 468468 480 468708 0 FreeSans 960 0 0 0 la_data_out[68]
port 381 nsew signal tristate
flabel metal2 s 527426 -960 527538 480 0 FreeSans 448 90 0 0 la_data_out[69]
port 382 nsew signal tristate
flabel metal3 s -960 537148 480 537388 0 FreeSans 960 0 0 0 la_data_out[6]
port 383 nsew signal tristate
flabel metal2 s 190614 703520 190726 704960 0 FreeSans 448 90 0 0 la_data_out[70]
port 384 nsew signal tristate
flabel metal3 s 583520 244748 584960 244988 0 FreeSans 960 0 0 0 la_data_out[71]
port 385 nsew signal tristate
flabel metal3 s 583520 184908 584960 185148 0 FreeSans 960 0 0 0 la_data_out[72]
port 386 nsew signal tristate
flabel metal2 s 318770 -960 318882 480 0 FreeSans 448 90 0 0 la_data_out[73]
port 387 nsew signal tristate
flabel metal2 s 474618 -960 474730 480 0 FreeSans 448 90 0 0 la_data_out[74]
port 388 nsew signal tristate
flabel metal2 s 246642 -960 246754 480 0 FreeSans 448 90 0 0 la_data_out[75]
port 389 nsew signal tristate
flabel metal2 s 437266 703520 437378 704960 0 FreeSans 448 90 0 0 la_data_out[76]
port 390 nsew signal tristate
flabel metal2 s 360630 -960 360742 480 0 FreeSans 448 90 0 0 la_data_out[77]
port 391 nsew signal tristate
flabel metal2 s 634 703520 746 704960 0 FreeSans 448 90 0 0 la_data_out[78]
port 392 nsew signal tristate
flabel metal3 s -960 460988 480 461228 0 FreeSans 960 0 0 0 la_data_out[79]
port 393 nsew signal tristate
flabel metal3 s -960 664988 480 665228 0 FreeSans 960 0 0 0 la_data_out[7]
port 394 nsew signal tristate
flabel metal3 s 583520 481388 584960 481628 0 FreeSans 960 0 0 0 la_data_out[80]
port 395 nsew signal tristate
flabel metal2 s 333582 -960 333694 480 0 FreeSans 448 90 0 0 la_data_out[81]
port 396 nsew signal tristate
flabel metal3 s 583520 152948 584960 153188 0 FreeSans 960 0 0 0 la_data_out[82]
port 397 nsew signal tristate
flabel metal3 s 583520 48228 584960 48468 0 FreeSans 960 0 0 0 la_data_out[83]
port 398 nsew signal tristate
flabel metal3 s 583520 237268 584960 237508 0 FreeSans 960 0 0 0 la_data_out[84]
port 399 nsew signal tristate
flabel metal3 s -960 569108 480 569348 0 FreeSans 960 0 0 0 la_data_out[85]
port 400 nsew signal tristate
flabel metal2 s 250506 -960 250618 480 0 FreeSans 448 90 0 0 la_data_out[86]
port 401 nsew signal tristate
flabel metal3 s -960 59788 480 60028 0 FreeSans 960 0 0 0 la_data_out[87]
port 402 nsew signal tristate
flabel metal2 s 466890 -960 467002 480 0 FreeSans 448 90 0 0 la_data_out[88]
port 403 nsew signal tristate
flabel metal2 s 513258 703520 513370 704960 0 FreeSans 448 90 0 0 la_data_out[89]
port 404 nsew signal tristate
flabel metal2 s 110758 703520 110870 704960 0 FreeSans 448 90 0 0 la_data_out[8]
port 405 nsew signal tristate
flabel metal3 s -960 280108 480 280348 0 FreeSans 960 0 0 0 la_data_out[90]
port 406 nsew signal tristate
flabel metal3 s -960 112148 480 112388 0 FreeSans 960 0 0 0 la_data_out[91]
port 407 nsew signal tristate
flabel metal3 s 583520 80868 584960 81108 0 FreeSans 960 0 0 0 la_data_out[92]
port 408 nsew signal tristate
flabel metal2 s 42494 703520 42606 704960 0 FreeSans 448 90 0 0 la_data_out[93]
port 409 nsew signal tristate
flabel metal2 s 220882 703520 220994 704960 0 FreeSans 448 90 0 0 la_data_out[94]
port 410 nsew signal tristate
flabel metal2 s 425030 -960 425142 480 0 FreeSans 448 90 0 0 la_data_out[95]
port 411 nsew signal tristate
flabel metal3 s -960 368508 480 368748 0 FreeSans 960 0 0 0 la_data_out[96]
port 412 nsew signal tristate
flabel metal3 s -960 208028 480 208268 0 FreeSans 960 0 0 0 la_data_out[97]
port 413 nsew signal tristate
flabel metal2 s 497158 -960 497270 480 0 FreeSans 448 90 0 0 la_data_out[98]
port 414 nsew signal tristate
flabel metal2 s 561558 -960 561670 480 0 FreeSans 448 90 0 0 la_data_out[99]
port 415 nsew signal tristate
flabel metal2 s 4498 703520 4610 704960 0 FreeSans 448 90 0 0 la_data_out[9]
port 416 nsew signal tristate
flabel metal2 s 76626 703520 76738 704960 0 FreeSans 448 90 0 0 la_oenb[0]
port 417 nsew signal input
flabel metal2 s 551254 703520 551366 704960 0 FreeSans 448 90 0 0 la_oenb[100]
port 418 nsew signal input
flabel metal2 s 515834 -960 515946 480 0 FreeSans 448 90 0 0 la_oenb[101]
port 419 nsew signal input
flabel metal2 s 12226 703520 12338 704960 0 FreeSans 448 90 0 0 la_oenb[102]
port 420 nsew signal input
flabel metal2 s 422454 703520 422566 704960 0 FreeSans 448 90 0 0 la_oenb[103]
port 421 nsew signal input
flabel metal2 s 403134 703520 403246 704960 0 FreeSans 448 90 0 0 la_oenb[104]
port 422 nsew signal input
flabel metal3 s -960 476628 480 476868 0 FreeSans 960 0 0 0 la_oenb[105]
port 423 nsew signal input
flabel metal2 s 299450 -960 299562 480 0 FreeSans 448 90 0 0 la_oenb[106]
port 424 nsew signal input
flabel metal2 s 352902 -960 353014 480 0 FreeSans 448 90 0 0 la_oenb[107]
port 425 nsew signal input
flabel metal2 s 532578 703520 532690 704960 0 FreeSans 448 90 0 0 la_oenb[108]
port 426 nsew signal input
flabel metal3 s 583520 164508 584960 164748 0 FreeSans 960 0 0 0 la_oenb[109]
port 427 nsew signal input
flabel metal2 s 418590 703520 418702 704960 0 FreeSans 448 90 0 0 la_oenb[10]
port 428 nsew signal input
flabel metal2 s 170650 -960 170762 480 0 FreeSans 448 90 0 0 la_oenb[110]
port 429 nsew signal input
flabel metal3 s 583520 473228 584960 473468 0 FreeSans 960 0 0 0 la_oenb[111]
port 430 nsew signal input
flabel metal2 s 171938 703520 172050 704960 0 FreeSans 448 90 0 0 la_oenb[112]
port 431 nsew signal input
flabel metal2 s 510038 703520 510150 704960 0 FreeSans 448 90 0 0 la_oenb[113]
port 432 nsew signal input
flabel metal2 s 137806 703520 137918 704960 0 FreeSans 448 90 0 0 la_oenb[114]
port 433 nsew signal input
flabel metal2 s 31546 703520 31658 704960 0 FreeSans 448 90 0 0 la_oenb[115]
port 434 nsew signal input
flabel metal2 s 380594 703520 380706 704960 0 FreeSans 448 90 0 0 la_oenb[116]
port 435 nsew signal input
flabel metal3 s -960 324308 480 324548 0 FreeSans 960 0 0 0 la_oenb[117]
port 436 nsew signal input
flabel metal3 s 583520 601748 584960 601988 0 FreeSans 960 0 0 0 la_oenb[118]
port 437 nsew signal input
flabel metal2 s 481702 -960 481814 480 0 FreeSans 448 90 0 0 la_oenb[119]
port 438 nsew signal input
flabel metal3 s 583520 437188 584960 437428 0 FreeSans 960 0 0 0 la_oenb[11]
port 439 nsew signal input
flabel metal2 s 124926 -960 125038 480 0 FreeSans 448 90 0 0 la_oenb[120]
port 440 nsew signal input
flabel metal3 s -960 79508 480 79748 0 FreeSans 960 0 0 0 la_oenb[121]
port 441 nsew signal input
flabel metal3 s -960 432428 480 432668 0 FreeSans 960 0 0 0 la_oenb[122]
port 442 nsew signal input
flabel metal2 s 341310 -960 341422 480 0 FreeSans 448 90 0 0 la_oenb[123]
port 443 nsew signal input
flabel metal2 s 558982 703520 559094 704960 0 FreeSans 448 90 0 0 la_oenb[124]
port 444 nsew signal input
flabel metal3 s -960 376668 480 376908 0 FreeSans 960 0 0 0 la_oenb[125]
port 445 nsew signal input
flabel metal3 s -960 336548 480 336788 0 FreeSans 960 0 0 0 la_oenb[126]
port 446 nsew signal input
flabel metal2 s 8362 703520 8474 704960 0 FreeSans 448 90 0 0 la_oenb[127]
port 447 nsew signal input
flabel metal2 s 46358 703520 46470 704960 0 FreeSans 448 90 0 0 la_oenb[12]
port 448 nsew signal input
flabel metal2 s 235050 -960 235162 480 0 FreeSans 448 90 0 0 la_oenb[13]
port 449 nsew signal input
flabel metal2 s 282062 703520 282174 704960 0 FreeSans 448 90 0 0 la_oenb[14]
port 450 nsew signal input
flabel metal3 s 583520 641868 584960 642108 0 FreeSans 960 0 0 0 la_oenb[15]
port 451 nsew signal input
flabel metal3 s 583520 305268 584960 305508 0 FreeSans 960 0 0 0 la_oenb[16]
port 452 nsew signal input
flabel metal3 s -960 316148 480 316388 0 FreeSans 960 0 0 0 la_oenb[17]
port 453 nsew signal input
flabel metal2 s 542882 -960 542994 480 0 FreeSans 448 90 0 0 la_oenb[18]
port 454 nsew signal input
flabel metal3 s 583520 248828 584960 249068 0 FreeSans 960 0 0 0 la_oenb[19]
port 455 nsew signal input
flabel metal3 s 583520 545988 584960 546228 0 FreeSans 960 0 0 0 la_oenb[1]
port 456 nsew signal input
flabel metal2 s 278198 703520 278310 704960 0 FreeSans 448 90 0 0 la_oenb[20]
port 457 nsew signal input
flabel metal3 s -960 152268 480 152508 0 FreeSans 960 0 0 0 la_oenb[21]
port 458 nsew signal input
flabel metal2 s 349038 -960 349150 480 0 FreeSans 448 90 0 0 la_oenb[22]
port 459 nsew signal input
flabel metal2 s 185462 -960 185574 480 0 FreeSans 448 90 0 0 la_oenb[23]
port 460 nsew signal input
flabel metal3 s 583520 193068 584960 193308 0 FreeSans 960 0 0 0 la_oenb[24]
port 461 nsew signal input
flabel metal2 s 41206 -960 41318 480 0 FreeSans 448 90 0 0 la_oenb[25]
port 462 nsew signal input
flabel metal2 s 193190 -960 193302 480 0 FreeSans 448 90 0 0 la_oenb[26]
port 463 nsew signal input
flabel metal3 s 583520 176748 584960 176988 0 FreeSans 960 0 0 0 la_oenb[27]
port 464 nsew signal input
flabel metal2 s 578302 703520 578414 704960 0 FreeSans 448 90 0 0 la_oenb[28]
port 465 nsew signal input
flabel metal3 s 583520 361028 584960 361268 0 FreeSans 960 0 0 0 la_oenb[29]
port 466 nsew signal input
flabel metal2 s 68254 -960 68366 480 0 FreeSans 448 90 0 0 la_oenb[2]
port 467 nsew signal input
flabel metal3 s -960 216188 480 216428 0 FreeSans 960 0 0 0 la_oenb[30]
port 468 nsew signal input
flabel metal3 s -960 15588 480 15828 0 FreeSans 960 0 0 0 la_oenb[31]
port 469 nsew signal input
flabel metal3 s -960 244068 480 244308 0 FreeSans 960 0 0 0 la_oenb[32]
port 470 nsew signal input
flabel metal2 s 421166 -960 421278 480 0 FreeSans 448 90 0 0 la_oenb[33]
port 471 nsew signal input
flabel metal3 s 583520 445348 584960 445588 0 FreeSans 960 0 0 0 la_oenb[34]
port 472 nsew signal input
flabel metal2 s 536442 703520 536554 704960 0 FreeSans 448 90 0 0 la_oenb[35]
port 473 nsew signal input
flabel metal3 s -960 596988 480 597228 0 FreeSans 960 0 0 0 la_oenb[36]
port 474 nsew signal input
flabel metal2 s 300738 703520 300850 704960 0 FreeSans 448 90 0 0 la_oenb[37]
port 475 nsew signal input
flabel metal2 s 544170 703520 544282 704960 0 FreeSans 448 90 0 0 la_oenb[38]
port 476 nsew signal input
flabel metal2 s 72762 703520 72874 704960 0 FreeSans 448 90 0 0 la_oenb[39]
port 477 nsew signal input
flabel metal3 s -960 300508 480 300748 0 FreeSans 960 0 0 0 la_oenb[3]
port 478 nsew signal input
flabel metal3 s 583520 116908 584960 117148 0 FreeSans 960 0 0 0 la_oenb[40]
port 479 nsew signal input
flabel metal3 s 583520 293028 584960 293268 0 FreeSans 960 0 0 0 la_oenb[41]
port 480 nsew signal input
flabel metal3 s 583520 465748 584960 465988 0 FreeSans 960 0 0 0 la_oenb[42]
port 481 nsew signal input
flabel metal2 s 209934 703520 210046 704960 0 FreeSans 448 90 0 0 la_oenb[43]
port 482 nsew signal input
flabel metal2 s 501022 -960 501134 480 0 FreeSans 448 90 0 0 la_oenb[44]
port 483 nsew signal input
flabel metal3 s -960 653428 480 653668 0 FreeSans 960 0 0 0 la_oenb[45]
port 484 nsew signal input
flabel metal3 s -960 99908 480 100148 0 FreeSans 960 0 0 0 la_oenb[46]
port 485 nsew signal input
flabel metal2 s 486854 703520 486966 704960 0 FreeSans 448 90 0 0 la_oenb[47]
port 486 nsew signal input
flabel metal3 s 583520 681988 584960 682228 0 FreeSans 960 0 0 0 la_oenb[48]
port 487 nsew signal input
flabel metal3 s 583520 20348 584960 20588 0 FreeSans 960 0 0 0 la_oenb[49]
port 488 nsew signal input
flabel metal3 s -960 11508 480 11748 0 FreeSans 960 0 0 0 la_oenb[4]
port 489 nsew signal input
flabel metal2 s 577014 -960 577126 480 0 FreeSans 448 90 0 0 la_oenb[50]
port 490 nsew signal input
flabel metal3 s 583520 112828 584960 113068 0 FreeSans 960 0 0 0 la_oenb[51]
port 491 nsew signal input
flabel metal2 s 117198 -960 117310 480 0 FreeSans 448 90 0 0 la_oenb[52]
port 492 nsew signal input
flabel metal2 s 178378 -960 178490 480 0 FreeSans 448 90 0 0 la_oenb[53]
port 493 nsew signal input
flabel metal3 s 583520 36668 584960 36908 0 FreeSans 960 0 0 0 la_oenb[54]
port 494 nsew signal input
flabel metal3 s 583520 273308 584960 273548 0 FreeSans 960 0 0 0 la_oenb[55]
port 495 nsew signal input
flabel metal3 s 583520 622148 584960 622388 0 FreeSans 960 0 0 0 la_oenb[56]
port 496 nsew signal input
flabel metal2 s 228610 703520 228722 704960 0 FreeSans 448 90 0 0 la_oenb[57]
port 497 nsew signal input
flabel metal2 s 202206 703520 202318 704960 0 FreeSans 448 90 0 0 la_oenb[58]
port 498 nsew signal input
flabel metal2 s 99810 703520 99922 704960 0 FreeSans 448 90 0 0 la_oenb[59]
port 499 nsew signal input
flabel metal2 s 220238 -960 220350 480 0 FreeSans 448 90 0 0 la_oenb[5]
port 500 nsew signal input
flabel metal3 s 583520 690148 584960 690388 0 FreeSans 960 0 0 0 la_oenb[60]
port 501 nsew signal input
flabel metal3 s -960 155668 480 155908 0 FreeSans 960 0 0 0 la_oenb[61]
port 502 nsew signal input
flabel metal2 s 65678 703520 65790 704960 0 FreeSans 448 90 0 0 la_oenb[62]
port 503 nsew signal input
flabel metal3 s -960 51628 480 51868 0 FreeSans 960 0 0 0 la_oenb[63]
port 504 nsew signal input
flabel metal3 s 583520 609908 584960 610148 0 FreeSans 960 0 0 0 la_oenb[64]
port 505 nsew signal input
flabel metal2 s 350326 703520 350438 704960 0 FreeSans 448 90 0 0 la_oenb[65]
port 506 nsew signal input
flabel metal2 s 312330 703520 312442 704960 0 FreeSans 448 90 0 0 la_oenb[66]
port 507 nsew signal input
flabel metal2 s 426318 703520 426430 704960 0 FreeSans 448 90 0 0 la_oenb[67]
port 508 nsew signal input
flabel metal2 s 460450 703520 460562 704960 0 FreeSans 448 90 0 0 la_oenb[68]
port 509 nsew signal input
flabel metal2 s 464314 703520 464426 704960 0 FreeSans 448 90 0 0 la_oenb[69]
port 510 nsew signal input
flabel metal3 s -960 252228 480 252468 0 FreeSans 960 0 0 0 la_oenb[6]
port 511 nsew signal input
flabel metal2 s 247930 703520 248042 704960 0 FreeSans 448 90 0 0 la_oenb[70]
port 512 nsew signal input
flabel metal3 s -960 224348 480 224588 0 FreeSans 960 0 0 0 la_oenb[71]
port 513 nsew signal input
flabel metal2 s 7074 -960 7186 480 0 FreeSans 448 90 0 0 la_oenb[72]
port 514 nsew signal input
flabel metal2 s 573150 -960 573262 480 0 FreeSans 448 90 0 0 la_oenb[73]
port 515 nsew signal input
flabel metal2 s 387034 -960 387146 480 0 FreeSans 448 90 0 0 la_oenb[74]
port 516 nsew signal input
flabel metal3 s 583520 200548 584960 200788 0 FreeSans 960 0 0 0 la_oenb[75]
port 517 nsew signal input
flabel metal2 s 316194 703520 316306 704960 0 FreeSans 448 90 0 0 la_oenb[76]
port 518 nsew signal input
flabel metal3 s 583520 265148 584960 265388 0 FreeSans 960 0 0 0 la_oenb[77]
port 519 nsew signal input
flabel metal3 s -960 581348 480 581588 0 FreeSans 960 0 0 0 la_oenb[78]
port 520 nsew signal input
flabel metal2 s 30258 -960 30370 480 0 FreeSans 448 90 0 0 la_oenb[79]
port 521 nsew signal input
flabel metal3 s -960 260388 480 260628 0 FreeSans 960 0 0 0 la_oenb[7]
port 522 nsew signal input
flabel metal3 s -960 171988 480 172228 0 FreeSans 960 0 0 0 la_oenb[80]
port 523 nsew signal input
flabel metal2 s 236338 703520 236450 704960 0 FreeSans 448 90 0 0 la_oenb[81]
port 524 nsew signal input
flabel metal3 s 583520 4708 584960 4948 0 FreeSans 960 0 0 0 la_oenb[82]
port 525 nsew signal input
flabel metal2 s 280774 -960 280886 480 0 FreeSans 448 90 0 0 la_oenb[83]
port 526 nsew signal input
flabel metal3 s -960 492948 480 493188 0 FreeSans 960 0 0 0 la_oenb[84]
port 527 nsew signal input
flabel metal3 s 583520 533748 584960 533988 0 FreeSans 960 0 0 0 la_oenb[85]
port 528 nsew signal input
flabel metal3 s 583520 669748 584960 669988 0 FreeSans 960 0 0 0 la_oenb[86]
port 529 nsew signal input
flabel metal2 s 565422 -960 565534 480 0 FreeSans 448 90 0 0 la_oenb[87]
port 530 nsew signal input
flabel metal3 s -960 584748 480 584988 0 FreeSans 960 0 0 0 la_oenb[88]
port 531 nsew signal input
flabel metal3 s -960 131868 480 132108 0 FreeSans 960 0 0 0 la_oenb[89]
port 532 nsew signal input
flabel metal3 s 583520 637788 584960 638028 0 FreeSans 960 0 0 0 la_oenb[8]
port 533 nsew signal input
flabel metal2 s 152618 703520 152730 704960 0 FreeSans 448 90 0 0 la_oenb[90]
port 534 nsew signal input
flabel metal3 s -960 39388 480 39628 0 FreeSans 960 0 0 0 la_oenb[91]
port 535 nsew signal input
flabel metal2 s 550610 -960 550722 480 0 FreeSans 448 90 0 0 la_oenb[92]
port 536 nsew signal input
flabel metal2 s 308466 703520 308578 704960 0 FreeSans 448 90 0 0 la_oenb[93]
port 537 nsew signal input
flabel metal3 s 583520 220948 584960 221188 0 FreeSans 960 0 0 0 la_oenb[94]
port 538 nsew signal input
flabel metal2 s 103674 703520 103786 704960 0 FreeSans 448 90 0 0 la_oenb[95]
port 539 nsew signal input
flabel metal3 s -960 372588 480 372828 0 FreeSans 960 0 0 0 la_oenb[96]
port 540 nsew signal input
flabel metal3 s -960 556868 480 557108 0 FreeSans 960 0 0 0 la_oenb[97]
port 541 nsew signal input
flabel metal2 s 90794 -960 90906 480 0 FreeSans 448 90 0 0 la_oenb[98]
port 542 nsew signal input
flabel metal3 s 583520 517428 584960 517668 0 FreeSans 960 0 0 0 la_oenb[99]
port 543 nsew signal input
flabel metal2 s 402490 -960 402602 480 0 FreeSans 448 90 0 0 la_oenb[9]
port 544 nsew signal input
flabel metal3 s -960 220268 480 220508 0 FreeSans 960 0 0 0 pxl_done
port 545 nsew signal tristate
flabel metal2 s 182242 -960 182354 480 0 FreeSans 448 90 0 0 pxl_start_in_path
port 546 nsew signal input
flabel metal3 s -960 292348 480 292588 0 FreeSans 960 0 0 0 pxl_start_out_path
port 547 nsew signal input
flabel metal3 s -960 613308 480 613548 0 FreeSans 960 0 0 0 serial_data_rlbp_out
port 548 nsew signal tristate
flabel metal2 s 320058 703520 320170 704960 0 FreeSans 448 90 0 0 user_clock2
port 549 nsew signal input
flabel metal3 s 583520 702388 584960 702628 0 FreeSans 960 0 0 0 user_irq[0]
port 550 nsew signal tristate
flabel metal3 s -960 592908 480 593148 0 FreeSans 960 0 0 0 user_irq[1]
port 551 nsew signal tristate
flabel metal3 s -960 660908 480 661148 0 FreeSans 960 0 0 0 user_irq[2]
port 552 nsew signal tristate
flabel metal4 s -2006 -934 -1386 704870 0 FreeSans 3840 90 0 0 vccd1
port 553 nsew power bidirectional
flabel metal5 s -2006 -934 585930 -314 0 FreeSans 2560 0 0 0 vccd1
port 553 nsew power bidirectional
flabel metal5 s -2006 704250 585930 704870 0 FreeSans 2560 0 0 0 vccd1
port 553 nsew power bidirectional
flabel metal4 s 585310 -934 585930 704870 0 FreeSans 3840 90 0 0 vccd1
port 553 nsew power bidirectional
flabel metal4 s 1794 -7654 2414 711590 0 FreeSans 3840 90 0 0 vccd1
port 553 nsew power bidirectional
flabel metal4 s 37794 -7654 38414 711590 0 FreeSans 3840 90 0 0 vccd1
port 553 nsew power bidirectional
flabel metal4 s 73794 -7654 74414 711590 0 FreeSans 3840 90 0 0 vccd1
port 553 nsew power bidirectional
flabel metal4 s 109794 -7654 110414 711590 0 FreeSans 3840 90 0 0 vccd1
port 553 nsew power bidirectional
flabel metal4 s 145794 -7654 146414 78000 0 FreeSans 3840 90 0 0 vccd1
port 553 nsew power bidirectional
flabel metal4 s 145794 142000 146414 198000 0 FreeSans 3840 90 0 0 vccd1
port 553 nsew power bidirectional
flabel metal4 s 145794 262000 146414 711590 0 FreeSans 3840 90 0 0 vccd1
port 553 nsew power bidirectional
flabel metal4 s 181794 -7654 182414 78000 0 FreeSans 3840 90 0 0 vccd1
port 553 nsew power bidirectional
flabel metal4 s 181794 142000 182414 198000 0 FreeSans 3840 90 0 0 vccd1
port 553 nsew power bidirectional
flabel metal4 s 181794 262000 182414 711590 0 FreeSans 3840 90 0 0 vccd1
port 553 nsew power bidirectional
flabel metal4 s 217794 -7654 218414 711590 0 FreeSans 3840 90 0 0 vccd1
port 553 nsew power bidirectional
flabel metal4 s 253794 -7654 254414 711590 0 FreeSans 3840 90 0 0 vccd1
port 553 nsew power bidirectional
flabel metal4 s 289794 -7654 290414 711590 0 FreeSans 3840 90 0 0 vccd1
port 553 nsew power bidirectional
flabel metal4 s 325794 -7654 326414 711590 0 FreeSans 3840 90 0 0 vccd1
port 553 nsew power bidirectional
flabel metal4 s 361794 -7654 362414 711590 0 FreeSans 3840 90 0 0 vccd1
port 553 nsew power bidirectional
flabel metal4 s 397794 -7654 398414 711590 0 FreeSans 3840 90 0 0 vccd1
port 553 nsew power bidirectional
flabel metal4 s 433794 -7654 434414 711590 0 FreeSans 3840 90 0 0 vccd1
port 553 nsew power bidirectional
flabel metal4 s 469794 -7654 470414 711590 0 FreeSans 3840 90 0 0 vccd1
port 553 nsew power bidirectional
flabel metal4 s 505794 -7654 506414 711590 0 FreeSans 3840 90 0 0 vccd1
port 553 nsew power bidirectional
flabel metal4 s 541794 -7654 542414 711590 0 FreeSans 3840 90 0 0 vccd1
port 553 nsew power bidirectional
flabel metal4 s 577794 -7654 578414 711590 0 FreeSans 3840 90 0 0 vccd1
port 553 nsew power bidirectional
flabel metal5 s -8726 2866 592650 3486 0 FreeSans 2560 0 0 0 vccd1
port 553 nsew power bidirectional
flabel metal5 s -8726 38866 592650 39486 0 FreeSans 2560 0 0 0 vccd1
port 553 nsew power bidirectional
flabel metal5 s -8726 74866 592650 75486 0 FreeSans 2560 0 0 0 vccd1
port 553 nsew power bidirectional
flabel metal5 s -8726 110866 592650 111486 0 FreeSans 2560 0 0 0 vccd1
port 553 nsew power bidirectional
flabel metal5 s -8726 146866 592650 147486 0 FreeSans 2560 0 0 0 vccd1
port 553 nsew power bidirectional
flabel metal5 s -8726 182866 592650 183486 0 FreeSans 2560 0 0 0 vccd1
port 553 nsew power bidirectional
flabel metal5 s -8726 218866 592650 219486 0 FreeSans 2560 0 0 0 vccd1
port 553 nsew power bidirectional
flabel metal5 s -8726 254866 592650 255486 0 FreeSans 2560 0 0 0 vccd1
port 553 nsew power bidirectional
flabel metal5 s -8726 290866 592650 291486 0 FreeSans 2560 0 0 0 vccd1
port 553 nsew power bidirectional
flabel metal5 s -8726 326866 592650 327486 0 FreeSans 2560 0 0 0 vccd1
port 553 nsew power bidirectional
flabel metal5 s -8726 362866 592650 363486 0 FreeSans 2560 0 0 0 vccd1
port 553 nsew power bidirectional
flabel metal5 s -8726 398866 592650 399486 0 FreeSans 2560 0 0 0 vccd1
port 553 nsew power bidirectional
flabel metal5 s -8726 434866 592650 435486 0 FreeSans 2560 0 0 0 vccd1
port 553 nsew power bidirectional
flabel metal5 s -8726 470866 592650 471486 0 FreeSans 2560 0 0 0 vccd1
port 553 nsew power bidirectional
flabel metal5 s -8726 506866 592650 507486 0 FreeSans 2560 0 0 0 vccd1
port 553 nsew power bidirectional
flabel metal5 s -8726 542866 592650 543486 0 FreeSans 2560 0 0 0 vccd1
port 553 nsew power bidirectional
flabel metal5 s -8726 578866 592650 579486 0 FreeSans 2560 0 0 0 vccd1
port 553 nsew power bidirectional
flabel metal5 s -8726 614866 592650 615486 0 FreeSans 2560 0 0 0 vccd1
port 553 nsew power bidirectional
flabel metal5 s -8726 650866 592650 651486 0 FreeSans 2560 0 0 0 vccd1
port 553 nsew power bidirectional
flabel metal5 s -8726 686866 592650 687486 0 FreeSans 2560 0 0 0 vccd1
port 553 nsew power bidirectional
flabel metal4 s -3926 -2854 -3306 706790 0 FreeSans 3840 90 0 0 vccd2
port 554 nsew power bidirectional
flabel metal5 s -3926 -2854 587850 -2234 0 FreeSans 2560 0 0 0 vccd2
port 554 nsew power bidirectional
flabel metal5 s -3926 706170 587850 706790 0 FreeSans 2560 0 0 0 vccd2
port 554 nsew power bidirectional
flabel metal4 s 587230 -2854 587850 706790 0 FreeSans 3840 90 0 0 vccd2
port 554 nsew power bidirectional
flabel metal4 s 10794 -7654 11414 711590 0 FreeSans 3840 90 0 0 vccd2
port 554 nsew power bidirectional
flabel metal4 s 46794 -7654 47414 711590 0 FreeSans 3840 90 0 0 vccd2
port 554 nsew power bidirectional
flabel metal4 s 82794 -7654 83414 711590 0 FreeSans 3840 90 0 0 vccd2
port 554 nsew power bidirectional
flabel metal4 s 118794 -7654 119414 78000 0 FreeSans 3840 90 0 0 vccd2
port 554 nsew power bidirectional
flabel metal4 s 118794 142000 119414 198000 0 FreeSans 3840 90 0 0 vccd2
port 554 nsew power bidirectional
flabel metal4 s 118794 262000 119414 711590 0 FreeSans 3840 90 0 0 vccd2
port 554 nsew power bidirectional
flabel metal4 s 154794 -7654 155414 78000 0 FreeSans 3840 90 0 0 vccd2
port 554 nsew power bidirectional
flabel metal4 s 154794 142000 155414 198000 0 FreeSans 3840 90 0 0 vccd2
port 554 nsew power bidirectional
flabel metal4 s 154794 262000 155414 711590 0 FreeSans 3840 90 0 0 vccd2
port 554 nsew power bidirectional
flabel metal4 s 190794 -7654 191414 78000 0 FreeSans 3840 90 0 0 vccd2
port 554 nsew power bidirectional
flabel metal4 s 190794 142000 191414 198000 0 FreeSans 3840 90 0 0 vccd2
port 554 nsew power bidirectional
flabel metal4 s 190794 262000 191414 711590 0 FreeSans 3840 90 0 0 vccd2
port 554 nsew power bidirectional
flabel metal4 s 226794 -7654 227414 711590 0 FreeSans 3840 90 0 0 vccd2
port 554 nsew power bidirectional
flabel metal4 s 262794 -7654 263414 711590 0 FreeSans 3840 90 0 0 vccd2
port 554 nsew power bidirectional
flabel metal4 s 298794 -7654 299414 711590 0 FreeSans 3840 90 0 0 vccd2
port 554 nsew power bidirectional
flabel metal4 s 334794 -7654 335414 711590 0 FreeSans 3840 90 0 0 vccd2
port 554 nsew power bidirectional
flabel metal4 s 370794 -7654 371414 711590 0 FreeSans 3840 90 0 0 vccd2
port 554 nsew power bidirectional
flabel metal4 s 406794 -7654 407414 711590 0 FreeSans 3840 90 0 0 vccd2
port 554 nsew power bidirectional
flabel metal4 s 442794 -7654 443414 711590 0 FreeSans 3840 90 0 0 vccd2
port 554 nsew power bidirectional
flabel metal4 s 478794 -7654 479414 711590 0 FreeSans 3840 90 0 0 vccd2
port 554 nsew power bidirectional
flabel metal4 s 514794 -7654 515414 711590 0 FreeSans 3840 90 0 0 vccd2
port 554 nsew power bidirectional
flabel metal4 s 550794 -7654 551414 711590 0 FreeSans 3840 90 0 0 vccd2
port 554 nsew power bidirectional
flabel metal5 s -8726 11866 592650 12486 0 FreeSans 2560 0 0 0 vccd2
port 554 nsew power bidirectional
flabel metal5 s -8726 47866 592650 48486 0 FreeSans 2560 0 0 0 vccd2
port 554 nsew power bidirectional
flabel metal5 s -8726 83866 592650 84486 0 FreeSans 2560 0 0 0 vccd2
port 554 nsew power bidirectional
flabel metal5 s -8726 119866 592650 120486 0 FreeSans 2560 0 0 0 vccd2
port 554 nsew power bidirectional
flabel metal5 s -8726 155866 592650 156486 0 FreeSans 2560 0 0 0 vccd2
port 554 nsew power bidirectional
flabel metal5 s -8726 191866 592650 192486 0 FreeSans 2560 0 0 0 vccd2
port 554 nsew power bidirectional
flabel metal5 s -8726 227866 592650 228486 0 FreeSans 2560 0 0 0 vccd2
port 554 nsew power bidirectional
flabel metal5 s -8726 263866 592650 264486 0 FreeSans 2560 0 0 0 vccd2
port 554 nsew power bidirectional
flabel metal5 s -8726 299866 592650 300486 0 FreeSans 2560 0 0 0 vccd2
port 554 nsew power bidirectional
flabel metal5 s -8726 335866 592650 336486 0 FreeSans 2560 0 0 0 vccd2
port 554 nsew power bidirectional
flabel metal5 s -8726 371866 592650 372486 0 FreeSans 2560 0 0 0 vccd2
port 554 nsew power bidirectional
flabel metal5 s -8726 407866 592650 408486 0 FreeSans 2560 0 0 0 vccd2
port 554 nsew power bidirectional
flabel metal5 s -8726 443866 592650 444486 0 FreeSans 2560 0 0 0 vccd2
port 554 nsew power bidirectional
flabel metal5 s -8726 479866 592650 480486 0 FreeSans 2560 0 0 0 vccd2
port 554 nsew power bidirectional
flabel metal5 s -8726 515866 592650 516486 0 FreeSans 2560 0 0 0 vccd2
port 554 nsew power bidirectional
flabel metal5 s -8726 551866 592650 552486 0 FreeSans 2560 0 0 0 vccd2
port 554 nsew power bidirectional
flabel metal5 s -8726 587866 592650 588486 0 FreeSans 2560 0 0 0 vccd2
port 554 nsew power bidirectional
flabel metal5 s -8726 623866 592650 624486 0 FreeSans 2560 0 0 0 vccd2
port 554 nsew power bidirectional
flabel metal5 s -8726 659866 592650 660486 0 FreeSans 2560 0 0 0 vccd2
port 554 nsew power bidirectional
flabel metal5 s -8726 695866 592650 696486 0 FreeSans 2560 0 0 0 vccd2
port 554 nsew power bidirectional
flabel metal4 s -5846 -4774 -5226 708710 0 FreeSans 3840 90 0 0 vdda1
port 555 nsew power bidirectional
flabel metal5 s -5846 -4774 589770 -4154 0 FreeSans 2560 0 0 0 vdda1
port 555 nsew power bidirectional
flabel metal5 s -5846 708090 589770 708710 0 FreeSans 2560 0 0 0 vdda1
port 555 nsew power bidirectional
flabel metal4 s 589150 -4774 589770 708710 0 FreeSans 3840 90 0 0 vdda1
port 555 nsew power bidirectional
flabel metal4 s 19794 -7654 20414 711590 0 FreeSans 3840 90 0 0 vdda1
port 555 nsew power bidirectional
flabel metal4 s 55794 -7654 56414 711590 0 FreeSans 3840 90 0 0 vdda1
port 555 nsew power bidirectional
flabel metal4 s 91794 -7654 92414 711590 0 FreeSans 3840 90 0 0 vdda1
port 555 nsew power bidirectional
flabel metal4 s 127794 -7654 128414 78000 0 FreeSans 3840 90 0 0 vdda1
port 555 nsew power bidirectional
flabel metal4 s 127794 262000 128414 711590 0 FreeSans 3840 90 0 0 vdda1
port 555 nsew power bidirectional
flabel metal4 s 163794 -7654 164414 78000 0 FreeSans 3840 90 0 0 vdda1
port 555 nsew power bidirectional
flabel metal4 s 163794 262000 164414 711590 0 FreeSans 3840 90 0 0 vdda1
port 555 nsew power bidirectional
flabel metal4 s 199794 -7654 200414 711590 0 FreeSans 3840 90 0 0 vdda1
port 555 nsew power bidirectional
flabel metal4 s 235794 -7654 236414 711590 0 FreeSans 3840 90 0 0 vdda1
port 555 nsew power bidirectional
flabel metal4 s 271794 -7654 272414 711590 0 FreeSans 3840 90 0 0 vdda1
port 555 nsew power bidirectional
flabel metal4 s 307794 -7654 308414 711590 0 FreeSans 3840 90 0 0 vdda1
port 555 nsew power bidirectional
flabel metal4 s 343794 -7654 344414 711590 0 FreeSans 3840 90 0 0 vdda1
port 555 nsew power bidirectional
flabel metal4 s 379794 -7654 380414 711590 0 FreeSans 3840 90 0 0 vdda1
port 555 nsew power bidirectional
flabel metal4 s 415794 -7654 416414 711590 0 FreeSans 3840 90 0 0 vdda1
port 555 nsew power bidirectional
flabel metal4 s 451794 -7654 452414 711590 0 FreeSans 3840 90 0 0 vdda1
port 555 nsew power bidirectional
flabel metal4 s 487794 -7654 488414 711590 0 FreeSans 3840 90 0 0 vdda1
port 555 nsew power bidirectional
flabel metal4 s 523794 -7654 524414 711590 0 FreeSans 3840 90 0 0 vdda1
port 555 nsew power bidirectional
flabel metal4 s 559794 -7654 560414 711590 0 FreeSans 3840 90 0 0 vdda1
port 555 nsew power bidirectional
flabel metal5 s -8726 20866 592650 21486 0 FreeSans 2560 0 0 0 vdda1
port 555 nsew power bidirectional
flabel metal5 s -8726 56866 592650 57486 0 FreeSans 2560 0 0 0 vdda1
port 555 nsew power bidirectional
flabel metal5 s -8726 92866 592650 93486 0 FreeSans 2560 0 0 0 vdda1
port 555 nsew power bidirectional
flabel metal5 s -8726 128866 592650 129486 0 FreeSans 2560 0 0 0 vdda1
port 555 nsew power bidirectional
flabel metal5 s -8726 164866 592650 165486 0 FreeSans 2560 0 0 0 vdda1
port 555 nsew power bidirectional
flabel metal5 s -8726 200866 592650 201486 0 FreeSans 2560 0 0 0 vdda1
port 555 nsew power bidirectional
flabel metal5 s -8726 236866 592650 237486 0 FreeSans 2560 0 0 0 vdda1
port 555 nsew power bidirectional
flabel metal5 s -8726 272866 592650 273486 0 FreeSans 2560 0 0 0 vdda1
port 555 nsew power bidirectional
flabel metal5 s -8726 308866 592650 309486 0 FreeSans 2560 0 0 0 vdda1
port 555 nsew power bidirectional
flabel metal5 s -8726 344866 592650 345486 0 FreeSans 2560 0 0 0 vdda1
port 555 nsew power bidirectional
flabel metal5 s -8726 380866 592650 381486 0 FreeSans 2560 0 0 0 vdda1
port 555 nsew power bidirectional
flabel metal5 s -8726 416866 592650 417486 0 FreeSans 2560 0 0 0 vdda1
port 555 nsew power bidirectional
flabel metal5 s -8726 452866 592650 453486 0 FreeSans 2560 0 0 0 vdda1
port 555 nsew power bidirectional
flabel metal5 s -8726 488866 592650 489486 0 FreeSans 2560 0 0 0 vdda1
port 555 nsew power bidirectional
flabel metal5 s -8726 524866 592650 525486 0 FreeSans 2560 0 0 0 vdda1
port 555 nsew power bidirectional
flabel metal5 s -8726 560866 592650 561486 0 FreeSans 2560 0 0 0 vdda1
port 555 nsew power bidirectional
flabel metal5 s -8726 596866 592650 597486 0 FreeSans 2560 0 0 0 vdda1
port 555 nsew power bidirectional
flabel metal5 s -8726 632866 592650 633486 0 FreeSans 2560 0 0 0 vdda1
port 555 nsew power bidirectional
flabel metal5 s -8726 668866 592650 669486 0 FreeSans 2560 0 0 0 vdda1
port 555 nsew power bidirectional
flabel metal4 s -7766 -6694 -7146 710630 0 FreeSans 3840 90 0 0 vdda2
port 556 nsew power bidirectional
flabel metal5 s -7766 -6694 591690 -6074 0 FreeSans 2560 0 0 0 vdda2
port 556 nsew power bidirectional
flabel metal5 s -7766 710010 591690 710630 0 FreeSans 2560 0 0 0 vdda2
port 556 nsew power bidirectional
flabel metal4 s 591070 -6694 591690 710630 0 FreeSans 3840 90 0 0 vdda2
port 556 nsew power bidirectional
flabel metal4 s 28794 -7654 29414 711590 0 FreeSans 3840 90 0 0 vdda2
port 556 nsew power bidirectional
flabel metal4 s 64794 -7654 65414 711590 0 FreeSans 3840 90 0 0 vdda2
port 556 nsew power bidirectional
flabel metal4 s 100794 -7654 101414 711590 0 FreeSans 3840 90 0 0 vdda2
port 556 nsew power bidirectional
flabel metal4 s 136794 -7654 137414 78000 0 FreeSans 3840 90 0 0 vdda2
port 556 nsew power bidirectional
flabel metal4 s 136794 262000 137414 711590 0 FreeSans 3840 90 0 0 vdda2
port 556 nsew power bidirectional
flabel metal4 s 172794 -7654 173414 78000 0 FreeSans 3840 90 0 0 vdda2
port 556 nsew power bidirectional
flabel metal4 s 172794 262000 173414 711590 0 FreeSans 3840 90 0 0 vdda2
port 556 nsew power bidirectional
flabel metal4 s 208794 -7654 209414 711590 0 FreeSans 3840 90 0 0 vdda2
port 556 nsew power bidirectional
flabel metal4 s 244794 -7654 245414 711590 0 FreeSans 3840 90 0 0 vdda2
port 556 nsew power bidirectional
flabel metal4 s 280794 -7654 281414 711590 0 FreeSans 3840 90 0 0 vdda2
port 556 nsew power bidirectional
flabel metal4 s 316794 -7654 317414 711590 0 FreeSans 3840 90 0 0 vdda2
port 556 nsew power bidirectional
flabel metal4 s 352794 -7654 353414 711590 0 FreeSans 3840 90 0 0 vdda2
port 556 nsew power bidirectional
flabel metal4 s 388794 -7654 389414 711590 0 FreeSans 3840 90 0 0 vdda2
port 556 nsew power bidirectional
flabel metal4 s 424794 -7654 425414 711590 0 FreeSans 3840 90 0 0 vdda2
port 556 nsew power bidirectional
flabel metal4 s 460794 -7654 461414 711590 0 FreeSans 3840 90 0 0 vdda2
port 556 nsew power bidirectional
flabel metal4 s 496794 -7654 497414 711590 0 FreeSans 3840 90 0 0 vdda2
port 556 nsew power bidirectional
flabel metal4 s 532794 -7654 533414 711590 0 FreeSans 3840 90 0 0 vdda2
port 556 nsew power bidirectional
flabel metal4 s 568794 -7654 569414 711590 0 FreeSans 3840 90 0 0 vdda2
port 556 nsew power bidirectional
flabel metal5 s -8726 29866 592650 30486 0 FreeSans 2560 0 0 0 vdda2
port 556 nsew power bidirectional
flabel metal5 s -8726 65866 592650 66486 0 FreeSans 2560 0 0 0 vdda2
port 556 nsew power bidirectional
flabel metal5 s -8726 101866 592650 102486 0 FreeSans 2560 0 0 0 vdda2
port 556 nsew power bidirectional
flabel metal5 s -8726 137866 592650 138486 0 FreeSans 2560 0 0 0 vdda2
port 556 nsew power bidirectional
flabel metal5 s -8726 173866 592650 174486 0 FreeSans 2560 0 0 0 vdda2
port 556 nsew power bidirectional
flabel metal5 s -8726 209866 592650 210486 0 FreeSans 2560 0 0 0 vdda2
port 556 nsew power bidirectional
flabel metal5 s -8726 245866 592650 246486 0 FreeSans 2560 0 0 0 vdda2
port 556 nsew power bidirectional
flabel metal5 s -8726 281866 592650 282486 0 FreeSans 2560 0 0 0 vdda2
port 556 nsew power bidirectional
flabel metal5 s -8726 317866 592650 318486 0 FreeSans 2560 0 0 0 vdda2
port 556 nsew power bidirectional
flabel metal5 s -8726 353866 592650 354486 0 FreeSans 2560 0 0 0 vdda2
port 556 nsew power bidirectional
flabel metal5 s -8726 389866 592650 390486 0 FreeSans 2560 0 0 0 vdda2
port 556 nsew power bidirectional
flabel metal5 s -8726 425866 592650 426486 0 FreeSans 2560 0 0 0 vdda2
port 556 nsew power bidirectional
flabel metal5 s -8726 461866 592650 462486 0 FreeSans 2560 0 0 0 vdda2
port 556 nsew power bidirectional
flabel metal5 s -8726 497866 592650 498486 0 FreeSans 2560 0 0 0 vdda2
port 556 nsew power bidirectional
flabel metal5 s -8726 533866 592650 534486 0 FreeSans 2560 0 0 0 vdda2
port 556 nsew power bidirectional
flabel metal5 s -8726 569866 592650 570486 0 FreeSans 2560 0 0 0 vdda2
port 556 nsew power bidirectional
flabel metal5 s -8726 605866 592650 606486 0 FreeSans 2560 0 0 0 vdda2
port 556 nsew power bidirectional
flabel metal5 s -8726 641866 592650 642486 0 FreeSans 2560 0 0 0 vdda2
port 556 nsew power bidirectional
flabel metal5 s -8726 677866 592650 678486 0 FreeSans 2560 0 0 0 vdda2
port 556 nsew power bidirectional
flabel metal4 s -6806 -5734 -6186 709670 0 FreeSans 3840 90 0 0 vssa1
port 557 nsew ground bidirectional
flabel metal5 s -6806 -5734 590730 -5114 0 FreeSans 2560 0 0 0 vssa1
port 557 nsew ground bidirectional
flabel metal5 s -6806 709050 590730 709670 0 FreeSans 2560 0 0 0 vssa1
port 557 nsew ground bidirectional
flabel metal4 s 590110 -5734 590730 709670 0 FreeSans 3840 90 0 0 vssa1
port 557 nsew ground bidirectional
flabel metal4 s 24294 -7654 24914 711590 0 FreeSans 3840 90 0 0 vssa1
port 557 nsew ground bidirectional
flabel metal4 s 60294 -7654 60914 711590 0 FreeSans 3840 90 0 0 vssa1
port 557 nsew ground bidirectional
flabel metal4 s 96294 -7654 96914 711590 0 FreeSans 3840 90 0 0 vssa1
port 557 nsew ground bidirectional
flabel metal4 s 132294 -7654 132914 78000 0 FreeSans 3840 90 0 0 vssa1
port 557 nsew ground bidirectional
flabel metal4 s 132294 262000 132914 711590 0 FreeSans 3840 90 0 0 vssa1
port 557 nsew ground bidirectional
flabel metal4 s 168294 -7654 168914 78000 0 FreeSans 3840 90 0 0 vssa1
port 557 nsew ground bidirectional
flabel metal4 s 168294 262000 168914 711590 0 FreeSans 3840 90 0 0 vssa1
port 557 nsew ground bidirectional
flabel metal4 s 204294 -7654 204914 711590 0 FreeSans 3840 90 0 0 vssa1
port 557 nsew ground bidirectional
flabel metal4 s 240294 -7654 240914 711590 0 FreeSans 3840 90 0 0 vssa1
port 557 nsew ground bidirectional
flabel metal4 s 276294 -7654 276914 711590 0 FreeSans 3840 90 0 0 vssa1
port 557 nsew ground bidirectional
flabel metal4 s 312294 -7654 312914 711590 0 FreeSans 3840 90 0 0 vssa1
port 557 nsew ground bidirectional
flabel metal4 s 348294 -7654 348914 711590 0 FreeSans 3840 90 0 0 vssa1
port 557 nsew ground bidirectional
flabel metal4 s 384294 -7654 384914 711590 0 FreeSans 3840 90 0 0 vssa1
port 557 nsew ground bidirectional
flabel metal4 s 420294 -7654 420914 711590 0 FreeSans 3840 90 0 0 vssa1
port 557 nsew ground bidirectional
flabel metal4 s 456294 -7654 456914 711590 0 FreeSans 3840 90 0 0 vssa1
port 557 nsew ground bidirectional
flabel metal4 s 492294 -7654 492914 711590 0 FreeSans 3840 90 0 0 vssa1
port 557 nsew ground bidirectional
flabel metal4 s 528294 -7654 528914 711590 0 FreeSans 3840 90 0 0 vssa1
port 557 nsew ground bidirectional
flabel metal4 s 564294 -7654 564914 711590 0 FreeSans 3840 90 0 0 vssa1
port 557 nsew ground bidirectional
flabel metal5 s -8726 25366 592650 25986 0 FreeSans 2560 0 0 0 vssa1
port 557 nsew ground bidirectional
flabel metal5 s -8726 61366 592650 61986 0 FreeSans 2560 0 0 0 vssa1
port 557 nsew ground bidirectional
flabel metal5 s -8726 97366 592650 97986 0 FreeSans 2560 0 0 0 vssa1
port 557 nsew ground bidirectional
flabel metal5 s -8726 133366 592650 133986 0 FreeSans 2560 0 0 0 vssa1
port 557 nsew ground bidirectional
flabel metal5 s -8726 169366 592650 169986 0 FreeSans 2560 0 0 0 vssa1
port 557 nsew ground bidirectional
flabel metal5 s -8726 205366 592650 205986 0 FreeSans 2560 0 0 0 vssa1
port 557 nsew ground bidirectional
flabel metal5 s -8726 241366 592650 241986 0 FreeSans 2560 0 0 0 vssa1
port 557 nsew ground bidirectional
flabel metal5 s -8726 277366 592650 277986 0 FreeSans 2560 0 0 0 vssa1
port 557 nsew ground bidirectional
flabel metal5 s -8726 313366 592650 313986 0 FreeSans 2560 0 0 0 vssa1
port 557 nsew ground bidirectional
flabel metal5 s -8726 349366 592650 349986 0 FreeSans 2560 0 0 0 vssa1
port 557 nsew ground bidirectional
flabel metal5 s -8726 385366 592650 385986 0 FreeSans 2560 0 0 0 vssa1
port 557 nsew ground bidirectional
flabel metal5 s -8726 421366 592650 421986 0 FreeSans 2560 0 0 0 vssa1
port 557 nsew ground bidirectional
flabel metal5 s -8726 457366 592650 457986 0 FreeSans 2560 0 0 0 vssa1
port 557 nsew ground bidirectional
flabel metal5 s -8726 493366 592650 493986 0 FreeSans 2560 0 0 0 vssa1
port 557 nsew ground bidirectional
flabel metal5 s -8726 529366 592650 529986 0 FreeSans 2560 0 0 0 vssa1
port 557 nsew ground bidirectional
flabel metal5 s -8726 565366 592650 565986 0 FreeSans 2560 0 0 0 vssa1
port 557 nsew ground bidirectional
flabel metal5 s -8726 601366 592650 601986 0 FreeSans 2560 0 0 0 vssa1
port 557 nsew ground bidirectional
flabel metal5 s -8726 637366 592650 637986 0 FreeSans 2560 0 0 0 vssa1
port 557 nsew ground bidirectional
flabel metal5 s -8726 673366 592650 673986 0 FreeSans 2560 0 0 0 vssa1
port 557 nsew ground bidirectional
flabel metal4 s -8726 -7654 -8106 711590 0 FreeSans 3840 90 0 0 vssa2
port 558 nsew ground bidirectional
flabel metal5 s -8726 -7654 592650 -7034 0 FreeSans 2560 0 0 0 vssa2
port 558 nsew ground bidirectional
flabel metal5 s -8726 710970 592650 711590 0 FreeSans 2560 0 0 0 vssa2
port 558 nsew ground bidirectional
flabel metal4 s 592030 -7654 592650 711590 0 FreeSans 3840 90 0 0 vssa2
port 558 nsew ground bidirectional
flabel metal4 s 33294 -7654 33914 711590 0 FreeSans 3840 90 0 0 vssa2
port 558 nsew ground bidirectional
flabel metal4 s 69294 -7654 69914 711590 0 FreeSans 3840 90 0 0 vssa2
port 558 nsew ground bidirectional
flabel metal4 s 105294 -7654 105914 711590 0 FreeSans 3840 90 0 0 vssa2
port 558 nsew ground bidirectional
flabel metal4 s 141294 -7654 141914 78000 0 FreeSans 3840 90 0 0 vssa2
port 558 nsew ground bidirectional
flabel metal4 s 141294 142000 141914 198000 0 FreeSans 3840 90 0 0 vssa2
port 558 nsew ground bidirectional
flabel metal4 s 141294 262000 141914 711590 0 FreeSans 3840 90 0 0 vssa2
port 558 nsew ground bidirectional
flabel metal4 s 177294 -7654 177914 78000 0 FreeSans 3840 90 0 0 vssa2
port 558 nsew ground bidirectional
flabel metal4 s 177294 142000 177914 198000 0 FreeSans 3840 90 0 0 vssa2
port 558 nsew ground bidirectional
flabel metal4 s 177294 262000 177914 711590 0 FreeSans 3840 90 0 0 vssa2
port 558 nsew ground bidirectional
flabel metal4 s 213294 -7654 213914 711590 0 FreeSans 3840 90 0 0 vssa2
port 558 nsew ground bidirectional
flabel metal4 s 249294 -7654 249914 711590 0 FreeSans 3840 90 0 0 vssa2
port 558 nsew ground bidirectional
flabel metal4 s 285294 -7654 285914 711590 0 FreeSans 3840 90 0 0 vssa2
port 558 nsew ground bidirectional
flabel metal4 s 321294 -7654 321914 711590 0 FreeSans 3840 90 0 0 vssa2
port 558 nsew ground bidirectional
flabel metal4 s 357294 -7654 357914 711590 0 FreeSans 3840 90 0 0 vssa2
port 558 nsew ground bidirectional
flabel metal4 s 393294 -7654 393914 711590 0 FreeSans 3840 90 0 0 vssa2
port 558 nsew ground bidirectional
flabel metal4 s 429294 -7654 429914 711590 0 FreeSans 3840 90 0 0 vssa2
port 558 nsew ground bidirectional
flabel metal4 s 465294 -7654 465914 711590 0 FreeSans 3840 90 0 0 vssa2
port 558 nsew ground bidirectional
flabel metal4 s 501294 -7654 501914 711590 0 FreeSans 3840 90 0 0 vssa2
port 558 nsew ground bidirectional
flabel metal4 s 537294 -7654 537914 711590 0 FreeSans 3840 90 0 0 vssa2
port 558 nsew ground bidirectional
flabel metal4 s 573294 -7654 573914 711590 0 FreeSans 3840 90 0 0 vssa2
port 558 nsew ground bidirectional
flabel metal5 s -8726 34366 592650 34986 0 FreeSans 2560 0 0 0 vssa2
port 558 nsew ground bidirectional
flabel metal5 s -8726 70366 592650 70986 0 FreeSans 2560 0 0 0 vssa2
port 558 nsew ground bidirectional
flabel metal5 s -8726 106366 592650 106986 0 FreeSans 2560 0 0 0 vssa2
port 558 nsew ground bidirectional
flabel metal5 s -8726 142366 592650 142986 0 FreeSans 2560 0 0 0 vssa2
port 558 nsew ground bidirectional
flabel metal5 s -8726 178366 592650 178986 0 FreeSans 2560 0 0 0 vssa2
port 558 nsew ground bidirectional
flabel metal5 s -8726 214366 592650 214986 0 FreeSans 2560 0 0 0 vssa2
port 558 nsew ground bidirectional
flabel metal5 s -8726 250366 592650 250986 0 FreeSans 2560 0 0 0 vssa2
port 558 nsew ground bidirectional
flabel metal5 s -8726 286366 592650 286986 0 FreeSans 2560 0 0 0 vssa2
port 558 nsew ground bidirectional
flabel metal5 s -8726 322366 592650 322986 0 FreeSans 2560 0 0 0 vssa2
port 558 nsew ground bidirectional
flabel metal5 s -8726 358366 592650 358986 0 FreeSans 2560 0 0 0 vssa2
port 558 nsew ground bidirectional
flabel metal5 s -8726 394366 592650 394986 0 FreeSans 2560 0 0 0 vssa2
port 558 nsew ground bidirectional
flabel metal5 s -8726 430366 592650 430986 0 FreeSans 2560 0 0 0 vssa2
port 558 nsew ground bidirectional
flabel metal5 s -8726 466366 592650 466986 0 FreeSans 2560 0 0 0 vssa2
port 558 nsew ground bidirectional
flabel metal5 s -8726 502366 592650 502986 0 FreeSans 2560 0 0 0 vssa2
port 558 nsew ground bidirectional
flabel metal5 s -8726 538366 592650 538986 0 FreeSans 2560 0 0 0 vssa2
port 558 nsew ground bidirectional
flabel metal5 s -8726 574366 592650 574986 0 FreeSans 2560 0 0 0 vssa2
port 558 nsew ground bidirectional
flabel metal5 s -8726 610366 592650 610986 0 FreeSans 2560 0 0 0 vssa2
port 558 nsew ground bidirectional
flabel metal5 s -8726 646366 592650 646986 0 FreeSans 2560 0 0 0 vssa2
port 558 nsew ground bidirectional
flabel metal5 s -8726 682366 592650 682986 0 FreeSans 2560 0 0 0 vssa2
port 558 nsew ground bidirectional
flabel metal4 s -2966 -1894 -2346 705830 0 FreeSans 3840 90 0 0 vssd1
port 559 nsew ground bidirectional
flabel metal5 s -2966 -1894 586890 -1274 0 FreeSans 2560 0 0 0 vssd1
port 559 nsew ground bidirectional
flabel metal5 s -2966 705210 586890 705830 0 FreeSans 2560 0 0 0 vssd1
port 559 nsew ground bidirectional
flabel metal4 s 586270 -1894 586890 705830 0 FreeSans 3840 90 0 0 vssd1
port 559 nsew ground bidirectional
flabel metal4 s 6294 -7654 6914 711590 0 FreeSans 3840 90 0 0 vssd1
port 559 nsew ground bidirectional
flabel metal4 s 42294 -7654 42914 711590 0 FreeSans 3840 90 0 0 vssd1
port 559 nsew ground bidirectional
flabel metal4 s 78294 -7654 78914 711590 0 FreeSans 3840 90 0 0 vssd1
port 559 nsew ground bidirectional
flabel metal4 s 114294 -7654 114914 711590 0 FreeSans 3840 90 0 0 vssd1
port 559 nsew ground bidirectional
flabel metal4 s 150294 -7654 150914 78000 0 FreeSans 3840 90 0 0 vssd1
port 559 nsew ground bidirectional
flabel metal4 s 150294 142000 150914 198000 0 FreeSans 3840 90 0 0 vssd1
port 559 nsew ground bidirectional
flabel metal4 s 150294 262000 150914 711590 0 FreeSans 3840 90 0 0 vssd1
port 559 nsew ground bidirectional
flabel metal4 s 186294 -7654 186914 78000 0 FreeSans 3840 90 0 0 vssd1
port 559 nsew ground bidirectional
flabel metal4 s 186294 142000 186914 198000 0 FreeSans 3840 90 0 0 vssd1
port 559 nsew ground bidirectional
flabel metal4 s 186294 262000 186914 711590 0 FreeSans 3840 90 0 0 vssd1
port 559 nsew ground bidirectional
flabel metal4 s 222294 -7654 222914 711590 0 FreeSans 3840 90 0 0 vssd1
port 559 nsew ground bidirectional
flabel metal4 s 258294 -7654 258914 711590 0 FreeSans 3840 90 0 0 vssd1
port 559 nsew ground bidirectional
flabel metal4 s 294294 -7654 294914 711590 0 FreeSans 3840 90 0 0 vssd1
port 559 nsew ground bidirectional
flabel metal4 s 330294 -7654 330914 711590 0 FreeSans 3840 90 0 0 vssd1
port 559 nsew ground bidirectional
flabel metal4 s 366294 -7654 366914 711590 0 FreeSans 3840 90 0 0 vssd1
port 559 nsew ground bidirectional
flabel metal4 s 402294 -7654 402914 711590 0 FreeSans 3840 90 0 0 vssd1
port 559 nsew ground bidirectional
flabel metal4 s 438294 -7654 438914 711590 0 FreeSans 3840 90 0 0 vssd1
port 559 nsew ground bidirectional
flabel metal4 s 474294 -7654 474914 711590 0 FreeSans 3840 90 0 0 vssd1
port 559 nsew ground bidirectional
flabel metal4 s 510294 -7654 510914 711590 0 FreeSans 3840 90 0 0 vssd1
port 559 nsew ground bidirectional
flabel metal4 s 546294 -7654 546914 711590 0 FreeSans 3840 90 0 0 vssd1
port 559 nsew ground bidirectional
flabel metal4 s 582294 -7654 582914 711590 0 FreeSans 3840 90 0 0 vssd1
port 559 nsew ground bidirectional
flabel metal5 s -8726 7366 592650 7986 0 FreeSans 2560 0 0 0 vssd1
port 559 nsew ground bidirectional
flabel metal5 s -8726 43366 592650 43986 0 FreeSans 2560 0 0 0 vssd1
port 559 nsew ground bidirectional
flabel metal5 s -8726 79366 592650 79986 0 FreeSans 2560 0 0 0 vssd1
port 559 nsew ground bidirectional
flabel metal5 s -8726 115366 592650 115986 0 FreeSans 2560 0 0 0 vssd1
port 559 nsew ground bidirectional
flabel metal5 s -8726 151366 592650 151986 0 FreeSans 2560 0 0 0 vssd1
port 559 nsew ground bidirectional
flabel metal5 s -8726 187366 592650 187986 0 FreeSans 2560 0 0 0 vssd1
port 559 nsew ground bidirectional
flabel metal5 s -8726 223366 592650 223986 0 FreeSans 2560 0 0 0 vssd1
port 559 nsew ground bidirectional
flabel metal5 s -8726 259366 592650 259986 0 FreeSans 2560 0 0 0 vssd1
port 559 nsew ground bidirectional
flabel metal5 s -8726 295366 592650 295986 0 FreeSans 2560 0 0 0 vssd1
port 559 nsew ground bidirectional
flabel metal5 s -8726 331366 592650 331986 0 FreeSans 2560 0 0 0 vssd1
port 559 nsew ground bidirectional
flabel metal5 s -8726 367366 592650 367986 0 FreeSans 2560 0 0 0 vssd1
port 559 nsew ground bidirectional
flabel metal5 s -8726 403366 592650 403986 0 FreeSans 2560 0 0 0 vssd1
port 559 nsew ground bidirectional
flabel metal5 s -8726 439366 592650 439986 0 FreeSans 2560 0 0 0 vssd1
port 559 nsew ground bidirectional
flabel metal5 s -8726 475366 592650 475986 0 FreeSans 2560 0 0 0 vssd1
port 559 nsew ground bidirectional
flabel metal5 s -8726 511366 592650 511986 0 FreeSans 2560 0 0 0 vssd1
port 559 nsew ground bidirectional
flabel metal5 s -8726 547366 592650 547986 0 FreeSans 2560 0 0 0 vssd1
port 559 nsew ground bidirectional
flabel metal5 s -8726 583366 592650 583986 0 FreeSans 2560 0 0 0 vssd1
port 559 nsew ground bidirectional
flabel metal5 s -8726 619366 592650 619986 0 FreeSans 2560 0 0 0 vssd1
port 559 nsew ground bidirectional
flabel metal5 s -8726 655366 592650 655986 0 FreeSans 2560 0 0 0 vssd1
port 559 nsew ground bidirectional
flabel metal5 s -8726 691366 592650 691986 0 FreeSans 2560 0 0 0 vssd1
port 559 nsew ground bidirectional
flabel metal4 s -4886 -3814 -4266 707750 0 FreeSans 3840 90 0 0 vssd2
port 560 nsew ground bidirectional
flabel metal5 s -4886 -3814 588810 -3194 0 FreeSans 2560 0 0 0 vssd2
port 560 nsew ground bidirectional
flabel metal5 s -4886 707130 588810 707750 0 FreeSans 2560 0 0 0 vssd2
port 560 nsew ground bidirectional
flabel metal4 s 588190 -3814 588810 707750 0 FreeSans 3840 90 0 0 vssd2
port 560 nsew ground bidirectional
flabel metal4 s 15294 -7654 15914 711590 0 FreeSans 3840 90 0 0 vssd2
port 560 nsew ground bidirectional
flabel metal4 s 51294 -7654 51914 711590 0 FreeSans 3840 90 0 0 vssd2
port 560 nsew ground bidirectional
flabel metal4 s 87294 -7654 87914 711590 0 FreeSans 3840 90 0 0 vssd2
port 560 nsew ground bidirectional
flabel metal4 s 123294 -7654 123914 78000 0 FreeSans 3840 90 0 0 vssd2
port 560 nsew ground bidirectional
flabel metal4 s 123294 142000 123914 198000 0 FreeSans 3840 90 0 0 vssd2
port 560 nsew ground bidirectional
flabel metal4 s 123294 262000 123914 711590 0 FreeSans 3840 90 0 0 vssd2
port 560 nsew ground bidirectional
flabel metal4 s 159294 -7654 159914 78000 0 FreeSans 3840 90 0 0 vssd2
port 560 nsew ground bidirectional
flabel metal4 s 159294 142000 159914 198000 0 FreeSans 3840 90 0 0 vssd2
port 560 nsew ground bidirectional
flabel metal4 s 159294 262000 159914 711590 0 FreeSans 3840 90 0 0 vssd2
port 560 nsew ground bidirectional
flabel metal4 s 195294 -7654 195914 711590 0 FreeSans 3840 90 0 0 vssd2
port 560 nsew ground bidirectional
flabel metal4 s 231294 -7654 231914 711590 0 FreeSans 3840 90 0 0 vssd2
port 560 nsew ground bidirectional
flabel metal4 s 267294 -7654 267914 711590 0 FreeSans 3840 90 0 0 vssd2
port 560 nsew ground bidirectional
flabel metal4 s 303294 -7654 303914 711590 0 FreeSans 3840 90 0 0 vssd2
port 560 nsew ground bidirectional
flabel metal4 s 339294 -7654 339914 711590 0 FreeSans 3840 90 0 0 vssd2
port 560 nsew ground bidirectional
flabel metal4 s 375294 -7654 375914 711590 0 FreeSans 3840 90 0 0 vssd2
port 560 nsew ground bidirectional
flabel metal4 s 411294 -7654 411914 711590 0 FreeSans 3840 90 0 0 vssd2
port 560 nsew ground bidirectional
flabel metal4 s 447294 -7654 447914 711590 0 FreeSans 3840 90 0 0 vssd2
port 560 nsew ground bidirectional
flabel metal4 s 483294 -7654 483914 711590 0 FreeSans 3840 90 0 0 vssd2
port 560 nsew ground bidirectional
flabel metal4 s 519294 -7654 519914 711590 0 FreeSans 3840 90 0 0 vssd2
port 560 nsew ground bidirectional
flabel metal4 s 555294 -7654 555914 711590 0 FreeSans 3840 90 0 0 vssd2
port 560 nsew ground bidirectional
flabel metal5 s -8726 16366 592650 16986 0 FreeSans 2560 0 0 0 vssd2
port 560 nsew ground bidirectional
flabel metal5 s -8726 52366 592650 52986 0 FreeSans 2560 0 0 0 vssd2
port 560 nsew ground bidirectional
flabel metal5 s -8726 88366 592650 88986 0 FreeSans 2560 0 0 0 vssd2
port 560 nsew ground bidirectional
flabel metal5 s -8726 124366 592650 124986 0 FreeSans 2560 0 0 0 vssd2
port 560 nsew ground bidirectional
flabel metal5 s -8726 160366 592650 160986 0 FreeSans 2560 0 0 0 vssd2
port 560 nsew ground bidirectional
flabel metal5 s -8726 196366 592650 196986 0 FreeSans 2560 0 0 0 vssd2
port 560 nsew ground bidirectional
flabel metal5 s -8726 232366 592650 232986 0 FreeSans 2560 0 0 0 vssd2
port 560 nsew ground bidirectional
flabel metal5 s -8726 268366 592650 268986 0 FreeSans 2560 0 0 0 vssd2
port 560 nsew ground bidirectional
flabel metal5 s -8726 304366 592650 304986 0 FreeSans 2560 0 0 0 vssd2
port 560 nsew ground bidirectional
flabel metal5 s -8726 340366 592650 340986 0 FreeSans 2560 0 0 0 vssd2
port 560 nsew ground bidirectional
flabel metal5 s -8726 376366 592650 376986 0 FreeSans 2560 0 0 0 vssd2
port 560 nsew ground bidirectional
flabel metal5 s -8726 412366 592650 412986 0 FreeSans 2560 0 0 0 vssd2
port 560 nsew ground bidirectional
flabel metal5 s -8726 448366 592650 448986 0 FreeSans 2560 0 0 0 vssd2
port 560 nsew ground bidirectional
flabel metal5 s -8726 484366 592650 484986 0 FreeSans 2560 0 0 0 vssd2
port 560 nsew ground bidirectional
flabel metal5 s -8726 520366 592650 520986 0 FreeSans 2560 0 0 0 vssd2
port 560 nsew ground bidirectional
flabel metal5 s -8726 556366 592650 556986 0 FreeSans 2560 0 0 0 vssd2
port 560 nsew ground bidirectional
flabel metal5 s -8726 592366 592650 592986 0 FreeSans 2560 0 0 0 vssd2
port 560 nsew ground bidirectional
flabel metal5 s -8726 628366 592650 628986 0 FreeSans 2560 0 0 0 vssd2
port 560 nsew ground bidirectional
flabel metal5 s -8726 664366 592650 664986 0 FreeSans 2560 0 0 0 vssd2
port 560 nsew ground bidirectional
flabel metal5 s -8726 700366 592650 700986 0 FreeSans 2560 0 0 0 vssd2
port 560 nsew ground bidirectional
flabel metal3 s 583520 256988 584960 257228 0 FreeSans 960 0 0 0 wb_clk_i
port 561 nsew signal input
flabel metal3 s -960 348788 480 349028 0 FreeSans 960 0 0 0 wb_rst_i
port 562 nsew signal input
flabel metal3 s 583520 385508 584960 385748 0 FreeSans 960 0 0 0 wbs_ack_o
port 563 nsew signal tristate
flabel metal2 s 198342 703520 198454 704960 0 FreeSans 448 90 0 0 wbs_adr_i[0]
port 564 nsew signal input
flabel metal2 s 54086 703520 54198 704960 0 FreeSans 448 90 0 0 wbs_adr_i[10]
port 565 nsew signal input
flabel metal3 s -960 472548 480 472788 0 FreeSans 960 0 0 0 wbs_adr_i[11]
port 566 nsew signal input
flabel metal2 s 64390 -960 64502 480 0 FreeSans 448 90 0 0 wbs_adr_i[12]
port 567 nsew signal input
flabel metal3 s -960 360348 480 360588 0 FreeSans 960 0 0 0 wbs_adr_i[13]
port 568 nsew signal input
flabel metal3 s 583520 662268 584960 662508 0 FreeSans 960 0 0 0 wbs_adr_i[14]
port 569 nsew signal input
flabel metal3 s 583520 613988 584960 614228 0 FreeSans 960 0 0 0 wbs_adr_i[15]
port 570 nsew signal input
flabel metal2 s 443706 -960 443818 480 0 FreeSans 448 90 0 0 wbs_adr_i[16]
port 571 nsew signal input
flabel metal3 s 583520 557548 584960 557788 0 FreeSans 960 0 0 0 wbs_adr_i[17]
port 572 nsew signal input
flabel metal3 s 583520 345388 584960 345628 0 FreeSans 960 0 0 0 wbs_adr_i[18]
port 573 nsew signal input
flabel metal3 s 583520 88348 584960 88588 0 FreeSans 960 0 0 0 wbs_adr_i[19]
port 574 nsew signal input
flabel metal2 s 206070 703520 206182 704960 0 FreeSans 448 90 0 0 wbs_adr_i[1]
port 575 nsew signal input
flabel metal2 s 406998 703520 407110 704960 0 FreeSans 448 90 0 0 wbs_adr_i[20]
port 576 nsew signal input
flabel metal2 s 390898 -960 391010 480 0 FreeSans 448 90 0 0 wbs_adr_i[21]
port 577 nsew signal input
flabel metal2 s 557694 -960 557806 480 0 FreeSans 448 90 0 0 wbs_adr_i[22]
port 578 nsew signal input
flabel metal3 s 583520 276708 584960 276948 0 FreeSans 960 0 0 0 wbs_adr_i[23]
port 579 nsew signal input
flabel metal3 s -960 552788 480 553028 0 FreeSans 960 0 0 0 wbs_adr_i[24]
port 580 nsew signal input
flabel metal2 s 375442 -960 375554 480 0 FreeSans 448 90 0 0 wbs_adr_i[25]
port 581 nsew signal input
flabel metal2 s 72118 -960 72230 480 0 FreeSans 448 90 0 0 wbs_adr_i[26]
port 582 nsew signal input
flabel metal3 s -960 19668 480 19908 0 FreeSans 960 0 0 0 wbs_adr_i[27]
port 583 nsew signal input
flabel metal3 s 583520 525588 584960 525828 0 FreeSans 960 0 0 0 wbs_adr_i[28]
port 584 nsew signal input
flabel metal2 s 498446 703520 498558 704960 0 FreeSans 448 90 0 0 wbs_adr_i[29]
port 585 nsew signal input
flabel metal2 s 265318 -960 265430 480 0 FreeSans 448 90 0 0 wbs_adr_i[2]
port 586 nsew signal input
flabel metal2 s 331006 703520 331118 704960 0 FreeSans 448 90 0 0 wbs_adr_i[30]
port 587 nsew signal input
flabel metal3 s 583520 405228 584960 405468 0 FreeSans 960 0 0 0 wbs_adr_i[31]
port 588 nsew signal input
flabel metal2 s 531290 -960 531402 480 0 FreeSans 448 90 0 0 wbs_adr_i[3]
port 589 nsew signal input
flabel metal2 s 323922 703520 324034 704960 0 FreeSans 448 90 0 0 wbs_adr_i[4]
port 590 nsew signal input
flabel metal3 s -960 108068 480 108308 0 FreeSans 960 0 0 0 wbs_adr_i[5]
port 591 nsew signal input
flabel metal2 s 216374 -960 216486 480 0 FreeSans 448 90 0 0 wbs_adr_i[6]
port 592 nsew signal input
flabel metal2 s 34122 -960 34234 480 0 FreeSans 448 90 0 0 wbs_adr_i[7]
port 593 nsew signal input
flabel metal3 s 583520 96508 584960 96748 0 FreeSans 960 0 0 0 wbs_adr_i[8]
port 594 nsew signal input
flabel metal3 s 583520 288948 584960 289188 0 FreeSans 960 0 0 0 wbs_adr_i[9]
port 595 nsew signal input
flabel metal2 s 27682 703520 27794 704960 0 FreeSans 448 90 0 0 wbs_cyc_i
port 596 nsew signal input
flabel metal2 s 574438 703520 574550 704960 0 FreeSans 448 90 0 0 wbs_dat_i[0]
port 597 nsew signal input
flabel metal3 s -960 356268 480 356508 0 FreeSans 960 0 0 0 wbs_dat_i[10]
port 598 nsew signal input
flabel metal3 s -960 408628 480 408868 0 FreeSans 960 0 0 0 wbs_dat_i[11]
port 599 nsew signal input
flabel metal3 s -960 388228 480 388468 0 FreeSans 960 0 0 0 wbs_dat_i[12]
port 600 nsew signal input
flabel metal2 s 26394 -960 26506 480 0 FreeSans 448 90 0 0 wbs_dat_i[13]
port 601 nsew signal input
flabel metal2 s 144246 -960 144358 480 0 FreeSans 448 90 0 0 wbs_dat_i[14]
port 602 nsew signal input
flabel metal3 s 583520 457588 584960 457828 0 FreeSans 960 0 0 0 wbs_dat_i[15]
port 603 nsew signal input
flabel metal3 s -960 43468 480 43708 0 FreeSans 960 0 0 0 wbs_dat_i[16]
port 604 nsew signal input
flabel metal2 s 293010 703520 293122 704960 0 FreeSans 448 90 0 0 wbs_dat_i[17]
port 605 nsew signal input
flabel metal2 s 456586 703520 456698 704960 0 FreeSans 448 90 0 0 wbs_dat_i[18]
port 606 nsew signal input
flabel metal3 s -960 577268 480 577508 0 FreeSans 960 0 0 0 wbs_dat_i[19]
port 607 nsew signal input
flabel metal2 s 102386 -960 102498 480 0 FreeSans 448 90 0 0 wbs_dat_i[1]
port 608 nsew signal input
flabel metal3 s 583520 505868 584960 506108 0 FreeSans 960 0 0 0 wbs_dat_i[20]
port 609 nsew signal input
flabel metal2 s 479126 703520 479238 704960 0 FreeSans 448 90 0 0 wbs_dat_i[21]
port 610 nsew signal input
flabel metal3 s -960 264468 480 264708 0 FreeSans 960 0 0 0 wbs_dat_i[22]
port 611 nsew signal input
flabel metal3 s 583520 629628 584960 629868 0 FreeSans 960 0 0 0 wbs_dat_i[23]
port 612 nsew signal input
flabel metal3 s 583520 309348 584960 309588 0 FreeSans 960 0 0 0 wbs_dat_i[24]
port 613 nsew signal input
flabel metal2 s 459162 -960 459274 480 0 FreeSans 448 90 0 0 wbs_dat_i[25]
port 614 nsew signal input
flabel metal2 s 410862 703520 410974 704960 0 FreeSans 448 90 0 0 wbs_dat_i[26]
port 615 nsew signal input
flabel metal2 s 19954 703520 20066 704960 0 FreeSans 448 90 0 0 wbs_dat_i[27]
port 616 nsew signal input
flabel metal2 s 208646 -960 208758 480 0 FreeSans 448 90 0 0 wbs_dat_i[28]
port 617 nsew signal input
flabel metal3 s 583520 497708 584960 497948 0 FreeSans 960 0 0 0 wbs_dat_i[29]
port 618 nsew signal input
flabel metal2 s 539018 -960 539130 480 0 FreeSans 448 90 0 0 wbs_dat_i[2]
port 619 nsew signal input
flabel metal3 s 583520 280788 584960 281028 0 FreeSans 960 0 0 0 wbs_dat_i[30]
port 620 nsew signal input
flabel metal3 s -960 248148 480 248388 0 FreeSans 960 0 0 0 wbs_dat_i[31]
port 621 nsew signal input
flabel metal3 s 583520 100588 584960 100828 0 FreeSans 960 0 0 0 wbs_dat_i[3]
port 622 nsew signal input
flabel metal2 s 106250 -960 106362 480 0 FreeSans 448 90 0 0 wbs_dat_i[4]
port 623 nsew signal input
flabel metal2 s 326498 -960 326610 480 0 FreeSans 448 90 0 0 wbs_dat_i[5]
port 624 nsew signal input
flabel metal3 s 583520 373268 584960 373508 0 FreeSans 960 0 0 0 wbs_dat_i[6]
port 625 nsew signal input
flabel metal2 s 399914 703520 400026 704960 0 FreeSans 448 90 0 0 wbs_dat_i[7]
port 626 nsew signal input
flabel metal3 s 583520 686068 584960 686308 0 FreeSans 960 0 0 0 wbs_dat_i[8]
port 627 nsew signal input
flabel metal3 s 583520 104668 584960 104908 0 FreeSans 960 0 0 0 wbs_dat_i[9]
port 628 nsew signal input
flabel metal2 s 52798 -960 52910 480 0 FreeSans 448 90 0 0 wbs_dat_o[0]
port 629 nsew signal tristate
flabel metal3 s 583520 461668 584960 461908 0 FreeSans 960 0 0 0 wbs_dat_o[10]
port 630 nsew signal tristate
flabel metal2 s 14802 -960 14914 480 0 FreeSans 448 90 0 0 wbs_dat_o[11]
port 631 nsew signal tristate
flabel metal3 s 583520 694228 584960 694468 0 FreeSans 960 0 0 0 wbs_dat_o[12]
port 632 nsew signal tristate
flabel metal2 s 384458 703520 384570 704960 0 FreeSans 448 90 0 0 wbs_dat_o[13]
port 633 nsew signal tristate
flabel metal3 s 583520 144788 584960 145028 0 FreeSans 960 0 0 0 wbs_dat_o[14]
port 634 nsew signal tristate
flabel metal2 s 365138 703520 365250 704960 0 FreeSans 448 90 0 0 wbs_dat_o[15]
port 635 nsew signal tristate
flabel metal2 s 436622 -960 436734 480 0 FreeSans 448 90 0 0 wbs_dat_o[16]
port 636 nsew signal tristate
flabel metal3 s -960 135948 480 136188 0 FreeSans 960 0 0 0 wbs_dat_o[17]
port 637 nsew signal tristate
flabel metal2 s 432758 -960 432870 480 0 FreeSans 448 90 0 0 wbs_dat_o[18]
port 638 nsew signal tristate
flabel metal2 s -10 -960 102 480 0 FreeSans 448 90 0 0 wbs_dat_o[19]
port 639 nsew signal tristate
flabel metal2 s 508750 -960 508862 480 0 FreeSans 448 90 0 0 wbs_dat_o[1]
port 640 nsew signal tristate
flabel metal3 s -960 256308 480 256548 0 FreeSans 960 0 0 0 wbs_dat_o[20]
port 641 nsew signal tristate
flabel metal3 s -960 524908 480 525148 0 FreeSans 960 0 0 0 wbs_dat_o[21]
port 642 nsew signal tristate
flabel metal2 s 92082 703520 92194 704960 0 FreeSans 448 90 0 0 wbs_dat_o[22]
port 643 nsew signal tristate
flabel metal3 s -960 167908 480 168148 0 FreeSans 960 0 0 0 wbs_dat_o[23]
port 644 nsew signal tristate
flabel metal2 s 132654 -960 132766 480 0 FreeSans 448 90 0 0 wbs_dat_o[24]
port 645 nsew signal tristate
flabel metal2 s 48934 -960 49046 480 0 FreeSans 448 90 0 0 wbs_dat_o[25]
port 646 nsew signal tristate
flabel metal2 s 255014 703520 255126 704960 0 FreeSans 448 90 0 0 wbs_dat_o[26]
port 647 nsew signal tristate
flabel metal2 s 114622 703520 114734 704960 0 FreeSans 448 90 0 0 wbs_dat_o[27]
port 648 nsew signal tristate
flabel metal2 s 345174 -960 345286 480 0 FreeSans 448 90 0 0 wbs_dat_o[28]
port 649 nsew signal tristate
flabel metal2 s 369002 703520 369114 704960 0 FreeSans 448 90 0 0 wbs_dat_o[29]
port 650 nsew signal tristate
flabel metal3 s 583520 240668 584960 240908 0 FreeSans 960 0 0 0 wbs_dat_o[2]
port 651 nsew signal tristate
flabel metal3 s -960 404548 480 404788 0 FreeSans 960 0 0 0 wbs_dat_o[30]
port 652 nsew signal tristate
flabel metal3 s 583520 569788 584960 570028 0 FreeSans 960 0 0 0 wbs_dat_o[31]
port 653 nsew signal tristate
flabel metal2 s 140382 -960 140494 480 0 FreeSans 448 90 0 0 wbs_dat_o[3]
port 654 nsew signal tristate
flabel metal2 s 242778 -960 242890 480 0 FreeSans 448 90 0 0 wbs_dat_o[4]
port 655 nsew signal tristate
flabel metal3 s -960 35988 480 36228 0 FreeSans 960 0 0 0 wbs_dat_o[5]
port 656 nsew signal tristate
flabel metal3 s 583520 541908 584960 542148 0 FreeSans 960 0 0 0 wbs_dat_o[6]
port 657 nsew signal tristate
flabel metal2 s 383170 -960 383282 480 0 FreeSans 448 90 0 0 wbs_dat_o[7]
port 658 nsew signal tristate
flabel metal2 s 358054 703520 358166 704960 0 FreeSans 448 90 0 0 wbs_dat_o[8]
port 659 nsew signal tristate
flabel metal2 s 354190 703520 354302 704960 0 FreeSans 448 90 0 0 wbs_dat_o[9]
port 660 nsew signal tristate
flabel metal3 s -960 601068 480 601308 0 FreeSans 960 0 0 0 wbs_sel_i[0]
port 661 nsew signal input
flabel metal2 s 16090 703520 16202 704960 0 FreeSans 448 90 0 0 wbs_sel_i[1]
port 662 nsew signal input
flabel metal2 s 455298 -960 455410 480 0 FreeSans 448 90 0 0 wbs_sel_i[2]
port 663 nsew signal input
flabel metal3 s -960 140028 480 140268 0 FreeSans 960 0 0 0 wbs_sel_i[3]
port 664 nsew signal input
flabel metal3 s -960 541228 480 541468 0 FreeSans 960 0 0 0 wbs_stb_i
port 665 nsew signal input
flabel metal3 s 583520 369188 584960 369428 0 FreeSans 960 0 0 0 wbs_we_i
port 666 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
